module basic_1000_10000_1500_10_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
xor U0 (N_0,In_739,In_948);
or U1 (N_1,In_509,In_589);
xnor U2 (N_2,In_639,In_823);
nor U3 (N_3,In_136,In_374);
xor U4 (N_4,In_531,In_395);
nor U5 (N_5,In_381,In_463);
and U6 (N_6,In_790,In_280);
or U7 (N_7,In_508,In_425);
nor U8 (N_8,In_500,In_227);
nand U9 (N_9,In_84,In_837);
xnor U10 (N_10,In_816,In_539);
xnor U11 (N_11,In_82,In_518);
xnor U12 (N_12,In_747,In_601);
nor U13 (N_13,In_950,In_768);
and U14 (N_14,In_669,In_77);
and U15 (N_15,In_255,In_822);
and U16 (N_16,In_880,In_346);
or U17 (N_17,In_157,In_792);
nand U18 (N_18,In_831,In_715);
nand U19 (N_19,In_905,In_414);
or U20 (N_20,In_783,In_545);
nor U21 (N_21,In_930,In_896);
or U22 (N_22,In_422,In_460);
nor U23 (N_23,In_844,In_690);
and U24 (N_24,In_989,In_288);
nor U25 (N_25,In_985,In_379);
xnor U26 (N_26,In_376,In_356);
or U27 (N_27,In_329,In_714);
and U28 (N_28,In_826,In_406);
or U29 (N_29,In_477,In_103);
nor U30 (N_30,In_26,In_527);
nand U31 (N_31,In_201,In_483);
or U32 (N_32,In_176,In_951);
or U33 (N_33,In_204,In_179);
xor U34 (N_34,In_563,In_383);
or U35 (N_35,In_752,In_11);
xor U36 (N_36,In_361,In_565);
and U37 (N_37,In_494,In_555);
nor U38 (N_38,In_40,In_855);
nand U39 (N_39,In_322,In_606);
and U40 (N_40,In_232,In_184);
nor U41 (N_41,In_264,In_666);
or U42 (N_42,In_964,In_932);
and U43 (N_43,In_338,In_403);
and U44 (N_44,In_526,In_110);
nand U45 (N_45,In_180,In_570);
or U46 (N_46,In_436,In_484);
and U47 (N_47,In_706,In_686);
nor U48 (N_48,In_482,In_640);
nor U49 (N_49,In_972,In_617);
nand U50 (N_50,In_865,In_623);
nand U51 (N_51,In_317,In_170);
nand U52 (N_52,In_7,In_210);
nor U53 (N_53,In_521,In_523);
and U54 (N_54,In_620,In_677);
nor U55 (N_55,In_126,In_995);
or U56 (N_56,In_140,In_707);
and U57 (N_57,In_24,In_743);
nor U58 (N_58,In_870,In_767);
nand U59 (N_59,In_986,In_828);
xor U60 (N_60,In_638,In_278);
and U61 (N_61,In_169,In_108);
nand U62 (N_62,In_630,In_18);
and U63 (N_63,In_943,In_242);
or U64 (N_64,In_773,In_475);
and U65 (N_65,In_207,In_37);
nor U66 (N_66,In_664,In_654);
or U67 (N_67,In_259,In_327);
or U68 (N_68,In_561,In_392);
and U69 (N_69,In_366,In_732);
and U70 (N_70,In_618,In_44);
nor U71 (N_71,In_312,In_745);
or U72 (N_72,In_716,In_344);
and U73 (N_73,In_293,In_340);
and U74 (N_74,In_770,In_848);
nand U75 (N_75,In_914,In_421);
nor U76 (N_76,In_78,In_240);
nor U77 (N_77,In_710,In_927);
or U78 (N_78,In_852,In_996);
xnor U79 (N_79,In_221,In_281);
xnor U80 (N_80,In_698,In_871);
xnor U81 (N_81,In_876,In_471);
nor U82 (N_82,In_467,In_54);
or U83 (N_83,In_622,In_564);
nand U84 (N_84,In_260,In_820);
and U85 (N_85,In_897,In_637);
xnor U86 (N_86,In_921,In_980);
nand U87 (N_87,In_287,In_998);
or U88 (N_88,In_696,In_94);
xnor U89 (N_89,In_311,In_16);
nor U90 (N_90,In_34,In_187);
xor U91 (N_91,In_434,In_629);
nor U92 (N_92,In_520,In_911);
xnor U93 (N_93,In_85,In_578);
nor U94 (N_94,In_970,In_528);
nand U95 (N_95,In_397,In_223);
nor U96 (N_96,In_411,In_358);
nor U97 (N_97,In_203,In_616);
and U98 (N_98,In_459,In_772);
and U99 (N_99,In_378,In_119);
and U100 (N_100,In_847,In_805);
and U101 (N_101,In_653,In_277);
nand U102 (N_102,In_367,In_824);
xnor U103 (N_103,In_702,In_314);
xor U104 (N_104,In_821,In_689);
xnor U105 (N_105,In_462,In_993);
and U106 (N_106,In_802,In_513);
nor U107 (N_107,In_579,In_257);
nand U108 (N_108,In_442,In_940);
and U109 (N_109,In_333,In_365);
xnor U110 (N_110,In_98,In_472);
xor U111 (N_111,In_735,In_107);
and U112 (N_112,In_440,In_857);
and U113 (N_113,In_685,In_969);
or U114 (N_114,In_214,In_355);
nor U115 (N_115,In_130,In_38);
and U116 (N_116,In_2,In_835);
nand U117 (N_117,In_321,In_572);
nand U118 (N_118,In_318,In_755);
and U119 (N_119,In_145,In_446);
nor U120 (N_120,In_774,In_49);
and U121 (N_121,In_731,In_953);
xnor U122 (N_122,In_580,In_784);
and U123 (N_123,In_218,In_448);
nand U124 (N_124,In_704,In_650);
or U125 (N_125,In_678,In_647);
nor U126 (N_126,In_62,In_430);
xnor U127 (N_127,In_974,In_920);
xor U128 (N_128,In_938,In_246);
nor U129 (N_129,In_213,In_765);
and U130 (N_130,In_568,In_152);
nor U131 (N_131,In_363,In_717);
nand U132 (N_132,In_931,In_503);
and U133 (N_133,In_804,In_88);
nor U134 (N_134,In_237,In_348);
or U135 (N_135,In_112,In_939);
xnor U136 (N_136,In_359,In_890);
nor U137 (N_137,In_819,In_688);
xor U138 (N_138,In_27,In_636);
nand U139 (N_139,In_189,In_727);
nand U140 (N_140,In_275,In_517);
and U141 (N_141,In_8,In_141);
nor U142 (N_142,In_615,In_611);
or U143 (N_143,In_86,In_682);
and U144 (N_144,In_901,In_25);
or U145 (N_145,In_510,In_265);
nor U146 (N_146,In_632,In_76);
xnor U147 (N_147,In_247,In_841);
nand U148 (N_148,In_429,In_538);
and U149 (N_149,In_658,In_282);
and U150 (N_150,In_14,In_352);
nor U151 (N_151,In_134,In_560);
nand U152 (N_152,In_933,In_780);
nand U153 (N_153,In_874,In_858);
xnor U154 (N_154,In_592,In_584);
nand U155 (N_155,In_43,In_760);
nor U156 (N_156,In_224,In_971);
and U157 (N_157,In_753,In_505);
xnor U158 (N_158,In_935,In_299);
nand U159 (N_159,In_612,In_489);
xnor U160 (N_160,In_591,In_51);
and U161 (N_161,In_104,In_36);
and U162 (N_162,In_233,In_769);
nand U163 (N_163,In_441,In_977);
nand U164 (N_164,In_574,In_91);
and U165 (N_165,In_480,In_127);
or U166 (N_166,In_663,In_6);
or U167 (N_167,In_501,In_334);
nor U168 (N_168,In_377,In_725);
nor U169 (N_169,In_909,In_32);
or U170 (N_170,In_241,In_335);
xor U171 (N_171,In_419,In_569);
and U172 (N_172,In_577,In_889);
and U173 (N_173,In_486,In_323);
nor U174 (N_174,In_786,In_634);
xnor U175 (N_175,In_324,In_478);
or U176 (N_176,In_499,In_468);
xnor U177 (N_177,In_785,In_173);
nand U178 (N_178,In_893,In_854);
nor U179 (N_179,In_779,In_956);
and U180 (N_180,In_39,In_600);
xor U181 (N_181,In_409,In_426);
or U182 (N_182,In_93,In_45);
xnor U183 (N_183,In_267,In_407);
or U184 (N_184,In_469,In_391);
nor U185 (N_185,In_530,In_557);
xnor U186 (N_186,In_982,In_33);
nor U187 (N_187,In_192,In_962);
nor U188 (N_188,In_481,In_608);
or U189 (N_189,In_882,In_149);
nand U190 (N_190,In_56,In_438);
and U191 (N_191,In_215,In_229);
nor U192 (N_192,In_125,In_929);
nand U193 (N_193,In_326,In_163);
nand U194 (N_194,In_23,In_479);
and U195 (N_195,In_867,In_793);
nor U196 (N_196,In_641,In_61);
xor U197 (N_197,In_684,In_511);
nand U198 (N_198,In_236,In_310);
nor U199 (N_199,In_28,In_162);
and U200 (N_200,In_129,In_394);
or U201 (N_201,In_263,In_271);
and U202 (N_202,In_963,In_303);
xor U203 (N_203,In_79,In_583);
nor U204 (N_204,In_270,In_529);
xor U205 (N_205,In_144,In_156);
nand U206 (N_206,In_946,In_535);
xor U207 (N_207,In_354,In_55);
xnor U208 (N_208,In_808,In_458);
nor U209 (N_209,In_945,In_47);
nand U210 (N_210,In_797,In_525);
nand U211 (N_211,In_674,In_595);
or U212 (N_212,In_633,In_991);
xnor U213 (N_213,In_984,In_840);
xor U214 (N_214,In_553,In_681);
and U215 (N_215,In_402,In_665);
nand U216 (N_216,In_659,In_506);
xnor U217 (N_217,In_728,In_566);
or U218 (N_218,In_700,In_197);
xnor U219 (N_219,In_50,In_74);
or U220 (N_220,In_3,In_485);
xor U221 (N_221,In_105,In_846);
xor U222 (N_222,In_185,In_514);
nor U223 (N_223,In_385,In_465);
nand U224 (N_224,In_992,In_164);
nand U225 (N_225,In_798,In_279);
nor U226 (N_226,In_268,In_498);
and U227 (N_227,In_853,In_541);
or U228 (N_228,In_596,In_843);
or U229 (N_229,In_777,In_139);
nand U230 (N_230,In_336,In_872);
nor U231 (N_231,In_69,In_80);
and U232 (N_232,In_290,In_540);
and U233 (N_233,In_137,In_524);
nand U234 (N_234,In_249,In_357);
and U235 (N_235,In_216,In_372);
nand U236 (N_236,In_220,In_234);
and U237 (N_237,In_894,In_48);
nand U238 (N_238,In_646,In_175);
xnor U239 (N_239,In_347,In_199);
nor U240 (N_240,In_362,In_627);
and U241 (N_241,In_159,In_315);
xor U242 (N_242,In_742,In_349);
xnor U243 (N_243,In_474,In_122);
and U244 (N_244,In_807,In_937);
and U245 (N_245,In_602,In_766);
xnor U246 (N_246,In_158,In_476);
nor U247 (N_247,In_544,In_941);
or U248 (N_248,In_67,In_427);
nor U249 (N_249,In_151,In_609);
and U250 (N_250,In_150,In_328);
nand U251 (N_251,In_918,In_965);
xor U252 (N_252,In_660,In_58);
nand U253 (N_253,In_21,In_902);
nor U254 (N_254,In_243,In_762);
nor U255 (N_255,In_624,In_202);
nor U256 (N_256,In_729,In_887);
nand U257 (N_257,In_92,In_331);
and U258 (N_258,In_269,In_694);
or U259 (N_259,In_863,In_188);
nand U260 (N_260,In_917,In_813);
nor U261 (N_261,In_764,In_680);
nor U262 (N_262,In_888,In_435);
and U263 (N_263,In_925,In_457);
nand U264 (N_264,In_389,In_17);
nor U265 (N_265,In_720,In_4);
nand U266 (N_266,In_955,In_988);
nand U267 (N_267,In_443,In_934);
or U268 (N_268,In_451,In_373);
nor U269 (N_269,In_226,In_292);
and U270 (N_270,In_597,In_235);
or U271 (N_271,In_748,In_492);
xor U272 (N_272,In_450,In_206);
nor U273 (N_273,In_285,In_502);
or U274 (N_274,In_364,In_416);
xor U275 (N_275,In_593,In_380);
nor U276 (N_276,In_59,In_668);
nand U277 (N_277,In_238,In_810);
nor U278 (N_278,In_705,In_360);
xor U279 (N_279,In_881,In_339);
nand U280 (N_280,In_947,In_75);
xnor U281 (N_281,In_212,In_211);
or U282 (N_282,In_532,In_744);
nor U283 (N_283,In_90,In_488);
xor U284 (N_284,In_398,In_771);
xor U285 (N_285,In_926,In_320);
or U286 (N_286,In_178,In_168);
nor U287 (N_287,In_598,In_730);
nand U288 (N_288,In_983,In_300);
nand U289 (N_289,In_936,In_519);
or U290 (N_290,In_63,In_657);
and U291 (N_291,In_154,In_504);
nand U292 (N_292,In_316,In_22);
and U293 (N_293,In_120,In_718);
or U294 (N_294,In_95,In_284);
nor U295 (N_295,In_309,In_547);
nand U296 (N_296,In_899,In_116);
and U297 (N_297,In_607,In_801);
nand U298 (N_298,In_928,In_691);
and U299 (N_299,In_845,In_332);
nor U300 (N_300,In_644,In_832);
nand U301 (N_301,In_849,In_57);
xor U302 (N_302,In_558,In_910);
xnor U303 (N_303,In_473,In_721);
or U304 (N_304,In_461,In_737);
xor U305 (N_305,In_573,In_800);
and U306 (N_306,In_746,In_975);
nand U307 (N_307,In_811,In_814);
xor U308 (N_308,In_976,In_997);
nand U309 (N_309,In_209,In_679);
nand U310 (N_310,In_759,In_952);
nor U311 (N_311,In_253,In_341);
nor U312 (N_312,In_493,In_628);
nor U313 (N_313,In_809,In_160);
or U314 (N_314,In_225,In_369);
nor U315 (N_315,In_10,In_827);
and U316 (N_316,In_726,In_262);
xor U317 (N_317,In_70,In_750);
or U318 (N_318,In_439,In_83);
nor U319 (N_319,In_683,In_671);
xnor U320 (N_320,In_307,In_432);
nor U321 (N_321,In_133,In_643);
or U322 (N_322,In_325,In_799);
xor U323 (N_323,In_304,In_878);
nand U324 (N_324,In_464,In_456);
or U325 (N_325,In_884,In_146);
nand U326 (N_326,In_46,In_635);
nor U327 (N_327,In_433,In_868);
nor U328 (N_328,In_960,In_205);
or U329 (N_329,In_834,In_537);
nand U330 (N_330,In_286,In_839);
and U331 (N_331,In_196,In_994);
or U332 (N_332,In_548,In_713);
and U333 (N_333,In_588,In_516);
or U334 (N_334,In_859,In_836);
nor U335 (N_335,In_128,In_533);
nand U336 (N_336,In_758,In_672);
nand U337 (N_337,In_812,In_455);
and U338 (N_338,In_576,In_289);
xnor U339 (N_339,In_231,In_195);
nand U340 (N_340,In_453,In_496);
nor U341 (N_341,In_631,In_490);
xor U342 (N_342,In_71,In_697);
or U343 (N_343,In_507,In_794);
and U344 (N_344,In_452,In_174);
xor U345 (N_345,In_515,In_454);
nor U346 (N_346,In_551,In_605);
and U347 (N_347,In_424,In_582);
nor U348 (N_348,In_171,In_661);
and U349 (N_349,In_850,In_979);
xor U350 (N_350,In_191,In_924);
or U351 (N_351,In_961,In_571);
or U352 (N_352,In_20,In_754);
nand U353 (N_353,In_9,In_15);
nor U354 (N_354,In_838,In_625);
and U355 (N_355,In_101,In_53);
or U356 (N_356,In_856,In_763);
nor U357 (N_357,In_873,In_692);
and U358 (N_358,In_19,In_554);
xor U359 (N_359,In_703,In_610);
nand U360 (N_360,In_399,In_353);
nand U361 (N_361,In_295,In_676);
xnor U362 (N_362,In_1,In_556);
or U363 (N_363,In_131,In_123);
nor U364 (N_364,In_981,In_308);
nand U365 (N_365,In_147,In_675);
and U366 (N_366,In_100,In_445);
nand U367 (N_367,In_603,In_586);
nor U368 (N_368,In_384,In_907);
or U369 (N_369,In_776,In_959);
nor U370 (N_370,In_172,In_673);
and U371 (N_371,In_791,In_978);
nor U372 (N_372,In_875,In_183);
or U373 (N_373,In_740,In_904);
nor U374 (N_374,In_388,In_670);
nand U375 (N_375,In_536,In_413);
and U376 (N_376,In_301,In_73);
xnor U377 (N_377,In_906,In_842);
nor U378 (N_378,In_655,In_552);
nand U379 (N_379,In_562,In_248);
or U380 (N_380,In_306,In_386);
nor U381 (N_381,In_41,In_512);
or U382 (N_382,In_417,In_250);
nor U383 (N_383,In_818,In_781);
nor U384 (N_384,In_782,In_298);
or U385 (N_385,In_115,In_118);
or U386 (N_386,In_102,In_420);
and U387 (N_387,In_567,In_177);
xnor U388 (N_388,In_751,In_651);
nand U389 (N_389,In_114,In_166);
and U390 (N_390,In_829,In_599);
and U391 (N_391,In_256,In_351);
and U392 (N_392,In_182,In_230);
nor U393 (N_393,In_866,In_757);
nor U394 (N_394,In_738,In_418);
xor U395 (N_395,In_594,In_276);
and U396 (N_396,In_550,In_198);
or U397 (N_397,In_109,In_415);
and U398 (N_398,In_313,In_319);
xor U399 (N_399,In_87,In_266);
xor U400 (N_400,In_968,In_879);
xnor U401 (N_401,In_862,In_778);
or U402 (N_402,In_795,In_656);
nor U403 (N_403,In_330,In_96);
nor U404 (N_404,In_957,In_13);
nor U405 (N_405,In_851,In_942);
and U406 (N_406,In_973,In_0);
or U407 (N_407,In_423,In_228);
xnor U408 (N_408,In_143,In_35);
nand U409 (N_409,In_111,In_65);
nand U410 (N_410,In_200,In_396);
xnor U411 (N_411,In_89,In_272);
and U412 (N_412,In_117,In_66);
nand U413 (N_413,In_756,In_546);
nor U414 (N_414,In_549,In_788);
and U415 (N_415,In_258,In_337);
nand U416 (N_416,In_590,In_273);
or U417 (N_417,In_194,In_291);
nor U418 (N_418,In_861,In_302);
xor U419 (N_419,In_701,In_648);
nand U420 (N_420,In_585,In_581);
and U421 (N_421,In_254,In_619);
nand U422 (N_422,In_741,In_186);
nand U423 (N_423,In_428,In_761);
or U424 (N_424,In_437,In_886);
nor U425 (N_425,In_891,In_400);
or U426 (N_426,In_587,In_401);
nand U427 (N_427,In_830,In_345);
and U428 (N_428,In_404,In_239);
nor U429 (N_429,In_903,In_900);
and U430 (N_430,In_495,In_52);
nand U431 (N_431,In_155,In_297);
nor U432 (N_432,In_375,In_864);
xor U433 (N_433,In_967,In_825);
xor U434 (N_434,In_723,In_898);
xor U435 (N_435,In_387,In_135);
nor U436 (N_436,In_722,In_719);
nor U437 (N_437,In_966,In_165);
xor U438 (N_438,In_412,In_491);
nand U439 (N_439,In_775,In_350);
nand U440 (N_440,In_817,In_405);
and U441 (N_441,In_113,In_121);
and U442 (N_442,In_294,In_181);
and U443 (N_443,In_787,In_885);
xor U444 (N_444,In_542,In_543);
nor U445 (N_445,In_693,In_408);
and U446 (N_446,In_190,In_711);
xor U447 (N_447,In_487,In_649);
and U448 (N_448,In_613,In_883);
nor U449 (N_449,In_916,In_106);
and U450 (N_450,In_42,In_915);
nor U451 (N_451,In_64,In_833);
nor U452 (N_452,In_958,In_662);
xor U453 (N_453,In_245,In_371);
xnor U454 (N_454,In_534,In_138);
nand U455 (N_455,In_447,In_990);
nand U456 (N_456,In_81,In_733);
nand U457 (N_457,In_431,In_217);
nor U458 (N_458,In_695,In_734);
and U459 (N_459,In_497,In_604);
xnor U460 (N_460,In_370,In_343);
xor U461 (N_461,In_390,In_193);
nand U462 (N_462,In_575,In_148);
nand U463 (N_463,In_559,In_382);
or U464 (N_464,In_803,In_30);
nand U465 (N_465,In_99,In_410);
nand U466 (N_466,In_869,In_97);
nor U467 (N_467,In_877,In_652);
nor U468 (N_468,In_614,In_470);
or U469 (N_469,In_949,In_153);
nand U470 (N_470,In_923,In_274);
nand U471 (N_471,In_305,In_796);
nor U472 (N_472,In_124,In_208);
and U473 (N_473,In_444,In_283);
and U474 (N_474,In_466,In_222);
nor U475 (N_475,In_72,In_642);
xnor U476 (N_476,In_987,In_522);
and U477 (N_477,In_29,In_132);
nand U478 (N_478,In_944,In_709);
xnor U479 (N_479,In_687,In_699);
nor U480 (N_480,In_68,In_749);
nand U481 (N_481,In_449,In_922);
or U482 (N_482,In_342,In_393);
nand U483 (N_483,In_708,In_219);
nor U484 (N_484,In_31,In_724);
and U485 (N_485,In_908,In_919);
xnor U486 (N_486,In_954,In_712);
and U487 (N_487,In_999,In_244);
xor U488 (N_488,In_368,In_296);
nor U489 (N_489,In_736,In_806);
xnor U490 (N_490,In_252,In_645);
and U491 (N_491,In_5,In_892);
nand U492 (N_492,In_251,In_60);
and U493 (N_493,In_167,In_860);
and U494 (N_494,In_895,In_161);
nand U495 (N_495,In_142,In_789);
or U496 (N_496,In_621,In_12);
or U497 (N_497,In_913,In_667);
nor U498 (N_498,In_815,In_261);
nand U499 (N_499,In_912,In_626);
xor U500 (N_500,In_118,In_854);
or U501 (N_501,In_449,In_271);
nor U502 (N_502,In_389,In_688);
and U503 (N_503,In_546,In_712);
or U504 (N_504,In_31,In_270);
xor U505 (N_505,In_305,In_979);
and U506 (N_506,In_855,In_467);
nor U507 (N_507,In_587,In_668);
nor U508 (N_508,In_851,In_319);
and U509 (N_509,In_97,In_528);
or U510 (N_510,In_419,In_676);
or U511 (N_511,In_995,In_146);
nand U512 (N_512,In_456,In_804);
and U513 (N_513,In_225,In_491);
and U514 (N_514,In_869,In_611);
nor U515 (N_515,In_611,In_344);
xnor U516 (N_516,In_180,In_995);
xnor U517 (N_517,In_449,In_367);
nor U518 (N_518,In_58,In_422);
xnor U519 (N_519,In_726,In_484);
or U520 (N_520,In_404,In_880);
or U521 (N_521,In_449,In_222);
nand U522 (N_522,In_951,In_39);
and U523 (N_523,In_682,In_391);
or U524 (N_524,In_29,In_169);
nand U525 (N_525,In_940,In_429);
xor U526 (N_526,In_409,In_614);
nand U527 (N_527,In_563,In_784);
xor U528 (N_528,In_801,In_159);
nand U529 (N_529,In_941,In_787);
nor U530 (N_530,In_387,In_955);
and U531 (N_531,In_37,In_539);
or U532 (N_532,In_47,In_563);
nor U533 (N_533,In_939,In_582);
xor U534 (N_534,In_328,In_426);
nor U535 (N_535,In_509,In_64);
nand U536 (N_536,In_469,In_324);
or U537 (N_537,In_661,In_800);
xnor U538 (N_538,In_347,In_865);
and U539 (N_539,In_796,In_755);
xor U540 (N_540,In_338,In_384);
nor U541 (N_541,In_552,In_436);
xnor U542 (N_542,In_626,In_159);
or U543 (N_543,In_686,In_23);
and U544 (N_544,In_915,In_302);
xnor U545 (N_545,In_367,In_168);
nor U546 (N_546,In_41,In_956);
xnor U547 (N_547,In_929,In_110);
xor U548 (N_548,In_657,In_233);
or U549 (N_549,In_297,In_878);
xor U550 (N_550,In_212,In_57);
nor U551 (N_551,In_244,In_28);
and U552 (N_552,In_819,In_217);
and U553 (N_553,In_991,In_607);
xor U554 (N_554,In_653,In_631);
nand U555 (N_555,In_239,In_996);
and U556 (N_556,In_254,In_402);
xor U557 (N_557,In_576,In_836);
or U558 (N_558,In_409,In_53);
xor U559 (N_559,In_2,In_48);
xnor U560 (N_560,In_989,In_66);
or U561 (N_561,In_102,In_112);
nand U562 (N_562,In_478,In_827);
or U563 (N_563,In_113,In_565);
or U564 (N_564,In_735,In_965);
nor U565 (N_565,In_196,In_829);
nand U566 (N_566,In_344,In_2);
or U567 (N_567,In_29,In_533);
and U568 (N_568,In_123,In_742);
nor U569 (N_569,In_414,In_967);
or U570 (N_570,In_28,In_952);
nand U571 (N_571,In_991,In_47);
xor U572 (N_572,In_591,In_303);
xor U573 (N_573,In_97,In_341);
and U574 (N_574,In_795,In_35);
and U575 (N_575,In_481,In_329);
and U576 (N_576,In_50,In_345);
nor U577 (N_577,In_541,In_929);
nor U578 (N_578,In_362,In_341);
and U579 (N_579,In_608,In_19);
and U580 (N_580,In_607,In_363);
nor U581 (N_581,In_842,In_518);
or U582 (N_582,In_736,In_987);
nand U583 (N_583,In_29,In_330);
nor U584 (N_584,In_207,In_983);
nor U585 (N_585,In_378,In_390);
or U586 (N_586,In_322,In_541);
xor U587 (N_587,In_334,In_849);
and U588 (N_588,In_42,In_341);
or U589 (N_589,In_326,In_851);
or U590 (N_590,In_299,In_209);
or U591 (N_591,In_3,In_679);
and U592 (N_592,In_353,In_473);
and U593 (N_593,In_215,In_564);
nand U594 (N_594,In_183,In_635);
nor U595 (N_595,In_226,In_849);
xnor U596 (N_596,In_644,In_615);
nor U597 (N_597,In_317,In_857);
nor U598 (N_598,In_930,In_685);
or U599 (N_599,In_86,In_854);
nor U600 (N_600,In_521,In_449);
and U601 (N_601,In_811,In_496);
or U602 (N_602,In_551,In_278);
nand U603 (N_603,In_778,In_103);
or U604 (N_604,In_657,In_148);
or U605 (N_605,In_320,In_384);
xor U606 (N_606,In_410,In_781);
and U607 (N_607,In_723,In_713);
nand U608 (N_608,In_210,In_551);
xor U609 (N_609,In_465,In_218);
nor U610 (N_610,In_783,In_670);
and U611 (N_611,In_748,In_942);
and U612 (N_612,In_383,In_914);
nand U613 (N_613,In_930,In_639);
xnor U614 (N_614,In_360,In_211);
and U615 (N_615,In_623,In_59);
and U616 (N_616,In_622,In_863);
and U617 (N_617,In_591,In_459);
nand U618 (N_618,In_771,In_183);
and U619 (N_619,In_755,In_403);
and U620 (N_620,In_644,In_563);
nor U621 (N_621,In_154,In_458);
and U622 (N_622,In_581,In_511);
nor U623 (N_623,In_395,In_102);
nor U624 (N_624,In_952,In_388);
and U625 (N_625,In_619,In_991);
and U626 (N_626,In_803,In_263);
nand U627 (N_627,In_465,In_430);
nand U628 (N_628,In_37,In_846);
and U629 (N_629,In_776,In_946);
nor U630 (N_630,In_668,In_636);
xor U631 (N_631,In_67,In_264);
xor U632 (N_632,In_686,In_196);
nor U633 (N_633,In_76,In_227);
xnor U634 (N_634,In_684,In_505);
xor U635 (N_635,In_35,In_934);
and U636 (N_636,In_801,In_87);
nor U637 (N_637,In_447,In_243);
nor U638 (N_638,In_564,In_42);
xor U639 (N_639,In_174,In_692);
nor U640 (N_640,In_508,In_455);
xnor U641 (N_641,In_223,In_913);
and U642 (N_642,In_715,In_467);
nand U643 (N_643,In_990,In_461);
or U644 (N_644,In_61,In_720);
nand U645 (N_645,In_138,In_112);
xnor U646 (N_646,In_739,In_252);
and U647 (N_647,In_506,In_305);
or U648 (N_648,In_672,In_247);
nor U649 (N_649,In_916,In_388);
and U650 (N_650,In_945,In_246);
nand U651 (N_651,In_490,In_628);
nand U652 (N_652,In_277,In_180);
or U653 (N_653,In_320,In_897);
or U654 (N_654,In_609,In_4);
and U655 (N_655,In_841,In_218);
nand U656 (N_656,In_684,In_138);
or U657 (N_657,In_994,In_995);
and U658 (N_658,In_449,In_285);
nand U659 (N_659,In_257,In_288);
xor U660 (N_660,In_127,In_209);
nand U661 (N_661,In_409,In_491);
and U662 (N_662,In_815,In_93);
and U663 (N_663,In_18,In_890);
or U664 (N_664,In_923,In_335);
and U665 (N_665,In_559,In_71);
nand U666 (N_666,In_227,In_510);
nand U667 (N_667,In_16,In_909);
xor U668 (N_668,In_520,In_986);
or U669 (N_669,In_765,In_837);
and U670 (N_670,In_563,In_586);
nand U671 (N_671,In_700,In_808);
and U672 (N_672,In_705,In_163);
nor U673 (N_673,In_798,In_568);
or U674 (N_674,In_683,In_29);
xnor U675 (N_675,In_509,In_229);
or U676 (N_676,In_675,In_419);
or U677 (N_677,In_888,In_318);
or U678 (N_678,In_431,In_956);
and U679 (N_679,In_274,In_828);
and U680 (N_680,In_220,In_771);
nor U681 (N_681,In_762,In_738);
xor U682 (N_682,In_196,In_264);
nand U683 (N_683,In_542,In_372);
nand U684 (N_684,In_883,In_286);
nand U685 (N_685,In_250,In_303);
or U686 (N_686,In_864,In_849);
xor U687 (N_687,In_67,In_202);
and U688 (N_688,In_815,In_502);
and U689 (N_689,In_991,In_691);
nor U690 (N_690,In_47,In_493);
and U691 (N_691,In_590,In_174);
xnor U692 (N_692,In_480,In_372);
or U693 (N_693,In_874,In_977);
and U694 (N_694,In_689,In_911);
nor U695 (N_695,In_561,In_831);
or U696 (N_696,In_806,In_892);
or U697 (N_697,In_891,In_597);
or U698 (N_698,In_820,In_646);
xor U699 (N_699,In_48,In_651);
nor U700 (N_700,In_609,In_937);
or U701 (N_701,In_148,In_658);
or U702 (N_702,In_296,In_117);
nand U703 (N_703,In_656,In_708);
nand U704 (N_704,In_822,In_701);
or U705 (N_705,In_965,In_688);
or U706 (N_706,In_298,In_834);
and U707 (N_707,In_184,In_458);
nand U708 (N_708,In_475,In_418);
or U709 (N_709,In_139,In_167);
nor U710 (N_710,In_983,In_22);
and U711 (N_711,In_419,In_602);
and U712 (N_712,In_847,In_102);
xor U713 (N_713,In_166,In_622);
nand U714 (N_714,In_779,In_859);
or U715 (N_715,In_386,In_575);
or U716 (N_716,In_444,In_618);
nor U717 (N_717,In_722,In_956);
and U718 (N_718,In_724,In_309);
xnor U719 (N_719,In_382,In_373);
xnor U720 (N_720,In_432,In_483);
nand U721 (N_721,In_789,In_136);
nor U722 (N_722,In_706,In_448);
nor U723 (N_723,In_135,In_622);
or U724 (N_724,In_98,In_825);
nand U725 (N_725,In_935,In_319);
and U726 (N_726,In_984,In_271);
and U727 (N_727,In_508,In_978);
nor U728 (N_728,In_898,In_103);
nand U729 (N_729,In_626,In_3);
and U730 (N_730,In_314,In_562);
xnor U731 (N_731,In_924,In_536);
nand U732 (N_732,In_340,In_892);
nor U733 (N_733,In_638,In_859);
nor U734 (N_734,In_405,In_114);
or U735 (N_735,In_752,In_496);
nor U736 (N_736,In_556,In_541);
nor U737 (N_737,In_364,In_219);
nand U738 (N_738,In_100,In_3);
or U739 (N_739,In_108,In_79);
and U740 (N_740,In_519,In_512);
nand U741 (N_741,In_908,In_530);
and U742 (N_742,In_430,In_515);
nand U743 (N_743,In_511,In_157);
or U744 (N_744,In_42,In_219);
xnor U745 (N_745,In_949,In_447);
nand U746 (N_746,In_901,In_133);
nand U747 (N_747,In_290,In_564);
or U748 (N_748,In_154,In_37);
nand U749 (N_749,In_154,In_125);
or U750 (N_750,In_550,In_601);
xor U751 (N_751,In_405,In_183);
nor U752 (N_752,In_663,In_292);
xor U753 (N_753,In_296,In_995);
xnor U754 (N_754,In_209,In_283);
nor U755 (N_755,In_500,In_480);
nand U756 (N_756,In_993,In_613);
nor U757 (N_757,In_661,In_878);
nand U758 (N_758,In_161,In_494);
nand U759 (N_759,In_584,In_304);
and U760 (N_760,In_595,In_485);
and U761 (N_761,In_992,In_279);
nand U762 (N_762,In_396,In_698);
and U763 (N_763,In_166,In_990);
nor U764 (N_764,In_397,In_713);
xnor U765 (N_765,In_502,In_58);
xnor U766 (N_766,In_991,In_788);
nor U767 (N_767,In_207,In_544);
and U768 (N_768,In_861,In_703);
nor U769 (N_769,In_200,In_36);
or U770 (N_770,In_874,In_246);
xor U771 (N_771,In_106,In_815);
nand U772 (N_772,In_667,In_834);
xnor U773 (N_773,In_109,In_859);
and U774 (N_774,In_517,In_542);
or U775 (N_775,In_673,In_44);
nand U776 (N_776,In_53,In_582);
xnor U777 (N_777,In_830,In_358);
or U778 (N_778,In_756,In_377);
nand U779 (N_779,In_953,In_568);
and U780 (N_780,In_660,In_213);
nor U781 (N_781,In_251,In_395);
xor U782 (N_782,In_887,In_273);
and U783 (N_783,In_955,In_4);
and U784 (N_784,In_724,In_751);
or U785 (N_785,In_77,In_113);
or U786 (N_786,In_950,In_540);
or U787 (N_787,In_380,In_371);
or U788 (N_788,In_8,In_201);
nor U789 (N_789,In_178,In_159);
nor U790 (N_790,In_748,In_145);
nor U791 (N_791,In_910,In_656);
xor U792 (N_792,In_470,In_475);
and U793 (N_793,In_434,In_59);
nand U794 (N_794,In_508,In_877);
and U795 (N_795,In_278,In_80);
and U796 (N_796,In_960,In_152);
xnor U797 (N_797,In_423,In_883);
or U798 (N_798,In_100,In_263);
xnor U799 (N_799,In_489,In_109);
xnor U800 (N_800,In_753,In_111);
and U801 (N_801,In_327,In_873);
xnor U802 (N_802,In_2,In_883);
xor U803 (N_803,In_71,In_357);
or U804 (N_804,In_720,In_708);
and U805 (N_805,In_12,In_905);
xnor U806 (N_806,In_743,In_935);
nor U807 (N_807,In_682,In_76);
or U808 (N_808,In_196,In_109);
or U809 (N_809,In_361,In_311);
or U810 (N_810,In_987,In_268);
nor U811 (N_811,In_859,In_641);
or U812 (N_812,In_846,In_30);
nor U813 (N_813,In_147,In_12);
or U814 (N_814,In_984,In_334);
nor U815 (N_815,In_717,In_660);
or U816 (N_816,In_806,In_872);
xor U817 (N_817,In_695,In_462);
or U818 (N_818,In_283,In_631);
or U819 (N_819,In_323,In_44);
or U820 (N_820,In_176,In_559);
nor U821 (N_821,In_208,In_393);
or U822 (N_822,In_13,In_455);
nand U823 (N_823,In_568,In_620);
or U824 (N_824,In_772,In_322);
or U825 (N_825,In_525,In_161);
nor U826 (N_826,In_185,In_72);
and U827 (N_827,In_749,In_391);
xor U828 (N_828,In_959,In_34);
xor U829 (N_829,In_315,In_160);
or U830 (N_830,In_558,In_829);
and U831 (N_831,In_910,In_550);
xor U832 (N_832,In_106,In_3);
or U833 (N_833,In_211,In_895);
nand U834 (N_834,In_528,In_621);
nor U835 (N_835,In_697,In_70);
nor U836 (N_836,In_863,In_582);
or U837 (N_837,In_602,In_620);
nand U838 (N_838,In_21,In_537);
or U839 (N_839,In_933,In_649);
xnor U840 (N_840,In_466,In_793);
xnor U841 (N_841,In_824,In_564);
xor U842 (N_842,In_746,In_322);
xnor U843 (N_843,In_851,In_740);
or U844 (N_844,In_298,In_602);
xor U845 (N_845,In_562,In_523);
xor U846 (N_846,In_811,In_906);
and U847 (N_847,In_608,In_929);
xor U848 (N_848,In_607,In_885);
or U849 (N_849,In_708,In_382);
nor U850 (N_850,In_584,In_758);
or U851 (N_851,In_16,In_836);
and U852 (N_852,In_838,In_699);
and U853 (N_853,In_347,In_910);
and U854 (N_854,In_544,In_668);
xnor U855 (N_855,In_383,In_616);
and U856 (N_856,In_567,In_641);
nor U857 (N_857,In_374,In_656);
nor U858 (N_858,In_360,In_155);
nor U859 (N_859,In_192,In_550);
and U860 (N_860,In_389,In_306);
nand U861 (N_861,In_699,In_633);
or U862 (N_862,In_597,In_984);
xnor U863 (N_863,In_392,In_506);
xnor U864 (N_864,In_478,In_975);
nand U865 (N_865,In_836,In_15);
nand U866 (N_866,In_88,In_799);
or U867 (N_867,In_706,In_161);
and U868 (N_868,In_8,In_407);
and U869 (N_869,In_215,In_290);
nor U870 (N_870,In_768,In_825);
nor U871 (N_871,In_414,In_172);
nand U872 (N_872,In_261,In_902);
nor U873 (N_873,In_200,In_286);
nand U874 (N_874,In_701,In_472);
nand U875 (N_875,In_94,In_215);
or U876 (N_876,In_875,In_592);
and U877 (N_877,In_947,In_941);
xor U878 (N_878,In_719,In_538);
nor U879 (N_879,In_21,In_860);
and U880 (N_880,In_360,In_748);
and U881 (N_881,In_391,In_822);
nand U882 (N_882,In_384,In_309);
nand U883 (N_883,In_418,In_80);
xnor U884 (N_884,In_588,In_871);
xnor U885 (N_885,In_925,In_693);
nand U886 (N_886,In_27,In_860);
or U887 (N_887,In_344,In_275);
nor U888 (N_888,In_811,In_202);
nand U889 (N_889,In_120,In_449);
xnor U890 (N_890,In_463,In_741);
or U891 (N_891,In_542,In_401);
nor U892 (N_892,In_991,In_37);
nor U893 (N_893,In_495,In_436);
or U894 (N_894,In_11,In_976);
xor U895 (N_895,In_187,In_442);
nor U896 (N_896,In_124,In_662);
or U897 (N_897,In_683,In_761);
nor U898 (N_898,In_314,In_749);
xnor U899 (N_899,In_928,In_524);
nand U900 (N_900,In_400,In_728);
nand U901 (N_901,In_208,In_234);
nand U902 (N_902,In_678,In_998);
or U903 (N_903,In_135,In_849);
xor U904 (N_904,In_624,In_540);
nand U905 (N_905,In_384,In_776);
and U906 (N_906,In_811,In_620);
and U907 (N_907,In_432,In_149);
xor U908 (N_908,In_630,In_994);
nor U909 (N_909,In_123,In_89);
and U910 (N_910,In_504,In_831);
nor U911 (N_911,In_345,In_429);
and U912 (N_912,In_610,In_134);
or U913 (N_913,In_60,In_852);
or U914 (N_914,In_126,In_992);
xor U915 (N_915,In_326,In_983);
and U916 (N_916,In_113,In_708);
nand U917 (N_917,In_244,In_611);
xor U918 (N_918,In_559,In_159);
or U919 (N_919,In_73,In_505);
nor U920 (N_920,In_232,In_972);
or U921 (N_921,In_327,In_441);
or U922 (N_922,In_914,In_9);
nor U923 (N_923,In_92,In_560);
or U924 (N_924,In_215,In_250);
and U925 (N_925,In_538,In_722);
or U926 (N_926,In_589,In_93);
or U927 (N_927,In_180,In_975);
and U928 (N_928,In_329,In_526);
or U929 (N_929,In_724,In_762);
xor U930 (N_930,In_153,In_401);
xor U931 (N_931,In_741,In_313);
and U932 (N_932,In_339,In_303);
xnor U933 (N_933,In_956,In_268);
and U934 (N_934,In_340,In_444);
and U935 (N_935,In_178,In_12);
xnor U936 (N_936,In_20,In_559);
xnor U937 (N_937,In_212,In_736);
or U938 (N_938,In_758,In_989);
and U939 (N_939,In_106,In_377);
and U940 (N_940,In_568,In_856);
nor U941 (N_941,In_120,In_700);
or U942 (N_942,In_677,In_809);
nor U943 (N_943,In_725,In_216);
or U944 (N_944,In_534,In_243);
and U945 (N_945,In_504,In_855);
xor U946 (N_946,In_725,In_27);
nand U947 (N_947,In_894,In_716);
xnor U948 (N_948,In_783,In_976);
nand U949 (N_949,In_549,In_786);
nand U950 (N_950,In_186,In_24);
and U951 (N_951,In_753,In_278);
nor U952 (N_952,In_86,In_824);
nor U953 (N_953,In_398,In_35);
or U954 (N_954,In_398,In_439);
nand U955 (N_955,In_716,In_646);
xor U956 (N_956,In_847,In_372);
or U957 (N_957,In_921,In_842);
or U958 (N_958,In_709,In_593);
nor U959 (N_959,In_763,In_269);
nand U960 (N_960,In_397,In_142);
xnor U961 (N_961,In_467,In_112);
nor U962 (N_962,In_319,In_857);
xnor U963 (N_963,In_38,In_973);
nand U964 (N_964,In_989,In_634);
nand U965 (N_965,In_555,In_674);
nor U966 (N_966,In_586,In_456);
or U967 (N_967,In_133,In_598);
or U968 (N_968,In_254,In_622);
or U969 (N_969,In_390,In_940);
nor U970 (N_970,In_447,In_974);
nand U971 (N_971,In_35,In_422);
nand U972 (N_972,In_172,In_439);
nor U973 (N_973,In_323,In_514);
xnor U974 (N_974,In_640,In_501);
nand U975 (N_975,In_357,In_565);
nor U976 (N_976,In_355,In_58);
and U977 (N_977,In_337,In_696);
and U978 (N_978,In_911,In_722);
nor U979 (N_979,In_320,In_722);
xnor U980 (N_980,In_280,In_630);
or U981 (N_981,In_297,In_379);
xor U982 (N_982,In_151,In_588);
xnor U983 (N_983,In_393,In_196);
xnor U984 (N_984,In_943,In_999);
xnor U985 (N_985,In_197,In_49);
nand U986 (N_986,In_520,In_623);
xor U987 (N_987,In_321,In_363);
nor U988 (N_988,In_705,In_316);
or U989 (N_989,In_295,In_434);
or U990 (N_990,In_889,In_143);
or U991 (N_991,In_359,In_437);
or U992 (N_992,In_682,In_631);
nand U993 (N_993,In_478,In_978);
nand U994 (N_994,In_821,In_559);
or U995 (N_995,In_469,In_844);
nand U996 (N_996,In_247,In_740);
and U997 (N_997,In_18,In_458);
xnor U998 (N_998,In_988,In_472);
nand U999 (N_999,In_495,In_203);
nor U1000 (N_1000,N_89,N_280);
nand U1001 (N_1001,N_438,N_743);
and U1002 (N_1002,N_856,N_433);
and U1003 (N_1003,N_57,N_481);
nor U1004 (N_1004,N_647,N_942);
xor U1005 (N_1005,N_722,N_936);
or U1006 (N_1006,N_712,N_126);
nor U1007 (N_1007,N_714,N_723);
xnor U1008 (N_1008,N_278,N_307);
xnor U1009 (N_1009,N_223,N_962);
xor U1010 (N_1010,N_678,N_716);
or U1011 (N_1011,N_948,N_197);
or U1012 (N_1012,N_19,N_950);
nor U1013 (N_1013,N_901,N_104);
xor U1014 (N_1014,N_116,N_83);
nor U1015 (N_1015,N_381,N_883);
nor U1016 (N_1016,N_398,N_885);
or U1017 (N_1017,N_400,N_189);
and U1018 (N_1018,N_734,N_1);
nor U1019 (N_1019,N_40,N_485);
xnor U1020 (N_1020,N_148,N_933);
or U1021 (N_1021,N_269,N_365);
nor U1022 (N_1022,N_429,N_87);
and U1023 (N_1023,N_477,N_984);
or U1024 (N_1024,N_426,N_855);
xnor U1025 (N_1025,N_501,N_779);
xnor U1026 (N_1026,N_699,N_820);
and U1027 (N_1027,N_389,N_26);
or U1028 (N_1028,N_548,N_739);
nand U1029 (N_1029,N_757,N_783);
or U1030 (N_1030,N_985,N_634);
xnor U1031 (N_1031,N_169,N_193);
nor U1032 (N_1032,N_931,N_82);
nor U1033 (N_1033,N_141,N_661);
nor U1034 (N_1034,N_164,N_685);
or U1035 (N_1035,N_778,N_997);
nor U1036 (N_1036,N_547,N_785);
xnor U1037 (N_1037,N_36,N_688);
and U1038 (N_1038,N_406,N_371);
nand U1039 (N_1039,N_875,N_515);
xor U1040 (N_1040,N_907,N_585);
xnor U1041 (N_1041,N_915,N_6);
nand U1042 (N_1042,N_848,N_562);
nor U1043 (N_1043,N_62,N_430);
nor U1044 (N_1044,N_495,N_940);
or U1045 (N_1045,N_965,N_608);
xnor U1046 (N_1046,N_420,N_506);
and U1047 (N_1047,N_640,N_409);
nor U1048 (N_1048,N_145,N_606);
xnor U1049 (N_1049,N_695,N_612);
and U1050 (N_1050,N_806,N_160);
nand U1051 (N_1051,N_241,N_7);
nor U1052 (N_1052,N_528,N_424);
nand U1053 (N_1053,N_541,N_527);
nand U1054 (N_1054,N_349,N_687);
or U1055 (N_1055,N_375,N_407);
and U1056 (N_1056,N_120,N_938);
or U1057 (N_1057,N_159,N_318);
or U1058 (N_1058,N_708,N_296);
and U1059 (N_1059,N_86,N_469);
xnor U1060 (N_1060,N_54,N_21);
nand U1061 (N_1061,N_799,N_232);
and U1062 (N_1062,N_403,N_761);
xnor U1063 (N_1063,N_786,N_298);
nor U1064 (N_1064,N_973,N_968);
xnor U1065 (N_1065,N_465,N_224);
and U1066 (N_1066,N_452,N_411);
xor U1067 (N_1067,N_720,N_509);
nor U1068 (N_1068,N_928,N_330);
and U1069 (N_1069,N_66,N_216);
or U1070 (N_1070,N_368,N_348);
nand U1071 (N_1071,N_233,N_168);
nor U1072 (N_1072,N_643,N_989);
or U1073 (N_1073,N_914,N_890);
or U1074 (N_1074,N_179,N_366);
xor U1075 (N_1075,N_898,N_98);
or U1076 (N_1076,N_815,N_762);
or U1077 (N_1077,N_203,N_602);
nor U1078 (N_1078,N_462,N_352);
or U1079 (N_1079,N_386,N_851);
or U1080 (N_1080,N_604,N_871);
xor U1081 (N_1081,N_442,N_844);
or U1082 (N_1082,N_570,N_759);
or U1083 (N_1083,N_839,N_670);
or U1084 (N_1084,N_102,N_443);
nand U1085 (N_1085,N_202,N_79);
and U1086 (N_1086,N_747,N_990);
xnor U1087 (N_1087,N_510,N_649);
nor U1088 (N_1088,N_118,N_291);
or U1089 (N_1089,N_282,N_52);
nand U1090 (N_1090,N_285,N_369);
or U1091 (N_1091,N_563,N_831);
nor U1092 (N_1092,N_693,N_618);
nor U1093 (N_1093,N_326,N_628);
and U1094 (N_1094,N_564,N_740);
xnor U1095 (N_1095,N_853,N_932);
or U1096 (N_1096,N_493,N_698);
nand U1097 (N_1097,N_674,N_12);
or U1098 (N_1098,N_733,N_467);
nand U1099 (N_1099,N_43,N_724);
nor U1100 (N_1100,N_484,N_713);
nor U1101 (N_1101,N_954,N_617);
or U1102 (N_1102,N_359,N_561);
or U1103 (N_1103,N_621,N_935);
nor U1104 (N_1104,N_391,N_921);
and U1105 (N_1105,N_867,N_217);
or U1106 (N_1106,N_721,N_152);
and U1107 (N_1107,N_434,N_696);
xnor U1108 (N_1108,N_309,N_669);
and U1109 (N_1109,N_502,N_525);
or U1110 (N_1110,N_227,N_73);
xor U1111 (N_1111,N_554,N_206);
and U1112 (N_1112,N_3,N_270);
xor U1113 (N_1113,N_956,N_777);
nand U1114 (N_1114,N_908,N_392);
nand U1115 (N_1115,N_792,N_150);
and U1116 (N_1116,N_81,N_646);
or U1117 (N_1117,N_922,N_824);
nand U1118 (N_1118,N_945,N_395);
nand U1119 (N_1119,N_814,N_436);
nor U1120 (N_1120,N_133,N_362);
nor U1121 (N_1121,N_313,N_966);
and U1122 (N_1122,N_245,N_847);
nand U1123 (N_1123,N_446,N_553);
or U1124 (N_1124,N_95,N_195);
nand U1125 (N_1125,N_300,N_252);
nand U1126 (N_1126,N_125,N_187);
and U1127 (N_1127,N_417,N_837);
nor U1128 (N_1128,N_995,N_219);
xnor U1129 (N_1129,N_297,N_742);
and U1130 (N_1130,N_85,N_648);
nor U1131 (N_1131,N_25,N_703);
and U1132 (N_1132,N_658,N_850);
nand U1133 (N_1133,N_346,N_673);
xnor U1134 (N_1134,N_741,N_97);
xnor U1135 (N_1135,N_801,N_876);
nand U1136 (N_1136,N_754,N_745);
or U1137 (N_1137,N_819,N_797);
xnor U1138 (N_1138,N_153,N_490);
xor U1139 (N_1139,N_939,N_751);
xnor U1140 (N_1140,N_170,N_644);
nor U1141 (N_1141,N_124,N_715);
nor U1142 (N_1142,N_225,N_412);
or U1143 (N_1143,N_770,N_51);
nor U1144 (N_1144,N_763,N_335);
or U1145 (N_1145,N_136,N_692);
nand U1146 (N_1146,N_384,N_635);
nor U1147 (N_1147,N_672,N_807);
and U1148 (N_1148,N_753,N_857);
xor U1149 (N_1149,N_657,N_457);
and U1150 (N_1150,N_190,N_926);
nor U1151 (N_1151,N_737,N_882);
nand U1152 (N_1152,N_677,N_222);
and U1153 (N_1153,N_70,N_828);
nor U1154 (N_1154,N_886,N_524);
or U1155 (N_1155,N_292,N_48);
nor U1156 (N_1156,N_394,N_47);
and U1157 (N_1157,N_415,N_286);
and U1158 (N_1158,N_378,N_571);
xor U1159 (N_1159,N_684,N_466);
and U1160 (N_1160,N_979,N_470);
and U1161 (N_1161,N_825,N_781);
nor U1162 (N_1162,N_479,N_100);
or U1163 (N_1163,N_860,N_147);
or U1164 (N_1164,N_315,N_611);
nand U1165 (N_1165,N_103,N_884);
nor U1166 (N_1166,N_870,N_271);
or U1167 (N_1167,N_772,N_513);
xnor U1168 (N_1168,N_877,N_499);
and U1169 (N_1169,N_631,N_239);
or U1170 (N_1170,N_846,N_607);
nand U1171 (N_1171,N_749,N_71);
nor U1172 (N_1172,N_755,N_795);
and U1173 (N_1173,N_30,N_836);
xnor U1174 (N_1174,N_555,N_887);
nor U1175 (N_1175,N_302,N_999);
and U1176 (N_1176,N_551,N_803);
and U1177 (N_1177,N_941,N_603);
nor U1178 (N_1178,N_538,N_530);
nor U1179 (N_1179,N_730,N_592);
and U1180 (N_1180,N_162,N_306);
nor U1181 (N_1181,N_128,N_199);
or U1182 (N_1182,N_172,N_651);
xnor U1183 (N_1183,N_702,N_72);
nor U1184 (N_1184,N_557,N_486);
or U1185 (N_1185,N_937,N_341);
nand U1186 (N_1186,N_192,N_154);
nand U1187 (N_1187,N_460,N_879);
or U1188 (N_1188,N_812,N_397);
nand U1189 (N_1189,N_257,N_494);
and U1190 (N_1190,N_68,N_28);
or U1191 (N_1191,N_333,N_709);
and U1192 (N_1192,N_188,N_44);
nand U1193 (N_1193,N_221,N_983);
xnor U1194 (N_1194,N_157,N_918);
and U1195 (N_1195,N_993,N_827);
or U1196 (N_1196,N_266,N_949);
and U1197 (N_1197,N_756,N_717);
and U1198 (N_1198,N_238,N_284);
nand U1199 (N_1199,N_858,N_235);
and U1200 (N_1200,N_67,N_580);
xor U1201 (N_1201,N_642,N_787);
xnor U1202 (N_1202,N_934,N_947);
nand U1203 (N_1203,N_960,N_959);
or U1204 (N_1204,N_975,N_101);
or U1205 (N_1205,N_500,N_166);
xnor U1206 (N_1206,N_121,N_322);
and U1207 (N_1207,N_23,N_872);
and U1208 (N_1208,N_393,N_289);
or U1209 (N_1209,N_881,N_22);
nand U1210 (N_1210,N_982,N_9);
nand U1211 (N_1211,N_594,N_171);
and U1212 (N_1212,N_957,N_588);
nand U1213 (N_1213,N_41,N_324);
xor U1214 (N_1214,N_295,N_789);
nand U1215 (N_1215,N_953,N_680);
xnor U1216 (N_1216,N_632,N_76);
xnor U1217 (N_1217,N_215,N_212);
nor U1218 (N_1218,N_345,N_458);
and U1219 (N_1219,N_483,N_109);
or U1220 (N_1220,N_589,N_182);
or U1221 (N_1221,N_784,N_732);
nand U1222 (N_1222,N_163,N_334);
xnor U1223 (N_1223,N_771,N_523);
or U1224 (N_1224,N_343,N_633);
nand U1225 (N_1225,N_60,N_609);
and U1226 (N_1226,N_913,N_808);
xnor U1227 (N_1227,N_361,N_288);
xnor U1228 (N_1228,N_559,N_177);
nor U1229 (N_1229,N_181,N_579);
xnor U1230 (N_1230,N_432,N_259);
nor U1231 (N_1231,N_536,N_868);
or U1232 (N_1232,N_310,N_521);
or U1233 (N_1233,N_593,N_277);
xnor U1234 (N_1234,N_208,N_888);
nor U1235 (N_1235,N_707,N_952);
nor U1236 (N_1236,N_809,N_645);
nor U1237 (N_1237,N_818,N_90);
nor U1238 (N_1238,N_437,N_262);
and U1239 (N_1239,N_210,N_201);
nand U1240 (N_1240,N_569,N_600);
or U1241 (N_1241,N_655,N_242);
xnor U1242 (N_1242,N_676,N_880);
or U1243 (N_1243,N_519,N_549);
nand U1244 (N_1244,N_878,N_294);
xor U1245 (N_1245,N_760,N_75);
nor U1246 (N_1246,N_186,N_834);
xnor U1247 (N_1247,N_823,N_654);
xnor U1248 (N_1248,N_69,N_613);
nand U1249 (N_1249,N_970,N_972);
nor U1250 (N_1250,N_767,N_805);
or U1251 (N_1251,N_574,N_32);
nand U1252 (N_1252,N_852,N_327);
or U1253 (N_1253,N_254,N_923);
or U1254 (N_1254,N_260,N_115);
xnor U1255 (N_1255,N_161,N_17);
or U1256 (N_1256,N_665,N_690);
and U1257 (N_1257,N_246,N_287);
nor U1258 (N_1258,N_314,N_447);
and U1259 (N_1259,N_376,N_336);
or U1260 (N_1260,N_273,N_796);
and U1261 (N_1261,N_813,N_987);
xor U1262 (N_1262,N_627,N_639);
nor U1263 (N_1263,N_545,N_976);
and U1264 (N_1264,N_800,N_453);
and U1265 (N_1265,N_92,N_573);
nor U1266 (N_1266,N_977,N_16);
or U1267 (N_1267,N_183,N_304);
and U1268 (N_1268,N_616,N_841);
and U1269 (N_1269,N_129,N_149);
or U1270 (N_1270,N_508,N_526);
xor U1271 (N_1271,N_427,N_146);
and U1272 (N_1272,N_917,N_782);
xnor U1273 (N_1273,N_961,N_862);
nand U1274 (N_1274,N_625,N_414);
nand U1275 (N_1275,N_546,N_752);
nand U1276 (N_1276,N_374,N_719);
or U1277 (N_1277,N_971,N_107);
or U1278 (N_1278,N_272,N_231);
and U1279 (N_1279,N_236,N_464);
nand U1280 (N_1280,N_487,N_401);
nor U1281 (N_1281,N_822,N_49);
xor U1282 (N_1282,N_283,N_463);
or U1283 (N_1283,N_736,N_590);
nor U1284 (N_1284,N_838,N_175);
nand U1285 (N_1285,N_380,N_893);
nor U1286 (N_1286,N_768,N_511);
or U1287 (N_1287,N_816,N_533);
nand U1288 (N_1288,N_110,N_725);
nor U1289 (N_1289,N_58,N_111);
nor U1290 (N_1290,N_379,N_731);
and U1291 (N_1291,N_200,N_728);
and U1292 (N_1292,N_354,N_583);
nor U1293 (N_1293,N_45,N_247);
xor U1294 (N_1294,N_675,N_587);
and U1295 (N_1295,N_980,N_8);
xnor U1296 (N_1296,N_710,N_958);
nand U1297 (N_1297,N_492,N_912);
and U1298 (N_1298,N_861,N_402);
and U1299 (N_1299,N_441,N_550);
xnor U1300 (N_1300,N_864,N_610);
and U1301 (N_1301,N_620,N_896);
nor U1302 (N_1302,N_531,N_951);
or U1303 (N_1303,N_764,N_165);
xor U1304 (N_1304,N_38,N_207);
or U1305 (N_1305,N_775,N_63);
nor U1306 (N_1306,N_735,N_11);
and U1307 (N_1307,N_205,N_944);
nor U1308 (N_1308,N_135,N_798);
and U1309 (N_1309,N_388,N_243);
nand U1310 (N_1310,N_84,N_817);
and U1311 (N_1311,N_15,N_840);
xnor U1312 (N_1312,N_566,N_355);
xnor U1313 (N_1313,N_14,N_105);
xnor U1314 (N_1314,N_694,N_347);
nand U1315 (N_1315,N_671,N_228);
or U1316 (N_1316,N_804,N_480);
or U1317 (N_1317,N_29,N_843);
nor U1318 (N_1318,N_577,N_320);
xor U1319 (N_1319,N_906,N_705);
xnor U1320 (N_1320,N_276,N_473);
xnor U1321 (N_1321,N_230,N_489);
xnor U1322 (N_1322,N_664,N_529);
or U1323 (N_1323,N_930,N_405);
xor U1324 (N_1324,N_176,N_444);
or U1325 (N_1325,N_399,N_601);
and U1326 (N_1326,N_404,N_614);
xor U1327 (N_1327,N_650,N_339);
nor U1328 (N_1328,N_24,N_211);
nand U1329 (N_1329,N_130,N_138);
and U1330 (N_1330,N_619,N_156);
and U1331 (N_1331,N_905,N_372);
nor U1332 (N_1332,N_543,N_660);
and U1333 (N_1333,N_899,N_475);
nor U1334 (N_1334,N_532,N_377);
or U1335 (N_1335,N_582,N_729);
xnor U1336 (N_1336,N_773,N_927);
nor U1337 (N_1337,N_383,N_849);
xnor U1338 (N_1338,N_516,N_65);
nand U1339 (N_1339,N_638,N_468);
and U1340 (N_1340,N_488,N_476);
and U1341 (N_1341,N_350,N_167);
nand U1342 (N_1342,N_209,N_630);
xnor U1343 (N_1343,N_367,N_988);
nor U1344 (N_1344,N_408,N_578);
xnor U1345 (N_1345,N_435,N_364);
nor U1346 (N_1346,N_268,N_251);
nor U1347 (N_1347,N_666,N_558);
and U1348 (N_1348,N_974,N_303);
and U1349 (N_1349,N_418,N_615);
and U1350 (N_1350,N_185,N_390);
nor U1351 (N_1351,N_679,N_869);
or U1352 (N_1352,N_535,N_652);
nor U1353 (N_1353,N_667,N_978);
nor U1354 (N_1354,N_910,N_833);
nand U1355 (N_1355,N_560,N_214);
nand U1356 (N_1356,N_27,N_450);
nand U1357 (N_1357,N_496,N_13);
xor U1358 (N_1358,N_832,N_39);
nand U1359 (N_1359,N_173,N_37);
and U1360 (N_1360,N_718,N_565);
nor U1361 (N_1361,N_338,N_991);
xnor U1362 (N_1362,N_80,N_174);
nor U1363 (N_1363,N_682,N_794);
nor U1364 (N_1364,N_963,N_512);
nor U1365 (N_1365,N_422,N_264);
and U1366 (N_1366,N_581,N_534);
or U1367 (N_1367,N_889,N_108);
or U1368 (N_1368,N_123,N_0);
xor U1369 (N_1369,N_842,N_440);
and U1370 (N_1370,N_498,N_293);
nor U1371 (N_1371,N_373,N_77);
xor U1372 (N_1372,N_213,N_586);
xnor U1373 (N_1373,N_88,N_605);
xor U1374 (N_1374,N_91,N_568);
nand U1375 (N_1375,N_131,N_419);
nand U1376 (N_1376,N_854,N_357);
or U1377 (N_1377,N_316,N_522);
and U1378 (N_1378,N_50,N_637);
nor U1379 (N_1379,N_964,N_311);
or U1380 (N_1380,N_358,N_503);
nor U1381 (N_1381,N_428,N_552);
xor U1382 (N_1382,N_916,N_994);
nand U1383 (N_1383,N_451,N_829);
nand U1384 (N_1384,N_758,N_55);
or U1385 (N_1385,N_117,N_790);
or U1386 (N_1386,N_598,N_668);
or U1387 (N_1387,N_356,N_727);
and U1388 (N_1388,N_31,N_659);
nor U1389 (N_1389,N_629,N_810);
xnor U1390 (N_1390,N_793,N_337);
nand U1391 (N_1391,N_226,N_929);
nor U1392 (N_1392,N_455,N_744);
and U1393 (N_1393,N_765,N_35);
or U1394 (N_1394,N_184,N_517);
and U1395 (N_1395,N_53,N_248);
nand U1396 (N_1396,N_2,N_396);
xnor U1397 (N_1397,N_701,N_955);
xor U1398 (N_1398,N_461,N_94);
nand U1399 (N_1399,N_151,N_416);
xnor U1400 (N_1400,N_865,N_328);
nor U1401 (N_1401,N_42,N_267);
nor U1402 (N_1402,N_774,N_471);
nor U1403 (N_1403,N_624,N_599);
or U1404 (N_1404,N_250,N_370);
nand U1405 (N_1405,N_290,N_265);
xor U1406 (N_1406,N_874,N_139);
nand U1407 (N_1407,N_454,N_218);
or U1408 (N_1408,N_491,N_902);
or U1409 (N_1409,N_738,N_360);
xor U1410 (N_1410,N_623,N_237);
nor U1411 (N_1411,N_113,N_726);
or U1412 (N_1412,N_256,N_96);
or U1413 (N_1413,N_788,N_497);
or U1414 (N_1414,N_700,N_5);
or U1415 (N_1415,N_132,N_308);
xnor U1416 (N_1416,N_776,N_340);
and U1417 (N_1417,N_969,N_329);
and U1418 (N_1418,N_750,N_894);
or U1419 (N_1419,N_46,N_998);
nand U1420 (N_1420,N_421,N_301);
nand U1421 (N_1421,N_382,N_279);
nor U1422 (N_1422,N_911,N_924);
nor U1423 (N_1423,N_540,N_996);
nor U1424 (N_1424,N_584,N_261);
xnor U1425 (N_1425,N_514,N_194);
nor U1426 (N_1426,N_683,N_255);
xor U1427 (N_1427,N_826,N_697);
xnor U1428 (N_1428,N_925,N_576);
xor U1429 (N_1429,N_992,N_689);
nand U1430 (N_1430,N_537,N_681);
or U1431 (N_1431,N_342,N_704);
nor U1432 (N_1432,N_472,N_119);
xnor U1433 (N_1433,N_410,N_263);
and U1434 (N_1434,N_281,N_572);
or U1435 (N_1435,N_691,N_539);
nand U1436 (N_1436,N_74,N_240);
nand U1437 (N_1437,N_321,N_198);
or U1438 (N_1438,N_114,N_802);
nor U1439 (N_1439,N_4,N_196);
nand U1440 (N_1440,N_413,N_791);
nor U1441 (N_1441,N_439,N_662);
nor U1442 (N_1442,N_542,N_20);
and U1443 (N_1443,N_748,N_122);
xnor U1444 (N_1444,N_137,N_895);
nor U1445 (N_1445,N_474,N_10);
nand U1446 (N_1446,N_61,N_423);
or U1447 (N_1447,N_332,N_449);
and U1448 (N_1448,N_835,N_686);
nor U1449 (N_1449,N_567,N_319);
xnor U1450 (N_1450,N_244,N_595);
nor U1451 (N_1451,N_305,N_18);
nor U1452 (N_1452,N_155,N_344);
nand U1453 (N_1453,N_920,N_178);
nor U1454 (N_1454,N_909,N_641);
nand U1455 (N_1455,N_597,N_981);
and U1456 (N_1456,N_191,N_143);
nor U1457 (N_1457,N_863,N_385);
xor U1458 (N_1458,N_919,N_158);
nor U1459 (N_1459,N_946,N_220);
or U1460 (N_1460,N_544,N_892);
xnor U1461 (N_1461,N_312,N_204);
nand U1462 (N_1462,N_866,N_591);
nor U1463 (N_1463,N_711,N_518);
and U1464 (N_1464,N_33,N_127);
and U1465 (N_1465,N_504,N_323);
xnor U1466 (N_1466,N_274,N_106);
xnor U1467 (N_1467,N_431,N_78);
nand U1468 (N_1468,N_325,N_520);
nand U1469 (N_1469,N_859,N_93);
nand U1470 (N_1470,N_112,N_766);
nor U1471 (N_1471,N_140,N_351);
nand U1472 (N_1472,N_811,N_636);
xor U1473 (N_1473,N_459,N_903);
xor U1474 (N_1474,N_656,N_425);
nor U1475 (N_1475,N_821,N_331);
xnor U1476 (N_1476,N_507,N_596);
nor U1477 (N_1477,N_897,N_448);
nor U1478 (N_1478,N_353,N_275);
nand U1479 (N_1479,N_622,N_904);
xor U1480 (N_1480,N_99,N_663);
or U1481 (N_1481,N_317,N_769);
nor U1482 (N_1482,N_626,N_229);
xor U1483 (N_1483,N_943,N_144);
or U1484 (N_1484,N_746,N_900);
and U1485 (N_1485,N_505,N_56);
nand U1486 (N_1486,N_134,N_234);
and U1487 (N_1487,N_456,N_253);
or U1488 (N_1488,N_180,N_653);
and U1489 (N_1489,N_830,N_706);
or U1490 (N_1490,N_249,N_258);
xnor U1491 (N_1491,N_556,N_967);
and U1492 (N_1492,N_575,N_34);
or U1493 (N_1493,N_845,N_363);
xor U1494 (N_1494,N_59,N_873);
xor U1495 (N_1495,N_142,N_891);
nor U1496 (N_1496,N_299,N_482);
nand U1497 (N_1497,N_387,N_445);
nor U1498 (N_1498,N_478,N_986);
nand U1499 (N_1499,N_780,N_64);
xor U1500 (N_1500,N_465,N_249);
nand U1501 (N_1501,N_596,N_752);
and U1502 (N_1502,N_993,N_762);
nand U1503 (N_1503,N_99,N_15);
xnor U1504 (N_1504,N_110,N_699);
and U1505 (N_1505,N_245,N_825);
and U1506 (N_1506,N_834,N_718);
xnor U1507 (N_1507,N_26,N_73);
nor U1508 (N_1508,N_353,N_756);
nor U1509 (N_1509,N_725,N_854);
and U1510 (N_1510,N_77,N_855);
nand U1511 (N_1511,N_29,N_94);
nand U1512 (N_1512,N_122,N_260);
or U1513 (N_1513,N_53,N_796);
and U1514 (N_1514,N_234,N_710);
or U1515 (N_1515,N_96,N_942);
nor U1516 (N_1516,N_248,N_269);
xor U1517 (N_1517,N_788,N_966);
nand U1518 (N_1518,N_723,N_621);
xnor U1519 (N_1519,N_388,N_662);
and U1520 (N_1520,N_907,N_567);
and U1521 (N_1521,N_382,N_564);
and U1522 (N_1522,N_974,N_555);
and U1523 (N_1523,N_564,N_468);
or U1524 (N_1524,N_749,N_3);
and U1525 (N_1525,N_141,N_758);
and U1526 (N_1526,N_295,N_628);
or U1527 (N_1527,N_647,N_891);
or U1528 (N_1528,N_67,N_249);
nor U1529 (N_1529,N_487,N_643);
xor U1530 (N_1530,N_135,N_185);
nor U1531 (N_1531,N_820,N_813);
and U1532 (N_1532,N_934,N_720);
or U1533 (N_1533,N_110,N_229);
xor U1534 (N_1534,N_159,N_611);
xor U1535 (N_1535,N_281,N_37);
or U1536 (N_1536,N_168,N_684);
xor U1537 (N_1537,N_715,N_689);
nand U1538 (N_1538,N_458,N_431);
xnor U1539 (N_1539,N_712,N_497);
and U1540 (N_1540,N_997,N_455);
nand U1541 (N_1541,N_159,N_99);
nor U1542 (N_1542,N_145,N_63);
nand U1543 (N_1543,N_196,N_587);
and U1544 (N_1544,N_581,N_96);
or U1545 (N_1545,N_626,N_764);
xor U1546 (N_1546,N_70,N_800);
or U1547 (N_1547,N_328,N_955);
and U1548 (N_1548,N_755,N_971);
xnor U1549 (N_1549,N_446,N_520);
nand U1550 (N_1550,N_854,N_115);
xor U1551 (N_1551,N_938,N_632);
nand U1552 (N_1552,N_673,N_657);
nor U1553 (N_1553,N_606,N_316);
xnor U1554 (N_1554,N_578,N_122);
nand U1555 (N_1555,N_150,N_237);
and U1556 (N_1556,N_509,N_525);
or U1557 (N_1557,N_713,N_204);
or U1558 (N_1558,N_82,N_124);
and U1559 (N_1559,N_677,N_100);
nor U1560 (N_1560,N_379,N_162);
and U1561 (N_1561,N_473,N_593);
and U1562 (N_1562,N_716,N_709);
xor U1563 (N_1563,N_556,N_175);
and U1564 (N_1564,N_878,N_677);
or U1565 (N_1565,N_541,N_694);
xnor U1566 (N_1566,N_228,N_825);
or U1567 (N_1567,N_717,N_388);
xor U1568 (N_1568,N_695,N_964);
nand U1569 (N_1569,N_379,N_930);
nand U1570 (N_1570,N_527,N_831);
nand U1571 (N_1571,N_571,N_26);
and U1572 (N_1572,N_716,N_223);
and U1573 (N_1573,N_587,N_637);
nand U1574 (N_1574,N_16,N_744);
and U1575 (N_1575,N_818,N_248);
and U1576 (N_1576,N_159,N_698);
and U1577 (N_1577,N_152,N_165);
xnor U1578 (N_1578,N_271,N_736);
nor U1579 (N_1579,N_105,N_907);
or U1580 (N_1580,N_290,N_825);
xnor U1581 (N_1581,N_671,N_616);
and U1582 (N_1582,N_198,N_194);
or U1583 (N_1583,N_124,N_398);
xor U1584 (N_1584,N_219,N_369);
xor U1585 (N_1585,N_400,N_134);
or U1586 (N_1586,N_724,N_676);
and U1587 (N_1587,N_807,N_787);
and U1588 (N_1588,N_69,N_546);
or U1589 (N_1589,N_391,N_216);
or U1590 (N_1590,N_957,N_199);
nand U1591 (N_1591,N_305,N_314);
nand U1592 (N_1592,N_773,N_215);
or U1593 (N_1593,N_887,N_435);
or U1594 (N_1594,N_582,N_746);
nand U1595 (N_1595,N_234,N_190);
nor U1596 (N_1596,N_57,N_680);
nor U1597 (N_1597,N_691,N_189);
nand U1598 (N_1598,N_980,N_875);
or U1599 (N_1599,N_127,N_208);
nor U1600 (N_1600,N_291,N_882);
or U1601 (N_1601,N_63,N_949);
nor U1602 (N_1602,N_676,N_328);
and U1603 (N_1603,N_601,N_60);
nand U1604 (N_1604,N_47,N_990);
nor U1605 (N_1605,N_843,N_427);
xor U1606 (N_1606,N_729,N_223);
xor U1607 (N_1607,N_729,N_830);
and U1608 (N_1608,N_534,N_177);
and U1609 (N_1609,N_692,N_117);
xnor U1610 (N_1610,N_944,N_323);
and U1611 (N_1611,N_903,N_110);
or U1612 (N_1612,N_209,N_130);
and U1613 (N_1613,N_168,N_492);
nor U1614 (N_1614,N_857,N_171);
nor U1615 (N_1615,N_197,N_633);
or U1616 (N_1616,N_108,N_234);
nand U1617 (N_1617,N_969,N_846);
and U1618 (N_1618,N_273,N_615);
or U1619 (N_1619,N_393,N_995);
nor U1620 (N_1620,N_175,N_102);
nor U1621 (N_1621,N_891,N_42);
nor U1622 (N_1622,N_179,N_796);
or U1623 (N_1623,N_700,N_984);
or U1624 (N_1624,N_863,N_815);
nand U1625 (N_1625,N_69,N_972);
nor U1626 (N_1626,N_839,N_237);
and U1627 (N_1627,N_304,N_588);
xor U1628 (N_1628,N_391,N_984);
xnor U1629 (N_1629,N_79,N_543);
nor U1630 (N_1630,N_39,N_948);
or U1631 (N_1631,N_279,N_569);
and U1632 (N_1632,N_937,N_825);
or U1633 (N_1633,N_825,N_211);
xnor U1634 (N_1634,N_760,N_529);
and U1635 (N_1635,N_654,N_362);
or U1636 (N_1636,N_69,N_770);
xor U1637 (N_1637,N_528,N_403);
xnor U1638 (N_1638,N_42,N_852);
nand U1639 (N_1639,N_794,N_995);
nor U1640 (N_1640,N_850,N_233);
or U1641 (N_1641,N_64,N_310);
or U1642 (N_1642,N_54,N_72);
nor U1643 (N_1643,N_381,N_605);
xnor U1644 (N_1644,N_392,N_955);
and U1645 (N_1645,N_106,N_808);
nand U1646 (N_1646,N_255,N_336);
nor U1647 (N_1647,N_740,N_576);
or U1648 (N_1648,N_999,N_562);
or U1649 (N_1649,N_800,N_293);
and U1650 (N_1650,N_762,N_699);
xor U1651 (N_1651,N_128,N_935);
nand U1652 (N_1652,N_706,N_301);
xnor U1653 (N_1653,N_753,N_815);
nor U1654 (N_1654,N_152,N_836);
or U1655 (N_1655,N_590,N_368);
nor U1656 (N_1656,N_226,N_273);
nand U1657 (N_1657,N_575,N_570);
nor U1658 (N_1658,N_838,N_158);
xnor U1659 (N_1659,N_330,N_289);
nor U1660 (N_1660,N_512,N_834);
xnor U1661 (N_1661,N_908,N_865);
and U1662 (N_1662,N_621,N_139);
and U1663 (N_1663,N_611,N_439);
xnor U1664 (N_1664,N_724,N_840);
xor U1665 (N_1665,N_468,N_959);
and U1666 (N_1666,N_41,N_55);
or U1667 (N_1667,N_423,N_702);
and U1668 (N_1668,N_974,N_923);
nand U1669 (N_1669,N_983,N_95);
xor U1670 (N_1670,N_136,N_752);
or U1671 (N_1671,N_68,N_172);
xnor U1672 (N_1672,N_500,N_400);
nor U1673 (N_1673,N_794,N_442);
xnor U1674 (N_1674,N_24,N_272);
xnor U1675 (N_1675,N_427,N_296);
xnor U1676 (N_1676,N_993,N_269);
xnor U1677 (N_1677,N_927,N_334);
and U1678 (N_1678,N_915,N_320);
nor U1679 (N_1679,N_990,N_16);
xnor U1680 (N_1680,N_556,N_718);
and U1681 (N_1681,N_319,N_818);
xnor U1682 (N_1682,N_580,N_909);
xnor U1683 (N_1683,N_401,N_471);
or U1684 (N_1684,N_483,N_66);
xnor U1685 (N_1685,N_416,N_725);
or U1686 (N_1686,N_534,N_342);
nand U1687 (N_1687,N_692,N_736);
nor U1688 (N_1688,N_987,N_401);
or U1689 (N_1689,N_604,N_798);
nand U1690 (N_1690,N_538,N_711);
nor U1691 (N_1691,N_238,N_821);
xor U1692 (N_1692,N_519,N_530);
xnor U1693 (N_1693,N_987,N_854);
or U1694 (N_1694,N_233,N_680);
and U1695 (N_1695,N_42,N_476);
xnor U1696 (N_1696,N_198,N_758);
or U1697 (N_1697,N_104,N_910);
xor U1698 (N_1698,N_684,N_609);
nor U1699 (N_1699,N_902,N_357);
nand U1700 (N_1700,N_410,N_348);
nand U1701 (N_1701,N_628,N_528);
xnor U1702 (N_1702,N_248,N_578);
and U1703 (N_1703,N_292,N_174);
or U1704 (N_1704,N_157,N_60);
xor U1705 (N_1705,N_180,N_636);
nand U1706 (N_1706,N_897,N_156);
nand U1707 (N_1707,N_54,N_830);
or U1708 (N_1708,N_462,N_55);
xnor U1709 (N_1709,N_20,N_663);
and U1710 (N_1710,N_292,N_886);
or U1711 (N_1711,N_683,N_166);
and U1712 (N_1712,N_241,N_332);
xor U1713 (N_1713,N_440,N_463);
xor U1714 (N_1714,N_802,N_119);
nor U1715 (N_1715,N_939,N_576);
or U1716 (N_1716,N_773,N_844);
nor U1717 (N_1717,N_876,N_910);
xnor U1718 (N_1718,N_612,N_7);
or U1719 (N_1719,N_811,N_648);
nor U1720 (N_1720,N_589,N_971);
xor U1721 (N_1721,N_369,N_772);
and U1722 (N_1722,N_92,N_721);
and U1723 (N_1723,N_533,N_380);
nor U1724 (N_1724,N_414,N_425);
or U1725 (N_1725,N_904,N_350);
xor U1726 (N_1726,N_433,N_550);
and U1727 (N_1727,N_962,N_337);
nand U1728 (N_1728,N_852,N_540);
and U1729 (N_1729,N_886,N_339);
xor U1730 (N_1730,N_515,N_376);
and U1731 (N_1731,N_733,N_36);
nand U1732 (N_1732,N_298,N_658);
and U1733 (N_1733,N_567,N_445);
nor U1734 (N_1734,N_37,N_224);
and U1735 (N_1735,N_440,N_152);
xor U1736 (N_1736,N_603,N_523);
nand U1737 (N_1737,N_529,N_847);
xnor U1738 (N_1738,N_362,N_843);
and U1739 (N_1739,N_492,N_495);
nor U1740 (N_1740,N_968,N_111);
and U1741 (N_1741,N_852,N_264);
xor U1742 (N_1742,N_809,N_89);
or U1743 (N_1743,N_46,N_212);
or U1744 (N_1744,N_154,N_144);
nor U1745 (N_1745,N_245,N_195);
nor U1746 (N_1746,N_918,N_765);
and U1747 (N_1747,N_100,N_3);
nand U1748 (N_1748,N_822,N_464);
xor U1749 (N_1749,N_422,N_768);
nor U1750 (N_1750,N_998,N_315);
or U1751 (N_1751,N_140,N_332);
and U1752 (N_1752,N_685,N_609);
or U1753 (N_1753,N_821,N_423);
nand U1754 (N_1754,N_479,N_956);
and U1755 (N_1755,N_740,N_874);
and U1756 (N_1756,N_115,N_23);
nor U1757 (N_1757,N_149,N_716);
nor U1758 (N_1758,N_644,N_10);
nor U1759 (N_1759,N_422,N_746);
nand U1760 (N_1760,N_288,N_928);
nor U1761 (N_1761,N_461,N_625);
xor U1762 (N_1762,N_505,N_589);
and U1763 (N_1763,N_862,N_617);
and U1764 (N_1764,N_645,N_225);
and U1765 (N_1765,N_807,N_730);
nand U1766 (N_1766,N_325,N_414);
xnor U1767 (N_1767,N_586,N_91);
or U1768 (N_1768,N_513,N_315);
or U1769 (N_1769,N_547,N_370);
xor U1770 (N_1770,N_952,N_56);
nand U1771 (N_1771,N_449,N_290);
xor U1772 (N_1772,N_175,N_409);
and U1773 (N_1773,N_273,N_299);
or U1774 (N_1774,N_909,N_42);
and U1775 (N_1775,N_59,N_131);
and U1776 (N_1776,N_90,N_26);
or U1777 (N_1777,N_227,N_850);
nor U1778 (N_1778,N_734,N_24);
nor U1779 (N_1779,N_656,N_245);
and U1780 (N_1780,N_43,N_296);
nand U1781 (N_1781,N_52,N_544);
and U1782 (N_1782,N_398,N_426);
nor U1783 (N_1783,N_37,N_862);
or U1784 (N_1784,N_756,N_706);
nor U1785 (N_1785,N_626,N_282);
nand U1786 (N_1786,N_128,N_383);
or U1787 (N_1787,N_830,N_385);
nand U1788 (N_1788,N_156,N_111);
nand U1789 (N_1789,N_442,N_891);
nand U1790 (N_1790,N_961,N_966);
nor U1791 (N_1791,N_926,N_630);
nor U1792 (N_1792,N_33,N_169);
nand U1793 (N_1793,N_41,N_588);
or U1794 (N_1794,N_293,N_329);
or U1795 (N_1795,N_993,N_950);
nor U1796 (N_1796,N_986,N_267);
or U1797 (N_1797,N_344,N_192);
or U1798 (N_1798,N_145,N_886);
and U1799 (N_1799,N_19,N_382);
xnor U1800 (N_1800,N_656,N_393);
nand U1801 (N_1801,N_440,N_753);
and U1802 (N_1802,N_981,N_335);
and U1803 (N_1803,N_950,N_48);
nand U1804 (N_1804,N_619,N_495);
and U1805 (N_1805,N_565,N_100);
or U1806 (N_1806,N_586,N_218);
or U1807 (N_1807,N_115,N_165);
xnor U1808 (N_1808,N_825,N_628);
xnor U1809 (N_1809,N_831,N_355);
and U1810 (N_1810,N_891,N_915);
or U1811 (N_1811,N_433,N_101);
and U1812 (N_1812,N_264,N_800);
nand U1813 (N_1813,N_969,N_946);
xor U1814 (N_1814,N_610,N_140);
and U1815 (N_1815,N_961,N_750);
nor U1816 (N_1816,N_88,N_246);
or U1817 (N_1817,N_188,N_117);
nor U1818 (N_1818,N_800,N_620);
or U1819 (N_1819,N_878,N_455);
nor U1820 (N_1820,N_837,N_499);
xor U1821 (N_1821,N_149,N_5);
nand U1822 (N_1822,N_26,N_499);
xor U1823 (N_1823,N_853,N_42);
and U1824 (N_1824,N_287,N_225);
and U1825 (N_1825,N_786,N_473);
nor U1826 (N_1826,N_322,N_726);
nor U1827 (N_1827,N_889,N_148);
or U1828 (N_1828,N_294,N_307);
nor U1829 (N_1829,N_160,N_150);
or U1830 (N_1830,N_282,N_16);
nand U1831 (N_1831,N_870,N_553);
and U1832 (N_1832,N_868,N_15);
xor U1833 (N_1833,N_929,N_81);
nand U1834 (N_1834,N_387,N_618);
and U1835 (N_1835,N_471,N_744);
or U1836 (N_1836,N_382,N_243);
nor U1837 (N_1837,N_702,N_460);
and U1838 (N_1838,N_891,N_737);
and U1839 (N_1839,N_862,N_35);
xnor U1840 (N_1840,N_832,N_424);
or U1841 (N_1841,N_48,N_947);
nor U1842 (N_1842,N_545,N_474);
or U1843 (N_1843,N_876,N_622);
xnor U1844 (N_1844,N_626,N_523);
nand U1845 (N_1845,N_824,N_771);
nor U1846 (N_1846,N_298,N_94);
xor U1847 (N_1847,N_474,N_979);
nor U1848 (N_1848,N_558,N_362);
and U1849 (N_1849,N_703,N_706);
or U1850 (N_1850,N_861,N_578);
nand U1851 (N_1851,N_327,N_545);
and U1852 (N_1852,N_989,N_460);
and U1853 (N_1853,N_202,N_835);
nand U1854 (N_1854,N_969,N_235);
xor U1855 (N_1855,N_273,N_149);
xnor U1856 (N_1856,N_545,N_635);
or U1857 (N_1857,N_685,N_956);
or U1858 (N_1858,N_723,N_903);
nor U1859 (N_1859,N_80,N_446);
nand U1860 (N_1860,N_735,N_711);
or U1861 (N_1861,N_309,N_454);
or U1862 (N_1862,N_337,N_632);
nor U1863 (N_1863,N_925,N_854);
and U1864 (N_1864,N_601,N_755);
and U1865 (N_1865,N_291,N_907);
xnor U1866 (N_1866,N_894,N_674);
and U1867 (N_1867,N_731,N_471);
or U1868 (N_1868,N_740,N_179);
or U1869 (N_1869,N_616,N_379);
or U1870 (N_1870,N_786,N_77);
or U1871 (N_1871,N_452,N_785);
xnor U1872 (N_1872,N_964,N_291);
nand U1873 (N_1873,N_346,N_587);
xor U1874 (N_1874,N_766,N_905);
and U1875 (N_1875,N_258,N_64);
xor U1876 (N_1876,N_67,N_941);
or U1877 (N_1877,N_511,N_959);
nand U1878 (N_1878,N_966,N_162);
xor U1879 (N_1879,N_663,N_201);
nand U1880 (N_1880,N_939,N_278);
xor U1881 (N_1881,N_40,N_748);
xor U1882 (N_1882,N_843,N_218);
nand U1883 (N_1883,N_651,N_831);
and U1884 (N_1884,N_100,N_376);
nor U1885 (N_1885,N_381,N_86);
and U1886 (N_1886,N_899,N_218);
nand U1887 (N_1887,N_887,N_702);
nor U1888 (N_1888,N_593,N_177);
nor U1889 (N_1889,N_801,N_630);
nor U1890 (N_1890,N_7,N_901);
xnor U1891 (N_1891,N_383,N_103);
xor U1892 (N_1892,N_596,N_992);
nand U1893 (N_1893,N_834,N_388);
nand U1894 (N_1894,N_645,N_357);
or U1895 (N_1895,N_298,N_665);
or U1896 (N_1896,N_40,N_235);
or U1897 (N_1897,N_134,N_926);
and U1898 (N_1898,N_835,N_384);
xnor U1899 (N_1899,N_925,N_408);
or U1900 (N_1900,N_400,N_787);
nor U1901 (N_1901,N_116,N_603);
or U1902 (N_1902,N_949,N_322);
nand U1903 (N_1903,N_45,N_486);
xnor U1904 (N_1904,N_408,N_226);
and U1905 (N_1905,N_73,N_282);
nand U1906 (N_1906,N_168,N_648);
nand U1907 (N_1907,N_144,N_720);
nor U1908 (N_1908,N_799,N_2);
nor U1909 (N_1909,N_720,N_567);
xor U1910 (N_1910,N_178,N_693);
nand U1911 (N_1911,N_480,N_662);
xnor U1912 (N_1912,N_595,N_558);
and U1913 (N_1913,N_342,N_103);
and U1914 (N_1914,N_426,N_785);
nand U1915 (N_1915,N_921,N_707);
and U1916 (N_1916,N_900,N_842);
and U1917 (N_1917,N_997,N_502);
or U1918 (N_1918,N_657,N_485);
nand U1919 (N_1919,N_691,N_222);
nand U1920 (N_1920,N_869,N_622);
nand U1921 (N_1921,N_456,N_871);
xnor U1922 (N_1922,N_459,N_157);
xor U1923 (N_1923,N_431,N_101);
xor U1924 (N_1924,N_765,N_33);
xnor U1925 (N_1925,N_476,N_47);
nand U1926 (N_1926,N_906,N_225);
nor U1927 (N_1927,N_720,N_221);
nand U1928 (N_1928,N_584,N_235);
nand U1929 (N_1929,N_938,N_590);
nor U1930 (N_1930,N_942,N_466);
nor U1931 (N_1931,N_467,N_314);
and U1932 (N_1932,N_192,N_700);
or U1933 (N_1933,N_10,N_963);
nand U1934 (N_1934,N_978,N_470);
nor U1935 (N_1935,N_584,N_115);
xor U1936 (N_1936,N_283,N_466);
or U1937 (N_1937,N_753,N_996);
or U1938 (N_1938,N_712,N_789);
or U1939 (N_1939,N_28,N_418);
and U1940 (N_1940,N_32,N_962);
and U1941 (N_1941,N_856,N_69);
nor U1942 (N_1942,N_30,N_333);
or U1943 (N_1943,N_290,N_140);
and U1944 (N_1944,N_239,N_729);
nor U1945 (N_1945,N_96,N_47);
and U1946 (N_1946,N_133,N_557);
and U1947 (N_1947,N_505,N_177);
xor U1948 (N_1948,N_682,N_107);
xor U1949 (N_1949,N_2,N_620);
or U1950 (N_1950,N_956,N_501);
nor U1951 (N_1951,N_638,N_713);
nor U1952 (N_1952,N_806,N_458);
or U1953 (N_1953,N_649,N_371);
nor U1954 (N_1954,N_139,N_497);
and U1955 (N_1955,N_100,N_109);
nor U1956 (N_1956,N_397,N_563);
nor U1957 (N_1957,N_287,N_844);
and U1958 (N_1958,N_902,N_931);
and U1959 (N_1959,N_826,N_430);
xnor U1960 (N_1960,N_777,N_187);
nand U1961 (N_1961,N_438,N_338);
nand U1962 (N_1962,N_898,N_872);
or U1963 (N_1963,N_191,N_431);
or U1964 (N_1964,N_928,N_113);
or U1965 (N_1965,N_417,N_616);
or U1966 (N_1966,N_409,N_784);
nor U1967 (N_1967,N_68,N_639);
nand U1968 (N_1968,N_166,N_170);
or U1969 (N_1969,N_22,N_297);
and U1970 (N_1970,N_85,N_907);
and U1971 (N_1971,N_393,N_323);
nor U1972 (N_1972,N_104,N_918);
nor U1973 (N_1973,N_812,N_478);
and U1974 (N_1974,N_197,N_3);
nor U1975 (N_1975,N_186,N_176);
or U1976 (N_1976,N_953,N_128);
or U1977 (N_1977,N_954,N_529);
xnor U1978 (N_1978,N_895,N_148);
and U1979 (N_1979,N_173,N_782);
nand U1980 (N_1980,N_641,N_6);
nand U1981 (N_1981,N_438,N_515);
nor U1982 (N_1982,N_421,N_617);
nand U1983 (N_1983,N_850,N_862);
nor U1984 (N_1984,N_914,N_840);
and U1985 (N_1985,N_180,N_2);
nand U1986 (N_1986,N_227,N_9);
or U1987 (N_1987,N_634,N_1);
or U1988 (N_1988,N_852,N_100);
nor U1989 (N_1989,N_966,N_936);
xnor U1990 (N_1990,N_632,N_820);
and U1991 (N_1991,N_845,N_771);
and U1992 (N_1992,N_376,N_847);
and U1993 (N_1993,N_62,N_433);
nand U1994 (N_1994,N_620,N_32);
and U1995 (N_1995,N_146,N_471);
xor U1996 (N_1996,N_872,N_80);
nand U1997 (N_1997,N_456,N_834);
xnor U1998 (N_1998,N_838,N_860);
xor U1999 (N_1999,N_754,N_221);
or U2000 (N_2000,N_1133,N_1726);
nand U2001 (N_2001,N_1320,N_1582);
nand U2002 (N_2002,N_1387,N_1712);
nand U2003 (N_2003,N_1772,N_1833);
xor U2004 (N_2004,N_1161,N_1944);
and U2005 (N_2005,N_1274,N_1023);
nor U2006 (N_2006,N_1733,N_1987);
nor U2007 (N_2007,N_1267,N_1044);
and U2008 (N_2008,N_1006,N_1301);
and U2009 (N_2009,N_1437,N_1426);
xnor U2010 (N_2010,N_1655,N_1538);
nand U2011 (N_2011,N_1674,N_1911);
or U2012 (N_2012,N_1839,N_1816);
or U2013 (N_2013,N_1366,N_1436);
nand U2014 (N_2014,N_1998,N_1590);
and U2015 (N_2015,N_1012,N_1572);
or U2016 (N_2016,N_1302,N_1790);
xor U2017 (N_2017,N_1996,N_1009);
nand U2018 (N_2018,N_1810,N_1725);
and U2019 (N_2019,N_1693,N_1865);
nor U2020 (N_2020,N_1030,N_1941);
xnor U2021 (N_2021,N_1187,N_1760);
nand U2022 (N_2022,N_1995,N_1908);
xnor U2023 (N_2023,N_1073,N_1668);
nor U2024 (N_2024,N_1936,N_1069);
xor U2025 (N_2025,N_1315,N_1993);
nor U2026 (N_2026,N_1515,N_1127);
xor U2027 (N_2027,N_1625,N_1978);
xor U2028 (N_2028,N_1679,N_1505);
and U2029 (N_2029,N_1076,N_1412);
or U2030 (N_2030,N_1094,N_1164);
and U2031 (N_2031,N_1016,N_1769);
nor U2032 (N_2032,N_1319,N_1165);
nand U2033 (N_2033,N_1308,N_1789);
nand U2034 (N_2034,N_1705,N_1932);
and U2035 (N_2035,N_1248,N_1162);
or U2036 (N_2036,N_1214,N_1869);
or U2037 (N_2037,N_1748,N_1672);
and U2038 (N_2038,N_1149,N_1395);
nand U2039 (N_2039,N_1128,N_1496);
or U2040 (N_2040,N_1943,N_1078);
or U2041 (N_2041,N_1380,N_1928);
and U2042 (N_2042,N_1844,N_1531);
nand U2043 (N_2043,N_1629,N_1153);
or U2044 (N_2044,N_1106,N_1322);
xor U2045 (N_2045,N_1517,N_1554);
and U2046 (N_2046,N_1093,N_1592);
nand U2047 (N_2047,N_1820,N_1438);
nor U2048 (N_2048,N_1120,N_1964);
xor U2049 (N_2049,N_1883,N_1049);
or U2050 (N_2050,N_1469,N_1776);
xnor U2051 (N_2051,N_1033,N_1229);
or U2052 (N_2052,N_1495,N_1367);
xnor U2053 (N_2053,N_1497,N_1738);
and U2054 (N_2054,N_1854,N_1491);
or U2055 (N_2055,N_1027,N_1986);
xnor U2056 (N_2056,N_1340,N_1291);
and U2057 (N_2057,N_1793,N_1130);
nor U2058 (N_2058,N_1018,N_1970);
and U2059 (N_2059,N_1186,N_1870);
or U2060 (N_2060,N_1107,N_1602);
nor U2061 (N_2061,N_1599,N_1206);
nor U2062 (N_2062,N_1604,N_1036);
xor U2063 (N_2063,N_1535,N_1550);
and U2064 (N_2064,N_1917,N_1935);
xor U2065 (N_2065,N_1266,N_1452);
nor U2066 (N_2066,N_1293,N_1193);
and U2067 (N_2067,N_1342,N_1798);
nor U2068 (N_2068,N_1905,N_1965);
nand U2069 (N_2069,N_1696,N_1887);
or U2070 (N_2070,N_1971,N_1851);
xnor U2071 (N_2071,N_1821,N_1809);
or U2072 (N_2072,N_1539,N_1290);
nor U2073 (N_2073,N_1191,N_1524);
nand U2074 (N_2074,N_1371,N_1551);
nand U2075 (N_2075,N_1796,N_1005);
nor U2076 (N_2076,N_1628,N_1251);
nand U2077 (N_2077,N_1516,N_1994);
xnor U2078 (N_2078,N_1203,N_1451);
and U2079 (N_2079,N_1511,N_1050);
or U2080 (N_2080,N_1972,N_1382);
nand U2081 (N_2081,N_1472,N_1202);
xnor U2082 (N_2082,N_1209,N_1278);
xnor U2083 (N_2083,N_1889,N_1638);
nand U2084 (N_2084,N_1727,N_1912);
xnor U2085 (N_2085,N_1415,N_1147);
and U2086 (N_2086,N_1091,N_1457);
or U2087 (N_2087,N_1349,N_1347);
and U2088 (N_2088,N_1878,N_1581);
nand U2089 (N_2089,N_1010,N_1873);
nand U2090 (N_2090,N_1823,N_1721);
or U2091 (N_2091,N_1242,N_1510);
nor U2092 (N_2092,N_1846,N_1985);
nor U2093 (N_2093,N_1700,N_1541);
or U2094 (N_2094,N_1653,N_1435);
xor U2095 (N_2095,N_1428,N_1609);
and U2096 (N_2096,N_1868,N_1766);
xor U2097 (N_2097,N_1453,N_1037);
nand U2098 (N_2098,N_1194,N_1190);
nand U2099 (N_2099,N_1683,N_1556);
and U2100 (N_2100,N_1463,N_1734);
and U2101 (N_2101,N_1362,N_1470);
nand U2102 (N_2102,N_1126,N_1975);
xor U2103 (N_2103,N_1396,N_1536);
nand U2104 (N_2104,N_1490,N_1228);
nor U2105 (N_2105,N_1205,N_1480);
xnor U2106 (N_2106,N_1068,N_1400);
or U2107 (N_2107,N_1794,N_1601);
nand U2108 (N_2108,N_1974,N_1560);
nand U2109 (N_2109,N_1719,N_1246);
nor U2110 (N_2110,N_1298,N_1060);
or U2111 (N_2111,N_1624,N_1166);
or U2112 (N_2112,N_1377,N_1421);
or U2113 (N_2113,N_1294,N_1742);
nand U2114 (N_2114,N_1717,N_1692);
xor U2115 (N_2115,N_1888,N_1462);
nor U2116 (N_2116,N_1355,N_1389);
or U2117 (N_2117,N_1019,N_1979);
xor U2118 (N_2118,N_1284,N_1432);
nand U2119 (N_2119,N_1427,N_1276);
nand U2120 (N_2120,N_1117,N_1782);
and U2121 (N_2121,N_1634,N_1695);
and U2122 (N_2122,N_1420,N_1336);
or U2123 (N_2123,N_1144,N_1761);
nor U2124 (N_2124,N_1927,N_1337);
and U2125 (N_2125,N_1441,N_1097);
xor U2126 (N_2126,N_1559,N_1578);
nor U2127 (N_2127,N_1157,N_1894);
nand U2128 (N_2128,N_1842,N_1408);
nor U2129 (N_2129,N_1805,N_1052);
nor U2130 (N_2130,N_1170,N_1208);
xor U2131 (N_2131,N_1759,N_1623);
nor U2132 (N_2132,N_1233,N_1813);
or U2133 (N_2133,N_1397,N_1989);
xnor U2134 (N_2134,N_1720,N_1746);
xnor U2135 (N_2135,N_1501,N_1652);
xor U2136 (N_2136,N_1607,N_1024);
nand U2137 (N_2137,N_1710,N_1825);
nor U2138 (N_2138,N_1200,N_1697);
and U2139 (N_2139,N_1473,N_1401);
xor U2140 (N_2140,N_1113,N_1788);
or U2141 (N_2141,N_1585,N_1708);
or U2142 (N_2142,N_1704,N_1882);
nor U2143 (N_2143,N_1022,N_1409);
nand U2144 (N_2144,N_1283,N_1500);
and U2145 (N_2145,N_1264,N_1521);
and U2146 (N_2146,N_1475,N_1178);
nor U2147 (N_2147,N_1771,N_1151);
nand U2148 (N_2148,N_1456,N_1621);
xor U2149 (N_2149,N_1573,N_1881);
nor U2150 (N_2150,N_1826,N_1923);
nand U2151 (N_2151,N_1552,N_1185);
xnor U2152 (N_2152,N_1534,N_1584);
and U2153 (N_2153,N_1474,N_1485);
nor U2154 (N_2154,N_1884,N_1433);
xnor U2155 (N_2155,N_1984,N_1583);
nand U2156 (N_2156,N_1523,N_1920);
xnor U2157 (N_2157,N_1612,N_1391);
xor U2158 (N_2158,N_1661,N_1890);
nor U2159 (N_2159,N_1952,N_1969);
and U2160 (N_2160,N_1632,N_1047);
nor U2161 (N_2161,N_1241,N_1425);
xnor U2162 (N_2162,N_1885,N_1353);
nor U2163 (N_2163,N_1945,N_1031);
nand U2164 (N_2164,N_1657,N_1177);
and U2165 (N_2165,N_1478,N_1174);
nand U2166 (N_2166,N_1611,N_1296);
and U2167 (N_2167,N_1747,N_1892);
and U2168 (N_2168,N_1137,N_1756);
nor U2169 (N_2169,N_1099,N_1508);
nor U2170 (N_2170,N_1083,N_1386);
or U2171 (N_2171,N_1728,N_1350);
xnor U2172 (N_2172,N_1758,N_1306);
or U2173 (N_2173,N_1188,N_1011);
xnor U2174 (N_2174,N_1731,N_1840);
nor U2175 (N_2175,N_1279,N_1953);
or U2176 (N_2176,N_1877,N_1393);
nor U2177 (N_2177,N_1215,N_1419);
or U2178 (N_2178,N_1297,N_1703);
or U2179 (N_2179,N_1730,N_1783);
nand U2180 (N_2180,N_1225,N_1981);
or U2181 (N_2181,N_1247,N_1256);
nand U2182 (N_2182,N_1848,N_1627);
and U2183 (N_2183,N_1586,N_1822);
or U2184 (N_2184,N_1471,N_1236);
and U2185 (N_2185,N_1930,N_1001);
and U2186 (N_2186,N_1828,N_1381);
and U2187 (N_2187,N_1836,N_1896);
xnor U2188 (N_2188,N_1218,N_1814);
and U2189 (N_2189,N_1614,N_1802);
nand U2190 (N_2190,N_1152,N_1392);
xnor U2191 (N_2191,N_1286,N_1711);
nor U2192 (N_2192,N_1980,N_1680);
xor U2193 (N_2193,N_1937,N_1767);
xnor U2194 (N_2194,N_1918,N_1707);
nor U2195 (N_2195,N_1316,N_1258);
and U2196 (N_2196,N_1785,N_1343);
or U2197 (N_2197,N_1647,N_1968);
xor U2198 (N_2198,N_1057,N_1588);
xnor U2199 (N_2199,N_1909,N_1253);
or U2200 (N_2200,N_1077,N_1555);
or U2201 (N_2201,N_1613,N_1872);
nor U2202 (N_2202,N_1558,N_1325);
and U2203 (N_2203,N_1014,N_1715);
and U2204 (N_2204,N_1212,N_1675);
xnor U2205 (N_2205,N_1548,N_1042);
and U2206 (N_2206,N_1459,N_1780);
nor U2207 (N_2207,N_1824,N_1956);
and U2208 (N_2208,N_1667,N_1455);
nand U2209 (N_2209,N_1633,N_1891);
xor U2210 (N_2210,N_1481,N_1313);
or U2211 (N_2211,N_1338,N_1189);
xnor U2212 (N_2212,N_1143,N_1095);
or U2213 (N_2213,N_1973,N_1673);
or U2214 (N_2214,N_1352,N_1509);
xnor U2215 (N_2215,N_1656,N_1866);
and U2216 (N_2216,N_1741,N_1394);
and U2217 (N_2217,N_1317,N_1196);
xnor U2218 (N_2218,N_1230,N_1440);
or U2219 (N_2219,N_1357,N_1285);
nor U2220 (N_2220,N_1053,N_1493);
nor U2221 (N_2221,N_1071,N_1811);
or U2222 (N_2222,N_1015,N_1026);
xor U2223 (N_2223,N_1346,N_1915);
and U2224 (N_2224,N_1684,N_1713);
and U2225 (N_2225,N_1874,N_1801);
and U2226 (N_2226,N_1950,N_1411);
or U2227 (N_2227,N_1959,N_1089);
and U2228 (N_2228,N_1931,N_1136);
nor U2229 (N_2229,N_1886,N_1533);
xor U2230 (N_2230,N_1863,N_1791);
nand U2231 (N_2231,N_1487,N_1605);
nand U2232 (N_2232,N_1983,N_1201);
nor U2233 (N_2233,N_1041,N_1365);
or U2234 (N_2234,N_1512,N_1879);
and U2235 (N_2235,N_1139,N_1620);
or U2236 (N_2236,N_1723,N_1942);
xor U2237 (N_2237,N_1379,N_1418);
and U2238 (N_2238,N_1775,N_1902);
and U2239 (N_2239,N_1477,N_1368);
and U2240 (N_2240,N_1402,N_1537);
nor U2241 (N_2241,N_1171,N_1580);
nand U2242 (N_2242,N_1341,N_1017);
nor U2243 (N_2243,N_1035,N_1806);
nand U2244 (N_2244,N_1563,N_1864);
and U2245 (N_2245,N_1145,N_1665);
and U2246 (N_2246,N_1792,N_1640);
nand U2247 (N_2247,N_1125,N_1948);
and U2248 (N_2248,N_1514,N_1378);
or U2249 (N_2249,N_1857,N_1079);
and U2250 (N_2250,N_1960,N_1739);
nand U2251 (N_2251,N_1195,N_1273);
or U2252 (N_2252,N_1255,N_1528);
nand U2253 (N_2253,N_1111,N_1797);
xor U2254 (N_2254,N_1483,N_1910);
or U2255 (N_2255,N_1765,N_1114);
or U2256 (N_2256,N_1641,N_1268);
or U2257 (N_2257,N_1764,N_1670);
or U2258 (N_2258,N_1630,N_1043);
nand U2259 (N_2259,N_1744,N_1450);
and U2260 (N_2260,N_1466,N_1770);
and U2261 (N_2261,N_1900,N_1321);
nor U2262 (N_2262,N_1754,N_1527);
xnor U2263 (N_2263,N_1694,N_1282);
or U2264 (N_2264,N_1413,N_1658);
xnor U2265 (N_2265,N_1992,N_1646);
or U2266 (N_2266,N_1217,N_1499);
xor U2267 (N_2267,N_1837,N_1061);
nor U2268 (N_2268,N_1300,N_1706);
or U2269 (N_2269,N_1880,N_1543);
nor U2270 (N_2270,N_1102,N_1988);
or U2271 (N_2271,N_1732,N_1654);
nand U2272 (N_2272,N_1399,N_1269);
nand U2273 (N_2273,N_1587,N_1309);
xor U2274 (N_2274,N_1360,N_1176);
nor U2275 (N_2275,N_1991,N_1688);
and U2276 (N_2276,N_1778,N_1498);
xnor U2277 (N_2277,N_1522,N_1561);
or U2278 (N_2278,N_1954,N_1940);
nand U2279 (N_2279,N_1351,N_1227);
nor U2280 (N_2280,N_1616,N_1687);
nand U2281 (N_2281,N_1664,N_1398);
and U2282 (N_2282,N_1540,N_1513);
xnor U2283 (N_2283,N_1048,N_1596);
and U2284 (N_2284,N_1461,N_1383);
xor U2285 (N_2285,N_1216,N_1446);
xnor U2286 (N_2286,N_1025,N_1179);
nand U2287 (N_2287,N_1210,N_1224);
nor U2288 (N_2288,N_1635,N_1299);
nand U2289 (N_2289,N_1239,N_1566);
or U2290 (N_2290,N_1310,N_1406);
nor U2291 (N_2291,N_1096,N_1831);
nand U2292 (N_2292,N_1807,N_1122);
xnor U2293 (N_2293,N_1020,N_1716);
nor U2294 (N_2294,N_1181,N_1682);
nand U2295 (N_2295,N_1547,N_1729);
and U2296 (N_2296,N_1407,N_1116);
or U2297 (N_2297,N_1356,N_1295);
xnor U2298 (N_2298,N_1649,N_1021);
nand U2299 (N_2299,N_1504,N_1118);
xnor U2300 (N_2300,N_1650,N_1849);
nand U2301 (N_2301,N_1618,N_1898);
nand U2302 (N_2302,N_1906,N_1861);
xor U2303 (N_2303,N_1372,N_1803);
nand U2304 (N_2304,N_1055,N_1331);
and U2305 (N_2305,N_1530,N_1799);
xnor U2306 (N_2306,N_1370,N_1226);
nor U2307 (N_2307,N_1159,N_1977);
nand U2308 (N_2308,N_1054,N_1324);
or U2309 (N_2309,N_1762,N_1800);
xnor U2310 (N_2310,N_1615,N_1752);
xor U2311 (N_2311,N_1345,N_1669);
nand U2312 (N_2312,N_1373,N_1678);
nand U2313 (N_2313,N_1997,N_1489);
or U2314 (N_2314,N_1569,N_1103);
xnor U2315 (N_2315,N_1326,N_1059);
or U2316 (N_2316,N_1087,N_1815);
nand U2317 (N_2317,N_1718,N_1492);
or U2318 (N_2318,N_1444,N_1867);
nand U2319 (N_2319,N_1924,N_1750);
and U2320 (N_2320,N_1819,N_1976);
and U2321 (N_2321,N_1062,N_1829);
xor U2322 (N_2322,N_1344,N_1467);
or U2323 (N_2323,N_1046,N_1709);
xnor U2324 (N_2324,N_1895,N_1781);
nand U2325 (N_2325,N_1135,N_1722);
xnor U2326 (N_2326,N_1173,N_1167);
nand U2327 (N_2327,N_1101,N_1198);
nor U2328 (N_2328,N_1631,N_1626);
and U2329 (N_2329,N_1271,N_1876);
nand U2330 (N_2330,N_1676,N_1967);
nand U2331 (N_2331,N_1850,N_1119);
nor U2332 (N_2332,N_1897,N_1422);
nand U2333 (N_2333,N_1132,N_1311);
nor U2334 (N_2334,N_1913,N_1827);
or U2335 (N_2335,N_1169,N_1180);
xor U2336 (N_2336,N_1545,N_1184);
nand U2337 (N_2337,N_1925,N_1464);
nor U2338 (N_2338,N_1150,N_1835);
nor U2339 (N_2339,N_1197,N_1098);
nor U2340 (N_2340,N_1237,N_1289);
nor U2341 (N_2341,N_1642,N_1375);
and U2342 (N_2342,N_1458,N_1774);
and U2343 (N_2343,N_1818,N_1949);
or U2344 (N_2344,N_1329,N_1335);
nor U2345 (N_2345,N_1926,N_1332);
nand U2346 (N_2346,N_1786,N_1595);
and U2347 (N_2347,N_1784,N_1105);
nand U2348 (N_2348,N_1086,N_1526);
xor U2349 (N_2349,N_1871,N_1568);
and U2350 (N_2350,N_1593,N_1243);
xor U2351 (N_2351,N_1841,N_1619);
or U2352 (N_2352,N_1529,N_1072);
nor U2353 (N_2353,N_1608,N_1235);
nor U2354 (N_2354,N_1429,N_1644);
xor U2355 (N_2355,N_1737,N_1817);
nand U2356 (N_2356,N_1305,N_1238);
nor U2357 (N_2357,N_1735,N_1115);
and U2358 (N_2358,N_1468,N_1749);
and U2359 (N_2359,N_1223,N_1685);
or U2360 (N_2360,N_1666,N_1454);
nand U2361 (N_2361,N_1431,N_1795);
xor U2362 (N_2362,N_1183,N_1104);
or U2363 (N_2363,N_1577,N_1755);
nand U2364 (N_2364,N_1339,N_1544);
xor U2365 (N_2365,N_1899,N_1081);
nand U2366 (N_2366,N_1124,N_1404);
xor U2367 (N_2367,N_1074,N_1999);
and U2368 (N_2368,N_1182,N_1736);
or U2369 (N_2369,N_1962,N_1121);
nand U2370 (N_2370,N_1946,N_1961);
or U2371 (N_2371,N_1525,N_1417);
xnor U2372 (N_2372,N_1449,N_1359);
nand U2373 (N_2373,N_1598,N_1610);
nand U2374 (N_2374,N_1403,N_1244);
nor U2375 (N_2375,N_1617,N_1287);
and U2376 (N_2376,N_1606,N_1192);
nor U2377 (N_2377,N_1808,N_1787);
xor U2378 (N_2378,N_1448,N_1576);
nor U2379 (N_2379,N_1064,N_1856);
and U2380 (N_2380,N_1963,N_1032);
and U2381 (N_2381,N_1066,N_1082);
xnor U2382 (N_2382,N_1919,N_1934);
xor U2383 (N_2383,N_1907,N_1123);
and U2384 (N_2384,N_1689,N_1270);
and U2385 (N_2385,N_1982,N_1260);
or U2386 (N_2386,N_1172,N_1855);
nor U2387 (N_2387,N_1249,N_1364);
or U2388 (N_2388,N_1029,N_1494);
nor U2389 (N_2389,N_1088,N_1063);
nor U2390 (N_2390,N_1384,N_1410);
xor U2391 (N_2391,N_1938,N_1643);
or U2392 (N_2392,N_1445,N_1859);
nor U2393 (N_2393,N_1532,N_1929);
nor U2394 (N_2394,N_1204,N_1385);
nand U2395 (N_2395,N_1699,N_1034);
or U2396 (N_2396,N_1507,N_1549);
nand U2397 (N_2397,N_1281,N_1482);
or U2398 (N_2398,N_1056,N_1565);
nor U2399 (N_2399,N_1659,N_1075);
and U2400 (N_2400,N_1405,N_1574);
or U2401 (N_2401,N_1259,N_1476);
xnor U2402 (N_2402,N_1753,N_1740);
and U2403 (N_2403,N_1328,N_1112);
xor U2404 (N_2404,N_1131,N_1757);
nor U2405 (N_2405,N_1245,N_1691);
xor U2406 (N_2406,N_1330,N_1168);
and U2407 (N_2407,N_1232,N_1363);
xnor U2408 (N_2408,N_1681,N_1348);
xnor U2409 (N_2409,N_1838,N_1951);
nor U2410 (N_2410,N_1231,N_1390);
and U2411 (N_2411,N_1140,N_1662);
nand U2412 (N_2412,N_1518,N_1488);
xor U2413 (N_2413,N_1318,N_1288);
xnor U2414 (N_2414,N_1416,N_1207);
xnor U2415 (N_2415,N_1213,N_1743);
xnor U2416 (N_2416,N_1155,N_1671);
nor U2417 (N_2417,N_1003,N_1698);
xnor U2418 (N_2418,N_1211,N_1220);
and U2419 (N_2419,N_1252,N_1254);
xor U2420 (N_2420,N_1520,N_1843);
and U2421 (N_2421,N_1564,N_1751);
nand U2422 (N_2422,N_1639,N_1008);
or U2423 (N_2423,N_1845,N_1110);
nand U2424 (N_2424,N_1376,N_1957);
nand U2425 (N_2425,N_1312,N_1636);
xor U2426 (N_2426,N_1142,N_1423);
nand U2427 (N_2427,N_1990,N_1439);
and U2428 (N_2428,N_1275,N_1603);
or U2429 (N_2429,N_1600,N_1257);
nand U2430 (N_2430,N_1853,N_1084);
nand U2431 (N_2431,N_1484,N_1645);
nor U2432 (N_2432,N_1070,N_1051);
and U2433 (N_2433,N_1442,N_1812);
nor U2434 (N_2434,N_1465,N_1893);
and U2435 (N_2435,N_1358,N_1327);
nor U2436 (N_2436,N_1460,N_1240);
nor U2437 (N_2437,N_1354,N_1447);
xor U2438 (N_2438,N_1277,N_1773);
xnor U2439 (N_2439,N_1109,N_1768);
and U2440 (N_2440,N_1690,N_1028);
xnor U2441 (N_2441,N_1922,N_1955);
nor U2442 (N_2442,N_1714,N_1663);
and U2443 (N_2443,N_1038,N_1303);
nand U2444 (N_2444,N_1272,N_1724);
or U2445 (N_2445,N_1002,N_1361);
or U2446 (N_2446,N_1065,N_1000);
and U2447 (N_2447,N_1007,N_1090);
nor U2448 (N_2448,N_1163,N_1160);
xnor U2449 (N_2449,N_1519,N_1660);
and U2450 (N_2450,N_1777,N_1129);
or U2451 (N_2451,N_1546,N_1369);
and U2452 (N_2452,N_1847,N_1199);
nand U2453 (N_2453,N_1916,N_1263);
nor U2454 (N_2454,N_1553,N_1939);
nor U2455 (N_2455,N_1579,N_1575);
and U2456 (N_2456,N_1702,N_1677);
nor U2457 (N_2457,N_1901,N_1443);
xor U2458 (N_2458,N_1314,N_1307);
xor U2459 (N_2459,N_1414,N_1333);
or U2460 (N_2460,N_1067,N_1221);
and U2461 (N_2461,N_1589,N_1486);
or U2462 (N_2462,N_1830,N_1903);
and U2463 (N_2463,N_1502,N_1134);
or U2464 (N_2464,N_1858,N_1804);
xor U2465 (N_2465,N_1424,N_1146);
and U2466 (N_2466,N_1100,N_1388);
xnor U2467 (N_2467,N_1280,N_1175);
nor U2468 (N_2468,N_1108,N_1651);
or U2469 (N_2469,N_1234,N_1304);
nor U2470 (N_2470,N_1141,N_1852);
or U2471 (N_2471,N_1058,N_1542);
nand U2472 (N_2472,N_1832,N_1222);
or U2473 (N_2473,N_1039,N_1570);
nand U2474 (N_2474,N_1763,N_1947);
or U2475 (N_2475,N_1933,N_1701);
nor U2476 (N_2476,N_1834,N_1158);
xnor U2477 (N_2477,N_1374,N_1148);
nand U2478 (N_2478,N_1571,N_1045);
nand U2479 (N_2479,N_1265,N_1745);
xor U2480 (N_2480,N_1557,N_1323);
xnor U2481 (N_2481,N_1262,N_1914);
and U2482 (N_2482,N_1138,N_1591);
or U2483 (N_2483,N_1648,N_1080);
xnor U2484 (N_2484,N_1779,N_1958);
nand U2485 (N_2485,N_1434,N_1154);
nand U2486 (N_2486,N_1637,N_1503);
nor U2487 (N_2487,N_1904,N_1506);
nor U2488 (N_2488,N_1040,N_1156);
nand U2489 (N_2489,N_1860,N_1686);
xor U2490 (N_2490,N_1292,N_1250);
or U2491 (N_2491,N_1261,N_1862);
xor U2492 (N_2492,N_1334,N_1013);
and U2493 (N_2493,N_1622,N_1004);
nor U2494 (N_2494,N_1567,N_1921);
nor U2495 (N_2495,N_1479,N_1092);
and U2496 (N_2496,N_1594,N_1430);
nor U2497 (N_2497,N_1085,N_1219);
or U2498 (N_2498,N_1597,N_1562);
nand U2499 (N_2499,N_1966,N_1875);
nor U2500 (N_2500,N_1257,N_1501);
nand U2501 (N_2501,N_1931,N_1161);
nor U2502 (N_2502,N_1179,N_1984);
nand U2503 (N_2503,N_1127,N_1970);
or U2504 (N_2504,N_1160,N_1058);
xnor U2505 (N_2505,N_1942,N_1105);
nor U2506 (N_2506,N_1442,N_1508);
or U2507 (N_2507,N_1835,N_1645);
nand U2508 (N_2508,N_1324,N_1920);
nor U2509 (N_2509,N_1245,N_1952);
or U2510 (N_2510,N_1299,N_1587);
nor U2511 (N_2511,N_1688,N_1351);
and U2512 (N_2512,N_1439,N_1039);
or U2513 (N_2513,N_1502,N_1852);
and U2514 (N_2514,N_1508,N_1388);
and U2515 (N_2515,N_1429,N_1919);
nand U2516 (N_2516,N_1660,N_1112);
nand U2517 (N_2517,N_1419,N_1036);
xnor U2518 (N_2518,N_1393,N_1640);
nor U2519 (N_2519,N_1876,N_1663);
or U2520 (N_2520,N_1597,N_1930);
xor U2521 (N_2521,N_1208,N_1095);
nand U2522 (N_2522,N_1603,N_1605);
or U2523 (N_2523,N_1088,N_1722);
nand U2524 (N_2524,N_1401,N_1779);
nand U2525 (N_2525,N_1211,N_1520);
nor U2526 (N_2526,N_1165,N_1569);
and U2527 (N_2527,N_1176,N_1085);
xor U2528 (N_2528,N_1720,N_1788);
and U2529 (N_2529,N_1432,N_1024);
or U2530 (N_2530,N_1025,N_1520);
or U2531 (N_2531,N_1469,N_1679);
nor U2532 (N_2532,N_1774,N_1740);
and U2533 (N_2533,N_1269,N_1258);
nand U2534 (N_2534,N_1063,N_1023);
xnor U2535 (N_2535,N_1781,N_1809);
and U2536 (N_2536,N_1435,N_1060);
and U2537 (N_2537,N_1879,N_1063);
xnor U2538 (N_2538,N_1559,N_1812);
and U2539 (N_2539,N_1771,N_1499);
and U2540 (N_2540,N_1506,N_1954);
nor U2541 (N_2541,N_1356,N_1310);
or U2542 (N_2542,N_1298,N_1354);
xnor U2543 (N_2543,N_1733,N_1789);
xor U2544 (N_2544,N_1726,N_1757);
or U2545 (N_2545,N_1947,N_1933);
or U2546 (N_2546,N_1595,N_1063);
or U2547 (N_2547,N_1070,N_1047);
or U2548 (N_2548,N_1768,N_1120);
or U2549 (N_2549,N_1441,N_1980);
and U2550 (N_2550,N_1302,N_1640);
nand U2551 (N_2551,N_1638,N_1893);
nand U2552 (N_2552,N_1243,N_1358);
nand U2553 (N_2553,N_1768,N_1444);
nand U2554 (N_2554,N_1295,N_1787);
and U2555 (N_2555,N_1241,N_1102);
or U2556 (N_2556,N_1467,N_1120);
or U2557 (N_2557,N_1909,N_1677);
nand U2558 (N_2558,N_1602,N_1733);
nand U2559 (N_2559,N_1368,N_1112);
xor U2560 (N_2560,N_1861,N_1490);
xnor U2561 (N_2561,N_1183,N_1835);
and U2562 (N_2562,N_1983,N_1563);
nor U2563 (N_2563,N_1199,N_1696);
nor U2564 (N_2564,N_1936,N_1850);
xor U2565 (N_2565,N_1395,N_1129);
xnor U2566 (N_2566,N_1778,N_1170);
nor U2567 (N_2567,N_1362,N_1610);
or U2568 (N_2568,N_1642,N_1362);
or U2569 (N_2569,N_1884,N_1366);
and U2570 (N_2570,N_1525,N_1773);
or U2571 (N_2571,N_1629,N_1410);
nand U2572 (N_2572,N_1283,N_1670);
or U2573 (N_2573,N_1313,N_1048);
and U2574 (N_2574,N_1850,N_1175);
xnor U2575 (N_2575,N_1857,N_1197);
xor U2576 (N_2576,N_1226,N_1321);
or U2577 (N_2577,N_1775,N_1565);
and U2578 (N_2578,N_1584,N_1811);
nand U2579 (N_2579,N_1454,N_1562);
and U2580 (N_2580,N_1202,N_1510);
and U2581 (N_2581,N_1761,N_1349);
nor U2582 (N_2582,N_1363,N_1333);
xnor U2583 (N_2583,N_1475,N_1161);
xor U2584 (N_2584,N_1187,N_1983);
xor U2585 (N_2585,N_1905,N_1798);
nor U2586 (N_2586,N_1180,N_1555);
and U2587 (N_2587,N_1611,N_1735);
xor U2588 (N_2588,N_1533,N_1987);
or U2589 (N_2589,N_1905,N_1840);
and U2590 (N_2590,N_1107,N_1609);
and U2591 (N_2591,N_1922,N_1196);
xor U2592 (N_2592,N_1762,N_1051);
and U2593 (N_2593,N_1411,N_1678);
or U2594 (N_2594,N_1713,N_1534);
nand U2595 (N_2595,N_1682,N_1932);
nand U2596 (N_2596,N_1557,N_1408);
nor U2597 (N_2597,N_1101,N_1250);
and U2598 (N_2598,N_1026,N_1363);
nor U2599 (N_2599,N_1186,N_1827);
nor U2600 (N_2600,N_1041,N_1846);
xor U2601 (N_2601,N_1117,N_1223);
nand U2602 (N_2602,N_1658,N_1480);
xor U2603 (N_2603,N_1215,N_1894);
nor U2604 (N_2604,N_1603,N_1840);
nor U2605 (N_2605,N_1278,N_1551);
nand U2606 (N_2606,N_1159,N_1183);
nor U2607 (N_2607,N_1082,N_1764);
and U2608 (N_2608,N_1114,N_1350);
and U2609 (N_2609,N_1545,N_1179);
xnor U2610 (N_2610,N_1778,N_1076);
nand U2611 (N_2611,N_1732,N_1972);
nand U2612 (N_2612,N_1486,N_1111);
xor U2613 (N_2613,N_1636,N_1457);
nand U2614 (N_2614,N_1266,N_1872);
nand U2615 (N_2615,N_1635,N_1987);
nor U2616 (N_2616,N_1995,N_1422);
or U2617 (N_2617,N_1172,N_1709);
or U2618 (N_2618,N_1500,N_1969);
nor U2619 (N_2619,N_1528,N_1439);
nand U2620 (N_2620,N_1470,N_1837);
xor U2621 (N_2621,N_1797,N_1705);
or U2622 (N_2622,N_1744,N_1266);
nor U2623 (N_2623,N_1638,N_1324);
nor U2624 (N_2624,N_1163,N_1583);
nand U2625 (N_2625,N_1326,N_1764);
or U2626 (N_2626,N_1490,N_1143);
nand U2627 (N_2627,N_1885,N_1368);
nand U2628 (N_2628,N_1783,N_1591);
nand U2629 (N_2629,N_1226,N_1150);
or U2630 (N_2630,N_1464,N_1640);
xnor U2631 (N_2631,N_1976,N_1001);
nor U2632 (N_2632,N_1925,N_1983);
xnor U2633 (N_2633,N_1752,N_1850);
nand U2634 (N_2634,N_1156,N_1384);
or U2635 (N_2635,N_1330,N_1107);
nand U2636 (N_2636,N_1678,N_1287);
nor U2637 (N_2637,N_1955,N_1298);
or U2638 (N_2638,N_1404,N_1853);
or U2639 (N_2639,N_1881,N_1278);
xor U2640 (N_2640,N_1032,N_1057);
nor U2641 (N_2641,N_1824,N_1463);
nand U2642 (N_2642,N_1175,N_1069);
or U2643 (N_2643,N_1256,N_1977);
nand U2644 (N_2644,N_1265,N_1895);
or U2645 (N_2645,N_1889,N_1004);
nand U2646 (N_2646,N_1902,N_1750);
nor U2647 (N_2647,N_1418,N_1930);
nor U2648 (N_2648,N_1287,N_1494);
and U2649 (N_2649,N_1819,N_1828);
or U2650 (N_2650,N_1325,N_1569);
nand U2651 (N_2651,N_1314,N_1813);
xor U2652 (N_2652,N_1397,N_1192);
nand U2653 (N_2653,N_1406,N_1097);
nand U2654 (N_2654,N_1130,N_1670);
or U2655 (N_2655,N_1962,N_1719);
or U2656 (N_2656,N_1774,N_1257);
nor U2657 (N_2657,N_1524,N_1413);
nor U2658 (N_2658,N_1642,N_1856);
or U2659 (N_2659,N_1249,N_1589);
nand U2660 (N_2660,N_1178,N_1497);
or U2661 (N_2661,N_1236,N_1763);
or U2662 (N_2662,N_1200,N_1143);
or U2663 (N_2663,N_1337,N_1529);
or U2664 (N_2664,N_1414,N_1800);
or U2665 (N_2665,N_1545,N_1618);
and U2666 (N_2666,N_1167,N_1937);
xor U2667 (N_2667,N_1329,N_1133);
and U2668 (N_2668,N_1108,N_1800);
and U2669 (N_2669,N_1505,N_1280);
or U2670 (N_2670,N_1686,N_1112);
nand U2671 (N_2671,N_1133,N_1813);
or U2672 (N_2672,N_1191,N_1149);
or U2673 (N_2673,N_1018,N_1804);
nor U2674 (N_2674,N_1079,N_1389);
xor U2675 (N_2675,N_1938,N_1400);
and U2676 (N_2676,N_1835,N_1416);
xor U2677 (N_2677,N_1348,N_1749);
and U2678 (N_2678,N_1742,N_1101);
or U2679 (N_2679,N_1616,N_1838);
or U2680 (N_2680,N_1825,N_1394);
nor U2681 (N_2681,N_1058,N_1177);
xor U2682 (N_2682,N_1372,N_1014);
nor U2683 (N_2683,N_1907,N_1771);
and U2684 (N_2684,N_1445,N_1636);
and U2685 (N_2685,N_1231,N_1540);
xor U2686 (N_2686,N_1481,N_1755);
nor U2687 (N_2687,N_1964,N_1138);
xor U2688 (N_2688,N_1461,N_1562);
xor U2689 (N_2689,N_1381,N_1055);
and U2690 (N_2690,N_1245,N_1128);
and U2691 (N_2691,N_1772,N_1703);
or U2692 (N_2692,N_1085,N_1808);
nor U2693 (N_2693,N_1440,N_1893);
nor U2694 (N_2694,N_1782,N_1639);
nand U2695 (N_2695,N_1434,N_1371);
nand U2696 (N_2696,N_1098,N_1779);
or U2697 (N_2697,N_1269,N_1219);
and U2698 (N_2698,N_1949,N_1483);
nand U2699 (N_2699,N_1665,N_1413);
nand U2700 (N_2700,N_1396,N_1862);
nor U2701 (N_2701,N_1048,N_1055);
xor U2702 (N_2702,N_1904,N_1173);
nand U2703 (N_2703,N_1470,N_1734);
xnor U2704 (N_2704,N_1400,N_1098);
and U2705 (N_2705,N_1098,N_1888);
and U2706 (N_2706,N_1856,N_1494);
nand U2707 (N_2707,N_1997,N_1425);
nor U2708 (N_2708,N_1734,N_1828);
nor U2709 (N_2709,N_1512,N_1801);
nand U2710 (N_2710,N_1621,N_1487);
nand U2711 (N_2711,N_1332,N_1598);
or U2712 (N_2712,N_1431,N_1695);
or U2713 (N_2713,N_1470,N_1181);
nand U2714 (N_2714,N_1719,N_1825);
or U2715 (N_2715,N_1228,N_1827);
or U2716 (N_2716,N_1447,N_1570);
xnor U2717 (N_2717,N_1424,N_1400);
nor U2718 (N_2718,N_1208,N_1690);
or U2719 (N_2719,N_1564,N_1735);
xor U2720 (N_2720,N_1077,N_1528);
or U2721 (N_2721,N_1755,N_1705);
and U2722 (N_2722,N_1083,N_1171);
and U2723 (N_2723,N_1945,N_1032);
and U2724 (N_2724,N_1921,N_1128);
xor U2725 (N_2725,N_1806,N_1245);
nand U2726 (N_2726,N_1454,N_1638);
nand U2727 (N_2727,N_1603,N_1215);
or U2728 (N_2728,N_1614,N_1486);
nand U2729 (N_2729,N_1131,N_1280);
nand U2730 (N_2730,N_1266,N_1118);
or U2731 (N_2731,N_1120,N_1492);
or U2732 (N_2732,N_1667,N_1391);
xnor U2733 (N_2733,N_1390,N_1930);
or U2734 (N_2734,N_1229,N_1628);
and U2735 (N_2735,N_1119,N_1244);
xnor U2736 (N_2736,N_1926,N_1910);
nand U2737 (N_2737,N_1538,N_1606);
nor U2738 (N_2738,N_1429,N_1545);
xnor U2739 (N_2739,N_1513,N_1023);
xnor U2740 (N_2740,N_1797,N_1823);
xor U2741 (N_2741,N_1676,N_1437);
nor U2742 (N_2742,N_1233,N_1663);
nor U2743 (N_2743,N_1174,N_1747);
and U2744 (N_2744,N_1759,N_1724);
nand U2745 (N_2745,N_1110,N_1505);
nor U2746 (N_2746,N_1734,N_1820);
nand U2747 (N_2747,N_1786,N_1697);
xor U2748 (N_2748,N_1492,N_1504);
and U2749 (N_2749,N_1946,N_1545);
or U2750 (N_2750,N_1085,N_1138);
or U2751 (N_2751,N_1249,N_1374);
and U2752 (N_2752,N_1094,N_1572);
nor U2753 (N_2753,N_1895,N_1434);
or U2754 (N_2754,N_1160,N_1452);
xnor U2755 (N_2755,N_1640,N_1241);
xnor U2756 (N_2756,N_1280,N_1830);
and U2757 (N_2757,N_1936,N_1743);
nor U2758 (N_2758,N_1039,N_1213);
and U2759 (N_2759,N_1638,N_1222);
xor U2760 (N_2760,N_1406,N_1673);
xor U2761 (N_2761,N_1538,N_1278);
and U2762 (N_2762,N_1926,N_1182);
and U2763 (N_2763,N_1622,N_1445);
or U2764 (N_2764,N_1547,N_1326);
nand U2765 (N_2765,N_1820,N_1495);
and U2766 (N_2766,N_1539,N_1203);
or U2767 (N_2767,N_1646,N_1817);
and U2768 (N_2768,N_1829,N_1005);
or U2769 (N_2769,N_1138,N_1108);
nor U2770 (N_2770,N_1489,N_1993);
xor U2771 (N_2771,N_1969,N_1668);
and U2772 (N_2772,N_1938,N_1536);
nor U2773 (N_2773,N_1303,N_1142);
and U2774 (N_2774,N_1046,N_1467);
nor U2775 (N_2775,N_1230,N_1994);
nor U2776 (N_2776,N_1229,N_1515);
and U2777 (N_2777,N_1371,N_1013);
nor U2778 (N_2778,N_1949,N_1573);
or U2779 (N_2779,N_1821,N_1955);
nor U2780 (N_2780,N_1780,N_1477);
nor U2781 (N_2781,N_1769,N_1216);
and U2782 (N_2782,N_1355,N_1098);
xor U2783 (N_2783,N_1704,N_1595);
or U2784 (N_2784,N_1454,N_1588);
xor U2785 (N_2785,N_1454,N_1462);
xor U2786 (N_2786,N_1055,N_1454);
nand U2787 (N_2787,N_1860,N_1088);
xor U2788 (N_2788,N_1113,N_1865);
and U2789 (N_2789,N_1541,N_1607);
xnor U2790 (N_2790,N_1777,N_1169);
or U2791 (N_2791,N_1765,N_1130);
or U2792 (N_2792,N_1094,N_1177);
nor U2793 (N_2793,N_1546,N_1041);
or U2794 (N_2794,N_1580,N_1854);
nand U2795 (N_2795,N_1044,N_1049);
xnor U2796 (N_2796,N_1620,N_1021);
nand U2797 (N_2797,N_1044,N_1633);
and U2798 (N_2798,N_1120,N_1907);
nor U2799 (N_2799,N_1446,N_1625);
or U2800 (N_2800,N_1391,N_1479);
nor U2801 (N_2801,N_1493,N_1403);
nand U2802 (N_2802,N_1293,N_1078);
nand U2803 (N_2803,N_1340,N_1652);
or U2804 (N_2804,N_1284,N_1311);
nand U2805 (N_2805,N_1697,N_1982);
nand U2806 (N_2806,N_1970,N_1164);
and U2807 (N_2807,N_1210,N_1602);
and U2808 (N_2808,N_1603,N_1897);
xor U2809 (N_2809,N_1003,N_1084);
nand U2810 (N_2810,N_1443,N_1940);
and U2811 (N_2811,N_1231,N_1226);
or U2812 (N_2812,N_1078,N_1977);
and U2813 (N_2813,N_1488,N_1132);
nor U2814 (N_2814,N_1365,N_1011);
nor U2815 (N_2815,N_1916,N_1249);
nand U2816 (N_2816,N_1261,N_1798);
or U2817 (N_2817,N_1368,N_1638);
xor U2818 (N_2818,N_1457,N_1209);
or U2819 (N_2819,N_1360,N_1900);
nand U2820 (N_2820,N_1743,N_1712);
and U2821 (N_2821,N_1072,N_1836);
nor U2822 (N_2822,N_1709,N_1603);
nand U2823 (N_2823,N_1796,N_1844);
xnor U2824 (N_2824,N_1904,N_1684);
xnor U2825 (N_2825,N_1417,N_1597);
xor U2826 (N_2826,N_1251,N_1870);
or U2827 (N_2827,N_1375,N_1784);
or U2828 (N_2828,N_1356,N_1023);
nand U2829 (N_2829,N_1926,N_1945);
nor U2830 (N_2830,N_1877,N_1397);
nand U2831 (N_2831,N_1814,N_1027);
or U2832 (N_2832,N_1585,N_1123);
or U2833 (N_2833,N_1541,N_1255);
xnor U2834 (N_2834,N_1098,N_1272);
xnor U2835 (N_2835,N_1023,N_1691);
and U2836 (N_2836,N_1676,N_1290);
and U2837 (N_2837,N_1149,N_1984);
and U2838 (N_2838,N_1879,N_1003);
or U2839 (N_2839,N_1956,N_1864);
or U2840 (N_2840,N_1519,N_1310);
nand U2841 (N_2841,N_1048,N_1395);
nor U2842 (N_2842,N_1460,N_1054);
or U2843 (N_2843,N_1955,N_1711);
and U2844 (N_2844,N_1164,N_1057);
nand U2845 (N_2845,N_1418,N_1900);
nor U2846 (N_2846,N_1428,N_1845);
nor U2847 (N_2847,N_1299,N_1598);
xnor U2848 (N_2848,N_1252,N_1174);
and U2849 (N_2849,N_1929,N_1753);
nand U2850 (N_2850,N_1560,N_1443);
xnor U2851 (N_2851,N_1497,N_1456);
xnor U2852 (N_2852,N_1909,N_1903);
nand U2853 (N_2853,N_1311,N_1714);
nand U2854 (N_2854,N_1347,N_1237);
nor U2855 (N_2855,N_1342,N_1905);
xnor U2856 (N_2856,N_1637,N_1416);
nand U2857 (N_2857,N_1302,N_1051);
nand U2858 (N_2858,N_1809,N_1421);
nor U2859 (N_2859,N_1832,N_1247);
and U2860 (N_2860,N_1462,N_1800);
and U2861 (N_2861,N_1215,N_1829);
or U2862 (N_2862,N_1839,N_1009);
nor U2863 (N_2863,N_1614,N_1315);
and U2864 (N_2864,N_1662,N_1834);
or U2865 (N_2865,N_1417,N_1586);
nand U2866 (N_2866,N_1246,N_1203);
nor U2867 (N_2867,N_1718,N_1137);
xor U2868 (N_2868,N_1311,N_1361);
nor U2869 (N_2869,N_1148,N_1396);
xnor U2870 (N_2870,N_1212,N_1346);
and U2871 (N_2871,N_1578,N_1781);
and U2872 (N_2872,N_1032,N_1144);
nand U2873 (N_2873,N_1307,N_1209);
or U2874 (N_2874,N_1306,N_1789);
or U2875 (N_2875,N_1853,N_1596);
and U2876 (N_2876,N_1298,N_1433);
nand U2877 (N_2877,N_1715,N_1336);
xor U2878 (N_2878,N_1867,N_1213);
or U2879 (N_2879,N_1399,N_1529);
or U2880 (N_2880,N_1258,N_1442);
and U2881 (N_2881,N_1984,N_1913);
and U2882 (N_2882,N_1326,N_1563);
nand U2883 (N_2883,N_1249,N_1529);
and U2884 (N_2884,N_1584,N_1451);
nand U2885 (N_2885,N_1673,N_1401);
xnor U2886 (N_2886,N_1690,N_1191);
nand U2887 (N_2887,N_1899,N_1890);
and U2888 (N_2888,N_1392,N_1531);
and U2889 (N_2889,N_1372,N_1025);
xnor U2890 (N_2890,N_1844,N_1806);
or U2891 (N_2891,N_1272,N_1083);
nand U2892 (N_2892,N_1902,N_1017);
or U2893 (N_2893,N_1146,N_1467);
xnor U2894 (N_2894,N_1712,N_1479);
or U2895 (N_2895,N_1817,N_1148);
or U2896 (N_2896,N_1730,N_1760);
or U2897 (N_2897,N_1485,N_1882);
or U2898 (N_2898,N_1169,N_1365);
nor U2899 (N_2899,N_1389,N_1518);
xnor U2900 (N_2900,N_1853,N_1784);
nor U2901 (N_2901,N_1429,N_1605);
or U2902 (N_2902,N_1449,N_1374);
xnor U2903 (N_2903,N_1556,N_1071);
xor U2904 (N_2904,N_1821,N_1517);
xor U2905 (N_2905,N_1206,N_1682);
nor U2906 (N_2906,N_1065,N_1976);
xnor U2907 (N_2907,N_1519,N_1960);
or U2908 (N_2908,N_1000,N_1390);
xnor U2909 (N_2909,N_1526,N_1262);
nand U2910 (N_2910,N_1451,N_1201);
xor U2911 (N_2911,N_1640,N_1113);
xor U2912 (N_2912,N_1829,N_1922);
or U2913 (N_2913,N_1180,N_1260);
xor U2914 (N_2914,N_1726,N_1072);
nor U2915 (N_2915,N_1163,N_1314);
or U2916 (N_2916,N_1430,N_1498);
or U2917 (N_2917,N_1497,N_1270);
nor U2918 (N_2918,N_1298,N_1898);
nand U2919 (N_2919,N_1105,N_1353);
nand U2920 (N_2920,N_1099,N_1487);
nand U2921 (N_2921,N_1540,N_1485);
xnor U2922 (N_2922,N_1467,N_1646);
nor U2923 (N_2923,N_1503,N_1521);
xnor U2924 (N_2924,N_1466,N_1293);
nor U2925 (N_2925,N_1745,N_1746);
xor U2926 (N_2926,N_1041,N_1732);
nor U2927 (N_2927,N_1863,N_1872);
nor U2928 (N_2928,N_1029,N_1922);
xnor U2929 (N_2929,N_1619,N_1673);
nand U2930 (N_2930,N_1931,N_1889);
and U2931 (N_2931,N_1867,N_1211);
nand U2932 (N_2932,N_1324,N_1567);
nor U2933 (N_2933,N_1045,N_1042);
or U2934 (N_2934,N_1126,N_1012);
and U2935 (N_2935,N_1908,N_1657);
nor U2936 (N_2936,N_1875,N_1776);
or U2937 (N_2937,N_1643,N_1039);
xnor U2938 (N_2938,N_1702,N_1772);
or U2939 (N_2939,N_1905,N_1812);
and U2940 (N_2940,N_1955,N_1365);
and U2941 (N_2941,N_1312,N_1331);
xor U2942 (N_2942,N_1787,N_1661);
or U2943 (N_2943,N_1140,N_1984);
nand U2944 (N_2944,N_1318,N_1778);
nor U2945 (N_2945,N_1722,N_1575);
and U2946 (N_2946,N_1447,N_1567);
xor U2947 (N_2947,N_1053,N_1320);
and U2948 (N_2948,N_1012,N_1348);
and U2949 (N_2949,N_1030,N_1431);
xor U2950 (N_2950,N_1151,N_1793);
and U2951 (N_2951,N_1780,N_1656);
or U2952 (N_2952,N_1565,N_1686);
or U2953 (N_2953,N_1489,N_1498);
xnor U2954 (N_2954,N_1424,N_1048);
nor U2955 (N_2955,N_1196,N_1894);
or U2956 (N_2956,N_1225,N_1507);
or U2957 (N_2957,N_1116,N_1594);
or U2958 (N_2958,N_1804,N_1159);
or U2959 (N_2959,N_1009,N_1813);
and U2960 (N_2960,N_1539,N_1435);
nor U2961 (N_2961,N_1634,N_1516);
and U2962 (N_2962,N_1571,N_1754);
nand U2963 (N_2963,N_1627,N_1615);
and U2964 (N_2964,N_1934,N_1338);
and U2965 (N_2965,N_1056,N_1070);
and U2966 (N_2966,N_1653,N_1113);
nand U2967 (N_2967,N_1365,N_1409);
nor U2968 (N_2968,N_1451,N_1963);
or U2969 (N_2969,N_1790,N_1543);
xor U2970 (N_2970,N_1397,N_1972);
nand U2971 (N_2971,N_1412,N_1577);
xor U2972 (N_2972,N_1604,N_1953);
nor U2973 (N_2973,N_1584,N_1383);
nand U2974 (N_2974,N_1945,N_1714);
or U2975 (N_2975,N_1313,N_1451);
nor U2976 (N_2976,N_1733,N_1011);
or U2977 (N_2977,N_1474,N_1600);
and U2978 (N_2978,N_1796,N_1599);
xnor U2979 (N_2979,N_1080,N_1489);
nor U2980 (N_2980,N_1361,N_1066);
and U2981 (N_2981,N_1667,N_1620);
nand U2982 (N_2982,N_1751,N_1935);
xor U2983 (N_2983,N_1816,N_1091);
nand U2984 (N_2984,N_1480,N_1061);
and U2985 (N_2985,N_1144,N_1960);
xnor U2986 (N_2986,N_1861,N_1281);
and U2987 (N_2987,N_1017,N_1030);
nor U2988 (N_2988,N_1739,N_1257);
or U2989 (N_2989,N_1206,N_1015);
and U2990 (N_2990,N_1201,N_1318);
and U2991 (N_2991,N_1302,N_1766);
and U2992 (N_2992,N_1002,N_1892);
nand U2993 (N_2993,N_1407,N_1386);
or U2994 (N_2994,N_1382,N_1432);
nand U2995 (N_2995,N_1229,N_1045);
nand U2996 (N_2996,N_1821,N_1242);
nor U2997 (N_2997,N_1213,N_1615);
xnor U2998 (N_2998,N_1416,N_1780);
xor U2999 (N_2999,N_1494,N_1321);
nor U3000 (N_3000,N_2136,N_2984);
and U3001 (N_3001,N_2525,N_2981);
nand U3002 (N_3002,N_2499,N_2797);
and U3003 (N_3003,N_2833,N_2449);
xnor U3004 (N_3004,N_2998,N_2747);
xnor U3005 (N_3005,N_2221,N_2047);
nand U3006 (N_3006,N_2544,N_2687);
or U3007 (N_3007,N_2300,N_2646);
xor U3008 (N_3008,N_2589,N_2590);
or U3009 (N_3009,N_2764,N_2683);
or U3010 (N_3010,N_2391,N_2636);
xor U3011 (N_3011,N_2814,N_2400);
xor U3012 (N_3012,N_2650,N_2176);
nand U3013 (N_3013,N_2293,N_2407);
or U3014 (N_3014,N_2695,N_2826);
nor U3015 (N_3015,N_2322,N_2754);
xnor U3016 (N_3016,N_2485,N_2691);
nand U3017 (N_3017,N_2884,N_2402);
xnor U3018 (N_3018,N_2375,N_2368);
nor U3019 (N_3019,N_2103,N_2704);
or U3020 (N_3020,N_2570,N_2721);
nor U3021 (N_3021,N_2673,N_2732);
nand U3022 (N_3022,N_2258,N_2278);
or U3023 (N_3023,N_2714,N_2528);
and U3024 (N_3024,N_2305,N_2999);
and U3025 (N_3025,N_2593,N_2444);
nand U3026 (N_3026,N_2017,N_2364);
xor U3027 (N_3027,N_2584,N_2566);
and U3028 (N_3028,N_2263,N_2940);
and U3029 (N_3029,N_2592,N_2643);
xor U3030 (N_3030,N_2203,N_2351);
or U3031 (N_3031,N_2064,N_2283);
nor U3032 (N_3032,N_2083,N_2448);
nor U3033 (N_3033,N_2843,N_2844);
nand U3034 (N_3034,N_2559,N_2717);
and U3035 (N_3035,N_2131,N_2072);
nand U3036 (N_3036,N_2168,N_2730);
or U3037 (N_3037,N_2378,N_2371);
or U3038 (N_3038,N_2688,N_2426);
nand U3039 (N_3039,N_2512,N_2233);
or U3040 (N_3040,N_2430,N_2259);
xnor U3041 (N_3041,N_2978,N_2581);
and U3042 (N_3042,N_2788,N_2343);
xor U3043 (N_3043,N_2308,N_2313);
xnor U3044 (N_3044,N_2824,N_2249);
nor U3045 (N_3045,N_2196,N_2873);
or U3046 (N_3046,N_2200,N_2401);
xnor U3047 (N_3047,N_2778,N_2193);
nand U3048 (N_3048,N_2409,N_2297);
nand U3049 (N_3049,N_2081,N_2447);
xor U3050 (N_3050,N_2519,N_2091);
nand U3051 (N_3051,N_2287,N_2423);
or U3052 (N_3052,N_2654,N_2336);
xnor U3053 (N_3053,N_2145,N_2334);
nor U3054 (N_3054,N_2161,N_2540);
or U3055 (N_3055,N_2063,N_2601);
xor U3056 (N_3056,N_2881,N_2903);
xnor U3057 (N_3057,N_2315,N_2163);
xor U3058 (N_3058,N_2492,N_2491);
nand U3059 (N_3059,N_2149,N_2555);
and U3060 (N_3060,N_2215,N_2619);
and U3061 (N_3061,N_2374,N_2562);
or U3062 (N_3062,N_2803,N_2908);
nor U3063 (N_3063,N_2112,N_2832);
xnor U3064 (N_3064,N_2373,N_2082);
nor U3065 (N_3065,N_2464,N_2338);
xnor U3066 (N_3066,N_2890,N_2395);
xor U3067 (N_3067,N_2777,N_2853);
nor U3068 (N_3068,N_2299,N_2446);
or U3069 (N_3069,N_2527,N_2858);
nor U3070 (N_3070,N_2523,N_2758);
nor U3071 (N_3071,N_2553,N_2694);
xor U3072 (N_3072,N_2950,N_2236);
or U3073 (N_3073,N_2791,N_2298);
and U3074 (N_3074,N_2756,N_2912);
nor U3075 (N_3075,N_2237,N_2275);
xor U3076 (N_3076,N_2554,N_2073);
and U3077 (N_3077,N_2975,N_2307);
nor U3078 (N_3078,N_2075,N_2744);
nand U3079 (N_3079,N_2792,N_2825);
xnor U3080 (N_3080,N_2326,N_2240);
nor U3081 (N_3081,N_2698,N_2970);
or U3082 (N_3082,N_2663,N_2214);
nand U3083 (N_3083,N_2610,N_2247);
and U3084 (N_3084,N_2035,N_2363);
or U3085 (N_3085,N_2757,N_2595);
or U3086 (N_3086,N_2591,N_2750);
xor U3087 (N_3087,N_2751,N_2005);
nor U3088 (N_3088,N_2501,N_2273);
nor U3089 (N_3089,N_2290,N_2040);
nand U3090 (N_3090,N_2996,N_2460);
xor U3091 (N_3091,N_2985,N_2805);
nand U3092 (N_3092,N_2626,N_2294);
xnor U3093 (N_3093,N_2852,N_2867);
xnor U3094 (N_3094,N_2011,N_2733);
and U3095 (N_3095,N_2889,N_2223);
nor U3096 (N_3096,N_2773,N_2494);
xor U3097 (N_3097,N_2945,N_2268);
nor U3098 (N_3098,N_2507,N_2573);
nand U3099 (N_3099,N_2874,N_2379);
nand U3100 (N_3100,N_2851,N_2471);
nand U3101 (N_3101,N_2693,N_2018);
nor U3102 (N_3102,N_2370,N_2349);
or U3103 (N_3103,N_2146,N_2863);
and U3104 (N_3104,N_2551,N_2675);
or U3105 (N_3105,N_2171,N_2250);
or U3106 (N_3106,N_2295,N_2895);
xor U3107 (N_3107,N_2183,N_2766);
and U3108 (N_3108,N_2986,N_2393);
nor U3109 (N_3109,N_2137,N_2353);
nor U3110 (N_3110,N_2265,N_2366);
nand U3111 (N_3111,N_2868,N_2316);
and U3112 (N_3112,N_2925,N_2835);
or U3113 (N_3113,N_2793,N_2222);
nand U3114 (N_3114,N_2154,N_2101);
nor U3115 (N_3115,N_2739,N_2845);
nor U3116 (N_3116,N_2454,N_2212);
nor U3117 (N_3117,N_2964,N_2888);
nand U3118 (N_3118,N_2552,N_2106);
xor U3119 (N_3119,N_2799,N_2779);
nand U3120 (N_3120,N_2417,N_2923);
nand U3121 (N_3121,N_2785,N_2541);
and U3122 (N_3122,N_2685,N_2927);
nor U3123 (N_3123,N_2088,N_2885);
nand U3124 (N_3124,N_2169,N_2569);
xnor U3125 (N_3125,N_2281,N_2919);
nand U3126 (N_3126,N_2804,N_2837);
nor U3127 (N_3127,N_2053,N_2008);
xnor U3128 (N_3128,N_2425,N_2948);
nand U3129 (N_3129,N_2253,N_2229);
xnor U3130 (N_3130,N_2352,N_2831);
or U3131 (N_3131,N_2960,N_2910);
nor U3132 (N_3132,N_2323,N_2410);
and U3133 (N_3133,N_2394,N_2734);
xnor U3134 (N_3134,N_2632,N_2406);
or U3135 (N_3135,N_2979,N_2955);
nand U3136 (N_3136,N_2434,N_2068);
xnor U3137 (N_3137,N_2529,N_2167);
nand U3138 (N_3138,N_2111,N_2576);
xor U3139 (N_3139,N_2561,N_2533);
and U3140 (N_3140,N_2711,N_2360);
nand U3141 (N_3141,N_2272,N_2361);
nand U3142 (N_3142,N_2127,N_2738);
and U3143 (N_3143,N_2857,N_2631);
and U3144 (N_3144,N_2291,N_2049);
or U3145 (N_3145,N_2085,N_2783);
nor U3146 (N_3146,N_2043,N_2669);
xnor U3147 (N_3147,N_2133,N_2204);
xnor U3148 (N_3148,N_2810,N_2725);
nand U3149 (N_3149,N_2860,N_2318);
or U3150 (N_3150,N_2380,N_2396);
nand U3151 (N_3151,N_2642,N_2288);
nor U3152 (N_3152,N_2697,N_2941);
nand U3153 (N_3153,N_2677,N_2344);
nand U3154 (N_3154,N_2197,N_2504);
nor U3155 (N_3155,N_2746,N_2547);
and U3156 (N_3156,N_2787,N_2019);
nand U3157 (N_3157,N_2050,N_2097);
or U3158 (N_3158,N_2206,N_2796);
or U3159 (N_3159,N_2661,N_2102);
nand U3160 (N_3160,N_2522,N_2384);
and U3161 (N_3161,N_2498,N_2871);
or U3162 (N_3162,N_2069,N_2560);
xor U3163 (N_3163,N_2658,N_2245);
or U3164 (N_3164,N_2164,N_2864);
or U3165 (N_3165,N_2440,N_2652);
nand U3166 (N_3166,N_2289,N_2475);
and U3167 (N_3167,N_2722,N_2938);
or U3168 (N_3168,N_2974,N_2473);
nand U3169 (N_3169,N_2060,N_2319);
nand U3170 (N_3170,N_2304,N_2893);
nor U3171 (N_3171,N_2850,N_2474);
or U3172 (N_3172,N_2213,N_2096);
xnor U3173 (N_3173,N_2246,N_2037);
or U3174 (N_3174,N_2546,N_2958);
and U3175 (N_3175,N_2033,N_2909);
xnor U3176 (N_3176,N_2862,N_2261);
or U3177 (N_3177,N_2823,N_2488);
and U3178 (N_3178,N_2680,N_2795);
nand U3179 (N_3179,N_2536,N_2624);
or U3180 (N_3180,N_2579,N_2761);
xnor U3181 (N_3181,N_2119,N_2412);
or U3182 (N_3182,N_2386,N_2630);
nor U3183 (N_3183,N_2269,N_2270);
nor U3184 (N_3184,N_2847,N_2915);
or U3185 (N_3185,N_2226,N_2728);
nor U3186 (N_3186,N_2550,N_2982);
or U3187 (N_3187,N_2752,N_2913);
or U3188 (N_3188,N_2937,N_2790);
xor U3189 (N_3189,N_2633,N_2388);
or U3190 (N_3190,N_2954,N_2645);
nor U3191 (N_3191,N_2710,N_2128);
and U3192 (N_3192,N_2381,N_2936);
and U3193 (N_3193,N_2794,N_2117);
nor U3194 (N_3194,N_2668,N_2230);
or U3195 (N_3195,N_2476,N_2113);
xor U3196 (N_3196,N_2122,N_2216);
xnor U3197 (N_3197,N_2095,N_2114);
xor U3198 (N_3198,N_2684,N_2170);
and U3199 (N_3199,N_2074,N_2178);
xor U3200 (N_3200,N_2849,N_2435);
or U3201 (N_3201,N_2963,N_2179);
nor U3202 (N_3202,N_2048,N_2034);
nor U3203 (N_3203,N_2548,N_2408);
nand U3204 (N_3204,N_2419,N_2439);
and U3205 (N_3205,N_2951,N_2662);
nor U3206 (N_3206,N_2451,N_2359);
xor U3207 (N_3207,N_2962,N_2134);
nand U3208 (N_3208,N_2956,N_2899);
nand U3209 (N_3209,N_2387,N_2003);
nor U3210 (N_3210,N_2883,N_2840);
nor U3211 (N_3211,N_2802,N_2462);
nor U3212 (N_3212,N_2225,N_2558);
nor U3213 (N_3213,N_2357,N_2012);
nand U3214 (N_3214,N_2207,N_2660);
and U3215 (N_3215,N_2953,N_2039);
xnor U3216 (N_3216,N_2526,N_2092);
or U3217 (N_3217,N_2354,N_2991);
nor U3218 (N_3218,N_2534,N_2071);
or U3219 (N_3219,N_2188,N_2789);
and U3220 (N_3220,N_2224,N_2467);
nor U3221 (N_3221,N_2716,N_2665);
or U3222 (N_3222,N_2775,N_2015);
nor U3223 (N_3223,N_2703,N_2967);
nor U3224 (N_3224,N_2699,N_2596);
nor U3225 (N_3225,N_2635,N_2531);
and U3226 (N_3226,N_2321,N_2465);
xnor U3227 (N_3227,N_2132,N_2489);
xor U3228 (N_3228,N_2198,N_2556);
and U3229 (N_3229,N_2199,N_2187);
nand U3230 (N_3230,N_2743,N_2922);
or U3231 (N_3231,N_2126,N_2618);
xnor U3232 (N_3232,N_2513,N_2980);
nor U3233 (N_3233,N_2995,N_2515);
xor U3234 (N_3234,N_2578,N_2543);
xor U3235 (N_3235,N_2463,N_2031);
and U3236 (N_3236,N_2538,N_2820);
nor U3237 (N_3237,N_2238,N_2718);
and U3238 (N_3238,N_2896,N_2104);
xnor U3239 (N_3239,N_2629,N_2495);
or U3240 (N_3240,N_2900,N_2928);
and U3241 (N_3241,N_2876,N_2159);
xnor U3242 (N_3242,N_2377,N_2487);
xnor U3243 (N_3243,N_2009,N_2597);
xor U3244 (N_3244,N_2563,N_2427);
nand U3245 (N_3245,N_2781,N_2234);
xor U3246 (N_3246,N_2369,N_2271);
or U3247 (N_3247,N_2254,N_2907);
or U3248 (N_3248,N_2416,N_2411);
or U3249 (N_3249,N_2517,N_2219);
xor U3250 (N_3250,N_2090,N_2854);
nor U3251 (N_3251,N_2320,N_2706);
nand U3252 (N_3252,N_2723,N_2162);
xnor U3253 (N_3253,N_2218,N_2933);
nand U3254 (N_3254,N_2022,N_2175);
or U3255 (N_3255,N_2046,N_2976);
nor U3256 (N_3256,N_2014,N_2959);
and U3257 (N_3257,N_2277,N_2262);
or U3258 (N_3258,N_2165,N_2839);
and U3259 (N_3259,N_2004,N_2030);
nand U3260 (N_3260,N_2514,N_2902);
or U3261 (N_3261,N_2657,N_2089);
nand U3262 (N_3262,N_2836,N_2413);
and U3263 (N_3263,N_2931,N_2220);
nor U3264 (N_3264,N_2911,N_2943);
or U3265 (N_3265,N_2585,N_2606);
xnor U3266 (N_3266,N_2302,N_2952);
nand U3267 (N_3267,N_2574,N_2510);
or U3268 (N_3268,N_2653,N_2634);
nand U3269 (N_3269,N_2520,N_2385);
or U3270 (N_3270,N_2604,N_2834);
xnor U3271 (N_3271,N_2770,N_2957);
nor U3272 (N_3272,N_2405,N_2006);
and U3273 (N_3273,N_2892,N_2026);
or U3274 (N_3274,N_2382,N_2692);
nor U3275 (N_3275,N_2838,N_2332);
xnor U3276 (N_3276,N_2067,N_2418);
xor U3277 (N_3277,N_2916,N_2649);
nand U3278 (N_3278,N_2568,N_2044);
nand U3279 (N_3279,N_2887,N_2621);
or U3280 (N_3280,N_2516,N_2612);
xor U3281 (N_3281,N_2765,N_2990);
nor U3282 (N_3282,N_2608,N_2174);
nand U3283 (N_3283,N_2740,N_2453);
and U3284 (N_3284,N_2142,N_2749);
xnor U3285 (N_3285,N_2116,N_2763);
nor U3286 (N_3286,N_2086,N_2603);
xor U3287 (N_3287,N_2780,N_2135);
or U3288 (N_3288,N_2392,N_2842);
or U3289 (N_3289,N_2762,N_2054);
and U3290 (N_3290,N_2811,N_2818);
or U3291 (N_3291,N_2333,N_2038);
nor U3292 (N_3292,N_2932,N_2613);
nor U3293 (N_3293,N_2689,N_2041);
or U3294 (N_3294,N_2490,N_2886);
and U3295 (N_3295,N_2007,N_2518);
nand U3296 (N_3296,N_2872,N_2317);
and U3297 (N_3297,N_2231,N_2856);
xnor U3298 (N_3298,N_2865,N_2042);
xnor U3299 (N_3299,N_2674,N_2098);
or U3300 (N_3300,N_2607,N_2355);
nor U3301 (N_3301,N_2808,N_2482);
nor U3302 (N_3302,N_2468,N_2483);
nor U3303 (N_3303,N_2929,N_2028);
xor U3304 (N_3304,N_2094,N_2904);
xor U3305 (N_3305,N_2942,N_2157);
nor U3306 (N_3306,N_2580,N_2422);
xnor U3307 (N_3307,N_2637,N_2855);
or U3308 (N_3308,N_2000,N_2994);
nand U3309 (N_3309,N_2324,N_2949);
nor U3310 (N_3310,N_2755,N_2079);
xor U3311 (N_3311,N_2784,N_2443);
nor U3312 (N_3312,N_2701,N_2917);
nor U3313 (N_3313,N_2737,N_2497);
nor U3314 (N_3314,N_2532,N_2898);
nand U3315 (N_3315,N_2615,N_2372);
and U3316 (N_3316,N_2731,N_2255);
xnor U3317 (N_3317,N_2347,N_2681);
xor U3318 (N_3318,N_2399,N_2753);
nor U3319 (N_3319,N_2726,N_2549);
or U3320 (N_3320,N_2702,N_2539);
and U3321 (N_3321,N_2565,N_2194);
xnor U3322 (N_3322,N_2358,N_2404);
xnor U3323 (N_3323,N_2328,N_2470);
xnor U3324 (N_3324,N_2924,N_2920);
nand U3325 (N_3325,N_2158,N_2878);
and U3326 (N_3326,N_2442,N_2870);
or U3327 (N_3327,N_2227,N_2997);
nand U3328 (N_3328,N_2208,N_2390);
nand U3329 (N_3329,N_2459,N_2506);
or U3330 (N_3330,N_2807,N_2724);
or U3331 (N_3331,N_2496,N_2228);
xnor U3332 (N_3332,N_2020,N_2700);
nand U3333 (N_3333,N_2690,N_2760);
or U3334 (N_3334,N_2666,N_2801);
xnor U3335 (N_3335,N_2016,N_2202);
nor U3336 (N_3336,N_2239,N_2182);
and U3337 (N_3337,N_2582,N_2640);
or U3338 (N_3338,N_2013,N_2616);
or U3339 (N_3339,N_2813,N_2274);
nor U3340 (N_3340,N_2189,N_2500);
nand U3341 (N_3341,N_2123,N_2027);
xnor U3342 (N_3342,N_2947,N_2311);
xor U3343 (N_3343,N_2428,N_2961);
xnor U3344 (N_3344,N_2679,N_2715);
nor U3345 (N_3345,N_2211,N_2664);
nor U3346 (N_3346,N_2882,N_2651);
xnor U3347 (N_3347,N_2583,N_2177);
xor U3348 (N_3348,N_2926,N_2152);
nor U3349 (N_3349,N_2080,N_2441);
nand U3350 (N_3350,N_2209,N_2901);
nand U3351 (N_3351,N_2966,N_2257);
nor U3352 (N_3352,N_2627,N_2348);
nor U3353 (N_3353,N_2798,N_2156);
and U3354 (N_3354,N_2545,N_2093);
and U3355 (N_3355,N_2639,N_2605);
nand U3356 (N_3356,N_2059,N_2341);
nor U3357 (N_3357,N_2125,N_2337);
and U3358 (N_3358,N_2232,N_2002);
xor U3359 (N_3359,N_2280,N_2458);
nand U3360 (N_3360,N_2946,N_2129);
nand U3361 (N_3361,N_2861,N_2481);
xor U3362 (N_3362,N_2148,N_2180);
nand U3363 (N_3363,N_2437,N_2415);
nor U3364 (N_3364,N_2429,N_2217);
nand U3365 (N_3365,N_2087,N_2445);
nor U3366 (N_3366,N_2535,N_2594);
xor U3367 (N_3367,N_2143,N_2350);
nor U3368 (N_3368,N_2151,N_2988);
nor U3369 (N_3369,N_2644,N_2078);
or U3370 (N_3370,N_2537,N_2301);
nand U3371 (N_3371,N_2772,N_2977);
and U3372 (N_3372,N_2502,N_2879);
xor U3373 (N_3373,N_2969,N_2939);
nor U3374 (N_3374,N_2735,N_2768);
nor U3375 (N_3375,N_2110,N_2330);
or U3376 (N_3376,N_2242,N_2848);
xor U3377 (N_3377,N_2598,N_2205);
nor U3378 (N_3378,N_2480,N_2477);
and U3379 (N_3379,N_2992,N_2252);
xnor U3380 (N_3380,N_2244,N_2622);
or U3381 (N_3381,N_2077,N_2897);
nand U3382 (N_3382,N_2010,N_2542);
nand U3383 (N_3383,N_2869,N_2181);
or U3384 (N_3384,N_2859,N_2256);
xnor U3385 (N_3385,N_2486,N_2120);
nor U3386 (N_3386,N_2024,N_2052);
nand U3387 (N_3387,N_2620,N_2100);
xnor U3388 (N_3388,N_2800,N_2479);
or U3389 (N_3389,N_2327,N_2172);
or U3390 (N_3390,N_2720,N_2748);
nand U3391 (N_3391,N_2609,N_2727);
nand U3392 (N_3392,N_2389,N_2184);
xor U3393 (N_3393,N_2173,N_2421);
or U3394 (N_3394,N_2306,N_2032);
xnor U3395 (N_3395,N_2987,N_2767);
or U3396 (N_3396,N_2331,N_2057);
or U3397 (N_3397,N_2973,N_2376);
or U3398 (N_3398,N_2201,N_2971);
and U3399 (N_3399,N_2235,N_2150);
and U3400 (N_3400,N_2587,N_2051);
or U3401 (N_3401,N_2934,N_2021);
nor U3402 (N_3402,N_2084,N_2638);
nand U3403 (N_3403,N_2736,N_2130);
and U3404 (N_3404,N_2771,N_2655);
nand U3405 (N_3405,N_2647,N_2906);
or U3406 (N_3406,N_2769,N_2025);
or U3407 (N_3407,N_2431,N_2108);
nor U3408 (N_3408,N_2118,N_2671);
nor U3409 (N_3409,N_2241,N_2841);
xnor U3410 (N_3410,N_2564,N_2894);
xnor U3411 (N_3411,N_2109,N_2866);
or U3412 (N_3412,N_2815,N_2509);
xor U3413 (N_3413,N_2141,N_2055);
nand U3414 (N_3414,N_2160,N_2676);
xor U3415 (N_3415,N_2806,N_2776);
or U3416 (N_3416,N_2628,N_2139);
nand U3417 (N_3417,N_2267,N_2107);
nor U3418 (N_3418,N_2782,N_2424);
and U3419 (N_3419,N_2105,N_2678);
nor U3420 (N_3420,N_2659,N_2403);
xnor U3421 (N_3421,N_2036,N_2670);
and U3422 (N_3422,N_2709,N_2989);
xor U3423 (N_3423,N_2484,N_2530);
xor U3424 (N_3424,N_2285,N_2367);
nor U3425 (N_3425,N_2812,N_2557);
and U3426 (N_3426,N_2493,N_2284);
xnor U3427 (N_3427,N_2819,N_2741);
xor U3428 (N_3428,N_2243,N_2076);
and U3429 (N_3429,N_2329,N_2809);
or U3430 (N_3430,N_2397,N_2588);
and U3431 (N_3431,N_2065,N_2286);
nand U3432 (N_3432,N_2266,N_2524);
nand U3433 (N_3433,N_2345,N_2586);
nor U3434 (N_3434,N_2166,N_2121);
nor U3435 (N_3435,N_2339,N_2875);
nand U3436 (N_3436,N_2759,N_2577);
nand U3437 (N_3437,N_2461,N_2877);
nor U3438 (N_3438,N_2045,N_2124);
nand U3439 (N_3439,N_2062,N_2667);
and U3440 (N_3440,N_2335,N_2891);
or U3441 (N_3441,N_2466,N_2452);
nor U3442 (N_3442,N_2296,N_2056);
nor U3443 (N_3443,N_2705,N_2186);
xor U3444 (N_3444,N_2190,N_2260);
xnor U3445 (N_3445,N_2567,N_2774);
or U3446 (N_3446,N_2503,N_2138);
and U3447 (N_3447,N_2648,N_2001);
or U3448 (N_3448,N_2070,N_2346);
or U3449 (N_3449,N_2325,N_2414);
nor U3450 (N_3450,N_2398,N_2029);
or U3451 (N_3451,N_2309,N_2195);
and U3452 (N_3452,N_2965,N_2153);
and U3453 (N_3453,N_2058,N_2436);
and U3454 (N_3454,N_2276,N_2696);
nor U3455 (N_3455,N_2115,N_2383);
and U3456 (N_3456,N_2438,N_2061);
xor U3457 (N_3457,N_2457,N_2944);
or U3458 (N_3458,N_2682,N_2905);
nor U3459 (N_3459,N_2935,N_2880);
nand U3460 (N_3460,N_2830,N_2786);
xnor U3461 (N_3461,N_2821,N_2279);
or U3462 (N_3462,N_2713,N_2433);
xnor U3463 (N_3463,N_2918,N_2575);
nor U3464 (N_3464,N_2822,N_2983);
nor U3465 (N_3465,N_2641,N_2817);
xor U3466 (N_3466,N_2672,N_2846);
nor U3467 (N_3467,N_2066,N_2656);
and U3468 (N_3468,N_2155,N_2686);
nor U3469 (N_3469,N_2310,N_2914);
nor U3470 (N_3470,N_2292,N_2147);
nor U3471 (N_3471,N_2719,N_2930);
nand U3472 (N_3472,N_2708,N_2023);
nor U3473 (N_3473,N_2342,N_2625);
or U3474 (N_3474,N_2185,N_2264);
nand U3475 (N_3475,N_2972,N_2829);
xor U3476 (N_3476,N_2456,N_2469);
and U3477 (N_3477,N_2478,N_2745);
xnor U3478 (N_3478,N_2472,N_2362);
or U3479 (N_3479,N_2450,N_2140);
or U3480 (N_3480,N_2602,N_2623);
and U3481 (N_3481,N_2707,N_2455);
and U3482 (N_3482,N_2511,N_2614);
nor U3483 (N_3483,N_2432,N_2191);
and U3484 (N_3484,N_2508,N_2729);
xnor U3485 (N_3485,N_2251,N_2571);
or U3486 (N_3486,N_2921,N_2282);
and U3487 (N_3487,N_2314,N_2742);
and U3488 (N_3488,N_2600,N_2521);
nand U3489 (N_3489,N_2712,N_2572);
nand U3490 (N_3490,N_2144,N_2816);
nor U3491 (N_3491,N_2340,N_2099);
or U3492 (N_3492,N_2599,N_2611);
nand U3493 (N_3493,N_2192,N_2505);
nor U3494 (N_3494,N_2968,N_2828);
or U3495 (N_3495,N_2617,N_2993);
or U3496 (N_3496,N_2210,N_2303);
nand U3497 (N_3497,N_2827,N_2248);
or U3498 (N_3498,N_2420,N_2356);
and U3499 (N_3499,N_2312,N_2365);
xor U3500 (N_3500,N_2344,N_2511);
and U3501 (N_3501,N_2230,N_2385);
and U3502 (N_3502,N_2908,N_2180);
or U3503 (N_3503,N_2352,N_2426);
nor U3504 (N_3504,N_2241,N_2318);
nand U3505 (N_3505,N_2941,N_2086);
xor U3506 (N_3506,N_2739,N_2749);
xnor U3507 (N_3507,N_2898,N_2080);
nand U3508 (N_3508,N_2722,N_2609);
xor U3509 (N_3509,N_2396,N_2882);
nor U3510 (N_3510,N_2770,N_2232);
nor U3511 (N_3511,N_2478,N_2770);
and U3512 (N_3512,N_2637,N_2922);
nand U3513 (N_3513,N_2212,N_2489);
nand U3514 (N_3514,N_2016,N_2699);
xnor U3515 (N_3515,N_2056,N_2317);
or U3516 (N_3516,N_2272,N_2289);
or U3517 (N_3517,N_2715,N_2728);
nand U3518 (N_3518,N_2366,N_2737);
xnor U3519 (N_3519,N_2901,N_2735);
and U3520 (N_3520,N_2984,N_2715);
nand U3521 (N_3521,N_2582,N_2392);
xor U3522 (N_3522,N_2555,N_2679);
nand U3523 (N_3523,N_2783,N_2079);
nand U3524 (N_3524,N_2100,N_2288);
or U3525 (N_3525,N_2697,N_2113);
or U3526 (N_3526,N_2764,N_2191);
or U3527 (N_3527,N_2675,N_2700);
and U3528 (N_3528,N_2828,N_2821);
nor U3529 (N_3529,N_2620,N_2273);
or U3530 (N_3530,N_2402,N_2089);
and U3531 (N_3531,N_2256,N_2234);
xor U3532 (N_3532,N_2006,N_2957);
nor U3533 (N_3533,N_2082,N_2862);
nor U3534 (N_3534,N_2308,N_2591);
or U3535 (N_3535,N_2925,N_2864);
and U3536 (N_3536,N_2354,N_2246);
nand U3537 (N_3537,N_2909,N_2138);
xor U3538 (N_3538,N_2936,N_2177);
and U3539 (N_3539,N_2044,N_2782);
xor U3540 (N_3540,N_2871,N_2466);
nand U3541 (N_3541,N_2219,N_2971);
xnor U3542 (N_3542,N_2470,N_2257);
or U3543 (N_3543,N_2065,N_2740);
nand U3544 (N_3544,N_2451,N_2638);
xor U3545 (N_3545,N_2708,N_2701);
and U3546 (N_3546,N_2421,N_2962);
nor U3547 (N_3547,N_2819,N_2311);
nor U3548 (N_3548,N_2060,N_2632);
and U3549 (N_3549,N_2116,N_2411);
and U3550 (N_3550,N_2189,N_2770);
or U3551 (N_3551,N_2035,N_2466);
and U3552 (N_3552,N_2314,N_2759);
nor U3553 (N_3553,N_2667,N_2270);
nor U3554 (N_3554,N_2501,N_2335);
or U3555 (N_3555,N_2927,N_2559);
xor U3556 (N_3556,N_2610,N_2604);
nor U3557 (N_3557,N_2812,N_2890);
or U3558 (N_3558,N_2888,N_2993);
nor U3559 (N_3559,N_2823,N_2619);
nand U3560 (N_3560,N_2923,N_2246);
or U3561 (N_3561,N_2519,N_2488);
nor U3562 (N_3562,N_2663,N_2046);
nand U3563 (N_3563,N_2377,N_2115);
nor U3564 (N_3564,N_2685,N_2469);
and U3565 (N_3565,N_2690,N_2653);
xor U3566 (N_3566,N_2663,N_2958);
and U3567 (N_3567,N_2973,N_2540);
xnor U3568 (N_3568,N_2179,N_2040);
nor U3569 (N_3569,N_2511,N_2551);
nand U3570 (N_3570,N_2946,N_2131);
xnor U3571 (N_3571,N_2511,N_2347);
nor U3572 (N_3572,N_2015,N_2302);
nand U3573 (N_3573,N_2204,N_2303);
and U3574 (N_3574,N_2973,N_2679);
and U3575 (N_3575,N_2785,N_2650);
nor U3576 (N_3576,N_2541,N_2669);
nand U3577 (N_3577,N_2498,N_2059);
or U3578 (N_3578,N_2086,N_2363);
nand U3579 (N_3579,N_2953,N_2564);
and U3580 (N_3580,N_2094,N_2302);
nand U3581 (N_3581,N_2034,N_2298);
or U3582 (N_3582,N_2220,N_2443);
and U3583 (N_3583,N_2392,N_2436);
or U3584 (N_3584,N_2367,N_2765);
and U3585 (N_3585,N_2563,N_2287);
or U3586 (N_3586,N_2839,N_2419);
nand U3587 (N_3587,N_2819,N_2728);
and U3588 (N_3588,N_2348,N_2750);
or U3589 (N_3589,N_2174,N_2437);
and U3590 (N_3590,N_2477,N_2553);
xnor U3591 (N_3591,N_2312,N_2183);
xnor U3592 (N_3592,N_2943,N_2330);
xnor U3593 (N_3593,N_2591,N_2978);
and U3594 (N_3594,N_2071,N_2925);
or U3595 (N_3595,N_2922,N_2781);
and U3596 (N_3596,N_2712,N_2498);
and U3597 (N_3597,N_2219,N_2397);
xor U3598 (N_3598,N_2333,N_2826);
and U3599 (N_3599,N_2407,N_2560);
nand U3600 (N_3600,N_2761,N_2951);
xor U3601 (N_3601,N_2467,N_2910);
and U3602 (N_3602,N_2249,N_2447);
and U3603 (N_3603,N_2962,N_2456);
nor U3604 (N_3604,N_2762,N_2551);
xor U3605 (N_3605,N_2747,N_2911);
and U3606 (N_3606,N_2101,N_2830);
or U3607 (N_3607,N_2628,N_2881);
nand U3608 (N_3608,N_2863,N_2371);
xor U3609 (N_3609,N_2219,N_2858);
or U3610 (N_3610,N_2814,N_2190);
xnor U3611 (N_3611,N_2588,N_2895);
and U3612 (N_3612,N_2622,N_2217);
xor U3613 (N_3613,N_2237,N_2141);
xor U3614 (N_3614,N_2302,N_2077);
or U3615 (N_3615,N_2523,N_2315);
nand U3616 (N_3616,N_2072,N_2245);
xor U3617 (N_3617,N_2888,N_2246);
or U3618 (N_3618,N_2670,N_2712);
xnor U3619 (N_3619,N_2181,N_2578);
nor U3620 (N_3620,N_2975,N_2017);
xnor U3621 (N_3621,N_2511,N_2582);
nand U3622 (N_3622,N_2108,N_2193);
or U3623 (N_3623,N_2336,N_2680);
nand U3624 (N_3624,N_2625,N_2774);
nor U3625 (N_3625,N_2666,N_2608);
or U3626 (N_3626,N_2318,N_2388);
xnor U3627 (N_3627,N_2074,N_2405);
or U3628 (N_3628,N_2440,N_2433);
nor U3629 (N_3629,N_2369,N_2609);
nand U3630 (N_3630,N_2450,N_2192);
nor U3631 (N_3631,N_2166,N_2750);
and U3632 (N_3632,N_2676,N_2977);
or U3633 (N_3633,N_2610,N_2831);
and U3634 (N_3634,N_2062,N_2484);
nand U3635 (N_3635,N_2559,N_2424);
nand U3636 (N_3636,N_2689,N_2278);
and U3637 (N_3637,N_2329,N_2649);
or U3638 (N_3638,N_2713,N_2964);
and U3639 (N_3639,N_2900,N_2843);
nor U3640 (N_3640,N_2119,N_2502);
nand U3641 (N_3641,N_2814,N_2967);
nor U3642 (N_3642,N_2046,N_2950);
nand U3643 (N_3643,N_2350,N_2865);
xnor U3644 (N_3644,N_2242,N_2801);
and U3645 (N_3645,N_2967,N_2332);
and U3646 (N_3646,N_2876,N_2802);
nand U3647 (N_3647,N_2251,N_2932);
xnor U3648 (N_3648,N_2359,N_2212);
xnor U3649 (N_3649,N_2357,N_2438);
and U3650 (N_3650,N_2920,N_2314);
and U3651 (N_3651,N_2034,N_2021);
nand U3652 (N_3652,N_2542,N_2731);
or U3653 (N_3653,N_2370,N_2936);
or U3654 (N_3654,N_2389,N_2867);
nor U3655 (N_3655,N_2038,N_2693);
and U3656 (N_3656,N_2170,N_2633);
and U3657 (N_3657,N_2456,N_2278);
xnor U3658 (N_3658,N_2069,N_2334);
and U3659 (N_3659,N_2062,N_2835);
nor U3660 (N_3660,N_2935,N_2085);
xnor U3661 (N_3661,N_2332,N_2697);
or U3662 (N_3662,N_2305,N_2632);
xor U3663 (N_3663,N_2687,N_2018);
nor U3664 (N_3664,N_2984,N_2935);
nor U3665 (N_3665,N_2764,N_2475);
and U3666 (N_3666,N_2211,N_2745);
nand U3667 (N_3667,N_2802,N_2867);
nor U3668 (N_3668,N_2335,N_2191);
nand U3669 (N_3669,N_2447,N_2762);
nor U3670 (N_3670,N_2836,N_2204);
nor U3671 (N_3671,N_2834,N_2219);
nor U3672 (N_3672,N_2897,N_2786);
or U3673 (N_3673,N_2449,N_2210);
nor U3674 (N_3674,N_2420,N_2864);
nand U3675 (N_3675,N_2376,N_2584);
nand U3676 (N_3676,N_2327,N_2334);
and U3677 (N_3677,N_2800,N_2564);
nand U3678 (N_3678,N_2851,N_2820);
and U3679 (N_3679,N_2476,N_2479);
nor U3680 (N_3680,N_2015,N_2944);
nand U3681 (N_3681,N_2887,N_2028);
xnor U3682 (N_3682,N_2895,N_2973);
xor U3683 (N_3683,N_2814,N_2520);
or U3684 (N_3684,N_2005,N_2298);
nand U3685 (N_3685,N_2374,N_2713);
and U3686 (N_3686,N_2620,N_2227);
or U3687 (N_3687,N_2687,N_2389);
nor U3688 (N_3688,N_2173,N_2340);
or U3689 (N_3689,N_2591,N_2841);
and U3690 (N_3690,N_2283,N_2631);
nand U3691 (N_3691,N_2674,N_2993);
and U3692 (N_3692,N_2558,N_2833);
nor U3693 (N_3693,N_2908,N_2480);
and U3694 (N_3694,N_2308,N_2928);
or U3695 (N_3695,N_2014,N_2193);
or U3696 (N_3696,N_2429,N_2288);
nand U3697 (N_3697,N_2473,N_2280);
xnor U3698 (N_3698,N_2251,N_2764);
and U3699 (N_3699,N_2817,N_2879);
nand U3700 (N_3700,N_2123,N_2984);
nand U3701 (N_3701,N_2176,N_2607);
or U3702 (N_3702,N_2503,N_2100);
and U3703 (N_3703,N_2968,N_2644);
nor U3704 (N_3704,N_2380,N_2232);
nor U3705 (N_3705,N_2860,N_2840);
xnor U3706 (N_3706,N_2160,N_2111);
nor U3707 (N_3707,N_2953,N_2559);
and U3708 (N_3708,N_2688,N_2365);
or U3709 (N_3709,N_2100,N_2233);
nor U3710 (N_3710,N_2171,N_2352);
xor U3711 (N_3711,N_2857,N_2908);
or U3712 (N_3712,N_2483,N_2359);
xnor U3713 (N_3713,N_2156,N_2506);
nand U3714 (N_3714,N_2244,N_2958);
nor U3715 (N_3715,N_2553,N_2727);
and U3716 (N_3716,N_2699,N_2085);
and U3717 (N_3717,N_2168,N_2681);
nand U3718 (N_3718,N_2000,N_2054);
xnor U3719 (N_3719,N_2587,N_2416);
nor U3720 (N_3720,N_2002,N_2014);
or U3721 (N_3721,N_2048,N_2966);
and U3722 (N_3722,N_2154,N_2510);
nand U3723 (N_3723,N_2280,N_2562);
nor U3724 (N_3724,N_2243,N_2627);
or U3725 (N_3725,N_2054,N_2091);
xor U3726 (N_3726,N_2082,N_2645);
nor U3727 (N_3727,N_2757,N_2419);
nand U3728 (N_3728,N_2394,N_2944);
xor U3729 (N_3729,N_2326,N_2560);
or U3730 (N_3730,N_2719,N_2430);
or U3731 (N_3731,N_2955,N_2705);
and U3732 (N_3732,N_2934,N_2235);
xor U3733 (N_3733,N_2879,N_2262);
or U3734 (N_3734,N_2278,N_2373);
or U3735 (N_3735,N_2739,N_2900);
and U3736 (N_3736,N_2542,N_2256);
xnor U3737 (N_3737,N_2760,N_2952);
nand U3738 (N_3738,N_2832,N_2855);
and U3739 (N_3739,N_2723,N_2404);
xnor U3740 (N_3740,N_2973,N_2225);
and U3741 (N_3741,N_2540,N_2868);
and U3742 (N_3742,N_2276,N_2446);
nor U3743 (N_3743,N_2593,N_2927);
or U3744 (N_3744,N_2928,N_2712);
xor U3745 (N_3745,N_2605,N_2877);
nand U3746 (N_3746,N_2916,N_2552);
nand U3747 (N_3747,N_2374,N_2734);
and U3748 (N_3748,N_2486,N_2503);
xor U3749 (N_3749,N_2898,N_2987);
xor U3750 (N_3750,N_2203,N_2328);
xor U3751 (N_3751,N_2761,N_2104);
nand U3752 (N_3752,N_2031,N_2415);
nand U3753 (N_3753,N_2004,N_2222);
nor U3754 (N_3754,N_2677,N_2816);
nor U3755 (N_3755,N_2650,N_2013);
nand U3756 (N_3756,N_2193,N_2795);
xnor U3757 (N_3757,N_2959,N_2217);
xor U3758 (N_3758,N_2142,N_2601);
nand U3759 (N_3759,N_2423,N_2197);
nand U3760 (N_3760,N_2082,N_2700);
or U3761 (N_3761,N_2161,N_2001);
nor U3762 (N_3762,N_2777,N_2840);
nor U3763 (N_3763,N_2625,N_2188);
and U3764 (N_3764,N_2817,N_2222);
xnor U3765 (N_3765,N_2229,N_2726);
nand U3766 (N_3766,N_2812,N_2341);
xnor U3767 (N_3767,N_2316,N_2441);
nor U3768 (N_3768,N_2975,N_2016);
nand U3769 (N_3769,N_2581,N_2271);
or U3770 (N_3770,N_2827,N_2703);
nor U3771 (N_3771,N_2785,N_2262);
and U3772 (N_3772,N_2124,N_2249);
nor U3773 (N_3773,N_2057,N_2682);
or U3774 (N_3774,N_2807,N_2823);
nand U3775 (N_3775,N_2562,N_2097);
or U3776 (N_3776,N_2602,N_2127);
nor U3777 (N_3777,N_2503,N_2175);
nor U3778 (N_3778,N_2026,N_2083);
and U3779 (N_3779,N_2229,N_2717);
xnor U3780 (N_3780,N_2903,N_2529);
nor U3781 (N_3781,N_2515,N_2366);
or U3782 (N_3782,N_2402,N_2541);
or U3783 (N_3783,N_2375,N_2850);
nand U3784 (N_3784,N_2805,N_2266);
and U3785 (N_3785,N_2762,N_2307);
nand U3786 (N_3786,N_2179,N_2021);
or U3787 (N_3787,N_2999,N_2883);
nand U3788 (N_3788,N_2024,N_2534);
and U3789 (N_3789,N_2632,N_2270);
nor U3790 (N_3790,N_2957,N_2141);
or U3791 (N_3791,N_2977,N_2937);
and U3792 (N_3792,N_2251,N_2286);
xor U3793 (N_3793,N_2931,N_2730);
nand U3794 (N_3794,N_2346,N_2908);
xor U3795 (N_3795,N_2656,N_2336);
nor U3796 (N_3796,N_2738,N_2425);
and U3797 (N_3797,N_2646,N_2963);
nand U3798 (N_3798,N_2278,N_2924);
and U3799 (N_3799,N_2983,N_2923);
or U3800 (N_3800,N_2808,N_2801);
xnor U3801 (N_3801,N_2641,N_2428);
or U3802 (N_3802,N_2440,N_2648);
or U3803 (N_3803,N_2479,N_2854);
nor U3804 (N_3804,N_2047,N_2655);
nand U3805 (N_3805,N_2506,N_2538);
or U3806 (N_3806,N_2962,N_2485);
nor U3807 (N_3807,N_2100,N_2830);
xor U3808 (N_3808,N_2958,N_2827);
nor U3809 (N_3809,N_2135,N_2723);
and U3810 (N_3810,N_2228,N_2355);
nor U3811 (N_3811,N_2976,N_2911);
or U3812 (N_3812,N_2338,N_2342);
nand U3813 (N_3813,N_2298,N_2792);
or U3814 (N_3814,N_2061,N_2670);
nand U3815 (N_3815,N_2063,N_2105);
nand U3816 (N_3816,N_2096,N_2306);
nor U3817 (N_3817,N_2477,N_2651);
and U3818 (N_3818,N_2581,N_2044);
or U3819 (N_3819,N_2551,N_2944);
or U3820 (N_3820,N_2191,N_2992);
or U3821 (N_3821,N_2587,N_2899);
nand U3822 (N_3822,N_2494,N_2934);
xor U3823 (N_3823,N_2967,N_2532);
xor U3824 (N_3824,N_2632,N_2478);
or U3825 (N_3825,N_2981,N_2415);
nand U3826 (N_3826,N_2104,N_2974);
or U3827 (N_3827,N_2239,N_2906);
xnor U3828 (N_3828,N_2759,N_2515);
or U3829 (N_3829,N_2080,N_2775);
nand U3830 (N_3830,N_2225,N_2087);
nor U3831 (N_3831,N_2344,N_2649);
xor U3832 (N_3832,N_2331,N_2046);
and U3833 (N_3833,N_2484,N_2969);
or U3834 (N_3834,N_2939,N_2878);
nand U3835 (N_3835,N_2539,N_2949);
nor U3836 (N_3836,N_2726,N_2625);
xnor U3837 (N_3837,N_2787,N_2775);
or U3838 (N_3838,N_2130,N_2452);
or U3839 (N_3839,N_2405,N_2822);
and U3840 (N_3840,N_2504,N_2982);
xor U3841 (N_3841,N_2576,N_2556);
nand U3842 (N_3842,N_2507,N_2032);
xnor U3843 (N_3843,N_2770,N_2538);
xnor U3844 (N_3844,N_2660,N_2436);
nand U3845 (N_3845,N_2108,N_2652);
xor U3846 (N_3846,N_2820,N_2034);
nand U3847 (N_3847,N_2349,N_2603);
xor U3848 (N_3848,N_2499,N_2369);
nor U3849 (N_3849,N_2479,N_2287);
xor U3850 (N_3850,N_2910,N_2248);
or U3851 (N_3851,N_2988,N_2590);
or U3852 (N_3852,N_2824,N_2439);
nor U3853 (N_3853,N_2379,N_2482);
and U3854 (N_3854,N_2275,N_2950);
nor U3855 (N_3855,N_2538,N_2482);
nor U3856 (N_3856,N_2164,N_2046);
xor U3857 (N_3857,N_2668,N_2988);
nor U3858 (N_3858,N_2892,N_2557);
or U3859 (N_3859,N_2193,N_2311);
and U3860 (N_3860,N_2836,N_2424);
and U3861 (N_3861,N_2237,N_2130);
nor U3862 (N_3862,N_2000,N_2633);
nor U3863 (N_3863,N_2801,N_2113);
nand U3864 (N_3864,N_2391,N_2129);
nor U3865 (N_3865,N_2603,N_2335);
nand U3866 (N_3866,N_2852,N_2889);
or U3867 (N_3867,N_2957,N_2829);
nand U3868 (N_3868,N_2685,N_2171);
nand U3869 (N_3869,N_2011,N_2138);
nor U3870 (N_3870,N_2225,N_2506);
xor U3871 (N_3871,N_2173,N_2424);
or U3872 (N_3872,N_2843,N_2015);
or U3873 (N_3873,N_2927,N_2729);
nand U3874 (N_3874,N_2644,N_2818);
or U3875 (N_3875,N_2701,N_2555);
xnor U3876 (N_3876,N_2099,N_2312);
nand U3877 (N_3877,N_2779,N_2658);
and U3878 (N_3878,N_2936,N_2249);
or U3879 (N_3879,N_2333,N_2087);
and U3880 (N_3880,N_2575,N_2904);
xnor U3881 (N_3881,N_2922,N_2867);
or U3882 (N_3882,N_2235,N_2297);
nor U3883 (N_3883,N_2719,N_2811);
or U3884 (N_3884,N_2085,N_2689);
or U3885 (N_3885,N_2521,N_2727);
nand U3886 (N_3886,N_2187,N_2117);
and U3887 (N_3887,N_2050,N_2305);
nand U3888 (N_3888,N_2746,N_2747);
or U3889 (N_3889,N_2054,N_2337);
and U3890 (N_3890,N_2848,N_2459);
and U3891 (N_3891,N_2704,N_2206);
and U3892 (N_3892,N_2644,N_2534);
nor U3893 (N_3893,N_2001,N_2284);
or U3894 (N_3894,N_2032,N_2835);
nor U3895 (N_3895,N_2825,N_2287);
or U3896 (N_3896,N_2527,N_2742);
nand U3897 (N_3897,N_2953,N_2526);
and U3898 (N_3898,N_2726,N_2913);
xnor U3899 (N_3899,N_2735,N_2682);
nor U3900 (N_3900,N_2353,N_2670);
xor U3901 (N_3901,N_2012,N_2870);
nor U3902 (N_3902,N_2848,N_2080);
or U3903 (N_3903,N_2503,N_2371);
nand U3904 (N_3904,N_2504,N_2100);
xnor U3905 (N_3905,N_2253,N_2849);
or U3906 (N_3906,N_2384,N_2041);
xor U3907 (N_3907,N_2082,N_2618);
or U3908 (N_3908,N_2653,N_2482);
and U3909 (N_3909,N_2189,N_2002);
or U3910 (N_3910,N_2920,N_2069);
nand U3911 (N_3911,N_2315,N_2117);
and U3912 (N_3912,N_2819,N_2813);
xnor U3913 (N_3913,N_2626,N_2371);
and U3914 (N_3914,N_2725,N_2757);
nor U3915 (N_3915,N_2402,N_2880);
or U3916 (N_3916,N_2383,N_2233);
nor U3917 (N_3917,N_2008,N_2354);
or U3918 (N_3918,N_2752,N_2877);
nor U3919 (N_3919,N_2687,N_2713);
and U3920 (N_3920,N_2628,N_2655);
or U3921 (N_3921,N_2071,N_2628);
or U3922 (N_3922,N_2613,N_2236);
or U3923 (N_3923,N_2009,N_2113);
xnor U3924 (N_3924,N_2802,N_2689);
and U3925 (N_3925,N_2842,N_2017);
xor U3926 (N_3926,N_2744,N_2559);
nor U3927 (N_3927,N_2844,N_2362);
or U3928 (N_3928,N_2448,N_2103);
nor U3929 (N_3929,N_2237,N_2064);
and U3930 (N_3930,N_2361,N_2556);
or U3931 (N_3931,N_2312,N_2238);
nor U3932 (N_3932,N_2351,N_2860);
or U3933 (N_3933,N_2115,N_2735);
nor U3934 (N_3934,N_2410,N_2779);
nor U3935 (N_3935,N_2173,N_2118);
nor U3936 (N_3936,N_2575,N_2104);
and U3937 (N_3937,N_2064,N_2331);
xor U3938 (N_3938,N_2868,N_2746);
nand U3939 (N_3939,N_2126,N_2713);
xnor U3940 (N_3940,N_2224,N_2115);
xor U3941 (N_3941,N_2309,N_2016);
nor U3942 (N_3942,N_2136,N_2341);
or U3943 (N_3943,N_2033,N_2768);
or U3944 (N_3944,N_2749,N_2753);
nand U3945 (N_3945,N_2754,N_2879);
and U3946 (N_3946,N_2766,N_2709);
or U3947 (N_3947,N_2893,N_2199);
or U3948 (N_3948,N_2840,N_2950);
nor U3949 (N_3949,N_2889,N_2611);
and U3950 (N_3950,N_2250,N_2209);
and U3951 (N_3951,N_2525,N_2513);
or U3952 (N_3952,N_2629,N_2319);
nand U3953 (N_3953,N_2508,N_2354);
and U3954 (N_3954,N_2980,N_2314);
and U3955 (N_3955,N_2501,N_2202);
nand U3956 (N_3956,N_2079,N_2573);
or U3957 (N_3957,N_2926,N_2660);
nor U3958 (N_3958,N_2265,N_2812);
nor U3959 (N_3959,N_2365,N_2926);
xor U3960 (N_3960,N_2254,N_2367);
nand U3961 (N_3961,N_2025,N_2683);
xor U3962 (N_3962,N_2423,N_2895);
nand U3963 (N_3963,N_2249,N_2652);
nand U3964 (N_3964,N_2288,N_2711);
or U3965 (N_3965,N_2017,N_2744);
or U3966 (N_3966,N_2549,N_2922);
nor U3967 (N_3967,N_2546,N_2392);
or U3968 (N_3968,N_2253,N_2134);
xor U3969 (N_3969,N_2799,N_2885);
nor U3970 (N_3970,N_2597,N_2983);
and U3971 (N_3971,N_2935,N_2129);
nor U3972 (N_3972,N_2425,N_2606);
and U3973 (N_3973,N_2720,N_2391);
nand U3974 (N_3974,N_2538,N_2167);
and U3975 (N_3975,N_2706,N_2445);
or U3976 (N_3976,N_2929,N_2290);
nor U3977 (N_3977,N_2665,N_2441);
nand U3978 (N_3978,N_2994,N_2771);
xor U3979 (N_3979,N_2239,N_2682);
nand U3980 (N_3980,N_2193,N_2906);
nor U3981 (N_3981,N_2942,N_2718);
nor U3982 (N_3982,N_2857,N_2636);
xnor U3983 (N_3983,N_2329,N_2083);
or U3984 (N_3984,N_2230,N_2986);
or U3985 (N_3985,N_2078,N_2809);
or U3986 (N_3986,N_2636,N_2971);
nand U3987 (N_3987,N_2405,N_2956);
xor U3988 (N_3988,N_2655,N_2969);
xor U3989 (N_3989,N_2863,N_2696);
or U3990 (N_3990,N_2737,N_2753);
and U3991 (N_3991,N_2795,N_2978);
nor U3992 (N_3992,N_2711,N_2832);
nand U3993 (N_3993,N_2880,N_2982);
or U3994 (N_3994,N_2067,N_2335);
nand U3995 (N_3995,N_2357,N_2416);
nor U3996 (N_3996,N_2682,N_2165);
or U3997 (N_3997,N_2343,N_2176);
or U3998 (N_3998,N_2832,N_2225);
and U3999 (N_3999,N_2174,N_2730);
or U4000 (N_4000,N_3558,N_3456);
xnor U4001 (N_4001,N_3934,N_3866);
or U4002 (N_4002,N_3875,N_3687);
nor U4003 (N_4003,N_3825,N_3364);
nand U4004 (N_4004,N_3893,N_3677);
nand U4005 (N_4005,N_3539,N_3272);
and U4006 (N_4006,N_3701,N_3997);
xor U4007 (N_4007,N_3975,N_3665);
nand U4008 (N_4008,N_3847,N_3546);
and U4009 (N_4009,N_3421,N_3391);
nand U4010 (N_4010,N_3280,N_3327);
and U4011 (N_4011,N_3348,N_3644);
nor U4012 (N_4012,N_3511,N_3037);
or U4013 (N_4013,N_3014,N_3968);
nor U4014 (N_4014,N_3297,N_3843);
or U4015 (N_4015,N_3463,N_3640);
nor U4016 (N_4016,N_3886,N_3300);
nor U4017 (N_4017,N_3424,N_3061);
or U4018 (N_4018,N_3897,N_3279);
nand U4019 (N_4019,N_3213,N_3122);
xnor U4020 (N_4020,N_3199,N_3151);
nand U4021 (N_4021,N_3774,N_3885);
nor U4022 (N_4022,N_3075,N_3654);
xnor U4023 (N_4023,N_3854,N_3492);
nor U4024 (N_4024,N_3859,N_3556);
nor U4025 (N_4025,N_3594,N_3167);
nand U4026 (N_4026,N_3807,N_3464);
and U4027 (N_4027,N_3024,N_3744);
nor U4028 (N_4028,N_3725,N_3781);
xnor U4029 (N_4029,N_3475,N_3451);
or U4030 (N_4030,N_3684,N_3366);
and U4031 (N_4031,N_3699,N_3597);
nand U4032 (N_4032,N_3084,N_3328);
or U4033 (N_4033,N_3661,N_3285);
or U4034 (N_4034,N_3347,N_3214);
and U4035 (N_4035,N_3462,N_3414);
and U4036 (N_4036,N_3979,N_3824);
or U4037 (N_4037,N_3604,N_3229);
and U4038 (N_4038,N_3933,N_3208);
or U4039 (N_4039,N_3560,N_3612);
nand U4040 (N_4040,N_3787,N_3956);
and U4041 (N_4041,N_3810,N_3380);
and U4042 (N_4042,N_3867,N_3652);
or U4043 (N_4043,N_3330,N_3466);
and U4044 (N_4044,N_3157,N_3430);
or U4045 (N_4045,N_3760,N_3868);
or U4046 (N_4046,N_3941,N_3888);
and U4047 (N_4047,N_3924,N_3153);
and U4048 (N_4048,N_3210,N_3853);
nand U4049 (N_4049,N_3282,N_3555);
xnor U4050 (N_4050,N_3026,N_3392);
nor U4051 (N_4051,N_3929,N_3336);
or U4052 (N_4052,N_3107,N_3925);
nor U4053 (N_4053,N_3653,N_3735);
and U4054 (N_4054,N_3458,N_3508);
or U4055 (N_4055,N_3568,N_3309);
nor U4056 (N_4056,N_3940,N_3574);
and U4057 (N_4057,N_3871,N_3756);
nor U4058 (N_4058,N_3133,N_3729);
and U4059 (N_4059,N_3720,N_3340);
nor U4060 (N_4060,N_3147,N_3104);
nand U4061 (N_4061,N_3668,N_3862);
nand U4062 (N_4062,N_3160,N_3187);
nor U4063 (N_4063,N_3532,N_3740);
nand U4064 (N_4064,N_3450,N_3799);
and U4065 (N_4065,N_3333,N_3426);
nor U4066 (N_4066,N_3381,N_3298);
and U4067 (N_4067,N_3087,N_3240);
nor U4068 (N_4068,N_3609,N_3733);
nor U4069 (N_4069,N_3454,N_3571);
and U4070 (N_4070,N_3714,N_3409);
or U4071 (N_4071,N_3023,N_3144);
nor U4072 (N_4072,N_3196,N_3999);
xor U4073 (N_4073,N_3388,N_3750);
nor U4074 (N_4074,N_3683,N_3792);
xor U4075 (N_4075,N_3072,N_3191);
xor U4076 (N_4076,N_3625,N_3387);
or U4077 (N_4077,N_3166,N_3531);
and U4078 (N_4078,N_3922,N_3861);
nor U4079 (N_4079,N_3360,N_3656);
nor U4080 (N_4080,N_3936,N_3883);
or U4081 (N_4081,N_3616,N_3727);
nand U4082 (N_4082,N_3887,N_3826);
and U4083 (N_4083,N_3065,N_3168);
and U4084 (N_4084,N_3752,N_3648);
nor U4085 (N_4085,N_3846,N_3903);
nor U4086 (N_4086,N_3707,N_3217);
xor U4087 (N_4087,N_3278,N_3769);
xor U4088 (N_4088,N_3811,N_3263);
xor U4089 (N_4089,N_3954,N_3221);
or U4090 (N_4090,N_3193,N_3749);
xnor U4091 (N_4091,N_3899,N_3273);
xor U4092 (N_4092,N_3322,N_3383);
nor U4093 (N_4093,N_3599,N_3165);
or U4094 (N_4094,N_3216,N_3434);
nor U4095 (N_4095,N_3980,N_3775);
and U4096 (N_4096,N_3211,N_3629);
or U4097 (N_4097,N_3692,N_3863);
and U4098 (N_4098,N_3894,N_3709);
nor U4099 (N_4099,N_3027,N_3461);
and U4100 (N_4100,N_3751,N_3314);
or U4101 (N_4101,N_3164,N_3148);
or U4102 (N_4102,N_3909,N_3129);
nand U4103 (N_4103,N_3848,N_3840);
and U4104 (N_4104,N_3386,N_3858);
xnor U4105 (N_4105,N_3784,N_3682);
or U4106 (N_4106,N_3739,N_3962);
and U4107 (N_4107,N_3379,N_3693);
nand U4108 (N_4108,N_3576,N_3407);
xor U4109 (N_4109,N_3354,N_3519);
nor U4110 (N_4110,N_3542,N_3504);
nor U4111 (N_4111,N_3713,N_3534);
nand U4112 (N_4112,N_3185,N_3577);
or U4113 (N_4113,N_3961,N_3710);
and U4114 (N_4114,N_3223,N_3865);
xnor U4115 (N_4115,N_3702,N_3538);
xor U4116 (N_4116,N_3331,N_3262);
nand U4117 (N_4117,N_3851,N_3737);
nand U4118 (N_4118,N_3988,N_3939);
nor U4119 (N_4119,N_3044,N_3841);
nand U4120 (N_4120,N_3112,N_3412);
xor U4121 (N_4121,N_3753,N_3494);
and U4122 (N_4122,N_3382,N_3425);
nand U4123 (N_4123,N_3788,N_3473);
or U4124 (N_4124,N_3238,N_3204);
xnor U4125 (N_4125,N_3042,N_3305);
xnor U4126 (N_4126,N_3192,N_3332);
or U4127 (N_4127,N_3949,N_3397);
or U4128 (N_4128,N_3628,N_3928);
nand U4129 (N_4129,N_3646,N_3172);
nand U4130 (N_4130,N_3978,N_3415);
or U4131 (N_4131,N_3819,N_3666);
nand U4132 (N_4132,N_3943,N_3317);
and U4133 (N_4133,N_3783,N_3265);
xnor U4134 (N_4134,N_3659,N_3679);
and U4135 (N_4135,N_3780,N_3130);
nand U4136 (N_4136,N_3872,N_3343);
xor U4137 (N_4137,N_3022,N_3290);
or U4138 (N_4138,N_3231,N_3131);
nor U4139 (N_4139,N_3830,N_3664);
or U4140 (N_4140,N_3174,N_3245);
and U4141 (N_4141,N_3398,N_3685);
xor U4142 (N_4142,N_3662,N_3306);
and U4143 (N_4143,N_3353,N_3528);
nand U4144 (N_4144,N_3796,N_3005);
and U4145 (N_4145,N_3622,N_3159);
nor U4146 (N_4146,N_3062,N_3141);
or U4147 (N_4147,N_3632,N_3944);
or U4148 (N_4148,N_3277,N_3161);
xnor U4149 (N_4149,N_3335,N_3708);
or U4150 (N_4150,N_3338,N_3967);
nand U4151 (N_4151,N_3877,N_3891);
xnor U4152 (N_4152,N_3806,N_3512);
and U4153 (N_4153,N_3960,N_3384);
or U4154 (N_4154,N_3237,N_3908);
and U4155 (N_4155,N_3312,N_3323);
or U4156 (N_4156,N_3764,N_3698);
nand U4157 (N_4157,N_3031,N_3110);
nand U4158 (N_4158,N_3446,N_3636);
or U4159 (N_4159,N_3948,N_3755);
nand U4160 (N_4160,N_3743,N_3390);
or U4161 (N_4161,N_3319,N_3073);
nand U4162 (N_4162,N_3986,N_3125);
and U4163 (N_4163,N_3015,N_3591);
nor U4164 (N_4164,N_3517,N_3581);
nand U4165 (N_4165,N_3809,N_3205);
nor U4166 (N_4166,N_3671,N_3155);
or U4167 (N_4167,N_3089,N_3003);
nor U4168 (N_4168,N_3186,N_3996);
nor U4169 (N_4169,N_3880,N_3097);
nor U4170 (N_4170,N_3991,N_3728);
or U4171 (N_4171,N_3584,N_3063);
nor U4172 (N_4172,N_3496,N_3578);
nand U4173 (N_4173,N_3918,N_3705);
xor U4174 (N_4174,N_3209,N_3010);
nand U4175 (N_4175,N_3823,N_3178);
or U4176 (N_4176,N_3109,N_3467);
nor U4177 (N_4177,N_3259,N_3931);
nand U4178 (N_4178,N_3495,N_3481);
xor U4179 (N_4179,N_3183,N_3719);
and U4180 (N_4180,N_3444,N_3429);
xnor U4181 (N_4181,N_3930,N_3953);
xnor U4182 (N_4182,N_3798,N_3499);
nor U4183 (N_4183,N_3198,N_3378);
nand U4184 (N_4184,N_3078,N_3852);
nand U4185 (N_4185,N_3175,N_3535);
and U4186 (N_4186,N_3189,N_3971);
or U4187 (N_4187,N_3945,N_3505);
or U4188 (N_4188,N_3431,N_3795);
nand U4189 (N_4189,N_3541,N_3289);
nand U4190 (N_4190,N_3470,N_3608);
nand U4191 (N_4191,N_3672,N_3907);
nand U4192 (N_4192,N_3566,N_3833);
nand U4193 (N_4193,N_3995,N_3474);
nor U4194 (N_4194,N_3012,N_3455);
nor U4195 (N_4195,N_3603,N_3762);
nand U4196 (N_4196,N_3572,N_3688);
or U4197 (N_4197,N_3201,N_3067);
xnor U4198 (N_4198,N_3812,N_3817);
nor U4199 (N_4199,N_3800,N_3086);
nand U4200 (N_4200,N_3308,N_3963);
nand U4201 (N_4201,N_3989,N_3476);
nand U4202 (N_4202,N_3520,N_3724);
and U4203 (N_4203,N_3605,N_3587);
and U4204 (N_4204,N_3870,N_3586);
or U4205 (N_4205,N_3435,N_3334);
nor U4206 (N_4206,N_3385,N_3049);
nor U4207 (N_4207,N_3983,N_3770);
and U4208 (N_4208,N_3040,N_3103);
nand U4209 (N_4209,N_3452,N_3139);
xor U4210 (N_4210,N_3651,N_3181);
xnor U4211 (N_4211,N_3527,N_3606);
or U4212 (N_4212,N_3892,N_3100);
nand U4213 (N_4213,N_3469,N_3879);
and U4214 (N_4214,N_3487,N_3038);
xnor U4215 (N_4215,N_3241,N_3310);
nand U4216 (N_4216,N_3946,N_3914);
nand U4217 (N_4217,N_3836,N_3620);
nand U4218 (N_4218,N_3526,N_3919);
and U4219 (N_4219,N_3889,N_3445);
nand U4220 (N_4220,N_3856,N_3916);
nand U4221 (N_4221,N_3745,N_3715);
or U4222 (N_4222,N_3436,N_3127);
nor U4223 (N_4223,N_3051,N_3401);
nor U4224 (N_4224,N_3182,N_3904);
nor U4225 (N_4225,N_3643,N_3544);
and U4226 (N_4226,N_3902,N_3017);
and U4227 (N_4227,N_3497,N_3607);
xor U4228 (N_4228,N_3686,N_3250);
nand U4229 (N_4229,N_3096,N_3070);
or U4230 (N_4230,N_3530,N_3099);
xor U4231 (N_4231,N_3261,N_3068);
or U4232 (N_4232,N_3785,N_3802);
xnor U4233 (N_4233,N_3345,N_3778);
and U4234 (N_4234,N_3649,N_3188);
or U4235 (N_4235,N_3838,N_3869);
nor U4236 (N_4236,N_3264,N_3140);
xor U4237 (N_4237,N_3410,N_3485);
nor U4238 (N_4238,N_3641,N_3993);
nor U4239 (N_4239,N_3171,N_3457);
or U4240 (N_4240,N_3082,N_3021);
nand U4241 (N_4241,N_3712,N_3920);
or U4242 (N_4242,N_3882,N_3395);
or U4243 (N_4243,N_3344,N_3521);
nand U4244 (N_4244,N_3580,N_3901);
and U4245 (N_4245,N_3090,N_3118);
xnor U4246 (N_4246,N_3176,N_3489);
nand U4247 (N_4247,N_3184,N_3066);
or U4248 (N_4248,N_3137,N_3835);
nand U4249 (N_4249,N_3681,N_3459);
and U4250 (N_4250,N_3486,N_3570);
nor U4251 (N_4251,N_3437,N_3367);
and U4252 (N_4252,N_3913,N_3906);
or U4253 (N_4253,N_3611,N_3617);
nor U4254 (N_4254,N_3375,N_3767);
or U4255 (N_4255,N_3478,N_3060);
xnor U4256 (N_4256,N_3376,N_3094);
nor U4257 (N_4257,N_3325,N_3736);
and U4258 (N_4258,N_3621,N_3311);
nor U4259 (N_4259,N_3923,N_3561);
xor U4260 (N_4260,N_3019,N_3896);
or U4261 (N_4261,N_3032,N_3195);
nand U4262 (N_4262,N_3471,N_3860);
nor U4263 (N_4263,N_3763,N_3490);
nand U4264 (N_4264,N_3001,N_3433);
xnor U4265 (N_4265,N_3674,N_3428);
xor U4266 (N_4266,N_3507,N_3647);
xnor U4267 (N_4267,N_3563,N_3955);
xnor U4268 (N_4268,N_3329,N_3083);
and U4269 (N_4269,N_3585,N_3514);
and U4270 (N_4270,N_3226,N_3533);
or U4271 (N_4271,N_3670,N_3910);
nand U4272 (N_4272,N_3855,N_3121);
xor U4273 (N_4273,N_3552,N_3123);
nor U4274 (N_4274,N_3222,N_3018);
or U4275 (N_4275,N_3299,N_3583);
nor U4276 (N_4276,N_3203,N_3927);
nand U4277 (N_4277,N_3441,N_3194);
nor U4278 (N_4278,N_3480,N_3905);
or U4279 (N_4279,N_3614,N_3623);
nand U4280 (N_4280,N_3857,N_3593);
or U4281 (N_4281,N_3844,N_3251);
xor U4282 (N_4282,N_3248,N_3700);
nor U4283 (N_4283,N_3247,N_3054);
nor U4284 (N_4284,N_3837,N_3116);
or U4285 (N_4285,N_3639,N_3368);
and U4286 (N_4286,N_3417,N_3408);
or U4287 (N_4287,N_3361,N_3794);
xor U4288 (N_4288,N_3219,N_3808);
nand U4289 (N_4289,N_3832,N_3275);
nand U4290 (N_4290,N_3270,N_3746);
or U4291 (N_4291,N_3255,N_3041);
and U4292 (N_4292,N_3977,N_3631);
or U4293 (N_4293,N_3150,N_3797);
and U4294 (N_4294,N_3726,N_3224);
and U4295 (N_4295,N_3105,N_3589);
nor U4296 (N_4296,N_3200,N_3921);
or U4297 (N_4297,N_3493,N_3722);
nand U4298 (N_4298,N_3113,N_3950);
nor U4299 (N_4299,N_3453,N_3281);
xnor U4300 (N_4300,N_3418,N_3827);
xnor U4301 (N_4301,N_3202,N_3180);
nand U4302 (N_4302,N_3258,N_3301);
or U4303 (N_4303,N_3814,N_3690);
and U4304 (N_4304,N_3994,N_3667);
nor U4305 (N_4305,N_3337,N_3575);
xor U4306 (N_4306,N_3399,N_3657);
nor U4307 (N_4307,N_3321,N_3220);
nor U4308 (N_4308,N_3691,N_3134);
or U4309 (N_4309,N_3935,N_3356);
or U4310 (N_4310,N_3973,N_3377);
and U4311 (N_4311,N_3663,N_3937);
xor U4312 (N_4312,N_3260,N_3030);
and U4313 (N_4313,N_3716,N_3269);
nor U4314 (N_4314,N_3029,N_3154);
and U4315 (N_4315,N_3972,N_3992);
and U4316 (N_4316,N_3420,N_3732);
or U4317 (N_4317,N_3293,N_3235);
or U4318 (N_4318,N_3350,N_3349);
nand U4319 (N_4319,N_3400,N_3128);
and U4320 (N_4320,N_3284,N_3645);
and U4321 (N_4321,N_3465,N_3839);
nor U4322 (N_4322,N_3624,N_3460);
nor U4323 (N_4323,N_3567,N_3942);
and U4324 (N_4324,N_3016,N_3829);
or U4325 (N_4325,N_3998,N_3138);
or U4326 (N_4326,N_3816,N_3320);
or U4327 (N_4327,N_3080,N_3025);
nor U4328 (N_4328,N_3215,N_3197);
nor U4329 (N_4329,N_3782,N_3633);
xor U4330 (N_4330,N_3790,N_3926);
nor U4331 (N_4331,N_3419,N_3286);
nor U4332 (N_4332,N_3355,N_3416);
xor U4333 (N_4333,N_3900,N_3747);
nor U4334 (N_4334,N_3177,N_3506);
or U4335 (N_4335,N_3227,N_3052);
or U4336 (N_4336,N_3502,N_3403);
xor U4337 (N_4337,N_3036,N_3267);
nand U4338 (N_4338,N_3634,N_3969);
xnor U4339 (N_4339,N_3064,N_3766);
and U4340 (N_4340,N_3190,N_3370);
or U4341 (N_4341,N_3615,N_3675);
nand U4342 (N_4342,N_3438,N_3912);
nor U4343 (N_4343,N_3126,N_3503);
and U4344 (N_4344,N_3283,N_3516);
and U4345 (N_4345,N_3136,N_3706);
nor U4346 (N_4346,N_3596,N_3404);
nand U4347 (N_4347,N_3079,N_3111);
xnor U4348 (N_4348,N_3818,N_3525);
nor U4349 (N_4349,N_3120,N_3890);
nor U4350 (N_4350,N_3553,N_3917);
xor U4351 (N_4351,N_3050,N_3595);
xor U4352 (N_4352,N_3976,N_3772);
nand U4353 (N_4353,N_3842,N_3045);
nor U4354 (N_4354,N_3515,N_3600);
nor U4355 (N_4355,N_3294,N_3947);
or U4356 (N_4356,N_3635,N_3501);
and U4357 (N_4357,N_3537,N_3974);
nor U4358 (N_4358,N_3828,N_3873);
or U4359 (N_4359,N_3831,N_3573);
nand U4360 (N_4360,N_3524,N_3440);
xor U4361 (N_4361,N_3413,N_3132);
xor U4362 (N_4362,N_3717,N_3058);
or U4363 (N_4363,N_3748,N_3365);
nor U4364 (N_4364,N_3773,N_3779);
or U4365 (N_4365,N_3696,N_3156);
or U4366 (N_4366,N_3723,N_3741);
or U4367 (N_4367,N_3849,N_3864);
xnor U4368 (N_4368,N_3468,N_3091);
and U4369 (N_4369,N_3369,N_3028);
nand U4370 (N_4370,N_3095,N_3225);
or U4371 (N_4371,N_3545,N_3821);
and U4372 (N_4372,N_3529,N_3152);
or U4373 (N_4373,N_3742,N_3915);
xnor U4374 (N_4374,N_3326,N_3757);
xnor U4375 (N_4375,N_3990,N_3271);
xnor U4376 (N_4376,N_3754,N_3730);
and U4377 (N_4377,N_3557,N_3093);
xnor U4378 (N_4378,N_3694,N_3479);
and U4379 (N_4379,N_3448,N_3046);
and U4380 (N_4380,N_3358,N_3145);
nor U4381 (N_4381,N_3218,N_3734);
xnor U4382 (N_4382,N_3878,N_3895);
xnor U4383 (N_4383,N_3362,N_3268);
nor U4384 (N_4384,N_3582,N_3339);
xor U4385 (N_4385,N_3296,N_3938);
nand U4386 (N_4386,N_3601,N_3815);
nor U4387 (N_4387,N_3630,N_3559);
nor U4388 (N_4388,N_3009,N_3371);
xor U4389 (N_4389,N_3731,N_3987);
nor U4390 (N_4390,N_3405,N_3483);
xor U4391 (N_4391,N_3964,N_3771);
nand U4392 (N_4392,N_3373,N_3958);
nand U4393 (N_4393,N_3363,N_3162);
or U4394 (N_4394,N_3721,N_3765);
nand U4395 (N_4395,N_3106,N_3253);
xnor U4396 (N_4396,N_3695,N_3179);
nor U4397 (N_4397,N_3035,N_3477);
nor U4398 (N_4398,N_3982,N_3389);
and U4399 (N_4399,N_3548,N_3484);
or U4400 (N_4400,N_3304,N_3443);
nor U4401 (N_4401,N_3033,N_3059);
nor U4402 (N_4402,N_3536,N_3540);
and U4403 (N_4403,N_3660,N_3981);
or U4404 (N_4404,N_3119,N_3678);
xnor U4405 (N_4405,N_3881,N_3590);
nor U4406 (N_4406,N_3549,N_3804);
xor U4407 (N_4407,N_3626,N_3143);
nor U4408 (N_4408,N_3315,N_3146);
and U4409 (N_4409,N_3249,N_3232);
nor U4410 (N_4410,N_3689,N_3098);
nand U4411 (N_4411,N_3491,N_3472);
or U4412 (N_4412,N_3242,N_3243);
nor U4413 (N_4413,N_3076,N_3233);
or U4414 (N_4414,N_3786,N_3598);
xor U4415 (N_4415,N_3911,N_3313);
or U4416 (N_4416,N_3423,N_3613);
or U4417 (N_4417,N_3758,N_3932);
xnor U4418 (N_4418,N_3820,N_3738);
nor U4419 (N_4419,N_3518,N_3074);
and U4420 (N_4420,N_3276,N_3346);
xor U4421 (N_4421,N_3985,N_3569);
and U4422 (N_4422,N_3173,N_3813);
nand U4423 (N_4423,N_3564,N_3959);
and U4424 (N_4424,N_3610,N_3007);
nand U4425 (N_4425,N_3008,N_3342);
nand U4426 (N_4426,N_3047,N_3718);
and U4427 (N_4427,N_3984,N_3422);
nand U4428 (N_4428,N_3697,N_3228);
and U4429 (N_4429,N_3966,N_3673);
nor U4430 (N_4430,N_3254,N_3352);
or U4431 (N_4431,N_3056,N_3638);
nand U4432 (N_4432,N_3011,N_3805);
nor U4433 (N_4433,N_3768,N_3884);
xor U4434 (N_4434,N_3565,N_3650);
or U4435 (N_4435,N_3013,N_3510);
nand U4436 (N_4436,N_3488,N_3246);
nand U4437 (N_4437,N_3302,N_3618);
nand U4438 (N_4438,N_3523,N_3170);
nand U4439 (N_4439,N_3149,N_3291);
nor U4440 (N_4440,N_3359,N_3239);
xnor U4441 (N_4441,N_3447,N_3256);
xnor U4442 (N_4442,N_3522,N_3845);
and U4443 (N_4443,N_3006,N_3158);
or U4444 (N_4444,N_3803,N_3550);
or U4445 (N_4445,N_3002,N_3547);
or U4446 (N_4446,N_3102,N_3244);
nand U4447 (N_4447,N_3658,N_3048);
nand U4448 (N_4448,N_3057,N_3406);
and U4449 (N_4449,N_3357,N_3449);
or U4450 (N_4450,N_3427,N_3711);
and U4451 (N_4451,N_3043,N_3341);
and U4452 (N_4452,N_3850,N_3500);
nor U4453 (N_4453,N_3055,N_3551);
and U4454 (N_4454,N_3898,N_3117);
xnor U4455 (N_4455,N_3206,N_3234);
or U4456 (N_4456,N_3509,N_3680);
or U4457 (N_4457,N_3704,N_3101);
nor U4458 (N_4458,N_3307,N_3351);
and U4459 (N_4459,N_3124,N_3034);
nand U4460 (N_4460,N_3020,N_3372);
or U4461 (N_4461,N_3142,N_3411);
nor U4462 (N_4462,N_3562,N_3236);
nor U4463 (N_4463,N_3834,N_3759);
nand U4464 (N_4464,N_3951,N_3053);
nor U4465 (N_4465,N_3252,N_3592);
nor U4466 (N_4466,N_3627,N_3088);
xnor U4467 (N_4467,N_3402,N_3374);
xor U4468 (N_4468,N_3163,N_3669);
or U4469 (N_4469,N_3081,N_3442);
or U4470 (N_4470,N_3482,N_3801);
nand U4471 (N_4471,N_3498,N_3303);
xnor U4472 (N_4472,N_3970,N_3135);
xor U4473 (N_4473,N_3965,N_3874);
or U4474 (N_4474,N_3642,N_3108);
or U4475 (N_4475,N_3169,N_3543);
or U4476 (N_4476,N_3396,N_3676);
and U4477 (N_4477,N_3637,N_3077);
and U4478 (N_4478,N_3274,N_3004);
nor U4479 (N_4479,N_3000,N_3092);
or U4480 (N_4480,N_3602,N_3439);
or U4481 (N_4481,N_3761,N_3295);
nand U4482 (N_4482,N_3777,N_3793);
nand U4483 (N_4483,N_3230,N_3394);
xnor U4484 (N_4484,N_3069,N_3085);
and U4485 (N_4485,N_3393,N_3957);
nor U4486 (N_4486,N_3115,N_3266);
nor U4487 (N_4487,N_3324,N_3619);
xor U4488 (N_4488,N_3554,N_3876);
nand U4489 (N_4489,N_3822,N_3071);
nand U4490 (N_4490,N_3207,N_3579);
nand U4491 (N_4491,N_3588,N_3952);
and U4492 (N_4492,N_3776,N_3789);
nand U4493 (N_4493,N_3703,N_3513);
or U4494 (N_4494,N_3791,N_3212);
nand U4495 (N_4495,N_3655,N_3432);
and U4496 (N_4496,N_3316,N_3287);
nand U4497 (N_4497,N_3292,N_3039);
and U4498 (N_4498,N_3288,N_3114);
or U4499 (N_4499,N_3257,N_3318);
nand U4500 (N_4500,N_3888,N_3116);
xor U4501 (N_4501,N_3934,N_3598);
nor U4502 (N_4502,N_3202,N_3962);
xnor U4503 (N_4503,N_3658,N_3998);
xnor U4504 (N_4504,N_3398,N_3996);
and U4505 (N_4505,N_3626,N_3772);
nor U4506 (N_4506,N_3723,N_3574);
xnor U4507 (N_4507,N_3147,N_3857);
xnor U4508 (N_4508,N_3031,N_3556);
or U4509 (N_4509,N_3904,N_3254);
and U4510 (N_4510,N_3566,N_3264);
nor U4511 (N_4511,N_3884,N_3440);
xnor U4512 (N_4512,N_3090,N_3987);
and U4513 (N_4513,N_3538,N_3234);
xnor U4514 (N_4514,N_3347,N_3439);
or U4515 (N_4515,N_3706,N_3128);
or U4516 (N_4516,N_3004,N_3919);
and U4517 (N_4517,N_3796,N_3313);
xor U4518 (N_4518,N_3815,N_3809);
and U4519 (N_4519,N_3277,N_3906);
and U4520 (N_4520,N_3819,N_3402);
nor U4521 (N_4521,N_3017,N_3148);
nor U4522 (N_4522,N_3615,N_3677);
or U4523 (N_4523,N_3099,N_3271);
and U4524 (N_4524,N_3533,N_3017);
xor U4525 (N_4525,N_3546,N_3649);
and U4526 (N_4526,N_3750,N_3329);
nor U4527 (N_4527,N_3884,N_3172);
nand U4528 (N_4528,N_3587,N_3857);
xor U4529 (N_4529,N_3458,N_3891);
or U4530 (N_4530,N_3309,N_3747);
nor U4531 (N_4531,N_3864,N_3120);
and U4532 (N_4532,N_3011,N_3945);
nand U4533 (N_4533,N_3440,N_3742);
nand U4534 (N_4534,N_3971,N_3146);
xor U4535 (N_4535,N_3413,N_3618);
and U4536 (N_4536,N_3325,N_3061);
xnor U4537 (N_4537,N_3122,N_3941);
or U4538 (N_4538,N_3319,N_3700);
and U4539 (N_4539,N_3146,N_3180);
and U4540 (N_4540,N_3711,N_3709);
and U4541 (N_4541,N_3281,N_3146);
and U4542 (N_4542,N_3736,N_3491);
and U4543 (N_4543,N_3173,N_3682);
and U4544 (N_4544,N_3926,N_3228);
nand U4545 (N_4545,N_3481,N_3205);
nor U4546 (N_4546,N_3845,N_3707);
nor U4547 (N_4547,N_3567,N_3982);
xnor U4548 (N_4548,N_3302,N_3701);
and U4549 (N_4549,N_3958,N_3080);
nand U4550 (N_4550,N_3446,N_3046);
and U4551 (N_4551,N_3458,N_3564);
and U4552 (N_4552,N_3776,N_3786);
nand U4553 (N_4553,N_3969,N_3749);
nand U4554 (N_4554,N_3697,N_3890);
nor U4555 (N_4555,N_3244,N_3969);
nand U4556 (N_4556,N_3047,N_3144);
nand U4557 (N_4557,N_3672,N_3326);
nand U4558 (N_4558,N_3850,N_3465);
nand U4559 (N_4559,N_3589,N_3553);
xor U4560 (N_4560,N_3222,N_3283);
or U4561 (N_4561,N_3143,N_3662);
nand U4562 (N_4562,N_3866,N_3945);
and U4563 (N_4563,N_3412,N_3991);
xor U4564 (N_4564,N_3485,N_3337);
nor U4565 (N_4565,N_3292,N_3230);
nand U4566 (N_4566,N_3039,N_3508);
or U4567 (N_4567,N_3657,N_3814);
or U4568 (N_4568,N_3887,N_3467);
nor U4569 (N_4569,N_3315,N_3765);
or U4570 (N_4570,N_3844,N_3287);
nor U4571 (N_4571,N_3216,N_3624);
or U4572 (N_4572,N_3286,N_3072);
or U4573 (N_4573,N_3671,N_3949);
and U4574 (N_4574,N_3099,N_3831);
xor U4575 (N_4575,N_3308,N_3775);
and U4576 (N_4576,N_3898,N_3951);
and U4577 (N_4577,N_3192,N_3185);
xor U4578 (N_4578,N_3524,N_3730);
or U4579 (N_4579,N_3198,N_3680);
or U4580 (N_4580,N_3704,N_3842);
xnor U4581 (N_4581,N_3306,N_3065);
or U4582 (N_4582,N_3624,N_3059);
nand U4583 (N_4583,N_3845,N_3230);
nand U4584 (N_4584,N_3742,N_3167);
nor U4585 (N_4585,N_3998,N_3396);
and U4586 (N_4586,N_3372,N_3237);
or U4587 (N_4587,N_3397,N_3120);
nand U4588 (N_4588,N_3560,N_3844);
xnor U4589 (N_4589,N_3416,N_3246);
or U4590 (N_4590,N_3059,N_3034);
and U4591 (N_4591,N_3463,N_3424);
or U4592 (N_4592,N_3127,N_3490);
nor U4593 (N_4593,N_3110,N_3221);
nor U4594 (N_4594,N_3067,N_3865);
nand U4595 (N_4595,N_3301,N_3827);
nand U4596 (N_4596,N_3187,N_3029);
or U4597 (N_4597,N_3823,N_3984);
or U4598 (N_4598,N_3233,N_3801);
and U4599 (N_4599,N_3518,N_3316);
nand U4600 (N_4600,N_3477,N_3295);
xor U4601 (N_4601,N_3440,N_3913);
nand U4602 (N_4602,N_3449,N_3049);
xnor U4603 (N_4603,N_3095,N_3002);
or U4604 (N_4604,N_3335,N_3978);
xnor U4605 (N_4605,N_3722,N_3136);
nand U4606 (N_4606,N_3888,N_3726);
nand U4607 (N_4607,N_3727,N_3883);
xnor U4608 (N_4608,N_3198,N_3934);
nand U4609 (N_4609,N_3734,N_3792);
and U4610 (N_4610,N_3652,N_3438);
nand U4611 (N_4611,N_3922,N_3309);
nand U4612 (N_4612,N_3818,N_3334);
and U4613 (N_4613,N_3534,N_3430);
nor U4614 (N_4614,N_3830,N_3332);
xor U4615 (N_4615,N_3998,N_3325);
or U4616 (N_4616,N_3237,N_3730);
xnor U4617 (N_4617,N_3293,N_3539);
and U4618 (N_4618,N_3527,N_3174);
or U4619 (N_4619,N_3767,N_3717);
or U4620 (N_4620,N_3209,N_3311);
nor U4621 (N_4621,N_3140,N_3591);
nand U4622 (N_4622,N_3184,N_3872);
and U4623 (N_4623,N_3961,N_3616);
xor U4624 (N_4624,N_3948,N_3503);
and U4625 (N_4625,N_3949,N_3693);
and U4626 (N_4626,N_3111,N_3856);
xnor U4627 (N_4627,N_3675,N_3256);
or U4628 (N_4628,N_3009,N_3883);
xor U4629 (N_4629,N_3488,N_3294);
nor U4630 (N_4630,N_3803,N_3047);
xnor U4631 (N_4631,N_3981,N_3441);
xnor U4632 (N_4632,N_3469,N_3877);
and U4633 (N_4633,N_3508,N_3693);
nor U4634 (N_4634,N_3604,N_3788);
or U4635 (N_4635,N_3359,N_3410);
xor U4636 (N_4636,N_3093,N_3967);
and U4637 (N_4637,N_3239,N_3073);
nand U4638 (N_4638,N_3627,N_3146);
nand U4639 (N_4639,N_3851,N_3199);
xor U4640 (N_4640,N_3076,N_3238);
xor U4641 (N_4641,N_3824,N_3829);
nor U4642 (N_4642,N_3012,N_3776);
xnor U4643 (N_4643,N_3605,N_3391);
and U4644 (N_4644,N_3106,N_3302);
or U4645 (N_4645,N_3596,N_3280);
or U4646 (N_4646,N_3470,N_3107);
nor U4647 (N_4647,N_3873,N_3505);
nand U4648 (N_4648,N_3749,N_3409);
nor U4649 (N_4649,N_3002,N_3294);
or U4650 (N_4650,N_3860,N_3402);
or U4651 (N_4651,N_3134,N_3674);
or U4652 (N_4652,N_3727,N_3744);
xnor U4653 (N_4653,N_3946,N_3641);
nand U4654 (N_4654,N_3893,N_3315);
nand U4655 (N_4655,N_3997,N_3357);
and U4656 (N_4656,N_3847,N_3602);
nand U4657 (N_4657,N_3106,N_3455);
xor U4658 (N_4658,N_3301,N_3772);
nor U4659 (N_4659,N_3620,N_3140);
and U4660 (N_4660,N_3615,N_3608);
xnor U4661 (N_4661,N_3217,N_3347);
and U4662 (N_4662,N_3420,N_3449);
and U4663 (N_4663,N_3099,N_3636);
xnor U4664 (N_4664,N_3898,N_3665);
nor U4665 (N_4665,N_3210,N_3953);
or U4666 (N_4666,N_3324,N_3609);
and U4667 (N_4667,N_3342,N_3370);
xnor U4668 (N_4668,N_3743,N_3302);
and U4669 (N_4669,N_3114,N_3883);
and U4670 (N_4670,N_3147,N_3368);
or U4671 (N_4671,N_3454,N_3698);
xor U4672 (N_4672,N_3548,N_3824);
and U4673 (N_4673,N_3127,N_3253);
nand U4674 (N_4674,N_3947,N_3093);
nand U4675 (N_4675,N_3693,N_3003);
nor U4676 (N_4676,N_3199,N_3305);
and U4677 (N_4677,N_3804,N_3622);
and U4678 (N_4678,N_3070,N_3019);
or U4679 (N_4679,N_3618,N_3010);
xnor U4680 (N_4680,N_3289,N_3657);
nor U4681 (N_4681,N_3287,N_3377);
and U4682 (N_4682,N_3103,N_3437);
or U4683 (N_4683,N_3465,N_3348);
xnor U4684 (N_4684,N_3771,N_3584);
and U4685 (N_4685,N_3273,N_3742);
or U4686 (N_4686,N_3788,N_3419);
and U4687 (N_4687,N_3983,N_3353);
and U4688 (N_4688,N_3546,N_3400);
and U4689 (N_4689,N_3647,N_3763);
and U4690 (N_4690,N_3395,N_3092);
nor U4691 (N_4691,N_3842,N_3808);
nand U4692 (N_4692,N_3464,N_3975);
or U4693 (N_4693,N_3256,N_3017);
xor U4694 (N_4694,N_3666,N_3496);
or U4695 (N_4695,N_3843,N_3681);
nor U4696 (N_4696,N_3345,N_3892);
xnor U4697 (N_4697,N_3879,N_3255);
nor U4698 (N_4698,N_3581,N_3835);
nand U4699 (N_4699,N_3264,N_3738);
nand U4700 (N_4700,N_3256,N_3789);
nor U4701 (N_4701,N_3825,N_3640);
nand U4702 (N_4702,N_3228,N_3918);
nand U4703 (N_4703,N_3417,N_3051);
xnor U4704 (N_4704,N_3005,N_3539);
and U4705 (N_4705,N_3389,N_3814);
nand U4706 (N_4706,N_3819,N_3721);
nand U4707 (N_4707,N_3877,N_3890);
and U4708 (N_4708,N_3942,N_3269);
or U4709 (N_4709,N_3280,N_3814);
nor U4710 (N_4710,N_3560,N_3765);
and U4711 (N_4711,N_3317,N_3608);
nor U4712 (N_4712,N_3618,N_3679);
or U4713 (N_4713,N_3764,N_3725);
and U4714 (N_4714,N_3169,N_3861);
nor U4715 (N_4715,N_3453,N_3105);
nand U4716 (N_4716,N_3714,N_3839);
xnor U4717 (N_4717,N_3586,N_3742);
nand U4718 (N_4718,N_3302,N_3206);
or U4719 (N_4719,N_3124,N_3161);
and U4720 (N_4720,N_3209,N_3720);
nor U4721 (N_4721,N_3997,N_3370);
or U4722 (N_4722,N_3944,N_3861);
or U4723 (N_4723,N_3814,N_3855);
and U4724 (N_4724,N_3195,N_3625);
xnor U4725 (N_4725,N_3395,N_3171);
xor U4726 (N_4726,N_3465,N_3291);
nor U4727 (N_4727,N_3254,N_3512);
and U4728 (N_4728,N_3903,N_3057);
xnor U4729 (N_4729,N_3161,N_3138);
nand U4730 (N_4730,N_3939,N_3464);
nor U4731 (N_4731,N_3113,N_3229);
xor U4732 (N_4732,N_3970,N_3439);
or U4733 (N_4733,N_3430,N_3982);
xnor U4734 (N_4734,N_3076,N_3720);
xnor U4735 (N_4735,N_3298,N_3157);
and U4736 (N_4736,N_3201,N_3054);
nand U4737 (N_4737,N_3664,N_3410);
nor U4738 (N_4738,N_3754,N_3565);
and U4739 (N_4739,N_3217,N_3256);
or U4740 (N_4740,N_3906,N_3898);
xor U4741 (N_4741,N_3651,N_3474);
and U4742 (N_4742,N_3326,N_3014);
xnor U4743 (N_4743,N_3617,N_3206);
and U4744 (N_4744,N_3798,N_3079);
xor U4745 (N_4745,N_3516,N_3015);
nor U4746 (N_4746,N_3691,N_3431);
nor U4747 (N_4747,N_3368,N_3845);
and U4748 (N_4748,N_3002,N_3290);
and U4749 (N_4749,N_3447,N_3569);
nand U4750 (N_4750,N_3612,N_3873);
xor U4751 (N_4751,N_3261,N_3762);
nor U4752 (N_4752,N_3571,N_3689);
nor U4753 (N_4753,N_3571,N_3838);
nand U4754 (N_4754,N_3098,N_3945);
and U4755 (N_4755,N_3186,N_3437);
xnor U4756 (N_4756,N_3613,N_3920);
or U4757 (N_4757,N_3194,N_3193);
and U4758 (N_4758,N_3490,N_3312);
xor U4759 (N_4759,N_3313,N_3391);
or U4760 (N_4760,N_3540,N_3469);
xor U4761 (N_4761,N_3455,N_3777);
and U4762 (N_4762,N_3307,N_3718);
or U4763 (N_4763,N_3376,N_3463);
xor U4764 (N_4764,N_3106,N_3371);
nor U4765 (N_4765,N_3139,N_3896);
and U4766 (N_4766,N_3903,N_3370);
nand U4767 (N_4767,N_3625,N_3005);
or U4768 (N_4768,N_3069,N_3582);
or U4769 (N_4769,N_3528,N_3177);
or U4770 (N_4770,N_3306,N_3327);
and U4771 (N_4771,N_3468,N_3590);
nand U4772 (N_4772,N_3596,N_3464);
xnor U4773 (N_4773,N_3484,N_3373);
nand U4774 (N_4774,N_3201,N_3444);
xor U4775 (N_4775,N_3408,N_3091);
or U4776 (N_4776,N_3333,N_3899);
and U4777 (N_4777,N_3269,N_3288);
nor U4778 (N_4778,N_3499,N_3090);
xnor U4779 (N_4779,N_3935,N_3780);
nor U4780 (N_4780,N_3679,N_3380);
and U4781 (N_4781,N_3722,N_3361);
xnor U4782 (N_4782,N_3168,N_3986);
or U4783 (N_4783,N_3792,N_3541);
xnor U4784 (N_4784,N_3896,N_3539);
nand U4785 (N_4785,N_3016,N_3472);
xnor U4786 (N_4786,N_3283,N_3590);
nand U4787 (N_4787,N_3394,N_3757);
or U4788 (N_4788,N_3353,N_3940);
nand U4789 (N_4789,N_3282,N_3333);
nor U4790 (N_4790,N_3015,N_3504);
and U4791 (N_4791,N_3551,N_3274);
or U4792 (N_4792,N_3882,N_3683);
xnor U4793 (N_4793,N_3550,N_3576);
nor U4794 (N_4794,N_3875,N_3039);
xnor U4795 (N_4795,N_3112,N_3833);
and U4796 (N_4796,N_3100,N_3140);
or U4797 (N_4797,N_3155,N_3430);
nand U4798 (N_4798,N_3044,N_3229);
or U4799 (N_4799,N_3936,N_3602);
nor U4800 (N_4800,N_3771,N_3750);
or U4801 (N_4801,N_3411,N_3408);
or U4802 (N_4802,N_3743,N_3644);
nand U4803 (N_4803,N_3819,N_3332);
nand U4804 (N_4804,N_3813,N_3733);
and U4805 (N_4805,N_3081,N_3974);
nor U4806 (N_4806,N_3602,N_3394);
or U4807 (N_4807,N_3988,N_3954);
xor U4808 (N_4808,N_3584,N_3926);
or U4809 (N_4809,N_3475,N_3399);
or U4810 (N_4810,N_3203,N_3321);
and U4811 (N_4811,N_3814,N_3759);
and U4812 (N_4812,N_3679,N_3757);
or U4813 (N_4813,N_3720,N_3728);
nor U4814 (N_4814,N_3845,N_3066);
nand U4815 (N_4815,N_3731,N_3895);
or U4816 (N_4816,N_3237,N_3960);
nor U4817 (N_4817,N_3530,N_3949);
nand U4818 (N_4818,N_3509,N_3639);
or U4819 (N_4819,N_3881,N_3915);
nor U4820 (N_4820,N_3133,N_3018);
xor U4821 (N_4821,N_3312,N_3894);
nor U4822 (N_4822,N_3969,N_3647);
and U4823 (N_4823,N_3734,N_3393);
xnor U4824 (N_4824,N_3403,N_3768);
nor U4825 (N_4825,N_3086,N_3255);
or U4826 (N_4826,N_3146,N_3787);
or U4827 (N_4827,N_3455,N_3493);
nor U4828 (N_4828,N_3191,N_3403);
nor U4829 (N_4829,N_3579,N_3391);
or U4830 (N_4830,N_3637,N_3131);
or U4831 (N_4831,N_3389,N_3026);
xnor U4832 (N_4832,N_3280,N_3056);
or U4833 (N_4833,N_3512,N_3738);
nand U4834 (N_4834,N_3674,N_3837);
nor U4835 (N_4835,N_3148,N_3130);
nand U4836 (N_4836,N_3158,N_3462);
or U4837 (N_4837,N_3403,N_3778);
and U4838 (N_4838,N_3575,N_3408);
nor U4839 (N_4839,N_3814,N_3916);
nand U4840 (N_4840,N_3637,N_3495);
and U4841 (N_4841,N_3015,N_3920);
and U4842 (N_4842,N_3926,N_3190);
nor U4843 (N_4843,N_3922,N_3663);
and U4844 (N_4844,N_3618,N_3889);
xnor U4845 (N_4845,N_3195,N_3225);
and U4846 (N_4846,N_3181,N_3616);
nor U4847 (N_4847,N_3965,N_3470);
or U4848 (N_4848,N_3526,N_3265);
nand U4849 (N_4849,N_3787,N_3817);
and U4850 (N_4850,N_3984,N_3016);
xnor U4851 (N_4851,N_3820,N_3055);
or U4852 (N_4852,N_3095,N_3142);
xnor U4853 (N_4853,N_3304,N_3689);
nand U4854 (N_4854,N_3806,N_3544);
or U4855 (N_4855,N_3781,N_3954);
or U4856 (N_4856,N_3168,N_3514);
or U4857 (N_4857,N_3115,N_3051);
or U4858 (N_4858,N_3956,N_3926);
nor U4859 (N_4859,N_3780,N_3510);
nand U4860 (N_4860,N_3552,N_3233);
or U4861 (N_4861,N_3316,N_3588);
nand U4862 (N_4862,N_3734,N_3656);
xnor U4863 (N_4863,N_3174,N_3639);
xor U4864 (N_4864,N_3333,N_3956);
nand U4865 (N_4865,N_3032,N_3735);
and U4866 (N_4866,N_3074,N_3825);
or U4867 (N_4867,N_3379,N_3307);
nand U4868 (N_4868,N_3576,N_3756);
nand U4869 (N_4869,N_3339,N_3824);
and U4870 (N_4870,N_3500,N_3512);
or U4871 (N_4871,N_3767,N_3262);
xnor U4872 (N_4872,N_3142,N_3491);
and U4873 (N_4873,N_3837,N_3893);
nand U4874 (N_4874,N_3614,N_3812);
nand U4875 (N_4875,N_3480,N_3578);
or U4876 (N_4876,N_3742,N_3329);
nor U4877 (N_4877,N_3338,N_3677);
nand U4878 (N_4878,N_3663,N_3120);
nor U4879 (N_4879,N_3734,N_3507);
nand U4880 (N_4880,N_3994,N_3403);
xnor U4881 (N_4881,N_3217,N_3353);
or U4882 (N_4882,N_3159,N_3315);
nor U4883 (N_4883,N_3501,N_3943);
xnor U4884 (N_4884,N_3824,N_3742);
or U4885 (N_4885,N_3503,N_3017);
and U4886 (N_4886,N_3690,N_3942);
or U4887 (N_4887,N_3781,N_3665);
xor U4888 (N_4888,N_3326,N_3046);
or U4889 (N_4889,N_3436,N_3885);
or U4890 (N_4890,N_3927,N_3122);
and U4891 (N_4891,N_3711,N_3626);
nand U4892 (N_4892,N_3980,N_3358);
and U4893 (N_4893,N_3100,N_3767);
xnor U4894 (N_4894,N_3307,N_3375);
and U4895 (N_4895,N_3281,N_3777);
xnor U4896 (N_4896,N_3858,N_3242);
or U4897 (N_4897,N_3449,N_3859);
and U4898 (N_4898,N_3197,N_3454);
and U4899 (N_4899,N_3759,N_3235);
and U4900 (N_4900,N_3717,N_3830);
nor U4901 (N_4901,N_3250,N_3769);
nor U4902 (N_4902,N_3544,N_3366);
xor U4903 (N_4903,N_3309,N_3338);
xnor U4904 (N_4904,N_3653,N_3929);
or U4905 (N_4905,N_3812,N_3297);
nand U4906 (N_4906,N_3010,N_3763);
nor U4907 (N_4907,N_3891,N_3561);
or U4908 (N_4908,N_3306,N_3254);
nor U4909 (N_4909,N_3237,N_3755);
nand U4910 (N_4910,N_3987,N_3464);
or U4911 (N_4911,N_3507,N_3636);
nor U4912 (N_4912,N_3749,N_3952);
and U4913 (N_4913,N_3387,N_3426);
and U4914 (N_4914,N_3528,N_3731);
or U4915 (N_4915,N_3547,N_3538);
and U4916 (N_4916,N_3215,N_3182);
and U4917 (N_4917,N_3211,N_3340);
xnor U4918 (N_4918,N_3224,N_3778);
xnor U4919 (N_4919,N_3372,N_3813);
or U4920 (N_4920,N_3895,N_3255);
xor U4921 (N_4921,N_3476,N_3215);
nand U4922 (N_4922,N_3977,N_3762);
xnor U4923 (N_4923,N_3758,N_3334);
nor U4924 (N_4924,N_3709,N_3744);
and U4925 (N_4925,N_3162,N_3569);
nand U4926 (N_4926,N_3199,N_3646);
nand U4927 (N_4927,N_3749,N_3660);
nor U4928 (N_4928,N_3174,N_3086);
and U4929 (N_4929,N_3311,N_3107);
nand U4930 (N_4930,N_3720,N_3404);
xor U4931 (N_4931,N_3379,N_3858);
xnor U4932 (N_4932,N_3346,N_3655);
nor U4933 (N_4933,N_3894,N_3151);
and U4934 (N_4934,N_3796,N_3001);
nand U4935 (N_4935,N_3988,N_3192);
and U4936 (N_4936,N_3085,N_3794);
nor U4937 (N_4937,N_3160,N_3176);
nand U4938 (N_4938,N_3269,N_3072);
nor U4939 (N_4939,N_3410,N_3291);
xnor U4940 (N_4940,N_3973,N_3469);
or U4941 (N_4941,N_3792,N_3344);
nand U4942 (N_4942,N_3423,N_3752);
xor U4943 (N_4943,N_3761,N_3427);
nand U4944 (N_4944,N_3047,N_3320);
and U4945 (N_4945,N_3706,N_3065);
nor U4946 (N_4946,N_3542,N_3816);
or U4947 (N_4947,N_3886,N_3891);
and U4948 (N_4948,N_3525,N_3180);
nor U4949 (N_4949,N_3105,N_3389);
nand U4950 (N_4950,N_3547,N_3562);
or U4951 (N_4951,N_3909,N_3978);
xor U4952 (N_4952,N_3413,N_3293);
or U4953 (N_4953,N_3715,N_3348);
nand U4954 (N_4954,N_3543,N_3646);
xnor U4955 (N_4955,N_3204,N_3022);
nor U4956 (N_4956,N_3449,N_3040);
and U4957 (N_4957,N_3951,N_3112);
or U4958 (N_4958,N_3808,N_3356);
xor U4959 (N_4959,N_3298,N_3460);
or U4960 (N_4960,N_3279,N_3479);
xor U4961 (N_4961,N_3329,N_3972);
or U4962 (N_4962,N_3634,N_3791);
nor U4963 (N_4963,N_3477,N_3927);
and U4964 (N_4964,N_3605,N_3284);
xor U4965 (N_4965,N_3587,N_3674);
xor U4966 (N_4966,N_3420,N_3743);
nor U4967 (N_4967,N_3338,N_3446);
or U4968 (N_4968,N_3221,N_3443);
or U4969 (N_4969,N_3386,N_3301);
and U4970 (N_4970,N_3787,N_3136);
xnor U4971 (N_4971,N_3284,N_3576);
xor U4972 (N_4972,N_3172,N_3609);
and U4973 (N_4973,N_3407,N_3919);
or U4974 (N_4974,N_3747,N_3375);
or U4975 (N_4975,N_3846,N_3652);
or U4976 (N_4976,N_3172,N_3638);
or U4977 (N_4977,N_3465,N_3679);
nor U4978 (N_4978,N_3698,N_3051);
nor U4979 (N_4979,N_3943,N_3472);
and U4980 (N_4980,N_3629,N_3304);
nor U4981 (N_4981,N_3303,N_3578);
xor U4982 (N_4982,N_3253,N_3450);
nand U4983 (N_4983,N_3332,N_3507);
or U4984 (N_4984,N_3756,N_3547);
nor U4985 (N_4985,N_3608,N_3602);
or U4986 (N_4986,N_3264,N_3365);
xor U4987 (N_4987,N_3788,N_3875);
nor U4988 (N_4988,N_3743,N_3173);
nor U4989 (N_4989,N_3321,N_3221);
or U4990 (N_4990,N_3422,N_3432);
or U4991 (N_4991,N_3504,N_3579);
xor U4992 (N_4992,N_3932,N_3154);
or U4993 (N_4993,N_3369,N_3725);
and U4994 (N_4994,N_3661,N_3168);
and U4995 (N_4995,N_3796,N_3732);
nor U4996 (N_4996,N_3708,N_3032);
or U4997 (N_4997,N_3597,N_3606);
or U4998 (N_4998,N_3440,N_3719);
xor U4999 (N_4999,N_3669,N_3592);
nor U5000 (N_5000,N_4308,N_4678);
xor U5001 (N_5001,N_4756,N_4215);
nor U5002 (N_5002,N_4398,N_4371);
xor U5003 (N_5003,N_4151,N_4345);
xnor U5004 (N_5004,N_4214,N_4944);
nor U5005 (N_5005,N_4180,N_4951);
nor U5006 (N_5006,N_4941,N_4010);
nand U5007 (N_5007,N_4240,N_4652);
nor U5008 (N_5008,N_4685,N_4131);
nor U5009 (N_5009,N_4182,N_4707);
and U5010 (N_5010,N_4419,N_4616);
and U5011 (N_5011,N_4237,N_4936);
or U5012 (N_5012,N_4093,N_4114);
nand U5013 (N_5013,N_4681,N_4003);
and U5014 (N_5014,N_4925,N_4055);
and U5015 (N_5015,N_4692,N_4425);
or U5016 (N_5016,N_4648,N_4897);
nand U5017 (N_5017,N_4289,N_4689);
or U5018 (N_5018,N_4317,N_4909);
nand U5019 (N_5019,N_4919,N_4447);
or U5020 (N_5020,N_4736,N_4143);
nand U5021 (N_5021,N_4133,N_4943);
nand U5022 (N_5022,N_4097,N_4588);
nor U5023 (N_5023,N_4474,N_4778);
nand U5024 (N_5024,N_4859,N_4987);
xnor U5025 (N_5025,N_4416,N_4740);
nand U5026 (N_5026,N_4406,N_4193);
xor U5027 (N_5027,N_4091,N_4614);
xor U5028 (N_5028,N_4053,N_4263);
nor U5029 (N_5029,N_4785,N_4860);
and U5030 (N_5030,N_4570,N_4499);
and U5031 (N_5031,N_4157,N_4332);
xor U5032 (N_5032,N_4280,N_4620);
nand U5033 (N_5033,N_4683,N_4144);
or U5034 (N_5034,N_4049,N_4099);
xnor U5035 (N_5035,N_4664,N_4449);
nor U5036 (N_5036,N_4950,N_4278);
nand U5037 (N_5037,N_4883,N_4313);
and U5038 (N_5038,N_4195,N_4154);
nand U5039 (N_5039,N_4495,N_4241);
and U5040 (N_5040,N_4621,N_4380);
and U5041 (N_5041,N_4760,N_4394);
and U5042 (N_5042,N_4567,N_4513);
xnor U5043 (N_5043,N_4617,N_4748);
or U5044 (N_5044,N_4638,N_4797);
and U5045 (N_5045,N_4119,N_4532);
or U5046 (N_5046,N_4338,N_4754);
nand U5047 (N_5047,N_4389,N_4693);
nor U5048 (N_5048,N_4908,N_4983);
or U5049 (N_5049,N_4939,N_4346);
xnor U5050 (N_5050,N_4159,N_4695);
nor U5051 (N_5051,N_4690,N_4836);
xor U5052 (N_5052,N_4098,N_4731);
nand U5053 (N_5053,N_4603,N_4976);
nand U5054 (N_5054,N_4312,N_4018);
nand U5055 (N_5055,N_4965,N_4669);
nor U5056 (N_5056,N_4155,N_4629);
and U5057 (N_5057,N_4032,N_4789);
and U5058 (N_5058,N_4675,N_4439);
or U5059 (N_5059,N_4888,N_4556);
and U5060 (N_5060,N_4504,N_4927);
nor U5061 (N_5061,N_4990,N_4014);
and U5062 (N_5062,N_4569,N_4016);
or U5063 (N_5063,N_4382,N_4628);
and U5064 (N_5064,N_4937,N_4135);
nor U5065 (N_5065,N_4732,N_4478);
xnor U5066 (N_5066,N_4694,N_4030);
and U5067 (N_5067,N_4720,N_4526);
or U5068 (N_5068,N_4670,N_4839);
nor U5069 (N_5069,N_4121,N_4814);
and U5070 (N_5070,N_4080,N_4101);
and U5071 (N_5071,N_4079,N_4216);
xnor U5072 (N_5072,N_4552,N_4626);
nand U5073 (N_5073,N_4776,N_4706);
nand U5074 (N_5074,N_4051,N_4535);
or U5075 (N_5075,N_4833,N_4691);
nand U5076 (N_5076,N_4120,N_4213);
nand U5077 (N_5077,N_4541,N_4273);
xor U5078 (N_5078,N_4550,N_4687);
nor U5079 (N_5079,N_4048,N_4129);
and U5080 (N_5080,N_4077,N_4660);
nor U5081 (N_5081,N_4333,N_4647);
xnor U5082 (N_5082,N_4530,N_4744);
and U5083 (N_5083,N_4822,N_4282);
nor U5084 (N_5084,N_4243,N_4701);
or U5085 (N_5085,N_4301,N_4659);
or U5086 (N_5086,N_4974,N_4715);
xor U5087 (N_5087,N_4635,N_4519);
nand U5088 (N_5088,N_4221,N_4432);
and U5089 (N_5089,N_4633,N_4174);
nor U5090 (N_5090,N_4654,N_4445);
nor U5091 (N_5091,N_4892,N_4370);
and U5092 (N_5092,N_4971,N_4163);
nor U5093 (N_5093,N_4323,N_4254);
or U5094 (N_5094,N_4733,N_4434);
and U5095 (N_5095,N_4959,N_4881);
or U5096 (N_5096,N_4742,N_4094);
and U5097 (N_5097,N_4999,N_4085);
xor U5098 (N_5098,N_4074,N_4817);
and U5099 (N_5099,N_4463,N_4642);
nor U5100 (N_5100,N_4782,N_4476);
nor U5101 (N_5101,N_4090,N_4824);
or U5102 (N_5102,N_4341,N_4861);
nand U5103 (N_5103,N_4327,N_4029);
or U5104 (N_5104,N_4725,N_4220);
and U5105 (N_5105,N_4103,N_4870);
and U5106 (N_5106,N_4108,N_4853);
xnor U5107 (N_5107,N_4525,N_4140);
nand U5108 (N_5108,N_4441,N_4735);
nand U5109 (N_5109,N_4516,N_4855);
and U5110 (N_5110,N_4679,N_4605);
and U5111 (N_5111,N_4915,N_4466);
or U5112 (N_5112,N_4258,N_4876);
and U5113 (N_5113,N_4724,N_4995);
nor U5114 (N_5114,N_4973,N_4739);
or U5115 (N_5115,N_4928,N_4623);
and U5116 (N_5116,N_4649,N_4627);
and U5117 (N_5117,N_4890,N_4835);
nor U5118 (N_5118,N_4012,N_4661);
nor U5119 (N_5119,N_4208,N_4092);
and U5120 (N_5120,N_4775,N_4767);
and U5121 (N_5121,N_4104,N_4584);
nand U5122 (N_5122,N_4038,N_4385);
xor U5123 (N_5123,N_4339,N_4217);
nand U5124 (N_5124,N_4684,N_4460);
or U5125 (N_5125,N_4127,N_4230);
nor U5126 (N_5126,N_4065,N_4819);
nor U5127 (N_5127,N_4381,N_4363);
or U5128 (N_5128,N_4924,N_4710);
nand U5129 (N_5129,N_4297,N_4471);
and U5130 (N_5130,N_4811,N_4395);
nand U5131 (N_5131,N_4904,N_4305);
or U5132 (N_5132,N_4089,N_4004);
xor U5133 (N_5133,N_4063,N_4162);
xor U5134 (N_5134,N_4444,N_4877);
nor U5135 (N_5135,N_4873,N_4458);
nand U5136 (N_5136,N_4759,N_4968);
and U5137 (N_5137,N_4268,N_4429);
xnor U5138 (N_5138,N_4290,N_4329);
and U5139 (N_5139,N_4576,N_4536);
and U5140 (N_5140,N_4910,N_4231);
nor U5141 (N_5141,N_4862,N_4618);
and U5142 (N_5142,N_4490,N_4244);
or U5143 (N_5143,N_4437,N_4544);
nand U5144 (N_5144,N_4422,N_4421);
and U5145 (N_5145,N_4903,N_4795);
or U5146 (N_5146,N_4637,N_4052);
nor U5147 (N_5147,N_4028,N_4455);
nor U5148 (N_5148,N_4820,N_4565);
nor U5149 (N_5149,N_4579,N_4377);
nand U5150 (N_5150,N_4431,N_4543);
nor U5151 (N_5151,N_4413,N_4967);
or U5152 (N_5152,N_4269,N_4804);
nand U5153 (N_5153,N_4537,N_4520);
or U5154 (N_5154,N_4325,N_4547);
and U5155 (N_5155,N_4790,N_4082);
xor U5156 (N_5156,N_4879,N_4171);
xor U5157 (N_5157,N_4600,N_4505);
or U5158 (N_5158,N_4450,N_4435);
nor U5159 (N_5159,N_4362,N_4858);
xnor U5160 (N_5160,N_4949,N_4923);
or U5161 (N_5161,N_4124,N_4643);
nand U5162 (N_5162,N_4470,N_4916);
nor U5163 (N_5163,N_4354,N_4777);
nand U5164 (N_5164,N_4272,N_4271);
nor U5165 (N_5165,N_4752,N_4769);
xnor U5166 (N_5166,N_4891,N_4930);
xor U5167 (N_5167,N_4745,N_4189);
nor U5168 (N_5168,N_4008,N_4299);
nand U5169 (N_5169,N_4266,N_4938);
nand U5170 (N_5170,N_4662,N_4319);
or U5171 (N_5171,N_4947,N_4986);
xor U5172 (N_5172,N_4946,N_4111);
and U5173 (N_5173,N_4674,N_4364);
nor U5174 (N_5174,N_4815,N_4728);
or U5175 (N_5175,N_4225,N_4264);
or U5176 (N_5176,N_4061,N_4784);
and U5177 (N_5177,N_4962,N_4798);
nand U5178 (N_5178,N_4456,N_4146);
nor U5179 (N_5179,N_4210,N_4343);
nand U5180 (N_5180,N_4911,N_4414);
and U5181 (N_5181,N_4601,N_4071);
nor U5182 (N_5182,N_4717,N_4852);
xor U5183 (N_5183,N_4296,N_4658);
or U5184 (N_5184,N_4042,N_4806);
nor U5185 (N_5185,N_4229,N_4046);
xor U5186 (N_5186,N_4430,N_4467);
nor U5187 (N_5187,N_4730,N_4178);
xnor U5188 (N_5188,N_4459,N_4084);
nor U5189 (N_5189,N_4529,N_4595);
nand U5190 (N_5190,N_4843,N_4921);
nand U5191 (N_5191,N_4677,N_4125);
xnor U5192 (N_5192,N_4578,N_4043);
xnor U5193 (N_5193,N_4224,N_4024);
nor U5194 (N_5194,N_4375,N_4598);
xnor U5195 (N_5195,N_4534,N_4391);
and U5196 (N_5196,N_4761,N_4792);
xnor U5197 (N_5197,N_4703,N_4992);
xor U5198 (N_5198,N_4234,N_4436);
or U5199 (N_5199,N_4321,N_4743);
xor U5200 (N_5200,N_4615,N_4123);
or U5201 (N_5201,N_4270,N_4207);
nand U5202 (N_5202,N_4166,N_4517);
nor U5203 (N_5203,N_4013,N_4383);
nor U5204 (N_5204,N_4580,N_4204);
nor U5205 (N_5205,N_4871,N_4068);
or U5206 (N_5206,N_4095,N_4137);
nand U5207 (N_5207,N_4233,N_4945);
nand U5208 (N_5208,N_4136,N_4002);
xnor U5209 (N_5209,N_4287,N_4011);
nor U5210 (N_5210,N_4842,N_4747);
nor U5211 (N_5211,N_4186,N_4110);
nand U5212 (N_5212,N_4845,N_4575);
and U5213 (N_5213,N_4036,N_4373);
and U5214 (N_5214,N_4105,N_4320);
xnor U5215 (N_5215,N_4721,N_4175);
nand U5216 (N_5216,N_4850,N_4359);
xnor U5217 (N_5217,N_4064,N_4005);
nand U5218 (N_5218,N_4676,N_4286);
nand U5219 (N_5219,N_4538,N_4086);
and U5220 (N_5220,N_4347,N_4274);
or U5221 (N_5221,N_4599,N_4737);
and U5222 (N_5222,N_4001,N_4582);
xor U5223 (N_5223,N_4961,N_4172);
nor U5224 (N_5224,N_4865,N_4956);
xnor U5225 (N_5225,N_4666,N_4142);
xor U5226 (N_5226,N_4893,N_4403);
xnor U5227 (N_5227,N_4348,N_4112);
or U5228 (N_5228,N_4610,N_4293);
nand U5229 (N_5229,N_4462,N_4920);
or U5230 (N_5230,N_4540,N_4411);
xor U5231 (N_5231,N_4118,N_4738);
nor U5232 (N_5232,N_4295,N_4896);
xor U5233 (N_5233,N_4805,N_4276);
nor U5234 (N_5234,N_4613,N_4807);
and U5235 (N_5235,N_4966,N_4846);
or U5236 (N_5236,N_4727,N_4746);
nor U5237 (N_5237,N_4309,N_4275);
or U5238 (N_5238,N_4755,N_4070);
and U5239 (N_5239,N_4557,N_4699);
xor U5240 (N_5240,N_4197,N_4590);
and U5241 (N_5241,N_4050,N_4841);
xnor U5242 (N_5242,N_4250,N_4181);
nor U5243 (N_5243,N_4889,N_4404);
or U5244 (N_5244,N_4772,N_4205);
or U5245 (N_5245,N_4632,N_4485);
xnor U5246 (N_5246,N_4672,N_4196);
and U5247 (N_5247,N_4953,N_4503);
and U5248 (N_5248,N_4957,N_4238);
or U5249 (N_5249,N_4473,N_4827);
and U5250 (N_5250,N_4033,N_4812);
nand U5251 (N_5251,N_4218,N_4192);
xor U5252 (N_5252,N_4650,N_4518);
nand U5253 (N_5253,N_4461,N_4787);
nand U5254 (N_5254,N_4549,N_4209);
and U5255 (N_5255,N_4088,N_4464);
or U5256 (N_5256,N_4982,N_4665);
nand U5257 (N_5257,N_4073,N_4996);
or U5258 (N_5258,N_4686,N_4794);
nor U5259 (N_5259,N_4542,N_4969);
and U5260 (N_5260,N_4863,N_4977);
or U5261 (N_5261,N_4799,N_4829);
nand U5262 (N_5262,N_4991,N_4867);
xnor U5263 (N_5263,N_4176,N_4899);
nand U5264 (N_5264,N_4239,N_4619);
nand U5265 (N_5265,N_4561,N_4480);
and U5266 (N_5266,N_4351,N_4041);
xor U5267 (N_5267,N_4634,N_4533);
xnor U5268 (N_5268,N_4830,N_4353);
or U5269 (N_5269,N_4496,N_4452);
and U5270 (N_5270,N_4378,N_4081);
nor U5271 (N_5271,N_4185,N_4342);
xor U5272 (N_5272,N_4591,N_4612);
nand U5273 (N_5273,N_4779,N_4837);
nor U5274 (N_5274,N_4281,N_4564);
nand U5275 (N_5275,N_4885,N_4279);
nand U5276 (N_5276,N_4438,N_4531);
xnor U5277 (N_5277,N_4497,N_4757);
and U5278 (N_5278,N_4487,N_4796);
nor U5279 (N_5279,N_4037,N_4479);
nand U5280 (N_5280,N_4849,N_4708);
or U5281 (N_5281,N_4765,N_4417);
xnor U5282 (N_5282,N_4384,N_4141);
and U5283 (N_5283,N_4884,N_4040);
nor U5284 (N_5284,N_4502,N_4132);
or U5285 (N_5285,N_4964,N_4465);
xor U5286 (N_5286,N_4006,N_4300);
and U5287 (N_5287,N_4696,N_4826);
and U5288 (N_5288,N_4644,N_4900);
xnor U5289 (N_5289,N_4498,N_4285);
and U5290 (N_5290,N_4963,N_4115);
nand U5291 (N_5291,N_4336,N_4408);
or U5292 (N_5292,N_4017,N_4337);
nand U5293 (N_5293,N_4026,N_4173);
nor U5294 (N_5294,N_4457,N_4393);
or U5295 (N_5295,N_4878,N_4688);
or U5296 (N_5296,N_4851,N_4023);
nor U5297 (N_5297,N_4506,N_4102);
xnor U5298 (N_5298,N_4770,N_4711);
and U5299 (N_5299,N_4087,N_4236);
and U5300 (N_5300,N_4907,N_4468);
nand U5301 (N_5301,N_4194,N_4673);
nand U5302 (N_5302,N_4880,N_4396);
xor U5303 (N_5303,N_4816,N_4454);
and U5304 (N_5304,N_4310,N_4405);
nor U5305 (N_5305,N_4369,N_4875);
xnor U5306 (N_5306,N_4009,N_4984);
and U5307 (N_5307,N_4545,N_4109);
nand U5308 (N_5308,N_4138,N_4232);
or U5309 (N_5309,N_4572,N_4527);
and U5310 (N_5310,N_4152,N_4402);
xor U5311 (N_5311,N_4872,N_4302);
or U5312 (N_5312,N_4451,N_4252);
and U5313 (N_5313,N_4357,N_4044);
xor U5314 (N_5314,N_4015,N_4107);
and U5315 (N_5315,N_4134,N_4762);
xor U5316 (N_5316,N_4078,N_4753);
nor U5317 (N_5317,N_4970,N_4453);
or U5318 (N_5318,N_4387,N_4262);
xor U5319 (N_5319,N_4303,N_4813);
or U5320 (N_5320,N_4161,N_4448);
xor U5321 (N_5321,N_4597,N_4246);
and U5322 (N_5322,N_4409,N_4840);
xnor U5323 (N_5323,N_4555,N_4682);
or U5324 (N_5324,N_4587,N_4223);
xor U5325 (N_5325,N_4399,N_4788);
nor U5326 (N_5326,N_4291,N_4156);
xnor U5327 (N_5327,N_4501,N_4019);
nor U5328 (N_5328,N_4318,N_4764);
xor U5329 (N_5329,N_4763,N_4235);
xnor U5330 (N_5330,N_4251,N_4698);
xnor U5331 (N_5331,N_4265,N_4407);
and U5332 (N_5332,N_4057,N_4802);
or U5333 (N_5333,N_4344,N_4574);
nand U5334 (N_5334,N_4905,N_4922);
nand U5335 (N_5335,N_4671,N_4428);
nor U5336 (N_5336,N_4021,N_4978);
xor U5337 (N_5337,N_4311,N_4488);
xor U5338 (N_5338,N_4994,N_4288);
nor U5339 (N_5339,N_4145,N_4420);
or U5340 (N_5340,N_4183,N_4523);
xor U5341 (N_5341,N_4334,N_4948);
nand U5342 (N_5342,N_4117,N_4734);
nand U5343 (N_5343,N_4810,N_4656);
nor U5344 (N_5344,N_4083,N_4592);
nor U5345 (N_5345,N_4979,N_4367);
or U5346 (N_5346,N_4314,N_4825);
xnor U5347 (N_5347,N_4722,N_4007);
nor U5348 (N_5348,N_4912,N_4573);
xor U5349 (N_5349,N_4169,N_4932);
xor U5350 (N_5350,N_4386,N_4955);
and U5351 (N_5351,N_4047,N_4153);
nor U5352 (N_5352,N_4298,N_4993);
and U5353 (N_5353,N_4940,N_4358);
nand U5354 (N_5354,N_4062,N_4147);
nand U5355 (N_5355,N_4716,N_4027);
xnor U5356 (N_5356,N_4934,N_4306);
and U5357 (N_5357,N_4149,N_4528);
xor U5358 (N_5358,N_4714,N_4242);
and U5359 (N_5359,N_4705,N_4589);
and U5360 (N_5360,N_4560,N_4653);
and U5361 (N_5361,N_4328,N_4292);
nor U5362 (N_5362,N_4284,N_4559);
nor U5363 (N_5363,N_4522,N_4397);
or U5364 (N_5364,N_4622,N_4718);
nand U5365 (N_5365,N_4602,N_4035);
nand U5366 (N_5366,N_4856,N_4267);
or U5367 (N_5367,N_4315,N_4486);
nor U5368 (N_5368,N_4700,N_4985);
or U5369 (N_5369,N_4139,N_4917);
nand U5370 (N_5370,N_4483,N_4585);
and U5371 (N_5371,N_4150,N_4713);
nand U5372 (N_5372,N_4607,N_4203);
nor U5373 (N_5373,N_4942,N_4593);
xor U5374 (N_5374,N_4418,N_4808);
nor U5375 (N_5375,N_4750,N_4493);
nor U5376 (N_5376,N_4360,N_4340);
and U5377 (N_5377,N_4130,N_4365);
xnor U5378 (N_5378,N_4160,N_4294);
nor U5379 (N_5379,N_4609,N_4212);
nand U5380 (N_5380,N_4834,N_4823);
and U5381 (N_5381,N_4423,N_4562);
xnor U5382 (N_5382,N_4630,N_4075);
or U5383 (N_5383,N_4645,N_4022);
nand U5384 (N_5384,N_4072,N_4067);
nand U5385 (N_5385,N_4256,N_4886);
and U5386 (N_5386,N_4514,N_4191);
and U5387 (N_5387,N_4000,N_4895);
nand U5388 (N_5388,N_4929,N_4882);
xor U5389 (N_5389,N_4553,N_4697);
or U5390 (N_5390,N_4539,N_4667);
xor U5391 (N_5391,N_4780,N_4307);
and U5392 (N_5392,N_4554,N_4277);
or U5393 (N_5393,N_4563,N_4100);
or U5394 (N_5394,N_4818,N_4355);
and U5395 (N_5395,N_4657,N_4472);
xnor U5396 (N_5396,N_4446,N_4509);
nand U5397 (N_5397,N_4704,N_4489);
or U5398 (N_5398,N_4952,N_4164);
xor U5399 (N_5399,N_4793,N_4521);
nor U5400 (N_5400,N_4443,N_4773);
xor U5401 (N_5401,N_4989,N_4020);
xnor U5402 (N_5402,N_4639,N_4039);
xnor U5403 (N_5403,N_4975,N_4228);
nor U5404 (N_5404,N_4577,N_4361);
and U5405 (N_5405,N_4206,N_4283);
nor U5406 (N_5406,N_4199,N_4606);
nor U5407 (N_5407,N_4261,N_4025);
nand U5408 (N_5408,N_4247,N_4249);
or U5409 (N_5409,N_4741,N_4781);
nor U5410 (N_5410,N_4848,N_4869);
nand U5411 (N_5411,N_4190,N_4749);
nor U5412 (N_5412,N_4401,N_4981);
or U5413 (N_5413,N_4596,N_4508);
nand U5414 (N_5414,N_4887,N_4608);
and U5415 (N_5415,N_4376,N_4838);
xnor U5416 (N_5416,N_4219,N_4116);
nand U5417 (N_5417,N_4477,N_4581);
xor U5418 (N_5418,N_4211,N_4729);
nor U5419 (N_5419,N_4170,N_4349);
and U5420 (N_5420,N_4202,N_4427);
nand U5421 (N_5421,N_4719,N_4158);
or U5422 (N_5422,N_4902,N_4641);
and U5423 (N_5423,N_4586,N_4059);
and U5424 (N_5424,N_4335,N_4512);
nor U5425 (N_5425,N_4188,N_4726);
nand U5426 (N_5426,N_4113,N_4410);
nor U5427 (N_5427,N_4165,N_4326);
xor U5428 (N_5428,N_4492,N_4854);
and U5429 (N_5429,N_4106,N_4201);
nand U5430 (N_5430,N_4255,N_4034);
or U5431 (N_5431,N_4954,N_4484);
xor U5432 (N_5432,N_4868,N_4894);
nand U5433 (N_5433,N_4374,N_4507);
xnor U5434 (N_5434,N_4786,N_4980);
and U5435 (N_5435,N_4500,N_4515);
and U5436 (N_5436,N_4388,N_4636);
or U5437 (N_5437,N_4646,N_4558);
nand U5438 (N_5438,N_4304,N_4611);
nor U5439 (N_5439,N_4651,N_4060);
nor U5440 (N_5440,N_4168,N_4198);
and U5441 (N_5441,N_4640,N_4958);
nor U5442 (N_5442,N_4723,N_4960);
or U5443 (N_5443,N_4551,N_4148);
or U5444 (N_5444,N_4844,N_4031);
and U5445 (N_5445,N_4906,N_4511);
nor U5446 (N_5446,N_4604,N_4200);
nor U5447 (N_5447,N_4482,N_4167);
nand U5448 (N_5448,N_4935,N_4997);
or U5449 (N_5449,N_4316,N_4433);
nand U5450 (N_5450,N_4774,N_4866);
xnor U5451 (N_5451,N_4475,N_4803);
nor U5452 (N_5452,N_4128,N_4758);
and U5453 (N_5453,N_4324,N_4972);
nor U5454 (N_5454,N_4809,N_4227);
nand U5455 (N_5455,N_4415,N_4821);
or U5456 (N_5456,N_4184,N_4122);
nand U5457 (N_5457,N_4783,N_4372);
nand U5458 (N_5458,N_4831,N_4322);
xnor U5459 (N_5459,N_4352,N_4392);
and U5460 (N_5460,N_4594,N_4177);
or U5461 (N_5461,N_4424,N_4379);
and U5462 (N_5462,N_4179,N_4926);
nor U5463 (N_5463,N_4847,N_4901);
nand U5464 (N_5464,N_4751,N_4766);
or U5465 (N_5465,N_4680,N_4768);
or U5466 (N_5466,N_4491,N_4469);
nor U5467 (N_5467,N_4226,N_4440);
xor U5468 (N_5468,N_4245,N_4350);
nor U5469 (N_5469,N_4187,N_4801);
or U5470 (N_5470,N_4546,N_4918);
nand U5471 (N_5471,N_4066,N_4702);
or U5472 (N_5472,N_4828,N_4045);
nand U5473 (N_5473,N_4913,N_4076);
nand U5474 (N_5474,N_4832,N_4253);
nor U5475 (N_5475,N_4260,N_4898);
and U5476 (N_5476,N_4931,N_4857);
or U5477 (N_5477,N_4494,N_4126);
nand U5478 (N_5478,N_4259,N_4624);
and U5479 (N_5479,N_4096,N_4524);
xnor U5480 (N_5480,N_4709,N_4583);
nor U5481 (N_5481,N_4566,N_4800);
nand U5482 (N_5482,N_4481,N_4933);
xor U5483 (N_5483,N_4442,N_4412);
and U5484 (N_5484,N_4791,N_4655);
and U5485 (N_5485,N_4330,N_4874);
nor U5486 (N_5486,N_4988,N_4998);
xor U5487 (N_5487,N_4331,N_4368);
xnor U5488 (N_5488,N_4668,N_4426);
or U5489 (N_5489,N_4366,N_4248);
xor U5490 (N_5490,N_4058,N_4257);
and U5491 (N_5491,N_4222,N_4631);
and U5492 (N_5492,N_4069,N_4914);
nor U5493 (N_5493,N_4054,N_4056);
or U5494 (N_5494,N_4400,N_4771);
or U5495 (N_5495,N_4625,N_4712);
and U5496 (N_5496,N_4663,N_4510);
nor U5497 (N_5497,N_4864,N_4548);
or U5498 (N_5498,N_4390,N_4568);
xnor U5499 (N_5499,N_4356,N_4571);
nand U5500 (N_5500,N_4431,N_4823);
xnor U5501 (N_5501,N_4449,N_4207);
nor U5502 (N_5502,N_4163,N_4359);
xnor U5503 (N_5503,N_4518,N_4728);
nor U5504 (N_5504,N_4477,N_4583);
nor U5505 (N_5505,N_4320,N_4551);
xor U5506 (N_5506,N_4769,N_4459);
xor U5507 (N_5507,N_4690,N_4798);
nor U5508 (N_5508,N_4866,N_4277);
xor U5509 (N_5509,N_4613,N_4535);
and U5510 (N_5510,N_4185,N_4242);
and U5511 (N_5511,N_4164,N_4379);
and U5512 (N_5512,N_4777,N_4683);
nand U5513 (N_5513,N_4113,N_4427);
and U5514 (N_5514,N_4202,N_4982);
nor U5515 (N_5515,N_4975,N_4106);
nor U5516 (N_5516,N_4929,N_4814);
and U5517 (N_5517,N_4062,N_4823);
nand U5518 (N_5518,N_4080,N_4540);
or U5519 (N_5519,N_4708,N_4035);
xnor U5520 (N_5520,N_4172,N_4289);
and U5521 (N_5521,N_4436,N_4559);
nand U5522 (N_5522,N_4790,N_4917);
or U5523 (N_5523,N_4887,N_4091);
or U5524 (N_5524,N_4091,N_4702);
xor U5525 (N_5525,N_4666,N_4645);
xnor U5526 (N_5526,N_4930,N_4454);
and U5527 (N_5527,N_4455,N_4432);
xor U5528 (N_5528,N_4785,N_4225);
xnor U5529 (N_5529,N_4495,N_4259);
nor U5530 (N_5530,N_4425,N_4734);
xor U5531 (N_5531,N_4829,N_4397);
nor U5532 (N_5532,N_4833,N_4560);
and U5533 (N_5533,N_4653,N_4455);
or U5534 (N_5534,N_4037,N_4432);
xnor U5535 (N_5535,N_4272,N_4140);
xnor U5536 (N_5536,N_4351,N_4837);
nor U5537 (N_5537,N_4796,N_4414);
nand U5538 (N_5538,N_4450,N_4881);
and U5539 (N_5539,N_4355,N_4500);
nand U5540 (N_5540,N_4070,N_4043);
and U5541 (N_5541,N_4858,N_4265);
xnor U5542 (N_5542,N_4158,N_4649);
nor U5543 (N_5543,N_4183,N_4092);
nand U5544 (N_5544,N_4305,N_4919);
nor U5545 (N_5545,N_4310,N_4865);
xnor U5546 (N_5546,N_4014,N_4011);
nand U5547 (N_5547,N_4126,N_4559);
nand U5548 (N_5548,N_4335,N_4608);
and U5549 (N_5549,N_4607,N_4460);
xnor U5550 (N_5550,N_4093,N_4679);
or U5551 (N_5551,N_4167,N_4847);
nand U5552 (N_5552,N_4802,N_4325);
or U5553 (N_5553,N_4157,N_4727);
nor U5554 (N_5554,N_4376,N_4454);
xor U5555 (N_5555,N_4438,N_4780);
and U5556 (N_5556,N_4586,N_4842);
and U5557 (N_5557,N_4609,N_4411);
nor U5558 (N_5558,N_4955,N_4233);
xnor U5559 (N_5559,N_4382,N_4754);
and U5560 (N_5560,N_4291,N_4985);
and U5561 (N_5561,N_4053,N_4701);
or U5562 (N_5562,N_4966,N_4314);
xor U5563 (N_5563,N_4675,N_4521);
nand U5564 (N_5564,N_4510,N_4943);
or U5565 (N_5565,N_4752,N_4448);
xnor U5566 (N_5566,N_4116,N_4609);
or U5567 (N_5567,N_4087,N_4364);
and U5568 (N_5568,N_4642,N_4193);
xor U5569 (N_5569,N_4476,N_4475);
nand U5570 (N_5570,N_4545,N_4638);
and U5571 (N_5571,N_4940,N_4095);
or U5572 (N_5572,N_4516,N_4217);
and U5573 (N_5573,N_4239,N_4833);
xnor U5574 (N_5574,N_4165,N_4270);
nor U5575 (N_5575,N_4890,N_4285);
xnor U5576 (N_5576,N_4162,N_4453);
nand U5577 (N_5577,N_4447,N_4353);
nand U5578 (N_5578,N_4182,N_4113);
nand U5579 (N_5579,N_4852,N_4024);
xnor U5580 (N_5580,N_4030,N_4742);
xor U5581 (N_5581,N_4154,N_4446);
nand U5582 (N_5582,N_4624,N_4547);
or U5583 (N_5583,N_4546,N_4193);
xnor U5584 (N_5584,N_4243,N_4454);
nor U5585 (N_5585,N_4810,N_4056);
nand U5586 (N_5586,N_4351,N_4076);
and U5587 (N_5587,N_4087,N_4814);
nand U5588 (N_5588,N_4065,N_4943);
and U5589 (N_5589,N_4534,N_4809);
and U5590 (N_5590,N_4062,N_4888);
xor U5591 (N_5591,N_4811,N_4506);
and U5592 (N_5592,N_4891,N_4394);
nor U5593 (N_5593,N_4882,N_4569);
xnor U5594 (N_5594,N_4877,N_4848);
or U5595 (N_5595,N_4758,N_4382);
nand U5596 (N_5596,N_4048,N_4894);
and U5597 (N_5597,N_4583,N_4860);
nor U5598 (N_5598,N_4507,N_4958);
and U5599 (N_5599,N_4179,N_4965);
xnor U5600 (N_5600,N_4417,N_4782);
and U5601 (N_5601,N_4221,N_4504);
xnor U5602 (N_5602,N_4742,N_4515);
xnor U5603 (N_5603,N_4416,N_4584);
xor U5604 (N_5604,N_4265,N_4563);
xnor U5605 (N_5605,N_4224,N_4310);
nor U5606 (N_5606,N_4584,N_4293);
nand U5607 (N_5607,N_4739,N_4759);
nor U5608 (N_5608,N_4259,N_4876);
nor U5609 (N_5609,N_4763,N_4409);
or U5610 (N_5610,N_4837,N_4065);
xnor U5611 (N_5611,N_4339,N_4583);
or U5612 (N_5612,N_4389,N_4960);
nor U5613 (N_5613,N_4895,N_4172);
nor U5614 (N_5614,N_4021,N_4504);
xnor U5615 (N_5615,N_4686,N_4846);
and U5616 (N_5616,N_4020,N_4081);
xnor U5617 (N_5617,N_4913,N_4685);
nand U5618 (N_5618,N_4074,N_4970);
and U5619 (N_5619,N_4987,N_4771);
or U5620 (N_5620,N_4922,N_4548);
nor U5621 (N_5621,N_4430,N_4619);
and U5622 (N_5622,N_4138,N_4294);
nor U5623 (N_5623,N_4065,N_4613);
or U5624 (N_5624,N_4788,N_4896);
nor U5625 (N_5625,N_4267,N_4081);
xnor U5626 (N_5626,N_4171,N_4367);
or U5627 (N_5627,N_4078,N_4711);
nand U5628 (N_5628,N_4578,N_4976);
or U5629 (N_5629,N_4495,N_4149);
or U5630 (N_5630,N_4762,N_4426);
nand U5631 (N_5631,N_4368,N_4431);
nand U5632 (N_5632,N_4182,N_4557);
or U5633 (N_5633,N_4497,N_4026);
or U5634 (N_5634,N_4152,N_4679);
nand U5635 (N_5635,N_4035,N_4677);
xnor U5636 (N_5636,N_4870,N_4945);
xor U5637 (N_5637,N_4860,N_4413);
or U5638 (N_5638,N_4466,N_4388);
nand U5639 (N_5639,N_4439,N_4497);
xor U5640 (N_5640,N_4676,N_4927);
xnor U5641 (N_5641,N_4777,N_4796);
and U5642 (N_5642,N_4976,N_4381);
or U5643 (N_5643,N_4727,N_4349);
and U5644 (N_5644,N_4907,N_4684);
and U5645 (N_5645,N_4550,N_4773);
and U5646 (N_5646,N_4418,N_4995);
or U5647 (N_5647,N_4746,N_4643);
xnor U5648 (N_5648,N_4161,N_4128);
nor U5649 (N_5649,N_4671,N_4076);
and U5650 (N_5650,N_4899,N_4089);
xnor U5651 (N_5651,N_4676,N_4353);
nand U5652 (N_5652,N_4805,N_4923);
and U5653 (N_5653,N_4569,N_4601);
nand U5654 (N_5654,N_4618,N_4583);
nand U5655 (N_5655,N_4015,N_4636);
nand U5656 (N_5656,N_4362,N_4467);
xnor U5657 (N_5657,N_4878,N_4015);
nor U5658 (N_5658,N_4171,N_4638);
nor U5659 (N_5659,N_4310,N_4443);
xor U5660 (N_5660,N_4770,N_4372);
nor U5661 (N_5661,N_4003,N_4511);
nand U5662 (N_5662,N_4835,N_4453);
nand U5663 (N_5663,N_4323,N_4312);
nor U5664 (N_5664,N_4681,N_4420);
xor U5665 (N_5665,N_4143,N_4215);
xor U5666 (N_5666,N_4655,N_4110);
nand U5667 (N_5667,N_4046,N_4794);
and U5668 (N_5668,N_4766,N_4057);
and U5669 (N_5669,N_4477,N_4711);
xnor U5670 (N_5670,N_4824,N_4569);
or U5671 (N_5671,N_4513,N_4441);
xnor U5672 (N_5672,N_4636,N_4764);
or U5673 (N_5673,N_4959,N_4893);
nand U5674 (N_5674,N_4617,N_4281);
or U5675 (N_5675,N_4991,N_4973);
or U5676 (N_5676,N_4962,N_4568);
xor U5677 (N_5677,N_4036,N_4564);
nand U5678 (N_5678,N_4786,N_4723);
or U5679 (N_5679,N_4719,N_4659);
nor U5680 (N_5680,N_4676,N_4838);
xor U5681 (N_5681,N_4269,N_4137);
nand U5682 (N_5682,N_4647,N_4351);
nor U5683 (N_5683,N_4375,N_4032);
nand U5684 (N_5684,N_4505,N_4546);
or U5685 (N_5685,N_4726,N_4812);
nand U5686 (N_5686,N_4127,N_4287);
and U5687 (N_5687,N_4244,N_4169);
nor U5688 (N_5688,N_4425,N_4108);
nand U5689 (N_5689,N_4649,N_4464);
nor U5690 (N_5690,N_4742,N_4540);
nor U5691 (N_5691,N_4754,N_4879);
nor U5692 (N_5692,N_4144,N_4278);
nand U5693 (N_5693,N_4941,N_4000);
xnor U5694 (N_5694,N_4561,N_4047);
nor U5695 (N_5695,N_4262,N_4253);
or U5696 (N_5696,N_4153,N_4932);
nand U5697 (N_5697,N_4447,N_4045);
nor U5698 (N_5698,N_4452,N_4212);
nand U5699 (N_5699,N_4006,N_4001);
nor U5700 (N_5700,N_4366,N_4785);
xor U5701 (N_5701,N_4331,N_4638);
nor U5702 (N_5702,N_4788,N_4513);
and U5703 (N_5703,N_4063,N_4279);
nor U5704 (N_5704,N_4138,N_4677);
xor U5705 (N_5705,N_4496,N_4248);
nor U5706 (N_5706,N_4034,N_4889);
or U5707 (N_5707,N_4246,N_4154);
nor U5708 (N_5708,N_4535,N_4824);
or U5709 (N_5709,N_4901,N_4414);
nand U5710 (N_5710,N_4412,N_4032);
or U5711 (N_5711,N_4436,N_4654);
and U5712 (N_5712,N_4432,N_4028);
and U5713 (N_5713,N_4848,N_4124);
nand U5714 (N_5714,N_4837,N_4815);
xor U5715 (N_5715,N_4813,N_4869);
nor U5716 (N_5716,N_4836,N_4161);
nand U5717 (N_5717,N_4936,N_4305);
nor U5718 (N_5718,N_4201,N_4587);
and U5719 (N_5719,N_4045,N_4889);
xnor U5720 (N_5720,N_4639,N_4795);
or U5721 (N_5721,N_4275,N_4157);
nor U5722 (N_5722,N_4029,N_4509);
and U5723 (N_5723,N_4193,N_4621);
or U5724 (N_5724,N_4321,N_4571);
nor U5725 (N_5725,N_4500,N_4378);
xor U5726 (N_5726,N_4811,N_4371);
and U5727 (N_5727,N_4281,N_4638);
nand U5728 (N_5728,N_4105,N_4707);
and U5729 (N_5729,N_4674,N_4075);
and U5730 (N_5730,N_4535,N_4812);
or U5731 (N_5731,N_4268,N_4351);
and U5732 (N_5732,N_4105,N_4300);
nor U5733 (N_5733,N_4173,N_4284);
xnor U5734 (N_5734,N_4134,N_4732);
nor U5735 (N_5735,N_4754,N_4266);
nand U5736 (N_5736,N_4753,N_4009);
xnor U5737 (N_5737,N_4907,N_4973);
xnor U5738 (N_5738,N_4047,N_4928);
and U5739 (N_5739,N_4307,N_4231);
and U5740 (N_5740,N_4102,N_4188);
and U5741 (N_5741,N_4934,N_4883);
and U5742 (N_5742,N_4981,N_4446);
xnor U5743 (N_5743,N_4741,N_4709);
nand U5744 (N_5744,N_4419,N_4256);
or U5745 (N_5745,N_4520,N_4273);
and U5746 (N_5746,N_4545,N_4451);
and U5747 (N_5747,N_4736,N_4238);
nor U5748 (N_5748,N_4632,N_4068);
xnor U5749 (N_5749,N_4354,N_4274);
nand U5750 (N_5750,N_4528,N_4619);
xnor U5751 (N_5751,N_4118,N_4820);
nand U5752 (N_5752,N_4293,N_4990);
nor U5753 (N_5753,N_4081,N_4769);
xor U5754 (N_5754,N_4500,N_4860);
nand U5755 (N_5755,N_4159,N_4520);
or U5756 (N_5756,N_4165,N_4825);
xnor U5757 (N_5757,N_4163,N_4691);
xor U5758 (N_5758,N_4568,N_4369);
nand U5759 (N_5759,N_4993,N_4574);
nand U5760 (N_5760,N_4910,N_4533);
xor U5761 (N_5761,N_4622,N_4723);
xor U5762 (N_5762,N_4101,N_4889);
and U5763 (N_5763,N_4767,N_4372);
nor U5764 (N_5764,N_4459,N_4337);
or U5765 (N_5765,N_4876,N_4184);
or U5766 (N_5766,N_4806,N_4647);
and U5767 (N_5767,N_4259,N_4957);
xnor U5768 (N_5768,N_4709,N_4976);
xnor U5769 (N_5769,N_4076,N_4532);
and U5770 (N_5770,N_4344,N_4800);
and U5771 (N_5771,N_4419,N_4917);
nand U5772 (N_5772,N_4802,N_4439);
and U5773 (N_5773,N_4811,N_4105);
or U5774 (N_5774,N_4707,N_4602);
and U5775 (N_5775,N_4177,N_4698);
or U5776 (N_5776,N_4828,N_4795);
or U5777 (N_5777,N_4520,N_4436);
xor U5778 (N_5778,N_4560,N_4251);
or U5779 (N_5779,N_4838,N_4792);
and U5780 (N_5780,N_4663,N_4299);
and U5781 (N_5781,N_4733,N_4149);
xor U5782 (N_5782,N_4178,N_4538);
or U5783 (N_5783,N_4913,N_4340);
nor U5784 (N_5784,N_4487,N_4124);
or U5785 (N_5785,N_4930,N_4318);
nor U5786 (N_5786,N_4428,N_4719);
nand U5787 (N_5787,N_4157,N_4647);
xor U5788 (N_5788,N_4235,N_4913);
and U5789 (N_5789,N_4810,N_4599);
nor U5790 (N_5790,N_4507,N_4782);
nor U5791 (N_5791,N_4403,N_4366);
xnor U5792 (N_5792,N_4114,N_4921);
and U5793 (N_5793,N_4756,N_4599);
or U5794 (N_5794,N_4627,N_4212);
and U5795 (N_5795,N_4346,N_4391);
xnor U5796 (N_5796,N_4806,N_4603);
xor U5797 (N_5797,N_4948,N_4452);
or U5798 (N_5798,N_4209,N_4521);
and U5799 (N_5799,N_4155,N_4727);
xor U5800 (N_5800,N_4287,N_4932);
and U5801 (N_5801,N_4172,N_4123);
xor U5802 (N_5802,N_4352,N_4452);
nor U5803 (N_5803,N_4744,N_4672);
nor U5804 (N_5804,N_4279,N_4445);
xor U5805 (N_5805,N_4374,N_4948);
or U5806 (N_5806,N_4668,N_4814);
nor U5807 (N_5807,N_4350,N_4365);
and U5808 (N_5808,N_4013,N_4717);
or U5809 (N_5809,N_4329,N_4940);
xor U5810 (N_5810,N_4004,N_4889);
nor U5811 (N_5811,N_4045,N_4739);
nor U5812 (N_5812,N_4362,N_4840);
and U5813 (N_5813,N_4386,N_4656);
nor U5814 (N_5814,N_4498,N_4361);
nand U5815 (N_5815,N_4993,N_4324);
xor U5816 (N_5816,N_4451,N_4298);
and U5817 (N_5817,N_4330,N_4327);
or U5818 (N_5818,N_4009,N_4809);
xnor U5819 (N_5819,N_4448,N_4397);
nand U5820 (N_5820,N_4376,N_4340);
and U5821 (N_5821,N_4712,N_4010);
xor U5822 (N_5822,N_4966,N_4755);
or U5823 (N_5823,N_4641,N_4375);
nor U5824 (N_5824,N_4992,N_4539);
or U5825 (N_5825,N_4971,N_4185);
or U5826 (N_5826,N_4895,N_4412);
nand U5827 (N_5827,N_4880,N_4099);
nand U5828 (N_5828,N_4297,N_4012);
xnor U5829 (N_5829,N_4940,N_4727);
xor U5830 (N_5830,N_4090,N_4962);
nor U5831 (N_5831,N_4113,N_4965);
xnor U5832 (N_5832,N_4756,N_4937);
or U5833 (N_5833,N_4456,N_4366);
xnor U5834 (N_5834,N_4317,N_4277);
xnor U5835 (N_5835,N_4685,N_4935);
or U5836 (N_5836,N_4692,N_4802);
and U5837 (N_5837,N_4235,N_4587);
xnor U5838 (N_5838,N_4653,N_4113);
nor U5839 (N_5839,N_4281,N_4672);
xnor U5840 (N_5840,N_4121,N_4246);
or U5841 (N_5841,N_4328,N_4295);
and U5842 (N_5842,N_4894,N_4816);
nor U5843 (N_5843,N_4919,N_4893);
and U5844 (N_5844,N_4510,N_4200);
xor U5845 (N_5845,N_4176,N_4643);
nand U5846 (N_5846,N_4338,N_4865);
nand U5847 (N_5847,N_4614,N_4877);
nand U5848 (N_5848,N_4527,N_4178);
and U5849 (N_5849,N_4603,N_4908);
and U5850 (N_5850,N_4671,N_4004);
nor U5851 (N_5851,N_4358,N_4910);
or U5852 (N_5852,N_4344,N_4696);
and U5853 (N_5853,N_4641,N_4766);
and U5854 (N_5854,N_4757,N_4204);
nand U5855 (N_5855,N_4037,N_4056);
xnor U5856 (N_5856,N_4625,N_4422);
or U5857 (N_5857,N_4368,N_4522);
nor U5858 (N_5858,N_4878,N_4157);
or U5859 (N_5859,N_4245,N_4685);
xnor U5860 (N_5860,N_4352,N_4687);
xor U5861 (N_5861,N_4003,N_4556);
nand U5862 (N_5862,N_4146,N_4797);
nor U5863 (N_5863,N_4494,N_4652);
and U5864 (N_5864,N_4111,N_4306);
and U5865 (N_5865,N_4246,N_4883);
and U5866 (N_5866,N_4344,N_4029);
nand U5867 (N_5867,N_4811,N_4828);
or U5868 (N_5868,N_4152,N_4928);
xnor U5869 (N_5869,N_4009,N_4101);
and U5870 (N_5870,N_4780,N_4422);
nand U5871 (N_5871,N_4311,N_4901);
nor U5872 (N_5872,N_4541,N_4413);
nor U5873 (N_5873,N_4657,N_4898);
and U5874 (N_5874,N_4512,N_4898);
nand U5875 (N_5875,N_4677,N_4618);
xnor U5876 (N_5876,N_4806,N_4615);
nand U5877 (N_5877,N_4768,N_4782);
or U5878 (N_5878,N_4050,N_4417);
xor U5879 (N_5879,N_4338,N_4955);
nor U5880 (N_5880,N_4178,N_4266);
nor U5881 (N_5881,N_4683,N_4898);
or U5882 (N_5882,N_4651,N_4423);
or U5883 (N_5883,N_4015,N_4831);
xnor U5884 (N_5884,N_4756,N_4701);
nand U5885 (N_5885,N_4110,N_4896);
and U5886 (N_5886,N_4256,N_4199);
nor U5887 (N_5887,N_4859,N_4965);
nand U5888 (N_5888,N_4724,N_4769);
or U5889 (N_5889,N_4374,N_4322);
xnor U5890 (N_5890,N_4191,N_4628);
nand U5891 (N_5891,N_4966,N_4281);
xor U5892 (N_5892,N_4666,N_4461);
nor U5893 (N_5893,N_4701,N_4723);
nand U5894 (N_5894,N_4999,N_4080);
xnor U5895 (N_5895,N_4519,N_4520);
xnor U5896 (N_5896,N_4116,N_4156);
nor U5897 (N_5897,N_4423,N_4468);
nor U5898 (N_5898,N_4752,N_4065);
and U5899 (N_5899,N_4248,N_4196);
nor U5900 (N_5900,N_4778,N_4008);
and U5901 (N_5901,N_4537,N_4375);
xnor U5902 (N_5902,N_4649,N_4647);
nor U5903 (N_5903,N_4943,N_4141);
nor U5904 (N_5904,N_4730,N_4645);
nand U5905 (N_5905,N_4630,N_4750);
nand U5906 (N_5906,N_4574,N_4486);
nor U5907 (N_5907,N_4346,N_4980);
and U5908 (N_5908,N_4344,N_4000);
nand U5909 (N_5909,N_4397,N_4066);
or U5910 (N_5910,N_4839,N_4516);
or U5911 (N_5911,N_4814,N_4256);
xor U5912 (N_5912,N_4958,N_4067);
and U5913 (N_5913,N_4875,N_4810);
xor U5914 (N_5914,N_4218,N_4891);
xnor U5915 (N_5915,N_4220,N_4797);
and U5916 (N_5916,N_4688,N_4208);
nand U5917 (N_5917,N_4696,N_4753);
nor U5918 (N_5918,N_4133,N_4636);
nor U5919 (N_5919,N_4021,N_4589);
nor U5920 (N_5920,N_4844,N_4505);
nor U5921 (N_5921,N_4222,N_4231);
nor U5922 (N_5922,N_4389,N_4647);
and U5923 (N_5923,N_4734,N_4849);
or U5924 (N_5924,N_4752,N_4432);
nor U5925 (N_5925,N_4379,N_4508);
nor U5926 (N_5926,N_4349,N_4419);
or U5927 (N_5927,N_4087,N_4529);
xnor U5928 (N_5928,N_4958,N_4243);
or U5929 (N_5929,N_4603,N_4563);
xnor U5930 (N_5930,N_4210,N_4960);
or U5931 (N_5931,N_4608,N_4258);
nor U5932 (N_5932,N_4946,N_4766);
nand U5933 (N_5933,N_4450,N_4780);
nor U5934 (N_5934,N_4666,N_4247);
and U5935 (N_5935,N_4948,N_4865);
nor U5936 (N_5936,N_4230,N_4306);
or U5937 (N_5937,N_4216,N_4272);
nor U5938 (N_5938,N_4351,N_4656);
nand U5939 (N_5939,N_4730,N_4104);
xor U5940 (N_5940,N_4730,N_4046);
nor U5941 (N_5941,N_4590,N_4692);
nand U5942 (N_5942,N_4339,N_4837);
and U5943 (N_5943,N_4656,N_4436);
nand U5944 (N_5944,N_4664,N_4456);
or U5945 (N_5945,N_4774,N_4133);
nand U5946 (N_5946,N_4897,N_4220);
nor U5947 (N_5947,N_4891,N_4326);
nor U5948 (N_5948,N_4073,N_4027);
xnor U5949 (N_5949,N_4239,N_4253);
nand U5950 (N_5950,N_4099,N_4590);
nand U5951 (N_5951,N_4416,N_4404);
and U5952 (N_5952,N_4382,N_4341);
nand U5953 (N_5953,N_4645,N_4129);
xor U5954 (N_5954,N_4500,N_4398);
xor U5955 (N_5955,N_4193,N_4842);
nor U5956 (N_5956,N_4187,N_4083);
nand U5957 (N_5957,N_4400,N_4615);
nand U5958 (N_5958,N_4534,N_4169);
and U5959 (N_5959,N_4174,N_4802);
nand U5960 (N_5960,N_4916,N_4738);
nand U5961 (N_5961,N_4918,N_4687);
xnor U5962 (N_5962,N_4882,N_4923);
xor U5963 (N_5963,N_4176,N_4256);
xor U5964 (N_5964,N_4104,N_4822);
and U5965 (N_5965,N_4387,N_4477);
xor U5966 (N_5966,N_4644,N_4694);
nor U5967 (N_5967,N_4632,N_4400);
xor U5968 (N_5968,N_4108,N_4124);
xor U5969 (N_5969,N_4175,N_4023);
nor U5970 (N_5970,N_4042,N_4212);
xor U5971 (N_5971,N_4370,N_4789);
and U5972 (N_5972,N_4331,N_4966);
xor U5973 (N_5973,N_4351,N_4670);
and U5974 (N_5974,N_4080,N_4254);
or U5975 (N_5975,N_4976,N_4046);
xnor U5976 (N_5976,N_4614,N_4687);
and U5977 (N_5977,N_4444,N_4552);
xnor U5978 (N_5978,N_4272,N_4998);
nor U5979 (N_5979,N_4493,N_4373);
or U5980 (N_5980,N_4311,N_4105);
nor U5981 (N_5981,N_4831,N_4573);
nand U5982 (N_5982,N_4981,N_4772);
nand U5983 (N_5983,N_4111,N_4445);
and U5984 (N_5984,N_4126,N_4470);
and U5985 (N_5985,N_4926,N_4707);
nor U5986 (N_5986,N_4659,N_4256);
nand U5987 (N_5987,N_4348,N_4730);
xor U5988 (N_5988,N_4872,N_4361);
nand U5989 (N_5989,N_4732,N_4655);
nor U5990 (N_5990,N_4986,N_4087);
and U5991 (N_5991,N_4099,N_4002);
or U5992 (N_5992,N_4249,N_4995);
nand U5993 (N_5993,N_4088,N_4276);
nor U5994 (N_5994,N_4982,N_4432);
nor U5995 (N_5995,N_4966,N_4244);
nand U5996 (N_5996,N_4772,N_4093);
nor U5997 (N_5997,N_4066,N_4462);
xor U5998 (N_5998,N_4006,N_4126);
nor U5999 (N_5999,N_4877,N_4103);
nor U6000 (N_6000,N_5224,N_5912);
or U6001 (N_6001,N_5620,N_5583);
nor U6002 (N_6002,N_5877,N_5593);
and U6003 (N_6003,N_5367,N_5412);
and U6004 (N_6004,N_5848,N_5437);
or U6005 (N_6005,N_5610,N_5594);
nor U6006 (N_6006,N_5673,N_5530);
nor U6007 (N_6007,N_5774,N_5989);
nor U6008 (N_6008,N_5028,N_5664);
xor U6009 (N_6009,N_5871,N_5637);
nand U6010 (N_6010,N_5266,N_5581);
and U6011 (N_6011,N_5371,N_5201);
and U6012 (N_6012,N_5343,N_5385);
xnor U6013 (N_6013,N_5159,N_5426);
nand U6014 (N_6014,N_5298,N_5809);
xor U6015 (N_6015,N_5926,N_5952);
nor U6016 (N_6016,N_5671,N_5644);
xnor U6017 (N_6017,N_5779,N_5528);
xor U6018 (N_6018,N_5012,N_5265);
and U6019 (N_6019,N_5626,N_5937);
nor U6020 (N_6020,N_5969,N_5837);
or U6021 (N_6021,N_5320,N_5271);
nand U6022 (N_6022,N_5206,N_5104);
or U6023 (N_6023,N_5796,N_5638);
nor U6024 (N_6024,N_5460,N_5380);
and U6025 (N_6025,N_5465,N_5325);
and U6026 (N_6026,N_5139,N_5330);
nand U6027 (N_6027,N_5504,N_5949);
xnor U6028 (N_6028,N_5427,N_5772);
and U6029 (N_6029,N_5732,N_5753);
nand U6030 (N_6030,N_5592,N_5014);
nand U6031 (N_6031,N_5097,N_5739);
or U6032 (N_6032,N_5329,N_5037);
or U6033 (N_6033,N_5857,N_5264);
nor U6034 (N_6034,N_5934,N_5270);
xnor U6035 (N_6035,N_5656,N_5721);
and U6036 (N_6036,N_5020,N_5398);
and U6037 (N_6037,N_5282,N_5834);
or U6038 (N_6038,N_5983,N_5900);
nand U6039 (N_6039,N_5150,N_5720);
or U6040 (N_6040,N_5500,N_5596);
or U6041 (N_6041,N_5497,N_5021);
and U6042 (N_6042,N_5411,N_5617);
nand U6043 (N_6043,N_5468,N_5029);
nor U6044 (N_6044,N_5584,N_5285);
or U6045 (N_6045,N_5095,N_5278);
or U6046 (N_6046,N_5030,N_5601);
and U6047 (N_6047,N_5185,N_5523);
or U6048 (N_6048,N_5519,N_5706);
nand U6049 (N_6049,N_5647,N_5561);
nand U6050 (N_6050,N_5140,N_5247);
and U6051 (N_6051,N_5651,N_5047);
xor U6052 (N_6052,N_5907,N_5710);
and U6053 (N_6053,N_5711,N_5612);
and U6054 (N_6054,N_5171,N_5082);
xnor U6055 (N_6055,N_5853,N_5220);
xor U6056 (N_6056,N_5641,N_5597);
nor U6057 (N_6057,N_5935,N_5554);
or U6058 (N_6058,N_5052,N_5440);
nor U6059 (N_6059,N_5203,N_5214);
xor U6060 (N_6060,N_5870,N_5954);
nand U6061 (N_6061,N_5568,N_5199);
nor U6062 (N_6062,N_5628,N_5881);
nor U6063 (N_6063,N_5101,N_5485);
nor U6064 (N_6064,N_5443,N_5024);
or U6065 (N_6065,N_5961,N_5393);
and U6066 (N_6066,N_5927,N_5086);
nand U6067 (N_6067,N_5256,N_5215);
nor U6068 (N_6068,N_5654,N_5396);
xor U6069 (N_6069,N_5856,N_5174);
nor U6070 (N_6070,N_5876,N_5223);
nand U6071 (N_6071,N_5035,N_5337);
xor U6072 (N_6072,N_5280,N_5525);
or U6073 (N_6073,N_5130,N_5589);
nor U6074 (N_6074,N_5194,N_5867);
nor U6075 (N_6075,N_5763,N_5317);
nor U6076 (N_6076,N_5992,N_5375);
xnor U6077 (N_6077,N_5948,N_5232);
nand U6078 (N_6078,N_5294,N_5313);
xnor U6079 (N_6079,N_5421,N_5734);
or U6080 (N_6080,N_5824,N_5459);
and U6081 (N_6081,N_5365,N_5209);
or U6082 (N_6082,N_5061,N_5026);
xor U6083 (N_6083,N_5198,N_5308);
nand U6084 (N_6084,N_5335,N_5669);
nand U6085 (N_6085,N_5558,N_5297);
nor U6086 (N_6086,N_5914,N_5361);
nand U6087 (N_6087,N_5376,N_5213);
nor U6088 (N_6088,N_5234,N_5183);
nand U6089 (N_6089,N_5689,N_5865);
and U6090 (N_6090,N_5841,N_5652);
nand U6091 (N_6091,N_5540,N_5341);
or U6092 (N_6092,N_5931,N_5891);
and U6093 (N_6093,N_5143,N_5895);
nor U6094 (N_6094,N_5686,N_5515);
xor U6095 (N_6095,N_5177,N_5321);
nor U6096 (N_6096,N_5535,N_5748);
or U6097 (N_6097,N_5036,N_5648);
or U6098 (N_6098,N_5559,N_5586);
or U6099 (N_6099,N_5822,N_5988);
nand U6100 (N_6100,N_5532,N_5251);
nand U6101 (N_6101,N_5507,N_5608);
and U6102 (N_6102,N_5768,N_5148);
xnor U6103 (N_6103,N_5263,N_5718);
nand U6104 (N_6104,N_5114,N_5433);
and U6105 (N_6105,N_5039,N_5392);
or U6106 (N_6106,N_5667,N_5805);
and U6107 (N_6107,N_5042,N_5843);
nor U6108 (N_6108,N_5484,N_5708);
nor U6109 (N_6109,N_5033,N_5410);
nand U6110 (N_6110,N_5635,N_5336);
and U6111 (N_6111,N_5453,N_5132);
nand U6112 (N_6112,N_5339,N_5879);
or U6113 (N_6113,N_5501,N_5991);
xnor U6114 (N_6114,N_5588,N_5046);
or U6115 (N_6115,N_5603,N_5788);
xnor U6116 (N_6116,N_5133,N_5115);
or U6117 (N_6117,N_5878,N_5546);
xnor U6118 (N_6118,N_5899,N_5245);
or U6119 (N_6119,N_5893,N_5757);
nor U6120 (N_6120,N_5678,N_5406);
nor U6121 (N_6121,N_5575,N_5126);
and U6122 (N_6122,N_5996,N_5063);
or U6123 (N_6123,N_5242,N_5823);
or U6124 (N_6124,N_5461,N_5769);
or U6125 (N_6125,N_5249,N_5828);
or U6126 (N_6126,N_5653,N_5346);
nor U6127 (N_6127,N_5383,N_5373);
and U6128 (N_6128,N_5547,N_5128);
or U6129 (N_6129,N_5882,N_5299);
or U6130 (N_6130,N_5331,N_5563);
xor U6131 (N_6131,N_5976,N_5925);
nor U6132 (N_6132,N_5636,N_5087);
xor U6133 (N_6133,N_5690,N_5704);
nand U6134 (N_6134,N_5463,N_5395);
and U6135 (N_6135,N_5211,N_5707);
nand U6136 (N_6136,N_5075,N_5181);
nand U6137 (N_6137,N_5422,N_5712);
nor U6138 (N_6138,N_5923,N_5808);
or U6139 (N_6139,N_5851,N_5434);
xnor U6140 (N_6140,N_5649,N_5387);
or U6141 (N_6141,N_5627,N_5386);
xor U6142 (N_6142,N_5423,N_5231);
and U6143 (N_6143,N_5038,N_5781);
xor U6144 (N_6144,N_5197,N_5378);
or U6145 (N_6145,N_5116,N_5633);
and U6146 (N_6146,N_5972,N_5910);
or U6147 (N_6147,N_5283,N_5844);
nor U6148 (N_6148,N_5227,N_5917);
xnor U6149 (N_6149,N_5741,N_5714);
nand U6150 (N_6150,N_5866,N_5802);
nand U6151 (N_6151,N_5573,N_5191);
nand U6152 (N_6152,N_5785,N_5318);
and U6153 (N_6153,N_5362,N_5725);
nor U6154 (N_6154,N_5713,N_5659);
and U6155 (N_6155,N_5112,N_5152);
xnor U6156 (N_6156,N_5897,N_5531);
nand U6157 (N_6157,N_5163,N_5344);
nand U6158 (N_6158,N_5254,N_5155);
nand U6159 (N_6159,N_5314,N_5011);
xnor U6160 (N_6160,N_5074,N_5319);
xor U6161 (N_6161,N_5252,N_5451);
nor U6162 (N_6162,N_5908,N_5599);
or U6163 (N_6163,N_5517,N_5567);
and U6164 (N_6164,N_5326,N_5773);
nor U6165 (N_6165,N_5640,N_5244);
or U6166 (N_6166,N_5994,N_5354);
nand U6167 (N_6167,N_5068,N_5993);
or U6168 (N_6168,N_5005,N_5787);
or U6169 (N_6169,N_5407,N_5486);
nand U6170 (N_6170,N_5302,N_5555);
xor U6171 (N_6171,N_5216,N_5915);
or U6172 (N_6172,N_5842,N_5552);
nand U6173 (N_6173,N_5668,N_5212);
xnor U6174 (N_6174,N_5932,N_5797);
nor U6175 (N_6175,N_5815,N_5289);
or U6176 (N_6176,N_5716,N_5259);
xnor U6177 (N_6177,N_5456,N_5488);
nand U6178 (N_6178,N_5040,N_5444);
xnor U6179 (N_6179,N_5863,N_5023);
nand U6180 (N_6180,N_5675,N_5722);
xor U6181 (N_6181,N_5536,N_5402);
xnor U6182 (N_6182,N_5147,N_5997);
nor U6183 (N_6183,N_5831,N_5469);
and U6184 (N_6184,N_5253,N_5292);
and U6185 (N_6185,N_5982,N_5793);
or U6186 (N_6186,N_5775,N_5417);
or U6187 (N_6187,N_5390,N_5303);
nor U6188 (N_6188,N_5006,N_5724);
or U6189 (N_6189,N_5450,N_5142);
nand U6190 (N_6190,N_5009,N_5027);
xor U6191 (N_6191,N_5248,N_5790);
nand U6192 (N_6192,N_5795,N_5565);
nor U6193 (N_6193,N_5701,N_5677);
nand U6194 (N_6194,N_5749,N_5609);
xor U6195 (N_6195,N_5505,N_5829);
xor U6196 (N_6196,N_5069,N_5845);
nand U6197 (N_6197,N_5307,N_5906);
xor U6198 (N_6198,N_5901,N_5578);
xnor U6199 (N_6199,N_5262,N_5408);
nand U6200 (N_6200,N_5804,N_5207);
nor U6201 (N_6201,N_5974,N_5055);
nand U6202 (N_6202,N_5058,N_5551);
nand U6203 (N_6203,N_5043,N_5958);
xor U6204 (N_6204,N_5065,N_5623);
xnor U6205 (N_6205,N_5777,N_5514);
xnor U6206 (N_6206,N_5728,N_5674);
xor U6207 (N_6207,N_5481,N_5650);
nand U6208 (N_6208,N_5146,N_5840);
xor U6209 (N_6209,N_5117,N_5111);
xnor U6210 (N_6210,N_5498,N_5400);
xnor U6211 (N_6211,N_5864,N_5975);
nor U6212 (N_6212,N_5642,N_5660);
nand U6213 (N_6213,N_5875,N_5685);
nor U6214 (N_6214,N_5222,N_5079);
xor U6215 (N_6215,N_5476,N_5295);
nor U6216 (N_6216,N_5416,N_5607);
nand U6217 (N_6217,N_5742,N_5090);
nand U6218 (N_6218,N_5987,N_5602);
and U6219 (N_6219,N_5105,N_5963);
nor U6220 (N_6220,N_5817,N_5816);
nand U6221 (N_6221,N_5141,N_5765);
nor U6222 (N_6222,N_5273,N_5170);
nor U6223 (N_6223,N_5301,N_5323);
or U6224 (N_6224,N_5358,N_5819);
xor U6225 (N_6225,N_5272,N_5801);
nand U6226 (N_6226,N_5814,N_5920);
nor U6227 (N_6227,N_5577,N_5533);
nand U6228 (N_6228,N_5000,N_5957);
nand U6229 (N_6229,N_5869,N_5740);
nand U6230 (N_6230,N_5986,N_5447);
xor U6231 (N_6231,N_5962,N_5850);
nand U6232 (N_6232,N_5670,N_5695);
or U6233 (N_6233,N_5059,N_5127);
xnor U6234 (N_6234,N_5665,N_5480);
nor U6235 (N_6235,N_5727,N_5008);
xnor U6236 (N_6236,N_5619,N_5233);
and U6237 (N_6237,N_5680,N_5334);
and U6238 (N_6238,N_5598,N_5499);
xnor U6239 (N_6239,N_5250,N_5316);
xor U6240 (N_6240,N_5646,N_5569);
or U6241 (N_6241,N_5328,N_5467);
or U6242 (N_6242,N_5364,N_5089);
xor U6243 (N_6243,N_5322,N_5257);
nor U6244 (N_6244,N_5836,N_5445);
nand U6245 (N_6245,N_5703,N_5529);
nand U6246 (N_6246,N_5643,N_5930);
nand U6247 (N_6247,N_5968,N_5807);
nor U6248 (N_6248,N_5770,N_5605);
and U6249 (N_6249,N_5747,N_5189);
and U6250 (N_6250,N_5911,N_5003);
or U6251 (N_6251,N_5939,N_5399);
nor U6252 (N_6252,N_5093,N_5345);
nand U6253 (N_6253,N_5521,N_5579);
or U6254 (N_6254,N_5696,N_5506);
and U6255 (N_6255,N_5372,N_5752);
and U6256 (N_6256,N_5418,N_5355);
xor U6257 (N_6257,N_5631,N_5004);
xor U6258 (N_6258,N_5066,N_5419);
xor U6259 (N_6259,N_5810,N_5990);
or U6260 (N_6260,N_5491,N_5928);
xor U6261 (N_6261,N_5760,N_5096);
xnor U6262 (N_6262,N_5032,N_5125);
nand U6263 (N_6263,N_5566,N_5639);
or U6264 (N_6264,N_5085,N_5943);
nand U6265 (N_6265,N_5771,N_5479);
and U6266 (N_6266,N_5384,N_5800);
xnor U6267 (N_6267,N_5634,N_5622);
xnor U6268 (N_6268,N_5092,N_5527);
and U6269 (N_6269,N_5119,N_5913);
or U6270 (N_6270,N_5791,N_5590);
nand U6271 (N_6271,N_5347,N_5662);
or U6272 (N_6272,N_5679,N_5945);
or U6273 (N_6273,N_5156,N_5274);
nor U6274 (N_6274,N_5258,N_5230);
and U6275 (N_6275,N_5124,N_5629);
or U6276 (N_6276,N_5109,N_5539);
or U6277 (N_6277,N_5697,N_5475);
and U6278 (N_6278,N_5905,N_5381);
nor U6279 (N_6279,N_5509,N_5726);
xnor U6280 (N_6280,N_5998,N_5144);
or U6281 (N_6281,N_5762,N_5276);
and U6282 (N_6282,N_5938,N_5067);
and U6283 (N_6283,N_5839,N_5903);
nor U6284 (N_6284,N_5600,N_5859);
or U6285 (N_6285,N_5979,N_5102);
nand U6286 (N_6286,N_5415,N_5936);
nand U6287 (N_6287,N_5574,N_5830);
and U6288 (N_6288,N_5333,N_5783);
or U6289 (N_6289,N_5776,N_5267);
nand U6290 (N_6290,N_5489,N_5496);
nor U6291 (N_6291,N_5894,N_5835);
nand U6292 (N_6292,N_5526,N_5464);
xor U6293 (N_6293,N_5977,N_5072);
nor U6294 (N_6294,N_5502,N_5077);
nand U6295 (N_6295,N_5162,N_5136);
or U6296 (N_6296,N_5572,N_5268);
nor U6297 (N_6297,N_5188,N_5129);
or U6298 (N_6298,N_5798,N_5730);
xnor U6299 (N_6299,N_5946,N_5955);
and U6300 (N_6300,N_5478,N_5855);
xnor U6301 (N_6301,N_5890,N_5431);
nand U6302 (N_6302,N_5582,N_5657);
and U6303 (N_6303,N_5511,N_5786);
and U6304 (N_6304,N_5432,N_5942);
xnor U6305 (N_6305,N_5424,N_5366);
or U6306 (N_6306,N_5293,N_5379);
or U6307 (N_6307,N_5246,N_5820);
nor U6308 (N_6308,N_5767,N_5754);
and U6309 (N_6309,N_5918,N_5113);
nand U6310 (N_6310,N_5350,N_5442);
and U6311 (N_6311,N_5107,N_5239);
or U6312 (N_6312,N_5363,N_5898);
xnor U6313 (N_6313,N_5548,N_5782);
xnor U6314 (N_6314,N_5108,N_5359);
and U6315 (N_6315,N_5663,N_5924);
nand U6316 (N_6316,N_5780,N_5311);
or U6317 (N_6317,N_5007,N_5508);
xnor U6318 (N_6318,N_5073,N_5862);
and U6319 (N_6319,N_5176,N_5922);
or U6320 (N_6320,N_5175,N_5715);
nand U6321 (N_6321,N_5057,N_5449);
and U6322 (N_6322,N_5013,N_5202);
nor U6323 (N_6323,N_5545,N_5645);
nand U6324 (N_6324,N_5557,N_5351);
nand U6325 (N_6325,N_5076,N_5094);
and U6326 (N_6326,N_5761,N_5312);
nor U6327 (N_6327,N_5340,N_5692);
xor U6328 (N_6328,N_5064,N_5070);
and U6329 (N_6329,N_5699,N_5374);
or U6330 (N_6330,N_5960,N_5970);
nand U6331 (N_6331,N_5241,N_5016);
xor U6332 (N_6332,N_5436,N_5847);
nor U6333 (N_6333,N_5041,N_5457);
or U6334 (N_6334,N_5737,N_5861);
nand U6335 (N_6335,N_5522,N_5495);
and U6336 (N_6336,N_5487,N_5022);
and U6337 (N_6337,N_5414,N_5173);
and U6338 (N_6338,N_5860,N_5613);
and U6339 (N_6339,N_5404,N_5138);
nand U6340 (N_6340,N_5389,N_5606);
xnor U6341 (N_6341,N_5624,N_5719);
and U6342 (N_6342,N_5980,N_5852);
or U6343 (N_6343,N_5219,N_5439);
nor U6344 (N_6344,N_5691,N_5435);
nor U6345 (N_6345,N_5360,N_5483);
nand U6346 (N_6346,N_5818,N_5492);
and U6347 (N_6347,N_5060,N_5315);
nand U6348 (N_6348,N_5929,N_5493);
and U6349 (N_6349,N_5338,N_5078);
nor U6350 (N_6350,N_5056,N_5287);
or U6351 (N_6351,N_5062,N_5179);
nand U6352 (N_6352,N_5904,N_5580);
xor U6353 (N_6353,N_5001,N_5698);
nor U6354 (N_6354,N_5812,N_5813);
and U6355 (N_6355,N_5332,N_5959);
xnor U6356 (N_6356,N_5615,N_5966);
nand U6357 (N_6357,N_5661,N_5953);
nor U6358 (N_6358,N_5121,N_5403);
or U6359 (N_6359,N_5981,N_5534);
and U6360 (N_6360,N_5088,N_5193);
nand U6361 (N_6361,N_5131,N_5357);
nand U6362 (N_6362,N_5441,N_5542);
nor U6363 (N_6363,N_5025,N_5208);
xnor U6364 (N_6364,N_5071,N_5100);
nand U6365 (N_6365,N_5755,N_5587);
nand U6366 (N_6366,N_5420,N_5053);
nand U6367 (N_6367,N_5083,N_5243);
and U6368 (N_6368,N_5145,N_5512);
xnor U6369 (N_6369,N_5688,N_5886);
nor U6370 (N_6370,N_5169,N_5585);
nor U6371 (N_6371,N_5304,N_5106);
nand U6372 (N_6372,N_5919,N_5494);
xor U6373 (N_6373,N_5799,N_5549);
and U6374 (N_6374,N_5458,N_5541);
nor U6375 (N_6375,N_5833,N_5228);
nor U6376 (N_6376,N_5591,N_5944);
nor U6377 (N_6377,N_5240,N_5611);
nor U6378 (N_6378,N_5448,N_5377);
nand U6379 (N_6379,N_5368,N_5570);
nand U6380 (N_6380,N_5401,N_5382);
nor U6381 (N_6381,N_5195,N_5310);
nor U6382 (N_6382,N_5178,N_5091);
nor U6383 (N_6383,N_5672,N_5160);
nor U6384 (N_6384,N_5999,N_5811);
and U6385 (N_6385,N_5562,N_5743);
xor U6386 (N_6386,N_5888,N_5482);
and U6387 (N_6387,N_5327,N_5868);
xor U6388 (N_6388,N_5034,N_5872);
nand U6389 (N_6389,N_5621,N_5172);
xor U6390 (N_6390,N_5909,N_5151);
and U6391 (N_6391,N_5655,N_5235);
and U6392 (N_6392,N_5275,N_5827);
xnor U6393 (N_6393,N_5700,N_5604);
or U6394 (N_6394,N_5054,N_5731);
nand U6395 (N_6395,N_5889,N_5683);
and U6396 (N_6396,N_5666,N_5744);
nand U6397 (N_6397,N_5658,N_5941);
xnor U6398 (N_6398,N_5348,N_5709);
or U6399 (N_6399,N_5503,N_5305);
nor U6400 (N_6400,N_5951,N_5735);
xnor U6401 (N_6401,N_5784,N_5123);
nand U6402 (N_6402,N_5550,N_5538);
nor U6403 (N_6403,N_5553,N_5269);
or U6404 (N_6404,N_5792,N_5759);
nor U6405 (N_6405,N_5225,N_5425);
xnor U6406 (N_6406,N_5324,N_5884);
nand U6407 (N_6407,N_5524,N_5099);
or U6408 (N_6408,N_5288,N_5751);
xor U6409 (N_6409,N_5520,N_5750);
nand U6410 (N_6410,N_5154,N_5940);
nor U6411 (N_6411,N_5002,N_5196);
and U6412 (N_6412,N_5756,N_5217);
and U6413 (N_6413,N_5806,N_5510);
or U6414 (N_6414,N_5702,N_5161);
or U6415 (N_6415,N_5564,N_5184);
xnor U6416 (N_6416,N_5238,N_5630);
nand U6417 (N_6417,N_5205,N_5736);
nor U6418 (N_6418,N_5764,N_5705);
xor U6419 (N_6419,N_5854,N_5513);
xor U6420 (N_6420,N_5164,N_5985);
or U6421 (N_6421,N_5103,N_5192);
nand U6422 (N_6422,N_5200,N_5738);
xor U6423 (N_6423,N_5284,N_5973);
or U6424 (N_6424,N_5044,N_5165);
nor U6425 (N_6425,N_5045,N_5694);
nand U6426 (N_6426,N_5281,N_5846);
nand U6427 (N_6427,N_5018,N_5356);
or U6428 (N_6428,N_5353,N_5153);
xor U6429 (N_6429,N_5186,N_5210);
nand U6430 (N_6430,N_5017,N_5682);
or U6431 (N_6431,N_5157,N_5237);
nor U6432 (N_6432,N_5995,N_5430);
or U6433 (N_6433,N_5556,N_5470);
nand U6434 (N_6434,N_5477,N_5277);
nor U6435 (N_6435,N_5428,N_5204);
and U6436 (N_6436,N_5286,N_5049);
nand U6437 (N_6437,N_5902,N_5964);
xnor U6438 (N_6438,N_5388,N_5462);
and U6439 (N_6439,N_5291,N_5454);
or U6440 (N_6440,N_5084,N_5723);
xnor U6441 (N_6441,N_5614,N_5618);
nand U6442 (N_6442,N_5978,N_5729);
nor U6443 (N_6443,N_5019,N_5544);
nor U6444 (N_6444,N_5352,N_5409);
nor U6445 (N_6445,N_5342,N_5050);
or U6446 (N_6446,N_5182,N_5733);
nor U6447 (N_6447,N_5838,N_5261);
nor U6448 (N_6448,N_5405,N_5825);
xor U6449 (N_6449,N_5221,N_5290);
nor U6450 (N_6450,N_5632,N_5168);
or U6451 (N_6451,N_5394,N_5789);
or U6452 (N_6452,N_5296,N_5516);
or U6453 (N_6453,N_5137,N_5260);
and U6454 (N_6454,N_5560,N_5950);
xnor U6455 (N_6455,N_5255,N_5167);
nor U6456 (N_6456,N_5180,N_5446);
nor U6457 (N_6457,N_5300,N_5933);
and U6458 (N_6458,N_5832,N_5616);
nand U6459 (N_6459,N_5874,N_5110);
or U6460 (N_6460,N_5120,N_5472);
and U6461 (N_6461,N_5821,N_5571);
nor U6462 (N_6462,N_5681,N_5826);
nor U6463 (N_6463,N_5693,N_5676);
nor U6464 (N_6464,N_5518,N_5391);
and U6465 (N_6465,N_5048,N_5947);
and U6466 (N_6466,N_5438,N_5218);
and U6467 (N_6467,N_5595,N_5803);
and U6468 (N_6468,N_5490,N_5122);
or U6469 (N_6469,N_5916,N_5537);
xor U6470 (N_6470,N_5397,N_5226);
nor U6471 (N_6471,N_5965,N_5455);
xor U6472 (N_6472,N_5031,N_5745);
and U6473 (N_6473,N_5717,N_5306);
nor U6474 (N_6474,N_5081,N_5885);
nor U6475 (N_6475,N_5051,N_5880);
or U6476 (N_6476,N_5625,N_5956);
and U6477 (N_6477,N_5984,N_5015);
nand U6478 (N_6478,N_5190,N_5766);
nand U6479 (N_6479,N_5474,N_5778);
or U6480 (N_6480,N_5187,N_5921);
nand U6481 (N_6481,N_5471,N_5429);
nor U6482 (N_6482,N_5746,N_5118);
and U6483 (N_6483,N_5971,N_5883);
and U6484 (N_6484,N_5158,N_5236);
nand U6485 (N_6485,N_5576,N_5349);
nand U6486 (N_6486,N_5080,N_5896);
xnor U6487 (N_6487,N_5279,N_5873);
or U6488 (N_6488,N_5010,N_5887);
or U6489 (N_6489,N_5413,N_5134);
or U6490 (N_6490,N_5166,N_5149);
nor U6491 (N_6491,N_5370,N_5135);
nor U6492 (N_6492,N_5967,N_5098);
xnor U6493 (N_6493,N_5229,N_5466);
nor U6494 (N_6494,N_5858,N_5794);
and U6495 (N_6495,N_5849,N_5687);
nor U6496 (N_6496,N_5543,N_5892);
and U6497 (N_6497,N_5309,N_5369);
nor U6498 (N_6498,N_5684,N_5452);
xor U6499 (N_6499,N_5473,N_5758);
and U6500 (N_6500,N_5480,N_5444);
xnor U6501 (N_6501,N_5054,N_5449);
xnor U6502 (N_6502,N_5659,N_5529);
nand U6503 (N_6503,N_5167,N_5966);
nand U6504 (N_6504,N_5235,N_5670);
or U6505 (N_6505,N_5417,N_5617);
nand U6506 (N_6506,N_5329,N_5706);
nand U6507 (N_6507,N_5280,N_5996);
xnor U6508 (N_6508,N_5897,N_5815);
nand U6509 (N_6509,N_5503,N_5620);
xnor U6510 (N_6510,N_5935,N_5572);
or U6511 (N_6511,N_5967,N_5596);
nand U6512 (N_6512,N_5906,N_5983);
or U6513 (N_6513,N_5417,N_5254);
or U6514 (N_6514,N_5056,N_5961);
xor U6515 (N_6515,N_5772,N_5370);
nand U6516 (N_6516,N_5006,N_5241);
or U6517 (N_6517,N_5495,N_5870);
or U6518 (N_6518,N_5171,N_5242);
xnor U6519 (N_6519,N_5399,N_5160);
nor U6520 (N_6520,N_5521,N_5998);
and U6521 (N_6521,N_5199,N_5894);
and U6522 (N_6522,N_5594,N_5801);
nand U6523 (N_6523,N_5133,N_5494);
or U6524 (N_6524,N_5108,N_5683);
nor U6525 (N_6525,N_5009,N_5930);
nor U6526 (N_6526,N_5609,N_5362);
nor U6527 (N_6527,N_5285,N_5677);
xor U6528 (N_6528,N_5674,N_5015);
xnor U6529 (N_6529,N_5977,N_5690);
or U6530 (N_6530,N_5541,N_5911);
nor U6531 (N_6531,N_5083,N_5840);
xnor U6532 (N_6532,N_5009,N_5432);
nand U6533 (N_6533,N_5300,N_5508);
or U6534 (N_6534,N_5274,N_5026);
and U6535 (N_6535,N_5694,N_5548);
xor U6536 (N_6536,N_5911,N_5567);
or U6537 (N_6537,N_5592,N_5786);
or U6538 (N_6538,N_5496,N_5038);
nor U6539 (N_6539,N_5719,N_5024);
and U6540 (N_6540,N_5503,N_5607);
and U6541 (N_6541,N_5611,N_5319);
nor U6542 (N_6542,N_5525,N_5582);
xor U6543 (N_6543,N_5088,N_5602);
and U6544 (N_6544,N_5180,N_5677);
nand U6545 (N_6545,N_5817,N_5155);
nand U6546 (N_6546,N_5294,N_5590);
nor U6547 (N_6547,N_5057,N_5893);
and U6548 (N_6548,N_5443,N_5889);
and U6549 (N_6549,N_5025,N_5245);
nand U6550 (N_6550,N_5563,N_5623);
and U6551 (N_6551,N_5267,N_5493);
and U6552 (N_6552,N_5927,N_5628);
or U6553 (N_6553,N_5152,N_5913);
and U6554 (N_6554,N_5430,N_5731);
nand U6555 (N_6555,N_5450,N_5898);
or U6556 (N_6556,N_5280,N_5824);
nand U6557 (N_6557,N_5272,N_5664);
xor U6558 (N_6558,N_5830,N_5336);
or U6559 (N_6559,N_5214,N_5720);
and U6560 (N_6560,N_5395,N_5681);
or U6561 (N_6561,N_5296,N_5446);
xnor U6562 (N_6562,N_5938,N_5530);
xor U6563 (N_6563,N_5992,N_5641);
and U6564 (N_6564,N_5590,N_5372);
or U6565 (N_6565,N_5001,N_5796);
and U6566 (N_6566,N_5541,N_5755);
or U6567 (N_6567,N_5720,N_5735);
nor U6568 (N_6568,N_5239,N_5486);
xnor U6569 (N_6569,N_5134,N_5983);
nand U6570 (N_6570,N_5841,N_5443);
or U6571 (N_6571,N_5622,N_5002);
or U6572 (N_6572,N_5368,N_5009);
or U6573 (N_6573,N_5325,N_5715);
or U6574 (N_6574,N_5021,N_5911);
nor U6575 (N_6575,N_5984,N_5937);
and U6576 (N_6576,N_5910,N_5187);
nand U6577 (N_6577,N_5471,N_5770);
xnor U6578 (N_6578,N_5246,N_5774);
or U6579 (N_6579,N_5044,N_5815);
xnor U6580 (N_6580,N_5273,N_5182);
and U6581 (N_6581,N_5143,N_5400);
and U6582 (N_6582,N_5449,N_5241);
xor U6583 (N_6583,N_5846,N_5090);
nand U6584 (N_6584,N_5227,N_5264);
nand U6585 (N_6585,N_5778,N_5300);
xor U6586 (N_6586,N_5489,N_5474);
xnor U6587 (N_6587,N_5232,N_5840);
or U6588 (N_6588,N_5871,N_5766);
and U6589 (N_6589,N_5656,N_5605);
nor U6590 (N_6590,N_5658,N_5344);
xnor U6591 (N_6591,N_5861,N_5250);
nor U6592 (N_6592,N_5189,N_5414);
or U6593 (N_6593,N_5344,N_5071);
or U6594 (N_6594,N_5936,N_5555);
or U6595 (N_6595,N_5567,N_5807);
nor U6596 (N_6596,N_5427,N_5654);
and U6597 (N_6597,N_5484,N_5976);
or U6598 (N_6598,N_5067,N_5270);
and U6599 (N_6599,N_5628,N_5227);
nor U6600 (N_6600,N_5509,N_5358);
xnor U6601 (N_6601,N_5116,N_5487);
nor U6602 (N_6602,N_5061,N_5271);
or U6603 (N_6603,N_5249,N_5112);
xor U6604 (N_6604,N_5706,N_5435);
xor U6605 (N_6605,N_5697,N_5229);
xor U6606 (N_6606,N_5641,N_5677);
or U6607 (N_6607,N_5799,N_5356);
and U6608 (N_6608,N_5841,N_5586);
xnor U6609 (N_6609,N_5239,N_5657);
nand U6610 (N_6610,N_5616,N_5716);
and U6611 (N_6611,N_5274,N_5455);
or U6612 (N_6612,N_5984,N_5431);
xor U6613 (N_6613,N_5076,N_5544);
and U6614 (N_6614,N_5462,N_5550);
nor U6615 (N_6615,N_5895,N_5514);
nor U6616 (N_6616,N_5436,N_5206);
xnor U6617 (N_6617,N_5333,N_5138);
nand U6618 (N_6618,N_5745,N_5412);
xor U6619 (N_6619,N_5270,N_5658);
nor U6620 (N_6620,N_5342,N_5143);
and U6621 (N_6621,N_5742,N_5953);
and U6622 (N_6622,N_5439,N_5371);
and U6623 (N_6623,N_5023,N_5807);
nor U6624 (N_6624,N_5709,N_5863);
xor U6625 (N_6625,N_5816,N_5716);
and U6626 (N_6626,N_5664,N_5070);
and U6627 (N_6627,N_5804,N_5425);
or U6628 (N_6628,N_5408,N_5976);
or U6629 (N_6629,N_5114,N_5205);
nor U6630 (N_6630,N_5305,N_5572);
or U6631 (N_6631,N_5187,N_5697);
or U6632 (N_6632,N_5383,N_5544);
or U6633 (N_6633,N_5920,N_5018);
xnor U6634 (N_6634,N_5899,N_5426);
xor U6635 (N_6635,N_5561,N_5648);
xnor U6636 (N_6636,N_5732,N_5989);
and U6637 (N_6637,N_5272,N_5127);
or U6638 (N_6638,N_5588,N_5665);
nand U6639 (N_6639,N_5995,N_5470);
and U6640 (N_6640,N_5082,N_5335);
or U6641 (N_6641,N_5941,N_5328);
nand U6642 (N_6642,N_5910,N_5487);
or U6643 (N_6643,N_5550,N_5328);
nand U6644 (N_6644,N_5096,N_5528);
or U6645 (N_6645,N_5851,N_5346);
nand U6646 (N_6646,N_5039,N_5184);
xor U6647 (N_6647,N_5328,N_5323);
or U6648 (N_6648,N_5654,N_5246);
nor U6649 (N_6649,N_5948,N_5942);
nor U6650 (N_6650,N_5846,N_5142);
nand U6651 (N_6651,N_5650,N_5629);
or U6652 (N_6652,N_5290,N_5449);
or U6653 (N_6653,N_5098,N_5331);
or U6654 (N_6654,N_5574,N_5399);
nand U6655 (N_6655,N_5763,N_5578);
nor U6656 (N_6656,N_5981,N_5548);
nor U6657 (N_6657,N_5286,N_5019);
or U6658 (N_6658,N_5188,N_5025);
or U6659 (N_6659,N_5036,N_5341);
nand U6660 (N_6660,N_5638,N_5349);
nor U6661 (N_6661,N_5796,N_5340);
nand U6662 (N_6662,N_5595,N_5893);
and U6663 (N_6663,N_5077,N_5261);
xnor U6664 (N_6664,N_5900,N_5455);
nand U6665 (N_6665,N_5664,N_5745);
xor U6666 (N_6666,N_5673,N_5325);
xor U6667 (N_6667,N_5515,N_5598);
and U6668 (N_6668,N_5170,N_5584);
nor U6669 (N_6669,N_5784,N_5807);
and U6670 (N_6670,N_5729,N_5345);
nor U6671 (N_6671,N_5386,N_5469);
or U6672 (N_6672,N_5373,N_5384);
and U6673 (N_6673,N_5028,N_5686);
or U6674 (N_6674,N_5876,N_5845);
nor U6675 (N_6675,N_5942,N_5211);
and U6676 (N_6676,N_5374,N_5195);
nand U6677 (N_6677,N_5929,N_5544);
nand U6678 (N_6678,N_5355,N_5948);
nor U6679 (N_6679,N_5362,N_5794);
and U6680 (N_6680,N_5550,N_5205);
xnor U6681 (N_6681,N_5136,N_5500);
or U6682 (N_6682,N_5227,N_5072);
or U6683 (N_6683,N_5719,N_5394);
nand U6684 (N_6684,N_5970,N_5666);
or U6685 (N_6685,N_5387,N_5130);
and U6686 (N_6686,N_5098,N_5731);
and U6687 (N_6687,N_5827,N_5154);
nor U6688 (N_6688,N_5738,N_5103);
and U6689 (N_6689,N_5291,N_5522);
xnor U6690 (N_6690,N_5820,N_5381);
nand U6691 (N_6691,N_5809,N_5755);
nor U6692 (N_6692,N_5923,N_5508);
xor U6693 (N_6693,N_5468,N_5293);
xor U6694 (N_6694,N_5745,N_5234);
or U6695 (N_6695,N_5802,N_5175);
and U6696 (N_6696,N_5265,N_5552);
or U6697 (N_6697,N_5823,N_5845);
or U6698 (N_6698,N_5180,N_5351);
or U6699 (N_6699,N_5468,N_5429);
or U6700 (N_6700,N_5324,N_5110);
and U6701 (N_6701,N_5368,N_5128);
nand U6702 (N_6702,N_5388,N_5354);
nand U6703 (N_6703,N_5944,N_5436);
or U6704 (N_6704,N_5722,N_5909);
and U6705 (N_6705,N_5564,N_5738);
nor U6706 (N_6706,N_5552,N_5512);
or U6707 (N_6707,N_5262,N_5978);
and U6708 (N_6708,N_5766,N_5354);
nand U6709 (N_6709,N_5209,N_5583);
nor U6710 (N_6710,N_5590,N_5667);
or U6711 (N_6711,N_5651,N_5779);
nand U6712 (N_6712,N_5130,N_5214);
nor U6713 (N_6713,N_5199,N_5824);
or U6714 (N_6714,N_5315,N_5988);
xor U6715 (N_6715,N_5293,N_5755);
or U6716 (N_6716,N_5140,N_5384);
or U6717 (N_6717,N_5440,N_5620);
xnor U6718 (N_6718,N_5715,N_5019);
xor U6719 (N_6719,N_5302,N_5603);
xnor U6720 (N_6720,N_5057,N_5433);
and U6721 (N_6721,N_5373,N_5431);
nor U6722 (N_6722,N_5499,N_5079);
nand U6723 (N_6723,N_5527,N_5722);
xor U6724 (N_6724,N_5616,N_5939);
and U6725 (N_6725,N_5778,N_5478);
nand U6726 (N_6726,N_5870,N_5278);
nor U6727 (N_6727,N_5419,N_5868);
nor U6728 (N_6728,N_5301,N_5690);
xnor U6729 (N_6729,N_5458,N_5938);
xnor U6730 (N_6730,N_5070,N_5816);
and U6731 (N_6731,N_5720,N_5063);
or U6732 (N_6732,N_5313,N_5955);
nor U6733 (N_6733,N_5477,N_5517);
and U6734 (N_6734,N_5040,N_5349);
nor U6735 (N_6735,N_5028,N_5763);
nand U6736 (N_6736,N_5539,N_5307);
nor U6737 (N_6737,N_5889,N_5399);
nor U6738 (N_6738,N_5077,N_5410);
xnor U6739 (N_6739,N_5671,N_5734);
or U6740 (N_6740,N_5459,N_5821);
or U6741 (N_6741,N_5675,N_5822);
nand U6742 (N_6742,N_5019,N_5492);
and U6743 (N_6743,N_5335,N_5734);
nor U6744 (N_6744,N_5746,N_5546);
nor U6745 (N_6745,N_5979,N_5098);
nand U6746 (N_6746,N_5527,N_5308);
nor U6747 (N_6747,N_5813,N_5059);
xor U6748 (N_6748,N_5073,N_5836);
or U6749 (N_6749,N_5499,N_5358);
xnor U6750 (N_6750,N_5350,N_5962);
nor U6751 (N_6751,N_5028,N_5669);
and U6752 (N_6752,N_5539,N_5240);
nand U6753 (N_6753,N_5371,N_5000);
nor U6754 (N_6754,N_5504,N_5438);
nand U6755 (N_6755,N_5755,N_5913);
or U6756 (N_6756,N_5956,N_5659);
or U6757 (N_6757,N_5244,N_5057);
and U6758 (N_6758,N_5212,N_5433);
nand U6759 (N_6759,N_5324,N_5456);
xnor U6760 (N_6760,N_5893,N_5724);
nand U6761 (N_6761,N_5056,N_5274);
and U6762 (N_6762,N_5679,N_5487);
nand U6763 (N_6763,N_5771,N_5816);
nor U6764 (N_6764,N_5017,N_5585);
or U6765 (N_6765,N_5571,N_5291);
nand U6766 (N_6766,N_5469,N_5756);
nand U6767 (N_6767,N_5672,N_5085);
nor U6768 (N_6768,N_5259,N_5895);
nand U6769 (N_6769,N_5728,N_5549);
nor U6770 (N_6770,N_5909,N_5347);
nor U6771 (N_6771,N_5040,N_5940);
or U6772 (N_6772,N_5759,N_5948);
nand U6773 (N_6773,N_5280,N_5075);
and U6774 (N_6774,N_5327,N_5980);
and U6775 (N_6775,N_5320,N_5824);
nor U6776 (N_6776,N_5917,N_5639);
and U6777 (N_6777,N_5547,N_5054);
xor U6778 (N_6778,N_5179,N_5002);
nor U6779 (N_6779,N_5156,N_5366);
xor U6780 (N_6780,N_5168,N_5491);
nand U6781 (N_6781,N_5320,N_5473);
nand U6782 (N_6782,N_5543,N_5353);
or U6783 (N_6783,N_5266,N_5623);
nand U6784 (N_6784,N_5888,N_5409);
nor U6785 (N_6785,N_5145,N_5147);
or U6786 (N_6786,N_5481,N_5489);
and U6787 (N_6787,N_5079,N_5596);
nor U6788 (N_6788,N_5213,N_5144);
nor U6789 (N_6789,N_5368,N_5380);
nand U6790 (N_6790,N_5292,N_5437);
nand U6791 (N_6791,N_5639,N_5474);
nand U6792 (N_6792,N_5328,N_5501);
nand U6793 (N_6793,N_5800,N_5049);
or U6794 (N_6794,N_5855,N_5306);
and U6795 (N_6795,N_5888,N_5488);
and U6796 (N_6796,N_5078,N_5349);
or U6797 (N_6797,N_5039,N_5582);
or U6798 (N_6798,N_5541,N_5671);
nand U6799 (N_6799,N_5576,N_5650);
nor U6800 (N_6800,N_5810,N_5043);
nand U6801 (N_6801,N_5997,N_5800);
and U6802 (N_6802,N_5889,N_5379);
nor U6803 (N_6803,N_5638,N_5663);
nand U6804 (N_6804,N_5587,N_5166);
nand U6805 (N_6805,N_5624,N_5831);
nand U6806 (N_6806,N_5418,N_5543);
nor U6807 (N_6807,N_5438,N_5324);
nand U6808 (N_6808,N_5143,N_5223);
nand U6809 (N_6809,N_5185,N_5308);
nand U6810 (N_6810,N_5203,N_5951);
nand U6811 (N_6811,N_5233,N_5550);
xor U6812 (N_6812,N_5483,N_5162);
and U6813 (N_6813,N_5796,N_5446);
nand U6814 (N_6814,N_5714,N_5713);
and U6815 (N_6815,N_5786,N_5938);
or U6816 (N_6816,N_5286,N_5550);
or U6817 (N_6817,N_5370,N_5663);
nor U6818 (N_6818,N_5450,N_5365);
nor U6819 (N_6819,N_5568,N_5112);
nand U6820 (N_6820,N_5528,N_5090);
or U6821 (N_6821,N_5230,N_5263);
and U6822 (N_6822,N_5071,N_5067);
xnor U6823 (N_6823,N_5406,N_5960);
xnor U6824 (N_6824,N_5711,N_5002);
nand U6825 (N_6825,N_5104,N_5272);
xor U6826 (N_6826,N_5978,N_5846);
nor U6827 (N_6827,N_5232,N_5346);
xor U6828 (N_6828,N_5111,N_5096);
and U6829 (N_6829,N_5762,N_5503);
and U6830 (N_6830,N_5262,N_5776);
nor U6831 (N_6831,N_5335,N_5530);
or U6832 (N_6832,N_5043,N_5748);
or U6833 (N_6833,N_5308,N_5528);
or U6834 (N_6834,N_5060,N_5554);
and U6835 (N_6835,N_5327,N_5736);
or U6836 (N_6836,N_5677,N_5544);
nor U6837 (N_6837,N_5830,N_5419);
nand U6838 (N_6838,N_5811,N_5365);
nand U6839 (N_6839,N_5236,N_5793);
xnor U6840 (N_6840,N_5968,N_5537);
or U6841 (N_6841,N_5920,N_5942);
and U6842 (N_6842,N_5752,N_5619);
nand U6843 (N_6843,N_5029,N_5837);
or U6844 (N_6844,N_5379,N_5394);
xor U6845 (N_6845,N_5309,N_5659);
nor U6846 (N_6846,N_5638,N_5406);
and U6847 (N_6847,N_5613,N_5009);
or U6848 (N_6848,N_5121,N_5874);
xor U6849 (N_6849,N_5770,N_5366);
nand U6850 (N_6850,N_5479,N_5279);
nand U6851 (N_6851,N_5988,N_5235);
and U6852 (N_6852,N_5365,N_5160);
xor U6853 (N_6853,N_5346,N_5784);
and U6854 (N_6854,N_5944,N_5549);
nor U6855 (N_6855,N_5573,N_5015);
nand U6856 (N_6856,N_5397,N_5489);
and U6857 (N_6857,N_5139,N_5585);
xnor U6858 (N_6858,N_5150,N_5471);
and U6859 (N_6859,N_5589,N_5566);
nor U6860 (N_6860,N_5081,N_5477);
nand U6861 (N_6861,N_5412,N_5986);
nor U6862 (N_6862,N_5711,N_5654);
xnor U6863 (N_6863,N_5439,N_5362);
and U6864 (N_6864,N_5962,N_5713);
nand U6865 (N_6865,N_5308,N_5272);
nor U6866 (N_6866,N_5840,N_5212);
and U6867 (N_6867,N_5978,N_5904);
and U6868 (N_6868,N_5299,N_5541);
nand U6869 (N_6869,N_5767,N_5513);
nand U6870 (N_6870,N_5759,N_5418);
xor U6871 (N_6871,N_5949,N_5742);
nor U6872 (N_6872,N_5040,N_5381);
nor U6873 (N_6873,N_5366,N_5579);
xor U6874 (N_6874,N_5556,N_5570);
nand U6875 (N_6875,N_5623,N_5456);
nand U6876 (N_6876,N_5708,N_5779);
nand U6877 (N_6877,N_5163,N_5296);
and U6878 (N_6878,N_5221,N_5156);
xor U6879 (N_6879,N_5002,N_5850);
nor U6880 (N_6880,N_5034,N_5660);
and U6881 (N_6881,N_5051,N_5020);
and U6882 (N_6882,N_5719,N_5418);
xor U6883 (N_6883,N_5003,N_5077);
nand U6884 (N_6884,N_5213,N_5761);
xor U6885 (N_6885,N_5709,N_5714);
xnor U6886 (N_6886,N_5128,N_5820);
or U6887 (N_6887,N_5226,N_5611);
nor U6888 (N_6888,N_5878,N_5165);
and U6889 (N_6889,N_5867,N_5433);
and U6890 (N_6890,N_5710,N_5295);
and U6891 (N_6891,N_5069,N_5087);
nand U6892 (N_6892,N_5028,N_5183);
xor U6893 (N_6893,N_5248,N_5178);
and U6894 (N_6894,N_5033,N_5403);
nand U6895 (N_6895,N_5096,N_5648);
or U6896 (N_6896,N_5440,N_5122);
nand U6897 (N_6897,N_5413,N_5182);
nand U6898 (N_6898,N_5493,N_5503);
or U6899 (N_6899,N_5362,N_5806);
nand U6900 (N_6900,N_5910,N_5412);
xnor U6901 (N_6901,N_5232,N_5265);
and U6902 (N_6902,N_5271,N_5235);
and U6903 (N_6903,N_5434,N_5950);
xor U6904 (N_6904,N_5988,N_5966);
or U6905 (N_6905,N_5921,N_5937);
xnor U6906 (N_6906,N_5791,N_5808);
and U6907 (N_6907,N_5759,N_5625);
or U6908 (N_6908,N_5504,N_5439);
nand U6909 (N_6909,N_5303,N_5882);
or U6910 (N_6910,N_5255,N_5550);
xor U6911 (N_6911,N_5682,N_5437);
nand U6912 (N_6912,N_5388,N_5147);
nand U6913 (N_6913,N_5323,N_5183);
xor U6914 (N_6914,N_5543,N_5969);
and U6915 (N_6915,N_5774,N_5351);
xor U6916 (N_6916,N_5122,N_5957);
nand U6917 (N_6917,N_5827,N_5139);
xor U6918 (N_6918,N_5154,N_5810);
xnor U6919 (N_6919,N_5305,N_5192);
and U6920 (N_6920,N_5325,N_5437);
nor U6921 (N_6921,N_5592,N_5398);
nor U6922 (N_6922,N_5351,N_5204);
or U6923 (N_6923,N_5348,N_5558);
xnor U6924 (N_6924,N_5423,N_5978);
and U6925 (N_6925,N_5635,N_5628);
or U6926 (N_6926,N_5149,N_5064);
and U6927 (N_6927,N_5970,N_5754);
xnor U6928 (N_6928,N_5087,N_5329);
and U6929 (N_6929,N_5465,N_5450);
and U6930 (N_6930,N_5785,N_5344);
nand U6931 (N_6931,N_5112,N_5182);
and U6932 (N_6932,N_5953,N_5932);
and U6933 (N_6933,N_5817,N_5749);
or U6934 (N_6934,N_5731,N_5798);
nand U6935 (N_6935,N_5783,N_5799);
nor U6936 (N_6936,N_5875,N_5681);
xnor U6937 (N_6937,N_5730,N_5043);
xor U6938 (N_6938,N_5254,N_5507);
and U6939 (N_6939,N_5985,N_5656);
or U6940 (N_6940,N_5425,N_5798);
xor U6941 (N_6941,N_5642,N_5847);
nor U6942 (N_6942,N_5071,N_5146);
nand U6943 (N_6943,N_5708,N_5555);
or U6944 (N_6944,N_5893,N_5380);
nand U6945 (N_6945,N_5071,N_5017);
nor U6946 (N_6946,N_5957,N_5302);
and U6947 (N_6947,N_5400,N_5696);
nand U6948 (N_6948,N_5059,N_5979);
nor U6949 (N_6949,N_5975,N_5630);
nand U6950 (N_6950,N_5909,N_5868);
xor U6951 (N_6951,N_5844,N_5757);
nor U6952 (N_6952,N_5779,N_5491);
or U6953 (N_6953,N_5994,N_5992);
nand U6954 (N_6954,N_5214,N_5235);
or U6955 (N_6955,N_5199,N_5421);
or U6956 (N_6956,N_5085,N_5894);
and U6957 (N_6957,N_5290,N_5003);
and U6958 (N_6958,N_5183,N_5899);
or U6959 (N_6959,N_5705,N_5595);
xor U6960 (N_6960,N_5066,N_5004);
or U6961 (N_6961,N_5903,N_5174);
and U6962 (N_6962,N_5869,N_5535);
nor U6963 (N_6963,N_5734,N_5286);
xnor U6964 (N_6964,N_5634,N_5956);
and U6965 (N_6965,N_5351,N_5087);
or U6966 (N_6966,N_5080,N_5629);
or U6967 (N_6967,N_5400,N_5497);
nor U6968 (N_6968,N_5987,N_5253);
nor U6969 (N_6969,N_5693,N_5123);
nor U6970 (N_6970,N_5613,N_5051);
xnor U6971 (N_6971,N_5910,N_5361);
or U6972 (N_6972,N_5858,N_5173);
xor U6973 (N_6973,N_5525,N_5334);
and U6974 (N_6974,N_5754,N_5775);
xor U6975 (N_6975,N_5351,N_5885);
nor U6976 (N_6976,N_5181,N_5521);
and U6977 (N_6977,N_5031,N_5964);
xor U6978 (N_6978,N_5547,N_5523);
nand U6979 (N_6979,N_5024,N_5396);
and U6980 (N_6980,N_5711,N_5766);
nand U6981 (N_6981,N_5051,N_5872);
and U6982 (N_6982,N_5376,N_5303);
nor U6983 (N_6983,N_5031,N_5938);
nand U6984 (N_6984,N_5316,N_5849);
nand U6985 (N_6985,N_5180,N_5589);
nor U6986 (N_6986,N_5412,N_5080);
nor U6987 (N_6987,N_5992,N_5164);
nand U6988 (N_6988,N_5266,N_5453);
and U6989 (N_6989,N_5658,N_5912);
xnor U6990 (N_6990,N_5479,N_5009);
nor U6991 (N_6991,N_5827,N_5343);
nor U6992 (N_6992,N_5344,N_5229);
nor U6993 (N_6993,N_5885,N_5224);
xor U6994 (N_6994,N_5595,N_5408);
or U6995 (N_6995,N_5525,N_5624);
nor U6996 (N_6996,N_5275,N_5637);
or U6997 (N_6997,N_5509,N_5948);
or U6998 (N_6998,N_5895,N_5978);
nor U6999 (N_6999,N_5997,N_5696);
and U7000 (N_7000,N_6058,N_6624);
nor U7001 (N_7001,N_6890,N_6255);
or U7002 (N_7002,N_6053,N_6463);
or U7003 (N_7003,N_6158,N_6082);
and U7004 (N_7004,N_6171,N_6126);
nor U7005 (N_7005,N_6691,N_6070);
nand U7006 (N_7006,N_6910,N_6172);
and U7007 (N_7007,N_6054,N_6840);
nand U7008 (N_7008,N_6297,N_6800);
xnor U7009 (N_7009,N_6168,N_6263);
xor U7010 (N_7010,N_6433,N_6372);
nand U7011 (N_7011,N_6667,N_6440);
or U7012 (N_7012,N_6909,N_6674);
nand U7013 (N_7013,N_6446,N_6280);
or U7014 (N_7014,N_6431,N_6285);
or U7015 (N_7015,N_6543,N_6309);
xor U7016 (N_7016,N_6369,N_6805);
nor U7017 (N_7017,N_6312,N_6872);
and U7018 (N_7018,N_6874,N_6103);
nand U7019 (N_7019,N_6899,N_6948);
xnor U7020 (N_7020,N_6024,N_6959);
nor U7021 (N_7021,N_6453,N_6019);
nand U7022 (N_7022,N_6476,N_6825);
xor U7023 (N_7023,N_6596,N_6497);
and U7024 (N_7024,N_6188,N_6376);
or U7025 (N_7025,N_6511,N_6278);
nand U7026 (N_7026,N_6966,N_6668);
xnor U7027 (N_7027,N_6830,N_6467);
xor U7028 (N_7028,N_6695,N_6965);
nor U7029 (N_7029,N_6514,N_6034);
xor U7030 (N_7030,N_6710,N_6223);
or U7031 (N_7031,N_6562,N_6527);
nand U7032 (N_7032,N_6300,N_6773);
xor U7033 (N_7033,N_6381,N_6995);
nand U7034 (N_7034,N_6443,N_6986);
nand U7035 (N_7035,N_6794,N_6895);
nand U7036 (N_7036,N_6603,N_6635);
nand U7037 (N_7037,N_6020,N_6326);
nand U7038 (N_7038,N_6235,N_6139);
or U7039 (N_7039,N_6161,N_6795);
nand U7040 (N_7040,N_6666,N_6083);
nor U7041 (N_7041,N_6332,N_6927);
nand U7042 (N_7042,N_6484,N_6799);
xnor U7043 (N_7043,N_6682,N_6980);
and U7044 (N_7044,N_6209,N_6379);
and U7045 (N_7045,N_6673,N_6227);
xnor U7046 (N_7046,N_6025,N_6652);
and U7047 (N_7047,N_6022,N_6958);
nand U7048 (N_7048,N_6204,N_6625);
and U7049 (N_7049,N_6566,N_6869);
xor U7050 (N_7050,N_6307,N_6190);
nor U7051 (N_7051,N_6665,N_6640);
nand U7052 (N_7052,N_6498,N_6677);
nand U7053 (N_7053,N_6616,N_6599);
and U7054 (N_7054,N_6117,N_6404);
and U7055 (N_7055,N_6137,N_6628);
or U7056 (N_7056,N_6915,N_6554);
nor U7057 (N_7057,N_6351,N_6120);
nor U7058 (N_7058,N_6397,N_6522);
nor U7059 (N_7059,N_6047,N_6760);
and U7060 (N_7060,N_6837,N_6253);
nor U7061 (N_7061,N_6279,N_6038);
nor U7062 (N_7062,N_6324,N_6731);
nor U7063 (N_7063,N_6122,N_6565);
nand U7064 (N_7064,N_6935,N_6924);
and U7065 (N_7065,N_6182,N_6454);
nor U7066 (N_7066,N_6239,N_6343);
or U7067 (N_7067,N_6193,N_6219);
nor U7068 (N_7068,N_6357,N_6481);
xor U7069 (N_7069,N_6807,N_6848);
nand U7070 (N_7070,N_6631,N_6932);
and U7071 (N_7071,N_6203,N_6246);
nand U7072 (N_7072,N_6000,N_6093);
nand U7073 (N_7073,N_6743,N_6437);
nor U7074 (N_7074,N_6736,N_6987);
xor U7075 (N_7075,N_6953,N_6189);
nor U7076 (N_7076,N_6764,N_6345);
nor U7077 (N_7077,N_6509,N_6270);
nor U7078 (N_7078,N_6237,N_6733);
and U7079 (N_7079,N_6809,N_6561);
and U7080 (N_7080,N_6559,N_6536);
nor U7081 (N_7081,N_6937,N_6205);
or U7082 (N_7082,N_6808,N_6289);
and U7083 (N_7083,N_6875,N_6845);
nor U7084 (N_7084,N_6755,N_6770);
and U7085 (N_7085,N_6500,N_6778);
xor U7086 (N_7086,N_6929,N_6810);
nor U7087 (N_7087,N_6546,N_6468);
nor U7088 (N_7088,N_6806,N_6521);
and U7089 (N_7089,N_6336,N_6542);
nor U7090 (N_7090,N_6916,N_6298);
nand U7091 (N_7091,N_6950,N_6415);
nor U7092 (N_7092,N_6659,N_6422);
and U7093 (N_7093,N_6634,N_6734);
nor U7094 (N_7094,N_6206,N_6076);
and U7095 (N_7095,N_6842,N_6132);
or U7096 (N_7096,N_6225,N_6811);
nor U7097 (N_7097,N_6064,N_6905);
xnor U7098 (N_7098,N_6207,N_6482);
and U7099 (N_7099,N_6823,N_6085);
and U7100 (N_7100,N_6316,N_6871);
and U7101 (N_7101,N_6098,N_6580);
xor U7102 (N_7102,N_6181,N_6311);
xor U7103 (N_7103,N_6793,N_6470);
nand U7104 (N_7104,N_6942,N_6886);
nand U7105 (N_7105,N_6897,N_6119);
nand U7106 (N_7106,N_6060,N_6664);
and U7107 (N_7107,N_6418,N_6244);
nor U7108 (N_7108,N_6475,N_6903);
nand U7109 (N_7109,N_6232,N_6409);
xnor U7110 (N_7110,N_6850,N_6902);
xnor U7111 (N_7111,N_6310,N_6104);
nor U7112 (N_7112,N_6146,N_6501);
nand U7113 (N_7113,N_6096,N_6164);
xor U7114 (N_7114,N_6593,N_6940);
xnor U7115 (N_7115,N_6982,N_6478);
or U7116 (N_7116,N_6140,N_6424);
nand U7117 (N_7117,N_6035,N_6354);
xor U7118 (N_7118,N_6169,N_6604);
xnor U7119 (N_7119,N_6928,N_6321);
xnor U7120 (N_7120,N_6314,N_6320);
nand U7121 (N_7121,N_6291,N_6273);
or U7122 (N_7122,N_6988,N_6271);
or U7123 (N_7123,N_6425,N_6390);
and U7124 (N_7124,N_6030,N_6220);
nand U7125 (N_7125,N_6647,N_6436);
xnor U7126 (N_7126,N_6907,N_6637);
nor U7127 (N_7127,N_6577,N_6663);
xor U7128 (N_7128,N_6486,N_6605);
or U7129 (N_7129,N_6394,N_6781);
nand U7130 (N_7130,N_6349,N_6589);
xor U7131 (N_7131,N_6547,N_6683);
nor U7132 (N_7132,N_6973,N_6346);
nor U7133 (N_7133,N_6044,N_6095);
nor U7134 (N_7134,N_6788,N_6059);
or U7135 (N_7135,N_6639,N_6857);
nand U7136 (N_7136,N_6487,N_6553);
and U7137 (N_7137,N_6308,N_6633);
nor U7138 (N_7138,N_6914,N_6541);
or U7139 (N_7139,N_6532,N_6090);
nor U7140 (N_7140,N_6116,N_6445);
nand U7141 (N_7141,N_6588,N_6177);
or U7142 (N_7142,N_6943,N_6365);
and U7143 (N_7143,N_6991,N_6693);
xor U7144 (N_7144,N_6643,N_6451);
xnor U7145 (N_7145,N_6334,N_6448);
nor U7146 (N_7146,N_6826,N_6075);
nand U7147 (N_7147,N_6912,N_6295);
nor U7148 (N_7148,N_6626,N_6597);
nor U7149 (N_7149,N_6983,N_6386);
and U7150 (N_7150,N_6769,N_6864);
or U7151 (N_7151,N_6758,N_6387);
nor U7152 (N_7152,N_6974,N_6776);
xor U7153 (N_7153,N_6411,N_6560);
and U7154 (N_7154,N_6496,N_6504);
nand U7155 (N_7155,N_6175,N_6893);
nor U7156 (N_7156,N_6153,N_6911);
and U7157 (N_7157,N_6266,N_6109);
or U7158 (N_7158,N_6144,N_6569);
or U7159 (N_7159,N_6131,N_6821);
nor U7160 (N_7160,N_6520,N_6630);
xnor U7161 (N_7161,N_6579,N_6018);
nand U7162 (N_7162,N_6032,N_6015);
xor U7163 (N_7163,N_6621,N_6105);
nor U7164 (N_7164,N_6787,N_6785);
or U7165 (N_7165,N_6563,N_6094);
and U7166 (N_7166,N_6452,N_6272);
or U7167 (N_7167,N_6614,N_6471);
or U7168 (N_7168,N_6660,N_6548);
or U7169 (N_7169,N_6523,N_6342);
nor U7170 (N_7170,N_6202,N_6011);
nor U7171 (N_7171,N_6277,N_6613);
nor U7172 (N_7172,N_6762,N_6551);
xnor U7173 (N_7173,N_6601,N_6706);
xor U7174 (N_7174,N_6642,N_6761);
nor U7175 (N_7175,N_6327,N_6858);
nand U7176 (N_7176,N_6378,N_6707);
and U7177 (N_7177,N_6748,N_6264);
nand U7178 (N_7178,N_6023,N_6495);
or U7179 (N_7179,N_6191,N_6675);
xnor U7180 (N_7180,N_6002,N_6347);
or U7181 (N_7181,N_6931,N_6441);
or U7182 (N_7182,N_6843,N_6281);
or U7183 (N_7183,N_6071,N_6184);
and U7184 (N_7184,N_6222,N_6240);
nand U7185 (N_7185,N_6210,N_6534);
xor U7186 (N_7186,N_6333,N_6533);
nor U7187 (N_7187,N_6215,N_6564);
xnor U7188 (N_7188,N_6641,N_6057);
xnor U7189 (N_7189,N_6335,N_6697);
and U7190 (N_7190,N_6091,N_6317);
and U7191 (N_7191,N_6692,N_6724);
nor U7192 (N_7192,N_6701,N_6473);
and U7193 (N_7193,N_6539,N_6792);
nor U7194 (N_7194,N_6696,N_6700);
and U7195 (N_7195,N_6363,N_6382);
or U7196 (N_7196,N_6961,N_6143);
xor U7197 (N_7197,N_6508,N_6557);
or U7198 (N_7198,N_6427,N_6728);
nand U7199 (N_7199,N_6714,N_6617);
xnor U7200 (N_7200,N_6051,N_6818);
nand U7201 (N_7201,N_6079,N_6938);
nand U7202 (N_7202,N_6881,N_6261);
and U7203 (N_7203,N_6155,N_6145);
nand U7204 (N_7204,N_6717,N_6407);
nand U7205 (N_7205,N_6978,N_6199);
nor U7206 (N_7206,N_6483,N_6888);
and U7207 (N_7207,N_6949,N_6322);
xnor U7208 (N_7208,N_6669,N_6535);
xor U7209 (N_7209,N_6477,N_6056);
xnor U7210 (N_7210,N_6195,N_6926);
and U7211 (N_7211,N_6672,N_6102);
xor U7212 (N_7212,N_6080,N_6606);
nor U7213 (N_7213,N_6439,N_6055);
and U7214 (N_7214,N_6824,N_6414);
or U7215 (N_7215,N_6331,N_6917);
and U7216 (N_7216,N_6494,N_6774);
nand U7217 (N_7217,N_6160,N_6248);
nand U7218 (N_7218,N_6353,N_6444);
or U7219 (N_7219,N_6513,N_6646);
or U7220 (N_7220,N_6670,N_6398);
or U7221 (N_7221,N_6505,N_6124);
nand U7222 (N_7222,N_6197,N_6703);
nor U7223 (N_7223,N_6726,N_6485);
xnor U7224 (N_7224,N_6866,N_6396);
nor U7225 (N_7225,N_6282,N_6662);
xnor U7226 (N_7226,N_6061,N_6999);
nand U7227 (N_7227,N_6048,N_6434);
and U7228 (N_7228,N_6885,N_6627);
or U7229 (N_7229,N_6720,N_6163);
or U7230 (N_7230,N_6592,N_6571);
and U7231 (N_7231,N_6016,N_6127);
nand U7232 (N_7232,N_6010,N_6419);
and U7233 (N_7233,N_6923,N_6620);
nor U7234 (N_7234,N_6360,N_6152);
or U7235 (N_7235,N_6786,N_6249);
or U7236 (N_7236,N_6366,N_6148);
and U7237 (N_7237,N_6582,N_6293);
nor U7238 (N_7238,N_6167,N_6087);
nand U7239 (N_7239,N_6361,N_6258);
nand U7240 (N_7240,N_6540,N_6012);
nor U7241 (N_7241,N_6106,N_6884);
nand U7242 (N_7242,N_6891,N_6086);
or U7243 (N_7243,N_6224,N_6142);
nand U7244 (N_7244,N_6068,N_6458);
and U7245 (N_7245,N_6233,N_6330);
and U7246 (N_7246,N_6783,N_6066);
nor U7247 (N_7247,N_6490,N_6186);
or U7248 (N_7248,N_6151,N_6713);
xnor U7249 (N_7249,N_6254,N_6684);
nand U7250 (N_7250,N_6969,N_6503);
nand U7251 (N_7251,N_6855,N_6108);
and U7252 (N_7252,N_6268,N_6591);
nor U7253 (N_7253,N_6529,N_6492);
and U7254 (N_7254,N_6516,N_6515);
or U7255 (N_7255,N_6413,N_6876);
xnor U7256 (N_7256,N_6636,N_6939);
nor U7257 (N_7257,N_6827,N_6882);
nor U7258 (N_7258,N_6650,N_6043);
nand U7259 (N_7259,N_6901,N_6801);
and U7260 (N_7260,N_6623,N_6288);
nand U7261 (N_7261,N_6198,N_6416);
nor U7262 (N_7262,N_6814,N_6506);
xnor U7263 (N_7263,N_6975,N_6052);
nand U7264 (N_7264,N_6303,N_6962);
nand U7265 (N_7265,N_6350,N_6704);
nand U7266 (N_7266,N_6461,N_6925);
or U7267 (N_7267,N_6649,N_6319);
nand U7268 (N_7268,N_6590,N_6567);
or U7269 (N_7269,N_6934,N_6073);
xnor U7270 (N_7270,N_6782,N_6658);
and U7271 (N_7271,N_6651,N_6970);
or U7272 (N_7272,N_6951,N_6392);
nand U7273 (N_7273,N_6746,N_6595);
xnor U7274 (N_7274,N_6517,N_6469);
nor U7275 (N_7275,N_6654,N_6399);
nor U7276 (N_7276,N_6180,N_6375);
nand U7277 (N_7277,N_6896,N_6723);
nor U7278 (N_7278,N_6290,N_6065);
or U7279 (N_7279,N_6196,N_6750);
and U7280 (N_7280,N_6526,N_6299);
or U7281 (N_7281,N_6072,N_6819);
xnor U7282 (N_7282,N_6853,N_6747);
nand U7283 (N_7283,N_6287,N_6217);
nand U7284 (N_7284,N_6989,N_6584);
nand U7285 (N_7285,N_6687,N_6829);
nand U7286 (N_7286,N_6370,N_6135);
and U7287 (N_7287,N_6883,N_6681);
or U7288 (N_7288,N_6302,N_6138);
and U7289 (N_7289,N_6766,N_6771);
xnor U7290 (N_7290,N_6420,N_6385);
xnor U7291 (N_7291,N_6763,N_6545);
or U7292 (N_7292,N_6552,N_6432);
nor U7293 (N_7293,N_6525,N_6252);
or U7294 (N_7294,N_6721,N_6136);
xor U7295 (N_7295,N_6472,N_6737);
nor U7296 (N_7296,N_6154,N_6046);
or U7297 (N_7297,N_6955,N_6100);
nor U7298 (N_7298,N_6039,N_6115);
nand U7299 (N_7299,N_6676,N_6849);
xor U7300 (N_7300,N_6130,N_6873);
or U7301 (N_7301,N_6229,N_6185);
or U7302 (N_7302,N_6259,N_6084);
and U7303 (N_7303,N_6007,N_6388);
nand U7304 (N_7304,N_6241,N_6945);
nand U7305 (N_7305,N_6709,N_6967);
or U7306 (N_7306,N_6306,N_6981);
nand U7307 (N_7307,N_6870,N_6518);
nor U7308 (N_7308,N_6679,N_6412);
and U7309 (N_7309,N_6752,N_6341);
nor U7310 (N_7310,N_6573,N_6097);
nand U7311 (N_7311,N_6921,N_6493);
nor U7312 (N_7312,N_6113,N_6648);
or U7313 (N_7313,N_6765,N_6170);
and U7314 (N_7314,N_6618,N_6732);
nand U7315 (N_7315,N_6339,N_6657);
nor U7316 (N_7316,N_6067,N_6549);
or U7317 (N_7317,N_6157,N_6256);
xnor U7318 (N_7318,N_6006,N_6519);
nand U7319 (N_7319,N_6283,N_6708);
nor U7320 (N_7320,N_6570,N_6753);
or U7321 (N_7321,N_6844,N_6653);
xor U7322 (N_7322,N_6898,N_6026);
xor U7323 (N_7323,N_6479,N_6622);
and U7324 (N_7324,N_6041,N_6125);
or U7325 (N_7325,N_6996,N_6262);
nand U7326 (N_7326,N_6005,N_6612);
nor U7327 (N_7327,N_6238,N_6491);
xor U7328 (N_7328,N_6465,N_6685);
or U7329 (N_7329,N_6833,N_6619);
or U7330 (N_7330,N_6865,N_6429);
xnor U7331 (N_7331,N_6174,N_6680);
or U7332 (N_7332,N_6460,N_6338);
and U7333 (N_7333,N_6009,N_6919);
nor U7334 (N_7334,N_6021,N_6822);
nor U7335 (N_7335,N_6946,N_6393);
nand U7336 (N_7336,N_6031,N_6798);
nor U7337 (N_7337,N_6194,N_6538);
and U7338 (N_7338,N_6267,N_6964);
or U7339 (N_7339,N_6231,N_6323);
or U7340 (N_7340,N_6014,N_6367);
or U7341 (N_7341,N_6908,N_6147);
nor U7342 (N_7342,N_6337,N_6128);
xor U7343 (N_7343,N_6852,N_6954);
or U7344 (N_7344,N_6963,N_6230);
or U7345 (N_7345,N_6629,N_6383);
nand U7346 (N_7346,N_6192,N_6305);
nand U7347 (N_7347,N_6112,N_6364);
nand U7348 (N_7348,N_6586,N_6742);
nor U7349 (N_7349,N_6555,N_6608);
and U7350 (N_7350,N_6466,N_6744);
nor U7351 (N_7351,N_6269,N_6201);
xor U7352 (N_7352,N_6159,N_6480);
xnor U7353 (N_7353,N_6401,N_6208);
nor U7354 (N_7354,N_6123,N_6069);
xnor U7355 (N_7355,N_6426,N_6528);
nand U7356 (N_7356,N_6089,N_6489);
nand U7357 (N_7357,N_6502,N_6328);
nor U7358 (N_7358,N_6245,N_6729);
nor U7359 (N_7359,N_6718,N_6110);
nand U7360 (N_7360,N_6550,N_6179);
xor U7361 (N_7361,N_6325,N_6671);
and U7362 (N_7362,N_6598,N_6968);
and U7363 (N_7363,N_6216,N_6141);
xor U7364 (N_7364,N_6049,N_6947);
nor U7365 (N_7365,N_6212,N_6234);
nand U7366 (N_7366,N_6735,N_6013);
nand U7367 (N_7367,N_6402,N_6027);
nand U7368 (N_7368,N_6329,N_6063);
and U7369 (N_7369,N_6941,N_6111);
nand U7370 (N_7370,N_6741,N_6854);
and U7371 (N_7371,N_6730,N_6400);
nand U7372 (N_7372,N_6183,N_6003);
xor U7373 (N_7373,N_6275,N_6558);
xnor U7374 (N_7374,N_6906,N_6040);
nand U7375 (N_7375,N_6847,N_6775);
and U7376 (N_7376,N_6133,N_6879);
or U7377 (N_7377,N_6575,N_6587);
nor U7378 (N_7378,N_6294,N_6754);
xnor U7379 (N_7379,N_6772,N_6149);
and U7380 (N_7380,N_6880,N_6979);
nor U7381 (N_7381,N_6831,N_6757);
and U7382 (N_7382,N_6738,N_6512);
nor U7383 (N_7383,N_6530,N_6352);
nand U7384 (N_7384,N_6221,N_6428);
nor U7385 (N_7385,N_6609,N_6074);
and U7386 (N_7386,N_6644,N_6162);
xnor U7387 (N_7387,N_6645,N_6745);
nand U7388 (N_7388,N_6286,N_6362);
nor U7389 (N_7389,N_6581,N_6944);
nand U7390 (N_7390,N_6856,N_6537);
xnor U7391 (N_7391,N_6992,N_6292);
xor U7392 (N_7392,N_6990,N_6768);
or U7393 (N_7393,N_6572,N_6779);
or U7394 (N_7394,N_6610,N_6789);
nor U7395 (N_7395,N_6711,N_6456);
and U7396 (N_7396,N_6442,N_6611);
nor U7397 (N_7397,N_6211,N_6062);
nor U7398 (N_7398,N_6348,N_6462);
nand U7399 (N_7399,N_6832,N_6839);
nand U7400 (N_7400,N_6423,N_6894);
and U7401 (N_7401,N_6088,N_6449);
nand U7402 (N_7402,N_6862,N_6421);
nor U7403 (N_7403,N_6340,N_6791);
and U7404 (N_7404,N_6384,N_6200);
xor U7405 (N_7405,N_6813,N_6033);
or U7406 (N_7406,N_6214,N_6816);
or U7407 (N_7407,N_6594,N_6218);
nand U7408 (N_7408,N_6820,N_6403);
xnor U7409 (N_7409,N_6719,N_6815);
or U7410 (N_7410,N_6344,N_6368);
nor U7411 (N_7411,N_6702,N_6276);
and U7412 (N_7412,N_6078,N_6892);
and U7413 (N_7413,N_6510,N_6930);
nand U7414 (N_7414,N_6107,N_6994);
xor U7415 (N_7415,N_6001,N_6689);
and U7416 (N_7416,N_6887,N_6661);
or U7417 (N_7417,N_6242,N_6756);
and U7418 (N_7418,N_6716,N_6568);
nand U7419 (N_7419,N_6972,N_6050);
or U7420 (N_7420,N_6796,N_6722);
nand U7421 (N_7421,N_6574,N_6835);
nor U7422 (N_7422,N_6638,N_6712);
nand U7423 (N_7423,N_6984,N_6812);
and U7424 (N_7424,N_6851,N_6410);
nand U7425 (N_7425,N_6993,N_6900);
nand U7426 (N_7426,N_6318,N_6828);
nor U7427 (N_7427,N_6867,N_6150);
xnor U7428 (N_7428,N_6173,N_6607);
and U7429 (N_7429,N_6099,N_6817);
nor U7430 (N_7430,N_6655,N_6129);
and U7431 (N_7431,N_6391,N_6698);
and U7432 (N_7432,N_6077,N_6725);
or U7433 (N_7433,N_6877,N_6101);
nor U7434 (N_7434,N_6260,N_6028);
xnor U7435 (N_7435,N_6956,N_6373);
xnor U7436 (N_7436,N_6374,N_6092);
and U7437 (N_7437,N_6438,N_6699);
nand U7438 (N_7438,N_6355,N_6187);
xnor U7439 (N_7439,N_6834,N_6380);
xor U7440 (N_7440,N_6838,N_6045);
and U7441 (N_7441,N_6081,N_6455);
xor U7442 (N_7442,N_6957,N_6134);
xor U7443 (N_7443,N_6166,N_6767);
xnor U7444 (N_7444,N_6008,N_6802);
and U7445 (N_7445,N_6952,N_6985);
nor U7446 (N_7446,N_6913,N_6447);
and U7447 (N_7447,N_6274,N_6417);
or U7448 (N_7448,N_6377,N_6578);
and U7449 (N_7449,N_6406,N_6474);
and U7450 (N_7450,N_6790,N_6236);
xnor U7451 (N_7451,N_6156,N_6836);
or U7452 (N_7452,N_6459,N_6408);
and U7453 (N_7453,N_6861,N_6017);
nor U7454 (N_7454,N_6960,N_6740);
nand U7455 (N_7455,N_6600,N_6936);
and U7456 (N_7456,N_6977,N_6265);
or U7457 (N_7457,N_6846,N_6036);
and U7458 (N_7458,N_6922,N_6751);
nor U7459 (N_7459,N_6859,N_6457);
nor U7460 (N_7460,N_6803,N_6920);
xor U7461 (N_7461,N_6739,N_6284);
or U7462 (N_7462,N_6583,N_6405);
xor U7463 (N_7463,N_6841,N_6114);
or U7464 (N_7464,N_6296,N_6998);
or U7465 (N_7465,N_6759,N_6933);
nor U7466 (N_7466,N_6615,N_6576);
and U7467 (N_7467,N_6435,N_6694);
or U7468 (N_7468,N_6727,N_6356);
and U7469 (N_7469,N_6804,N_6971);
nand U7470 (N_7470,N_6690,N_6688);
xnor U7471 (N_7471,N_6868,N_6524);
nand U7472 (N_7472,N_6585,N_6450);
nor U7473 (N_7473,N_6780,N_6632);
nor U7474 (N_7474,N_6257,N_6247);
nand U7475 (N_7475,N_6004,N_6371);
xor U7476 (N_7476,N_6556,N_6749);
and U7477 (N_7477,N_6889,N_6042);
nand U7478 (N_7478,N_6250,N_6029);
or U7479 (N_7479,N_6784,N_6395);
nor U7480 (N_7480,N_6656,N_6226);
and U7481 (N_7481,N_6464,N_6304);
nor U7482 (N_7482,N_6678,N_6213);
nor U7483 (N_7483,N_6507,N_6118);
or U7484 (N_7484,N_6165,N_6997);
xnor U7485 (N_7485,N_6178,N_6037);
or U7486 (N_7486,N_6176,N_6878);
nor U7487 (N_7487,N_6430,N_6863);
nand U7488 (N_7488,N_6531,N_6715);
or U7489 (N_7489,N_6904,N_6301);
nand U7490 (N_7490,N_6686,N_6797);
nor U7491 (N_7491,N_6976,N_6243);
and U7492 (N_7492,N_6251,N_6389);
and U7493 (N_7493,N_6121,N_6228);
xnor U7494 (N_7494,N_6315,N_6358);
nand U7495 (N_7495,N_6705,N_6602);
nand U7496 (N_7496,N_6918,N_6313);
xor U7497 (N_7497,N_6860,N_6359);
xnor U7498 (N_7498,N_6777,N_6488);
and U7499 (N_7499,N_6499,N_6544);
and U7500 (N_7500,N_6306,N_6230);
xor U7501 (N_7501,N_6912,N_6653);
nand U7502 (N_7502,N_6460,N_6985);
xnor U7503 (N_7503,N_6830,N_6863);
nor U7504 (N_7504,N_6665,N_6060);
xnor U7505 (N_7505,N_6435,N_6426);
xnor U7506 (N_7506,N_6209,N_6350);
nand U7507 (N_7507,N_6131,N_6246);
and U7508 (N_7508,N_6422,N_6691);
xnor U7509 (N_7509,N_6742,N_6877);
nand U7510 (N_7510,N_6842,N_6908);
and U7511 (N_7511,N_6373,N_6669);
and U7512 (N_7512,N_6589,N_6781);
xnor U7513 (N_7513,N_6207,N_6677);
or U7514 (N_7514,N_6686,N_6679);
and U7515 (N_7515,N_6274,N_6884);
xnor U7516 (N_7516,N_6347,N_6849);
nor U7517 (N_7517,N_6432,N_6059);
nand U7518 (N_7518,N_6565,N_6780);
xor U7519 (N_7519,N_6586,N_6384);
xnor U7520 (N_7520,N_6652,N_6636);
or U7521 (N_7521,N_6648,N_6200);
and U7522 (N_7522,N_6655,N_6929);
and U7523 (N_7523,N_6002,N_6130);
and U7524 (N_7524,N_6997,N_6833);
nor U7525 (N_7525,N_6952,N_6688);
and U7526 (N_7526,N_6768,N_6184);
xnor U7527 (N_7527,N_6241,N_6378);
or U7528 (N_7528,N_6337,N_6962);
or U7529 (N_7529,N_6366,N_6816);
or U7530 (N_7530,N_6956,N_6288);
xnor U7531 (N_7531,N_6754,N_6050);
nor U7532 (N_7532,N_6292,N_6197);
or U7533 (N_7533,N_6762,N_6851);
or U7534 (N_7534,N_6448,N_6386);
and U7535 (N_7535,N_6439,N_6436);
nand U7536 (N_7536,N_6673,N_6472);
xor U7537 (N_7537,N_6791,N_6917);
xor U7538 (N_7538,N_6063,N_6966);
and U7539 (N_7539,N_6326,N_6225);
and U7540 (N_7540,N_6767,N_6667);
nand U7541 (N_7541,N_6362,N_6224);
xnor U7542 (N_7542,N_6393,N_6652);
nor U7543 (N_7543,N_6409,N_6173);
and U7544 (N_7544,N_6489,N_6235);
xnor U7545 (N_7545,N_6783,N_6836);
xor U7546 (N_7546,N_6284,N_6777);
or U7547 (N_7547,N_6896,N_6145);
nand U7548 (N_7548,N_6007,N_6041);
nor U7549 (N_7549,N_6582,N_6422);
nor U7550 (N_7550,N_6536,N_6611);
nor U7551 (N_7551,N_6320,N_6897);
nand U7552 (N_7552,N_6431,N_6922);
xor U7553 (N_7553,N_6152,N_6079);
nor U7554 (N_7554,N_6264,N_6343);
nand U7555 (N_7555,N_6816,N_6985);
nor U7556 (N_7556,N_6508,N_6330);
nand U7557 (N_7557,N_6548,N_6288);
nor U7558 (N_7558,N_6378,N_6555);
nor U7559 (N_7559,N_6224,N_6585);
nand U7560 (N_7560,N_6418,N_6024);
or U7561 (N_7561,N_6049,N_6995);
nor U7562 (N_7562,N_6599,N_6706);
nor U7563 (N_7563,N_6253,N_6284);
nand U7564 (N_7564,N_6566,N_6577);
and U7565 (N_7565,N_6804,N_6039);
and U7566 (N_7566,N_6609,N_6944);
nor U7567 (N_7567,N_6835,N_6818);
nand U7568 (N_7568,N_6998,N_6103);
nand U7569 (N_7569,N_6106,N_6589);
nor U7570 (N_7570,N_6855,N_6134);
or U7571 (N_7571,N_6947,N_6060);
and U7572 (N_7572,N_6119,N_6475);
and U7573 (N_7573,N_6553,N_6390);
nand U7574 (N_7574,N_6181,N_6335);
or U7575 (N_7575,N_6189,N_6820);
xnor U7576 (N_7576,N_6892,N_6484);
xnor U7577 (N_7577,N_6650,N_6898);
and U7578 (N_7578,N_6965,N_6030);
xnor U7579 (N_7579,N_6255,N_6083);
or U7580 (N_7580,N_6427,N_6086);
nor U7581 (N_7581,N_6632,N_6608);
xor U7582 (N_7582,N_6607,N_6678);
nand U7583 (N_7583,N_6959,N_6508);
nor U7584 (N_7584,N_6384,N_6086);
xnor U7585 (N_7585,N_6472,N_6118);
and U7586 (N_7586,N_6564,N_6707);
nand U7587 (N_7587,N_6819,N_6692);
or U7588 (N_7588,N_6842,N_6593);
or U7589 (N_7589,N_6785,N_6479);
xor U7590 (N_7590,N_6472,N_6583);
and U7591 (N_7591,N_6415,N_6145);
and U7592 (N_7592,N_6618,N_6185);
and U7593 (N_7593,N_6685,N_6734);
nand U7594 (N_7594,N_6280,N_6398);
and U7595 (N_7595,N_6682,N_6874);
nor U7596 (N_7596,N_6857,N_6444);
nand U7597 (N_7597,N_6648,N_6286);
xnor U7598 (N_7598,N_6396,N_6353);
nor U7599 (N_7599,N_6921,N_6666);
and U7600 (N_7600,N_6952,N_6517);
nor U7601 (N_7601,N_6426,N_6967);
nor U7602 (N_7602,N_6912,N_6951);
nor U7603 (N_7603,N_6756,N_6722);
nor U7604 (N_7604,N_6689,N_6819);
xnor U7605 (N_7605,N_6977,N_6711);
nand U7606 (N_7606,N_6074,N_6924);
and U7607 (N_7607,N_6906,N_6701);
or U7608 (N_7608,N_6289,N_6655);
nand U7609 (N_7609,N_6935,N_6098);
and U7610 (N_7610,N_6749,N_6807);
or U7611 (N_7611,N_6484,N_6589);
nand U7612 (N_7612,N_6846,N_6207);
xor U7613 (N_7613,N_6900,N_6868);
xor U7614 (N_7614,N_6270,N_6635);
nand U7615 (N_7615,N_6819,N_6605);
xor U7616 (N_7616,N_6348,N_6756);
xnor U7617 (N_7617,N_6373,N_6905);
or U7618 (N_7618,N_6831,N_6747);
or U7619 (N_7619,N_6868,N_6709);
nor U7620 (N_7620,N_6197,N_6753);
nor U7621 (N_7621,N_6541,N_6154);
xnor U7622 (N_7622,N_6294,N_6846);
or U7623 (N_7623,N_6020,N_6314);
and U7624 (N_7624,N_6312,N_6896);
nor U7625 (N_7625,N_6766,N_6586);
nor U7626 (N_7626,N_6697,N_6319);
or U7627 (N_7627,N_6920,N_6400);
or U7628 (N_7628,N_6202,N_6713);
xnor U7629 (N_7629,N_6307,N_6673);
nand U7630 (N_7630,N_6455,N_6116);
and U7631 (N_7631,N_6919,N_6824);
nand U7632 (N_7632,N_6119,N_6220);
nand U7633 (N_7633,N_6806,N_6781);
nor U7634 (N_7634,N_6399,N_6524);
or U7635 (N_7635,N_6154,N_6459);
nand U7636 (N_7636,N_6779,N_6450);
xor U7637 (N_7637,N_6984,N_6014);
nand U7638 (N_7638,N_6674,N_6508);
and U7639 (N_7639,N_6526,N_6518);
nor U7640 (N_7640,N_6296,N_6923);
and U7641 (N_7641,N_6249,N_6920);
nor U7642 (N_7642,N_6075,N_6918);
nor U7643 (N_7643,N_6040,N_6165);
nand U7644 (N_7644,N_6861,N_6050);
xnor U7645 (N_7645,N_6958,N_6792);
nand U7646 (N_7646,N_6157,N_6025);
and U7647 (N_7647,N_6484,N_6950);
nor U7648 (N_7648,N_6888,N_6142);
nand U7649 (N_7649,N_6758,N_6551);
and U7650 (N_7650,N_6231,N_6273);
nor U7651 (N_7651,N_6053,N_6486);
or U7652 (N_7652,N_6620,N_6312);
nor U7653 (N_7653,N_6565,N_6160);
or U7654 (N_7654,N_6467,N_6680);
nor U7655 (N_7655,N_6245,N_6009);
xor U7656 (N_7656,N_6013,N_6714);
nor U7657 (N_7657,N_6669,N_6901);
nand U7658 (N_7658,N_6470,N_6862);
nand U7659 (N_7659,N_6930,N_6717);
nor U7660 (N_7660,N_6031,N_6948);
nor U7661 (N_7661,N_6557,N_6883);
or U7662 (N_7662,N_6682,N_6365);
and U7663 (N_7663,N_6231,N_6275);
xnor U7664 (N_7664,N_6196,N_6489);
and U7665 (N_7665,N_6632,N_6404);
and U7666 (N_7666,N_6111,N_6021);
or U7667 (N_7667,N_6257,N_6292);
and U7668 (N_7668,N_6910,N_6604);
or U7669 (N_7669,N_6741,N_6590);
and U7670 (N_7670,N_6261,N_6636);
or U7671 (N_7671,N_6167,N_6923);
nor U7672 (N_7672,N_6984,N_6849);
nand U7673 (N_7673,N_6040,N_6096);
or U7674 (N_7674,N_6588,N_6661);
or U7675 (N_7675,N_6210,N_6614);
xor U7676 (N_7676,N_6574,N_6410);
nand U7677 (N_7677,N_6347,N_6692);
and U7678 (N_7678,N_6182,N_6622);
nand U7679 (N_7679,N_6728,N_6322);
or U7680 (N_7680,N_6957,N_6174);
xor U7681 (N_7681,N_6248,N_6780);
or U7682 (N_7682,N_6084,N_6758);
xor U7683 (N_7683,N_6000,N_6096);
xor U7684 (N_7684,N_6553,N_6070);
nor U7685 (N_7685,N_6835,N_6290);
xor U7686 (N_7686,N_6762,N_6880);
nor U7687 (N_7687,N_6914,N_6016);
or U7688 (N_7688,N_6579,N_6388);
and U7689 (N_7689,N_6387,N_6229);
xnor U7690 (N_7690,N_6638,N_6835);
or U7691 (N_7691,N_6781,N_6631);
or U7692 (N_7692,N_6966,N_6590);
nand U7693 (N_7693,N_6298,N_6279);
nor U7694 (N_7694,N_6123,N_6788);
xor U7695 (N_7695,N_6294,N_6991);
and U7696 (N_7696,N_6026,N_6133);
nand U7697 (N_7697,N_6086,N_6807);
and U7698 (N_7698,N_6192,N_6377);
or U7699 (N_7699,N_6962,N_6150);
nor U7700 (N_7700,N_6500,N_6719);
or U7701 (N_7701,N_6524,N_6222);
or U7702 (N_7702,N_6822,N_6263);
and U7703 (N_7703,N_6723,N_6988);
xnor U7704 (N_7704,N_6341,N_6982);
nor U7705 (N_7705,N_6384,N_6293);
nor U7706 (N_7706,N_6158,N_6369);
or U7707 (N_7707,N_6842,N_6001);
or U7708 (N_7708,N_6882,N_6417);
xnor U7709 (N_7709,N_6366,N_6184);
and U7710 (N_7710,N_6234,N_6073);
nand U7711 (N_7711,N_6878,N_6383);
xor U7712 (N_7712,N_6078,N_6951);
or U7713 (N_7713,N_6518,N_6030);
nand U7714 (N_7714,N_6793,N_6959);
nor U7715 (N_7715,N_6879,N_6890);
and U7716 (N_7716,N_6183,N_6489);
nor U7717 (N_7717,N_6814,N_6053);
nand U7718 (N_7718,N_6217,N_6541);
and U7719 (N_7719,N_6389,N_6844);
or U7720 (N_7720,N_6814,N_6148);
or U7721 (N_7721,N_6362,N_6688);
nand U7722 (N_7722,N_6326,N_6713);
nor U7723 (N_7723,N_6938,N_6093);
and U7724 (N_7724,N_6786,N_6044);
nor U7725 (N_7725,N_6365,N_6356);
and U7726 (N_7726,N_6493,N_6001);
nor U7727 (N_7727,N_6835,N_6365);
nand U7728 (N_7728,N_6894,N_6118);
and U7729 (N_7729,N_6150,N_6536);
or U7730 (N_7730,N_6864,N_6878);
nand U7731 (N_7731,N_6679,N_6242);
nor U7732 (N_7732,N_6598,N_6977);
nor U7733 (N_7733,N_6170,N_6703);
xor U7734 (N_7734,N_6515,N_6340);
nand U7735 (N_7735,N_6328,N_6759);
nor U7736 (N_7736,N_6631,N_6864);
and U7737 (N_7737,N_6824,N_6790);
xnor U7738 (N_7738,N_6503,N_6632);
xor U7739 (N_7739,N_6906,N_6570);
and U7740 (N_7740,N_6945,N_6941);
nand U7741 (N_7741,N_6436,N_6381);
or U7742 (N_7742,N_6833,N_6984);
nor U7743 (N_7743,N_6200,N_6718);
nand U7744 (N_7744,N_6622,N_6231);
xor U7745 (N_7745,N_6133,N_6842);
nand U7746 (N_7746,N_6228,N_6111);
and U7747 (N_7747,N_6917,N_6377);
or U7748 (N_7748,N_6018,N_6930);
xor U7749 (N_7749,N_6640,N_6094);
and U7750 (N_7750,N_6136,N_6515);
nand U7751 (N_7751,N_6170,N_6821);
or U7752 (N_7752,N_6394,N_6445);
or U7753 (N_7753,N_6647,N_6796);
or U7754 (N_7754,N_6265,N_6803);
and U7755 (N_7755,N_6731,N_6070);
or U7756 (N_7756,N_6801,N_6198);
or U7757 (N_7757,N_6523,N_6874);
nor U7758 (N_7758,N_6763,N_6092);
and U7759 (N_7759,N_6345,N_6581);
xnor U7760 (N_7760,N_6801,N_6460);
or U7761 (N_7761,N_6081,N_6830);
nor U7762 (N_7762,N_6411,N_6001);
or U7763 (N_7763,N_6455,N_6339);
nor U7764 (N_7764,N_6179,N_6582);
or U7765 (N_7765,N_6359,N_6888);
or U7766 (N_7766,N_6631,N_6192);
nor U7767 (N_7767,N_6041,N_6652);
xnor U7768 (N_7768,N_6778,N_6128);
and U7769 (N_7769,N_6332,N_6279);
nand U7770 (N_7770,N_6130,N_6936);
or U7771 (N_7771,N_6243,N_6479);
nor U7772 (N_7772,N_6177,N_6233);
nand U7773 (N_7773,N_6359,N_6981);
nor U7774 (N_7774,N_6745,N_6885);
nand U7775 (N_7775,N_6782,N_6899);
nand U7776 (N_7776,N_6220,N_6028);
nand U7777 (N_7777,N_6784,N_6417);
nand U7778 (N_7778,N_6315,N_6423);
xor U7779 (N_7779,N_6314,N_6493);
nand U7780 (N_7780,N_6070,N_6613);
or U7781 (N_7781,N_6366,N_6349);
nand U7782 (N_7782,N_6468,N_6665);
or U7783 (N_7783,N_6394,N_6355);
nand U7784 (N_7784,N_6564,N_6177);
or U7785 (N_7785,N_6199,N_6729);
or U7786 (N_7786,N_6114,N_6780);
or U7787 (N_7787,N_6189,N_6375);
or U7788 (N_7788,N_6191,N_6111);
nand U7789 (N_7789,N_6244,N_6293);
and U7790 (N_7790,N_6246,N_6708);
xnor U7791 (N_7791,N_6189,N_6601);
xnor U7792 (N_7792,N_6782,N_6679);
and U7793 (N_7793,N_6979,N_6631);
and U7794 (N_7794,N_6337,N_6130);
or U7795 (N_7795,N_6109,N_6816);
nor U7796 (N_7796,N_6905,N_6599);
nor U7797 (N_7797,N_6592,N_6329);
and U7798 (N_7798,N_6606,N_6000);
nand U7799 (N_7799,N_6635,N_6634);
nor U7800 (N_7800,N_6323,N_6736);
xnor U7801 (N_7801,N_6725,N_6460);
and U7802 (N_7802,N_6685,N_6182);
and U7803 (N_7803,N_6028,N_6179);
or U7804 (N_7804,N_6380,N_6479);
nor U7805 (N_7805,N_6038,N_6161);
nor U7806 (N_7806,N_6922,N_6397);
nand U7807 (N_7807,N_6600,N_6756);
nor U7808 (N_7808,N_6665,N_6682);
or U7809 (N_7809,N_6493,N_6908);
nand U7810 (N_7810,N_6192,N_6113);
nor U7811 (N_7811,N_6645,N_6699);
nor U7812 (N_7812,N_6635,N_6364);
and U7813 (N_7813,N_6022,N_6433);
nor U7814 (N_7814,N_6333,N_6900);
nand U7815 (N_7815,N_6613,N_6581);
xor U7816 (N_7816,N_6164,N_6149);
nor U7817 (N_7817,N_6533,N_6497);
or U7818 (N_7818,N_6611,N_6143);
nor U7819 (N_7819,N_6596,N_6246);
xnor U7820 (N_7820,N_6146,N_6921);
xor U7821 (N_7821,N_6946,N_6632);
nand U7822 (N_7822,N_6911,N_6991);
nor U7823 (N_7823,N_6002,N_6047);
nand U7824 (N_7824,N_6920,N_6898);
or U7825 (N_7825,N_6151,N_6307);
xnor U7826 (N_7826,N_6181,N_6291);
or U7827 (N_7827,N_6839,N_6118);
nand U7828 (N_7828,N_6868,N_6119);
xnor U7829 (N_7829,N_6700,N_6537);
and U7830 (N_7830,N_6577,N_6036);
and U7831 (N_7831,N_6059,N_6458);
nor U7832 (N_7832,N_6229,N_6330);
and U7833 (N_7833,N_6604,N_6262);
or U7834 (N_7834,N_6236,N_6891);
nand U7835 (N_7835,N_6850,N_6990);
nor U7836 (N_7836,N_6830,N_6274);
nand U7837 (N_7837,N_6309,N_6674);
nor U7838 (N_7838,N_6652,N_6614);
and U7839 (N_7839,N_6957,N_6301);
nand U7840 (N_7840,N_6082,N_6162);
nor U7841 (N_7841,N_6867,N_6523);
xnor U7842 (N_7842,N_6649,N_6222);
xor U7843 (N_7843,N_6680,N_6140);
nand U7844 (N_7844,N_6478,N_6782);
and U7845 (N_7845,N_6207,N_6928);
or U7846 (N_7846,N_6796,N_6599);
xor U7847 (N_7847,N_6768,N_6629);
nor U7848 (N_7848,N_6145,N_6296);
xor U7849 (N_7849,N_6804,N_6645);
nand U7850 (N_7850,N_6500,N_6818);
xnor U7851 (N_7851,N_6594,N_6392);
or U7852 (N_7852,N_6926,N_6318);
nand U7853 (N_7853,N_6458,N_6484);
xor U7854 (N_7854,N_6678,N_6039);
xor U7855 (N_7855,N_6126,N_6794);
or U7856 (N_7856,N_6373,N_6578);
xor U7857 (N_7857,N_6248,N_6325);
and U7858 (N_7858,N_6052,N_6776);
xor U7859 (N_7859,N_6490,N_6967);
and U7860 (N_7860,N_6913,N_6550);
nand U7861 (N_7861,N_6309,N_6362);
and U7862 (N_7862,N_6973,N_6171);
nand U7863 (N_7863,N_6797,N_6043);
nand U7864 (N_7864,N_6768,N_6836);
xnor U7865 (N_7865,N_6198,N_6942);
nor U7866 (N_7866,N_6553,N_6207);
xor U7867 (N_7867,N_6431,N_6963);
nor U7868 (N_7868,N_6025,N_6533);
and U7869 (N_7869,N_6925,N_6051);
nor U7870 (N_7870,N_6079,N_6329);
nand U7871 (N_7871,N_6385,N_6880);
and U7872 (N_7872,N_6972,N_6390);
nand U7873 (N_7873,N_6402,N_6238);
xnor U7874 (N_7874,N_6756,N_6919);
nand U7875 (N_7875,N_6080,N_6574);
nor U7876 (N_7876,N_6325,N_6699);
nor U7877 (N_7877,N_6687,N_6256);
nor U7878 (N_7878,N_6722,N_6508);
and U7879 (N_7879,N_6998,N_6927);
nand U7880 (N_7880,N_6999,N_6429);
nor U7881 (N_7881,N_6900,N_6577);
xnor U7882 (N_7882,N_6485,N_6192);
and U7883 (N_7883,N_6123,N_6839);
or U7884 (N_7884,N_6492,N_6322);
nand U7885 (N_7885,N_6359,N_6566);
xor U7886 (N_7886,N_6514,N_6919);
or U7887 (N_7887,N_6363,N_6754);
xor U7888 (N_7888,N_6066,N_6462);
nand U7889 (N_7889,N_6484,N_6474);
or U7890 (N_7890,N_6065,N_6035);
nor U7891 (N_7891,N_6382,N_6587);
nor U7892 (N_7892,N_6723,N_6377);
nor U7893 (N_7893,N_6537,N_6840);
nand U7894 (N_7894,N_6595,N_6483);
nor U7895 (N_7895,N_6741,N_6754);
xnor U7896 (N_7896,N_6532,N_6242);
or U7897 (N_7897,N_6296,N_6818);
nand U7898 (N_7898,N_6259,N_6615);
xor U7899 (N_7899,N_6914,N_6695);
or U7900 (N_7900,N_6883,N_6105);
xnor U7901 (N_7901,N_6646,N_6737);
xnor U7902 (N_7902,N_6391,N_6488);
or U7903 (N_7903,N_6477,N_6821);
nand U7904 (N_7904,N_6525,N_6661);
nand U7905 (N_7905,N_6870,N_6166);
or U7906 (N_7906,N_6085,N_6945);
nand U7907 (N_7907,N_6644,N_6278);
nand U7908 (N_7908,N_6783,N_6916);
xor U7909 (N_7909,N_6070,N_6972);
nor U7910 (N_7910,N_6351,N_6526);
nand U7911 (N_7911,N_6481,N_6254);
nand U7912 (N_7912,N_6128,N_6985);
xor U7913 (N_7913,N_6071,N_6414);
nand U7914 (N_7914,N_6380,N_6720);
nor U7915 (N_7915,N_6217,N_6521);
nand U7916 (N_7916,N_6223,N_6808);
and U7917 (N_7917,N_6541,N_6605);
nand U7918 (N_7918,N_6946,N_6778);
xor U7919 (N_7919,N_6671,N_6042);
and U7920 (N_7920,N_6085,N_6943);
nor U7921 (N_7921,N_6926,N_6035);
or U7922 (N_7922,N_6042,N_6378);
nor U7923 (N_7923,N_6695,N_6355);
and U7924 (N_7924,N_6343,N_6245);
and U7925 (N_7925,N_6632,N_6680);
nor U7926 (N_7926,N_6353,N_6467);
and U7927 (N_7927,N_6129,N_6977);
nand U7928 (N_7928,N_6756,N_6605);
nand U7929 (N_7929,N_6954,N_6040);
or U7930 (N_7930,N_6162,N_6269);
nand U7931 (N_7931,N_6728,N_6995);
nor U7932 (N_7932,N_6763,N_6713);
xnor U7933 (N_7933,N_6871,N_6122);
or U7934 (N_7934,N_6995,N_6481);
nand U7935 (N_7935,N_6213,N_6560);
nor U7936 (N_7936,N_6890,N_6028);
nor U7937 (N_7937,N_6753,N_6675);
or U7938 (N_7938,N_6203,N_6397);
nand U7939 (N_7939,N_6304,N_6747);
nand U7940 (N_7940,N_6727,N_6937);
nand U7941 (N_7941,N_6569,N_6365);
xnor U7942 (N_7942,N_6974,N_6624);
nor U7943 (N_7943,N_6169,N_6222);
or U7944 (N_7944,N_6737,N_6005);
and U7945 (N_7945,N_6830,N_6373);
nand U7946 (N_7946,N_6748,N_6761);
or U7947 (N_7947,N_6735,N_6707);
or U7948 (N_7948,N_6883,N_6183);
or U7949 (N_7949,N_6762,N_6720);
and U7950 (N_7950,N_6163,N_6614);
nand U7951 (N_7951,N_6297,N_6793);
nor U7952 (N_7952,N_6498,N_6434);
nor U7953 (N_7953,N_6983,N_6399);
nand U7954 (N_7954,N_6099,N_6848);
or U7955 (N_7955,N_6322,N_6698);
and U7956 (N_7956,N_6817,N_6877);
xnor U7957 (N_7957,N_6579,N_6706);
xor U7958 (N_7958,N_6285,N_6974);
nor U7959 (N_7959,N_6882,N_6903);
nor U7960 (N_7960,N_6511,N_6675);
nand U7961 (N_7961,N_6287,N_6007);
and U7962 (N_7962,N_6421,N_6949);
nor U7963 (N_7963,N_6700,N_6262);
nor U7964 (N_7964,N_6230,N_6239);
nor U7965 (N_7965,N_6207,N_6222);
and U7966 (N_7966,N_6691,N_6372);
or U7967 (N_7967,N_6995,N_6157);
nor U7968 (N_7968,N_6962,N_6609);
nand U7969 (N_7969,N_6835,N_6115);
and U7970 (N_7970,N_6782,N_6100);
xor U7971 (N_7971,N_6800,N_6214);
or U7972 (N_7972,N_6046,N_6081);
or U7973 (N_7973,N_6046,N_6857);
or U7974 (N_7974,N_6745,N_6727);
or U7975 (N_7975,N_6892,N_6984);
xnor U7976 (N_7976,N_6028,N_6555);
or U7977 (N_7977,N_6875,N_6208);
nand U7978 (N_7978,N_6648,N_6687);
nand U7979 (N_7979,N_6914,N_6998);
nor U7980 (N_7980,N_6271,N_6447);
and U7981 (N_7981,N_6762,N_6532);
and U7982 (N_7982,N_6175,N_6131);
nor U7983 (N_7983,N_6032,N_6374);
xor U7984 (N_7984,N_6008,N_6482);
and U7985 (N_7985,N_6311,N_6699);
nor U7986 (N_7986,N_6483,N_6488);
and U7987 (N_7987,N_6077,N_6046);
nand U7988 (N_7988,N_6706,N_6360);
and U7989 (N_7989,N_6280,N_6680);
and U7990 (N_7990,N_6243,N_6724);
nand U7991 (N_7991,N_6631,N_6646);
nor U7992 (N_7992,N_6212,N_6089);
xor U7993 (N_7993,N_6760,N_6765);
or U7994 (N_7994,N_6274,N_6948);
or U7995 (N_7995,N_6990,N_6755);
or U7996 (N_7996,N_6732,N_6237);
xor U7997 (N_7997,N_6538,N_6392);
xor U7998 (N_7998,N_6161,N_6559);
nor U7999 (N_7999,N_6005,N_6894);
or U8000 (N_8000,N_7281,N_7527);
and U8001 (N_8001,N_7242,N_7896);
and U8002 (N_8002,N_7118,N_7171);
nor U8003 (N_8003,N_7056,N_7279);
or U8004 (N_8004,N_7961,N_7410);
or U8005 (N_8005,N_7563,N_7862);
and U8006 (N_8006,N_7052,N_7869);
xnor U8007 (N_8007,N_7111,N_7224);
nor U8008 (N_8008,N_7227,N_7036);
xor U8009 (N_8009,N_7349,N_7311);
nand U8010 (N_8010,N_7409,N_7807);
nor U8011 (N_8011,N_7871,N_7496);
xnor U8012 (N_8012,N_7136,N_7123);
xnor U8013 (N_8013,N_7680,N_7492);
nor U8014 (N_8014,N_7288,N_7423);
xnor U8015 (N_8015,N_7889,N_7587);
and U8016 (N_8016,N_7940,N_7247);
nand U8017 (N_8017,N_7248,N_7933);
or U8018 (N_8018,N_7882,N_7829);
or U8019 (N_8019,N_7449,N_7385);
and U8020 (N_8020,N_7086,N_7342);
nor U8021 (N_8021,N_7365,N_7571);
and U8022 (N_8022,N_7361,N_7647);
or U8023 (N_8023,N_7939,N_7820);
nand U8024 (N_8024,N_7812,N_7946);
nor U8025 (N_8025,N_7074,N_7969);
and U8026 (N_8026,N_7468,N_7355);
or U8027 (N_8027,N_7285,N_7107);
xor U8028 (N_8028,N_7033,N_7740);
nand U8029 (N_8029,N_7474,N_7816);
nand U8030 (N_8030,N_7175,N_7044);
and U8031 (N_8031,N_7536,N_7794);
nand U8032 (N_8032,N_7234,N_7637);
nor U8033 (N_8033,N_7935,N_7394);
xor U8034 (N_8034,N_7280,N_7225);
and U8035 (N_8035,N_7879,N_7324);
nor U8036 (N_8036,N_7913,N_7800);
and U8037 (N_8037,N_7199,N_7110);
xor U8038 (N_8038,N_7024,N_7244);
nor U8039 (N_8039,N_7340,N_7153);
or U8040 (N_8040,N_7992,N_7648);
nand U8041 (N_8041,N_7343,N_7263);
nand U8042 (N_8042,N_7608,N_7284);
or U8043 (N_8043,N_7641,N_7152);
and U8044 (N_8044,N_7019,N_7654);
nor U8045 (N_8045,N_7835,N_7254);
nor U8046 (N_8046,N_7016,N_7352);
and U8047 (N_8047,N_7389,N_7728);
nand U8048 (N_8048,N_7575,N_7318);
nor U8049 (N_8049,N_7709,N_7834);
nand U8050 (N_8050,N_7738,N_7660);
or U8051 (N_8051,N_7774,N_7450);
nand U8052 (N_8052,N_7336,N_7158);
nor U8053 (N_8053,N_7549,N_7895);
and U8054 (N_8054,N_7170,N_7290);
nand U8055 (N_8055,N_7307,N_7704);
nor U8056 (N_8056,N_7934,N_7184);
xor U8057 (N_8057,N_7106,N_7327);
or U8058 (N_8058,N_7228,N_7950);
nor U8059 (N_8059,N_7076,N_7168);
and U8060 (N_8060,N_7770,N_7194);
and U8061 (N_8061,N_7141,N_7497);
nand U8062 (N_8062,N_7192,N_7500);
nand U8063 (N_8063,N_7518,N_7880);
xor U8064 (N_8064,N_7154,N_7005);
nor U8065 (N_8065,N_7018,N_7268);
xor U8066 (N_8066,N_7951,N_7588);
or U8067 (N_8067,N_7428,N_7900);
xnor U8068 (N_8068,N_7229,N_7029);
and U8069 (N_8069,N_7870,N_7581);
xnor U8070 (N_8070,N_7661,N_7269);
xnor U8071 (N_8071,N_7475,N_7180);
or U8072 (N_8072,N_7677,N_7217);
nand U8073 (N_8073,N_7705,N_7273);
and U8074 (N_8074,N_7972,N_7923);
xnor U8075 (N_8075,N_7981,N_7758);
or U8076 (N_8076,N_7090,N_7424);
or U8077 (N_8077,N_7299,N_7725);
and U8078 (N_8078,N_7069,N_7119);
and U8079 (N_8079,N_7208,N_7730);
nand U8080 (N_8080,N_7039,N_7464);
nand U8081 (N_8081,N_7767,N_7821);
or U8082 (N_8082,N_7792,N_7121);
and U8083 (N_8083,N_7407,N_7116);
xor U8084 (N_8084,N_7542,N_7043);
nand U8085 (N_8085,N_7852,N_7746);
or U8086 (N_8086,N_7393,N_7957);
xnor U8087 (N_8087,N_7734,N_7973);
nor U8088 (N_8088,N_7965,N_7133);
xor U8089 (N_8089,N_7521,N_7867);
nor U8090 (N_8090,N_7253,N_7543);
xnor U8091 (N_8091,N_7235,N_7621);
and U8092 (N_8092,N_7126,N_7260);
nor U8093 (N_8093,N_7038,N_7264);
xor U8094 (N_8094,N_7833,N_7777);
or U8095 (N_8095,N_7541,N_7522);
nand U8096 (N_8096,N_7566,N_7860);
nand U8097 (N_8097,N_7538,N_7723);
and U8098 (N_8098,N_7875,N_7696);
xnor U8099 (N_8099,N_7837,N_7788);
nor U8100 (N_8100,N_7432,N_7130);
xor U8101 (N_8101,N_7367,N_7544);
or U8102 (N_8102,N_7612,N_7613);
nor U8103 (N_8103,N_7380,N_7586);
nor U8104 (N_8104,N_7062,N_7427);
or U8105 (N_8105,N_7089,N_7552);
or U8106 (N_8106,N_7178,N_7291);
and U8107 (N_8107,N_7551,N_7784);
and U8108 (N_8108,N_7562,N_7966);
or U8109 (N_8109,N_7855,N_7422);
xor U8110 (N_8110,N_7490,N_7331);
nor U8111 (N_8111,N_7322,N_7341);
and U8112 (N_8112,N_7021,N_7907);
and U8113 (N_8113,N_7716,N_7143);
nand U8114 (N_8114,N_7173,N_7467);
or U8115 (N_8115,N_7849,N_7809);
nand U8116 (N_8116,N_7582,N_7053);
nor U8117 (N_8117,N_7321,N_7674);
nor U8118 (N_8118,N_7292,N_7081);
nor U8119 (N_8119,N_7145,N_7459);
and U8120 (N_8120,N_7615,N_7499);
or U8121 (N_8121,N_7131,N_7553);
or U8122 (N_8122,N_7993,N_7437);
or U8123 (N_8123,N_7640,N_7616);
nor U8124 (N_8124,N_7537,N_7569);
nor U8125 (N_8125,N_7902,N_7667);
and U8126 (N_8126,N_7020,N_7446);
nor U8127 (N_8127,N_7762,N_7669);
nand U8128 (N_8128,N_7839,N_7822);
nand U8129 (N_8129,N_7572,N_7642);
or U8130 (N_8130,N_7323,N_7914);
and U8131 (N_8131,N_7397,N_7597);
xnor U8132 (N_8132,N_7238,N_7398);
nand U8133 (N_8133,N_7547,N_7160);
nand U8134 (N_8134,N_7692,N_7930);
nor U8135 (N_8135,N_7007,N_7887);
xor U8136 (N_8136,N_7294,N_7431);
and U8137 (N_8137,N_7611,N_7811);
xnor U8138 (N_8138,N_7023,N_7626);
or U8139 (N_8139,N_7334,N_7656);
xnor U8140 (N_8140,N_7333,N_7994);
nor U8141 (N_8141,N_7986,N_7694);
or U8142 (N_8142,N_7798,N_7655);
or U8143 (N_8143,N_7519,N_7658);
xnor U8144 (N_8144,N_7713,N_7167);
nor U8145 (N_8145,N_7147,N_7139);
or U8146 (N_8146,N_7604,N_7146);
and U8147 (N_8147,N_7594,N_7975);
xnor U8148 (N_8148,N_7861,N_7371);
nand U8149 (N_8149,N_7463,N_7698);
xnor U8150 (N_8150,N_7980,N_7006);
and U8151 (N_8151,N_7348,N_7164);
and U8152 (N_8152,N_7003,N_7243);
xnor U8153 (N_8153,N_7873,N_7046);
nor U8154 (N_8154,N_7634,N_7567);
xnor U8155 (N_8155,N_7737,N_7109);
or U8156 (N_8156,N_7561,N_7216);
nor U8157 (N_8157,N_7351,N_7138);
nand U8158 (N_8158,N_7583,N_7874);
xor U8159 (N_8159,N_7967,N_7577);
nor U8160 (N_8160,N_7927,N_7771);
xnor U8161 (N_8161,N_7293,N_7652);
nand U8162 (N_8162,N_7451,N_7898);
and U8163 (N_8163,N_7245,N_7987);
nor U8164 (N_8164,N_7638,N_7205);
and U8165 (N_8165,N_7721,N_7908);
or U8166 (N_8166,N_7193,N_7388);
or U8167 (N_8167,N_7974,N_7050);
nor U8168 (N_8168,N_7712,N_7511);
or U8169 (N_8169,N_7761,N_7357);
nor U8170 (N_8170,N_7752,N_7347);
xnor U8171 (N_8171,N_7607,N_7922);
xnor U8172 (N_8172,N_7941,N_7990);
xnor U8173 (N_8173,N_7962,N_7828);
or U8174 (N_8174,N_7404,N_7296);
xnor U8175 (N_8175,N_7488,N_7295);
nand U8176 (N_8176,N_7448,N_7883);
or U8177 (N_8177,N_7071,N_7316);
nor U8178 (N_8178,N_7618,N_7134);
or U8179 (N_8179,N_7097,N_7491);
nor U8180 (N_8180,N_7257,N_7457);
and U8181 (N_8181,N_7915,N_7643);
or U8182 (N_8182,N_7010,N_7310);
or U8183 (N_8183,N_7191,N_7379);
xnor U8184 (N_8184,N_7665,N_7486);
nand U8185 (N_8185,N_7048,N_7255);
xnor U8186 (N_8186,N_7970,N_7102);
xor U8187 (N_8187,N_7345,N_7113);
or U8188 (N_8188,N_7445,N_7949);
and U8189 (N_8189,N_7403,N_7354);
nand U8190 (N_8190,N_7516,N_7865);
nor U8191 (N_8191,N_7789,N_7631);
and U8192 (N_8192,N_7818,N_7906);
and U8193 (N_8193,N_7531,N_7937);
and U8194 (N_8194,N_7122,N_7406);
nor U8195 (N_8195,N_7309,N_7719);
or U8196 (N_8196,N_7429,N_7539);
and U8197 (N_8197,N_7091,N_7057);
and U8198 (N_8198,N_7493,N_7142);
and U8199 (N_8199,N_7441,N_7101);
xnor U8200 (N_8200,N_7484,N_7905);
nor U8201 (N_8201,N_7742,N_7578);
or U8202 (N_8202,N_7999,N_7619);
nor U8203 (N_8203,N_7399,N_7769);
nand U8204 (N_8204,N_7751,N_7392);
or U8205 (N_8205,N_7502,N_7979);
nor U8206 (N_8206,N_7465,N_7997);
and U8207 (N_8207,N_7899,N_7787);
or U8208 (N_8208,N_7300,N_7720);
nor U8209 (N_8209,N_7370,N_7884);
or U8210 (N_8210,N_7435,N_7535);
nor U8211 (N_8211,N_7213,N_7120);
nand U8212 (N_8212,N_7666,N_7104);
nand U8213 (N_8213,N_7218,N_7476);
nor U8214 (N_8214,N_7657,N_7162);
or U8215 (N_8215,N_7825,N_7190);
nand U8216 (N_8216,N_7037,N_7159);
and U8217 (N_8217,N_7282,N_7198);
and U8218 (N_8218,N_7453,N_7289);
or U8219 (N_8219,N_7786,N_7550);
or U8220 (N_8220,N_7517,N_7329);
nand U8221 (N_8221,N_7030,N_7344);
and U8222 (N_8222,N_7169,N_7002);
and U8223 (N_8223,N_7649,N_7651);
or U8224 (N_8224,N_7301,N_7795);
and U8225 (N_8225,N_7850,N_7757);
nor U8226 (N_8226,N_7374,N_7181);
nand U8227 (N_8227,N_7554,N_7904);
xnor U8228 (N_8228,N_7505,N_7420);
nor U8229 (N_8229,N_7506,N_7948);
nand U8230 (N_8230,N_7212,N_7080);
and U8231 (N_8231,N_7901,N_7886);
nand U8232 (N_8232,N_7068,N_7186);
xor U8233 (N_8233,N_7826,N_7419);
and U8234 (N_8234,N_7614,N_7697);
xor U8235 (N_8235,N_7646,N_7456);
nand U8236 (N_8236,N_7629,N_7840);
nand U8237 (N_8237,N_7878,N_7000);
xnor U8238 (N_8238,N_7481,N_7338);
xnor U8239 (N_8239,N_7592,N_7004);
xor U8240 (N_8240,N_7768,N_7715);
or U8241 (N_8241,N_7266,N_7312);
and U8242 (N_8242,N_7998,N_7326);
or U8243 (N_8243,N_7765,N_7636);
xor U8244 (N_8244,N_7412,N_7434);
nor U8245 (N_8245,N_7185,N_7617);
xnor U8246 (N_8246,N_7804,N_7405);
and U8247 (N_8247,N_7686,N_7890);
and U8248 (N_8248,N_7054,N_7699);
or U8249 (N_8249,N_7202,N_7396);
nor U8250 (N_8250,N_7909,N_7673);
and U8251 (N_8251,N_7356,N_7797);
or U8252 (N_8252,N_7778,N_7013);
nor U8253 (N_8253,N_7084,N_7042);
xnor U8254 (N_8254,N_7847,N_7953);
and U8255 (N_8255,N_7671,N_7681);
and U8256 (N_8256,N_7859,N_7172);
and U8257 (N_8257,N_7286,N_7596);
nand U8258 (N_8258,N_7524,N_7386);
nand U8259 (N_8259,N_7830,N_7200);
and U8260 (N_8260,N_7960,N_7622);
nand U8261 (N_8261,N_7092,N_7605);
nand U8262 (N_8262,N_7954,N_7876);
xor U8263 (N_8263,N_7026,N_7534);
xnor U8264 (N_8264,N_7440,N_7576);
and U8265 (N_8265,N_7383,N_7087);
or U8266 (N_8266,N_7017,N_7603);
xor U8267 (N_8267,N_7401,N_7853);
xor U8268 (N_8268,N_7472,N_7841);
nor U8269 (N_8269,N_7791,N_7796);
or U8270 (N_8270,N_7144,N_7776);
nand U8271 (N_8271,N_7827,N_7670);
nor U8272 (N_8272,N_7230,N_7805);
or U8273 (N_8273,N_7942,N_7773);
and U8274 (N_8274,N_7358,N_7221);
xnor U8275 (N_8275,N_7595,N_7921);
and U8276 (N_8276,N_7189,N_7801);
nor U8277 (N_8277,N_7645,N_7512);
or U8278 (N_8278,N_7846,N_7894);
nand U8279 (N_8279,N_7529,N_7179);
nand U8280 (N_8280,N_7732,N_7851);
xnor U8281 (N_8281,N_7350,N_7706);
nand U8282 (N_8282,N_7599,N_7701);
or U8283 (N_8283,N_7968,N_7702);
xnor U8284 (N_8284,N_7461,N_7868);
nand U8285 (N_8285,N_7078,N_7215);
and U8286 (N_8286,N_7635,N_7609);
nor U8287 (N_8287,N_7377,N_7843);
nand U8288 (N_8288,N_7944,N_7947);
nand U8289 (N_8289,N_7127,N_7685);
nand U8290 (N_8290,N_7584,N_7240);
and U8291 (N_8291,N_7077,N_7653);
or U8292 (N_8292,N_7772,N_7022);
xnor U8293 (N_8293,N_7753,N_7320);
xor U8294 (N_8294,N_7633,N_7700);
nor U8295 (N_8295,N_7304,N_7443);
and U8296 (N_8296,N_7418,N_7411);
and U8297 (N_8297,N_7362,N_7863);
nand U8298 (N_8298,N_7375,N_7408);
or U8299 (N_8299,N_7856,N_7750);
nor U8300 (N_8300,N_7460,N_7462);
xor U8301 (N_8301,N_7032,N_7688);
nand U8302 (N_8302,N_7112,N_7079);
and U8303 (N_8303,N_7919,N_7689);
nand U8304 (N_8304,N_7366,N_7368);
or U8305 (N_8305,N_7479,N_7684);
and U8306 (N_8306,N_7735,N_7210);
and U8307 (N_8307,N_7378,N_7231);
nor U8308 (N_8308,N_7495,N_7278);
nor U8309 (N_8309,N_7008,N_7739);
xnor U8310 (N_8310,N_7936,N_7478);
or U8311 (N_8311,N_7025,N_7482);
and U8312 (N_8312,N_7070,N_7525);
or U8313 (N_8313,N_7780,N_7831);
and U8314 (N_8314,N_7067,N_7306);
nand U8315 (N_8315,N_7187,N_7748);
nand U8316 (N_8316,N_7731,N_7040);
or U8317 (N_8317,N_7135,N_7838);
nand U8318 (N_8318,N_7978,N_7384);
xnor U8319 (N_8319,N_7845,N_7815);
and U8320 (N_8320,N_7682,N_7832);
or U8321 (N_8321,N_7063,N_7755);
xnor U8322 (N_8322,N_7402,N_7031);
nand U8323 (N_8323,N_7252,N_7964);
and U8324 (N_8324,N_7466,N_7760);
xnor U8325 (N_8325,N_7082,N_7911);
xnor U8326 (N_8326,N_7219,N_7246);
or U8327 (N_8327,N_7319,N_7503);
and U8328 (N_8328,N_7630,N_7687);
nor U8329 (N_8329,N_7854,N_7745);
nand U8330 (N_8330,N_7724,N_7802);
xor U8331 (N_8331,N_7557,N_7664);
xnor U8332 (N_8332,N_7014,N_7675);
xor U8333 (N_8333,N_7672,N_7211);
nand U8334 (N_8334,N_7754,N_7775);
nand U8335 (N_8335,N_7452,N_7659);
nand U8336 (N_8336,N_7444,N_7494);
xnor U8337 (N_8337,N_7372,N_7220);
and U8338 (N_8338,N_7893,N_7925);
nor U8339 (N_8339,N_7241,N_7416);
nor U8340 (N_8340,N_7736,N_7650);
and U8341 (N_8341,N_7259,N_7580);
or U8342 (N_8342,N_7625,N_7382);
nor U8343 (N_8343,N_7691,N_7881);
nand U8344 (N_8344,N_7996,N_7117);
nor U8345 (N_8345,N_7806,N_7223);
nand U8346 (N_8346,N_7163,N_7764);
nor U8347 (N_8347,N_7955,N_7785);
nand U8348 (N_8348,N_7012,N_7783);
nor U8349 (N_8349,N_7564,N_7848);
nor U8350 (N_8350,N_7509,N_7381);
nand U8351 (N_8351,N_7679,N_7100);
xnor U8352 (N_8352,N_7693,N_7498);
nand U8353 (N_8353,N_7639,N_7707);
xnor U8354 (N_8354,N_7001,N_7628);
nand U8355 (N_8355,N_7251,N_7819);
nand U8356 (N_8356,N_7644,N_7556);
or U8357 (N_8357,N_7710,N_7620);
xnor U8358 (N_8358,N_7176,N_7364);
or U8359 (N_8359,N_7376,N_7489);
nand U8360 (N_8360,N_7132,N_7236);
or U8361 (N_8361,N_7150,N_7565);
nand U8362 (N_8362,N_7239,N_7124);
xnor U8363 (N_8363,N_7857,N_7515);
and U8364 (N_8364,N_7533,N_7601);
and U8365 (N_8365,N_7066,N_7781);
nor U8366 (N_8366,N_7958,N_7073);
nor U8367 (N_8367,N_7471,N_7924);
nand U8368 (N_8368,N_7454,N_7574);
nand U8369 (N_8369,N_7415,N_7864);
or U8370 (N_8370,N_7678,N_7174);
nand U8371 (N_8371,N_7346,N_7041);
or U8372 (N_8372,N_7083,N_7442);
and U8373 (N_8373,N_7988,N_7610);
nor U8374 (N_8374,N_7283,N_7866);
nand U8375 (N_8375,N_7233,N_7548);
or U8376 (N_8376,N_7747,N_7714);
nor U8377 (N_8377,N_7058,N_7064);
or U8378 (N_8378,N_7214,N_7526);
or U8379 (N_8379,N_7600,N_7718);
xnor U8380 (N_8380,N_7125,N_7166);
xor U8381 (N_8381,N_7756,N_7177);
xnor U8382 (N_8382,N_7302,N_7267);
or U8383 (N_8383,N_7803,N_7983);
nand U8384 (N_8384,N_7872,N_7417);
or U8385 (N_8385,N_7918,N_7209);
xnor U8386 (N_8386,N_7337,N_7989);
or U8387 (N_8387,N_7182,N_7413);
xor U8388 (N_8388,N_7985,N_7157);
xnor U8389 (N_8389,N_7274,N_7275);
nand U8390 (N_8390,N_7095,N_7059);
or U8391 (N_8391,N_7061,N_7808);
xor U8392 (N_8392,N_7470,N_7888);
nor U8393 (N_8393,N_7155,N_7115);
and U8394 (N_8394,N_7910,N_7624);
nand U8395 (N_8395,N_7045,N_7313);
or U8396 (N_8396,N_7959,N_7128);
and U8397 (N_8397,N_7325,N_7265);
nand U8398 (N_8398,N_7513,N_7779);
nand U8399 (N_8399,N_7991,N_7814);
or U8400 (N_8400,N_7262,N_7314);
xor U8401 (N_8401,N_7929,N_7353);
xnor U8402 (N_8402,N_7717,N_7627);
nor U8403 (N_8403,N_7877,N_7799);
or U8404 (N_8404,N_7733,N_7328);
nor U8405 (N_8405,N_7335,N_7027);
nor U8406 (N_8406,N_7051,N_7477);
xor U8407 (N_8407,N_7072,N_7984);
xor U8408 (N_8408,N_7555,N_7183);
or U8409 (N_8409,N_7270,N_7956);
xnor U8410 (N_8410,N_7226,N_7060);
or U8411 (N_8411,N_7096,N_7824);
nor U8412 (N_8412,N_7237,N_7485);
or U8413 (N_8413,N_7823,N_7891);
nor U8414 (N_8414,N_7703,N_7011);
nor U8415 (N_8415,N_7690,N_7726);
nand U8416 (N_8416,N_7560,N_7129);
or U8417 (N_8417,N_7507,N_7743);
nor U8418 (N_8418,N_7207,N_7222);
nand U8419 (N_8419,N_7501,N_7836);
and U8420 (N_8420,N_7897,N_7593);
nand U8421 (N_8421,N_7813,N_7085);
nor U8422 (N_8422,N_7075,N_7196);
or U8423 (N_8423,N_7579,N_7400);
nand U8424 (N_8424,N_7663,N_7585);
and U8425 (N_8425,N_7149,N_7912);
and U8426 (N_8426,N_7952,N_7945);
and U8427 (N_8427,N_7360,N_7510);
and U8428 (N_8428,N_7928,N_7250);
or U8429 (N_8429,N_7683,N_7623);
and U8430 (N_8430,N_7395,N_7369);
nor U8431 (N_8431,N_7249,N_7793);
and U8432 (N_8432,N_7103,N_7483);
nor U8433 (N_8433,N_7662,N_7790);
and U8434 (N_8434,N_7035,N_7421);
or U8435 (N_8435,N_7436,N_7590);
nor U8436 (N_8436,N_7390,N_7099);
xnor U8437 (N_8437,N_7932,N_7447);
nand U8438 (N_8438,N_7009,N_7744);
or U8439 (N_8439,N_7188,N_7598);
nor U8440 (N_8440,N_7559,N_7148);
or U8441 (N_8441,N_7414,N_7810);
xor U8442 (N_8442,N_7156,N_7916);
nor U8443 (N_8443,N_7602,N_7487);
xor U8444 (N_8444,N_7523,N_7256);
nor U8445 (N_8445,N_7455,N_7098);
nor U8446 (N_8446,N_7976,N_7568);
nand U8447 (N_8447,N_7433,N_7201);
and U8448 (N_8448,N_7094,N_7332);
and U8449 (N_8449,N_7330,N_7151);
or U8450 (N_8450,N_7589,N_7931);
nand U8451 (N_8451,N_7546,N_7232);
nor U8452 (N_8452,N_7926,N_7520);
or U8453 (N_8453,N_7276,N_7308);
xnor U8454 (N_8454,N_7430,N_7920);
nand U8455 (N_8455,N_7844,N_7028);
nand U8456 (N_8456,N_7741,N_7258);
nand U8457 (N_8457,N_7763,N_7858);
nand U8458 (N_8458,N_7817,N_7711);
or U8459 (N_8459,N_7206,N_7903);
nand U8460 (N_8460,N_7047,N_7315);
nand U8461 (N_8461,N_7297,N_7439);
nor U8462 (N_8462,N_7514,N_7426);
xor U8463 (N_8463,N_7277,N_7759);
and U8464 (N_8464,N_7065,N_7458);
or U8465 (N_8465,N_7425,N_7545);
nor U8466 (N_8466,N_7943,N_7885);
and U8467 (N_8467,N_7938,N_7530);
nand U8468 (N_8468,N_7504,N_7303);
nand U8469 (N_8469,N_7298,N_7995);
nand U8470 (N_8470,N_7917,N_7708);
xor U8471 (N_8471,N_7558,N_7971);
nor U8472 (N_8472,N_7093,N_7197);
xnor U8473 (N_8473,N_7676,N_7204);
xor U8474 (N_8474,N_7387,N_7532);
nand U8475 (N_8475,N_7359,N_7049);
nor U8476 (N_8476,N_7034,N_7508);
nand U8477 (N_8477,N_7722,N_7305);
or U8478 (N_8478,N_7261,N_7695);
and U8479 (N_8479,N_7287,N_7161);
or U8480 (N_8480,N_7480,N_7140);
or U8481 (N_8481,N_7573,N_7591);
and U8482 (N_8482,N_7105,N_7271);
or U8483 (N_8483,N_7114,N_7088);
and U8484 (N_8484,N_7339,N_7469);
or U8485 (N_8485,N_7668,N_7842);
xnor U8486 (N_8486,N_7977,N_7363);
nor U8487 (N_8487,N_7963,N_7165);
or U8488 (N_8488,N_7982,N_7137);
and U8489 (N_8489,N_7438,N_7317);
or U8490 (N_8490,N_7373,N_7015);
nor U8491 (N_8491,N_7606,N_7528);
or U8492 (N_8492,N_7782,N_7729);
nor U8493 (N_8493,N_7203,N_7892);
nor U8494 (N_8494,N_7749,N_7570);
or U8495 (N_8495,N_7272,N_7632);
and U8496 (N_8496,N_7391,N_7727);
xor U8497 (N_8497,N_7473,N_7055);
xor U8498 (N_8498,N_7195,N_7108);
xnor U8499 (N_8499,N_7540,N_7766);
nor U8500 (N_8500,N_7815,N_7489);
or U8501 (N_8501,N_7062,N_7354);
and U8502 (N_8502,N_7076,N_7767);
and U8503 (N_8503,N_7466,N_7563);
and U8504 (N_8504,N_7837,N_7552);
and U8505 (N_8505,N_7040,N_7958);
and U8506 (N_8506,N_7163,N_7019);
nand U8507 (N_8507,N_7507,N_7863);
nor U8508 (N_8508,N_7046,N_7273);
and U8509 (N_8509,N_7224,N_7148);
or U8510 (N_8510,N_7951,N_7802);
or U8511 (N_8511,N_7736,N_7824);
xnor U8512 (N_8512,N_7213,N_7330);
xnor U8513 (N_8513,N_7271,N_7807);
xnor U8514 (N_8514,N_7572,N_7821);
or U8515 (N_8515,N_7370,N_7532);
xor U8516 (N_8516,N_7877,N_7000);
nand U8517 (N_8517,N_7442,N_7014);
xnor U8518 (N_8518,N_7676,N_7628);
and U8519 (N_8519,N_7598,N_7543);
and U8520 (N_8520,N_7306,N_7469);
nor U8521 (N_8521,N_7748,N_7357);
nand U8522 (N_8522,N_7517,N_7920);
nor U8523 (N_8523,N_7503,N_7392);
or U8524 (N_8524,N_7074,N_7575);
and U8525 (N_8525,N_7313,N_7558);
nand U8526 (N_8526,N_7203,N_7254);
xnor U8527 (N_8527,N_7740,N_7905);
xnor U8528 (N_8528,N_7106,N_7889);
nor U8529 (N_8529,N_7219,N_7649);
nor U8530 (N_8530,N_7109,N_7114);
or U8531 (N_8531,N_7957,N_7111);
or U8532 (N_8532,N_7670,N_7442);
nor U8533 (N_8533,N_7717,N_7402);
nor U8534 (N_8534,N_7343,N_7813);
nor U8535 (N_8535,N_7637,N_7173);
or U8536 (N_8536,N_7095,N_7088);
or U8537 (N_8537,N_7887,N_7503);
nor U8538 (N_8538,N_7789,N_7765);
nor U8539 (N_8539,N_7778,N_7473);
or U8540 (N_8540,N_7228,N_7648);
nor U8541 (N_8541,N_7964,N_7956);
and U8542 (N_8542,N_7932,N_7349);
xor U8543 (N_8543,N_7139,N_7492);
xor U8544 (N_8544,N_7283,N_7059);
xnor U8545 (N_8545,N_7255,N_7858);
or U8546 (N_8546,N_7485,N_7404);
or U8547 (N_8547,N_7106,N_7282);
or U8548 (N_8548,N_7135,N_7734);
xnor U8549 (N_8549,N_7165,N_7356);
nor U8550 (N_8550,N_7368,N_7291);
nand U8551 (N_8551,N_7049,N_7438);
xnor U8552 (N_8552,N_7287,N_7659);
and U8553 (N_8553,N_7416,N_7854);
or U8554 (N_8554,N_7121,N_7678);
or U8555 (N_8555,N_7363,N_7463);
and U8556 (N_8556,N_7842,N_7196);
nand U8557 (N_8557,N_7406,N_7519);
nand U8558 (N_8558,N_7851,N_7326);
nand U8559 (N_8559,N_7035,N_7754);
xor U8560 (N_8560,N_7787,N_7755);
and U8561 (N_8561,N_7634,N_7485);
and U8562 (N_8562,N_7604,N_7545);
nor U8563 (N_8563,N_7934,N_7699);
nand U8564 (N_8564,N_7970,N_7302);
and U8565 (N_8565,N_7880,N_7904);
and U8566 (N_8566,N_7644,N_7420);
xor U8567 (N_8567,N_7512,N_7555);
xor U8568 (N_8568,N_7033,N_7282);
and U8569 (N_8569,N_7690,N_7308);
nand U8570 (N_8570,N_7976,N_7351);
and U8571 (N_8571,N_7312,N_7679);
and U8572 (N_8572,N_7313,N_7965);
or U8573 (N_8573,N_7989,N_7793);
xor U8574 (N_8574,N_7182,N_7109);
or U8575 (N_8575,N_7811,N_7650);
or U8576 (N_8576,N_7445,N_7966);
xor U8577 (N_8577,N_7664,N_7302);
nor U8578 (N_8578,N_7543,N_7217);
or U8579 (N_8579,N_7001,N_7261);
nand U8580 (N_8580,N_7844,N_7614);
nor U8581 (N_8581,N_7414,N_7410);
or U8582 (N_8582,N_7706,N_7795);
nor U8583 (N_8583,N_7084,N_7539);
or U8584 (N_8584,N_7467,N_7613);
or U8585 (N_8585,N_7430,N_7549);
and U8586 (N_8586,N_7337,N_7224);
nand U8587 (N_8587,N_7701,N_7814);
or U8588 (N_8588,N_7506,N_7322);
nand U8589 (N_8589,N_7557,N_7850);
or U8590 (N_8590,N_7529,N_7246);
nor U8591 (N_8591,N_7842,N_7034);
nor U8592 (N_8592,N_7276,N_7509);
nor U8593 (N_8593,N_7951,N_7258);
nor U8594 (N_8594,N_7716,N_7215);
or U8595 (N_8595,N_7915,N_7333);
nand U8596 (N_8596,N_7154,N_7653);
nand U8597 (N_8597,N_7912,N_7885);
nor U8598 (N_8598,N_7105,N_7895);
nand U8599 (N_8599,N_7417,N_7559);
or U8600 (N_8600,N_7393,N_7423);
nand U8601 (N_8601,N_7886,N_7505);
or U8602 (N_8602,N_7035,N_7923);
nor U8603 (N_8603,N_7249,N_7454);
and U8604 (N_8604,N_7819,N_7610);
nand U8605 (N_8605,N_7029,N_7927);
and U8606 (N_8606,N_7522,N_7883);
nor U8607 (N_8607,N_7979,N_7383);
xnor U8608 (N_8608,N_7732,N_7002);
nor U8609 (N_8609,N_7243,N_7014);
or U8610 (N_8610,N_7550,N_7018);
nor U8611 (N_8611,N_7164,N_7032);
or U8612 (N_8612,N_7126,N_7657);
and U8613 (N_8613,N_7867,N_7810);
or U8614 (N_8614,N_7345,N_7243);
nand U8615 (N_8615,N_7939,N_7585);
or U8616 (N_8616,N_7513,N_7207);
nand U8617 (N_8617,N_7784,N_7168);
nor U8618 (N_8618,N_7516,N_7251);
nand U8619 (N_8619,N_7269,N_7816);
xor U8620 (N_8620,N_7115,N_7017);
or U8621 (N_8621,N_7875,N_7944);
xor U8622 (N_8622,N_7628,N_7250);
nor U8623 (N_8623,N_7514,N_7531);
and U8624 (N_8624,N_7715,N_7730);
nor U8625 (N_8625,N_7035,N_7037);
xor U8626 (N_8626,N_7563,N_7509);
nand U8627 (N_8627,N_7194,N_7589);
or U8628 (N_8628,N_7632,N_7278);
nand U8629 (N_8629,N_7154,N_7495);
nand U8630 (N_8630,N_7679,N_7271);
nand U8631 (N_8631,N_7921,N_7850);
or U8632 (N_8632,N_7825,N_7320);
or U8633 (N_8633,N_7128,N_7019);
nor U8634 (N_8634,N_7498,N_7048);
and U8635 (N_8635,N_7607,N_7481);
or U8636 (N_8636,N_7235,N_7229);
xnor U8637 (N_8637,N_7968,N_7640);
nor U8638 (N_8638,N_7205,N_7702);
or U8639 (N_8639,N_7044,N_7891);
nand U8640 (N_8640,N_7805,N_7673);
nand U8641 (N_8641,N_7266,N_7100);
nor U8642 (N_8642,N_7009,N_7261);
and U8643 (N_8643,N_7657,N_7508);
nand U8644 (N_8644,N_7105,N_7642);
nand U8645 (N_8645,N_7879,N_7409);
xnor U8646 (N_8646,N_7736,N_7450);
or U8647 (N_8647,N_7153,N_7027);
and U8648 (N_8648,N_7659,N_7363);
nand U8649 (N_8649,N_7059,N_7540);
nand U8650 (N_8650,N_7440,N_7860);
and U8651 (N_8651,N_7960,N_7643);
nor U8652 (N_8652,N_7406,N_7612);
or U8653 (N_8653,N_7126,N_7656);
nor U8654 (N_8654,N_7613,N_7174);
xnor U8655 (N_8655,N_7735,N_7060);
or U8656 (N_8656,N_7453,N_7448);
nand U8657 (N_8657,N_7247,N_7385);
or U8658 (N_8658,N_7663,N_7257);
nor U8659 (N_8659,N_7563,N_7828);
xnor U8660 (N_8660,N_7699,N_7616);
xor U8661 (N_8661,N_7847,N_7473);
nor U8662 (N_8662,N_7660,N_7771);
nor U8663 (N_8663,N_7478,N_7506);
or U8664 (N_8664,N_7512,N_7966);
and U8665 (N_8665,N_7325,N_7374);
xnor U8666 (N_8666,N_7831,N_7681);
nor U8667 (N_8667,N_7171,N_7922);
or U8668 (N_8668,N_7576,N_7761);
xnor U8669 (N_8669,N_7540,N_7132);
xor U8670 (N_8670,N_7466,N_7409);
and U8671 (N_8671,N_7025,N_7193);
xnor U8672 (N_8672,N_7392,N_7203);
and U8673 (N_8673,N_7906,N_7705);
nor U8674 (N_8674,N_7192,N_7652);
nand U8675 (N_8675,N_7027,N_7499);
and U8676 (N_8676,N_7553,N_7986);
nand U8677 (N_8677,N_7245,N_7547);
xnor U8678 (N_8678,N_7158,N_7828);
or U8679 (N_8679,N_7788,N_7629);
and U8680 (N_8680,N_7641,N_7694);
or U8681 (N_8681,N_7554,N_7855);
and U8682 (N_8682,N_7640,N_7341);
xor U8683 (N_8683,N_7254,N_7543);
or U8684 (N_8684,N_7117,N_7588);
and U8685 (N_8685,N_7632,N_7446);
and U8686 (N_8686,N_7757,N_7551);
nor U8687 (N_8687,N_7174,N_7790);
or U8688 (N_8688,N_7900,N_7502);
or U8689 (N_8689,N_7445,N_7057);
nor U8690 (N_8690,N_7658,N_7207);
nand U8691 (N_8691,N_7868,N_7371);
nor U8692 (N_8692,N_7984,N_7100);
or U8693 (N_8693,N_7760,N_7379);
and U8694 (N_8694,N_7289,N_7096);
nor U8695 (N_8695,N_7621,N_7690);
or U8696 (N_8696,N_7619,N_7572);
and U8697 (N_8697,N_7130,N_7858);
or U8698 (N_8698,N_7255,N_7038);
nor U8699 (N_8699,N_7390,N_7412);
nand U8700 (N_8700,N_7289,N_7953);
and U8701 (N_8701,N_7328,N_7365);
nand U8702 (N_8702,N_7284,N_7524);
nor U8703 (N_8703,N_7961,N_7500);
nor U8704 (N_8704,N_7775,N_7063);
xor U8705 (N_8705,N_7356,N_7317);
nor U8706 (N_8706,N_7373,N_7028);
nand U8707 (N_8707,N_7485,N_7469);
nand U8708 (N_8708,N_7378,N_7154);
nand U8709 (N_8709,N_7301,N_7609);
xor U8710 (N_8710,N_7294,N_7003);
nand U8711 (N_8711,N_7960,N_7038);
or U8712 (N_8712,N_7211,N_7539);
xnor U8713 (N_8713,N_7700,N_7116);
nor U8714 (N_8714,N_7883,N_7007);
xnor U8715 (N_8715,N_7831,N_7218);
nand U8716 (N_8716,N_7957,N_7212);
nand U8717 (N_8717,N_7567,N_7069);
or U8718 (N_8718,N_7328,N_7307);
and U8719 (N_8719,N_7853,N_7146);
nand U8720 (N_8720,N_7091,N_7349);
or U8721 (N_8721,N_7593,N_7506);
xnor U8722 (N_8722,N_7970,N_7019);
or U8723 (N_8723,N_7752,N_7686);
and U8724 (N_8724,N_7297,N_7323);
nor U8725 (N_8725,N_7885,N_7020);
nand U8726 (N_8726,N_7907,N_7317);
and U8727 (N_8727,N_7269,N_7282);
xnor U8728 (N_8728,N_7747,N_7628);
xnor U8729 (N_8729,N_7932,N_7744);
nor U8730 (N_8730,N_7241,N_7697);
and U8731 (N_8731,N_7058,N_7363);
nand U8732 (N_8732,N_7312,N_7696);
nor U8733 (N_8733,N_7121,N_7978);
nor U8734 (N_8734,N_7182,N_7198);
xor U8735 (N_8735,N_7439,N_7950);
and U8736 (N_8736,N_7776,N_7470);
nand U8737 (N_8737,N_7669,N_7405);
and U8738 (N_8738,N_7629,N_7698);
or U8739 (N_8739,N_7172,N_7147);
or U8740 (N_8740,N_7749,N_7828);
nor U8741 (N_8741,N_7693,N_7502);
nor U8742 (N_8742,N_7949,N_7871);
or U8743 (N_8743,N_7275,N_7692);
or U8744 (N_8744,N_7370,N_7852);
xnor U8745 (N_8745,N_7633,N_7679);
xnor U8746 (N_8746,N_7080,N_7252);
and U8747 (N_8747,N_7714,N_7520);
and U8748 (N_8748,N_7311,N_7864);
or U8749 (N_8749,N_7922,N_7964);
or U8750 (N_8750,N_7994,N_7565);
xor U8751 (N_8751,N_7308,N_7186);
nor U8752 (N_8752,N_7655,N_7957);
nor U8753 (N_8753,N_7650,N_7430);
or U8754 (N_8754,N_7130,N_7544);
nand U8755 (N_8755,N_7486,N_7110);
nor U8756 (N_8756,N_7746,N_7949);
and U8757 (N_8757,N_7593,N_7298);
and U8758 (N_8758,N_7296,N_7133);
or U8759 (N_8759,N_7008,N_7373);
or U8760 (N_8760,N_7889,N_7039);
nand U8761 (N_8761,N_7800,N_7480);
nand U8762 (N_8762,N_7781,N_7222);
nand U8763 (N_8763,N_7910,N_7485);
nand U8764 (N_8764,N_7774,N_7926);
nand U8765 (N_8765,N_7756,N_7861);
and U8766 (N_8766,N_7520,N_7250);
or U8767 (N_8767,N_7428,N_7851);
or U8768 (N_8768,N_7456,N_7930);
and U8769 (N_8769,N_7797,N_7669);
nor U8770 (N_8770,N_7536,N_7326);
and U8771 (N_8771,N_7883,N_7983);
nor U8772 (N_8772,N_7859,N_7707);
xor U8773 (N_8773,N_7642,N_7744);
nand U8774 (N_8774,N_7956,N_7685);
nor U8775 (N_8775,N_7615,N_7368);
and U8776 (N_8776,N_7576,N_7670);
xor U8777 (N_8777,N_7849,N_7928);
and U8778 (N_8778,N_7284,N_7081);
xnor U8779 (N_8779,N_7869,N_7984);
or U8780 (N_8780,N_7681,N_7130);
nand U8781 (N_8781,N_7302,N_7394);
and U8782 (N_8782,N_7231,N_7819);
and U8783 (N_8783,N_7161,N_7586);
and U8784 (N_8784,N_7701,N_7343);
nand U8785 (N_8785,N_7264,N_7291);
xnor U8786 (N_8786,N_7439,N_7723);
nand U8787 (N_8787,N_7579,N_7236);
nand U8788 (N_8788,N_7003,N_7249);
nand U8789 (N_8789,N_7661,N_7889);
nand U8790 (N_8790,N_7834,N_7638);
nand U8791 (N_8791,N_7515,N_7911);
nor U8792 (N_8792,N_7602,N_7955);
and U8793 (N_8793,N_7326,N_7683);
xnor U8794 (N_8794,N_7895,N_7842);
or U8795 (N_8795,N_7699,N_7867);
xor U8796 (N_8796,N_7071,N_7704);
xor U8797 (N_8797,N_7760,N_7727);
xnor U8798 (N_8798,N_7598,N_7876);
or U8799 (N_8799,N_7854,N_7938);
and U8800 (N_8800,N_7087,N_7662);
or U8801 (N_8801,N_7216,N_7609);
nor U8802 (N_8802,N_7221,N_7736);
and U8803 (N_8803,N_7449,N_7725);
and U8804 (N_8804,N_7944,N_7808);
xor U8805 (N_8805,N_7579,N_7452);
nand U8806 (N_8806,N_7201,N_7331);
nor U8807 (N_8807,N_7239,N_7628);
nand U8808 (N_8808,N_7542,N_7299);
nand U8809 (N_8809,N_7208,N_7443);
and U8810 (N_8810,N_7735,N_7832);
or U8811 (N_8811,N_7228,N_7074);
nor U8812 (N_8812,N_7935,N_7145);
xor U8813 (N_8813,N_7588,N_7657);
nor U8814 (N_8814,N_7657,N_7115);
nand U8815 (N_8815,N_7904,N_7507);
nand U8816 (N_8816,N_7399,N_7649);
and U8817 (N_8817,N_7123,N_7535);
xnor U8818 (N_8818,N_7578,N_7472);
or U8819 (N_8819,N_7866,N_7553);
nor U8820 (N_8820,N_7507,N_7177);
nor U8821 (N_8821,N_7890,N_7427);
nand U8822 (N_8822,N_7371,N_7795);
nand U8823 (N_8823,N_7720,N_7345);
nor U8824 (N_8824,N_7606,N_7222);
nor U8825 (N_8825,N_7006,N_7435);
nand U8826 (N_8826,N_7598,N_7407);
nand U8827 (N_8827,N_7815,N_7622);
or U8828 (N_8828,N_7014,N_7614);
nand U8829 (N_8829,N_7574,N_7877);
and U8830 (N_8830,N_7335,N_7986);
xor U8831 (N_8831,N_7745,N_7020);
nand U8832 (N_8832,N_7581,N_7645);
and U8833 (N_8833,N_7726,N_7728);
xor U8834 (N_8834,N_7096,N_7556);
xnor U8835 (N_8835,N_7692,N_7021);
and U8836 (N_8836,N_7991,N_7910);
xnor U8837 (N_8837,N_7205,N_7620);
nand U8838 (N_8838,N_7472,N_7759);
and U8839 (N_8839,N_7608,N_7246);
nor U8840 (N_8840,N_7139,N_7250);
xor U8841 (N_8841,N_7953,N_7254);
nor U8842 (N_8842,N_7886,N_7006);
xnor U8843 (N_8843,N_7924,N_7235);
or U8844 (N_8844,N_7447,N_7779);
xnor U8845 (N_8845,N_7904,N_7627);
xor U8846 (N_8846,N_7151,N_7469);
xnor U8847 (N_8847,N_7671,N_7973);
nand U8848 (N_8848,N_7633,N_7151);
xor U8849 (N_8849,N_7645,N_7519);
or U8850 (N_8850,N_7489,N_7054);
or U8851 (N_8851,N_7975,N_7837);
xor U8852 (N_8852,N_7494,N_7368);
nand U8853 (N_8853,N_7386,N_7392);
and U8854 (N_8854,N_7821,N_7865);
nand U8855 (N_8855,N_7737,N_7431);
nand U8856 (N_8856,N_7166,N_7821);
nand U8857 (N_8857,N_7450,N_7981);
or U8858 (N_8858,N_7947,N_7030);
nand U8859 (N_8859,N_7174,N_7321);
nand U8860 (N_8860,N_7834,N_7517);
xnor U8861 (N_8861,N_7577,N_7886);
or U8862 (N_8862,N_7512,N_7653);
xnor U8863 (N_8863,N_7606,N_7532);
and U8864 (N_8864,N_7097,N_7687);
and U8865 (N_8865,N_7885,N_7378);
and U8866 (N_8866,N_7460,N_7332);
and U8867 (N_8867,N_7143,N_7844);
nor U8868 (N_8868,N_7721,N_7829);
nor U8869 (N_8869,N_7415,N_7003);
xor U8870 (N_8870,N_7716,N_7709);
xor U8871 (N_8871,N_7097,N_7854);
xor U8872 (N_8872,N_7565,N_7867);
nand U8873 (N_8873,N_7070,N_7184);
and U8874 (N_8874,N_7970,N_7969);
nand U8875 (N_8875,N_7414,N_7736);
xor U8876 (N_8876,N_7540,N_7541);
and U8877 (N_8877,N_7915,N_7546);
or U8878 (N_8878,N_7251,N_7117);
or U8879 (N_8879,N_7324,N_7477);
and U8880 (N_8880,N_7971,N_7459);
or U8881 (N_8881,N_7310,N_7423);
nand U8882 (N_8882,N_7975,N_7683);
nand U8883 (N_8883,N_7022,N_7106);
and U8884 (N_8884,N_7030,N_7888);
or U8885 (N_8885,N_7691,N_7786);
xnor U8886 (N_8886,N_7658,N_7210);
or U8887 (N_8887,N_7592,N_7995);
and U8888 (N_8888,N_7167,N_7128);
or U8889 (N_8889,N_7617,N_7333);
and U8890 (N_8890,N_7307,N_7566);
and U8891 (N_8891,N_7117,N_7909);
and U8892 (N_8892,N_7790,N_7518);
xor U8893 (N_8893,N_7279,N_7558);
xor U8894 (N_8894,N_7723,N_7678);
and U8895 (N_8895,N_7217,N_7453);
and U8896 (N_8896,N_7433,N_7248);
nor U8897 (N_8897,N_7798,N_7103);
or U8898 (N_8898,N_7907,N_7879);
and U8899 (N_8899,N_7078,N_7327);
nor U8900 (N_8900,N_7015,N_7605);
nand U8901 (N_8901,N_7598,N_7104);
xnor U8902 (N_8902,N_7970,N_7818);
nand U8903 (N_8903,N_7360,N_7602);
nand U8904 (N_8904,N_7914,N_7345);
nand U8905 (N_8905,N_7204,N_7281);
or U8906 (N_8906,N_7157,N_7078);
nor U8907 (N_8907,N_7654,N_7805);
nor U8908 (N_8908,N_7128,N_7636);
nand U8909 (N_8909,N_7528,N_7206);
nand U8910 (N_8910,N_7654,N_7316);
xor U8911 (N_8911,N_7164,N_7497);
and U8912 (N_8912,N_7151,N_7878);
and U8913 (N_8913,N_7031,N_7670);
or U8914 (N_8914,N_7032,N_7829);
nor U8915 (N_8915,N_7710,N_7793);
nor U8916 (N_8916,N_7560,N_7162);
nand U8917 (N_8917,N_7718,N_7175);
or U8918 (N_8918,N_7573,N_7666);
nand U8919 (N_8919,N_7089,N_7713);
or U8920 (N_8920,N_7293,N_7670);
and U8921 (N_8921,N_7366,N_7429);
nor U8922 (N_8922,N_7150,N_7853);
nor U8923 (N_8923,N_7224,N_7760);
and U8924 (N_8924,N_7345,N_7507);
nor U8925 (N_8925,N_7433,N_7335);
nor U8926 (N_8926,N_7348,N_7805);
or U8927 (N_8927,N_7588,N_7613);
xor U8928 (N_8928,N_7271,N_7701);
nand U8929 (N_8929,N_7460,N_7975);
nor U8930 (N_8930,N_7324,N_7853);
nand U8931 (N_8931,N_7448,N_7260);
and U8932 (N_8932,N_7978,N_7272);
nand U8933 (N_8933,N_7959,N_7850);
xor U8934 (N_8934,N_7144,N_7794);
nor U8935 (N_8935,N_7829,N_7463);
xnor U8936 (N_8936,N_7229,N_7497);
or U8937 (N_8937,N_7251,N_7578);
and U8938 (N_8938,N_7715,N_7151);
nor U8939 (N_8939,N_7272,N_7808);
nand U8940 (N_8940,N_7384,N_7052);
and U8941 (N_8941,N_7696,N_7772);
nand U8942 (N_8942,N_7469,N_7324);
xnor U8943 (N_8943,N_7413,N_7582);
nor U8944 (N_8944,N_7475,N_7725);
xnor U8945 (N_8945,N_7488,N_7779);
and U8946 (N_8946,N_7851,N_7661);
or U8947 (N_8947,N_7127,N_7137);
and U8948 (N_8948,N_7472,N_7750);
and U8949 (N_8949,N_7363,N_7672);
nor U8950 (N_8950,N_7549,N_7469);
xor U8951 (N_8951,N_7427,N_7664);
xor U8952 (N_8952,N_7403,N_7295);
nor U8953 (N_8953,N_7730,N_7127);
nor U8954 (N_8954,N_7270,N_7670);
nor U8955 (N_8955,N_7081,N_7704);
and U8956 (N_8956,N_7861,N_7924);
xor U8957 (N_8957,N_7676,N_7486);
nor U8958 (N_8958,N_7237,N_7774);
and U8959 (N_8959,N_7783,N_7066);
xnor U8960 (N_8960,N_7554,N_7990);
nand U8961 (N_8961,N_7764,N_7304);
and U8962 (N_8962,N_7656,N_7613);
xor U8963 (N_8963,N_7391,N_7590);
or U8964 (N_8964,N_7524,N_7720);
nor U8965 (N_8965,N_7427,N_7326);
nor U8966 (N_8966,N_7966,N_7944);
or U8967 (N_8967,N_7129,N_7040);
nand U8968 (N_8968,N_7416,N_7105);
or U8969 (N_8969,N_7166,N_7430);
nor U8970 (N_8970,N_7353,N_7708);
nor U8971 (N_8971,N_7743,N_7607);
or U8972 (N_8972,N_7327,N_7428);
or U8973 (N_8973,N_7956,N_7537);
nand U8974 (N_8974,N_7461,N_7252);
or U8975 (N_8975,N_7426,N_7028);
xnor U8976 (N_8976,N_7894,N_7861);
or U8977 (N_8977,N_7634,N_7554);
nor U8978 (N_8978,N_7206,N_7092);
xor U8979 (N_8979,N_7592,N_7700);
nand U8980 (N_8980,N_7074,N_7176);
or U8981 (N_8981,N_7509,N_7801);
nand U8982 (N_8982,N_7881,N_7478);
or U8983 (N_8983,N_7147,N_7388);
nor U8984 (N_8984,N_7273,N_7641);
nand U8985 (N_8985,N_7533,N_7042);
nor U8986 (N_8986,N_7982,N_7511);
or U8987 (N_8987,N_7515,N_7662);
xnor U8988 (N_8988,N_7692,N_7079);
or U8989 (N_8989,N_7040,N_7669);
or U8990 (N_8990,N_7238,N_7566);
nand U8991 (N_8991,N_7816,N_7285);
nand U8992 (N_8992,N_7398,N_7983);
and U8993 (N_8993,N_7655,N_7833);
or U8994 (N_8994,N_7517,N_7661);
or U8995 (N_8995,N_7741,N_7774);
or U8996 (N_8996,N_7537,N_7853);
xor U8997 (N_8997,N_7720,N_7840);
nand U8998 (N_8998,N_7104,N_7618);
and U8999 (N_8999,N_7849,N_7961);
xnor U9000 (N_9000,N_8048,N_8562);
or U9001 (N_9001,N_8682,N_8230);
xnor U9002 (N_9002,N_8716,N_8880);
and U9003 (N_9003,N_8406,N_8264);
nand U9004 (N_9004,N_8885,N_8610);
nor U9005 (N_9005,N_8514,N_8888);
or U9006 (N_9006,N_8666,N_8619);
and U9007 (N_9007,N_8799,N_8893);
nand U9008 (N_9008,N_8464,N_8824);
or U9009 (N_9009,N_8227,N_8652);
nor U9010 (N_9010,N_8973,N_8910);
xor U9011 (N_9011,N_8509,N_8575);
and U9012 (N_9012,N_8774,N_8403);
nor U9013 (N_9013,N_8906,N_8879);
nand U9014 (N_9014,N_8827,N_8712);
or U9015 (N_9015,N_8083,N_8595);
xor U9016 (N_9016,N_8840,N_8030);
nor U9017 (N_9017,N_8484,N_8536);
nand U9018 (N_9018,N_8203,N_8684);
nor U9019 (N_9019,N_8686,N_8458);
nor U9020 (N_9020,N_8635,N_8640);
xor U9021 (N_9021,N_8551,N_8463);
xnor U9022 (N_9022,N_8984,N_8991);
and U9023 (N_9023,N_8376,N_8363);
nor U9024 (N_9024,N_8802,N_8672);
nand U9025 (N_9025,N_8498,N_8823);
nor U9026 (N_9026,N_8947,N_8432);
or U9027 (N_9027,N_8470,N_8095);
and U9028 (N_9028,N_8106,N_8953);
or U9029 (N_9029,N_8613,N_8298);
nor U9030 (N_9030,N_8164,N_8373);
nor U9031 (N_9031,N_8356,N_8244);
and U9032 (N_9032,N_8820,N_8162);
nand U9033 (N_9033,N_8936,N_8590);
nand U9034 (N_9034,N_8100,N_8121);
nor U9035 (N_9035,N_8168,N_8513);
nor U9036 (N_9036,N_8833,N_8070);
nand U9037 (N_9037,N_8239,N_8690);
and U9038 (N_9038,N_8300,N_8451);
xor U9039 (N_9039,N_8648,N_8517);
xor U9040 (N_9040,N_8954,N_8715);
nand U9041 (N_9041,N_8014,N_8500);
xor U9042 (N_9042,N_8612,N_8388);
nand U9043 (N_9043,N_8204,N_8145);
xor U9044 (N_9044,N_8235,N_8579);
xnor U9045 (N_9045,N_8891,N_8767);
xor U9046 (N_9046,N_8442,N_8567);
xnor U9047 (N_9047,N_8104,N_8131);
nor U9048 (N_9048,N_8588,N_8995);
or U9049 (N_9049,N_8245,N_8537);
and U9050 (N_9050,N_8211,N_8952);
and U9051 (N_9051,N_8812,N_8553);
nor U9052 (N_9052,N_8294,N_8447);
and U9053 (N_9053,N_8266,N_8364);
nor U9054 (N_9054,N_8871,N_8308);
nor U9055 (N_9055,N_8876,N_8003);
nor U9056 (N_9056,N_8383,N_8582);
nand U9057 (N_9057,N_8071,N_8404);
xor U9058 (N_9058,N_8696,N_8511);
nand U9059 (N_9059,N_8902,N_8545);
and U9060 (N_9060,N_8217,N_8315);
or U9061 (N_9061,N_8645,N_8603);
and U9062 (N_9062,N_8276,N_8624);
or U9063 (N_9063,N_8172,N_8223);
nand U9064 (N_9064,N_8042,N_8787);
nand U9065 (N_9065,N_8604,N_8477);
nand U9066 (N_9066,N_8560,N_8756);
nand U9067 (N_9067,N_8117,N_8055);
and U9068 (N_9068,N_8249,N_8207);
nor U9069 (N_9069,N_8368,N_8546);
nor U9070 (N_9070,N_8163,N_8704);
nor U9071 (N_9071,N_8053,N_8597);
or U9072 (N_9072,N_8994,N_8090);
and U9073 (N_9073,N_8748,N_8114);
and U9074 (N_9074,N_8968,N_8135);
nand U9075 (N_9075,N_8804,N_8656);
and U9076 (N_9076,N_8448,N_8602);
xnor U9077 (N_9077,N_8864,N_8620);
nor U9078 (N_9078,N_8739,N_8675);
xor U9079 (N_9079,N_8858,N_8830);
nor U9080 (N_9080,N_8951,N_8760);
or U9081 (N_9081,N_8355,N_8969);
and U9082 (N_9082,N_8371,N_8596);
xor U9083 (N_9083,N_8129,N_8111);
nand U9084 (N_9084,N_8169,N_8655);
or U9085 (N_9085,N_8989,N_8002);
xor U9086 (N_9086,N_8057,N_8310);
nand U9087 (N_9087,N_8395,N_8544);
or U9088 (N_9088,N_8870,N_8197);
and U9089 (N_9089,N_8073,N_8487);
or U9090 (N_9090,N_8784,N_8324);
and U9091 (N_9091,N_8456,N_8428);
and U9092 (N_9092,N_8076,N_8261);
nand U9093 (N_9093,N_8307,N_8068);
and U9094 (N_9094,N_8977,N_8455);
nor U9095 (N_9095,N_8279,N_8216);
or U9096 (N_9096,N_8291,N_8650);
nor U9097 (N_9097,N_8846,N_8228);
xor U9098 (N_9098,N_8843,N_8981);
nand U9099 (N_9099,N_8342,N_8155);
nor U9100 (N_9100,N_8658,N_8829);
nor U9101 (N_9101,N_8459,N_8157);
and U9102 (N_9102,N_8637,N_8093);
nor U9103 (N_9103,N_8174,N_8797);
or U9104 (N_9104,N_8584,N_8399);
nand U9105 (N_9105,N_8181,N_8124);
or U9106 (N_9106,N_8443,N_8636);
and U9107 (N_9107,N_8616,N_8894);
and U9108 (N_9108,N_8810,N_8427);
nand U9109 (N_9109,N_8020,N_8743);
or U9110 (N_9110,N_8144,N_8499);
nand U9111 (N_9111,N_8297,N_8109);
xnor U9112 (N_9112,N_8009,N_8449);
xor U9113 (N_9113,N_8015,N_8421);
and U9114 (N_9114,N_8186,N_8420);
xor U9115 (N_9115,N_8099,N_8836);
nor U9116 (N_9116,N_8205,N_8738);
and U9117 (N_9117,N_8761,N_8159);
and U9118 (N_9118,N_8419,N_8081);
nand U9119 (N_9119,N_8401,N_8215);
xor U9120 (N_9120,N_8548,N_8729);
or U9121 (N_9121,N_8505,N_8151);
nand U9122 (N_9122,N_8614,N_8445);
and U9123 (N_9123,N_8054,N_8385);
xor U9124 (N_9124,N_8842,N_8601);
nand U9125 (N_9125,N_8831,N_8328);
and U9126 (N_9126,N_8295,N_8265);
xor U9127 (N_9127,N_8460,N_8576);
xnor U9128 (N_9128,N_8592,N_8961);
nor U9129 (N_9129,N_8649,N_8224);
xnor U9130 (N_9130,N_8097,N_8685);
and U9131 (N_9131,N_8360,N_8754);
nor U9132 (N_9132,N_8632,N_8381);
and U9133 (N_9133,N_8734,N_8524);
nor U9134 (N_9134,N_8102,N_8242);
nor U9135 (N_9135,N_8890,N_8755);
nor U9136 (N_9136,N_8282,N_8200);
and U9137 (N_9137,N_8450,N_8148);
nand U9138 (N_9138,N_8563,N_8764);
and U9139 (N_9139,N_8486,N_8338);
nor U9140 (N_9140,N_8542,N_8859);
or U9141 (N_9141,N_8017,N_8789);
or U9142 (N_9142,N_8949,N_8241);
xnor U9143 (N_9143,N_8865,N_8749);
nor U9144 (N_9144,N_8416,N_8247);
and U9145 (N_9145,N_8886,N_8790);
nand U9146 (N_9146,N_8633,N_8374);
and U9147 (N_9147,N_8158,N_8365);
xor U9148 (N_9148,N_8327,N_8492);
nand U9149 (N_9149,N_8034,N_8725);
nand U9150 (N_9150,N_8944,N_8309);
nor U9151 (N_9151,N_8722,N_8191);
xor U9152 (N_9152,N_8429,N_8663);
nand U9153 (N_9153,N_8924,N_8897);
xnor U9154 (N_9154,N_8084,N_8518);
nand U9155 (N_9155,N_8251,N_8869);
xor U9156 (N_9156,N_8950,N_8958);
or U9157 (N_9157,N_8867,N_8232);
nor U9158 (N_9158,N_8847,N_8999);
xor U9159 (N_9159,N_8063,N_8165);
or U9160 (N_9160,N_8819,N_8642);
nand U9161 (N_9161,N_8959,N_8290);
or U9162 (N_9162,N_8611,N_8801);
or U9163 (N_9163,N_8454,N_8676);
xnor U9164 (N_9164,N_8577,N_8758);
and U9165 (N_9165,N_8007,N_8744);
or U9166 (N_9166,N_8516,N_8378);
xor U9167 (N_9167,N_8439,N_8422);
nand U9168 (N_9168,N_8664,N_8201);
or U9169 (N_9169,N_8120,N_8390);
nand U9170 (N_9170,N_8411,N_8851);
nor U9171 (N_9171,N_8268,N_8948);
nor U9172 (N_9172,N_8293,N_8335);
and U9173 (N_9173,N_8280,N_8219);
or U9174 (N_9174,N_8726,N_8909);
xor U9175 (N_9175,N_8221,N_8461);
and U9176 (N_9176,N_8127,N_8641);
and U9177 (N_9177,N_8375,N_8646);
nor U9178 (N_9178,N_8934,N_8913);
nor U9179 (N_9179,N_8468,N_8092);
nand U9180 (N_9180,N_8581,N_8709);
nand U9181 (N_9181,N_8118,N_8314);
and U9182 (N_9182,N_8996,N_8875);
or U9183 (N_9183,N_8483,N_8036);
or U9184 (N_9184,N_8510,N_8698);
xnor U9185 (N_9185,N_8639,N_8260);
nand U9186 (N_9186,N_8258,N_8096);
or U9187 (N_9187,N_8139,N_8193);
or U9188 (N_9188,N_8705,N_8004);
or U9189 (N_9189,N_8103,N_8688);
nor U9190 (N_9190,N_8476,N_8872);
nand U9191 (N_9191,N_8839,N_8113);
or U9192 (N_9192,N_8182,N_8920);
nand U9193 (N_9193,N_8380,N_8137);
and U9194 (N_9194,N_8019,N_8653);
nand U9195 (N_9195,N_8627,N_8868);
nand U9196 (N_9196,N_8326,N_8933);
and U9197 (N_9197,N_8539,N_8176);
nor U9198 (N_9198,N_8571,N_8010);
xor U9199 (N_9199,N_8707,N_8351);
xor U9200 (N_9200,N_8248,N_8817);
xnor U9201 (N_9201,N_8850,N_8062);
xnor U9202 (N_9202,N_8852,N_8692);
or U9203 (N_9203,N_8552,N_8702);
xor U9204 (N_9204,N_8918,N_8564);
or U9205 (N_9205,N_8803,N_8029);
nand U9206 (N_9206,N_8992,N_8384);
and U9207 (N_9207,N_8046,N_8150);
or U9208 (N_9208,N_8408,N_8878);
nor U9209 (N_9209,N_8252,N_8605);
and U9210 (N_9210,N_8382,N_8533);
nor U9211 (N_9211,N_8337,N_8444);
nand U9212 (N_9212,N_8059,N_8033);
nor U9213 (N_9213,N_8067,N_8853);
xnor U9214 (N_9214,N_8522,N_8066);
xor U9215 (N_9215,N_8208,N_8344);
nor U9216 (N_9216,N_8023,N_8188);
and U9217 (N_9217,N_8462,N_8006);
or U9218 (N_9218,N_8405,N_8746);
xnor U9219 (N_9219,N_8039,N_8431);
nand U9220 (N_9220,N_8914,N_8480);
nand U9221 (N_9221,N_8013,N_8243);
or U9222 (N_9222,N_8695,N_8946);
xnor U9223 (N_9223,N_8369,N_8689);
nand U9224 (N_9224,N_8849,N_8618);
and U9225 (N_9225,N_8674,N_8892);
nor U9226 (N_9226,N_8267,N_8128);
nand U9227 (N_9227,N_8555,N_8359);
or U9228 (N_9228,N_8651,N_8394);
or U9229 (N_9229,N_8400,N_8430);
and U9230 (N_9230,N_8808,N_8474);
nor U9231 (N_9231,N_8680,N_8668);
or U9232 (N_9232,N_8608,N_8926);
xnor U9233 (N_9233,N_8331,N_8643);
or U9234 (N_9234,N_8759,N_8467);
and U9235 (N_9235,N_8209,N_8098);
xor U9236 (N_9236,N_8848,N_8863);
nor U9237 (N_9237,N_8935,N_8506);
xnor U9238 (N_9238,N_8110,N_8001);
and U9239 (N_9239,N_8940,N_8296);
nor U9240 (N_9240,N_8213,N_8101);
nor U9241 (N_9241,N_8329,N_8591);
and U9242 (N_9242,N_8634,N_8358);
xor U9243 (N_9243,N_8805,N_8901);
xor U9244 (N_9244,N_8550,N_8000);
nand U9245 (N_9245,N_8785,N_8983);
nand U9246 (N_9246,N_8900,N_8838);
and U9247 (N_9247,N_8903,N_8418);
nand U9248 (N_9248,N_8987,N_8943);
nor U9249 (N_9249,N_8132,N_8923);
xnor U9250 (N_9250,N_8237,N_8069);
nor U9251 (N_9251,N_8587,N_8183);
nor U9252 (N_9252,N_8975,N_8501);
nand U9253 (N_9253,N_8304,N_8669);
and U9254 (N_9254,N_8153,N_8857);
nor U9255 (N_9255,N_8569,N_8485);
nor U9256 (N_9256,N_8905,N_8038);
xnor U9257 (N_9257,N_8278,N_8222);
nor U9258 (N_9258,N_8299,N_8800);
or U9259 (N_9259,N_8717,N_8319);
nor U9260 (N_9260,N_8889,N_8166);
xnor U9261 (N_9261,N_8988,N_8040);
and U9262 (N_9262,N_8770,N_8154);
and U9263 (N_9263,N_8256,N_8490);
nor U9264 (N_9264,N_8736,N_8077);
and U9265 (N_9265,N_8964,N_8687);
nor U9266 (N_9266,N_8438,N_8021);
nor U9267 (N_9267,N_8465,N_8414);
or U9268 (N_9268,N_8538,N_8731);
and U9269 (N_9269,N_8187,N_8479);
and U9270 (N_9270,N_8678,N_8779);
xor U9271 (N_9271,N_8728,N_8273);
xor U9272 (N_9272,N_8583,N_8044);
xnor U9273 (N_9273,N_8481,N_8482);
or U9274 (N_9274,N_8966,N_8788);
xnor U9275 (N_9275,N_8271,N_8478);
nor U9276 (N_9276,N_8541,N_8711);
nand U9277 (N_9277,N_8699,N_8332);
nor U9278 (N_9278,N_8841,N_8970);
and U9279 (N_9279,N_8737,N_8697);
xor U9280 (N_9280,N_8740,N_8031);
xnor U9281 (N_9281,N_8343,N_8527);
nand U9282 (N_9282,N_8976,N_8339);
or U9283 (N_9283,N_8286,N_8058);
or U9284 (N_9284,N_8446,N_8231);
and U9285 (N_9285,N_8189,N_8349);
or U9286 (N_9286,N_8320,N_8703);
xnor U9287 (N_9287,N_8361,N_8277);
and U9288 (N_9288,N_8845,N_8809);
or U9289 (N_9289,N_8396,N_8520);
or U9290 (N_9290,N_8556,N_8075);
and U9291 (N_9291,N_8362,N_8491);
nand U9292 (N_9292,N_8557,N_8783);
nand U9293 (N_9293,N_8194,N_8771);
nor U9294 (N_9294,N_8367,N_8967);
nor U9295 (N_9295,N_8156,N_8352);
nor U9296 (N_9296,N_8091,N_8125);
nor U9297 (N_9297,N_8469,N_8321);
and U9298 (N_9298,N_8167,N_8873);
nor U9299 (N_9299,N_8519,N_8238);
xnor U9300 (N_9300,N_8775,N_8724);
nand U9301 (N_9301,N_8960,N_8730);
nand U9302 (N_9302,N_8565,N_8255);
or U9303 (N_9303,N_8119,N_8441);
and U9304 (N_9304,N_8559,N_8171);
and U9305 (N_9305,N_8065,N_8939);
nand U9306 (N_9306,N_8932,N_8005);
xnor U9307 (N_9307,N_8741,N_8621);
nand U9308 (N_9308,N_8079,N_8883);
xor U9309 (N_9309,N_8389,N_8617);
xnor U9310 (N_9310,N_8026,N_8670);
and U9311 (N_9311,N_8306,N_8495);
xnor U9312 (N_9312,N_8660,N_8765);
nand U9313 (N_9313,N_8152,N_8625);
nand U9314 (N_9314,N_8622,N_8440);
xor U9315 (N_9315,N_8270,N_8535);
or U9316 (N_9316,N_8757,N_8735);
nor U9317 (N_9317,N_8195,N_8811);
and U9318 (N_9318,N_8078,N_8022);
nand U9319 (N_9319,N_8884,N_8543);
or U9320 (N_9320,N_8473,N_8777);
xnor U9321 (N_9321,N_8816,N_8250);
nor U9322 (N_9322,N_8496,N_8896);
and U9323 (N_9323,N_8629,N_8190);
and U9324 (N_9324,N_8701,N_8866);
or U9325 (N_9325,N_8855,N_8986);
nor U9326 (N_9326,N_8503,N_8654);
and U9327 (N_9327,N_8745,N_8832);
nand U9328 (N_9328,N_8292,N_8844);
xnor U9329 (N_9329,N_8210,N_8313);
and U9330 (N_9330,N_8529,N_8175);
nand U9331 (N_9331,N_8693,N_8628);
nor U9332 (N_9332,N_8435,N_8494);
and U9333 (N_9333,N_8782,N_8115);
nor U9334 (N_9334,N_8379,N_8862);
and U9335 (N_9335,N_8140,N_8028);
and U9336 (N_9336,N_8821,N_8773);
nor U9337 (N_9337,N_8037,N_8957);
and U9338 (N_9338,N_8018,N_8667);
xor U9339 (N_9339,N_8357,N_8087);
and U9340 (N_9340,N_8558,N_8471);
nor U9341 (N_9341,N_8257,N_8874);
and U9342 (N_9342,N_8723,N_8796);
nor U9343 (N_9343,N_8956,N_8061);
nor U9344 (N_9344,N_8919,N_8965);
and U9345 (N_9345,N_8263,N_8554);
xnor U9346 (N_9346,N_8860,N_8887);
and U9347 (N_9347,N_8727,N_8072);
nor U9348 (N_9348,N_8353,N_8751);
nor U9349 (N_9349,N_8283,N_8768);
and U9350 (N_9350,N_8594,N_8915);
xnor U9351 (N_9351,N_8781,N_8142);
xnor U9352 (N_9352,N_8985,N_8206);
nand U9353 (N_9353,N_8807,N_8713);
nor U9354 (N_9354,N_8272,N_8212);
xnor U9355 (N_9355,N_8572,N_8254);
nor U9356 (N_9356,N_8512,N_8185);
or U9357 (N_9357,N_8170,N_8828);
xnor U9358 (N_9358,N_8346,N_8665);
nor U9359 (N_9359,N_8671,N_8990);
xnor U9360 (N_9360,N_8122,N_8130);
nand U9361 (N_9361,N_8141,N_8599);
or U9362 (N_9362,N_8573,N_8942);
and U9363 (N_9363,N_8334,N_8178);
xor U9364 (N_9364,N_8123,N_8963);
nor U9365 (N_9365,N_8927,N_8236);
nand U9366 (N_9366,N_8303,N_8861);
nand U9367 (N_9367,N_8644,N_8045);
xnor U9368 (N_9368,N_8615,N_8762);
and U9369 (N_9369,N_8094,N_8146);
or U9370 (N_9370,N_8753,N_8791);
nand U9371 (N_9371,N_8978,N_8082);
nand U9372 (N_9372,N_8436,N_8532);
or U9373 (N_9373,N_8136,N_8837);
nor U9374 (N_9374,N_8945,N_8147);
xnor U9375 (N_9375,N_8568,N_8218);
nand U9376 (N_9376,N_8877,N_8972);
nand U9377 (N_9377,N_8413,N_8631);
nor U9378 (N_9378,N_8772,N_8229);
nor U9379 (N_9379,N_8600,N_8074);
nor U9380 (N_9380,N_8080,N_8366);
or U9381 (N_9381,N_8708,N_8377);
nand U9382 (N_9382,N_8489,N_8750);
nor U9383 (N_9383,N_8105,N_8997);
and U9384 (N_9384,N_8126,N_8763);
nor U9385 (N_9385,N_8417,N_8302);
xor U9386 (N_9386,N_8931,N_8143);
or U9387 (N_9387,N_8177,N_8035);
nor U9388 (N_9388,N_8856,N_8025);
xor U9389 (N_9389,N_8806,N_8008);
xor U9390 (N_9390,N_8116,N_8694);
or U9391 (N_9391,N_8345,N_8412);
nand U9392 (N_9392,N_8908,N_8240);
xnor U9393 (N_9393,N_8024,N_8312);
nor U9394 (N_9394,N_8180,N_8027);
and U9395 (N_9395,N_8904,N_8937);
xnor U9396 (N_9396,N_8493,N_8160);
nand U9397 (N_9397,N_8769,N_8980);
xor U9398 (N_9398,N_8630,N_8998);
and U9399 (N_9399,N_8882,N_8452);
xnor U9400 (N_9400,N_8198,N_8993);
nor U9401 (N_9401,N_8488,N_8011);
nor U9402 (N_9402,N_8370,N_8246);
nand U9403 (N_9403,N_8971,N_8881);
and U9404 (N_9404,N_8916,N_8792);
or U9405 (N_9405,N_8928,N_8659);
and U9406 (N_9406,N_8391,N_8813);
xnor U9407 (N_9407,N_8393,N_8415);
xor U9408 (N_9408,N_8714,N_8609);
xnor U9409 (N_9409,N_8929,N_8794);
xor U9410 (N_9410,N_8386,N_8525);
and U9411 (N_9411,N_8289,N_8173);
xnor U9412 (N_9412,N_8134,N_8220);
or U9413 (N_9413,N_8284,N_8161);
xor U9414 (N_9414,N_8398,N_8340);
nand U9415 (N_9415,N_8281,N_8107);
nor U9416 (N_9416,N_8043,N_8262);
nand U9417 (N_9417,N_8917,N_8508);
or U9418 (N_9418,N_8259,N_8347);
nor U9419 (N_9419,N_8409,N_8333);
xnor U9420 (N_9420,N_8834,N_8673);
nand U9421 (N_9421,N_8350,N_8798);
nor U9422 (N_9422,N_8088,N_8912);
or U9423 (N_9423,N_8911,N_8607);
or U9424 (N_9424,N_8531,N_8497);
xor U9425 (N_9425,N_8234,N_8606);
and U9426 (N_9426,N_8287,N_8457);
nor U9427 (N_9427,N_8433,N_8051);
or U9428 (N_9428,N_8330,N_8822);
or U9429 (N_9429,N_8835,N_8434);
or U9430 (N_9430,N_8311,N_8086);
and U9431 (N_9431,N_8895,N_8196);
nor U9432 (N_9432,N_8534,N_8016);
xor U9433 (N_9433,N_8305,N_8528);
nand U9434 (N_9434,N_8700,N_8089);
xnor U9435 (N_9435,N_8184,N_8192);
xor U9436 (N_9436,N_8348,N_8341);
or U9437 (N_9437,N_8566,N_8778);
nor U9438 (N_9438,N_8854,N_8226);
and U9439 (N_9439,N_8032,N_8706);
or U9440 (N_9440,N_8392,N_8780);
and U9441 (N_9441,N_8372,N_8275);
nand U9442 (N_9442,N_8472,N_8199);
and U9443 (N_9443,N_8225,N_8410);
and U9444 (N_9444,N_8626,N_8683);
and U9445 (N_9445,N_8056,N_8776);
nand U9446 (N_9446,N_8589,N_8826);
nand U9447 (N_9447,N_8719,N_8732);
or U9448 (N_9448,N_8504,N_8586);
or U9449 (N_9449,N_8766,N_8955);
and U9450 (N_9450,N_8317,N_8540);
nor U9451 (N_9451,N_8064,N_8747);
nand U9452 (N_9452,N_8336,N_8941);
xor U9453 (N_9453,N_8233,N_8325);
or U9454 (N_9454,N_8530,N_8424);
or U9455 (N_9455,N_8814,N_8466);
and U9456 (N_9456,N_8523,N_8285);
xnor U9457 (N_9457,N_8052,N_8301);
nand U9458 (N_9458,N_8561,N_8982);
nor U9459 (N_9459,N_8407,N_8657);
and U9460 (N_9460,N_8108,N_8681);
or U9461 (N_9461,N_8752,N_8580);
nor U9462 (N_9462,N_8638,N_8149);
or U9463 (N_9463,N_8085,N_8041);
and U9464 (N_9464,N_8047,N_8049);
nand U9465 (N_9465,N_8138,N_8974);
nand U9466 (N_9466,N_8718,N_8930);
or U9467 (N_9467,N_8316,N_8733);
nor U9468 (N_9468,N_8721,N_8274);
nor U9469 (N_9469,N_8214,N_8526);
and U9470 (N_9470,N_8507,N_8426);
nand U9471 (N_9471,N_8521,N_8898);
nand U9472 (N_9472,N_8179,N_8815);
xnor U9473 (N_9473,N_8318,N_8437);
nand U9474 (N_9474,N_8547,N_8962);
nand U9475 (N_9475,N_8720,N_8679);
xnor U9476 (N_9476,N_8133,N_8742);
nand U9477 (N_9477,N_8578,N_8202);
and U9478 (N_9478,N_8397,N_8050);
or U9479 (N_9479,N_8585,N_8549);
nor U9480 (N_9480,N_8677,N_8574);
nor U9481 (N_9481,N_8593,N_8402);
and U9482 (N_9482,N_8795,N_8899);
and U9483 (N_9483,N_8818,N_8922);
nor U9484 (N_9484,N_8662,N_8323);
and U9485 (N_9485,N_8288,N_8012);
xor U9486 (N_9486,N_8423,N_8387);
nand U9487 (N_9487,N_8907,N_8661);
and U9488 (N_9488,N_8475,N_8425);
and U9489 (N_9489,N_8979,N_8786);
or U9490 (N_9490,N_8938,N_8570);
and U9491 (N_9491,N_8502,N_8925);
and U9492 (N_9492,N_8453,N_8710);
nand U9493 (N_9493,N_8112,N_8623);
and U9494 (N_9494,N_8691,N_8825);
xnor U9495 (N_9495,N_8253,N_8647);
or U9496 (N_9496,N_8269,N_8921);
and U9497 (N_9497,N_8598,N_8354);
and U9498 (N_9498,N_8322,N_8515);
or U9499 (N_9499,N_8793,N_8060);
nor U9500 (N_9500,N_8591,N_8446);
nor U9501 (N_9501,N_8506,N_8171);
or U9502 (N_9502,N_8218,N_8471);
nor U9503 (N_9503,N_8042,N_8166);
or U9504 (N_9504,N_8359,N_8088);
xor U9505 (N_9505,N_8185,N_8315);
nand U9506 (N_9506,N_8576,N_8163);
nor U9507 (N_9507,N_8938,N_8482);
nor U9508 (N_9508,N_8600,N_8384);
xor U9509 (N_9509,N_8145,N_8687);
nor U9510 (N_9510,N_8031,N_8221);
nand U9511 (N_9511,N_8183,N_8075);
nor U9512 (N_9512,N_8828,N_8144);
xor U9513 (N_9513,N_8645,N_8929);
or U9514 (N_9514,N_8057,N_8506);
nand U9515 (N_9515,N_8327,N_8391);
and U9516 (N_9516,N_8246,N_8828);
nand U9517 (N_9517,N_8733,N_8889);
or U9518 (N_9518,N_8440,N_8866);
or U9519 (N_9519,N_8254,N_8256);
or U9520 (N_9520,N_8698,N_8416);
nor U9521 (N_9521,N_8888,N_8407);
nand U9522 (N_9522,N_8910,N_8624);
nand U9523 (N_9523,N_8079,N_8597);
and U9524 (N_9524,N_8818,N_8891);
xor U9525 (N_9525,N_8394,N_8479);
xor U9526 (N_9526,N_8730,N_8545);
nor U9527 (N_9527,N_8238,N_8912);
and U9528 (N_9528,N_8667,N_8536);
xor U9529 (N_9529,N_8900,N_8922);
nand U9530 (N_9530,N_8777,N_8933);
nand U9531 (N_9531,N_8471,N_8191);
xnor U9532 (N_9532,N_8982,N_8249);
xnor U9533 (N_9533,N_8138,N_8553);
or U9534 (N_9534,N_8866,N_8544);
or U9535 (N_9535,N_8021,N_8556);
nor U9536 (N_9536,N_8610,N_8979);
xor U9537 (N_9537,N_8358,N_8324);
and U9538 (N_9538,N_8122,N_8256);
or U9539 (N_9539,N_8158,N_8498);
nand U9540 (N_9540,N_8999,N_8348);
xnor U9541 (N_9541,N_8385,N_8320);
xor U9542 (N_9542,N_8980,N_8981);
and U9543 (N_9543,N_8593,N_8059);
and U9544 (N_9544,N_8770,N_8293);
xnor U9545 (N_9545,N_8212,N_8576);
or U9546 (N_9546,N_8687,N_8654);
or U9547 (N_9547,N_8186,N_8742);
or U9548 (N_9548,N_8502,N_8556);
xnor U9549 (N_9549,N_8628,N_8094);
and U9550 (N_9550,N_8943,N_8981);
or U9551 (N_9551,N_8828,N_8490);
nor U9552 (N_9552,N_8667,N_8677);
xor U9553 (N_9553,N_8800,N_8458);
xor U9554 (N_9554,N_8871,N_8688);
nand U9555 (N_9555,N_8630,N_8632);
or U9556 (N_9556,N_8159,N_8597);
and U9557 (N_9557,N_8164,N_8194);
xor U9558 (N_9558,N_8825,N_8444);
and U9559 (N_9559,N_8826,N_8986);
nand U9560 (N_9560,N_8382,N_8904);
nand U9561 (N_9561,N_8279,N_8435);
xnor U9562 (N_9562,N_8339,N_8953);
nor U9563 (N_9563,N_8545,N_8094);
xnor U9564 (N_9564,N_8501,N_8286);
or U9565 (N_9565,N_8880,N_8236);
nand U9566 (N_9566,N_8137,N_8822);
nor U9567 (N_9567,N_8298,N_8238);
and U9568 (N_9568,N_8222,N_8717);
nand U9569 (N_9569,N_8863,N_8676);
and U9570 (N_9570,N_8312,N_8158);
or U9571 (N_9571,N_8939,N_8543);
nand U9572 (N_9572,N_8725,N_8963);
nand U9573 (N_9573,N_8885,N_8438);
nor U9574 (N_9574,N_8331,N_8794);
or U9575 (N_9575,N_8993,N_8494);
and U9576 (N_9576,N_8776,N_8917);
nand U9577 (N_9577,N_8834,N_8573);
or U9578 (N_9578,N_8569,N_8588);
and U9579 (N_9579,N_8747,N_8877);
and U9580 (N_9580,N_8530,N_8109);
or U9581 (N_9581,N_8425,N_8545);
nor U9582 (N_9582,N_8285,N_8930);
and U9583 (N_9583,N_8625,N_8832);
xnor U9584 (N_9584,N_8670,N_8201);
nand U9585 (N_9585,N_8796,N_8193);
or U9586 (N_9586,N_8379,N_8922);
nand U9587 (N_9587,N_8374,N_8841);
nand U9588 (N_9588,N_8474,N_8332);
nor U9589 (N_9589,N_8663,N_8745);
xor U9590 (N_9590,N_8134,N_8320);
or U9591 (N_9591,N_8139,N_8336);
nand U9592 (N_9592,N_8478,N_8704);
nor U9593 (N_9593,N_8935,N_8167);
nand U9594 (N_9594,N_8069,N_8285);
or U9595 (N_9595,N_8503,N_8636);
and U9596 (N_9596,N_8814,N_8380);
nand U9597 (N_9597,N_8592,N_8965);
nor U9598 (N_9598,N_8476,N_8329);
nor U9599 (N_9599,N_8849,N_8121);
or U9600 (N_9600,N_8043,N_8430);
xor U9601 (N_9601,N_8282,N_8851);
and U9602 (N_9602,N_8750,N_8430);
nand U9603 (N_9603,N_8189,N_8661);
nor U9604 (N_9604,N_8546,N_8374);
and U9605 (N_9605,N_8042,N_8484);
nand U9606 (N_9606,N_8683,N_8467);
or U9607 (N_9607,N_8350,N_8147);
or U9608 (N_9608,N_8222,N_8554);
nand U9609 (N_9609,N_8603,N_8375);
xor U9610 (N_9610,N_8800,N_8688);
or U9611 (N_9611,N_8663,N_8305);
and U9612 (N_9612,N_8154,N_8735);
nor U9613 (N_9613,N_8410,N_8084);
and U9614 (N_9614,N_8208,N_8611);
or U9615 (N_9615,N_8417,N_8079);
nor U9616 (N_9616,N_8437,N_8604);
or U9617 (N_9617,N_8778,N_8453);
or U9618 (N_9618,N_8917,N_8550);
xor U9619 (N_9619,N_8450,N_8558);
nand U9620 (N_9620,N_8858,N_8007);
nor U9621 (N_9621,N_8805,N_8798);
nand U9622 (N_9622,N_8873,N_8048);
xnor U9623 (N_9623,N_8725,N_8490);
and U9624 (N_9624,N_8104,N_8892);
or U9625 (N_9625,N_8965,N_8944);
nand U9626 (N_9626,N_8716,N_8372);
and U9627 (N_9627,N_8735,N_8869);
nand U9628 (N_9628,N_8571,N_8584);
or U9629 (N_9629,N_8781,N_8298);
and U9630 (N_9630,N_8781,N_8669);
and U9631 (N_9631,N_8177,N_8189);
xor U9632 (N_9632,N_8987,N_8273);
xor U9633 (N_9633,N_8668,N_8740);
or U9634 (N_9634,N_8696,N_8978);
nand U9635 (N_9635,N_8364,N_8520);
or U9636 (N_9636,N_8987,N_8934);
xnor U9637 (N_9637,N_8301,N_8594);
nor U9638 (N_9638,N_8083,N_8277);
and U9639 (N_9639,N_8440,N_8346);
nand U9640 (N_9640,N_8830,N_8926);
and U9641 (N_9641,N_8144,N_8649);
xor U9642 (N_9642,N_8743,N_8779);
or U9643 (N_9643,N_8087,N_8106);
nand U9644 (N_9644,N_8046,N_8622);
nor U9645 (N_9645,N_8269,N_8828);
or U9646 (N_9646,N_8279,N_8398);
nor U9647 (N_9647,N_8182,N_8046);
and U9648 (N_9648,N_8933,N_8165);
or U9649 (N_9649,N_8573,N_8712);
xnor U9650 (N_9650,N_8646,N_8990);
or U9651 (N_9651,N_8948,N_8805);
nand U9652 (N_9652,N_8992,N_8863);
nor U9653 (N_9653,N_8094,N_8040);
and U9654 (N_9654,N_8708,N_8852);
nand U9655 (N_9655,N_8628,N_8833);
or U9656 (N_9656,N_8827,N_8947);
nor U9657 (N_9657,N_8010,N_8045);
xnor U9658 (N_9658,N_8244,N_8930);
nand U9659 (N_9659,N_8007,N_8548);
nor U9660 (N_9660,N_8900,N_8813);
xnor U9661 (N_9661,N_8601,N_8117);
or U9662 (N_9662,N_8398,N_8288);
nand U9663 (N_9663,N_8042,N_8581);
and U9664 (N_9664,N_8658,N_8605);
xnor U9665 (N_9665,N_8824,N_8754);
nand U9666 (N_9666,N_8979,N_8229);
nor U9667 (N_9667,N_8381,N_8650);
nor U9668 (N_9668,N_8765,N_8871);
nor U9669 (N_9669,N_8095,N_8740);
nor U9670 (N_9670,N_8181,N_8250);
xnor U9671 (N_9671,N_8169,N_8918);
nand U9672 (N_9672,N_8679,N_8816);
or U9673 (N_9673,N_8235,N_8468);
nand U9674 (N_9674,N_8771,N_8815);
xor U9675 (N_9675,N_8494,N_8715);
nand U9676 (N_9676,N_8726,N_8930);
and U9677 (N_9677,N_8446,N_8196);
or U9678 (N_9678,N_8708,N_8819);
and U9679 (N_9679,N_8708,N_8884);
nor U9680 (N_9680,N_8342,N_8338);
or U9681 (N_9681,N_8687,N_8871);
nand U9682 (N_9682,N_8589,N_8458);
xnor U9683 (N_9683,N_8525,N_8654);
xor U9684 (N_9684,N_8421,N_8816);
and U9685 (N_9685,N_8824,N_8859);
nand U9686 (N_9686,N_8246,N_8481);
xor U9687 (N_9687,N_8057,N_8270);
and U9688 (N_9688,N_8879,N_8510);
or U9689 (N_9689,N_8106,N_8854);
xor U9690 (N_9690,N_8310,N_8397);
or U9691 (N_9691,N_8507,N_8340);
or U9692 (N_9692,N_8187,N_8050);
or U9693 (N_9693,N_8686,N_8901);
or U9694 (N_9694,N_8941,N_8978);
or U9695 (N_9695,N_8500,N_8194);
xnor U9696 (N_9696,N_8533,N_8039);
nand U9697 (N_9697,N_8459,N_8970);
or U9698 (N_9698,N_8898,N_8697);
or U9699 (N_9699,N_8403,N_8222);
nor U9700 (N_9700,N_8448,N_8003);
xnor U9701 (N_9701,N_8658,N_8471);
nand U9702 (N_9702,N_8907,N_8041);
and U9703 (N_9703,N_8656,N_8464);
nor U9704 (N_9704,N_8499,N_8932);
and U9705 (N_9705,N_8289,N_8271);
nor U9706 (N_9706,N_8770,N_8103);
nor U9707 (N_9707,N_8164,N_8076);
xnor U9708 (N_9708,N_8135,N_8794);
nor U9709 (N_9709,N_8890,N_8562);
or U9710 (N_9710,N_8250,N_8890);
and U9711 (N_9711,N_8040,N_8775);
or U9712 (N_9712,N_8866,N_8538);
xor U9713 (N_9713,N_8537,N_8254);
xor U9714 (N_9714,N_8669,N_8473);
nor U9715 (N_9715,N_8279,N_8336);
nor U9716 (N_9716,N_8309,N_8924);
and U9717 (N_9717,N_8079,N_8304);
nand U9718 (N_9718,N_8161,N_8098);
nand U9719 (N_9719,N_8014,N_8854);
xnor U9720 (N_9720,N_8915,N_8647);
nand U9721 (N_9721,N_8318,N_8555);
xnor U9722 (N_9722,N_8135,N_8554);
xnor U9723 (N_9723,N_8198,N_8328);
xor U9724 (N_9724,N_8298,N_8561);
or U9725 (N_9725,N_8946,N_8574);
nand U9726 (N_9726,N_8669,N_8977);
and U9727 (N_9727,N_8486,N_8299);
nand U9728 (N_9728,N_8551,N_8990);
nand U9729 (N_9729,N_8620,N_8826);
xnor U9730 (N_9730,N_8719,N_8377);
nand U9731 (N_9731,N_8145,N_8746);
xor U9732 (N_9732,N_8245,N_8017);
and U9733 (N_9733,N_8887,N_8324);
nand U9734 (N_9734,N_8541,N_8122);
xnor U9735 (N_9735,N_8096,N_8836);
nor U9736 (N_9736,N_8825,N_8445);
and U9737 (N_9737,N_8508,N_8979);
nand U9738 (N_9738,N_8743,N_8267);
or U9739 (N_9739,N_8585,N_8358);
or U9740 (N_9740,N_8554,N_8086);
nand U9741 (N_9741,N_8182,N_8265);
xor U9742 (N_9742,N_8929,N_8110);
xor U9743 (N_9743,N_8141,N_8686);
nand U9744 (N_9744,N_8184,N_8839);
nand U9745 (N_9745,N_8293,N_8320);
and U9746 (N_9746,N_8260,N_8595);
xor U9747 (N_9747,N_8625,N_8217);
and U9748 (N_9748,N_8507,N_8368);
and U9749 (N_9749,N_8265,N_8236);
or U9750 (N_9750,N_8193,N_8120);
or U9751 (N_9751,N_8226,N_8317);
nor U9752 (N_9752,N_8980,N_8305);
and U9753 (N_9753,N_8167,N_8883);
nand U9754 (N_9754,N_8400,N_8877);
or U9755 (N_9755,N_8441,N_8763);
and U9756 (N_9756,N_8304,N_8744);
and U9757 (N_9757,N_8439,N_8773);
nor U9758 (N_9758,N_8388,N_8282);
xor U9759 (N_9759,N_8379,N_8109);
xor U9760 (N_9760,N_8571,N_8117);
xor U9761 (N_9761,N_8035,N_8215);
and U9762 (N_9762,N_8334,N_8720);
nand U9763 (N_9763,N_8529,N_8070);
nand U9764 (N_9764,N_8637,N_8665);
and U9765 (N_9765,N_8735,N_8850);
nand U9766 (N_9766,N_8571,N_8375);
nor U9767 (N_9767,N_8116,N_8178);
xor U9768 (N_9768,N_8275,N_8775);
or U9769 (N_9769,N_8564,N_8210);
and U9770 (N_9770,N_8390,N_8799);
nor U9771 (N_9771,N_8064,N_8032);
and U9772 (N_9772,N_8967,N_8262);
or U9773 (N_9773,N_8206,N_8309);
and U9774 (N_9774,N_8377,N_8753);
or U9775 (N_9775,N_8214,N_8904);
nand U9776 (N_9776,N_8034,N_8710);
and U9777 (N_9777,N_8430,N_8745);
nand U9778 (N_9778,N_8949,N_8087);
xor U9779 (N_9779,N_8931,N_8575);
nand U9780 (N_9780,N_8056,N_8113);
xor U9781 (N_9781,N_8988,N_8710);
nor U9782 (N_9782,N_8186,N_8324);
nor U9783 (N_9783,N_8532,N_8843);
xnor U9784 (N_9784,N_8377,N_8000);
nor U9785 (N_9785,N_8615,N_8998);
nand U9786 (N_9786,N_8307,N_8128);
nor U9787 (N_9787,N_8021,N_8728);
nor U9788 (N_9788,N_8117,N_8852);
xnor U9789 (N_9789,N_8680,N_8613);
or U9790 (N_9790,N_8298,N_8072);
and U9791 (N_9791,N_8533,N_8182);
nor U9792 (N_9792,N_8125,N_8598);
or U9793 (N_9793,N_8369,N_8392);
nor U9794 (N_9794,N_8835,N_8356);
or U9795 (N_9795,N_8565,N_8658);
and U9796 (N_9796,N_8234,N_8552);
xnor U9797 (N_9797,N_8951,N_8241);
or U9798 (N_9798,N_8889,N_8078);
or U9799 (N_9799,N_8532,N_8846);
and U9800 (N_9800,N_8985,N_8676);
nand U9801 (N_9801,N_8196,N_8001);
nor U9802 (N_9802,N_8933,N_8970);
nand U9803 (N_9803,N_8496,N_8503);
nor U9804 (N_9804,N_8024,N_8672);
and U9805 (N_9805,N_8943,N_8656);
or U9806 (N_9806,N_8305,N_8780);
and U9807 (N_9807,N_8897,N_8829);
and U9808 (N_9808,N_8705,N_8362);
xor U9809 (N_9809,N_8376,N_8413);
or U9810 (N_9810,N_8420,N_8735);
nand U9811 (N_9811,N_8470,N_8151);
nand U9812 (N_9812,N_8404,N_8793);
xor U9813 (N_9813,N_8832,N_8428);
nor U9814 (N_9814,N_8507,N_8423);
nor U9815 (N_9815,N_8508,N_8974);
and U9816 (N_9816,N_8543,N_8809);
nor U9817 (N_9817,N_8623,N_8019);
and U9818 (N_9818,N_8714,N_8509);
or U9819 (N_9819,N_8871,N_8064);
xnor U9820 (N_9820,N_8427,N_8930);
nor U9821 (N_9821,N_8915,N_8096);
nand U9822 (N_9822,N_8717,N_8047);
nor U9823 (N_9823,N_8463,N_8757);
nand U9824 (N_9824,N_8825,N_8697);
xor U9825 (N_9825,N_8806,N_8995);
nand U9826 (N_9826,N_8415,N_8198);
nor U9827 (N_9827,N_8118,N_8161);
xnor U9828 (N_9828,N_8487,N_8244);
nand U9829 (N_9829,N_8760,N_8917);
or U9830 (N_9830,N_8364,N_8987);
xnor U9831 (N_9831,N_8714,N_8591);
nand U9832 (N_9832,N_8870,N_8363);
nor U9833 (N_9833,N_8536,N_8312);
nor U9834 (N_9834,N_8858,N_8443);
and U9835 (N_9835,N_8640,N_8287);
nor U9836 (N_9836,N_8510,N_8455);
nand U9837 (N_9837,N_8264,N_8193);
nor U9838 (N_9838,N_8360,N_8373);
xor U9839 (N_9839,N_8352,N_8727);
nor U9840 (N_9840,N_8409,N_8195);
nand U9841 (N_9841,N_8113,N_8376);
xor U9842 (N_9842,N_8341,N_8441);
or U9843 (N_9843,N_8581,N_8562);
or U9844 (N_9844,N_8149,N_8428);
and U9845 (N_9845,N_8551,N_8794);
or U9846 (N_9846,N_8962,N_8376);
xnor U9847 (N_9847,N_8920,N_8651);
xor U9848 (N_9848,N_8754,N_8369);
and U9849 (N_9849,N_8843,N_8396);
xor U9850 (N_9850,N_8082,N_8894);
and U9851 (N_9851,N_8570,N_8364);
nand U9852 (N_9852,N_8352,N_8077);
nor U9853 (N_9853,N_8750,N_8302);
and U9854 (N_9854,N_8283,N_8541);
and U9855 (N_9855,N_8021,N_8977);
and U9856 (N_9856,N_8779,N_8260);
nand U9857 (N_9857,N_8069,N_8527);
and U9858 (N_9858,N_8745,N_8457);
nand U9859 (N_9859,N_8297,N_8598);
or U9860 (N_9860,N_8247,N_8053);
xnor U9861 (N_9861,N_8778,N_8708);
and U9862 (N_9862,N_8956,N_8290);
nor U9863 (N_9863,N_8474,N_8377);
nand U9864 (N_9864,N_8545,N_8228);
xor U9865 (N_9865,N_8318,N_8439);
and U9866 (N_9866,N_8620,N_8676);
and U9867 (N_9867,N_8174,N_8967);
xnor U9868 (N_9868,N_8338,N_8907);
and U9869 (N_9869,N_8284,N_8179);
and U9870 (N_9870,N_8378,N_8679);
nor U9871 (N_9871,N_8380,N_8387);
or U9872 (N_9872,N_8796,N_8850);
or U9873 (N_9873,N_8382,N_8437);
and U9874 (N_9874,N_8446,N_8015);
nor U9875 (N_9875,N_8878,N_8641);
and U9876 (N_9876,N_8155,N_8224);
nand U9877 (N_9877,N_8610,N_8611);
nor U9878 (N_9878,N_8769,N_8071);
xor U9879 (N_9879,N_8802,N_8479);
or U9880 (N_9880,N_8382,N_8571);
or U9881 (N_9881,N_8525,N_8642);
or U9882 (N_9882,N_8587,N_8382);
or U9883 (N_9883,N_8657,N_8677);
and U9884 (N_9884,N_8494,N_8019);
nand U9885 (N_9885,N_8050,N_8029);
xor U9886 (N_9886,N_8284,N_8173);
nand U9887 (N_9887,N_8054,N_8928);
xnor U9888 (N_9888,N_8850,N_8748);
or U9889 (N_9889,N_8073,N_8443);
xnor U9890 (N_9890,N_8406,N_8693);
and U9891 (N_9891,N_8258,N_8705);
xor U9892 (N_9892,N_8331,N_8618);
nor U9893 (N_9893,N_8566,N_8698);
nor U9894 (N_9894,N_8801,N_8564);
xnor U9895 (N_9895,N_8603,N_8581);
nor U9896 (N_9896,N_8773,N_8431);
and U9897 (N_9897,N_8442,N_8483);
xor U9898 (N_9898,N_8540,N_8815);
nor U9899 (N_9899,N_8400,N_8323);
nor U9900 (N_9900,N_8488,N_8199);
xnor U9901 (N_9901,N_8478,N_8187);
or U9902 (N_9902,N_8099,N_8042);
nor U9903 (N_9903,N_8753,N_8863);
and U9904 (N_9904,N_8548,N_8580);
nor U9905 (N_9905,N_8022,N_8828);
nand U9906 (N_9906,N_8625,N_8171);
nor U9907 (N_9907,N_8250,N_8919);
nor U9908 (N_9908,N_8989,N_8969);
nor U9909 (N_9909,N_8720,N_8961);
or U9910 (N_9910,N_8252,N_8446);
and U9911 (N_9911,N_8729,N_8295);
xor U9912 (N_9912,N_8309,N_8081);
or U9913 (N_9913,N_8597,N_8612);
or U9914 (N_9914,N_8738,N_8292);
and U9915 (N_9915,N_8208,N_8328);
xnor U9916 (N_9916,N_8091,N_8611);
xor U9917 (N_9917,N_8298,N_8818);
or U9918 (N_9918,N_8120,N_8123);
and U9919 (N_9919,N_8250,N_8783);
xnor U9920 (N_9920,N_8665,N_8930);
nand U9921 (N_9921,N_8959,N_8898);
or U9922 (N_9922,N_8627,N_8794);
xnor U9923 (N_9923,N_8488,N_8052);
xor U9924 (N_9924,N_8528,N_8977);
and U9925 (N_9925,N_8829,N_8423);
xor U9926 (N_9926,N_8717,N_8938);
nand U9927 (N_9927,N_8128,N_8359);
nand U9928 (N_9928,N_8018,N_8127);
nor U9929 (N_9929,N_8338,N_8985);
and U9930 (N_9930,N_8464,N_8318);
and U9931 (N_9931,N_8653,N_8480);
nand U9932 (N_9932,N_8396,N_8884);
nand U9933 (N_9933,N_8912,N_8231);
nand U9934 (N_9934,N_8180,N_8366);
nor U9935 (N_9935,N_8936,N_8239);
xnor U9936 (N_9936,N_8623,N_8295);
and U9937 (N_9937,N_8143,N_8753);
or U9938 (N_9938,N_8176,N_8748);
xnor U9939 (N_9939,N_8352,N_8942);
and U9940 (N_9940,N_8189,N_8439);
nand U9941 (N_9941,N_8507,N_8471);
xor U9942 (N_9942,N_8603,N_8405);
or U9943 (N_9943,N_8264,N_8479);
and U9944 (N_9944,N_8556,N_8878);
nor U9945 (N_9945,N_8984,N_8611);
nand U9946 (N_9946,N_8265,N_8462);
xor U9947 (N_9947,N_8919,N_8764);
nor U9948 (N_9948,N_8435,N_8892);
xor U9949 (N_9949,N_8600,N_8254);
nor U9950 (N_9950,N_8269,N_8528);
or U9951 (N_9951,N_8930,N_8931);
nor U9952 (N_9952,N_8281,N_8395);
or U9953 (N_9953,N_8345,N_8238);
nand U9954 (N_9954,N_8810,N_8508);
xor U9955 (N_9955,N_8415,N_8686);
nand U9956 (N_9956,N_8208,N_8520);
nand U9957 (N_9957,N_8300,N_8303);
or U9958 (N_9958,N_8132,N_8658);
nor U9959 (N_9959,N_8176,N_8165);
xor U9960 (N_9960,N_8887,N_8062);
nor U9961 (N_9961,N_8192,N_8518);
nor U9962 (N_9962,N_8491,N_8048);
or U9963 (N_9963,N_8138,N_8050);
nand U9964 (N_9964,N_8743,N_8692);
and U9965 (N_9965,N_8775,N_8867);
and U9966 (N_9966,N_8126,N_8637);
or U9967 (N_9967,N_8871,N_8069);
nand U9968 (N_9968,N_8665,N_8977);
xnor U9969 (N_9969,N_8409,N_8857);
or U9970 (N_9970,N_8268,N_8774);
xnor U9971 (N_9971,N_8008,N_8427);
nor U9972 (N_9972,N_8092,N_8165);
nor U9973 (N_9973,N_8239,N_8523);
xor U9974 (N_9974,N_8279,N_8901);
and U9975 (N_9975,N_8198,N_8201);
nand U9976 (N_9976,N_8431,N_8256);
and U9977 (N_9977,N_8024,N_8311);
nor U9978 (N_9978,N_8475,N_8668);
nor U9979 (N_9979,N_8929,N_8428);
and U9980 (N_9980,N_8196,N_8862);
and U9981 (N_9981,N_8618,N_8641);
nand U9982 (N_9982,N_8051,N_8973);
xor U9983 (N_9983,N_8026,N_8545);
nor U9984 (N_9984,N_8024,N_8100);
and U9985 (N_9985,N_8312,N_8123);
nand U9986 (N_9986,N_8183,N_8166);
xnor U9987 (N_9987,N_8951,N_8837);
nand U9988 (N_9988,N_8549,N_8543);
or U9989 (N_9989,N_8522,N_8435);
nand U9990 (N_9990,N_8272,N_8039);
nor U9991 (N_9991,N_8409,N_8710);
and U9992 (N_9992,N_8807,N_8626);
or U9993 (N_9993,N_8812,N_8123);
nand U9994 (N_9994,N_8797,N_8343);
or U9995 (N_9995,N_8636,N_8958);
nor U9996 (N_9996,N_8807,N_8860);
nand U9997 (N_9997,N_8605,N_8631);
nand U9998 (N_9998,N_8564,N_8966);
xnor U9999 (N_9999,N_8785,N_8499);
nand UO_0 (O_0,N_9942,N_9032);
xor UO_1 (O_1,N_9462,N_9479);
nand UO_2 (O_2,N_9584,N_9577);
nor UO_3 (O_3,N_9294,N_9896);
and UO_4 (O_4,N_9389,N_9680);
xor UO_5 (O_5,N_9227,N_9533);
and UO_6 (O_6,N_9417,N_9947);
nand UO_7 (O_7,N_9373,N_9642);
nand UO_8 (O_8,N_9137,N_9847);
and UO_9 (O_9,N_9837,N_9254);
xor UO_10 (O_10,N_9511,N_9025);
or UO_11 (O_11,N_9496,N_9284);
xor UO_12 (O_12,N_9201,N_9569);
nor UO_13 (O_13,N_9517,N_9629);
or UO_14 (O_14,N_9066,N_9377);
or UO_15 (O_15,N_9428,N_9492);
xor UO_16 (O_16,N_9572,N_9676);
nand UO_17 (O_17,N_9897,N_9898);
or UO_18 (O_18,N_9705,N_9369);
or UO_19 (O_19,N_9279,N_9784);
or UO_20 (O_20,N_9114,N_9487);
or UO_21 (O_21,N_9594,N_9667);
or UO_22 (O_22,N_9356,N_9693);
nand UO_23 (O_23,N_9931,N_9925);
or UO_24 (O_24,N_9226,N_9042);
nand UO_25 (O_25,N_9790,N_9502);
or UO_26 (O_26,N_9873,N_9368);
or UO_27 (O_27,N_9851,N_9240);
or UO_28 (O_28,N_9628,N_9478);
or UO_29 (O_29,N_9688,N_9681);
or UO_30 (O_30,N_9384,N_9600);
xnor UO_31 (O_31,N_9349,N_9080);
and UO_32 (O_32,N_9464,N_9340);
and UO_33 (O_33,N_9625,N_9235);
or UO_34 (O_34,N_9855,N_9123);
or UO_35 (O_35,N_9909,N_9923);
xor UO_36 (O_36,N_9028,N_9434);
and UO_37 (O_37,N_9692,N_9454);
or UO_38 (O_38,N_9878,N_9485);
or UO_39 (O_39,N_9437,N_9414);
nand UO_40 (O_40,N_9514,N_9475);
nand UO_41 (O_41,N_9551,N_9871);
nand UO_42 (O_42,N_9887,N_9776);
and UO_43 (O_43,N_9506,N_9883);
and UO_44 (O_44,N_9242,N_9756);
or UO_45 (O_45,N_9009,N_9044);
nand UO_46 (O_46,N_9574,N_9622);
nand UO_47 (O_47,N_9059,N_9314);
or UO_48 (O_48,N_9682,N_9877);
and UO_49 (O_49,N_9341,N_9166);
or UO_50 (O_50,N_9094,N_9103);
nor UO_51 (O_51,N_9905,N_9449);
nor UO_52 (O_52,N_9231,N_9396);
and UO_53 (O_53,N_9081,N_9627);
nand UO_54 (O_54,N_9272,N_9968);
and UO_55 (O_55,N_9952,N_9438);
or UO_56 (O_56,N_9380,N_9662);
nand UO_57 (O_57,N_9697,N_9199);
nor UO_58 (O_58,N_9904,N_9355);
xor UO_59 (O_59,N_9063,N_9530);
or UO_60 (O_60,N_9943,N_9171);
xnor UO_61 (O_61,N_9385,N_9788);
and UO_62 (O_62,N_9860,N_9169);
and UO_63 (O_63,N_9580,N_9656);
and UO_64 (O_64,N_9099,N_9609);
nand UO_65 (O_65,N_9160,N_9175);
nand UO_66 (O_66,N_9838,N_9586);
nor UO_67 (O_67,N_9433,N_9445);
or UO_68 (O_68,N_9415,N_9113);
nand UO_69 (O_69,N_9538,N_9229);
nor UO_70 (O_70,N_9830,N_9631);
and UO_71 (O_71,N_9687,N_9819);
and UO_72 (O_72,N_9779,N_9616);
nand UO_73 (O_73,N_9089,N_9397);
or UO_74 (O_74,N_9601,N_9016);
nor UO_75 (O_75,N_9352,N_9273);
nand UO_76 (O_76,N_9889,N_9398);
or UO_77 (O_77,N_9865,N_9178);
nor UO_78 (O_78,N_9177,N_9549);
nand UO_79 (O_79,N_9222,N_9769);
or UO_80 (O_80,N_9712,N_9739);
nor UO_81 (O_81,N_9466,N_9306);
and UO_82 (O_82,N_9996,N_9026);
and UO_83 (O_83,N_9154,N_9218);
or UO_84 (O_84,N_9948,N_9277);
nor UO_85 (O_85,N_9181,N_9679);
nor UO_86 (O_86,N_9164,N_9092);
or UO_87 (O_87,N_9363,N_9072);
xnor UO_88 (O_88,N_9258,N_9471);
xnor UO_89 (O_89,N_9076,N_9095);
nor UO_90 (O_90,N_9815,N_9468);
and UO_91 (O_91,N_9321,N_9215);
or UO_92 (O_92,N_9288,N_9949);
and UO_93 (O_93,N_9536,N_9035);
xnor UO_94 (O_94,N_9375,N_9040);
xor UO_95 (O_95,N_9357,N_9835);
and UO_96 (O_96,N_9490,N_9304);
xnor UO_97 (O_97,N_9988,N_9209);
nand UO_98 (O_98,N_9309,N_9358);
nor UO_99 (O_99,N_9208,N_9736);
or UO_100 (O_100,N_9722,N_9900);
nor UO_101 (O_101,N_9192,N_9527);
or UO_102 (O_102,N_9322,N_9771);
nand UO_103 (O_103,N_9960,N_9684);
or UO_104 (O_104,N_9421,N_9402);
nand UO_105 (O_105,N_9390,N_9796);
or UO_106 (O_106,N_9271,N_9732);
or UO_107 (O_107,N_9578,N_9180);
and UO_108 (O_108,N_9023,N_9470);
or UO_109 (O_109,N_9100,N_9070);
or UO_110 (O_110,N_9685,N_9108);
nor UO_111 (O_111,N_9136,N_9150);
nand UO_112 (O_112,N_9486,N_9173);
nand UO_113 (O_113,N_9084,N_9686);
and UO_114 (O_114,N_9840,N_9650);
and UO_115 (O_115,N_9128,N_9014);
xor UO_116 (O_116,N_9579,N_9954);
xnor UO_117 (O_117,N_9747,N_9512);
nand UO_118 (O_118,N_9800,N_9236);
and UO_119 (O_119,N_9046,N_9864);
and UO_120 (O_120,N_9104,N_9391);
and UO_121 (O_121,N_9246,N_9316);
nand UO_122 (O_122,N_9690,N_9899);
xnor UO_123 (O_123,N_9383,N_9412);
xor UO_124 (O_124,N_9621,N_9978);
nor UO_125 (O_125,N_9921,N_9648);
xnor UO_126 (O_126,N_9153,N_9633);
or UO_127 (O_127,N_9351,N_9214);
nor UO_128 (O_128,N_9221,N_9327);
nor UO_129 (O_129,N_9786,N_9759);
nor UO_130 (O_130,N_9561,N_9976);
nand UO_131 (O_131,N_9731,N_9430);
and UO_132 (O_132,N_9927,N_9834);
nand UO_133 (O_133,N_9303,N_9553);
nor UO_134 (O_134,N_9587,N_9854);
nand UO_135 (O_135,N_9720,N_9179);
and UO_136 (O_136,N_9073,N_9989);
nor UO_137 (O_137,N_9733,N_9255);
nand UO_138 (O_138,N_9754,N_9879);
nand UO_139 (O_139,N_9301,N_9291);
nand UO_140 (O_140,N_9593,N_9090);
nand UO_141 (O_141,N_9155,N_9802);
and UO_142 (O_142,N_9265,N_9945);
xor UO_143 (O_143,N_9822,N_9852);
and UO_144 (O_144,N_9596,N_9052);
or UO_145 (O_145,N_9110,N_9312);
nand UO_146 (O_146,N_9426,N_9264);
nand UO_147 (O_147,N_9888,N_9183);
nor UO_148 (O_148,N_9443,N_9489);
or UO_149 (O_149,N_9957,N_9472);
nor UO_150 (O_150,N_9983,N_9406);
or UO_151 (O_151,N_9290,N_9121);
or UO_152 (O_152,N_9504,N_9268);
nor UO_153 (O_153,N_9620,N_9047);
and UO_154 (O_154,N_9962,N_9330);
xor UO_155 (O_155,N_9233,N_9342);
and UO_156 (O_156,N_9152,N_9567);
nand UO_157 (O_157,N_9575,N_9400);
or UO_158 (O_158,N_9311,N_9666);
nand UO_159 (O_159,N_9710,N_9995);
or UO_160 (O_160,N_9262,N_9432);
xor UO_161 (O_161,N_9148,N_9022);
xor UO_162 (O_162,N_9672,N_9683);
xnor UO_163 (O_163,N_9033,N_9938);
and UO_164 (O_164,N_9045,N_9523);
and UO_165 (O_165,N_9757,N_9528);
or UO_166 (O_166,N_9477,N_9058);
or UO_167 (O_167,N_9785,N_9381);
nand UO_168 (O_168,N_9250,N_9420);
xnor UO_169 (O_169,N_9869,N_9839);
or UO_170 (O_170,N_9409,N_9547);
xor UO_171 (O_171,N_9135,N_9071);
xor UO_172 (O_172,N_9207,N_9275);
nand UO_173 (O_173,N_9501,N_9808);
xor UO_174 (O_174,N_9370,N_9663);
nor UO_175 (O_175,N_9156,N_9168);
nor UO_176 (O_176,N_9297,N_9917);
nand UO_177 (O_177,N_9941,N_9555);
xor UO_178 (O_178,N_9185,N_9787);
nand UO_179 (O_179,N_9726,N_9661);
nor UO_180 (O_180,N_9362,N_9919);
nand UO_181 (O_181,N_9678,N_9918);
xnor UO_182 (O_182,N_9818,N_9308);
xnor UO_183 (O_183,N_9767,N_9816);
xor UO_184 (O_184,N_9737,N_9143);
xnor UO_185 (O_185,N_9098,N_9162);
nand UO_186 (O_186,N_9734,N_9556);
nand UO_187 (O_187,N_9323,N_9797);
and UO_188 (O_188,N_9429,N_9660);
nand UO_189 (O_189,N_9243,N_9458);
nor UO_190 (O_190,N_9670,N_9866);
xor UO_191 (O_191,N_9760,N_9752);
xnor UO_192 (O_192,N_9345,N_9324);
nand UO_193 (O_193,N_9077,N_9654);
xor UO_194 (O_194,N_9427,N_9335);
nand UO_195 (O_195,N_9846,N_9457);
nor UO_196 (O_196,N_9467,N_9120);
or UO_197 (O_197,N_9951,N_9749);
xnor UO_198 (O_198,N_9936,N_9038);
or UO_199 (O_199,N_9955,N_9086);
nor UO_200 (O_200,N_9619,N_9149);
or UO_201 (O_201,N_9425,N_9542);
nand UO_202 (O_202,N_9003,N_9163);
or UO_203 (O_203,N_9051,N_9346);
xnor UO_204 (O_204,N_9701,N_9758);
nor UO_205 (O_205,N_9134,N_9336);
or UO_206 (O_206,N_9407,N_9144);
or UO_207 (O_207,N_9891,N_9975);
and UO_208 (O_208,N_9903,N_9966);
nand UO_209 (O_209,N_9484,N_9172);
nor UO_210 (O_210,N_9001,N_9704);
or UO_211 (O_211,N_9768,N_9354);
nor UO_212 (O_212,N_9789,N_9010);
and UO_213 (O_213,N_9245,N_9244);
and UO_214 (O_214,N_9651,N_9576);
xor UO_215 (O_215,N_9302,N_9392);
and UO_216 (O_216,N_9206,N_9497);
and UO_217 (O_217,N_9102,N_9266);
xor UO_218 (O_218,N_9285,N_9890);
or UO_219 (O_219,N_9859,N_9982);
nand UO_220 (O_220,N_9333,N_9805);
nand UO_221 (O_221,N_9278,N_9069);
and UO_222 (O_222,N_9248,N_9435);
nor UO_223 (O_223,N_9807,N_9940);
xor UO_224 (O_224,N_9640,N_9826);
and UO_225 (O_225,N_9524,N_9002);
xnor UO_226 (O_226,N_9465,N_9934);
nand UO_227 (O_227,N_9519,N_9500);
nand UO_228 (O_228,N_9617,N_9447);
xor UO_229 (O_229,N_9196,N_9958);
xnor UO_230 (O_230,N_9770,N_9850);
and UO_231 (O_231,N_9085,N_9034);
nor UO_232 (O_232,N_9111,N_9612);
nor UO_233 (O_233,N_9118,N_9992);
xor UO_234 (O_234,N_9188,N_9766);
xnor UO_235 (O_235,N_9933,N_9801);
and UO_236 (O_236,N_9863,N_9446);
xnor UO_237 (O_237,N_9823,N_9703);
nor UO_238 (O_238,N_9334,N_9115);
nand UO_239 (O_239,N_9965,N_9295);
nor UO_240 (O_240,N_9743,N_9283);
nor UO_241 (O_241,N_9591,N_9928);
nor UO_242 (O_242,N_9774,N_9473);
nand UO_243 (O_243,N_9773,N_9371);
or UO_244 (O_244,N_9444,N_9386);
nor UO_245 (O_245,N_9376,N_9083);
and UO_246 (O_246,N_9105,N_9986);
nor UO_247 (O_247,N_9219,N_9378);
xor UO_248 (O_248,N_9509,N_9442);
and UO_249 (O_249,N_9963,N_9521);
nor UO_250 (O_250,N_9117,N_9597);
nor UO_251 (O_251,N_9119,N_9483);
nand UO_252 (O_252,N_9013,N_9939);
xnor UO_253 (O_253,N_9915,N_9583);
or UO_254 (O_254,N_9723,N_9459);
xnor UO_255 (O_255,N_9671,N_9474);
xnor UO_256 (O_256,N_9745,N_9132);
xnor UO_257 (O_257,N_9831,N_9270);
and UO_258 (O_258,N_9924,N_9698);
nor UO_259 (O_259,N_9061,N_9006);
xor UO_260 (O_260,N_9836,N_9418);
nor UO_261 (O_261,N_9062,N_9653);
nand UO_262 (O_262,N_9318,N_9636);
nand UO_263 (O_263,N_9643,N_9618);
nor UO_264 (O_264,N_9189,N_9510);
xor UO_265 (O_265,N_9505,N_9867);
and UO_266 (O_266,N_9541,N_9293);
nor UO_267 (O_267,N_9037,N_9008);
xnor UO_268 (O_268,N_9861,N_9298);
nand UO_269 (O_269,N_9885,N_9259);
or UO_270 (O_270,N_9204,N_9015);
and UO_271 (O_271,N_9646,N_9706);
xor UO_272 (O_272,N_9582,N_9570);
or UO_273 (O_273,N_9315,N_9937);
xor UO_274 (O_274,N_9049,N_9526);
or UO_275 (O_275,N_9267,N_9916);
nor UO_276 (O_276,N_9507,N_9953);
nor UO_277 (O_277,N_9605,N_9408);
xor UO_278 (O_278,N_9170,N_9495);
nand UO_279 (O_279,N_9018,N_9431);
nand UO_280 (O_280,N_9844,N_9050);
nor UO_281 (O_281,N_9223,N_9211);
nand UO_282 (O_282,N_9848,N_9738);
and UO_283 (O_283,N_9730,N_9423);
or UO_284 (O_284,N_9453,N_9320);
nor UO_285 (O_285,N_9987,N_9101);
xnor UO_286 (O_286,N_9907,N_9969);
xor UO_287 (O_287,N_9599,N_9803);
nand UO_288 (O_288,N_9491,N_9659);
and UO_289 (O_289,N_9534,N_9959);
nand UO_290 (O_290,N_9263,N_9498);
nand UO_291 (O_291,N_9515,N_9652);
or UO_292 (O_292,N_9884,N_9325);
nand UO_293 (O_293,N_9048,N_9213);
nand UO_294 (O_294,N_9724,N_9571);
or UO_295 (O_295,N_9299,N_9598);
and UO_296 (O_296,N_9344,N_9901);
or UO_297 (O_297,N_9623,N_9870);
nor UO_298 (O_298,N_9590,N_9332);
or UO_299 (O_299,N_9482,N_9716);
or UO_300 (O_300,N_9632,N_9508);
or UO_301 (O_301,N_9935,N_9820);
or UO_302 (O_302,N_9020,N_9696);
nand UO_303 (O_303,N_9481,N_9727);
and UO_304 (O_304,N_9190,N_9748);
xor UO_305 (O_305,N_9125,N_9130);
nand UO_306 (O_306,N_9565,N_9212);
and UO_307 (O_307,N_9030,N_9795);
xor UO_308 (O_308,N_9602,N_9326);
xnor UO_309 (O_309,N_9289,N_9133);
nand UO_310 (O_310,N_9395,N_9405);
nor UO_311 (O_311,N_9140,N_9416);
nor UO_312 (O_312,N_9343,N_9637);
xnor UO_313 (O_313,N_9399,N_9630);
and UO_314 (O_314,N_9544,N_9012);
nor UO_315 (O_315,N_9281,N_9305);
or UO_316 (O_316,N_9106,N_9804);
xnor UO_317 (O_317,N_9261,N_9564);
xor UO_318 (O_318,N_9488,N_9990);
nand UO_319 (O_319,N_9107,N_9588);
nor UO_320 (O_320,N_9060,N_9568);
nor UO_321 (O_321,N_9592,N_9753);
nand UO_322 (O_322,N_9127,N_9634);
nand UO_323 (O_323,N_9019,N_9589);
nand UO_324 (O_324,N_9853,N_9451);
xnor UO_325 (O_325,N_9360,N_9200);
nor UO_326 (O_326,N_9984,N_9087);
nand UO_327 (O_327,N_9658,N_9142);
xor UO_328 (O_328,N_9893,N_9053);
and UO_329 (O_329,N_9735,N_9476);
and UO_330 (O_330,N_9292,N_9313);
and UO_331 (O_331,N_9361,N_9635);
nand UO_332 (O_332,N_9922,N_9751);
nand UO_333 (O_333,N_9857,N_9639);
xor UO_334 (O_334,N_9902,N_9041);
nand UO_335 (O_335,N_9296,N_9210);
and UO_336 (O_336,N_9469,N_9765);
xnor UO_337 (O_337,N_9310,N_9694);
xor UO_338 (O_338,N_9991,N_9202);
and UO_339 (O_339,N_9525,N_9401);
or UO_340 (O_340,N_9145,N_9876);
and UO_341 (O_341,N_9174,N_9367);
and UO_342 (O_342,N_9056,N_9338);
nand UO_343 (O_343,N_9980,N_9886);
or UO_344 (O_344,N_9728,N_9974);
nor UO_345 (O_345,N_9755,N_9827);
nor UO_346 (O_346,N_9404,N_9715);
nand UO_347 (O_347,N_9424,N_9999);
and UO_348 (O_348,N_9097,N_9906);
nor UO_349 (O_349,N_9131,N_9455);
or UO_350 (O_350,N_9224,N_9543);
xor UO_351 (O_351,N_9610,N_9998);
nor UO_352 (O_352,N_9764,N_9708);
xor UO_353 (O_353,N_9719,N_9926);
nand UO_354 (O_354,N_9146,N_9141);
or UO_355 (O_355,N_9828,N_9868);
xnor UO_356 (O_356,N_9778,N_9328);
and UO_357 (O_357,N_9783,N_9535);
xor UO_358 (O_358,N_9282,N_9895);
and UO_359 (O_359,N_9930,N_9811);
nor UO_360 (O_360,N_9742,N_9116);
nand UO_361 (O_361,N_9970,N_9065);
and UO_362 (O_362,N_9994,N_9039);
xnor UO_363 (O_363,N_9036,N_9088);
and UO_364 (O_364,N_9329,N_9516);
and UO_365 (O_365,N_9882,N_9856);
or UO_366 (O_366,N_9122,N_9337);
or UO_367 (O_367,N_9379,N_9096);
nor UO_368 (O_368,N_9159,N_9456);
nand UO_369 (O_369,N_9460,N_9480);
nand UO_370 (O_370,N_9387,N_9810);
or UO_371 (O_371,N_9027,N_9910);
or UO_372 (O_372,N_9920,N_9566);
xnor UO_373 (O_373,N_9366,N_9641);
or UO_374 (O_374,N_9545,N_9608);
nand UO_375 (O_375,N_9806,N_9675);
and UO_376 (O_376,N_9809,N_9985);
nor UO_377 (O_377,N_9531,N_9411);
xor UO_378 (O_378,N_9862,N_9031);
nand UO_379 (O_379,N_9972,N_9585);
or UO_380 (O_380,N_9167,N_9522);
nand UO_381 (O_381,N_9821,N_9624);
xor UO_382 (O_382,N_9664,N_9912);
nand UO_383 (O_383,N_9956,N_9950);
and UO_384 (O_384,N_9503,N_9559);
xor UO_385 (O_385,N_9908,N_9064);
nor UO_386 (O_386,N_9611,N_9638);
xor UO_387 (O_387,N_9439,N_9317);
xnor UO_388 (O_388,N_9237,N_9613);
nor UO_389 (O_389,N_9817,N_9126);
nand UO_390 (O_390,N_9011,N_9082);
xnor UO_391 (O_391,N_9091,N_9410);
or UO_392 (O_392,N_9286,N_9394);
and UO_393 (O_393,N_9005,N_9721);
or UO_394 (O_394,N_9763,N_9225);
xnor UO_395 (O_395,N_9713,N_9252);
nand UO_396 (O_396,N_9257,N_9832);
or UO_397 (O_397,N_9674,N_9881);
and UO_398 (O_398,N_9929,N_9824);
nor UO_399 (O_399,N_9669,N_9203);
or UO_400 (O_400,N_9191,N_9665);
nor UO_401 (O_401,N_9198,N_9024);
nand UO_402 (O_402,N_9021,N_9550);
and UO_403 (O_403,N_9825,N_9781);
and UO_404 (O_404,N_9269,N_9403);
nand UO_405 (O_405,N_9532,N_9043);
nor UO_406 (O_406,N_9017,N_9746);
and UO_407 (O_407,N_9772,N_9388);
or UO_408 (O_408,N_9762,N_9799);
or UO_409 (O_409,N_9230,N_9777);
nor UO_410 (O_410,N_9782,N_9812);
nor UO_411 (O_411,N_9829,N_9780);
and UO_412 (O_412,N_9382,N_9093);
xor UO_413 (O_413,N_9184,N_9695);
xor UO_414 (O_414,N_9725,N_9655);
xor UO_415 (O_415,N_9353,N_9798);
or UO_416 (O_416,N_9699,N_9274);
nand UO_417 (O_417,N_9463,N_9581);
or UO_418 (O_418,N_9793,N_9539);
xor UO_419 (O_419,N_9461,N_9702);
nand UO_420 (O_420,N_9932,N_9186);
xnor UO_421 (O_421,N_9339,N_9109);
nor UO_422 (O_422,N_9744,N_9247);
or UO_423 (O_423,N_9165,N_9450);
or UO_424 (O_424,N_9436,N_9161);
xnor UO_425 (O_425,N_9374,N_9964);
or UO_426 (O_426,N_9792,N_9718);
xor UO_427 (O_427,N_9858,N_9452);
nand UO_428 (O_428,N_9775,N_9193);
or UO_429 (O_429,N_9158,N_9139);
or UO_430 (O_430,N_9372,N_9573);
xor UO_431 (O_431,N_9843,N_9276);
nand UO_432 (O_432,N_9228,N_9518);
or UO_433 (O_433,N_9493,N_9997);
or UO_434 (O_434,N_9606,N_9709);
and UO_435 (O_435,N_9078,N_9157);
and UO_436 (O_436,N_9359,N_9241);
xnor UO_437 (O_437,N_9689,N_9552);
nor UO_438 (O_438,N_9700,N_9300);
nand UO_439 (O_439,N_9112,N_9075);
and UO_440 (O_440,N_9614,N_9849);
nand UO_441 (O_441,N_9260,N_9971);
or UO_442 (O_442,N_9287,N_9147);
nor UO_443 (O_443,N_9499,N_9741);
nor UO_444 (O_444,N_9626,N_9238);
or UO_445 (O_445,N_9714,N_9413);
or UO_446 (O_446,N_9707,N_9419);
or UO_447 (O_447,N_9546,N_9711);
and UO_448 (O_448,N_9548,N_9068);
or UO_449 (O_449,N_9347,N_9007);
nor UO_450 (O_450,N_9604,N_9253);
nand UO_451 (O_451,N_9029,N_9892);
xor UO_452 (O_452,N_9946,N_9560);
nor UO_453 (O_453,N_9331,N_9645);
nor UO_454 (O_454,N_9761,N_9513);
nand UO_455 (O_455,N_9603,N_9057);
or UO_456 (O_456,N_9067,N_9649);
nand UO_457 (O_457,N_9607,N_9205);
or UO_458 (O_458,N_9677,N_9079);
xnor UO_459 (O_459,N_9647,N_9691);
nand UO_460 (O_460,N_9563,N_9977);
nor UO_461 (O_461,N_9673,N_9422);
xnor UO_462 (O_462,N_9729,N_9365);
nand UO_463 (O_463,N_9914,N_9494);
and UO_464 (O_464,N_9740,N_9393);
nand UO_465 (O_465,N_9880,N_9348);
or UO_466 (O_466,N_9138,N_9000);
xor UO_467 (O_467,N_9441,N_9845);
xor UO_468 (O_468,N_9529,N_9872);
nand UO_469 (O_469,N_9216,N_9814);
and UO_470 (O_470,N_9054,N_9197);
and UO_471 (O_471,N_9842,N_9595);
and UO_472 (O_472,N_9220,N_9794);
xor UO_473 (O_473,N_9562,N_9875);
xor UO_474 (O_474,N_9448,N_9791);
xor UO_475 (O_475,N_9644,N_9979);
or UO_476 (O_476,N_9151,N_9537);
xnor UO_477 (O_477,N_9176,N_9961);
xor UO_478 (O_478,N_9841,N_9217);
nor UO_479 (O_479,N_9554,N_9124);
nor UO_480 (O_480,N_9717,N_9232);
xor UO_481 (O_481,N_9307,N_9074);
nor UO_482 (O_482,N_9187,N_9833);
or UO_483 (O_483,N_9350,N_9256);
nor UO_484 (O_484,N_9364,N_9194);
or UO_485 (O_485,N_9280,N_9234);
or UO_486 (O_486,N_9993,N_9129);
or UO_487 (O_487,N_9319,N_9239);
xnor UO_488 (O_488,N_9911,N_9944);
xnor UO_489 (O_489,N_9750,N_9981);
and UO_490 (O_490,N_9894,N_9520);
and UO_491 (O_491,N_9004,N_9055);
nand UO_492 (O_492,N_9249,N_9251);
nor UO_493 (O_493,N_9558,N_9973);
and UO_494 (O_494,N_9657,N_9874);
xnor UO_495 (O_495,N_9615,N_9540);
nor UO_496 (O_496,N_9557,N_9668);
xor UO_497 (O_497,N_9182,N_9967);
nand UO_498 (O_498,N_9813,N_9195);
nor UO_499 (O_499,N_9913,N_9440);
nand UO_500 (O_500,N_9327,N_9208);
nor UO_501 (O_501,N_9495,N_9684);
nand UO_502 (O_502,N_9528,N_9202);
xor UO_503 (O_503,N_9625,N_9437);
nand UO_504 (O_504,N_9312,N_9186);
xor UO_505 (O_505,N_9468,N_9391);
xor UO_506 (O_506,N_9413,N_9040);
nand UO_507 (O_507,N_9210,N_9287);
or UO_508 (O_508,N_9966,N_9988);
and UO_509 (O_509,N_9580,N_9261);
nor UO_510 (O_510,N_9477,N_9965);
and UO_511 (O_511,N_9069,N_9610);
or UO_512 (O_512,N_9940,N_9372);
and UO_513 (O_513,N_9250,N_9660);
xnor UO_514 (O_514,N_9120,N_9794);
and UO_515 (O_515,N_9716,N_9352);
and UO_516 (O_516,N_9369,N_9079);
xor UO_517 (O_517,N_9396,N_9513);
nor UO_518 (O_518,N_9565,N_9460);
or UO_519 (O_519,N_9203,N_9277);
xnor UO_520 (O_520,N_9178,N_9770);
nor UO_521 (O_521,N_9886,N_9293);
nor UO_522 (O_522,N_9774,N_9534);
nand UO_523 (O_523,N_9552,N_9193);
xor UO_524 (O_524,N_9265,N_9546);
xnor UO_525 (O_525,N_9615,N_9277);
or UO_526 (O_526,N_9055,N_9627);
and UO_527 (O_527,N_9615,N_9196);
xnor UO_528 (O_528,N_9487,N_9958);
or UO_529 (O_529,N_9033,N_9613);
or UO_530 (O_530,N_9028,N_9659);
nand UO_531 (O_531,N_9299,N_9293);
and UO_532 (O_532,N_9556,N_9385);
nor UO_533 (O_533,N_9536,N_9465);
nor UO_534 (O_534,N_9043,N_9966);
nand UO_535 (O_535,N_9103,N_9397);
nand UO_536 (O_536,N_9023,N_9797);
nor UO_537 (O_537,N_9144,N_9722);
nor UO_538 (O_538,N_9674,N_9811);
and UO_539 (O_539,N_9612,N_9038);
nand UO_540 (O_540,N_9538,N_9287);
or UO_541 (O_541,N_9436,N_9167);
nor UO_542 (O_542,N_9090,N_9216);
nor UO_543 (O_543,N_9340,N_9320);
and UO_544 (O_544,N_9138,N_9208);
or UO_545 (O_545,N_9473,N_9695);
and UO_546 (O_546,N_9220,N_9621);
nand UO_547 (O_547,N_9359,N_9580);
nor UO_548 (O_548,N_9033,N_9312);
xor UO_549 (O_549,N_9415,N_9676);
nor UO_550 (O_550,N_9399,N_9109);
nor UO_551 (O_551,N_9628,N_9059);
nor UO_552 (O_552,N_9987,N_9440);
and UO_553 (O_553,N_9905,N_9137);
nor UO_554 (O_554,N_9111,N_9726);
xnor UO_555 (O_555,N_9911,N_9406);
and UO_556 (O_556,N_9280,N_9037);
or UO_557 (O_557,N_9050,N_9235);
xor UO_558 (O_558,N_9388,N_9773);
and UO_559 (O_559,N_9238,N_9897);
nand UO_560 (O_560,N_9137,N_9160);
nand UO_561 (O_561,N_9411,N_9135);
or UO_562 (O_562,N_9980,N_9101);
and UO_563 (O_563,N_9909,N_9336);
nor UO_564 (O_564,N_9634,N_9946);
nand UO_565 (O_565,N_9841,N_9828);
nor UO_566 (O_566,N_9331,N_9235);
or UO_567 (O_567,N_9581,N_9982);
nand UO_568 (O_568,N_9525,N_9509);
and UO_569 (O_569,N_9065,N_9837);
xor UO_570 (O_570,N_9267,N_9962);
or UO_571 (O_571,N_9512,N_9493);
nor UO_572 (O_572,N_9833,N_9368);
nand UO_573 (O_573,N_9855,N_9220);
nor UO_574 (O_574,N_9317,N_9035);
and UO_575 (O_575,N_9844,N_9129);
nand UO_576 (O_576,N_9809,N_9422);
and UO_577 (O_577,N_9943,N_9572);
or UO_578 (O_578,N_9912,N_9310);
and UO_579 (O_579,N_9028,N_9934);
or UO_580 (O_580,N_9332,N_9367);
nand UO_581 (O_581,N_9118,N_9622);
and UO_582 (O_582,N_9084,N_9239);
xnor UO_583 (O_583,N_9876,N_9831);
xnor UO_584 (O_584,N_9167,N_9570);
and UO_585 (O_585,N_9862,N_9850);
nor UO_586 (O_586,N_9618,N_9492);
or UO_587 (O_587,N_9132,N_9185);
xor UO_588 (O_588,N_9846,N_9638);
xnor UO_589 (O_589,N_9218,N_9852);
or UO_590 (O_590,N_9877,N_9519);
and UO_591 (O_591,N_9173,N_9382);
nor UO_592 (O_592,N_9379,N_9090);
nor UO_593 (O_593,N_9785,N_9837);
and UO_594 (O_594,N_9234,N_9798);
nor UO_595 (O_595,N_9205,N_9389);
and UO_596 (O_596,N_9174,N_9754);
xor UO_597 (O_597,N_9666,N_9523);
and UO_598 (O_598,N_9153,N_9532);
xor UO_599 (O_599,N_9138,N_9658);
xnor UO_600 (O_600,N_9976,N_9403);
xnor UO_601 (O_601,N_9389,N_9959);
xnor UO_602 (O_602,N_9588,N_9780);
or UO_603 (O_603,N_9185,N_9785);
nand UO_604 (O_604,N_9097,N_9627);
nor UO_605 (O_605,N_9178,N_9986);
nand UO_606 (O_606,N_9259,N_9219);
and UO_607 (O_607,N_9743,N_9060);
nor UO_608 (O_608,N_9221,N_9697);
and UO_609 (O_609,N_9120,N_9612);
xnor UO_610 (O_610,N_9737,N_9847);
or UO_611 (O_611,N_9964,N_9824);
xnor UO_612 (O_612,N_9776,N_9615);
nand UO_613 (O_613,N_9940,N_9850);
xnor UO_614 (O_614,N_9351,N_9456);
and UO_615 (O_615,N_9512,N_9592);
and UO_616 (O_616,N_9334,N_9058);
xor UO_617 (O_617,N_9149,N_9207);
and UO_618 (O_618,N_9576,N_9783);
nand UO_619 (O_619,N_9849,N_9312);
nand UO_620 (O_620,N_9058,N_9039);
nand UO_621 (O_621,N_9131,N_9512);
xor UO_622 (O_622,N_9852,N_9467);
xor UO_623 (O_623,N_9147,N_9553);
xnor UO_624 (O_624,N_9930,N_9628);
xnor UO_625 (O_625,N_9556,N_9031);
xor UO_626 (O_626,N_9220,N_9491);
or UO_627 (O_627,N_9009,N_9317);
nor UO_628 (O_628,N_9097,N_9851);
nor UO_629 (O_629,N_9403,N_9539);
or UO_630 (O_630,N_9336,N_9804);
nand UO_631 (O_631,N_9335,N_9947);
nand UO_632 (O_632,N_9862,N_9707);
or UO_633 (O_633,N_9205,N_9070);
xnor UO_634 (O_634,N_9944,N_9662);
nor UO_635 (O_635,N_9570,N_9987);
and UO_636 (O_636,N_9133,N_9135);
nand UO_637 (O_637,N_9548,N_9681);
and UO_638 (O_638,N_9562,N_9063);
or UO_639 (O_639,N_9121,N_9636);
xnor UO_640 (O_640,N_9742,N_9944);
xnor UO_641 (O_641,N_9114,N_9680);
xnor UO_642 (O_642,N_9943,N_9420);
and UO_643 (O_643,N_9719,N_9097);
xor UO_644 (O_644,N_9249,N_9648);
or UO_645 (O_645,N_9222,N_9069);
nand UO_646 (O_646,N_9271,N_9141);
nand UO_647 (O_647,N_9379,N_9659);
nand UO_648 (O_648,N_9382,N_9790);
xor UO_649 (O_649,N_9227,N_9094);
or UO_650 (O_650,N_9161,N_9916);
xnor UO_651 (O_651,N_9767,N_9789);
or UO_652 (O_652,N_9588,N_9989);
nand UO_653 (O_653,N_9328,N_9133);
xnor UO_654 (O_654,N_9397,N_9892);
and UO_655 (O_655,N_9278,N_9275);
xor UO_656 (O_656,N_9208,N_9977);
nand UO_657 (O_657,N_9203,N_9940);
and UO_658 (O_658,N_9327,N_9748);
nor UO_659 (O_659,N_9554,N_9939);
and UO_660 (O_660,N_9606,N_9273);
nand UO_661 (O_661,N_9418,N_9119);
xnor UO_662 (O_662,N_9674,N_9831);
xnor UO_663 (O_663,N_9740,N_9706);
xor UO_664 (O_664,N_9960,N_9319);
nor UO_665 (O_665,N_9005,N_9088);
or UO_666 (O_666,N_9246,N_9414);
and UO_667 (O_667,N_9952,N_9786);
xor UO_668 (O_668,N_9108,N_9079);
nand UO_669 (O_669,N_9226,N_9315);
nor UO_670 (O_670,N_9036,N_9849);
nand UO_671 (O_671,N_9434,N_9441);
and UO_672 (O_672,N_9586,N_9548);
nor UO_673 (O_673,N_9508,N_9763);
nor UO_674 (O_674,N_9684,N_9189);
or UO_675 (O_675,N_9519,N_9757);
nand UO_676 (O_676,N_9197,N_9521);
nor UO_677 (O_677,N_9974,N_9679);
nor UO_678 (O_678,N_9430,N_9059);
and UO_679 (O_679,N_9232,N_9595);
nor UO_680 (O_680,N_9044,N_9807);
nand UO_681 (O_681,N_9580,N_9236);
and UO_682 (O_682,N_9098,N_9317);
and UO_683 (O_683,N_9145,N_9255);
nand UO_684 (O_684,N_9134,N_9564);
and UO_685 (O_685,N_9039,N_9367);
xnor UO_686 (O_686,N_9594,N_9982);
nor UO_687 (O_687,N_9048,N_9026);
nand UO_688 (O_688,N_9818,N_9341);
nand UO_689 (O_689,N_9350,N_9769);
nand UO_690 (O_690,N_9175,N_9580);
nand UO_691 (O_691,N_9670,N_9749);
or UO_692 (O_692,N_9095,N_9975);
nor UO_693 (O_693,N_9091,N_9774);
and UO_694 (O_694,N_9955,N_9981);
or UO_695 (O_695,N_9683,N_9453);
nor UO_696 (O_696,N_9068,N_9264);
or UO_697 (O_697,N_9518,N_9366);
nand UO_698 (O_698,N_9402,N_9891);
or UO_699 (O_699,N_9390,N_9244);
xnor UO_700 (O_700,N_9370,N_9493);
xnor UO_701 (O_701,N_9021,N_9007);
xor UO_702 (O_702,N_9626,N_9255);
nor UO_703 (O_703,N_9977,N_9690);
and UO_704 (O_704,N_9723,N_9533);
xnor UO_705 (O_705,N_9792,N_9952);
nor UO_706 (O_706,N_9030,N_9483);
or UO_707 (O_707,N_9434,N_9989);
nand UO_708 (O_708,N_9156,N_9487);
and UO_709 (O_709,N_9777,N_9757);
and UO_710 (O_710,N_9605,N_9455);
and UO_711 (O_711,N_9948,N_9890);
xnor UO_712 (O_712,N_9406,N_9589);
nor UO_713 (O_713,N_9802,N_9977);
xnor UO_714 (O_714,N_9207,N_9028);
nor UO_715 (O_715,N_9195,N_9081);
nor UO_716 (O_716,N_9962,N_9802);
nand UO_717 (O_717,N_9446,N_9519);
xnor UO_718 (O_718,N_9531,N_9309);
or UO_719 (O_719,N_9581,N_9673);
nand UO_720 (O_720,N_9277,N_9911);
or UO_721 (O_721,N_9086,N_9456);
nand UO_722 (O_722,N_9724,N_9179);
nand UO_723 (O_723,N_9318,N_9317);
nand UO_724 (O_724,N_9580,N_9267);
nor UO_725 (O_725,N_9256,N_9138);
nor UO_726 (O_726,N_9145,N_9121);
or UO_727 (O_727,N_9737,N_9695);
xnor UO_728 (O_728,N_9057,N_9351);
nor UO_729 (O_729,N_9852,N_9454);
and UO_730 (O_730,N_9932,N_9193);
xor UO_731 (O_731,N_9142,N_9537);
xnor UO_732 (O_732,N_9930,N_9354);
xor UO_733 (O_733,N_9792,N_9873);
xnor UO_734 (O_734,N_9323,N_9852);
xnor UO_735 (O_735,N_9464,N_9884);
and UO_736 (O_736,N_9715,N_9299);
xnor UO_737 (O_737,N_9084,N_9415);
nor UO_738 (O_738,N_9123,N_9349);
nand UO_739 (O_739,N_9910,N_9627);
or UO_740 (O_740,N_9411,N_9462);
nor UO_741 (O_741,N_9085,N_9197);
nand UO_742 (O_742,N_9125,N_9958);
nor UO_743 (O_743,N_9026,N_9330);
xnor UO_744 (O_744,N_9227,N_9631);
and UO_745 (O_745,N_9546,N_9164);
xor UO_746 (O_746,N_9004,N_9727);
xor UO_747 (O_747,N_9733,N_9560);
or UO_748 (O_748,N_9584,N_9078);
xnor UO_749 (O_749,N_9864,N_9967);
or UO_750 (O_750,N_9053,N_9178);
and UO_751 (O_751,N_9570,N_9018);
xnor UO_752 (O_752,N_9657,N_9225);
nand UO_753 (O_753,N_9358,N_9544);
and UO_754 (O_754,N_9776,N_9047);
xor UO_755 (O_755,N_9302,N_9399);
or UO_756 (O_756,N_9667,N_9487);
xor UO_757 (O_757,N_9305,N_9622);
nand UO_758 (O_758,N_9541,N_9939);
xor UO_759 (O_759,N_9257,N_9925);
nor UO_760 (O_760,N_9468,N_9120);
or UO_761 (O_761,N_9534,N_9018);
nor UO_762 (O_762,N_9327,N_9949);
nand UO_763 (O_763,N_9138,N_9444);
or UO_764 (O_764,N_9529,N_9404);
xnor UO_765 (O_765,N_9281,N_9490);
nor UO_766 (O_766,N_9252,N_9439);
nand UO_767 (O_767,N_9421,N_9039);
or UO_768 (O_768,N_9800,N_9913);
nor UO_769 (O_769,N_9404,N_9898);
xor UO_770 (O_770,N_9263,N_9134);
xor UO_771 (O_771,N_9193,N_9737);
and UO_772 (O_772,N_9803,N_9109);
xor UO_773 (O_773,N_9873,N_9434);
nor UO_774 (O_774,N_9232,N_9700);
or UO_775 (O_775,N_9958,N_9167);
nand UO_776 (O_776,N_9703,N_9965);
and UO_777 (O_777,N_9831,N_9333);
nor UO_778 (O_778,N_9225,N_9432);
and UO_779 (O_779,N_9219,N_9830);
nor UO_780 (O_780,N_9689,N_9397);
and UO_781 (O_781,N_9150,N_9558);
and UO_782 (O_782,N_9681,N_9129);
nor UO_783 (O_783,N_9691,N_9315);
or UO_784 (O_784,N_9261,N_9318);
xor UO_785 (O_785,N_9191,N_9976);
and UO_786 (O_786,N_9109,N_9048);
or UO_787 (O_787,N_9073,N_9530);
nand UO_788 (O_788,N_9370,N_9870);
nand UO_789 (O_789,N_9019,N_9521);
xnor UO_790 (O_790,N_9515,N_9167);
nand UO_791 (O_791,N_9655,N_9720);
and UO_792 (O_792,N_9754,N_9084);
nor UO_793 (O_793,N_9038,N_9650);
nor UO_794 (O_794,N_9143,N_9694);
nand UO_795 (O_795,N_9373,N_9744);
and UO_796 (O_796,N_9387,N_9978);
or UO_797 (O_797,N_9365,N_9865);
nand UO_798 (O_798,N_9492,N_9610);
nand UO_799 (O_799,N_9760,N_9078);
xnor UO_800 (O_800,N_9383,N_9965);
nand UO_801 (O_801,N_9227,N_9761);
nor UO_802 (O_802,N_9052,N_9041);
or UO_803 (O_803,N_9368,N_9463);
and UO_804 (O_804,N_9895,N_9749);
or UO_805 (O_805,N_9068,N_9289);
nand UO_806 (O_806,N_9794,N_9647);
and UO_807 (O_807,N_9973,N_9579);
nand UO_808 (O_808,N_9742,N_9227);
or UO_809 (O_809,N_9003,N_9195);
nand UO_810 (O_810,N_9288,N_9222);
or UO_811 (O_811,N_9593,N_9141);
or UO_812 (O_812,N_9000,N_9448);
or UO_813 (O_813,N_9380,N_9019);
nor UO_814 (O_814,N_9749,N_9032);
or UO_815 (O_815,N_9661,N_9753);
and UO_816 (O_816,N_9869,N_9105);
nand UO_817 (O_817,N_9553,N_9397);
xor UO_818 (O_818,N_9191,N_9529);
nor UO_819 (O_819,N_9099,N_9626);
and UO_820 (O_820,N_9494,N_9030);
and UO_821 (O_821,N_9061,N_9001);
nand UO_822 (O_822,N_9253,N_9773);
and UO_823 (O_823,N_9529,N_9003);
and UO_824 (O_824,N_9355,N_9456);
nor UO_825 (O_825,N_9031,N_9543);
nor UO_826 (O_826,N_9417,N_9280);
nor UO_827 (O_827,N_9910,N_9480);
or UO_828 (O_828,N_9708,N_9049);
nand UO_829 (O_829,N_9633,N_9109);
or UO_830 (O_830,N_9228,N_9486);
or UO_831 (O_831,N_9918,N_9751);
nand UO_832 (O_832,N_9048,N_9173);
or UO_833 (O_833,N_9279,N_9617);
nor UO_834 (O_834,N_9297,N_9921);
or UO_835 (O_835,N_9537,N_9716);
and UO_836 (O_836,N_9187,N_9626);
and UO_837 (O_837,N_9606,N_9100);
xnor UO_838 (O_838,N_9601,N_9197);
and UO_839 (O_839,N_9867,N_9606);
nor UO_840 (O_840,N_9958,N_9717);
or UO_841 (O_841,N_9634,N_9058);
xnor UO_842 (O_842,N_9340,N_9122);
nor UO_843 (O_843,N_9651,N_9050);
nand UO_844 (O_844,N_9723,N_9458);
nand UO_845 (O_845,N_9860,N_9560);
nor UO_846 (O_846,N_9657,N_9852);
or UO_847 (O_847,N_9921,N_9415);
xor UO_848 (O_848,N_9144,N_9682);
nor UO_849 (O_849,N_9742,N_9881);
and UO_850 (O_850,N_9682,N_9601);
and UO_851 (O_851,N_9242,N_9149);
nand UO_852 (O_852,N_9572,N_9115);
nand UO_853 (O_853,N_9819,N_9670);
nor UO_854 (O_854,N_9891,N_9840);
xnor UO_855 (O_855,N_9499,N_9811);
or UO_856 (O_856,N_9748,N_9375);
nor UO_857 (O_857,N_9916,N_9829);
xnor UO_858 (O_858,N_9156,N_9488);
and UO_859 (O_859,N_9639,N_9065);
xor UO_860 (O_860,N_9194,N_9252);
and UO_861 (O_861,N_9080,N_9759);
nand UO_862 (O_862,N_9314,N_9927);
or UO_863 (O_863,N_9145,N_9618);
and UO_864 (O_864,N_9252,N_9994);
nand UO_865 (O_865,N_9900,N_9329);
or UO_866 (O_866,N_9225,N_9207);
nand UO_867 (O_867,N_9672,N_9639);
nor UO_868 (O_868,N_9706,N_9992);
xnor UO_869 (O_869,N_9727,N_9500);
and UO_870 (O_870,N_9204,N_9171);
xnor UO_871 (O_871,N_9761,N_9957);
and UO_872 (O_872,N_9183,N_9730);
or UO_873 (O_873,N_9679,N_9617);
and UO_874 (O_874,N_9381,N_9430);
or UO_875 (O_875,N_9001,N_9020);
nand UO_876 (O_876,N_9784,N_9800);
and UO_877 (O_877,N_9695,N_9081);
nand UO_878 (O_878,N_9383,N_9728);
or UO_879 (O_879,N_9688,N_9350);
xor UO_880 (O_880,N_9332,N_9319);
xor UO_881 (O_881,N_9517,N_9940);
and UO_882 (O_882,N_9920,N_9736);
and UO_883 (O_883,N_9939,N_9915);
nor UO_884 (O_884,N_9631,N_9482);
nor UO_885 (O_885,N_9750,N_9949);
nor UO_886 (O_886,N_9301,N_9722);
and UO_887 (O_887,N_9477,N_9316);
and UO_888 (O_888,N_9495,N_9758);
and UO_889 (O_889,N_9592,N_9526);
xnor UO_890 (O_890,N_9618,N_9871);
nor UO_891 (O_891,N_9514,N_9932);
xnor UO_892 (O_892,N_9497,N_9929);
and UO_893 (O_893,N_9191,N_9490);
or UO_894 (O_894,N_9809,N_9322);
xor UO_895 (O_895,N_9234,N_9958);
nand UO_896 (O_896,N_9957,N_9670);
and UO_897 (O_897,N_9418,N_9867);
nor UO_898 (O_898,N_9772,N_9904);
nand UO_899 (O_899,N_9119,N_9761);
xnor UO_900 (O_900,N_9980,N_9215);
nand UO_901 (O_901,N_9562,N_9584);
and UO_902 (O_902,N_9230,N_9806);
nand UO_903 (O_903,N_9459,N_9335);
and UO_904 (O_904,N_9511,N_9136);
xor UO_905 (O_905,N_9742,N_9743);
xnor UO_906 (O_906,N_9732,N_9377);
xnor UO_907 (O_907,N_9921,N_9424);
nor UO_908 (O_908,N_9214,N_9104);
and UO_909 (O_909,N_9046,N_9212);
nor UO_910 (O_910,N_9744,N_9219);
xor UO_911 (O_911,N_9517,N_9763);
and UO_912 (O_912,N_9179,N_9661);
nor UO_913 (O_913,N_9746,N_9627);
nand UO_914 (O_914,N_9804,N_9391);
nor UO_915 (O_915,N_9563,N_9896);
nand UO_916 (O_916,N_9823,N_9661);
nor UO_917 (O_917,N_9091,N_9558);
and UO_918 (O_918,N_9398,N_9106);
or UO_919 (O_919,N_9568,N_9621);
or UO_920 (O_920,N_9039,N_9166);
xnor UO_921 (O_921,N_9464,N_9524);
nor UO_922 (O_922,N_9034,N_9227);
xor UO_923 (O_923,N_9544,N_9049);
or UO_924 (O_924,N_9879,N_9299);
nand UO_925 (O_925,N_9908,N_9344);
nand UO_926 (O_926,N_9864,N_9791);
nor UO_927 (O_927,N_9784,N_9993);
xnor UO_928 (O_928,N_9070,N_9125);
and UO_929 (O_929,N_9717,N_9246);
nand UO_930 (O_930,N_9651,N_9451);
and UO_931 (O_931,N_9598,N_9448);
or UO_932 (O_932,N_9690,N_9242);
and UO_933 (O_933,N_9642,N_9685);
nand UO_934 (O_934,N_9942,N_9582);
xnor UO_935 (O_935,N_9107,N_9776);
and UO_936 (O_936,N_9676,N_9853);
xnor UO_937 (O_937,N_9108,N_9288);
xor UO_938 (O_938,N_9607,N_9643);
nor UO_939 (O_939,N_9858,N_9422);
and UO_940 (O_940,N_9403,N_9444);
or UO_941 (O_941,N_9438,N_9296);
or UO_942 (O_942,N_9979,N_9599);
nor UO_943 (O_943,N_9838,N_9842);
xor UO_944 (O_944,N_9231,N_9624);
and UO_945 (O_945,N_9242,N_9923);
or UO_946 (O_946,N_9493,N_9750);
nor UO_947 (O_947,N_9817,N_9818);
or UO_948 (O_948,N_9761,N_9654);
and UO_949 (O_949,N_9455,N_9688);
or UO_950 (O_950,N_9735,N_9972);
nor UO_951 (O_951,N_9658,N_9424);
xnor UO_952 (O_952,N_9860,N_9437);
nand UO_953 (O_953,N_9704,N_9047);
nor UO_954 (O_954,N_9166,N_9773);
nand UO_955 (O_955,N_9014,N_9439);
and UO_956 (O_956,N_9160,N_9120);
nor UO_957 (O_957,N_9539,N_9246);
xor UO_958 (O_958,N_9713,N_9992);
and UO_959 (O_959,N_9472,N_9891);
xor UO_960 (O_960,N_9050,N_9028);
or UO_961 (O_961,N_9703,N_9260);
or UO_962 (O_962,N_9987,N_9851);
nand UO_963 (O_963,N_9879,N_9840);
nor UO_964 (O_964,N_9595,N_9169);
or UO_965 (O_965,N_9243,N_9141);
and UO_966 (O_966,N_9109,N_9912);
and UO_967 (O_967,N_9744,N_9465);
or UO_968 (O_968,N_9468,N_9295);
or UO_969 (O_969,N_9513,N_9524);
nand UO_970 (O_970,N_9851,N_9243);
nor UO_971 (O_971,N_9299,N_9247);
xnor UO_972 (O_972,N_9717,N_9345);
or UO_973 (O_973,N_9101,N_9159);
nand UO_974 (O_974,N_9671,N_9826);
xor UO_975 (O_975,N_9641,N_9829);
xnor UO_976 (O_976,N_9727,N_9884);
nand UO_977 (O_977,N_9872,N_9627);
and UO_978 (O_978,N_9483,N_9520);
and UO_979 (O_979,N_9912,N_9918);
or UO_980 (O_980,N_9180,N_9177);
and UO_981 (O_981,N_9905,N_9422);
xnor UO_982 (O_982,N_9592,N_9278);
and UO_983 (O_983,N_9277,N_9014);
nand UO_984 (O_984,N_9379,N_9835);
xor UO_985 (O_985,N_9129,N_9765);
nor UO_986 (O_986,N_9807,N_9700);
nand UO_987 (O_987,N_9367,N_9600);
and UO_988 (O_988,N_9058,N_9928);
or UO_989 (O_989,N_9250,N_9220);
xnor UO_990 (O_990,N_9385,N_9506);
xnor UO_991 (O_991,N_9506,N_9991);
and UO_992 (O_992,N_9135,N_9643);
xnor UO_993 (O_993,N_9891,N_9152);
xor UO_994 (O_994,N_9010,N_9530);
and UO_995 (O_995,N_9688,N_9273);
or UO_996 (O_996,N_9731,N_9949);
nand UO_997 (O_997,N_9487,N_9446);
nor UO_998 (O_998,N_9123,N_9644);
or UO_999 (O_999,N_9855,N_9151);
nand UO_1000 (O_1000,N_9936,N_9783);
and UO_1001 (O_1001,N_9689,N_9352);
nand UO_1002 (O_1002,N_9951,N_9803);
and UO_1003 (O_1003,N_9262,N_9332);
and UO_1004 (O_1004,N_9825,N_9506);
nor UO_1005 (O_1005,N_9449,N_9592);
or UO_1006 (O_1006,N_9424,N_9633);
and UO_1007 (O_1007,N_9231,N_9288);
xnor UO_1008 (O_1008,N_9934,N_9548);
nor UO_1009 (O_1009,N_9203,N_9663);
or UO_1010 (O_1010,N_9971,N_9261);
and UO_1011 (O_1011,N_9965,N_9458);
xor UO_1012 (O_1012,N_9886,N_9530);
or UO_1013 (O_1013,N_9487,N_9093);
and UO_1014 (O_1014,N_9751,N_9912);
nor UO_1015 (O_1015,N_9869,N_9321);
nor UO_1016 (O_1016,N_9015,N_9611);
xor UO_1017 (O_1017,N_9046,N_9568);
nor UO_1018 (O_1018,N_9473,N_9087);
xor UO_1019 (O_1019,N_9597,N_9799);
or UO_1020 (O_1020,N_9314,N_9260);
xnor UO_1021 (O_1021,N_9388,N_9254);
or UO_1022 (O_1022,N_9741,N_9073);
and UO_1023 (O_1023,N_9191,N_9174);
nand UO_1024 (O_1024,N_9128,N_9560);
xor UO_1025 (O_1025,N_9502,N_9470);
xnor UO_1026 (O_1026,N_9085,N_9577);
nand UO_1027 (O_1027,N_9045,N_9964);
and UO_1028 (O_1028,N_9468,N_9591);
or UO_1029 (O_1029,N_9487,N_9582);
xor UO_1030 (O_1030,N_9769,N_9655);
nand UO_1031 (O_1031,N_9872,N_9716);
nor UO_1032 (O_1032,N_9884,N_9491);
or UO_1033 (O_1033,N_9986,N_9963);
nor UO_1034 (O_1034,N_9203,N_9975);
and UO_1035 (O_1035,N_9806,N_9410);
xnor UO_1036 (O_1036,N_9791,N_9608);
nor UO_1037 (O_1037,N_9901,N_9426);
or UO_1038 (O_1038,N_9396,N_9027);
nand UO_1039 (O_1039,N_9129,N_9883);
and UO_1040 (O_1040,N_9928,N_9392);
and UO_1041 (O_1041,N_9099,N_9659);
xnor UO_1042 (O_1042,N_9867,N_9630);
nor UO_1043 (O_1043,N_9414,N_9750);
xor UO_1044 (O_1044,N_9365,N_9866);
or UO_1045 (O_1045,N_9008,N_9592);
nand UO_1046 (O_1046,N_9868,N_9921);
nand UO_1047 (O_1047,N_9073,N_9343);
nand UO_1048 (O_1048,N_9964,N_9212);
nand UO_1049 (O_1049,N_9274,N_9786);
nor UO_1050 (O_1050,N_9836,N_9168);
xor UO_1051 (O_1051,N_9125,N_9686);
nand UO_1052 (O_1052,N_9089,N_9253);
and UO_1053 (O_1053,N_9836,N_9241);
xnor UO_1054 (O_1054,N_9930,N_9571);
nor UO_1055 (O_1055,N_9091,N_9869);
nand UO_1056 (O_1056,N_9342,N_9623);
nor UO_1057 (O_1057,N_9941,N_9195);
or UO_1058 (O_1058,N_9813,N_9933);
and UO_1059 (O_1059,N_9930,N_9724);
nand UO_1060 (O_1060,N_9887,N_9061);
and UO_1061 (O_1061,N_9906,N_9521);
and UO_1062 (O_1062,N_9312,N_9255);
xor UO_1063 (O_1063,N_9179,N_9374);
or UO_1064 (O_1064,N_9580,N_9472);
nor UO_1065 (O_1065,N_9278,N_9954);
nor UO_1066 (O_1066,N_9578,N_9838);
or UO_1067 (O_1067,N_9513,N_9950);
nor UO_1068 (O_1068,N_9916,N_9861);
nor UO_1069 (O_1069,N_9374,N_9408);
and UO_1070 (O_1070,N_9236,N_9793);
nor UO_1071 (O_1071,N_9256,N_9897);
nor UO_1072 (O_1072,N_9408,N_9571);
nor UO_1073 (O_1073,N_9775,N_9325);
nor UO_1074 (O_1074,N_9470,N_9483);
and UO_1075 (O_1075,N_9739,N_9823);
xnor UO_1076 (O_1076,N_9346,N_9769);
nand UO_1077 (O_1077,N_9499,N_9549);
nor UO_1078 (O_1078,N_9538,N_9432);
nand UO_1079 (O_1079,N_9637,N_9051);
and UO_1080 (O_1080,N_9994,N_9588);
nor UO_1081 (O_1081,N_9940,N_9544);
and UO_1082 (O_1082,N_9246,N_9873);
or UO_1083 (O_1083,N_9232,N_9569);
nand UO_1084 (O_1084,N_9463,N_9165);
xor UO_1085 (O_1085,N_9646,N_9053);
nand UO_1086 (O_1086,N_9595,N_9221);
or UO_1087 (O_1087,N_9289,N_9083);
nand UO_1088 (O_1088,N_9117,N_9378);
and UO_1089 (O_1089,N_9376,N_9787);
and UO_1090 (O_1090,N_9360,N_9314);
or UO_1091 (O_1091,N_9548,N_9886);
or UO_1092 (O_1092,N_9457,N_9463);
or UO_1093 (O_1093,N_9233,N_9953);
xor UO_1094 (O_1094,N_9688,N_9466);
nand UO_1095 (O_1095,N_9224,N_9886);
or UO_1096 (O_1096,N_9876,N_9522);
or UO_1097 (O_1097,N_9952,N_9979);
nand UO_1098 (O_1098,N_9331,N_9435);
nand UO_1099 (O_1099,N_9886,N_9464);
nor UO_1100 (O_1100,N_9402,N_9300);
nor UO_1101 (O_1101,N_9113,N_9727);
xor UO_1102 (O_1102,N_9147,N_9618);
nand UO_1103 (O_1103,N_9135,N_9472);
nand UO_1104 (O_1104,N_9105,N_9206);
nand UO_1105 (O_1105,N_9050,N_9219);
nand UO_1106 (O_1106,N_9092,N_9032);
or UO_1107 (O_1107,N_9838,N_9631);
nand UO_1108 (O_1108,N_9909,N_9693);
nor UO_1109 (O_1109,N_9463,N_9961);
or UO_1110 (O_1110,N_9832,N_9950);
xnor UO_1111 (O_1111,N_9141,N_9897);
nand UO_1112 (O_1112,N_9008,N_9574);
and UO_1113 (O_1113,N_9469,N_9821);
and UO_1114 (O_1114,N_9806,N_9877);
xnor UO_1115 (O_1115,N_9902,N_9376);
and UO_1116 (O_1116,N_9018,N_9595);
xor UO_1117 (O_1117,N_9676,N_9529);
nand UO_1118 (O_1118,N_9650,N_9347);
xnor UO_1119 (O_1119,N_9404,N_9151);
nand UO_1120 (O_1120,N_9351,N_9108);
xnor UO_1121 (O_1121,N_9857,N_9098);
nor UO_1122 (O_1122,N_9038,N_9454);
or UO_1123 (O_1123,N_9243,N_9809);
or UO_1124 (O_1124,N_9161,N_9338);
or UO_1125 (O_1125,N_9608,N_9951);
nand UO_1126 (O_1126,N_9343,N_9957);
xor UO_1127 (O_1127,N_9910,N_9945);
xor UO_1128 (O_1128,N_9747,N_9372);
nor UO_1129 (O_1129,N_9918,N_9264);
or UO_1130 (O_1130,N_9509,N_9653);
or UO_1131 (O_1131,N_9063,N_9273);
xnor UO_1132 (O_1132,N_9629,N_9302);
and UO_1133 (O_1133,N_9458,N_9013);
or UO_1134 (O_1134,N_9465,N_9642);
and UO_1135 (O_1135,N_9988,N_9381);
nor UO_1136 (O_1136,N_9355,N_9103);
or UO_1137 (O_1137,N_9377,N_9863);
and UO_1138 (O_1138,N_9190,N_9428);
nor UO_1139 (O_1139,N_9529,N_9591);
nand UO_1140 (O_1140,N_9812,N_9413);
nand UO_1141 (O_1141,N_9769,N_9229);
xnor UO_1142 (O_1142,N_9342,N_9063);
xnor UO_1143 (O_1143,N_9955,N_9925);
or UO_1144 (O_1144,N_9051,N_9851);
nor UO_1145 (O_1145,N_9711,N_9112);
nand UO_1146 (O_1146,N_9678,N_9229);
nand UO_1147 (O_1147,N_9158,N_9148);
xnor UO_1148 (O_1148,N_9128,N_9517);
nand UO_1149 (O_1149,N_9752,N_9737);
nand UO_1150 (O_1150,N_9621,N_9980);
or UO_1151 (O_1151,N_9875,N_9125);
nand UO_1152 (O_1152,N_9001,N_9658);
xor UO_1153 (O_1153,N_9690,N_9573);
nand UO_1154 (O_1154,N_9901,N_9584);
or UO_1155 (O_1155,N_9777,N_9671);
and UO_1156 (O_1156,N_9020,N_9205);
nand UO_1157 (O_1157,N_9404,N_9299);
nand UO_1158 (O_1158,N_9826,N_9527);
and UO_1159 (O_1159,N_9398,N_9417);
or UO_1160 (O_1160,N_9351,N_9568);
nor UO_1161 (O_1161,N_9598,N_9384);
and UO_1162 (O_1162,N_9963,N_9444);
xnor UO_1163 (O_1163,N_9228,N_9936);
and UO_1164 (O_1164,N_9251,N_9026);
and UO_1165 (O_1165,N_9837,N_9695);
nand UO_1166 (O_1166,N_9121,N_9276);
nand UO_1167 (O_1167,N_9578,N_9134);
nor UO_1168 (O_1168,N_9423,N_9725);
nand UO_1169 (O_1169,N_9295,N_9513);
and UO_1170 (O_1170,N_9777,N_9238);
nor UO_1171 (O_1171,N_9157,N_9716);
nand UO_1172 (O_1172,N_9895,N_9159);
nand UO_1173 (O_1173,N_9327,N_9830);
or UO_1174 (O_1174,N_9021,N_9460);
nor UO_1175 (O_1175,N_9955,N_9056);
nand UO_1176 (O_1176,N_9290,N_9087);
and UO_1177 (O_1177,N_9315,N_9486);
xnor UO_1178 (O_1178,N_9328,N_9584);
nand UO_1179 (O_1179,N_9999,N_9802);
xnor UO_1180 (O_1180,N_9964,N_9432);
or UO_1181 (O_1181,N_9141,N_9325);
nand UO_1182 (O_1182,N_9954,N_9463);
nand UO_1183 (O_1183,N_9424,N_9200);
or UO_1184 (O_1184,N_9897,N_9779);
xor UO_1185 (O_1185,N_9909,N_9160);
nor UO_1186 (O_1186,N_9586,N_9897);
and UO_1187 (O_1187,N_9030,N_9916);
or UO_1188 (O_1188,N_9454,N_9533);
or UO_1189 (O_1189,N_9561,N_9988);
or UO_1190 (O_1190,N_9719,N_9913);
and UO_1191 (O_1191,N_9775,N_9595);
nor UO_1192 (O_1192,N_9149,N_9648);
or UO_1193 (O_1193,N_9098,N_9244);
nand UO_1194 (O_1194,N_9971,N_9422);
and UO_1195 (O_1195,N_9711,N_9673);
xor UO_1196 (O_1196,N_9097,N_9448);
or UO_1197 (O_1197,N_9626,N_9682);
and UO_1198 (O_1198,N_9959,N_9539);
or UO_1199 (O_1199,N_9803,N_9482);
xnor UO_1200 (O_1200,N_9785,N_9302);
and UO_1201 (O_1201,N_9371,N_9878);
nor UO_1202 (O_1202,N_9339,N_9540);
and UO_1203 (O_1203,N_9089,N_9769);
and UO_1204 (O_1204,N_9354,N_9926);
nand UO_1205 (O_1205,N_9974,N_9771);
nor UO_1206 (O_1206,N_9110,N_9186);
nand UO_1207 (O_1207,N_9181,N_9002);
nand UO_1208 (O_1208,N_9981,N_9873);
and UO_1209 (O_1209,N_9792,N_9080);
and UO_1210 (O_1210,N_9263,N_9671);
nand UO_1211 (O_1211,N_9748,N_9966);
and UO_1212 (O_1212,N_9403,N_9060);
or UO_1213 (O_1213,N_9768,N_9209);
nor UO_1214 (O_1214,N_9662,N_9613);
nor UO_1215 (O_1215,N_9601,N_9337);
xor UO_1216 (O_1216,N_9082,N_9253);
nor UO_1217 (O_1217,N_9455,N_9393);
or UO_1218 (O_1218,N_9000,N_9574);
or UO_1219 (O_1219,N_9582,N_9766);
xor UO_1220 (O_1220,N_9059,N_9053);
nand UO_1221 (O_1221,N_9457,N_9802);
nor UO_1222 (O_1222,N_9642,N_9456);
nand UO_1223 (O_1223,N_9588,N_9720);
xor UO_1224 (O_1224,N_9003,N_9213);
xor UO_1225 (O_1225,N_9043,N_9801);
xor UO_1226 (O_1226,N_9189,N_9927);
xor UO_1227 (O_1227,N_9726,N_9522);
nor UO_1228 (O_1228,N_9565,N_9965);
nand UO_1229 (O_1229,N_9723,N_9937);
or UO_1230 (O_1230,N_9301,N_9473);
xor UO_1231 (O_1231,N_9409,N_9237);
and UO_1232 (O_1232,N_9425,N_9809);
or UO_1233 (O_1233,N_9674,N_9998);
nor UO_1234 (O_1234,N_9692,N_9712);
nand UO_1235 (O_1235,N_9311,N_9332);
xor UO_1236 (O_1236,N_9468,N_9739);
and UO_1237 (O_1237,N_9420,N_9450);
or UO_1238 (O_1238,N_9220,N_9979);
nand UO_1239 (O_1239,N_9191,N_9352);
xnor UO_1240 (O_1240,N_9192,N_9154);
nor UO_1241 (O_1241,N_9643,N_9100);
nand UO_1242 (O_1242,N_9910,N_9294);
nand UO_1243 (O_1243,N_9320,N_9529);
xnor UO_1244 (O_1244,N_9219,N_9959);
or UO_1245 (O_1245,N_9909,N_9471);
nand UO_1246 (O_1246,N_9661,N_9273);
nor UO_1247 (O_1247,N_9895,N_9655);
and UO_1248 (O_1248,N_9751,N_9172);
or UO_1249 (O_1249,N_9580,N_9856);
nand UO_1250 (O_1250,N_9046,N_9300);
nand UO_1251 (O_1251,N_9564,N_9872);
nor UO_1252 (O_1252,N_9498,N_9130);
xor UO_1253 (O_1253,N_9362,N_9081);
nand UO_1254 (O_1254,N_9064,N_9790);
nor UO_1255 (O_1255,N_9613,N_9644);
nand UO_1256 (O_1256,N_9612,N_9350);
nor UO_1257 (O_1257,N_9145,N_9644);
xor UO_1258 (O_1258,N_9647,N_9616);
nand UO_1259 (O_1259,N_9627,N_9571);
xnor UO_1260 (O_1260,N_9561,N_9718);
nand UO_1261 (O_1261,N_9348,N_9871);
or UO_1262 (O_1262,N_9592,N_9511);
or UO_1263 (O_1263,N_9869,N_9297);
and UO_1264 (O_1264,N_9503,N_9580);
nor UO_1265 (O_1265,N_9584,N_9285);
or UO_1266 (O_1266,N_9146,N_9536);
nand UO_1267 (O_1267,N_9372,N_9491);
nor UO_1268 (O_1268,N_9466,N_9629);
or UO_1269 (O_1269,N_9327,N_9457);
xor UO_1270 (O_1270,N_9700,N_9153);
xnor UO_1271 (O_1271,N_9499,N_9519);
and UO_1272 (O_1272,N_9287,N_9572);
xnor UO_1273 (O_1273,N_9217,N_9116);
xor UO_1274 (O_1274,N_9296,N_9680);
nand UO_1275 (O_1275,N_9961,N_9447);
nand UO_1276 (O_1276,N_9392,N_9876);
and UO_1277 (O_1277,N_9317,N_9169);
xor UO_1278 (O_1278,N_9957,N_9476);
and UO_1279 (O_1279,N_9814,N_9412);
nor UO_1280 (O_1280,N_9447,N_9869);
nand UO_1281 (O_1281,N_9953,N_9028);
nor UO_1282 (O_1282,N_9240,N_9508);
nand UO_1283 (O_1283,N_9853,N_9818);
or UO_1284 (O_1284,N_9979,N_9781);
nand UO_1285 (O_1285,N_9861,N_9144);
xnor UO_1286 (O_1286,N_9412,N_9346);
and UO_1287 (O_1287,N_9063,N_9366);
nor UO_1288 (O_1288,N_9765,N_9226);
xnor UO_1289 (O_1289,N_9337,N_9743);
xor UO_1290 (O_1290,N_9381,N_9412);
nor UO_1291 (O_1291,N_9569,N_9084);
and UO_1292 (O_1292,N_9086,N_9387);
and UO_1293 (O_1293,N_9266,N_9599);
and UO_1294 (O_1294,N_9247,N_9606);
and UO_1295 (O_1295,N_9950,N_9348);
nor UO_1296 (O_1296,N_9828,N_9668);
or UO_1297 (O_1297,N_9322,N_9626);
or UO_1298 (O_1298,N_9584,N_9422);
xnor UO_1299 (O_1299,N_9609,N_9049);
or UO_1300 (O_1300,N_9483,N_9295);
nand UO_1301 (O_1301,N_9570,N_9982);
and UO_1302 (O_1302,N_9840,N_9835);
xnor UO_1303 (O_1303,N_9444,N_9054);
or UO_1304 (O_1304,N_9400,N_9131);
and UO_1305 (O_1305,N_9697,N_9856);
and UO_1306 (O_1306,N_9548,N_9082);
or UO_1307 (O_1307,N_9856,N_9970);
nor UO_1308 (O_1308,N_9925,N_9653);
or UO_1309 (O_1309,N_9738,N_9766);
nand UO_1310 (O_1310,N_9085,N_9891);
and UO_1311 (O_1311,N_9281,N_9234);
and UO_1312 (O_1312,N_9589,N_9585);
and UO_1313 (O_1313,N_9099,N_9702);
and UO_1314 (O_1314,N_9677,N_9451);
or UO_1315 (O_1315,N_9357,N_9481);
or UO_1316 (O_1316,N_9144,N_9014);
and UO_1317 (O_1317,N_9866,N_9683);
and UO_1318 (O_1318,N_9119,N_9530);
or UO_1319 (O_1319,N_9261,N_9026);
nor UO_1320 (O_1320,N_9069,N_9562);
and UO_1321 (O_1321,N_9288,N_9646);
nand UO_1322 (O_1322,N_9945,N_9553);
nand UO_1323 (O_1323,N_9405,N_9723);
nor UO_1324 (O_1324,N_9840,N_9619);
xor UO_1325 (O_1325,N_9295,N_9838);
xor UO_1326 (O_1326,N_9065,N_9000);
and UO_1327 (O_1327,N_9083,N_9702);
nor UO_1328 (O_1328,N_9885,N_9686);
xor UO_1329 (O_1329,N_9725,N_9659);
nor UO_1330 (O_1330,N_9992,N_9744);
nand UO_1331 (O_1331,N_9505,N_9075);
and UO_1332 (O_1332,N_9041,N_9705);
or UO_1333 (O_1333,N_9605,N_9978);
xnor UO_1334 (O_1334,N_9878,N_9461);
xnor UO_1335 (O_1335,N_9298,N_9532);
and UO_1336 (O_1336,N_9830,N_9135);
nand UO_1337 (O_1337,N_9199,N_9213);
and UO_1338 (O_1338,N_9128,N_9233);
xor UO_1339 (O_1339,N_9899,N_9741);
nor UO_1340 (O_1340,N_9482,N_9456);
nor UO_1341 (O_1341,N_9608,N_9105);
and UO_1342 (O_1342,N_9380,N_9286);
nand UO_1343 (O_1343,N_9283,N_9201);
xnor UO_1344 (O_1344,N_9064,N_9267);
nand UO_1345 (O_1345,N_9021,N_9245);
xor UO_1346 (O_1346,N_9730,N_9898);
nand UO_1347 (O_1347,N_9057,N_9937);
nor UO_1348 (O_1348,N_9983,N_9937);
or UO_1349 (O_1349,N_9891,N_9861);
or UO_1350 (O_1350,N_9196,N_9370);
or UO_1351 (O_1351,N_9862,N_9008);
nand UO_1352 (O_1352,N_9521,N_9802);
nor UO_1353 (O_1353,N_9133,N_9485);
and UO_1354 (O_1354,N_9210,N_9983);
nand UO_1355 (O_1355,N_9574,N_9277);
nand UO_1356 (O_1356,N_9829,N_9400);
and UO_1357 (O_1357,N_9166,N_9184);
xor UO_1358 (O_1358,N_9498,N_9800);
nor UO_1359 (O_1359,N_9552,N_9762);
or UO_1360 (O_1360,N_9216,N_9435);
nor UO_1361 (O_1361,N_9419,N_9941);
nand UO_1362 (O_1362,N_9868,N_9465);
nand UO_1363 (O_1363,N_9895,N_9206);
and UO_1364 (O_1364,N_9244,N_9649);
or UO_1365 (O_1365,N_9962,N_9605);
xor UO_1366 (O_1366,N_9603,N_9467);
nand UO_1367 (O_1367,N_9139,N_9172);
nand UO_1368 (O_1368,N_9448,N_9107);
nand UO_1369 (O_1369,N_9821,N_9549);
xor UO_1370 (O_1370,N_9655,N_9458);
or UO_1371 (O_1371,N_9415,N_9680);
nor UO_1372 (O_1372,N_9122,N_9134);
nand UO_1373 (O_1373,N_9784,N_9298);
xor UO_1374 (O_1374,N_9302,N_9972);
or UO_1375 (O_1375,N_9739,N_9106);
nand UO_1376 (O_1376,N_9505,N_9757);
or UO_1377 (O_1377,N_9062,N_9913);
or UO_1378 (O_1378,N_9965,N_9312);
nand UO_1379 (O_1379,N_9038,N_9188);
nand UO_1380 (O_1380,N_9378,N_9568);
and UO_1381 (O_1381,N_9265,N_9833);
nor UO_1382 (O_1382,N_9996,N_9712);
xnor UO_1383 (O_1383,N_9157,N_9115);
xor UO_1384 (O_1384,N_9645,N_9008);
nand UO_1385 (O_1385,N_9300,N_9950);
nand UO_1386 (O_1386,N_9565,N_9853);
or UO_1387 (O_1387,N_9845,N_9435);
or UO_1388 (O_1388,N_9946,N_9983);
nor UO_1389 (O_1389,N_9518,N_9098);
xor UO_1390 (O_1390,N_9468,N_9352);
or UO_1391 (O_1391,N_9491,N_9219);
xnor UO_1392 (O_1392,N_9331,N_9152);
and UO_1393 (O_1393,N_9938,N_9290);
or UO_1394 (O_1394,N_9864,N_9367);
and UO_1395 (O_1395,N_9244,N_9439);
and UO_1396 (O_1396,N_9534,N_9977);
nor UO_1397 (O_1397,N_9404,N_9992);
or UO_1398 (O_1398,N_9157,N_9580);
nand UO_1399 (O_1399,N_9862,N_9477);
and UO_1400 (O_1400,N_9001,N_9355);
nand UO_1401 (O_1401,N_9797,N_9745);
or UO_1402 (O_1402,N_9528,N_9505);
nor UO_1403 (O_1403,N_9475,N_9887);
nor UO_1404 (O_1404,N_9188,N_9991);
nor UO_1405 (O_1405,N_9659,N_9493);
nand UO_1406 (O_1406,N_9937,N_9321);
nor UO_1407 (O_1407,N_9153,N_9816);
or UO_1408 (O_1408,N_9833,N_9142);
nand UO_1409 (O_1409,N_9687,N_9195);
or UO_1410 (O_1410,N_9282,N_9012);
xor UO_1411 (O_1411,N_9349,N_9883);
nor UO_1412 (O_1412,N_9499,N_9261);
nor UO_1413 (O_1413,N_9826,N_9209);
nand UO_1414 (O_1414,N_9861,N_9374);
nand UO_1415 (O_1415,N_9520,N_9809);
and UO_1416 (O_1416,N_9652,N_9096);
nand UO_1417 (O_1417,N_9637,N_9752);
and UO_1418 (O_1418,N_9244,N_9773);
and UO_1419 (O_1419,N_9595,N_9352);
nand UO_1420 (O_1420,N_9692,N_9320);
nand UO_1421 (O_1421,N_9361,N_9268);
or UO_1422 (O_1422,N_9228,N_9187);
and UO_1423 (O_1423,N_9209,N_9834);
and UO_1424 (O_1424,N_9730,N_9184);
or UO_1425 (O_1425,N_9005,N_9786);
nand UO_1426 (O_1426,N_9839,N_9799);
nor UO_1427 (O_1427,N_9247,N_9046);
and UO_1428 (O_1428,N_9525,N_9060);
or UO_1429 (O_1429,N_9287,N_9402);
or UO_1430 (O_1430,N_9310,N_9901);
xor UO_1431 (O_1431,N_9427,N_9565);
or UO_1432 (O_1432,N_9048,N_9920);
xnor UO_1433 (O_1433,N_9652,N_9361);
or UO_1434 (O_1434,N_9558,N_9518);
xnor UO_1435 (O_1435,N_9553,N_9189);
or UO_1436 (O_1436,N_9396,N_9234);
xor UO_1437 (O_1437,N_9023,N_9621);
nand UO_1438 (O_1438,N_9450,N_9690);
nor UO_1439 (O_1439,N_9715,N_9919);
and UO_1440 (O_1440,N_9740,N_9530);
nor UO_1441 (O_1441,N_9158,N_9761);
xnor UO_1442 (O_1442,N_9079,N_9526);
nor UO_1443 (O_1443,N_9988,N_9244);
nand UO_1444 (O_1444,N_9525,N_9491);
xor UO_1445 (O_1445,N_9501,N_9064);
xor UO_1446 (O_1446,N_9714,N_9474);
nand UO_1447 (O_1447,N_9992,N_9011);
nor UO_1448 (O_1448,N_9703,N_9376);
nor UO_1449 (O_1449,N_9652,N_9011);
or UO_1450 (O_1450,N_9309,N_9951);
and UO_1451 (O_1451,N_9706,N_9158);
or UO_1452 (O_1452,N_9789,N_9521);
or UO_1453 (O_1453,N_9922,N_9149);
or UO_1454 (O_1454,N_9779,N_9365);
or UO_1455 (O_1455,N_9785,N_9870);
or UO_1456 (O_1456,N_9589,N_9933);
or UO_1457 (O_1457,N_9048,N_9293);
xor UO_1458 (O_1458,N_9907,N_9269);
or UO_1459 (O_1459,N_9227,N_9382);
nor UO_1460 (O_1460,N_9796,N_9041);
or UO_1461 (O_1461,N_9545,N_9361);
xor UO_1462 (O_1462,N_9702,N_9489);
nor UO_1463 (O_1463,N_9594,N_9547);
xor UO_1464 (O_1464,N_9667,N_9734);
and UO_1465 (O_1465,N_9414,N_9280);
xor UO_1466 (O_1466,N_9272,N_9138);
nand UO_1467 (O_1467,N_9716,N_9856);
or UO_1468 (O_1468,N_9897,N_9051);
xor UO_1469 (O_1469,N_9953,N_9271);
and UO_1470 (O_1470,N_9797,N_9851);
and UO_1471 (O_1471,N_9383,N_9150);
nor UO_1472 (O_1472,N_9122,N_9303);
nor UO_1473 (O_1473,N_9714,N_9525);
nand UO_1474 (O_1474,N_9568,N_9126);
and UO_1475 (O_1475,N_9890,N_9963);
and UO_1476 (O_1476,N_9445,N_9817);
nand UO_1477 (O_1477,N_9865,N_9675);
nand UO_1478 (O_1478,N_9816,N_9722);
and UO_1479 (O_1479,N_9460,N_9675);
or UO_1480 (O_1480,N_9806,N_9006);
or UO_1481 (O_1481,N_9470,N_9603);
and UO_1482 (O_1482,N_9995,N_9694);
or UO_1483 (O_1483,N_9066,N_9402);
xnor UO_1484 (O_1484,N_9024,N_9116);
or UO_1485 (O_1485,N_9879,N_9545);
xor UO_1486 (O_1486,N_9838,N_9987);
and UO_1487 (O_1487,N_9647,N_9302);
or UO_1488 (O_1488,N_9622,N_9587);
nand UO_1489 (O_1489,N_9057,N_9039);
or UO_1490 (O_1490,N_9133,N_9259);
nor UO_1491 (O_1491,N_9806,N_9571);
nand UO_1492 (O_1492,N_9476,N_9006);
nor UO_1493 (O_1493,N_9995,N_9554);
xnor UO_1494 (O_1494,N_9222,N_9367);
xor UO_1495 (O_1495,N_9264,N_9897);
nor UO_1496 (O_1496,N_9147,N_9252);
xor UO_1497 (O_1497,N_9246,N_9842);
xnor UO_1498 (O_1498,N_9883,N_9977);
nand UO_1499 (O_1499,N_9727,N_9714);
endmodule