module basic_2000_20000_2500_10_levels_5xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nor U0 (N_0,In_989,In_1933);
and U1 (N_1,In_1881,In_1066);
or U2 (N_2,In_174,In_111);
nand U3 (N_3,In_948,In_598);
or U4 (N_4,In_797,In_708);
and U5 (N_5,In_1857,In_1316);
nor U6 (N_6,In_823,In_1051);
xnor U7 (N_7,In_201,In_557);
nor U8 (N_8,In_536,In_810);
or U9 (N_9,In_51,In_1766);
nand U10 (N_10,In_11,In_864);
xnor U11 (N_11,In_1809,In_1624);
nand U12 (N_12,In_356,In_22);
and U13 (N_13,In_894,In_326);
nand U14 (N_14,In_1210,In_1107);
and U15 (N_15,In_1799,In_1685);
xor U16 (N_16,In_149,In_995);
or U17 (N_17,In_1007,In_712);
and U18 (N_18,In_173,In_1805);
xnor U19 (N_19,In_583,In_1558);
nand U20 (N_20,In_1348,In_628);
nand U21 (N_21,In_58,In_1431);
nand U22 (N_22,In_167,In_1560);
xnor U23 (N_23,In_368,In_771);
and U24 (N_24,In_455,In_451);
or U25 (N_25,In_231,In_1890);
nand U26 (N_26,In_1669,In_1607);
nand U27 (N_27,In_124,In_669);
nor U28 (N_28,In_460,In_905);
and U29 (N_29,In_125,In_103);
or U30 (N_30,In_1276,In_1787);
nor U31 (N_31,In_280,In_172);
and U32 (N_32,In_1729,In_640);
and U33 (N_33,In_139,In_1580);
nor U34 (N_34,In_24,In_959);
nand U35 (N_35,In_644,In_1676);
nor U36 (N_36,In_886,In_256);
and U37 (N_37,In_1855,In_1414);
and U38 (N_38,In_1073,In_1067);
nor U39 (N_39,In_129,In_316);
nand U40 (N_40,In_1760,In_90);
xor U41 (N_41,In_182,In_93);
or U42 (N_42,In_377,In_1842);
and U43 (N_43,In_1606,In_1437);
xor U44 (N_44,In_1812,In_1638);
nand U45 (N_45,In_1869,In_1736);
and U46 (N_46,In_1938,In_1806);
or U47 (N_47,In_1042,In_867);
nor U48 (N_48,In_1070,In_1002);
and U49 (N_49,In_909,In_1053);
nor U50 (N_50,In_384,In_100);
nor U51 (N_51,In_1514,In_219);
xnor U52 (N_52,In_1436,In_1557);
nand U53 (N_53,In_1555,In_1103);
nor U54 (N_54,In_117,In_791);
or U55 (N_55,In_786,In_1292);
nor U56 (N_56,In_1953,In_1393);
nand U57 (N_57,In_458,In_321);
nand U58 (N_58,In_1033,In_1159);
or U59 (N_59,In_136,In_802);
nor U60 (N_60,In_1291,In_1728);
nor U61 (N_61,In_1228,In_928);
nand U62 (N_62,In_1828,In_1678);
nand U63 (N_63,In_169,In_1388);
nand U64 (N_64,In_1029,In_1453);
and U65 (N_65,In_666,In_574);
nand U66 (N_66,In_1982,In_1796);
and U67 (N_67,In_1046,In_1548);
xor U68 (N_68,In_1961,In_497);
and U69 (N_69,In_302,In_1776);
and U70 (N_70,In_829,In_880);
and U71 (N_71,In_578,In_725);
nor U72 (N_72,In_713,In_1127);
nor U73 (N_73,In_32,In_661);
nor U74 (N_74,In_422,In_199);
and U75 (N_75,In_1145,In_1894);
or U76 (N_76,In_1625,In_1352);
xor U77 (N_77,In_1720,In_593);
or U78 (N_78,In_1732,In_1820);
and U79 (N_79,In_1011,In_314);
or U80 (N_80,In_1079,In_275);
nor U81 (N_81,In_1199,In_261);
nor U82 (N_82,In_1153,In_1602);
xor U83 (N_83,In_1130,In_1251);
and U84 (N_84,In_505,In_648);
or U85 (N_85,In_507,In_335);
nand U86 (N_86,In_859,In_1919);
and U87 (N_87,In_134,In_571);
nand U88 (N_88,In_1432,In_917);
and U89 (N_89,In_9,In_843);
or U90 (N_90,In_1775,In_346);
and U91 (N_91,In_1567,In_34);
and U92 (N_92,In_1986,In_1731);
nand U93 (N_93,In_936,In_60);
and U94 (N_94,In_370,In_127);
nand U95 (N_95,In_1659,In_25);
nor U96 (N_96,In_1257,In_194);
nand U97 (N_97,In_1464,In_555);
nand U98 (N_98,In_271,In_307);
nor U99 (N_99,In_535,In_1407);
nor U100 (N_100,In_1412,In_1394);
or U101 (N_101,In_1928,In_1670);
and U102 (N_102,In_1610,In_728);
nor U103 (N_103,In_1131,In_1296);
nor U104 (N_104,In_509,In_387);
nor U105 (N_105,In_1654,In_1517);
nor U106 (N_106,In_733,In_643);
xor U107 (N_107,In_793,In_1113);
nand U108 (N_108,In_964,In_230);
or U109 (N_109,In_1510,In_308);
and U110 (N_110,In_1402,In_228);
or U111 (N_111,In_39,In_1429);
xnor U112 (N_112,In_1120,In_626);
xnor U113 (N_113,In_372,In_1149);
and U114 (N_114,In_1154,In_1155);
and U115 (N_115,In_1507,In_778);
nor U116 (N_116,In_1613,In_545);
nor U117 (N_117,In_1768,In_1868);
or U118 (N_118,In_1588,In_1318);
nor U119 (N_119,In_343,In_1460);
and U120 (N_120,In_727,In_1197);
nand U121 (N_121,In_1069,In_160);
xnor U122 (N_122,In_1821,In_1789);
nand U123 (N_123,In_1048,In_896);
nor U124 (N_124,In_763,In_629);
nor U125 (N_125,In_144,In_907);
or U126 (N_126,In_1382,In_1955);
nand U127 (N_127,In_1322,In_1829);
and U128 (N_128,In_1288,In_1977);
or U129 (N_129,In_1188,In_652);
and U130 (N_130,In_488,In_1234);
nor U131 (N_131,In_526,In_130);
xor U132 (N_132,In_1765,In_937);
nor U133 (N_133,In_893,In_1173);
or U134 (N_134,In_722,In_1981);
and U135 (N_135,In_1932,In_1827);
nand U136 (N_136,In_804,In_1274);
xor U137 (N_137,In_576,In_1744);
or U138 (N_138,In_1930,In_1494);
xor U139 (N_139,In_1873,In_1049);
nor U140 (N_140,In_825,In_296);
and U141 (N_141,In_1823,In_255);
or U142 (N_142,In_1704,In_195);
or U143 (N_143,In_133,In_1600);
nor U144 (N_144,In_1405,In_1245);
nand U145 (N_145,In_1506,In_1802);
nor U146 (N_146,In_1942,In_1550);
and U147 (N_147,In_73,In_1608);
and U148 (N_148,In_1644,In_599);
or U149 (N_149,In_105,In_516);
nand U150 (N_150,In_945,In_1254);
and U151 (N_151,In_756,In_1259);
and U152 (N_152,In_1944,In_438);
xor U153 (N_153,In_1653,In_1293);
or U154 (N_154,In_600,In_883);
nor U155 (N_155,In_863,In_597);
nor U156 (N_156,In_243,In_339);
xnor U157 (N_157,In_1878,In_519);
nand U158 (N_158,In_664,In_118);
and U159 (N_159,In_1454,In_879);
and U160 (N_160,In_987,In_374);
or U161 (N_161,In_1660,In_608);
and U162 (N_162,In_1770,In_785);
and U163 (N_163,In_483,In_476);
nand U164 (N_164,In_425,In_1939);
or U165 (N_165,In_1618,In_1998);
nor U166 (N_166,In_1110,In_1343);
nor U167 (N_167,In_417,In_913);
nand U168 (N_168,In_567,In_1418);
nor U169 (N_169,In_703,In_1512);
nor U170 (N_170,In_482,In_313);
nand U171 (N_171,In_1683,In_1708);
and U172 (N_172,In_1746,In_1834);
or U173 (N_173,In_1723,In_1673);
nor U174 (N_174,In_1469,In_1688);
nand U175 (N_175,In_614,In_1022);
and U176 (N_176,In_632,In_1275);
nand U177 (N_177,In_480,In_116);
and U178 (N_178,In_768,In_143);
nor U179 (N_179,In_932,In_1907);
nand U180 (N_180,In_457,In_1526);
nor U181 (N_181,In_1417,In_1208);
nand U182 (N_182,In_1895,In_348);
or U183 (N_183,In_1767,In_889);
or U184 (N_184,In_1097,In_579);
nor U185 (N_185,In_1725,In_1129);
and U186 (N_186,In_657,In_1957);
nand U187 (N_187,In_1219,In_427);
and U188 (N_188,In_1747,In_1573);
nor U189 (N_189,In_341,In_1969);
nand U190 (N_190,In_1397,In_1190);
nand U191 (N_191,In_122,In_1287);
or U192 (N_192,In_215,In_43);
and U193 (N_193,In_1643,In_1075);
nor U194 (N_194,In_1759,In_289);
or U195 (N_195,In_847,In_630);
nor U196 (N_196,In_1546,In_973);
nor U197 (N_197,In_1439,In_1327);
nor U198 (N_198,In_991,In_393);
or U199 (N_199,In_151,In_115);
nor U200 (N_200,In_415,In_1310);
or U201 (N_201,In_1456,In_150);
nand U202 (N_202,In_826,In_1222);
nor U203 (N_203,In_1739,In_52);
xnor U204 (N_204,In_1921,In_753);
nand U205 (N_205,In_464,In_101);
or U206 (N_206,In_1909,In_1380);
nor U207 (N_207,In_1658,In_1628);
nor U208 (N_208,In_1603,In_984);
xor U209 (N_209,In_463,In_200);
or U210 (N_210,In_1003,In_446);
or U211 (N_211,In_1699,In_342);
nor U212 (N_212,In_546,In_1248);
nor U213 (N_213,In_426,In_752);
or U214 (N_214,In_1421,In_359);
and U215 (N_215,In_919,In_809);
or U216 (N_216,In_774,In_240);
nor U217 (N_217,In_962,In_1693);
nand U218 (N_218,In_1164,In_158);
nor U219 (N_219,In_1238,In_975);
or U220 (N_220,In_564,In_1966);
or U221 (N_221,In_259,In_503);
or U222 (N_222,In_1843,In_1636);
and U223 (N_223,In_999,In_1064);
xnor U224 (N_224,In_156,In_27);
xnor U225 (N_225,In_450,In_747);
nand U226 (N_226,In_1779,In_495);
nand U227 (N_227,In_755,In_1118);
or U228 (N_228,In_1370,In_94);
nor U229 (N_229,In_554,In_462);
nand U230 (N_230,In_1195,In_327);
or U231 (N_231,In_606,In_508);
xor U232 (N_232,In_1888,In_1390);
nor U233 (N_233,In_16,In_469);
nand U234 (N_234,In_1232,In_246);
nand U235 (N_235,In_1124,In_189);
nand U236 (N_236,In_1443,In_1183);
nand U237 (N_237,In_1849,In_796);
nand U238 (N_238,In_954,In_1745);
and U239 (N_239,In_266,In_1386);
or U240 (N_240,In_1213,In_1698);
nand U241 (N_241,In_254,In_155);
or U242 (N_242,In_330,In_741);
nand U243 (N_243,In_1534,In_104);
and U244 (N_244,In_1467,In_588);
or U245 (N_245,In_846,In_1383);
and U246 (N_246,In_382,In_1959);
nor U247 (N_247,In_1312,In_1950);
nor U248 (N_248,In_1055,In_988);
or U249 (N_249,In_328,In_1952);
and U250 (N_250,In_977,In_336);
or U251 (N_251,In_279,In_1750);
nand U252 (N_252,In_1810,In_1413);
nor U253 (N_253,In_402,In_0);
or U254 (N_254,In_398,In_636);
nor U255 (N_255,In_1169,In_448);
and U256 (N_256,In_258,In_452);
xnor U257 (N_257,In_1020,In_1143);
nand U258 (N_258,In_1611,In_1269);
xor U259 (N_259,In_1754,In_761);
nand U260 (N_260,In_1984,In_968);
and U261 (N_261,In_474,In_1419);
and U262 (N_262,In_20,In_709);
xnor U263 (N_263,In_1672,In_1114);
nor U264 (N_264,In_1740,In_381);
nor U265 (N_265,In_1062,In_720);
nor U266 (N_266,In_1844,In_1374);
nor U267 (N_267,In_1911,In_613);
or U268 (N_268,In_1864,In_62);
xor U269 (N_269,In_1160,In_515);
xnor U270 (N_270,In_1784,In_544);
nor U271 (N_271,In_1426,In_929);
nand U272 (N_272,In_1924,In_1264);
or U273 (N_273,In_585,In_1043);
or U274 (N_274,In_1572,In_1449);
nand U275 (N_275,In_409,In_758);
nand U276 (N_276,In_1323,In_852);
nor U277 (N_277,In_1218,In_1866);
and U278 (N_278,In_420,In_89);
nand U279 (N_279,In_26,In_815);
or U280 (N_280,In_1294,In_924);
nor U281 (N_281,In_1462,In_877);
and U282 (N_282,In_860,In_1363);
nand U283 (N_283,In_850,In_1076);
and U284 (N_284,In_1031,In_1123);
and U285 (N_285,In_1531,In_1349);
and U286 (N_286,In_1757,In_1427);
xor U287 (N_287,In_888,In_1639);
nor U288 (N_288,In_357,In_1781);
nor U289 (N_289,In_1622,In_1176);
and U290 (N_290,In_1023,In_1202);
and U291 (N_291,In_1927,In_1121);
nand U292 (N_292,In_107,In_524);
nand U293 (N_293,In_742,In_1201);
nor U294 (N_294,In_1267,In_1299);
and U295 (N_295,In_938,In_1451);
and U296 (N_296,In_542,In_1326);
nor U297 (N_297,In_1904,In_1461);
nand U298 (N_298,In_290,In_354);
nor U299 (N_299,In_565,In_1148);
or U300 (N_300,In_40,In_1224);
xnor U301 (N_301,In_186,In_1306);
xor U302 (N_302,In_1956,In_1320);
nand U303 (N_303,In_787,In_1655);
nor U304 (N_304,In_449,In_112);
xor U305 (N_305,In_903,In_83);
or U306 (N_306,In_349,In_908);
nand U307 (N_307,In_649,In_589);
nor U308 (N_308,In_247,In_715);
xnor U309 (N_309,In_487,In_334);
nor U310 (N_310,In_1015,In_874);
or U311 (N_311,In_910,In_273);
and U312 (N_312,In_1398,In_1499);
or U313 (N_313,In_770,In_414);
nand U314 (N_314,In_734,In_695);
or U315 (N_315,In_1205,In_744);
nand U316 (N_316,In_878,In_1008);
or U317 (N_317,In_244,In_548);
nand U318 (N_318,In_220,In_759);
and U319 (N_319,In_876,In_260);
and U320 (N_320,In_216,In_871);
or U321 (N_321,In_1063,In_670);
and U322 (N_322,In_499,In_739);
and U323 (N_323,In_1778,In_625);
or U324 (N_324,In_413,In_206);
nor U325 (N_325,In_1415,In_942);
or U326 (N_326,In_1865,In_940);
and U327 (N_327,In_963,In_1543);
nor U328 (N_328,In_830,In_504);
and U329 (N_329,In_1112,In_1798);
and U330 (N_330,In_1595,In_803);
or U331 (N_331,In_1214,In_1695);
nand U332 (N_332,In_310,In_424);
or U333 (N_333,In_538,In_1652);
and U334 (N_334,In_1125,In_6);
and U335 (N_335,In_396,In_193);
or U336 (N_336,In_239,In_673);
nand U337 (N_337,In_743,In_1255);
xor U338 (N_338,In_1917,In_137);
or U339 (N_339,In_1883,In_808);
or U340 (N_340,In_1491,In_85);
or U341 (N_341,In_453,In_479);
nand U342 (N_342,In_1646,In_935);
xnor U343 (N_343,In_1111,In_559);
or U344 (N_344,In_1925,In_1045);
and U345 (N_345,In_659,In_1592);
and U346 (N_346,In_1715,In_1330);
nor U347 (N_347,In_1701,In_1762);
nor U348 (N_348,In_895,In_1408);
or U349 (N_349,In_784,In_660);
xor U350 (N_350,In_135,In_1285);
and U351 (N_351,In_1447,In_1086);
nor U352 (N_352,In_202,In_865);
nand U353 (N_353,In_461,In_371);
nor U354 (N_354,In_1325,In_510);
xor U355 (N_355,In_534,In_750);
or U356 (N_356,In_835,In_1501);
and U357 (N_357,In_99,In_543);
nor U358 (N_358,In_798,In_1138);
nand U359 (N_359,In_217,In_1900);
nand U360 (N_360,In_306,In_33);
nor U361 (N_361,In_1337,In_408);
or U362 (N_362,In_87,In_1231);
and U363 (N_363,In_286,In_179);
or U364 (N_364,In_74,In_1818);
or U365 (N_365,In_1424,In_1428);
and U366 (N_366,In_1877,In_1584);
or U367 (N_367,In_1711,In_28);
xnor U368 (N_368,In_378,In_854);
nor U369 (N_369,In_1266,In_1885);
nor U370 (N_370,In_572,In_320);
nor U371 (N_371,In_868,In_1975);
nand U372 (N_372,In_1331,In_1466);
or U373 (N_373,In_272,In_944);
or U374 (N_374,In_1458,In_1940);
nand U375 (N_375,In_1052,In_914);
or U376 (N_376,In_573,In_1126);
and U377 (N_377,In_1246,In_1498);
nand U378 (N_378,In_57,In_208);
or U379 (N_379,In_916,In_1479);
or U380 (N_380,In_1241,In_1553);
or U381 (N_381,In_1662,In_533);
nor U382 (N_382,In_442,In_1175);
or U383 (N_383,In_584,In_178);
or U384 (N_384,In_655,In_605);
or U385 (N_385,In_485,In_1375);
nand U386 (N_386,In_1936,In_1242);
or U387 (N_387,In_570,In_1283);
nor U388 (N_388,In_1356,In_958);
or U389 (N_389,In_1128,In_1170);
xor U390 (N_390,In_1085,In_1511);
and U391 (N_391,In_211,In_61);
nand U392 (N_392,In_1867,In_783);
and U393 (N_393,In_1490,In_1263);
and U394 (N_394,In_501,In_1005);
nand U395 (N_395,In_1184,In_762);
xnor U396 (N_396,In_15,In_1240);
nor U397 (N_397,In_1152,In_300);
and U398 (N_398,In_1935,In_1100);
nand U399 (N_399,In_1281,In_807);
or U400 (N_400,In_1099,In_706);
and U401 (N_401,In_775,In_1528);
and U402 (N_402,In_1562,In_1362);
and U403 (N_403,In_701,In_729);
nand U404 (N_404,In_1619,In_1492);
nor U405 (N_405,In_407,In_1139);
or U406 (N_406,In_490,In_410);
xnor U407 (N_407,In_1633,In_665);
nor U408 (N_408,In_899,In_748);
and U409 (N_409,In_1756,In_1438);
or U410 (N_410,In_79,In_1420);
nand U411 (N_411,In_882,In_383);
or U412 (N_412,In_325,In_1722);
or U413 (N_413,In_994,In_1645);
or U414 (N_414,In_1786,In_245);
nor U415 (N_415,In_1792,In_920);
nor U416 (N_416,In_1230,In_185);
xor U417 (N_417,In_4,In_1682);
xnor U418 (N_418,In_885,In_1972);
and U419 (N_419,In_745,In_819);
nor U420 (N_420,In_820,In_177);
nor U421 (N_421,In_1340,In_1997);
or U422 (N_422,In_517,In_514);
and U423 (N_423,In_806,In_738);
or U424 (N_424,In_1171,In_257);
nand U425 (N_425,In_1634,In_154);
nand U426 (N_426,In_1880,In_1568);
nor U427 (N_427,In_454,In_672);
nor U428 (N_428,In_162,In_1385);
and U429 (N_429,In_1477,In_140);
nor U430 (N_430,In_1674,In_401);
or U431 (N_431,In_1496,In_1830);
and U432 (N_432,In_612,In_1694);
nand U433 (N_433,In_223,In_1596);
nor U434 (N_434,In_1065,In_1247);
or U435 (N_435,In_1017,In_840);
nor U436 (N_436,In_1117,In_262);
xor U437 (N_437,In_1379,In_692);
nor U438 (N_438,In_653,In_355);
xor U439 (N_439,In_1481,In_971);
or U440 (N_440,In_468,In_965);
nor U441 (N_441,In_780,In_931);
xnor U442 (N_442,In_925,In_203);
nor U443 (N_443,In_1886,In_858);
nand U444 (N_444,In_813,In_278);
nand U445 (N_445,In_891,In_1870);
nand U446 (N_446,In_1423,In_1132);
nand U447 (N_447,In_1301,In_56);
and U448 (N_448,In_631,In_88);
and U449 (N_449,In_724,In_1627);
and U450 (N_450,In_1353,In_855);
nor U451 (N_451,In_1027,In_210);
nand U452 (N_452,In_1513,In_1430);
and U453 (N_453,In_71,In_431);
nor U454 (N_454,In_1000,In_961);
and U455 (N_455,In_176,In_941);
nor U456 (N_456,In_1785,In_765);
nor U457 (N_457,In_904,In_63);
xnor U458 (N_458,In_1180,In_1090);
or U459 (N_459,In_1119,In_1875);
nand U460 (N_460,In_1036,In_1142);
xnor U461 (N_461,In_654,In_736);
nand U462 (N_462,In_1707,In_1300);
and U463 (N_463,In_1813,In_1297);
and U464 (N_464,In_596,In_1915);
nand U465 (N_465,In_1542,In_721);
and U466 (N_466,In_754,In_1667);
and U467 (N_467,In_873,In_1450);
nand U468 (N_468,In_1743,In_1157);
or U469 (N_469,In_209,In_592);
nand U470 (N_470,In_1657,In_1135);
nor U471 (N_471,In_1001,In_486);
or U472 (N_472,In_1544,In_651);
and U473 (N_473,In_418,In_1500);
nor U474 (N_474,In_1578,In_168);
nor U475 (N_475,In_238,In_1617);
or U476 (N_476,In_1705,In_998);
or U477 (N_477,In_1605,In_1012);
nor U478 (N_478,In_1249,In_817);
and U479 (N_479,In_1913,In_697);
nor U480 (N_480,In_1755,In_856);
xnor U481 (N_481,In_1282,In_184);
or U482 (N_482,In_1575,In_556);
nand U483 (N_483,In_1091,In_1474);
nand U484 (N_484,In_1772,In_506);
or U485 (N_485,In_686,In_1223);
nand U486 (N_486,In_687,In_1037);
nand U487 (N_487,In_638,In_831);
nor U488 (N_488,In_428,In_1751);
and U489 (N_489,In_1763,In_939);
nand U490 (N_490,In_49,In_1044);
nor U491 (N_491,In_166,In_465);
or U492 (N_492,In_126,In_478);
xnor U493 (N_493,In_601,In_365);
nor U494 (N_494,In_1172,In_952);
xnor U495 (N_495,In_1808,In_1105);
and U496 (N_496,In_790,In_1010);
or U497 (N_497,In_749,In_1116);
nand U498 (N_498,In_433,In_1404);
or U499 (N_499,In_329,In_818);
nand U500 (N_500,In_1523,In_1258);
and U501 (N_501,In_1978,In_1906);
or U502 (N_502,In_119,In_1571);
or U503 (N_503,In_1753,In_1963);
xnor U504 (N_504,In_492,In_624);
or U505 (N_505,In_389,In_1182);
or U506 (N_506,In_1509,In_1435);
nor U507 (N_507,In_5,In_72);
or U508 (N_508,In_493,In_1156);
and U509 (N_509,In_972,In_1752);
nor U510 (N_510,In_473,In_1167);
or U511 (N_511,In_1177,In_1522);
or U512 (N_512,In_207,In_1376);
and U513 (N_513,In_1604,In_429);
nand U514 (N_514,In_782,In_1059);
nor U515 (N_515,In_662,In_1533);
or U516 (N_516,In_645,In_1358);
or U517 (N_517,In_1615,In_441);
or U518 (N_518,In_1268,In_1191);
or U519 (N_519,In_1648,In_985);
nor U520 (N_520,In_658,In_1516);
nand U521 (N_521,In_1087,In_707);
xnor U522 (N_522,In_236,In_769);
nand U523 (N_523,In_1315,In_1215);
and U524 (N_524,In_1361,In_1561);
and U525 (N_525,In_1040,In_323);
and U526 (N_526,In_694,In_730);
or U527 (N_527,In_974,In_1505);
or U528 (N_528,In_293,In_214);
and U529 (N_529,In_1220,In_1943);
or U530 (N_530,In_529,In_682);
or U531 (N_531,In_301,In_1713);
and U532 (N_532,In_1317,In_699);
xnor U533 (N_533,In_1656,In_97);
nor U534 (N_534,In_1058,In_59);
nand U535 (N_535,In_406,In_322);
or U536 (N_536,In_1816,In_277);
nand U537 (N_537,In_575,In_607);
nor U538 (N_538,In_1692,In_267);
and U539 (N_539,In_1244,In_1920);
and U540 (N_540,In_1179,In_1614);
nand U541 (N_541,In_1077,In_1710);
xor U542 (N_542,In_558,In_1651);
or U543 (N_543,In_1271,In_1861);
or U544 (N_544,In_1389,In_1009);
nand U545 (N_545,In_1194,In_1668);
and U546 (N_546,In_1050,In_1366);
nand U547 (N_547,In_1529,In_319);
or U548 (N_548,In_1444,In_956);
or U549 (N_549,In_312,In_29);
or U550 (N_550,In_547,In_362);
nor U551 (N_551,In_1239,In_95);
and U552 (N_552,In_656,In_911);
nand U553 (N_553,In_1583,In_1166);
nor U554 (N_554,In_153,In_1289);
nand U555 (N_555,In_1525,In_581);
and U556 (N_556,In_1872,In_718);
and U557 (N_557,In_1161,In_1344);
nor U558 (N_558,In_1937,In_76);
nand U559 (N_559,In_496,In_1902);
nand U560 (N_560,In_1082,In_960);
nand U561 (N_561,In_617,In_1021);
and U562 (N_562,In_1028,In_1137);
or U563 (N_563,In_1503,In_1313);
nor U564 (N_564,In_1764,In_1863);
nand U565 (N_565,In_1780,In_1996);
and U566 (N_566,In_1089,In_1758);
or U567 (N_567,In_1630,In_901);
or U568 (N_568,In_108,In_990);
or U569 (N_569,In_1095,In_367);
and U570 (N_570,In_264,In_1733);
nor U571 (N_571,In_477,In_1054);
nand U572 (N_572,In_1585,In_1594);
nor U573 (N_573,In_252,In_67);
and U574 (N_574,In_1187,In_1338);
or U575 (N_575,In_224,In_890);
nor U576 (N_576,In_623,In_688);
nand U577 (N_577,In_435,In_1931);
nor U578 (N_578,In_55,In_80);
or U579 (N_579,In_849,In_1341);
nand U580 (N_580,In_434,In_1463);
nand U581 (N_581,In_1712,In_1473);
nand U582 (N_582,In_353,In_197);
or U583 (N_583,In_1941,In_1250);
nor U584 (N_584,In_142,In_110);
xnor U585 (N_585,In_1748,In_838);
xnor U586 (N_586,In_1593,In_45);
nor U587 (N_587,In_502,In_1101);
or U588 (N_588,In_1039,In_951);
and U589 (N_589,In_1236,In_520);
nor U590 (N_590,In_421,In_1206);
nand U591 (N_591,In_1068,In_3);
and U592 (N_592,In_1721,In_950);
nor U593 (N_593,In_304,In_731);
and U594 (N_594,In_128,In_1504);
or U595 (N_595,In_96,In_1273);
and U596 (N_596,In_539,In_1677);
xnor U597 (N_597,In_811,In_1518);
or U598 (N_598,In_603,In_416);
and U599 (N_599,In_1227,In_1416);
nor U600 (N_600,In_21,In_1783);
or U601 (N_601,In_1845,In_622);
and U602 (N_602,In_1217,In_1032);
or U603 (N_603,In_1144,In_1189);
nor U604 (N_604,In_1749,In_440);
and U605 (N_605,In_1047,In_1899);
or U606 (N_606,In_248,In_1400);
nor U607 (N_607,In_569,In_1801);
or U608 (N_608,In_121,In_746);
nand U609 (N_609,In_726,In_1335);
and U610 (N_610,In_1631,In_1581);
nor U611 (N_611,In_1104,In_1409);
or U612 (N_612,In_1468,In_1976);
and U613 (N_613,In_1832,In_171);
xnor U614 (N_614,In_351,In_132);
nand U615 (N_615,In_1235,In_30);
or U616 (N_616,In_347,In_1489);
or U617 (N_617,In_253,In_799);
or U618 (N_618,In_970,In_1387);
and U619 (N_619,In_48,In_735);
nand U620 (N_620,In_1597,In_1472);
and U621 (N_621,In_1262,In_620);
or U622 (N_622,In_1256,In_1284);
and U623 (N_623,In_1401,In_553);
or U624 (N_624,In_1378,In_376);
or U625 (N_625,In_1871,In_1280);
or U626 (N_626,In_7,In_698);
and U627 (N_627,In_997,In_1345);
nand U628 (N_628,In_1837,In_1056);
nor U629 (N_629,In_345,In_364);
nor U630 (N_630,In_540,In_1570);
nand U631 (N_631,In_1488,In_1874);
xor U632 (N_632,In_957,In_537);
and U633 (N_633,In_1493,In_1470);
nor U634 (N_634,In_1396,In_1689);
and U635 (N_635,In_494,In_1162);
nor U636 (N_636,In_164,In_943);
nand U637 (N_637,In_1502,In_205);
nor U638 (N_638,In_305,In_311);
and U639 (N_639,In_1434,In_737);
or U640 (N_640,In_1229,In_1314);
or U641 (N_641,In_1916,In_776);
and U642 (N_642,In_1882,In_1838);
and U643 (N_643,In_646,In_380);
nand U644 (N_644,In_902,In_1333);
xor U645 (N_645,In_616,In_1072);
xnor U646 (N_646,In_1847,In_432);
and U647 (N_647,In_1302,In_862);
or U648 (N_648,In_1038,In_1270);
and U649 (N_649,In_1535,In_1980);
xor U650 (N_650,In_647,In_1949);
nand U651 (N_651,In_1369,In_221);
or U652 (N_652,In_1853,In_1181);
nor U653 (N_653,In_1918,In_906);
and U654 (N_654,In_148,In_1025);
nand U655 (N_655,In_1856,In_1962);
or U656 (N_656,In_1665,In_513);
and U657 (N_657,In_1486,In_1);
and U658 (N_658,In_1988,In_1859);
and U659 (N_659,In_609,In_1876);
nor U660 (N_660,In_1679,In_333);
nand U661 (N_661,In_795,In_1372);
or U662 (N_662,In_1616,In_1260);
nor U663 (N_663,In_824,In_1591);
and U664 (N_664,In_930,In_602);
nand U665 (N_665,In_1730,In_781);
or U666 (N_666,In_1532,In_566);
nand U667 (N_667,In_1342,In_77);
and U668 (N_668,In_1286,In_397);
xor U669 (N_669,In_532,In_1084);
xnor U670 (N_670,In_618,In_1716);
and U671 (N_671,In_1092,In_1237);
xor U672 (N_672,In_857,In_1018);
or U673 (N_673,In_1680,In_1265);
or U674 (N_674,In_1841,In_1146);
nand U675 (N_675,In_1515,In_1034);
and U676 (N_676,In_1442,In_1440);
nor U677 (N_677,In_1696,In_705);
nor U678 (N_678,In_1989,In_404);
or U679 (N_679,In_1016,In_227);
and U680 (N_680,In_1307,In_915);
xor U681 (N_681,In_1621,In_1649);
or U682 (N_682,In_779,In_1411);
nor U683 (N_683,In_1556,In_777);
and U684 (N_684,In_1093,In_352);
xor U685 (N_685,In_1253,In_218);
nand U686 (N_686,In_690,In_1800);
or U687 (N_687,In_1738,In_212);
nand U688 (N_688,In_577,In_1860);
nand U689 (N_689,In_1094,In_717);
and U690 (N_690,In_949,In_1803);
xnor U691 (N_691,In_1967,In_1186);
and U692 (N_692,In_641,In_180);
and U693 (N_693,In_385,In_552);
and U694 (N_694,In_927,In_269);
or U695 (N_695,In_828,In_268);
xor U696 (N_696,In_1774,In_98);
nand U697 (N_697,In_1360,In_1934);
nor U698 (N_698,In_1455,In_1083);
nor U699 (N_699,In_1965,In_1623);
nor U700 (N_700,In_190,In_1946);
nor U701 (N_701,In_853,In_183);
nand U702 (N_702,In_563,In_604);
nand U703 (N_703,In_1994,In_550);
xnor U704 (N_704,In_1332,In_1026);
nand U705 (N_705,In_922,In_38);
xor U706 (N_706,In_832,In_317);
nand U707 (N_707,In_1311,In_716);
nor U708 (N_708,In_1471,In_1520);
nand U709 (N_709,In_222,In_1852);
and U710 (N_710,In_1487,In_684);
nand U711 (N_711,In_419,In_1226);
and U712 (N_712,In_1368,In_1457);
and U713 (N_713,In_213,In_1850);
and U714 (N_714,In_1006,In_91);
or U715 (N_715,In_1912,In_1737);
nor U716 (N_716,In_1632,In_447);
nor U717 (N_717,In_1537,In_299);
nand U718 (N_718,In_1599,In_993);
nand U719 (N_719,In_437,In_923);
nand U720 (N_720,In_1303,In_1794);
or U721 (N_721,In_1354,In_456);
or U722 (N_722,In_1339,In_1185);
nor U723 (N_723,In_1706,In_1565);
and U724 (N_724,In_1999,In_634);
nand U725 (N_725,In_285,In_1204);
nor U726 (N_726,In_375,In_926);
and U727 (N_727,In_1484,In_751);
and U728 (N_728,In_1041,In_521);
and U729 (N_729,In_1364,In_475);
nand U730 (N_730,In_318,In_1071);
nand U731 (N_731,In_131,In_287);
and U732 (N_732,In_1433,In_773);
nor U733 (N_733,In_1403,In_610);
nand U734 (N_734,In_1547,In_1252);
and U735 (N_735,In_1703,In_812);
and U736 (N_736,In_1862,In_881);
and U737 (N_737,In_1109,In_1081);
xnor U738 (N_738,In_642,In_897);
or U739 (N_739,In_884,In_1495);
nand U740 (N_740,In_303,In_412);
xnor U741 (N_741,In_714,In_443);
or U742 (N_742,In_861,In_1141);
or U743 (N_743,In_511,In_337);
nor U744 (N_744,In_527,In_1441);
or U745 (N_745,In_366,In_530);
and U746 (N_746,In_291,In_918);
nor U747 (N_747,In_106,In_175);
nor U748 (N_748,In_1970,In_912);
nand U749 (N_749,In_2,In_181);
or U750 (N_750,In_1687,In_872);
nand U751 (N_751,In_992,In_1979);
nor U752 (N_752,In_594,In_1192);
nor U753 (N_753,In_350,In_251);
nor U754 (N_754,In_54,In_123);
nand U755 (N_755,In_561,In_1777);
nor U756 (N_756,In_390,In_1350);
or U757 (N_757,In_1824,In_1908);
nand U758 (N_758,In_141,In_1671);
nand U759 (N_759,In_392,In_42);
nand U760 (N_760,In_1150,In_1884);
or U761 (N_761,In_1102,In_1914);
or U762 (N_762,In_1207,In_225);
or U763 (N_763,In_1395,In_66);
and U764 (N_764,In_288,In_466);
and U765 (N_765,In_31,In_1321);
xnor U766 (N_766,In_788,In_822);
nor U767 (N_767,In_518,In_582);
or U768 (N_768,In_400,In_1193);
and U769 (N_769,In_1620,In_1035);
xor U770 (N_770,In_1684,In_1609);
nor U771 (N_771,In_1563,In_84);
nor U772 (N_772,In_498,In_981);
and U773 (N_773,In_1840,In_1700);
nor U774 (N_774,In_1586,In_1848);
or U775 (N_775,In_1717,In_1158);
and U776 (N_776,In_1367,In_161);
nor U777 (N_777,In_675,In_1964);
or U778 (N_778,In_1697,In_1973);
xnor U779 (N_779,In_1661,In_237);
or U780 (N_780,In_1278,In_562);
or U781 (N_781,In_1140,In_138);
nor U782 (N_782,In_983,In_146);
or U783 (N_783,In_1922,In_551);
or U784 (N_784,In_1216,In_980);
and U785 (N_785,In_800,In_276);
nand U786 (N_786,In_1483,In_794);
nor U787 (N_787,In_1903,In_1272);
or U788 (N_788,In_1521,In_1196);
and U789 (N_789,In_1566,In_1108);
and U790 (N_790,In_679,In_309);
and U791 (N_791,In_633,In_1815);
or U792 (N_792,In_187,In_1541);
xor U793 (N_793,In_361,In_1650);
or U794 (N_794,In_379,In_668);
nor U795 (N_795,In_946,In_1410);
and U796 (N_796,In_836,In_120);
nand U797 (N_797,In_1030,In_191);
and U798 (N_798,In_1735,In_405);
nor U799 (N_799,In_619,In_1098);
nand U800 (N_800,In_232,In_102);
or U801 (N_801,In_1839,In_979);
nor U802 (N_802,In_1896,In_1719);
or U803 (N_803,In_821,In_373);
xor U804 (N_804,In_1726,In_1795);
and U805 (N_805,In_1552,In_1825);
and U806 (N_806,In_283,In_436);
nand U807 (N_807,In_47,In_833);
nand U808 (N_808,In_953,In_113);
nand U809 (N_809,In_766,In_723);
nor U810 (N_810,In_281,In_531);
nor U811 (N_811,In_159,In_163);
and U812 (N_812,In_978,In_1681);
nand U813 (N_813,In_1835,In_145);
nand U814 (N_814,In_1061,In_680);
nor U815 (N_815,In_1954,In_1019);
nand U816 (N_816,In_1947,In_1891);
or U817 (N_817,In_1373,In_1577);
nand U818 (N_818,In_467,In_1209);
and U819 (N_819,In_1836,In_1995);
and U820 (N_820,In_1351,In_500);
or U821 (N_821,In_1524,In_472);
nand U822 (N_822,In_1243,In_250);
xnor U823 (N_823,In_1347,In_621);
or U824 (N_824,In_1465,In_226);
nor U825 (N_825,In_1826,In_1277);
nor U826 (N_826,In_188,In_512);
xnor U827 (N_827,In_445,In_1951);
nand U828 (N_828,In_580,In_1549);
or U829 (N_829,In_1324,In_23);
nor U830 (N_830,In_1889,In_444);
or U831 (N_831,In_1508,In_64);
nor U832 (N_832,In_152,In_1626);
nor U833 (N_833,In_242,In_394);
nor U834 (N_834,In_674,In_92);
xnor U835 (N_835,In_1392,In_827);
nor U836 (N_836,In_704,In_792);
nand U837 (N_837,In_639,In_423);
xor U838 (N_838,In_1929,In_386);
and U839 (N_839,In_635,In_541);
nor U840 (N_840,In_1926,In_1305);
nand U841 (N_841,In_1355,In_1290);
nor U842 (N_842,In_1629,In_1203);
nand U843 (N_843,In_1788,In_439);
and U844 (N_844,In_1391,In_1948);
nor U845 (N_845,In_615,In_1406);
or U846 (N_846,In_1635,In_801);
xnor U847 (N_847,In_1452,In_1359);
nand U848 (N_848,In_1446,In_1480);
nand U849 (N_849,In_1168,In_1905);
and U850 (N_850,In_1459,In_297);
nand U851 (N_851,In_1790,In_1530);
and U852 (N_852,In_1846,In_1576);
nand U853 (N_853,In_1147,In_1163);
or U854 (N_854,In_839,In_1734);
or U855 (N_855,In_851,In_549);
nand U856 (N_856,In_68,In_1992);
nor U857 (N_857,In_192,In_369);
nand U858 (N_858,In_1309,In_1819);
or U859 (N_859,In_1211,In_681);
and U860 (N_860,In_595,In_53);
and U861 (N_861,In_1718,In_1174);
nand U862 (N_862,In_663,In_1080);
xor U863 (N_863,In_1334,In_1096);
nor U864 (N_864,In_147,In_1691);
nand U865 (N_865,In_1178,In_898);
or U866 (N_866,In_332,In_1709);
or U867 (N_867,In_676,In_834);
or U868 (N_868,In_996,In_1365);
or U869 (N_869,In_37,In_109);
nor U870 (N_870,In_671,In_1991);
and U871 (N_871,In_955,In_1329);
nor U872 (N_872,In_1641,In_982);
xor U873 (N_873,In_298,In_331);
nand U874 (N_874,In_1381,In_81);
nor U875 (N_875,In_1782,In_1690);
and U876 (N_876,In_841,In_1115);
nor U877 (N_877,In_764,In_360);
nand U878 (N_878,In_1898,In_1640);
and U879 (N_879,In_1990,In_587);
nor U880 (N_880,In_282,In_1761);
or U881 (N_881,In_50,In_165);
nand U882 (N_882,In_1551,In_1811);
and U883 (N_883,In_1887,In_481);
nand U884 (N_884,In_1822,In_1974);
or U885 (N_885,In_933,In_757);
or U886 (N_886,In_114,In_845);
or U887 (N_887,In_395,In_1582);
and U888 (N_888,In_1793,In_1536);
or U889 (N_889,In_693,In_1817);
or U890 (N_890,In_1014,In_969);
nor U891 (N_891,In_1233,In_1304);
or U892 (N_892,In_842,In_528);
and U893 (N_893,In_1225,In_1590);
nand U894 (N_894,In_814,In_702);
nand U895 (N_895,In_1074,In_1945);
xnor U896 (N_896,In_523,In_934);
xnor U897 (N_897,In_484,In_459);
or U898 (N_898,In_892,In_1666);
nand U899 (N_899,In_44,In_1346);
and U900 (N_900,In_1165,In_263);
and U901 (N_901,In_233,In_611);
nand U902 (N_902,In_1519,In_1742);
nand U903 (N_903,In_1024,In_1198);
or U904 (N_904,In_1425,In_470);
and U905 (N_905,In_844,In_1298);
nor U906 (N_906,In_1814,In_1261);
nor U907 (N_907,In_1642,In_489);
xor U908 (N_908,In_586,In_677);
nand U909 (N_909,In_1399,In_1983);
xnor U910 (N_910,In_1371,In_650);
nand U911 (N_911,In_887,In_875);
and U912 (N_912,In_1797,In_900);
nor U913 (N_913,In_1057,In_789);
nor U914 (N_914,In_344,In_627);
nor U915 (N_915,In_338,In_86);
nor U916 (N_916,In_1647,In_249);
or U917 (N_917,In_869,In_315);
and U918 (N_918,In_198,In_391);
or U919 (N_919,In_1136,In_711);
and U920 (N_920,In_767,In_1106);
nor U921 (N_921,In_491,In_1554);
nand U922 (N_922,In_1727,In_430);
nand U923 (N_923,In_1308,In_1336);
nand U924 (N_924,In_740,In_1569);
nand U925 (N_925,In_13,In_590);
xnor U926 (N_926,In_691,In_1637);
or U927 (N_927,In_1985,In_1773);
and U928 (N_928,In_1587,In_1476);
or U929 (N_929,In_1319,In_870);
nor U930 (N_930,In_986,In_36);
and U931 (N_931,In_1539,In_1212);
xnor U932 (N_932,In_65,In_1833);
and U933 (N_933,In_710,In_1923);
nand U934 (N_934,In_1663,In_732);
xor U935 (N_935,In_678,In_685);
nand U936 (N_936,In_837,In_403);
nor U937 (N_937,In_1851,In_1538);
nor U938 (N_938,In_1769,In_1675);
or U939 (N_939,In_1482,In_1445);
and U940 (N_940,In_1422,In_411);
and U941 (N_941,In_14,In_683);
nand U942 (N_942,In_204,In_1497);
xor U943 (N_943,In_560,In_1485);
nand U944 (N_944,In_1134,In_234);
nor U945 (N_945,In_1897,In_1078);
and U946 (N_946,In_324,In_78);
nor U947 (N_947,In_18,In_1741);
nor U948 (N_948,In_525,In_772);
nand U949 (N_949,In_229,In_1377);
or U950 (N_950,In_719,In_1686);
nor U951 (N_951,In_1831,In_591);
nor U952 (N_952,In_69,In_46);
nand U953 (N_953,In_689,In_1791);
nor U954 (N_954,In_1540,In_1892);
or U955 (N_955,In_1601,In_295);
nand U956 (N_956,In_12,In_292);
xor U957 (N_957,In_1968,In_1893);
or U958 (N_958,In_805,In_241);
or U959 (N_959,In_816,In_75);
nor U960 (N_960,In_696,In_1478);
or U961 (N_961,In_866,In_1545);
nand U962 (N_962,In_170,In_1910);
and U963 (N_963,In_921,In_35);
nor U964 (N_964,In_157,In_1702);
nand U965 (N_965,In_363,In_1013);
nor U966 (N_966,In_1200,In_1357);
nor U967 (N_967,In_1804,In_265);
nor U968 (N_968,In_41,In_1612);
xor U969 (N_969,In_196,In_1574);
and U970 (N_970,In_1724,In_637);
and U971 (N_971,In_667,In_235);
nand U972 (N_972,In_1133,In_1714);
and U973 (N_973,In_1448,In_70);
or U974 (N_974,In_294,In_1295);
nor U975 (N_975,In_1559,In_1004);
nand U976 (N_976,In_1598,In_1579);
nor U977 (N_977,In_471,In_1328);
nor U978 (N_978,In_947,In_284);
xor U979 (N_979,In_976,In_17);
nand U980 (N_980,In_760,In_274);
nand U981 (N_981,In_1854,In_1384);
and U982 (N_982,In_10,In_1221);
nor U983 (N_983,In_568,In_358);
or U984 (N_984,In_399,In_270);
nor U985 (N_985,In_1589,In_1564);
or U986 (N_986,In_1993,In_82);
and U987 (N_987,In_8,In_1987);
nand U988 (N_988,In_1971,In_388);
nor U989 (N_989,In_848,In_1958);
or U990 (N_990,In_1527,In_1475);
nand U991 (N_991,In_1664,In_1807);
nand U992 (N_992,In_522,In_1858);
nand U993 (N_993,In_967,In_1879);
nand U994 (N_994,In_700,In_1771);
nor U995 (N_995,In_19,In_1151);
nand U996 (N_996,In_1901,In_1960);
nor U997 (N_997,In_1088,In_1060);
xor U998 (N_998,In_1279,In_1122);
and U999 (N_999,In_340,In_966);
and U1000 (N_1000,In_1359,In_1274);
xor U1001 (N_1001,In_1648,In_170);
nor U1002 (N_1002,In_993,In_1838);
nor U1003 (N_1003,In_1343,In_208);
nand U1004 (N_1004,In_825,In_1631);
or U1005 (N_1005,In_1608,In_405);
or U1006 (N_1006,In_301,In_735);
xor U1007 (N_1007,In_155,In_1361);
nand U1008 (N_1008,In_821,In_746);
nor U1009 (N_1009,In_967,In_1512);
nand U1010 (N_1010,In_396,In_1803);
nor U1011 (N_1011,In_798,In_1144);
xor U1012 (N_1012,In_1412,In_503);
or U1013 (N_1013,In_1607,In_130);
and U1014 (N_1014,In_413,In_176);
xnor U1015 (N_1015,In_175,In_1177);
and U1016 (N_1016,In_1280,In_760);
nand U1017 (N_1017,In_479,In_1441);
nor U1018 (N_1018,In_352,In_1009);
nand U1019 (N_1019,In_332,In_1736);
nand U1020 (N_1020,In_625,In_1889);
or U1021 (N_1021,In_52,In_320);
or U1022 (N_1022,In_1586,In_1823);
xor U1023 (N_1023,In_503,In_1344);
or U1024 (N_1024,In_952,In_1836);
or U1025 (N_1025,In_1449,In_268);
or U1026 (N_1026,In_504,In_399);
nor U1027 (N_1027,In_1337,In_754);
and U1028 (N_1028,In_1275,In_690);
nor U1029 (N_1029,In_1543,In_506);
or U1030 (N_1030,In_1422,In_1704);
xnor U1031 (N_1031,In_446,In_739);
nand U1032 (N_1032,In_236,In_439);
nand U1033 (N_1033,In_1277,In_800);
nor U1034 (N_1034,In_931,In_334);
and U1035 (N_1035,In_810,In_847);
nand U1036 (N_1036,In_1729,In_1479);
and U1037 (N_1037,In_424,In_789);
nor U1038 (N_1038,In_432,In_212);
nand U1039 (N_1039,In_1154,In_521);
nand U1040 (N_1040,In_1720,In_8);
nor U1041 (N_1041,In_1451,In_848);
nand U1042 (N_1042,In_1288,In_1046);
xnor U1043 (N_1043,In_1081,In_1931);
or U1044 (N_1044,In_525,In_321);
xor U1045 (N_1045,In_108,In_720);
or U1046 (N_1046,In_188,In_503);
and U1047 (N_1047,In_1627,In_825);
and U1048 (N_1048,In_1850,In_1208);
or U1049 (N_1049,In_1542,In_1646);
and U1050 (N_1050,In_779,In_1283);
nor U1051 (N_1051,In_1567,In_727);
nor U1052 (N_1052,In_1717,In_668);
or U1053 (N_1053,In_1509,In_949);
or U1054 (N_1054,In_820,In_598);
or U1055 (N_1055,In_1855,In_897);
and U1056 (N_1056,In_956,In_1077);
and U1057 (N_1057,In_1902,In_1584);
nand U1058 (N_1058,In_115,In_1708);
or U1059 (N_1059,In_448,In_1905);
or U1060 (N_1060,In_1493,In_1471);
and U1061 (N_1061,In_1727,In_1788);
or U1062 (N_1062,In_1460,In_156);
and U1063 (N_1063,In_1081,In_1843);
or U1064 (N_1064,In_468,In_949);
or U1065 (N_1065,In_210,In_1806);
or U1066 (N_1066,In_149,In_1941);
nor U1067 (N_1067,In_401,In_1049);
xor U1068 (N_1068,In_834,In_311);
nand U1069 (N_1069,In_1768,In_1163);
and U1070 (N_1070,In_1805,In_862);
nor U1071 (N_1071,In_1273,In_1837);
or U1072 (N_1072,In_1641,In_495);
xor U1073 (N_1073,In_240,In_1766);
nand U1074 (N_1074,In_428,In_1487);
and U1075 (N_1075,In_1923,In_714);
and U1076 (N_1076,In_121,In_212);
nor U1077 (N_1077,In_1866,In_1619);
xnor U1078 (N_1078,In_345,In_118);
xnor U1079 (N_1079,In_703,In_1016);
and U1080 (N_1080,In_555,In_1483);
or U1081 (N_1081,In_1665,In_1914);
nor U1082 (N_1082,In_33,In_1695);
nor U1083 (N_1083,In_454,In_973);
or U1084 (N_1084,In_130,In_1368);
or U1085 (N_1085,In_495,In_249);
xnor U1086 (N_1086,In_1201,In_902);
and U1087 (N_1087,In_803,In_317);
nor U1088 (N_1088,In_492,In_1127);
and U1089 (N_1089,In_1946,In_950);
or U1090 (N_1090,In_1602,In_1144);
or U1091 (N_1091,In_765,In_1826);
nand U1092 (N_1092,In_356,In_376);
or U1093 (N_1093,In_511,In_206);
xor U1094 (N_1094,In_1363,In_1839);
nand U1095 (N_1095,In_614,In_712);
nand U1096 (N_1096,In_230,In_827);
and U1097 (N_1097,In_1533,In_1710);
and U1098 (N_1098,In_1001,In_597);
nand U1099 (N_1099,In_1934,In_503);
xor U1100 (N_1100,In_503,In_343);
or U1101 (N_1101,In_317,In_1602);
xnor U1102 (N_1102,In_407,In_1555);
or U1103 (N_1103,In_680,In_1041);
or U1104 (N_1104,In_801,In_1440);
xnor U1105 (N_1105,In_1754,In_498);
nor U1106 (N_1106,In_957,In_961);
nand U1107 (N_1107,In_152,In_193);
or U1108 (N_1108,In_597,In_1279);
nor U1109 (N_1109,In_155,In_1704);
or U1110 (N_1110,In_122,In_60);
or U1111 (N_1111,In_1798,In_1362);
nor U1112 (N_1112,In_176,In_281);
and U1113 (N_1113,In_152,In_471);
nand U1114 (N_1114,In_900,In_391);
nand U1115 (N_1115,In_1563,In_224);
and U1116 (N_1116,In_885,In_576);
or U1117 (N_1117,In_531,In_563);
and U1118 (N_1118,In_1990,In_1292);
nand U1119 (N_1119,In_967,In_1152);
nor U1120 (N_1120,In_941,In_1564);
and U1121 (N_1121,In_1420,In_822);
nor U1122 (N_1122,In_1226,In_1906);
or U1123 (N_1123,In_425,In_1305);
and U1124 (N_1124,In_1264,In_582);
nor U1125 (N_1125,In_1753,In_592);
nand U1126 (N_1126,In_897,In_726);
nand U1127 (N_1127,In_797,In_1063);
nand U1128 (N_1128,In_441,In_872);
nor U1129 (N_1129,In_1985,In_1721);
xor U1130 (N_1130,In_1651,In_1743);
nor U1131 (N_1131,In_1606,In_1054);
or U1132 (N_1132,In_1323,In_888);
nor U1133 (N_1133,In_35,In_330);
or U1134 (N_1134,In_426,In_83);
nand U1135 (N_1135,In_280,In_1546);
and U1136 (N_1136,In_442,In_1164);
and U1137 (N_1137,In_1181,In_73);
nor U1138 (N_1138,In_90,In_1159);
nand U1139 (N_1139,In_1608,In_172);
nor U1140 (N_1140,In_47,In_1366);
nand U1141 (N_1141,In_209,In_638);
or U1142 (N_1142,In_862,In_1845);
nand U1143 (N_1143,In_1825,In_1353);
nand U1144 (N_1144,In_1874,In_449);
or U1145 (N_1145,In_1233,In_748);
and U1146 (N_1146,In_1916,In_184);
xnor U1147 (N_1147,In_1062,In_1965);
nand U1148 (N_1148,In_915,In_256);
nand U1149 (N_1149,In_1445,In_629);
nor U1150 (N_1150,In_1269,In_1197);
and U1151 (N_1151,In_1236,In_20);
or U1152 (N_1152,In_1754,In_1968);
nor U1153 (N_1153,In_1740,In_1363);
or U1154 (N_1154,In_837,In_1482);
nor U1155 (N_1155,In_1910,In_398);
or U1156 (N_1156,In_1204,In_1863);
or U1157 (N_1157,In_268,In_977);
nand U1158 (N_1158,In_1609,In_704);
nor U1159 (N_1159,In_1005,In_1243);
nand U1160 (N_1160,In_353,In_990);
nand U1161 (N_1161,In_646,In_1571);
or U1162 (N_1162,In_362,In_759);
or U1163 (N_1163,In_236,In_1371);
nor U1164 (N_1164,In_426,In_1400);
or U1165 (N_1165,In_1216,In_549);
nor U1166 (N_1166,In_1920,In_118);
nor U1167 (N_1167,In_1177,In_1180);
or U1168 (N_1168,In_480,In_543);
nor U1169 (N_1169,In_1108,In_460);
nand U1170 (N_1170,In_1968,In_1736);
and U1171 (N_1171,In_774,In_1942);
or U1172 (N_1172,In_1830,In_1595);
and U1173 (N_1173,In_552,In_792);
xnor U1174 (N_1174,In_549,In_264);
and U1175 (N_1175,In_1684,In_1492);
nand U1176 (N_1176,In_908,In_223);
xor U1177 (N_1177,In_685,In_888);
nor U1178 (N_1178,In_910,In_1343);
xnor U1179 (N_1179,In_223,In_505);
or U1180 (N_1180,In_1907,In_1034);
and U1181 (N_1181,In_1508,In_396);
xnor U1182 (N_1182,In_1302,In_459);
and U1183 (N_1183,In_1948,In_338);
and U1184 (N_1184,In_306,In_1433);
nand U1185 (N_1185,In_44,In_1624);
or U1186 (N_1186,In_114,In_1166);
nand U1187 (N_1187,In_284,In_869);
and U1188 (N_1188,In_621,In_1985);
or U1189 (N_1189,In_1967,In_1880);
or U1190 (N_1190,In_256,In_559);
xnor U1191 (N_1191,In_67,In_206);
nor U1192 (N_1192,In_1101,In_517);
nor U1193 (N_1193,In_1929,In_1603);
nand U1194 (N_1194,In_805,In_539);
nand U1195 (N_1195,In_1345,In_1998);
xnor U1196 (N_1196,In_1299,In_549);
and U1197 (N_1197,In_778,In_336);
nor U1198 (N_1198,In_847,In_72);
nand U1199 (N_1199,In_1477,In_1147);
and U1200 (N_1200,In_947,In_201);
nor U1201 (N_1201,In_682,In_1513);
xor U1202 (N_1202,In_1250,In_1493);
and U1203 (N_1203,In_1444,In_1595);
or U1204 (N_1204,In_255,In_1827);
nand U1205 (N_1205,In_1237,In_1404);
nand U1206 (N_1206,In_613,In_1402);
nand U1207 (N_1207,In_266,In_780);
nor U1208 (N_1208,In_105,In_287);
nor U1209 (N_1209,In_171,In_1357);
nor U1210 (N_1210,In_1040,In_1313);
or U1211 (N_1211,In_351,In_1010);
or U1212 (N_1212,In_584,In_1723);
nor U1213 (N_1213,In_156,In_1869);
xnor U1214 (N_1214,In_1233,In_1584);
or U1215 (N_1215,In_476,In_625);
or U1216 (N_1216,In_1743,In_108);
and U1217 (N_1217,In_1817,In_1469);
xor U1218 (N_1218,In_1252,In_1307);
nor U1219 (N_1219,In_318,In_1409);
nand U1220 (N_1220,In_931,In_1079);
or U1221 (N_1221,In_965,In_1151);
nor U1222 (N_1222,In_1147,In_1463);
nor U1223 (N_1223,In_154,In_56);
or U1224 (N_1224,In_76,In_708);
or U1225 (N_1225,In_960,In_1693);
or U1226 (N_1226,In_546,In_1782);
nor U1227 (N_1227,In_255,In_1525);
or U1228 (N_1228,In_305,In_1968);
xnor U1229 (N_1229,In_1508,In_1970);
and U1230 (N_1230,In_311,In_693);
nand U1231 (N_1231,In_1044,In_418);
and U1232 (N_1232,In_1782,In_1615);
or U1233 (N_1233,In_671,In_949);
and U1234 (N_1234,In_1940,In_1646);
or U1235 (N_1235,In_71,In_1884);
and U1236 (N_1236,In_181,In_1580);
and U1237 (N_1237,In_584,In_1583);
and U1238 (N_1238,In_1318,In_1985);
nor U1239 (N_1239,In_1674,In_1316);
xnor U1240 (N_1240,In_773,In_1839);
or U1241 (N_1241,In_1076,In_183);
nor U1242 (N_1242,In_279,In_251);
and U1243 (N_1243,In_446,In_1575);
or U1244 (N_1244,In_1438,In_1347);
or U1245 (N_1245,In_511,In_293);
nand U1246 (N_1246,In_1984,In_1474);
and U1247 (N_1247,In_1675,In_1639);
or U1248 (N_1248,In_473,In_529);
or U1249 (N_1249,In_1234,In_791);
nand U1250 (N_1250,In_318,In_390);
nand U1251 (N_1251,In_1645,In_902);
nor U1252 (N_1252,In_757,In_181);
or U1253 (N_1253,In_913,In_554);
nor U1254 (N_1254,In_720,In_438);
or U1255 (N_1255,In_1545,In_1252);
and U1256 (N_1256,In_1734,In_1244);
and U1257 (N_1257,In_56,In_1466);
nand U1258 (N_1258,In_1059,In_464);
xor U1259 (N_1259,In_658,In_1804);
xnor U1260 (N_1260,In_1781,In_1872);
or U1261 (N_1261,In_1439,In_1795);
nor U1262 (N_1262,In_175,In_1266);
or U1263 (N_1263,In_302,In_1072);
nand U1264 (N_1264,In_1995,In_830);
and U1265 (N_1265,In_1805,In_438);
and U1266 (N_1266,In_1076,In_1717);
or U1267 (N_1267,In_121,In_1658);
nand U1268 (N_1268,In_1412,In_51);
and U1269 (N_1269,In_692,In_88);
nor U1270 (N_1270,In_424,In_1523);
nor U1271 (N_1271,In_5,In_905);
or U1272 (N_1272,In_1303,In_1015);
nand U1273 (N_1273,In_1086,In_1089);
xnor U1274 (N_1274,In_1643,In_564);
nand U1275 (N_1275,In_574,In_1978);
or U1276 (N_1276,In_1159,In_1418);
nor U1277 (N_1277,In_879,In_792);
xnor U1278 (N_1278,In_1478,In_765);
nand U1279 (N_1279,In_1858,In_383);
nor U1280 (N_1280,In_1345,In_677);
nor U1281 (N_1281,In_797,In_812);
nor U1282 (N_1282,In_431,In_405);
nor U1283 (N_1283,In_1603,In_1549);
and U1284 (N_1284,In_838,In_949);
or U1285 (N_1285,In_810,In_645);
or U1286 (N_1286,In_632,In_1740);
or U1287 (N_1287,In_284,In_375);
and U1288 (N_1288,In_1173,In_1370);
or U1289 (N_1289,In_150,In_565);
or U1290 (N_1290,In_1874,In_1621);
and U1291 (N_1291,In_1523,In_871);
nand U1292 (N_1292,In_1550,In_437);
nor U1293 (N_1293,In_671,In_565);
or U1294 (N_1294,In_1059,In_1332);
nor U1295 (N_1295,In_483,In_1502);
or U1296 (N_1296,In_869,In_1355);
or U1297 (N_1297,In_730,In_704);
and U1298 (N_1298,In_1428,In_1477);
nor U1299 (N_1299,In_1636,In_362);
and U1300 (N_1300,In_521,In_466);
nand U1301 (N_1301,In_910,In_216);
or U1302 (N_1302,In_1380,In_1604);
and U1303 (N_1303,In_799,In_1790);
nor U1304 (N_1304,In_426,In_262);
or U1305 (N_1305,In_302,In_1946);
nor U1306 (N_1306,In_1632,In_493);
nand U1307 (N_1307,In_439,In_1460);
nand U1308 (N_1308,In_1889,In_687);
nand U1309 (N_1309,In_714,In_882);
nand U1310 (N_1310,In_1877,In_606);
or U1311 (N_1311,In_396,In_579);
and U1312 (N_1312,In_681,In_412);
xnor U1313 (N_1313,In_1929,In_952);
nor U1314 (N_1314,In_977,In_1416);
and U1315 (N_1315,In_789,In_66);
and U1316 (N_1316,In_1603,In_1948);
or U1317 (N_1317,In_888,In_1097);
or U1318 (N_1318,In_1852,In_1293);
xor U1319 (N_1319,In_994,In_131);
nor U1320 (N_1320,In_355,In_936);
and U1321 (N_1321,In_893,In_1865);
nor U1322 (N_1322,In_1266,In_295);
or U1323 (N_1323,In_1799,In_175);
nand U1324 (N_1324,In_1090,In_83);
or U1325 (N_1325,In_543,In_829);
nand U1326 (N_1326,In_313,In_40);
nor U1327 (N_1327,In_483,In_1362);
xor U1328 (N_1328,In_1085,In_292);
nand U1329 (N_1329,In_50,In_1974);
nand U1330 (N_1330,In_1427,In_670);
or U1331 (N_1331,In_297,In_240);
or U1332 (N_1332,In_1178,In_937);
nand U1333 (N_1333,In_499,In_653);
or U1334 (N_1334,In_1222,In_1601);
or U1335 (N_1335,In_978,In_920);
nor U1336 (N_1336,In_791,In_1551);
and U1337 (N_1337,In_1886,In_724);
and U1338 (N_1338,In_870,In_674);
or U1339 (N_1339,In_594,In_430);
or U1340 (N_1340,In_995,In_96);
nand U1341 (N_1341,In_662,In_1419);
or U1342 (N_1342,In_275,In_1694);
nor U1343 (N_1343,In_1861,In_643);
and U1344 (N_1344,In_1001,In_929);
nor U1345 (N_1345,In_469,In_491);
and U1346 (N_1346,In_865,In_1653);
nand U1347 (N_1347,In_1443,In_1711);
nand U1348 (N_1348,In_759,In_267);
or U1349 (N_1349,In_1019,In_1379);
nor U1350 (N_1350,In_1228,In_1837);
nor U1351 (N_1351,In_988,In_921);
xor U1352 (N_1352,In_1920,In_1782);
and U1353 (N_1353,In_1698,In_25);
nand U1354 (N_1354,In_1694,In_1963);
and U1355 (N_1355,In_898,In_815);
or U1356 (N_1356,In_1642,In_778);
and U1357 (N_1357,In_5,In_1758);
or U1358 (N_1358,In_1539,In_141);
nand U1359 (N_1359,In_1075,In_1939);
nand U1360 (N_1360,In_700,In_116);
nand U1361 (N_1361,In_717,In_1006);
or U1362 (N_1362,In_1167,In_356);
nor U1363 (N_1363,In_1943,In_1964);
and U1364 (N_1364,In_1920,In_672);
or U1365 (N_1365,In_1811,In_42);
xor U1366 (N_1366,In_1289,In_1346);
nand U1367 (N_1367,In_1606,In_1127);
or U1368 (N_1368,In_1887,In_339);
nand U1369 (N_1369,In_475,In_1483);
or U1370 (N_1370,In_357,In_132);
nand U1371 (N_1371,In_328,In_269);
nand U1372 (N_1372,In_1943,In_124);
or U1373 (N_1373,In_696,In_1479);
and U1374 (N_1374,In_680,In_245);
xnor U1375 (N_1375,In_159,In_75);
or U1376 (N_1376,In_1069,In_599);
and U1377 (N_1377,In_188,In_1486);
nor U1378 (N_1378,In_207,In_1344);
xor U1379 (N_1379,In_1738,In_576);
and U1380 (N_1380,In_1642,In_1972);
nor U1381 (N_1381,In_38,In_1526);
and U1382 (N_1382,In_738,In_635);
xor U1383 (N_1383,In_1264,In_1758);
nand U1384 (N_1384,In_1972,In_1065);
xnor U1385 (N_1385,In_1619,In_1902);
nand U1386 (N_1386,In_102,In_1549);
and U1387 (N_1387,In_1082,In_66);
or U1388 (N_1388,In_1021,In_1055);
and U1389 (N_1389,In_921,In_807);
and U1390 (N_1390,In_957,In_1342);
nand U1391 (N_1391,In_343,In_798);
nor U1392 (N_1392,In_439,In_1135);
and U1393 (N_1393,In_444,In_1993);
or U1394 (N_1394,In_1830,In_1373);
nand U1395 (N_1395,In_1322,In_288);
nand U1396 (N_1396,In_922,In_1802);
nor U1397 (N_1397,In_921,In_1519);
or U1398 (N_1398,In_879,In_973);
or U1399 (N_1399,In_732,In_677);
nand U1400 (N_1400,In_796,In_111);
and U1401 (N_1401,In_1534,In_33);
or U1402 (N_1402,In_1905,In_348);
and U1403 (N_1403,In_1751,In_315);
nand U1404 (N_1404,In_1782,In_1851);
and U1405 (N_1405,In_1741,In_223);
or U1406 (N_1406,In_1873,In_375);
nor U1407 (N_1407,In_1139,In_1152);
and U1408 (N_1408,In_1194,In_1091);
nand U1409 (N_1409,In_451,In_1192);
and U1410 (N_1410,In_1076,In_451);
xor U1411 (N_1411,In_489,In_1196);
nor U1412 (N_1412,In_997,In_240);
nand U1413 (N_1413,In_743,In_65);
nand U1414 (N_1414,In_654,In_828);
xor U1415 (N_1415,In_780,In_1884);
nand U1416 (N_1416,In_1918,In_225);
nor U1417 (N_1417,In_1780,In_231);
nand U1418 (N_1418,In_1154,In_1870);
nand U1419 (N_1419,In_1955,In_1526);
nor U1420 (N_1420,In_156,In_157);
nand U1421 (N_1421,In_356,In_626);
and U1422 (N_1422,In_653,In_1480);
or U1423 (N_1423,In_1752,In_1734);
nand U1424 (N_1424,In_514,In_1064);
nor U1425 (N_1425,In_279,In_782);
or U1426 (N_1426,In_1646,In_1134);
or U1427 (N_1427,In_175,In_969);
xnor U1428 (N_1428,In_370,In_316);
or U1429 (N_1429,In_1894,In_1379);
nand U1430 (N_1430,In_43,In_1961);
nor U1431 (N_1431,In_1473,In_37);
nor U1432 (N_1432,In_233,In_266);
or U1433 (N_1433,In_645,In_1943);
nand U1434 (N_1434,In_439,In_1859);
nor U1435 (N_1435,In_885,In_1645);
nand U1436 (N_1436,In_1682,In_246);
nor U1437 (N_1437,In_1090,In_1608);
nor U1438 (N_1438,In_483,In_1026);
nand U1439 (N_1439,In_1492,In_1861);
and U1440 (N_1440,In_470,In_1809);
and U1441 (N_1441,In_552,In_559);
xnor U1442 (N_1442,In_1384,In_642);
nand U1443 (N_1443,In_1812,In_903);
nand U1444 (N_1444,In_20,In_1502);
xnor U1445 (N_1445,In_560,In_1241);
or U1446 (N_1446,In_252,In_61);
nor U1447 (N_1447,In_1710,In_265);
xor U1448 (N_1448,In_1387,In_1860);
xnor U1449 (N_1449,In_1852,In_1723);
xnor U1450 (N_1450,In_1603,In_1820);
nor U1451 (N_1451,In_1129,In_959);
nand U1452 (N_1452,In_160,In_574);
and U1453 (N_1453,In_1228,In_1845);
and U1454 (N_1454,In_527,In_289);
nor U1455 (N_1455,In_1648,In_1975);
nand U1456 (N_1456,In_946,In_1777);
and U1457 (N_1457,In_1151,In_1495);
nand U1458 (N_1458,In_1225,In_75);
nand U1459 (N_1459,In_1740,In_1993);
or U1460 (N_1460,In_626,In_1173);
nor U1461 (N_1461,In_1085,In_1691);
and U1462 (N_1462,In_1591,In_691);
or U1463 (N_1463,In_745,In_929);
or U1464 (N_1464,In_1163,In_945);
and U1465 (N_1465,In_660,In_77);
nor U1466 (N_1466,In_254,In_1835);
xnor U1467 (N_1467,In_1869,In_432);
and U1468 (N_1468,In_1295,In_535);
xor U1469 (N_1469,In_87,In_466);
nor U1470 (N_1470,In_991,In_1861);
xor U1471 (N_1471,In_335,In_1747);
nor U1472 (N_1472,In_906,In_636);
or U1473 (N_1473,In_422,In_1058);
nor U1474 (N_1474,In_1948,In_1813);
or U1475 (N_1475,In_1727,In_548);
nand U1476 (N_1476,In_1892,In_1429);
nand U1477 (N_1477,In_312,In_1765);
and U1478 (N_1478,In_572,In_757);
and U1479 (N_1479,In_719,In_724);
nor U1480 (N_1480,In_713,In_843);
and U1481 (N_1481,In_17,In_1624);
nand U1482 (N_1482,In_1723,In_1306);
nor U1483 (N_1483,In_1469,In_458);
or U1484 (N_1484,In_1631,In_1580);
and U1485 (N_1485,In_830,In_1829);
or U1486 (N_1486,In_758,In_1842);
nor U1487 (N_1487,In_1100,In_1616);
and U1488 (N_1488,In_804,In_1254);
nand U1489 (N_1489,In_951,In_100);
nor U1490 (N_1490,In_1505,In_728);
or U1491 (N_1491,In_847,In_1339);
xor U1492 (N_1492,In_563,In_1130);
nor U1493 (N_1493,In_1617,In_486);
and U1494 (N_1494,In_447,In_407);
and U1495 (N_1495,In_1059,In_731);
or U1496 (N_1496,In_1991,In_1150);
xnor U1497 (N_1497,In_783,In_220);
and U1498 (N_1498,In_39,In_1395);
or U1499 (N_1499,In_668,In_349);
nor U1500 (N_1500,In_122,In_1416);
or U1501 (N_1501,In_1954,In_423);
and U1502 (N_1502,In_1980,In_528);
and U1503 (N_1503,In_319,In_453);
or U1504 (N_1504,In_1999,In_261);
or U1505 (N_1505,In_1157,In_1934);
nor U1506 (N_1506,In_897,In_840);
nor U1507 (N_1507,In_281,In_1730);
xor U1508 (N_1508,In_895,In_1761);
nor U1509 (N_1509,In_1587,In_1094);
xnor U1510 (N_1510,In_1009,In_1681);
nor U1511 (N_1511,In_13,In_507);
nor U1512 (N_1512,In_1175,In_559);
nand U1513 (N_1513,In_1293,In_1593);
and U1514 (N_1514,In_1482,In_748);
nor U1515 (N_1515,In_541,In_1468);
xor U1516 (N_1516,In_955,In_1403);
nand U1517 (N_1517,In_490,In_1425);
and U1518 (N_1518,In_740,In_1810);
nor U1519 (N_1519,In_1752,In_657);
or U1520 (N_1520,In_1495,In_1184);
or U1521 (N_1521,In_1517,In_1054);
and U1522 (N_1522,In_1555,In_974);
nor U1523 (N_1523,In_1326,In_1009);
or U1524 (N_1524,In_1889,In_1115);
or U1525 (N_1525,In_1287,In_1569);
nor U1526 (N_1526,In_560,In_1460);
and U1527 (N_1527,In_1871,In_1295);
nor U1528 (N_1528,In_677,In_1481);
and U1529 (N_1529,In_1448,In_1025);
nand U1530 (N_1530,In_1630,In_1304);
nor U1531 (N_1531,In_246,In_654);
xnor U1532 (N_1532,In_1166,In_323);
and U1533 (N_1533,In_1146,In_1197);
and U1534 (N_1534,In_610,In_1141);
xor U1535 (N_1535,In_821,In_119);
nand U1536 (N_1536,In_698,In_1218);
nand U1537 (N_1537,In_288,In_1548);
and U1538 (N_1538,In_1888,In_1612);
or U1539 (N_1539,In_874,In_395);
and U1540 (N_1540,In_1363,In_1692);
and U1541 (N_1541,In_1993,In_1931);
xnor U1542 (N_1542,In_147,In_1147);
or U1543 (N_1543,In_1105,In_603);
nand U1544 (N_1544,In_1096,In_1791);
nand U1545 (N_1545,In_1156,In_363);
nand U1546 (N_1546,In_381,In_761);
nor U1547 (N_1547,In_1980,In_1971);
nand U1548 (N_1548,In_118,In_1738);
nand U1549 (N_1549,In_278,In_1143);
or U1550 (N_1550,In_1985,In_257);
and U1551 (N_1551,In_1682,In_1355);
or U1552 (N_1552,In_1149,In_981);
and U1553 (N_1553,In_198,In_814);
nand U1554 (N_1554,In_1993,In_774);
nor U1555 (N_1555,In_376,In_801);
nand U1556 (N_1556,In_1162,In_471);
nor U1557 (N_1557,In_1562,In_1419);
or U1558 (N_1558,In_1732,In_879);
and U1559 (N_1559,In_1230,In_1956);
or U1560 (N_1560,In_20,In_1807);
or U1561 (N_1561,In_313,In_775);
and U1562 (N_1562,In_598,In_1726);
and U1563 (N_1563,In_822,In_857);
or U1564 (N_1564,In_1561,In_664);
nor U1565 (N_1565,In_1447,In_1033);
xnor U1566 (N_1566,In_249,In_1724);
and U1567 (N_1567,In_49,In_389);
xor U1568 (N_1568,In_1783,In_141);
and U1569 (N_1569,In_595,In_617);
or U1570 (N_1570,In_868,In_415);
nand U1571 (N_1571,In_1720,In_692);
and U1572 (N_1572,In_935,In_1406);
nand U1573 (N_1573,In_482,In_101);
nor U1574 (N_1574,In_584,In_1923);
and U1575 (N_1575,In_1781,In_713);
nand U1576 (N_1576,In_1326,In_874);
nor U1577 (N_1577,In_155,In_850);
or U1578 (N_1578,In_1468,In_906);
nor U1579 (N_1579,In_1633,In_787);
or U1580 (N_1580,In_1851,In_136);
and U1581 (N_1581,In_585,In_1184);
nor U1582 (N_1582,In_1973,In_903);
xnor U1583 (N_1583,In_279,In_988);
nand U1584 (N_1584,In_1482,In_542);
or U1585 (N_1585,In_0,In_1098);
nand U1586 (N_1586,In_783,In_1697);
nand U1587 (N_1587,In_1092,In_595);
or U1588 (N_1588,In_1595,In_584);
nor U1589 (N_1589,In_531,In_1146);
nand U1590 (N_1590,In_1824,In_304);
or U1591 (N_1591,In_568,In_1029);
nor U1592 (N_1592,In_1996,In_33);
and U1593 (N_1593,In_1128,In_92);
or U1594 (N_1594,In_1466,In_1940);
nor U1595 (N_1595,In_1053,In_1768);
and U1596 (N_1596,In_1536,In_1885);
nor U1597 (N_1597,In_232,In_19);
nor U1598 (N_1598,In_800,In_1363);
nor U1599 (N_1599,In_1451,In_170);
nand U1600 (N_1600,In_1048,In_1817);
nand U1601 (N_1601,In_15,In_1856);
nor U1602 (N_1602,In_1496,In_277);
and U1603 (N_1603,In_1244,In_1605);
or U1604 (N_1604,In_1371,In_1610);
nand U1605 (N_1605,In_1010,In_949);
or U1606 (N_1606,In_215,In_1448);
or U1607 (N_1607,In_890,In_1770);
or U1608 (N_1608,In_1833,In_1791);
or U1609 (N_1609,In_54,In_456);
or U1610 (N_1610,In_641,In_1122);
nor U1611 (N_1611,In_577,In_1508);
and U1612 (N_1612,In_940,In_1143);
or U1613 (N_1613,In_1707,In_1757);
xnor U1614 (N_1614,In_1695,In_1137);
nor U1615 (N_1615,In_1851,In_1728);
and U1616 (N_1616,In_669,In_481);
or U1617 (N_1617,In_1114,In_649);
and U1618 (N_1618,In_62,In_1861);
and U1619 (N_1619,In_1361,In_1566);
nand U1620 (N_1620,In_1044,In_690);
nor U1621 (N_1621,In_1700,In_205);
or U1622 (N_1622,In_589,In_1897);
nand U1623 (N_1623,In_1532,In_1432);
or U1624 (N_1624,In_50,In_1247);
nor U1625 (N_1625,In_1887,In_1037);
xor U1626 (N_1626,In_1779,In_1151);
xor U1627 (N_1627,In_547,In_935);
nor U1628 (N_1628,In_113,In_1379);
and U1629 (N_1629,In_1392,In_734);
xnor U1630 (N_1630,In_699,In_287);
nand U1631 (N_1631,In_630,In_1175);
nand U1632 (N_1632,In_834,In_960);
nor U1633 (N_1633,In_1298,In_1644);
nand U1634 (N_1634,In_1998,In_1660);
or U1635 (N_1635,In_1650,In_1605);
and U1636 (N_1636,In_1986,In_29);
nor U1637 (N_1637,In_452,In_635);
or U1638 (N_1638,In_529,In_840);
nor U1639 (N_1639,In_1066,In_1617);
nand U1640 (N_1640,In_229,In_788);
nand U1641 (N_1641,In_1630,In_823);
nand U1642 (N_1642,In_1238,In_675);
or U1643 (N_1643,In_1120,In_152);
and U1644 (N_1644,In_239,In_745);
xor U1645 (N_1645,In_650,In_722);
and U1646 (N_1646,In_1021,In_1855);
nor U1647 (N_1647,In_1038,In_856);
nand U1648 (N_1648,In_536,In_1937);
or U1649 (N_1649,In_1801,In_200);
nor U1650 (N_1650,In_1544,In_1789);
nor U1651 (N_1651,In_626,In_1159);
nor U1652 (N_1652,In_240,In_1616);
or U1653 (N_1653,In_1578,In_238);
nor U1654 (N_1654,In_166,In_555);
nor U1655 (N_1655,In_109,In_1508);
and U1656 (N_1656,In_274,In_768);
nor U1657 (N_1657,In_270,In_706);
and U1658 (N_1658,In_56,In_599);
or U1659 (N_1659,In_1721,In_690);
nor U1660 (N_1660,In_1083,In_766);
nand U1661 (N_1661,In_9,In_1191);
xor U1662 (N_1662,In_1742,In_1364);
nor U1663 (N_1663,In_1068,In_1862);
or U1664 (N_1664,In_1496,In_1292);
nor U1665 (N_1665,In_1753,In_172);
and U1666 (N_1666,In_569,In_1927);
nor U1667 (N_1667,In_907,In_1454);
nor U1668 (N_1668,In_1567,In_543);
and U1669 (N_1669,In_159,In_1050);
and U1670 (N_1670,In_1992,In_1751);
and U1671 (N_1671,In_1394,In_1302);
and U1672 (N_1672,In_963,In_1789);
nand U1673 (N_1673,In_836,In_744);
xnor U1674 (N_1674,In_374,In_1603);
nand U1675 (N_1675,In_1632,In_1772);
nand U1676 (N_1676,In_1244,In_1653);
xor U1677 (N_1677,In_770,In_381);
or U1678 (N_1678,In_699,In_272);
nand U1679 (N_1679,In_1052,In_403);
nor U1680 (N_1680,In_230,In_26);
and U1681 (N_1681,In_1177,In_1931);
nor U1682 (N_1682,In_561,In_1657);
nor U1683 (N_1683,In_1752,In_29);
nand U1684 (N_1684,In_64,In_1219);
nand U1685 (N_1685,In_1316,In_1588);
or U1686 (N_1686,In_750,In_1474);
or U1687 (N_1687,In_1135,In_964);
or U1688 (N_1688,In_1447,In_987);
nand U1689 (N_1689,In_284,In_180);
and U1690 (N_1690,In_701,In_400);
and U1691 (N_1691,In_340,In_1529);
nand U1692 (N_1692,In_1180,In_702);
or U1693 (N_1693,In_1392,In_465);
and U1694 (N_1694,In_828,In_1356);
and U1695 (N_1695,In_1730,In_1582);
nor U1696 (N_1696,In_255,In_217);
and U1697 (N_1697,In_1004,In_40);
or U1698 (N_1698,In_988,In_1544);
nor U1699 (N_1699,In_172,In_603);
or U1700 (N_1700,In_1990,In_935);
and U1701 (N_1701,In_285,In_1335);
nand U1702 (N_1702,In_945,In_388);
and U1703 (N_1703,In_292,In_0);
nor U1704 (N_1704,In_1004,In_365);
or U1705 (N_1705,In_1958,In_1615);
and U1706 (N_1706,In_176,In_1476);
nor U1707 (N_1707,In_581,In_697);
and U1708 (N_1708,In_992,In_1552);
nand U1709 (N_1709,In_828,In_429);
nor U1710 (N_1710,In_1088,In_1419);
nand U1711 (N_1711,In_1078,In_1991);
or U1712 (N_1712,In_1753,In_327);
nor U1713 (N_1713,In_763,In_717);
and U1714 (N_1714,In_1897,In_1883);
or U1715 (N_1715,In_266,In_258);
and U1716 (N_1716,In_1820,In_1639);
nor U1717 (N_1717,In_1765,In_315);
and U1718 (N_1718,In_228,In_1810);
nor U1719 (N_1719,In_1643,In_1427);
nand U1720 (N_1720,In_1668,In_1742);
nand U1721 (N_1721,In_1083,In_1146);
or U1722 (N_1722,In_1223,In_1640);
or U1723 (N_1723,In_1848,In_657);
or U1724 (N_1724,In_889,In_985);
nor U1725 (N_1725,In_1150,In_1535);
nor U1726 (N_1726,In_505,In_1261);
nor U1727 (N_1727,In_527,In_1302);
or U1728 (N_1728,In_112,In_54);
or U1729 (N_1729,In_1981,In_279);
and U1730 (N_1730,In_554,In_157);
and U1731 (N_1731,In_1950,In_1695);
nor U1732 (N_1732,In_836,In_14);
nor U1733 (N_1733,In_204,In_581);
nor U1734 (N_1734,In_1700,In_789);
or U1735 (N_1735,In_723,In_1665);
and U1736 (N_1736,In_1504,In_1676);
nor U1737 (N_1737,In_1981,In_1609);
nor U1738 (N_1738,In_769,In_343);
nor U1739 (N_1739,In_480,In_436);
nand U1740 (N_1740,In_1110,In_1017);
nand U1741 (N_1741,In_221,In_1345);
nand U1742 (N_1742,In_531,In_1847);
nor U1743 (N_1743,In_1174,In_432);
nand U1744 (N_1744,In_1805,In_694);
nor U1745 (N_1745,In_283,In_1113);
and U1746 (N_1746,In_1057,In_586);
nand U1747 (N_1747,In_1044,In_1396);
nor U1748 (N_1748,In_222,In_120);
nand U1749 (N_1749,In_723,In_1031);
or U1750 (N_1750,In_405,In_521);
or U1751 (N_1751,In_962,In_97);
and U1752 (N_1752,In_991,In_466);
nor U1753 (N_1753,In_1263,In_940);
and U1754 (N_1754,In_1163,In_507);
or U1755 (N_1755,In_1488,In_1909);
nor U1756 (N_1756,In_1498,In_1405);
and U1757 (N_1757,In_1773,In_192);
or U1758 (N_1758,In_1632,In_251);
xor U1759 (N_1759,In_428,In_1328);
nor U1760 (N_1760,In_1031,In_1010);
nand U1761 (N_1761,In_334,In_856);
and U1762 (N_1762,In_1909,In_1368);
and U1763 (N_1763,In_658,In_1103);
and U1764 (N_1764,In_832,In_754);
nor U1765 (N_1765,In_1938,In_579);
nand U1766 (N_1766,In_385,In_836);
xor U1767 (N_1767,In_1916,In_1898);
nand U1768 (N_1768,In_188,In_1229);
or U1769 (N_1769,In_1579,In_800);
nor U1770 (N_1770,In_947,In_1145);
nand U1771 (N_1771,In_1945,In_1320);
or U1772 (N_1772,In_1898,In_457);
or U1773 (N_1773,In_1096,In_1120);
or U1774 (N_1774,In_1917,In_816);
or U1775 (N_1775,In_943,In_888);
or U1776 (N_1776,In_1218,In_1944);
nor U1777 (N_1777,In_805,In_1603);
xor U1778 (N_1778,In_637,In_5);
xnor U1779 (N_1779,In_1271,In_1777);
and U1780 (N_1780,In_1481,In_107);
nor U1781 (N_1781,In_1087,In_1517);
or U1782 (N_1782,In_1230,In_1423);
nor U1783 (N_1783,In_1937,In_1763);
nand U1784 (N_1784,In_1640,In_1454);
nor U1785 (N_1785,In_434,In_729);
and U1786 (N_1786,In_1479,In_1113);
nor U1787 (N_1787,In_850,In_124);
nor U1788 (N_1788,In_307,In_1347);
and U1789 (N_1789,In_34,In_140);
and U1790 (N_1790,In_1426,In_1390);
and U1791 (N_1791,In_1496,In_171);
or U1792 (N_1792,In_1035,In_737);
nand U1793 (N_1793,In_1160,In_1433);
nor U1794 (N_1794,In_1226,In_1913);
nor U1795 (N_1795,In_1434,In_1170);
nor U1796 (N_1796,In_1405,In_353);
nand U1797 (N_1797,In_1907,In_693);
or U1798 (N_1798,In_376,In_1589);
nand U1799 (N_1799,In_985,In_1524);
nor U1800 (N_1800,In_908,In_1501);
or U1801 (N_1801,In_656,In_1418);
xnor U1802 (N_1802,In_1745,In_1689);
or U1803 (N_1803,In_137,In_1075);
and U1804 (N_1804,In_715,In_404);
nor U1805 (N_1805,In_313,In_1738);
nor U1806 (N_1806,In_222,In_292);
nor U1807 (N_1807,In_39,In_1867);
and U1808 (N_1808,In_652,In_861);
nor U1809 (N_1809,In_843,In_703);
and U1810 (N_1810,In_781,In_1008);
and U1811 (N_1811,In_752,In_1245);
and U1812 (N_1812,In_788,In_1939);
and U1813 (N_1813,In_114,In_472);
or U1814 (N_1814,In_1650,In_858);
nor U1815 (N_1815,In_1093,In_927);
or U1816 (N_1816,In_605,In_1367);
nand U1817 (N_1817,In_1316,In_1315);
nor U1818 (N_1818,In_1798,In_121);
xnor U1819 (N_1819,In_651,In_1054);
nor U1820 (N_1820,In_969,In_703);
and U1821 (N_1821,In_330,In_1707);
nand U1822 (N_1822,In_358,In_1139);
and U1823 (N_1823,In_1472,In_523);
or U1824 (N_1824,In_1261,In_594);
and U1825 (N_1825,In_260,In_1551);
xnor U1826 (N_1826,In_838,In_712);
or U1827 (N_1827,In_706,In_72);
xnor U1828 (N_1828,In_831,In_934);
nor U1829 (N_1829,In_628,In_886);
and U1830 (N_1830,In_1723,In_944);
or U1831 (N_1831,In_1694,In_1894);
and U1832 (N_1832,In_744,In_693);
nand U1833 (N_1833,In_1706,In_88);
nor U1834 (N_1834,In_1020,In_1529);
nand U1835 (N_1835,In_1589,In_1838);
or U1836 (N_1836,In_967,In_1103);
nor U1837 (N_1837,In_511,In_1819);
nor U1838 (N_1838,In_1521,In_1567);
and U1839 (N_1839,In_1070,In_1436);
xnor U1840 (N_1840,In_1228,In_752);
or U1841 (N_1841,In_878,In_408);
nor U1842 (N_1842,In_1555,In_912);
or U1843 (N_1843,In_1089,In_1794);
and U1844 (N_1844,In_367,In_1164);
nor U1845 (N_1845,In_981,In_278);
or U1846 (N_1846,In_1353,In_190);
or U1847 (N_1847,In_1691,In_405);
xnor U1848 (N_1848,In_470,In_7);
or U1849 (N_1849,In_1739,In_90);
nor U1850 (N_1850,In_1248,In_1831);
nand U1851 (N_1851,In_283,In_236);
or U1852 (N_1852,In_616,In_859);
and U1853 (N_1853,In_1915,In_385);
and U1854 (N_1854,In_1169,In_113);
nor U1855 (N_1855,In_60,In_93);
nand U1856 (N_1856,In_1306,In_807);
and U1857 (N_1857,In_556,In_1229);
and U1858 (N_1858,In_1735,In_1025);
nor U1859 (N_1859,In_1089,In_124);
nand U1860 (N_1860,In_90,In_955);
or U1861 (N_1861,In_1604,In_340);
nor U1862 (N_1862,In_1013,In_1656);
xor U1863 (N_1863,In_1903,In_10);
or U1864 (N_1864,In_957,In_647);
and U1865 (N_1865,In_530,In_1726);
or U1866 (N_1866,In_704,In_125);
or U1867 (N_1867,In_1785,In_228);
or U1868 (N_1868,In_424,In_1211);
nor U1869 (N_1869,In_1194,In_459);
nor U1870 (N_1870,In_342,In_803);
and U1871 (N_1871,In_1004,In_1235);
or U1872 (N_1872,In_133,In_1924);
and U1873 (N_1873,In_134,In_389);
nand U1874 (N_1874,In_1454,In_701);
nor U1875 (N_1875,In_280,In_22);
and U1876 (N_1876,In_779,In_679);
nand U1877 (N_1877,In_71,In_1439);
nand U1878 (N_1878,In_873,In_988);
and U1879 (N_1879,In_790,In_123);
nand U1880 (N_1880,In_930,In_643);
or U1881 (N_1881,In_504,In_123);
and U1882 (N_1882,In_1817,In_1591);
or U1883 (N_1883,In_1845,In_1744);
nor U1884 (N_1884,In_817,In_644);
nand U1885 (N_1885,In_1652,In_939);
or U1886 (N_1886,In_549,In_966);
xnor U1887 (N_1887,In_480,In_672);
and U1888 (N_1888,In_1874,In_326);
and U1889 (N_1889,In_1984,In_1819);
or U1890 (N_1890,In_1712,In_166);
nand U1891 (N_1891,In_6,In_1633);
nand U1892 (N_1892,In_888,In_1853);
and U1893 (N_1893,In_618,In_1369);
nand U1894 (N_1894,In_1762,In_391);
nand U1895 (N_1895,In_1641,In_151);
and U1896 (N_1896,In_1414,In_1000);
and U1897 (N_1897,In_726,In_1855);
or U1898 (N_1898,In_156,In_1644);
or U1899 (N_1899,In_614,In_1328);
and U1900 (N_1900,In_994,In_436);
nand U1901 (N_1901,In_591,In_812);
or U1902 (N_1902,In_2,In_1890);
nand U1903 (N_1903,In_1105,In_1750);
and U1904 (N_1904,In_1580,In_1691);
or U1905 (N_1905,In_1395,In_1614);
or U1906 (N_1906,In_229,In_1435);
or U1907 (N_1907,In_664,In_1341);
or U1908 (N_1908,In_1405,In_1776);
and U1909 (N_1909,In_1285,In_517);
nand U1910 (N_1910,In_314,In_850);
nor U1911 (N_1911,In_608,In_129);
and U1912 (N_1912,In_651,In_1729);
nor U1913 (N_1913,In_1878,In_1201);
xor U1914 (N_1914,In_1823,In_149);
and U1915 (N_1915,In_1650,In_1644);
nor U1916 (N_1916,In_1804,In_822);
nor U1917 (N_1917,In_225,In_113);
nand U1918 (N_1918,In_107,In_760);
or U1919 (N_1919,In_1827,In_225);
or U1920 (N_1920,In_398,In_1222);
nor U1921 (N_1921,In_1394,In_1658);
and U1922 (N_1922,In_1402,In_1942);
and U1923 (N_1923,In_724,In_833);
or U1924 (N_1924,In_286,In_1541);
or U1925 (N_1925,In_262,In_430);
nand U1926 (N_1926,In_733,In_1451);
and U1927 (N_1927,In_1731,In_100);
nor U1928 (N_1928,In_1212,In_133);
nand U1929 (N_1929,In_1952,In_667);
and U1930 (N_1930,In_1935,In_1678);
and U1931 (N_1931,In_701,In_525);
nand U1932 (N_1932,In_1203,In_1868);
xnor U1933 (N_1933,In_1029,In_1454);
nand U1934 (N_1934,In_218,In_1536);
nand U1935 (N_1935,In_1993,In_1853);
nand U1936 (N_1936,In_1245,In_1898);
or U1937 (N_1937,In_579,In_351);
and U1938 (N_1938,In_1924,In_1133);
nor U1939 (N_1939,In_133,In_925);
nand U1940 (N_1940,In_1343,In_230);
or U1941 (N_1941,In_1528,In_996);
or U1942 (N_1942,In_9,In_960);
or U1943 (N_1943,In_17,In_1963);
nor U1944 (N_1944,In_658,In_127);
or U1945 (N_1945,In_1027,In_541);
nand U1946 (N_1946,In_1110,In_1240);
xnor U1947 (N_1947,In_1408,In_1310);
nor U1948 (N_1948,In_912,In_1650);
or U1949 (N_1949,In_1255,In_1617);
nor U1950 (N_1950,In_1140,In_1763);
or U1951 (N_1951,In_1971,In_491);
xor U1952 (N_1952,In_1719,In_1384);
or U1953 (N_1953,In_972,In_514);
and U1954 (N_1954,In_371,In_1579);
nand U1955 (N_1955,In_1308,In_355);
or U1956 (N_1956,In_808,In_1167);
or U1957 (N_1957,In_908,In_1812);
nand U1958 (N_1958,In_180,In_497);
nor U1959 (N_1959,In_936,In_1620);
and U1960 (N_1960,In_1055,In_1573);
nand U1961 (N_1961,In_1360,In_1236);
or U1962 (N_1962,In_474,In_1571);
and U1963 (N_1963,In_1807,In_872);
and U1964 (N_1964,In_567,In_1200);
and U1965 (N_1965,In_203,In_977);
nor U1966 (N_1966,In_336,In_33);
nand U1967 (N_1967,In_1244,In_1904);
nand U1968 (N_1968,In_1012,In_1049);
and U1969 (N_1969,In_1254,In_1956);
nor U1970 (N_1970,In_602,In_1673);
xnor U1971 (N_1971,In_1480,In_328);
nor U1972 (N_1972,In_1971,In_1551);
or U1973 (N_1973,In_1484,In_1476);
nor U1974 (N_1974,In_51,In_1610);
or U1975 (N_1975,In_1514,In_670);
and U1976 (N_1976,In_1909,In_781);
nor U1977 (N_1977,In_1744,In_950);
or U1978 (N_1978,In_0,In_696);
or U1979 (N_1979,In_544,In_661);
or U1980 (N_1980,In_801,In_1397);
nor U1981 (N_1981,In_863,In_635);
or U1982 (N_1982,In_211,In_423);
or U1983 (N_1983,In_196,In_403);
nand U1984 (N_1984,In_232,In_1868);
and U1985 (N_1985,In_1816,In_490);
nor U1986 (N_1986,In_462,In_924);
nor U1987 (N_1987,In_521,In_1465);
or U1988 (N_1988,In_756,In_1959);
or U1989 (N_1989,In_1145,In_331);
and U1990 (N_1990,In_1921,In_140);
nor U1991 (N_1991,In_1948,In_1673);
xnor U1992 (N_1992,In_1956,In_1219);
nor U1993 (N_1993,In_1998,In_955);
xnor U1994 (N_1994,In_558,In_1261);
nor U1995 (N_1995,In_1397,In_1538);
and U1996 (N_1996,In_1772,In_280);
or U1997 (N_1997,In_856,In_344);
nor U1998 (N_1998,In_776,In_1523);
nand U1999 (N_1999,In_1041,In_1222);
nor U2000 (N_2000,N_1343,N_977);
and U2001 (N_2001,N_103,N_280);
nor U2002 (N_2002,N_1985,N_712);
nor U2003 (N_2003,N_1934,N_210);
and U2004 (N_2004,N_1122,N_1052);
or U2005 (N_2005,N_1534,N_849);
xor U2006 (N_2006,N_909,N_1062);
or U2007 (N_2007,N_1184,N_1508);
nand U2008 (N_2008,N_193,N_1223);
or U2009 (N_2009,N_1522,N_1279);
nor U2010 (N_2010,N_1780,N_425);
nand U2011 (N_2011,N_510,N_1300);
and U2012 (N_2012,N_1472,N_1526);
or U2013 (N_2013,N_982,N_1877);
or U2014 (N_2014,N_950,N_685);
or U2015 (N_2015,N_873,N_1267);
nor U2016 (N_2016,N_1627,N_1630);
nand U2017 (N_2017,N_88,N_1161);
and U2018 (N_2018,N_611,N_1225);
and U2019 (N_2019,N_1140,N_1853);
nand U2020 (N_2020,N_642,N_600);
nand U2021 (N_2021,N_388,N_449);
nand U2022 (N_2022,N_780,N_31);
nand U2023 (N_2023,N_184,N_864);
or U2024 (N_2024,N_1255,N_79);
and U2025 (N_2025,N_1682,N_1128);
xor U2026 (N_2026,N_1552,N_1382);
or U2027 (N_2027,N_317,N_1289);
or U2028 (N_2028,N_586,N_1330);
nor U2029 (N_2029,N_1355,N_1070);
or U2030 (N_2030,N_1925,N_1669);
or U2031 (N_2031,N_254,N_1432);
xnor U2032 (N_2032,N_466,N_1708);
xor U2033 (N_2033,N_12,N_1843);
xor U2034 (N_2034,N_108,N_485);
nand U2035 (N_2035,N_89,N_8);
nor U2036 (N_2036,N_1318,N_1668);
or U2037 (N_2037,N_1322,N_1480);
nor U2038 (N_2038,N_1380,N_918);
nand U2039 (N_2039,N_375,N_1915);
nand U2040 (N_2040,N_1453,N_1109);
or U2041 (N_2041,N_1118,N_1248);
and U2042 (N_2042,N_1023,N_771);
nor U2043 (N_2043,N_319,N_1944);
nand U2044 (N_2044,N_1547,N_7);
nand U2045 (N_2045,N_1990,N_387);
or U2046 (N_2046,N_1196,N_251);
and U2047 (N_2047,N_721,N_838);
or U2048 (N_2048,N_1660,N_1638);
or U2049 (N_2049,N_875,N_1164);
or U2050 (N_2050,N_1670,N_1914);
nor U2051 (N_2051,N_1895,N_1737);
xnor U2052 (N_2052,N_947,N_1600);
nand U2053 (N_2053,N_117,N_111);
xnor U2054 (N_2054,N_1976,N_659);
nor U2055 (N_2055,N_63,N_1878);
xor U2056 (N_2056,N_716,N_850);
or U2057 (N_2057,N_1507,N_1405);
nor U2058 (N_2058,N_306,N_393);
nand U2059 (N_2059,N_772,N_618);
or U2060 (N_2060,N_1617,N_818);
and U2061 (N_2061,N_1845,N_1779);
nand U2062 (N_2062,N_952,N_755);
or U2063 (N_2063,N_1932,N_1422);
or U2064 (N_2064,N_135,N_1957);
and U2065 (N_2065,N_311,N_788);
and U2066 (N_2066,N_1723,N_1285);
or U2067 (N_2067,N_1221,N_1215);
and U2068 (N_2068,N_284,N_1363);
nor U2069 (N_2069,N_1703,N_105);
nor U2070 (N_2070,N_444,N_1387);
nand U2071 (N_2071,N_1603,N_261);
nor U2072 (N_2072,N_462,N_1830);
and U2073 (N_2073,N_645,N_1975);
nor U2074 (N_2074,N_1991,N_252);
nand U2075 (N_2075,N_1209,N_890);
and U2076 (N_2076,N_792,N_1414);
nand U2077 (N_2077,N_382,N_914);
xor U2078 (N_2078,N_763,N_781);
or U2079 (N_2079,N_963,N_499);
or U2080 (N_2080,N_623,N_1523);
and U2081 (N_2081,N_1212,N_200);
nand U2082 (N_2082,N_406,N_112);
nand U2083 (N_2083,N_1046,N_514);
xor U2084 (N_2084,N_226,N_1130);
nand U2085 (N_2085,N_643,N_1888);
nor U2086 (N_2086,N_1439,N_824);
nand U2087 (N_2087,N_351,N_1698);
or U2088 (N_2088,N_23,N_422);
nand U2089 (N_2089,N_334,N_1981);
nand U2090 (N_2090,N_324,N_750);
or U2091 (N_2091,N_903,N_895);
nor U2092 (N_2092,N_1871,N_1494);
nor U2093 (N_2093,N_1873,N_744);
or U2094 (N_2094,N_1378,N_1012);
nor U2095 (N_2095,N_1763,N_1655);
and U2096 (N_2096,N_1483,N_1689);
or U2097 (N_2097,N_424,N_497);
or U2098 (N_2098,N_708,N_1226);
nor U2099 (N_2099,N_907,N_1538);
nand U2100 (N_2100,N_486,N_1063);
nand U2101 (N_2101,N_1415,N_1531);
nand U2102 (N_2102,N_411,N_1098);
and U2103 (N_2103,N_1272,N_1589);
or U2104 (N_2104,N_741,N_1276);
nand U2105 (N_2105,N_367,N_1358);
or U2106 (N_2106,N_1806,N_925);
or U2107 (N_2107,N_1851,N_1762);
nand U2108 (N_2108,N_1585,N_1704);
nor U2109 (N_2109,N_1574,N_511);
nor U2110 (N_2110,N_37,N_1119);
nor U2111 (N_2111,N_1263,N_143);
nor U2112 (N_2112,N_1919,N_292);
nor U2113 (N_2113,N_1352,N_1312);
xnor U2114 (N_2114,N_274,N_121);
and U2115 (N_2115,N_1163,N_1902);
nand U2116 (N_2116,N_1528,N_1211);
or U2117 (N_2117,N_1738,N_1974);
and U2118 (N_2118,N_126,N_598);
and U2119 (N_2119,N_1373,N_919);
or U2120 (N_2120,N_546,N_186);
nand U2121 (N_2121,N_144,N_561);
and U2122 (N_2122,N_910,N_1139);
nand U2123 (N_2123,N_1836,N_1733);
or U2124 (N_2124,N_1470,N_1258);
or U2125 (N_2125,N_854,N_619);
or U2126 (N_2126,N_348,N_141);
xnor U2127 (N_2127,N_1755,N_1306);
nand U2128 (N_2128,N_1663,N_752);
nand U2129 (N_2129,N_1581,N_521);
or U2130 (N_2130,N_1464,N_764);
and U2131 (N_2131,N_1634,N_188);
xor U2132 (N_2132,N_515,N_427);
and U2133 (N_2133,N_1813,N_1728);
or U2134 (N_2134,N_1781,N_1736);
nor U2135 (N_2135,N_962,N_1434);
nand U2136 (N_2136,N_1511,N_701);
nand U2137 (N_2137,N_1087,N_529);
or U2138 (N_2138,N_1691,N_1942);
and U2139 (N_2139,N_451,N_358);
nand U2140 (N_2140,N_1371,N_522);
or U2141 (N_2141,N_1980,N_735);
nor U2142 (N_2142,N_1407,N_509);
nand U2143 (N_2143,N_1699,N_520);
or U2144 (N_2144,N_756,N_1560);
and U2145 (N_2145,N_1461,N_92);
or U2146 (N_2146,N_1410,N_765);
or U2147 (N_2147,N_1165,N_1103);
or U2148 (N_2148,N_981,N_1541);
and U2149 (N_2149,N_187,N_174);
nor U2150 (N_2150,N_336,N_1427);
and U2151 (N_2151,N_1249,N_636);
or U2152 (N_2152,N_953,N_1961);
or U2153 (N_2153,N_917,N_1860);
nand U2154 (N_2154,N_615,N_550);
and U2155 (N_2155,N_1107,N_318);
or U2156 (N_2156,N_1295,N_214);
nor U2157 (N_2157,N_1462,N_965);
nor U2158 (N_2158,N_1654,N_68);
xnor U2159 (N_2159,N_1984,N_1852);
and U2160 (N_2160,N_423,N_1084);
nand U2161 (N_2161,N_582,N_342);
nor U2162 (N_2162,N_937,N_1190);
nand U2163 (N_2163,N_1594,N_1108);
and U2164 (N_2164,N_32,N_552);
and U2165 (N_2165,N_524,N_898);
nand U2166 (N_2166,N_244,N_1767);
nand U2167 (N_2167,N_1963,N_834);
nand U2168 (N_2168,N_1346,N_531);
nor U2169 (N_2169,N_39,N_1183);
nor U2170 (N_2170,N_535,N_1316);
nand U2171 (N_2171,N_227,N_124);
nand U2172 (N_2172,N_846,N_458);
nand U2173 (N_2173,N_1156,N_1452);
or U2174 (N_2174,N_1442,N_1816);
and U2175 (N_2175,N_626,N_1093);
and U2176 (N_2176,N_1003,N_748);
xnor U2177 (N_2177,N_1179,N_1734);
or U2178 (N_2178,N_1236,N_1490);
nand U2179 (N_2179,N_961,N_624);
or U2180 (N_2180,N_1768,N_1141);
nand U2181 (N_2181,N_305,N_443);
and U2182 (N_2182,N_276,N_1809);
or U2183 (N_2183,N_1092,N_1444);
and U2184 (N_2184,N_973,N_1497);
nor U2185 (N_2185,N_352,N_1310);
and U2186 (N_2186,N_1034,N_1078);
and U2187 (N_2187,N_452,N_1158);
xor U2188 (N_2188,N_1269,N_1596);
and U2189 (N_2189,N_1181,N_882);
and U2190 (N_2190,N_198,N_1198);
or U2191 (N_2191,N_421,N_663);
and U2192 (N_2192,N_1495,N_248);
or U2193 (N_2193,N_1745,N_1533);
and U2194 (N_2194,N_1232,N_585);
and U2195 (N_2195,N_1074,N_776);
xnor U2196 (N_2196,N_253,N_923);
nand U2197 (N_2197,N_177,N_1868);
or U2198 (N_2198,N_385,N_1941);
or U2199 (N_2199,N_1930,N_494);
nor U2200 (N_2200,N_145,N_817);
or U2201 (N_2201,N_402,N_1235);
nor U2202 (N_2202,N_110,N_312);
or U2203 (N_2203,N_418,N_1799);
nor U2204 (N_2204,N_1121,N_361);
nor U2205 (N_2205,N_1896,N_1067);
and U2206 (N_2206,N_1842,N_852);
or U2207 (N_2207,N_971,N_1825);
and U2208 (N_2208,N_264,N_1123);
and U2209 (N_2209,N_197,N_1862);
and U2210 (N_2210,N_58,N_1501);
nand U2211 (N_2211,N_1820,N_323);
and U2212 (N_2212,N_243,N_1839);
xor U2213 (N_2213,N_1337,N_1571);
or U2214 (N_2214,N_749,N_308);
and U2215 (N_2215,N_1396,N_1688);
and U2216 (N_2216,N_1135,N_80);
nand U2217 (N_2217,N_593,N_1374);
nand U2218 (N_2218,N_676,N_332);
nand U2219 (N_2219,N_1629,N_1955);
and U2220 (N_2220,N_1653,N_1129);
and U2221 (N_2221,N_83,N_167);
and U2222 (N_2222,N_534,N_1372);
nor U2223 (N_2223,N_1020,N_557);
nand U2224 (N_2224,N_941,N_616);
xor U2225 (N_2225,N_1567,N_934);
and U2226 (N_2226,N_596,N_1426);
nand U2227 (N_2227,N_1649,N_831);
nand U2228 (N_2228,N_1364,N_1091);
and U2229 (N_2229,N_1344,N_1000);
and U2230 (N_2230,N_1752,N_123);
nand U2231 (N_2231,N_128,N_1982);
xor U2232 (N_2232,N_660,N_1283);
xor U2233 (N_2233,N_1641,N_258);
nand U2234 (N_2234,N_500,N_389);
nand U2235 (N_2235,N_1770,N_1720);
nand U2236 (N_2236,N_1706,N_1419);
nand U2237 (N_2237,N_766,N_938);
xnor U2238 (N_2238,N_1025,N_1076);
and U2239 (N_2239,N_1385,N_1402);
nand U2240 (N_2240,N_313,N_1005);
or U2241 (N_2241,N_265,N_944);
nand U2242 (N_2242,N_1582,N_1929);
xnor U2243 (N_2243,N_1808,N_498);
and U2244 (N_2244,N_987,N_1124);
and U2245 (N_2245,N_1448,N_431);
xnor U2246 (N_2246,N_872,N_1615);
or U2247 (N_2247,N_1307,N_150);
nand U2248 (N_2248,N_863,N_349);
or U2249 (N_2249,N_827,N_1166);
or U2250 (N_2250,N_885,N_842);
or U2251 (N_2251,N_225,N_1220);
nand U2252 (N_2252,N_999,N_1502);
nand U2253 (N_2253,N_1521,N_779);
nor U2254 (N_2254,N_1889,N_1599);
and U2255 (N_2255,N_853,N_806);
and U2256 (N_2256,N_1401,N_906);
nor U2257 (N_2257,N_1875,N_574);
nand U2258 (N_2258,N_1867,N_1317);
or U2259 (N_2259,N_1788,N_986);
xnor U2260 (N_2260,N_413,N_76);
xor U2261 (N_2261,N_249,N_1758);
or U2262 (N_2262,N_1805,N_374);
and U2263 (N_2263,N_1536,N_18);
xor U2264 (N_2264,N_1692,N_1579);
and U2265 (N_2265,N_289,N_670);
or U2266 (N_2266,N_858,N_1381);
nor U2267 (N_2267,N_711,N_1077);
and U2268 (N_2268,N_1887,N_1553);
nand U2269 (N_2269,N_713,N_1550);
or U2270 (N_2270,N_213,N_905);
or U2271 (N_2271,N_1493,N_683);
or U2272 (N_2272,N_14,N_745);
nor U2273 (N_2273,N_206,N_1142);
nor U2274 (N_2274,N_353,N_271);
nand U2275 (N_2275,N_231,N_591);
nor U2276 (N_2276,N_983,N_1783);
nor U2277 (N_2277,N_1790,N_841);
xor U2278 (N_2278,N_1213,N_669);
and U2279 (N_2279,N_1619,N_82);
nand U2280 (N_2280,N_476,N_1241);
nand U2281 (N_2281,N_237,N_53);
xor U2282 (N_2282,N_1506,N_437);
or U2283 (N_2283,N_1133,N_828);
or U2284 (N_2284,N_69,N_114);
xnor U2285 (N_2285,N_1262,N_1614);
or U2286 (N_2286,N_1999,N_653);
and U2287 (N_2287,N_355,N_115);
nor U2288 (N_2288,N_1886,N_26);
and U2289 (N_2289,N_1265,N_803);
nor U2290 (N_2290,N_1510,N_1154);
or U2291 (N_2291,N_296,N_246);
nor U2292 (N_2292,N_816,N_1345);
nor U2293 (N_2293,N_714,N_1195);
or U2294 (N_2294,N_1840,N_65);
or U2295 (N_2295,N_1082,N_975);
nor U2296 (N_2296,N_1080,N_1075);
nand U2297 (N_2297,N_1822,N_1527);
or U2298 (N_2298,N_928,N_884);
nand U2299 (N_2299,N_1002,N_571);
xnor U2300 (N_2300,N_608,N_450);
nor U2301 (N_2301,N_1741,N_1509);
nor U2302 (N_2302,N_1719,N_467);
nand U2303 (N_2303,N_625,N_688);
and U2304 (N_2304,N_1988,N_1701);
nor U2305 (N_2305,N_844,N_1050);
nor U2306 (N_2306,N_1465,N_516);
nor U2307 (N_2307,N_1045,N_201);
nor U2308 (N_2308,N_1443,N_1053);
or U2309 (N_2309,N_517,N_166);
and U2310 (N_2310,N_1037,N_1714);
and U2311 (N_2311,N_1650,N_392);
and U2312 (N_2312,N_1469,N_1543);
nor U2313 (N_2313,N_560,N_929);
nand U2314 (N_2314,N_1548,N_930);
nand U2315 (N_2315,N_547,N_960);
and U2316 (N_2316,N_1308,N_597);
and U2317 (N_2317,N_1,N_5);
nor U2318 (N_2318,N_675,N_897);
or U2319 (N_2319,N_924,N_1782);
nor U2320 (N_2320,N_835,N_1881);
nor U2321 (N_2321,N_1416,N_1049);
or U2322 (N_2322,N_1819,N_1759);
xor U2323 (N_2323,N_232,N_1943);
or U2324 (N_2324,N_799,N_1847);
or U2325 (N_2325,N_922,N_456);
nor U2326 (N_2326,N_178,N_1369);
or U2327 (N_2327,N_1150,N_380);
and U2328 (N_2328,N_562,N_1970);
and U2329 (N_2329,N_568,N_980);
and U2330 (N_2330,N_1335,N_1673);
nand U2331 (N_2331,N_1244,N_646);
or U2332 (N_2332,N_1892,N_1962);
nand U2333 (N_2333,N_551,N_1127);
nor U2334 (N_2334,N_1171,N_221);
or U2335 (N_2335,N_813,N_822);
nand U2336 (N_2336,N_541,N_782);
nor U2337 (N_2337,N_696,N_1144);
or U2338 (N_2338,N_1390,N_1643);
and U2339 (N_2339,N_478,N_1972);
nor U2340 (N_2340,N_757,N_840);
xor U2341 (N_2341,N_403,N_286);
and U2342 (N_2342,N_902,N_268);
and U2343 (N_2343,N_321,N_1716);
nor U2344 (N_2344,N_281,N_1858);
nor U2345 (N_2345,N_1284,N_940);
nor U2346 (N_2346,N_698,N_359);
and U2347 (N_2347,N_1239,N_339);
or U2348 (N_2348,N_350,N_1712);
and U2349 (N_2349,N_156,N_1340);
nor U2350 (N_2350,N_576,N_1570);
or U2351 (N_2351,N_1217,N_484);
or U2352 (N_2352,N_1173,N_273);
xnor U2353 (N_2353,N_1910,N_943);
and U2354 (N_2354,N_77,N_310);
nand U2355 (N_2355,N_979,N_993);
nand U2356 (N_2356,N_1447,N_790);
or U2357 (N_2357,N_1288,N_1286);
and U2358 (N_2358,N_687,N_722);
and U2359 (N_2359,N_257,N_1750);
xor U2360 (N_2360,N_893,N_1879);
or U2361 (N_2361,N_1515,N_732);
and U2362 (N_2362,N_1298,N_996);
nand U2363 (N_2363,N_93,N_1730);
and U2364 (N_2364,N_131,N_584);
or U2365 (N_2365,N_935,N_33);
nand U2366 (N_2366,N_595,N_1246);
or U2367 (N_2367,N_1609,N_1998);
nor U2368 (N_2368,N_1398,N_1281);
nor U2369 (N_2369,N_1132,N_459);
nor U2370 (N_2370,N_1167,N_1519);
or U2371 (N_2371,N_445,N_915);
nand U2372 (N_2372,N_1940,N_1496);
nor U2373 (N_2373,N_1702,N_1019);
and U2374 (N_2374,N_1097,N_995);
nand U2375 (N_2375,N_1197,N_668);
nand U2376 (N_2376,N_1696,N_1802);
or U2377 (N_2377,N_1601,N_238);
nor U2378 (N_2378,N_1967,N_481);
and U2379 (N_2379,N_285,N_678);
and U2380 (N_2380,N_775,N_338);
or U2381 (N_2381,N_1551,N_344);
nor U2382 (N_2382,N_203,N_38);
nor U2383 (N_2383,N_211,N_1690);
or U2384 (N_2384,N_1893,N_212);
nor U2385 (N_2385,N_800,N_163);
nand U2386 (N_2386,N_224,N_345);
nand U2387 (N_2387,N_1834,N_1558);
nor U2388 (N_2388,N_1463,N_832);
and U2389 (N_2389,N_1408,N_573);
or U2390 (N_2390,N_1185,N_1458);
or U2391 (N_2391,N_240,N_648);
and U2392 (N_2392,N_287,N_1577);
xor U2393 (N_2393,N_40,N_1923);
or U2394 (N_2394,N_815,N_1032);
nor U2395 (N_2395,N_1951,N_43);
and U2396 (N_2396,N_1791,N_1437);
nand U2397 (N_2397,N_808,N_804);
xor U2398 (N_2398,N_1376,N_1718);
xor U2399 (N_2399,N_1593,N_635);
nand U2400 (N_2400,N_892,N_1817);
nand U2401 (N_2401,N_739,N_1922);
or U2402 (N_2402,N_632,N_833);
and U2403 (N_2403,N_1573,N_1769);
and U2404 (N_2404,N_1611,N_1977);
and U2405 (N_2405,N_1633,N_830);
and U2406 (N_2406,N_661,N_1661);
xor U2407 (N_2407,N_1801,N_230);
or U2408 (N_2408,N_705,N_1992);
or U2409 (N_2409,N_394,N_223);
nor U2410 (N_2410,N_519,N_731);
and U2411 (N_2411,N_233,N_297);
or U2412 (N_2412,N_1586,N_1821);
nand U2413 (N_2413,N_1987,N_183);
and U2414 (N_2414,N_1028,N_1064);
or U2415 (N_2415,N_1347,N_523);
or U2416 (N_2416,N_113,N_1754);
or U2417 (N_2417,N_506,N_1530);
or U2418 (N_2418,N_894,N_1200);
nand U2419 (N_2419,N_74,N_327);
nor U2420 (N_2420,N_1639,N_1178);
xor U2421 (N_2421,N_888,N_490);
or U2422 (N_2422,N_753,N_1027);
or U2423 (N_2423,N_404,N_137);
nand U2424 (N_2424,N_829,N_1489);
or U2425 (N_2425,N_60,N_335);
or U2426 (N_2426,N_1810,N_1208);
and U2427 (N_2427,N_369,N_988);
nor U2428 (N_2428,N_1377,N_347);
nor U2429 (N_2429,N_340,N_1245);
and U2430 (N_2430,N_761,N_530);
nor U2431 (N_2431,N_3,N_138);
xnor U2432 (N_2432,N_797,N_1112);
or U2433 (N_2433,N_1549,N_472);
xor U2434 (N_2434,N_569,N_447);
nand U2435 (N_2435,N_1412,N_290);
and U2436 (N_2436,N_677,N_1646);
xnor U2437 (N_2437,N_955,N_1604);
nor U2438 (N_2438,N_1058,N_1833);
or U2439 (N_2439,N_1039,N_1254);
or U2440 (N_2440,N_182,N_1438);
nor U2441 (N_2441,N_471,N_1116);
and U2442 (N_2442,N_1400,N_1499);
nand U2443 (N_2443,N_1349,N_837);
or U2444 (N_2444,N_1787,N_1882);
or U2445 (N_2445,N_1815,N_52);
nor U2446 (N_2446,N_398,N_159);
and U2447 (N_2447,N_770,N_158);
or U2448 (N_2448,N_630,N_1468);
nand U2449 (N_2449,N_1911,N_259);
nand U2450 (N_2450,N_1467,N_1939);
nor U2451 (N_2451,N_1906,N_189);
and U2452 (N_2452,N_633,N_1773);
nor U2453 (N_2453,N_1338,N_501);
and U2454 (N_2454,N_1683,N_185);
or U2455 (N_2455,N_370,N_878);
and U2456 (N_2456,N_508,N_868);
nand U2457 (N_2457,N_487,N_976);
and U2458 (N_2458,N_526,N_879);
and U2459 (N_2459,N_1360,N_1218);
and U2460 (N_2460,N_639,N_1435);
nand U2461 (N_2461,N_542,N_587);
nand U2462 (N_2462,N_1379,N_978);
nand U2463 (N_2463,N_638,N_1937);
nand U2464 (N_2464,N_1749,N_16);
nand U2465 (N_2465,N_738,N_1610);
nor U2466 (N_2466,N_1341,N_95);
nor U2467 (N_2467,N_371,N_656);
nor U2468 (N_2468,N_362,N_843);
nor U2469 (N_2469,N_991,N_1658);
or U2470 (N_2470,N_1433,N_1389);
xnor U2471 (N_2471,N_409,N_1162);
nor U2472 (N_2472,N_733,N_690);
xor U2473 (N_2473,N_658,N_19);
and U2474 (N_2474,N_1137,N_473);
or U2475 (N_2475,N_1562,N_845);
nor U2476 (N_2476,N_1993,N_657);
nand U2477 (N_2477,N_1675,N_62);
and U2478 (N_2478,N_565,N_1313);
nand U2479 (N_2479,N_1777,N_1384);
and U2480 (N_2480,N_614,N_1041);
nand U2481 (N_2481,N_759,N_699);
nand U2482 (N_2482,N_1789,N_1829);
or U2483 (N_2483,N_1818,N_1479);
or U2484 (N_2484,N_325,N_1841);
or U2485 (N_2485,N_162,N_1066);
xor U2486 (N_2486,N_1138,N_1863);
nand U2487 (N_2487,N_381,N_220);
nand U2488 (N_2488,N_164,N_1648);
or U2489 (N_2489,N_1030,N_951);
and U2490 (N_2490,N_865,N_1846);
or U2491 (N_2491,N_1812,N_1177);
or U2492 (N_2492,N_773,N_354);
or U2493 (N_2493,N_1492,N_1153);
nand U2494 (N_2494,N_94,N_1476);
and U2495 (N_2495,N_320,N_577);
nand U2496 (N_2496,N_768,N_417);
and U2497 (N_2497,N_1238,N_1071);
nand U2498 (N_2498,N_465,N_146);
or U2499 (N_2499,N_649,N_1252);
xor U2500 (N_2500,N_1440,N_1228);
and U2501 (N_2501,N_527,N_1631);
and U2502 (N_2502,N_691,N_1015);
nor U2503 (N_2503,N_365,N_1938);
nor U2504 (N_2504,N_533,N_1933);
xnor U2505 (N_2505,N_1169,N_537);
or U2506 (N_2506,N_73,N_15);
nand U2507 (N_2507,N_496,N_877);
xor U2508 (N_2508,N_118,N_1952);
nor U2509 (N_2509,N_309,N_674);
nor U2510 (N_2510,N_729,N_703);
or U2511 (N_2511,N_1884,N_400);
and U2512 (N_2512,N_1676,N_555);
and U2513 (N_2513,N_260,N_505);
or U2514 (N_2514,N_1303,N_1418);
or U2515 (N_2515,N_1029,N_1456);
nand U2516 (N_2516,N_1193,N_333);
and U2517 (N_2517,N_1848,N_1293);
and U2518 (N_2518,N_383,N_277);
nor U2519 (N_2519,N_559,N_168);
xor U2520 (N_2520,N_1216,N_1399);
xnor U2521 (N_2521,N_1155,N_789);
nor U2522 (N_2522,N_1986,N_30);
and U2523 (N_2523,N_647,N_122);
nand U2524 (N_2524,N_1595,N_363);
or U2525 (N_2525,N_1243,N_71);
nor U2526 (N_2526,N_432,N_997);
and U2527 (N_2527,N_1997,N_725);
and U2528 (N_2528,N_820,N_44);
or U2529 (N_2529,N_1561,N_777);
and U2530 (N_2530,N_970,N_440);
and U2531 (N_2531,N_1516,N_891);
and U2532 (N_2532,N_219,N_1455);
nand U2533 (N_2533,N_1684,N_1057);
nor U2534 (N_2534,N_1203,N_1575);
nand U2535 (N_2535,N_1257,N_572);
xor U2536 (N_2536,N_1931,N_1885);
and U2537 (N_2537,N_298,N_1563);
and U2538 (N_2538,N_454,N_106);
nand U2539 (N_2539,N_1251,N_1110);
nor U2540 (N_2540,N_720,N_315);
and U2541 (N_2541,N_1291,N_543);
nand U2542 (N_2542,N_1386,N_1705);
nor U2543 (N_2543,N_1824,N_1430);
or U2544 (N_2544,N_899,N_1036);
or U2545 (N_2545,N_1857,N_1271);
or U2546 (N_2546,N_629,N_479);
nand U2547 (N_2547,N_554,N_1814);
nor U2548 (N_2548,N_1336,N_1564);
nand U2549 (N_2549,N_1644,N_441);
nand U2550 (N_2550,N_876,N_1827);
nand U2551 (N_2551,N_1026,N_1207);
or U2552 (N_2552,N_1055,N_634);
nor U2553 (N_2553,N_1866,N_1230);
xor U2554 (N_2554,N_1735,N_1375);
and U2555 (N_2555,N_45,N_1010);
and U2556 (N_2556,N_662,N_116);
nor U2557 (N_2557,N_819,N_463);
nor U2558 (N_2558,N_1792,N_378);
nand U2559 (N_2559,N_96,N_959);
nand U2560 (N_2560,N_746,N_405);
xor U2561 (N_2561,N_1278,N_1651);
or U2562 (N_2562,N_889,N_1726);
nand U2563 (N_2563,N_946,N_1160);
and U2564 (N_2564,N_704,N_1978);
or U2565 (N_2565,N_1008,N_75);
xor U2566 (N_2566,N_426,N_1832);
and U2567 (N_2567,N_1449,N_316);
nand U2568 (N_2568,N_1157,N_504);
or U2569 (N_2569,N_870,N_1192);
nor U2570 (N_2570,N_730,N_307);
xor U2571 (N_2571,N_70,N_1765);
and U2572 (N_2572,N_109,N_628);
and U2573 (N_2573,N_811,N_1302);
nor U2574 (N_2574,N_439,N_825);
nand U2575 (N_2575,N_1233,N_1918);
xor U2576 (N_2576,N_1016,N_1088);
or U2577 (N_2577,N_1457,N_48);
xnor U2578 (N_2578,N_1305,N_857);
nand U2579 (N_2579,N_1069,N_1831);
nor U2580 (N_2580,N_682,N_563);
nand U2581 (N_2581,N_1557,N_132);
nor U2582 (N_2582,N_1994,N_1920);
and U2583 (N_2583,N_1473,N_627);
and U2584 (N_2584,N_98,N_1778);
nor U2585 (N_2585,N_171,N_1849);
or U2586 (N_2586,N_1441,N_1391);
xnor U2587 (N_2587,N_1693,N_1451);
or U2588 (N_2588,N_823,N_1428);
nor U2589 (N_2589,N_826,N_267);
nand U2590 (N_2590,N_583,N_196);
or U2591 (N_2591,N_489,N_740);
or U2592 (N_2592,N_356,N_1409);
nand U2593 (N_2593,N_1421,N_1598);
and U2594 (N_2594,N_886,N_1011);
or U2595 (N_2595,N_602,N_1870);
nand U2596 (N_2596,N_1174,N_1366);
xor U2597 (N_2597,N_1844,N_793);
or U2598 (N_2598,N_862,N_1040);
nor U2599 (N_2599,N_1007,N_1623);
nand U2600 (N_2600,N_241,N_100);
nand U2601 (N_2601,N_1756,N_1960);
or U2602 (N_2602,N_1309,N_322);
nor U2603 (N_2603,N_153,N_107);
xnor U2604 (N_2604,N_1280,N_99);
or U2605 (N_2605,N_1106,N_612);
nor U2606 (N_2606,N_1478,N_1393);
xor U2607 (N_2607,N_1068,N_1250);
xor U2608 (N_2608,N_1540,N_896);
and U2609 (N_2609,N_1270,N_1539);
xnor U2610 (N_2610,N_1392,N_190);
nor U2611 (N_2611,N_176,N_967);
or U2612 (N_2612,N_1319,N_1104);
or U2613 (N_2613,N_1081,N_742);
nand U2614 (N_2614,N_1898,N_1089);
nand U2615 (N_2615,N_255,N_707);
nor U2616 (N_2616,N_968,N_1147);
nand U2617 (N_2617,N_1370,N_1202);
or U2618 (N_2618,N_1065,N_715);
and U2619 (N_2619,N_566,N_1724);
nand U2620 (N_2620,N_589,N_130);
nor U2621 (N_2621,N_1176,N_809);
xor U2622 (N_2622,N_1912,N_860);
nand U2623 (N_2623,N_1194,N_1743);
and U2624 (N_2624,N_758,N_949);
nor U2625 (N_2625,N_1707,N_1013);
or U2626 (N_2626,N_1182,N_1354);
nor U2627 (N_2627,N_651,N_1126);
and U2628 (N_2628,N_357,N_536);
and U2629 (N_2629,N_1722,N_855);
nand U2630 (N_2630,N_1620,N_1983);
and U2631 (N_2631,N_640,N_1090);
or U2632 (N_2632,N_1460,N_710);
nor U2633 (N_2633,N_942,N_379);
and U2634 (N_2634,N_1713,N_1628);
nor U2635 (N_2635,N_1175,N_1956);
nor U2636 (N_2636,N_1512,N_1913);
nand U2637 (N_2637,N_1766,N_1214);
and U2638 (N_2638,N_637,N_266);
nor U2639 (N_2639,N_360,N_429);
nand U2640 (N_2640,N_140,N_460);
xnor U2641 (N_2641,N_1314,N_548);
xnor U2642 (N_2642,N_412,N_1517);
nand U2643 (N_2643,N_29,N_35);
and U2644 (N_2644,N_1880,N_1260);
xor U2645 (N_2645,N_1612,N_1785);
or U2646 (N_2646,N_165,N_1024);
or U2647 (N_2647,N_477,N_1657);
xnor U2648 (N_2648,N_1056,N_364);
nor U2649 (N_2649,N_784,N_1261);
nand U2650 (N_2650,N_180,N_1608);
or U2651 (N_2651,N_807,N_1229);
xnor U2652 (N_2652,N_1796,N_1275);
and U2653 (N_2653,N_61,N_1954);
xnor U2654 (N_2654,N_1367,N_588);
nor U2655 (N_2655,N_1085,N_681);
nand U2656 (N_2656,N_346,N_1290);
nor U2657 (N_2657,N_1383,N_461);
xor U2658 (N_2658,N_139,N_1775);
or U2659 (N_2659,N_1237,N_1921);
nand U2660 (N_2660,N_1397,N_1436);
or U2661 (N_2661,N_1647,N_920);
and U2662 (N_2662,N_1488,N_1640);
nor U2663 (N_2663,N_64,N_672);
and U2664 (N_2664,N_1545,N_1328);
or U2665 (N_2665,N_1578,N_700);
or U2666 (N_2666,N_912,N_512);
nor U2667 (N_2667,N_1227,N_901);
nand U2668 (N_2668,N_686,N_28);
nand U2669 (N_2669,N_1945,N_9);
nand U2670 (N_2670,N_1872,N_607);
and U2671 (N_2671,N_1664,N_692);
xor U2672 (N_2672,N_1725,N_847);
or U2673 (N_2673,N_926,N_1964);
xnor U2674 (N_2674,N_610,N_578);
xor U2675 (N_2675,N_1231,N_1856);
or U2676 (N_2676,N_594,N_331);
xnor U2677 (N_2677,N_985,N_81);
nor U2678 (N_2678,N_1823,N_709);
nand U2679 (N_2679,N_377,N_839);
and U2680 (N_2680,N_1727,N_1869);
nor U2681 (N_2681,N_1331,N_1111);
xnor U2682 (N_2682,N_1188,N_256);
nor U2683 (N_2683,N_1021,N_718);
nand U2684 (N_2684,N_1224,N_434);
and U2685 (N_2685,N_1277,N_1905);
and U2686 (N_2686,N_1546,N_1001);
nor U2687 (N_2687,N_396,N_1753);
and U2688 (N_2688,N_989,N_613);
nand U2689 (N_2689,N_181,N_415);
or U2690 (N_2690,N_783,N_397);
nand U2691 (N_2691,N_1356,N_1061);
nor U2692 (N_2692,N_1148,N_272);
or U2693 (N_2693,N_1597,N_664);
nor U2694 (N_2694,N_482,N_127);
nand U2695 (N_2695,N_1950,N_1253);
and U2696 (N_2696,N_1742,N_419);
and U2697 (N_2697,N_1900,N_549);
or U2698 (N_2698,N_101,N_457);
or U2699 (N_2699,N_160,N_1423);
nand U2700 (N_2700,N_1047,N_1296);
nor U2701 (N_2701,N_693,N_133);
nand U2702 (N_2702,N_1031,N_939);
or U2703 (N_2703,N_1351,N_1446);
or U2704 (N_2704,N_97,N_1006);
and U2705 (N_2705,N_1861,N_1187);
xor U2706 (N_2706,N_1191,N_410);
nand U2707 (N_2707,N_1083,N_337);
or U2708 (N_2708,N_134,N_723);
or U2709 (N_2709,N_1907,N_282);
and U2710 (N_2710,N_1004,N_288);
or U2711 (N_2711,N_620,N_1583);
or U2712 (N_2712,N_974,N_395);
and U2713 (N_2713,N_697,N_1477);
xnor U2714 (N_2714,N_204,N_1899);
or U2715 (N_2715,N_326,N_1324);
nand U2716 (N_2716,N_278,N_1429);
or U2717 (N_2717,N_812,N_673);
or U2718 (N_2718,N_767,N_1927);
nor U2719 (N_2719,N_617,N_438);
and U2720 (N_2720,N_1099,N_11);
nor U2721 (N_2721,N_998,N_1606);
nor U2722 (N_2722,N_1079,N_57);
nor U2723 (N_2723,N_1301,N_694);
nor U2724 (N_2724,N_215,N_936);
nand U2725 (N_2725,N_373,N_900);
nand U2726 (N_2726,N_1095,N_1917);
nor U2727 (N_2727,N_1795,N_1266);
nor U2728 (N_2728,N_1311,N_908);
and U2729 (N_2729,N_368,N_291);
and U2730 (N_2730,N_760,N_518);
xor U2731 (N_2731,N_726,N_1120);
nor U2732 (N_2732,N_1935,N_1968);
xor U2733 (N_2733,N_1592,N_667);
xnor U2734 (N_2734,N_1803,N_1761);
or U2735 (N_2735,N_719,N_469);
or U2736 (N_2736,N_590,N_25);
xor U2737 (N_2737,N_1326,N_1100);
and U2738 (N_2738,N_1555,N_1491);
or U2739 (N_2739,N_1949,N_1159);
and U2740 (N_2740,N_234,N_46);
xor U2741 (N_2741,N_1798,N_407);
and U2742 (N_2742,N_1897,N_91);
or U2743 (N_2743,N_1924,N_270);
nor U2744 (N_2744,N_1580,N_1883);
nand U2745 (N_2745,N_604,N_1678);
nor U2746 (N_2746,N_666,N_1222);
nand U2747 (N_2747,N_59,N_87);
nor U2748 (N_2748,N_199,N_1757);
nor U2749 (N_2749,N_575,N_1746);
nor U2750 (N_2750,N_1125,N_1838);
nor U2751 (N_2751,N_866,N_1835);
nor U2752 (N_2752,N_250,N_1514);
nand U2753 (N_2753,N_1315,N_1971);
nand U2754 (N_2754,N_957,N_921);
and U2755 (N_2755,N_480,N_433);
nor U2756 (N_2756,N_263,N_283);
nor U2757 (N_2757,N_1264,N_1891);
xnor U2758 (N_2758,N_245,N_1569);
nand U2759 (N_2759,N_229,N_247);
nor U2760 (N_2760,N_17,N_1048);
or U2761 (N_2761,N_1748,N_474);
xnor U2762 (N_2762,N_1947,N_1804);
nand U2763 (N_2763,N_1017,N_796);
nand U2764 (N_2764,N_172,N_1717);
nor U2765 (N_2765,N_1424,N_1665);
nand U2766 (N_2766,N_558,N_1959);
nor U2767 (N_2767,N_601,N_650);
nor U2768 (N_2768,N_1096,N_671);
nor U2769 (N_2769,N_1544,N_366);
nor U2770 (N_2770,N_507,N_102);
and U2771 (N_2771,N_1953,N_737);
and U2772 (N_2772,N_1584,N_136);
xor U2773 (N_2773,N_1687,N_1680);
nand U2774 (N_2774,N_856,N_1180);
or U2775 (N_2775,N_390,N_1686);
nand U2776 (N_2776,N_1454,N_1556);
nand U2777 (N_2777,N_119,N_4);
or U2778 (N_2778,N_1850,N_599);
and U2779 (N_2779,N_1321,N_1625);
and U2780 (N_2780,N_1450,N_1710);
nand U2781 (N_2781,N_1325,N_1559);
nor U2782 (N_2782,N_525,N_493);
nand U2783 (N_2783,N_1094,N_275);
and U2784 (N_2784,N_1903,N_149);
nand U2785 (N_2785,N_1890,N_727);
nand U2786 (N_2786,N_1323,N_1537);
nor U2787 (N_2787,N_1826,N_1909);
nor U2788 (N_2788,N_1711,N_1388);
nor U2789 (N_2789,N_54,N_931);
nor U2790 (N_2790,N_927,N_805);
or U2791 (N_2791,N_859,N_239);
nor U2792 (N_2792,N_1685,N_216);
and U2793 (N_2793,N_1874,N_1073);
and U2794 (N_2794,N_964,N_836);
and U2795 (N_2795,N_222,N_1168);
nand U2796 (N_2796,N_142,N_581);
nor U2797 (N_2797,N_314,N_1022);
nor U2798 (N_2798,N_1481,N_774);
and U2799 (N_2799,N_762,N_1334);
nand U2800 (N_2800,N_874,N_279);
or U2801 (N_2801,N_72,N_861);
nor U2802 (N_2802,N_1667,N_329);
nand U2803 (N_2803,N_399,N_1287);
nand U2804 (N_2804,N_1828,N_1042);
and U2805 (N_2805,N_1113,N_1149);
nor U2806 (N_2806,N_202,N_1044);
or U2807 (N_2807,N_706,N_1486);
nor U2808 (N_2808,N_242,N_448);
nand U2809 (N_2809,N_702,N_169);
nand U2810 (N_2810,N_990,N_236);
xnor U2811 (N_2811,N_1626,N_84);
or U2812 (N_2812,N_994,N_302);
and U2813 (N_2813,N_1320,N_468);
and U2814 (N_2814,N_1359,N_1350);
and U2815 (N_2815,N_20,N_1086);
nor U2816 (N_2816,N_1206,N_1672);
nand U2817 (N_2817,N_1855,N_304);
nor U2818 (N_2818,N_430,N_1590);
or U2819 (N_2819,N_1695,N_1425);
nand U2820 (N_2820,N_293,N_341);
or U2821 (N_2821,N_1652,N_1786);
xnor U2822 (N_2822,N_1764,N_455);
and U2823 (N_2823,N_564,N_553);
or U2824 (N_2824,N_1500,N_1294);
nor U2825 (N_2825,N_1186,N_1715);
and U2826 (N_2826,N_954,N_376);
and U2827 (N_2827,N_769,N_1666);
nor U2828 (N_2828,N_401,N_622);
nand U2829 (N_2829,N_1622,N_1189);
xor U2830 (N_2830,N_24,N_194);
nor U2831 (N_2831,N_1172,N_1431);
and U2832 (N_2832,N_217,N_1115);
nor U2833 (N_2833,N_717,N_1807);
or U2834 (N_2834,N_372,N_191);
xnor U2835 (N_2835,N_1700,N_1417);
nand U2836 (N_2836,N_956,N_147);
and U2837 (N_2837,N_1072,N_475);
nand U2838 (N_2838,N_1256,N_1529);
nand U2839 (N_2839,N_1674,N_1525);
nand U2840 (N_2840,N_945,N_1487);
nand U2841 (N_2841,N_751,N_1259);
nand U2842 (N_2842,N_1339,N_1136);
xor U2843 (N_2843,N_992,N_179);
or U2844 (N_2844,N_0,N_343);
and U2845 (N_2845,N_736,N_1060);
nand U2846 (N_2846,N_1681,N_1505);
or U2847 (N_2847,N_1043,N_262);
or U2848 (N_2848,N_170,N_503);
nor U2849 (N_2849,N_652,N_1504);
nor U2850 (N_2850,N_801,N_1989);
nand U2851 (N_2851,N_1542,N_814);
nor U2852 (N_2852,N_1904,N_1482);
nand U2853 (N_2853,N_680,N_34);
and U2854 (N_2854,N_1170,N_1772);
and U2855 (N_2855,N_1901,N_1613);
nand U2856 (N_2856,N_1794,N_747);
or U2857 (N_2857,N_1353,N_1102);
nand U2858 (N_2858,N_1709,N_786);
or U2859 (N_2859,N_78,N_1966);
xor U2860 (N_2860,N_1624,N_1797);
nand U2861 (N_2861,N_1679,N_50);
nor U2862 (N_2862,N_1740,N_540);
nand U2863 (N_2863,N_958,N_1268);
or U2864 (N_2864,N_1776,N_207);
nor U2865 (N_2865,N_125,N_1471);
nand U2866 (N_2866,N_90,N_299);
and U2867 (N_2867,N_1632,N_1744);
nor U2868 (N_2868,N_1739,N_603);
and U2869 (N_2869,N_1908,N_1327);
nand U2870 (N_2870,N_1299,N_1205);
nor U2871 (N_2871,N_1282,N_1771);
nor U2872 (N_2872,N_966,N_556);
nor U2873 (N_2873,N_1014,N_1524);
nand U2874 (N_2874,N_442,N_785);
nand U2875 (N_2875,N_1051,N_1059);
or U2876 (N_2876,N_1973,N_609);
or U2877 (N_2877,N_1729,N_416);
and U2878 (N_2878,N_1995,N_66);
or U2879 (N_2879,N_1605,N_1498);
and U2880 (N_2880,N_1420,N_86);
xnor U2881 (N_2881,N_1240,N_1273);
nand U2882 (N_2882,N_1747,N_802);
nand U2883 (N_2883,N_294,N_295);
and U2884 (N_2884,N_1009,N_1865);
xnor U2885 (N_2885,N_1131,N_1199);
and U2886 (N_2886,N_435,N_1928);
nor U2887 (N_2887,N_1576,N_1694);
nor U2888 (N_2888,N_1635,N_205);
nor U2889 (N_2889,N_933,N_1946);
nand U2890 (N_2890,N_1554,N_161);
nand U2891 (N_2891,N_1242,N_436);
or U2892 (N_2892,N_1361,N_1936);
nor U2893 (N_2893,N_192,N_384);
nand U2894 (N_2894,N_810,N_1357);
xor U2895 (N_2895,N_1588,N_173);
nand U2896 (N_2896,N_606,N_984);
nor U2897 (N_2897,N_218,N_209);
nor U2898 (N_2898,N_228,N_1800);
xnor U2899 (N_2899,N_1969,N_679);
xnor U2900 (N_2900,N_21,N_1342);
nor U2901 (N_2901,N_175,N_1774);
and U2902 (N_2902,N_1403,N_67);
or U2903 (N_2903,N_913,N_1332);
nor U2904 (N_2904,N_969,N_464);
nand U2905 (N_2905,N_129,N_754);
or U2906 (N_2906,N_328,N_1837);
and U2907 (N_2907,N_689,N_269);
or U2908 (N_2908,N_605,N_152);
and U2909 (N_2909,N_154,N_867);
and U2910 (N_2910,N_654,N_545);
nand U2911 (N_2911,N_1105,N_794);
xnor U2912 (N_2912,N_1114,N_470);
and U2913 (N_2913,N_155,N_1143);
nor U2914 (N_2914,N_492,N_1365);
nor U2915 (N_2915,N_55,N_27);
xor U2916 (N_2916,N_1394,N_1151);
nand U2917 (N_2917,N_1656,N_1297);
and U2918 (N_2918,N_22,N_1965);
or U2919 (N_2919,N_580,N_1134);
and U2920 (N_2920,N_1234,N_538);
and U2921 (N_2921,N_1572,N_1018);
and U2922 (N_2922,N_1304,N_1751);
or U2923 (N_2923,N_532,N_1731);
nand U2924 (N_2924,N_13,N_916);
nand U2925 (N_2925,N_1671,N_684);
or U2926 (N_2926,N_528,N_1518);
nor U2927 (N_2927,N_798,N_871);
or U2928 (N_2928,N_1926,N_1894);
and U2929 (N_2929,N_1996,N_56);
xnor U2930 (N_2930,N_1636,N_1645);
xor U2931 (N_2931,N_1348,N_972);
nor U2932 (N_2932,N_728,N_303);
nand U2933 (N_2933,N_120,N_41);
nand U2934 (N_2934,N_724,N_1038);
or U2935 (N_2935,N_948,N_1395);
or U2936 (N_2936,N_1732,N_1292);
and U2937 (N_2937,N_495,N_195);
nor U2938 (N_2938,N_644,N_1485);
and U2939 (N_2939,N_1760,N_787);
and U2940 (N_2940,N_1274,N_1568);
and U2941 (N_2941,N_848,N_386);
nor U2942 (N_2942,N_881,N_665);
and U2943 (N_2943,N_2,N_1117);
and U2944 (N_2944,N_1784,N_49);
nor U2945 (N_2945,N_1204,N_1854);
nand U2946 (N_2946,N_1474,N_1618);
or U2947 (N_2947,N_1219,N_1602);
xnor U2948 (N_2948,N_880,N_420);
xnor U2949 (N_2949,N_1368,N_1201);
or U2950 (N_2950,N_791,N_695);
nor U2951 (N_2951,N_1035,N_301);
and U2952 (N_2952,N_1662,N_10);
and U2953 (N_2953,N_1793,N_1145);
nor U2954 (N_2954,N_1565,N_1591);
and U2955 (N_2955,N_1948,N_1466);
nand U2956 (N_2956,N_734,N_208);
nor U2957 (N_2957,N_869,N_235);
nor U2958 (N_2958,N_592,N_1607);
or U2959 (N_2959,N_414,N_904);
and U2960 (N_2960,N_491,N_151);
xnor U2961 (N_2961,N_1721,N_887);
and U2962 (N_2962,N_1621,N_743);
nor U2963 (N_2963,N_157,N_579);
xor U2964 (N_2964,N_1864,N_300);
and U2965 (N_2965,N_1637,N_446);
nand U2966 (N_2966,N_883,N_483);
nand U2967 (N_2967,N_1979,N_641);
and U2968 (N_2968,N_391,N_36);
or U2969 (N_2969,N_1054,N_47);
and U2970 (N_2970,N_1404,N_795);
nor U2971 (N_2971,N_1503,N_1958);
or U2972 (N_2972,N_1210,N_1677);
and U2973 (N_2973,N_1535,N_539);
or U2974 (N_2974,N_655,N_621);
nor U2975 (N_2975,N_851,N_502);
and U2976 (N_2976,N_408,N_1406);
and U2977 (N_2977,N_1033,N_513);
and U2978 (N_2978,N_1362,N_453);
nor U2979 (N_2979,N_544,N_1616);
nor U2980 (N_2980,N_1859,N_1459);
nor U2981 (N_2981,N_932,N_330);
nand U2982 (N_2982,N_1513,N_148);
nand U2983 (N_2983,N_570,N_1101);
nand U2984 (N_2984,N_42,N_1876);
xor U2985 (N_2985,N_911,N_1247);
nand U2986 (N_2986,N_1475,N_1566);
and U2987 (N_2987,N_1445,N_1484);
xnor U2988 (N_2988,N_1659,N_567);
and U2989 (N_2989,N_488,N_85);
or U2990 (N_2990,N_1520,N_778);
or U2991 (N_2991,N_1413,N_1587);
nand U2992 (N_2992,N_1642,N_51);
nand U2993 (N_2993,N_1329,N_1697);
or U2994 (N_2994,N_1411,N_1532);
nand U2995 (N_2995,N_104,N_1916);
nand U2996 (N_2996,N_1333,N_6);
or U2997 (N_2997,N_428,N_821);
or U2998 (N_2998,N_1152,N_1811);
or U2999 (N_2999,N_1146,N_631);
nor U3000 (N_3000,N_310,N_1649);
or U3001 (N_3001,N_139,N_1210);
or U3002 (N_3002,N_1725,N_1514);
xor U3003 (N_3003,N_781,N_765);
nand U3004 (N_3004,N_320,N_1103);
and U3005 (N_3005,N_1939,N_294);
nor U3006 (N_3006,N_1681,N_207);
nor U3007 (N_3007,N_1734,N_1465);
nor U3008 (N_3008,N_1318,N_597);
or U3009 (N_3009,N_1721,N_1977);
or U3010 (N_3010,N_1266,N_1216);
or U3011 (N_3011,N_1888,N_1669);
nor U3012 (N_3012,N_1684,N_1501);
nand U3013 (N_3013,N_766,N_1722);
and U3014 (N_3014,N_1992,N_1243);
and U3015 (N_3015,N_1764,N_695);
xnor U3016 (N_3016,N_546,N_1272);
and U3017 (N_3017,N_1269,N_1334);
nor U3018 (N_3018,N_1231,N_405);
nand U3019 (N_3019,N_195,N_1330);
and U3020 (N_3020,N_145,N_223);
and U3021 (N_3021,N_1540,N_1978);
nand U3022 (N_3022,N_740,N_560);
nor U3023 (N_3023,N_689,N_641);
nand U3024 (N_3024,N_1787,N_1540);
nand U3025 (N_3025,N_274,N_239);
or U3026 (N_3026,N_1953,N_118);
xnor U3027 (N_3027,N_1794,N_1708);
nand U3028 (N_3028,N_637,N_1671);
and U3029 (N_3029,N_1822,N_1787);
and U3030 (N_3030,N_1402,N_1739);
or U3031 (N_3031,N_745,N_1614);
or U3032 (N_3032,N_912,N_803);
xor U3033 (N_3033,N_21,N_1257);
nor U3034 (N_3034,N_188,N_492);
nand U3035 (N_3035,N_1625,N_72);
nand U3036 (N_3036,N_579,N_144);
or U3037 (N_3037,N_540,N_598);
nor U3038 (N_3038,N_184,N_1766);
or U3039 (N_3039,N_1161,N_740);
or U3040 (N_3040,N_853,N_1120);
and U3041 (N_3041,N_1160,N_1656);
nor U3042 (N_3042,N_1575,N_276);
nor U3043 (N_3043,N_782,N_1645);
nor U3044 (N_3044,N_1168,N_850);
nor U3045 (N_3045,N_488,N_464);
or U3046 (N_3046,N_465,N_1781);
and U3047 (N_3047,N_1266,N_738);
xor U3048 (N_3048,N_505,N_418);
or U3049 (N_3049,N_249,N_923);
nand U3050 (N_3050,N_122,N_1484);
and U3051 (N_3051,N_1245,N_920);
xnor U3052 (N_3052,N_1022,N_931);
nand U3053 (N_3053,N_1658,N_1196);
or U3054 (N_3054,N_1904,N_693);
or U3055 (N_3055,N_954,N_1444);
or U3056 (N_3056,N_1121,N_1378);
or U3057 (N_3057,N_1559,N_1199);
or U3058 (N_3058,N_344,N_190);
nand U3059 (N_3059,N_851,N_263);
xor U3060 (N_3060,N_1699,N_1311);
or U3061 (N_3061,N_215,N_1158);
or U3062 (N_3062,N_1443,N_1585);
and U3063 (N_3063,N_694,N_1441);
or U3064 (N_3064,N_68,N_20);
and U3065 (N_3065,N_1292,N_1028);
and U3066 (N_3066,N_204,N_1680);
or U3067 (N_3067,N_731,N_328);
nor U3068 (N_3068,N_137,N_567);
nor U3069 (N_3069,N_703,N_254);
nand U3070 (N_3070,N_1994,N_1604);
or U3071 (N_3071,N_1929,N_654);
nor U3072 (N_3072,N_583,N_603);
and U3073 (N_3073,N_1003,N_408);
xnor U3074 (N_3074,N_355,N_1658);
and U3075 (N_3075,N_611,N_1384);
xnor U3076 (N_3076,N_1996,N_1141);
nand U3077 (N_3077,N_325,N_1538);
or U3078 (N_3078,N_492,N_940);
or U3079 (N_3079,N_1217,N_1237);
nand U3080 (N_3080,N_1728,N_1100);
nand U3081 (N_3081,N_1623,N_1750);
or U3082 (N_3082,N_503,N_1345);
nand U3083 (N_3083,N_1803,N_181);
nor U3084 (N_3084,N_55,N_301);
or U3085 (N_3085,N_1403,N_1467);
or U3086 (N_3086,N_887,N_1518);
or U3087 (N_3087,N_214,N_1443);
xnor U3088 (N_3088,N_409,N_1434);
nand U3089 (N_3089,N_727,N_1622);
and U3090 (N_3090,N_979,N_227);
or U3091 (N_3091,N_779,N_129);
or U3092 (N_3092,N_468,N_1970);
or U3093 (N_3093,N_982,N_1618);
nand U3094 (N_3094,N_1750,N_1044);
nand U3095 (N_3095,N_1910,N_432);
and U3096 (N_3096,N_581,N_660);
nor U3097 (N_3097,N_1470,N_459);
nor U3098 (N_3098,N_1755,N_540);
xnor U3099 (N_3099,N_1235,N_682);
and U3100 (N_3100,N_678,N_1978);
xnor U3101 (N_3101,N_1937,N_1749);
nor U3102 (N_3102,N_1388,N_852);
nand U3103 (N_3103,N_963,N_1181);
xor U3104 (N_3104,N_466,N_1531);
nand U3105 (N_3105,N_267,N_55);
and U3106 (N_3106,N_1077,N_1468);
nand U3107 (N_3107,N_1205,N_1115);
nand U3108 (N_3108,N_695,N_79);
and U3109 (N_3109,N_1654,N_226);
nor U3110 (N_3110,N_1788,N_1550);
and U3111 (N_3111,N_361,N_526);
or U3112 (N_3112,N_1472,N_1318);
or U3113 (N_3113,N_1371,N_1719);
nand U3114 (N_3114,N_347,N_514);
nor U3115 (N_3115,N_1199,N_914);
or U3116 (N_3116,N_1104,N_3);
xor U3117 (N_3117,N_1147,N_850);
nand U3118 (N_3118,N_215,N_1629);
and U3119 (N_3119,N_1776,N_1789);
nand U3120 (N_3120,N_1036,N_1931);
or U3121 (N_3121,N_390,N_102);
and U3122 (N_3122,N_1311,N_108);
or U3123 (N_3123,N_568,N_208);
nand U3124 (N_3124,N_1139,N_893);
and U3125 (N_3125,N_272,N_620);
or U3126 (N_3126,N_1651,N_17);
nor U3127 (N_3127,N_1244,N_975);
nor U3128 (N_3128,N_1772,N_1970);
nand U3129 (N_3129,N_1219,N_964);
and U3130 (N_3130,N_118,N_389);
and U3131 (N_3131,N_1977,N_941);
nand U3132 (N_3132,N_1266,N_742);
nor U3133 (N_3133,N_1097,N_1182);
nor U3134 (N_3134,N_304,N_790);
nor U3135 (N_3135,N_1960,N_534);
or U3136 (N_3136,N_997,N_155);
or U3137 (N_3137,N_1404,N_567);
and U3138 (N_3138,N_1635,N_226);
nor U3139 (N_3139,N_804,N_211);
and U3140 (N_3140,N_1938,N_333);
or U3141 (N_3141,N_776,N_1180);
nand U3142 (N_3142,N_1348,N_757);
or U3143 (N_3143,N_1889,N_574);
nand U3144 (N_3144,N_755,N_526);
or U3145 (N_3145,N_1729,N_1042);
or U3146 (N_3146,N_248,N_261);
or U3147 (N_3147,N_43,N_642);
nand U3148 (N_3148,N_1698,N_134);
nor U3149 (N_3149,N_1438,N_1876);
nand U3150 (N_3150,N_1073,N_1060);
nor U3151 (N_3151,N_270,N_1716);
nor U3152 (N_3152,N_1683,N_673);
nor U3153 (N_3153,N_96,N_1399);
or U3154 (N_3154,N_860,N_230);
nor U3155 (N_3155,N_981,N_176);
xor U3156 (N_3156,N_775,N_1356);
or U3157 (N_3157,N_271,N_724);
and U3158 (N_3158,N_1747,N_1340);
nor U3159 (N_3159,N_1882,N_1460);
and U3160 (N_3160,N_525,N_1363);
nor U3161 (N_3161,N_860,N_1117);
xnor U3162 (N_3162,N_565,N_1738);
and U3163 (N_3163,N_1271,N_1097);
nor U3164 (N_3164,N_1920,N_855);
nor U3165 (N_3165,N_312,N_174);
or U3166 (N_3166,N_872,N_1610);
nand U3167 (N_3167,N_521,N_1750);
nand U3168 (N_3168,N_556,N_1754);
and U3169 (N_3169,N_1525,N_1877);
xor U3170 (N_3170,N_608,N_534);
xnor U3171 (N_3171,N_1437,N_212);
or U3172 (N_3172,N_624,N_778);
xor U3173 (N_3173,N_34,N_686);
xnor U3174 (N_3174,N_1309,N_1344);
nand U3175 (N_3175,N_1461,N_631);
nor U3176 (N_3176,N_970,N_1746);
nand U3177 (N_3177,N_1389,N_1742);
or U3178 (N_3178,N_991,N_69);
or U3179 (N_3179,N_1257,N_208);
nor U3180 (N_3180,N_1604,N_1785);
and U3181 (N_3181,N_969,N_1421);
and U3182 (N_3182,N_850,N_1314);
nor U3183 (N_3183,N_1932,N_578);
nor U3184 (N_3184,N_1173,N_1668);
nand U3185 (N_3185,N_192,N_307);
nand U3186 (N_3186,N_1672,N_1020);
nor U3187 (N_3187,N_242,N_900);
or U3188 (N_3188,N_1209,N_1704);
or U3189 (N_3189,N_1843,N_743);
nor U3190 (N_3190,N_180,N_1009);
nand U3191 (N_3191,N_653,N_834);
nor U3192 (N_3192,N_1757,N_203);
nand U3193 (N_3193,N_1134,N_1437);
nand U3194 (N_3194,N_568,N_1664);
nor U3195 (N_3195,N_648,N_1413);
nand U3196 (N_3196,N_416,N_1408);
nor U3197 (N_3197,N_435,N_1104);
or U3198 (N_3198,N_1286,N_239);
and U3199 (N_3199,N_980,N_756);
nand U3200 (N_3200,N_1478,N_943);
nand U3201 (N_3201,N_782,N_360);
nor U3202 (N_3202,N_1720,N_579);
nand U3203 (N_3203,N_662,N_850);
nand U3204 (N_3204,N_132,N_1736);
or U3205 (N_3205,N_1579,N_43);
xor U3206 (N_3206,N_581,N_1401);
nor U3207 (N_3207,N_936,N_579);
or U3208 (N_3208,N_61,N_442);
nand U3209 (N_3209,N_974,N_583);
nand U3210 (N_3210,N_267,N_139);
or U3211 (N_3211,N_241,N_372);
nand U3212 (N_3212,N_833,N_710);
or U3213 (N_3213,N_955,N_915);
nand U3214 (N_3214,N_287,N_1689);
or U3215 (N_3215,N_759,N_700);
nand U3216 (N_3216,N_696,N_1829);
and U3217 (N_3217,N_1779,N_435);
nand U3218 (N_3218,N_1321,N_296);
or U3219 (N_3219,N_769,N_894);
nand U3220 (N_3220,N_1264,N_446);
nand U3221 (N_3221,N_864,N_1478);
and U3222 (N_3222,N_357,N_1308);
and U3223 (N_3223,N_937,N_1057);
nand U3224 (N_3224,N_1984,N_902);
xor U3225 (N_3225,N_712,N_1662);
nor U3226 (N_3226,N_1078,N_1110);
xnor U3227 (N_3227,N_1091,N_1172);
nor U3228 (N_3228,N_347,N_1206);
nor U3229 (N_3229,N_875,N_145);
nand U3230 (N_3230,N_1571,N_808);
nand U3231 (N_3231,N_39,N_1109);
or U3232 (N_3232,N_1101,N_300);
nand U3233 (N_3233,N_138,N_1952);
and U3234 (N_3234,N_1324,N_77);
or U3235 (N_3235,N_67,N_1534);
and U3236 (N_3236,N_1509,N_114);
nand U3237 (N_3237,N_1514,N_1440);
nor U3238 (N_3238,N_927,N_196);
or U3239 (N_3239,N_308,N_795);
and U3240 (N_3240,N_835,N_1627);
nor U3241 (N_3241,N_68,N_1081);
and U3242 (N_3242,N_1225,N_1999);
nor U3243 (N_3243,N_169,N_402);
and U3244 (N_3244,N_1934,N_1314);
nor U3245 (N_3245,N_1886,N_1469);
nor U3246 (N_3246,N_1189,N_298);
or U3247 (N_3247,N_959,N_1125);
and U3248 (N_3248,N_271,N_1131);
or U3249 (N_3249,N_856,N_1542);
or U3250 (N_3250,N_359,N_1841);
nor U3251 (N_3251,N_491,N_402);
and U3252 (N_3252,N_1850,N_1420);
and U3253 (N_3253,N_402,N_1898);
nand U3254 (N_3254,N_941,N_749);
and U3255 (N_3255,N_1874,N_1714);
nor U3256 (N_3256,N_1716,N_335);
and U3257 (N_3257,N_218,N_1671);
xor U3258 (N_3258,N_1078,N_1746);
xor U3259 (N_3259,N_931,N_183);
or U3260 (N_3260,N_407,N_1102);
or U3261 (N_3261,N_1144,N_934);
and U3262 (N_3262,N_1921,N_1973);
or U3263 (N_3263,N_1534,N_1879);
nand U3264 (N_3264,N_1956,N_260);
or U3265 (N_3265,N_451,N_1804);
or U3266 (N_3266,N_372,N_0);
or U3267 (N_3267,N_1497,N_622);
and U3268 (N_3268,N_500,N_833);
nand U3269 (N_3269,N_936,N_221);
or U3270 (N_3270,N_195,N_688);
and U3271 (N_3271,N_1790,N_536);
nor U3272 (N_3272,N_1689,N_817);
nor U3273 (N_3273,N_631,N_3);
nand U3274 (N_3274,N_342,N_461);
nor U3275 (N_3275,N_1316,N_724);
xor U3276 (N_3276,N_955,N_1472);
nor U3277 (N_3277,N_1448,N_900);
xor U3278 (N_3278,N_1806,N_1298);
nor U3279 (N_3279,N_1506,N_224);
or U3280 (N_3280,N_57,N_1229);
nand U3281 (N_3281,N_1324,N_1145);
nor U3282 (N_3282,N_28,N_86);
nor U3283 (N_3283,N_1408,N_1002);
and U3284 (N_3284,N_171,N_1652);
and U3285 (N_3285,N_472,N_88);
xnor U3286 (N_3286,N_1808,N_24);
nand U3287 (N_3287,N_1213,N_1394);
nand U3288 (N_3288,N_1464,N_563);
nand U3289 (N_3289,N_1949,N_1618);
nand U3290 (N_3290,N_536,N_421);
or U3291 (N_3291,N_1855,N_1423);
nor U3292 (N_3292,N_73,N_1319);
or U3293 (N_3293,N_1012,N_1715);
nor U3294 (N_3294,N_148,N_1741);
nand U3295 (N_3295,N_665,N_1683);
and U3296 (N_3296,N_1825,N_1338);
and U3297 (N_3297,N_1197,N_369);
nor U3298 (N_3298,N_1909,N_988);
nor U3299 (N_3299,N_1018,N_1407);
or U3300 (N_3300,N_1228,N_66);
nand U3301 (N_3301,N_683,N_1998);
nand U3302 (N_3302,N_980,N_527);
nor U3303 (N_3303,N_1731,N_222);
nor U3304 (N_3304,N_371,N_530);
nor U3305 (N_3305,N_1116,N_1547);
xnor U3306 (N_3306,N_1886,N_1829);
nand U3307 (N_3307,N_1555,N_763);
or U3308 (N_3308,N_1278,N_1757);
nor U3309 (N_3309,N_318,N_1372);
nor U3310 (N_3310,N_1873,N_1695);
and U3311 (N_3311,N_1709,N_160);
nor U3312 (N_3312,N_1960,N_847);
or U3313 (N_3313,N_1846,N_158);
or U3314 (N_3314,N_72,N_836);
nand U3315 (N_3315,N_1519,N_1259);
and U3316 (N_3316,N_1111,N_161);
or U3317 (N_3317,N_1728,N_590);
and U3318 (N_3318,N_1221,N_1349);
nand U3319 (N_3319,N_1730,N_24);
nor U3320 (N_3320,N_1913,N_47);
nor U3321 (N_3321,N_28,N_425);
xnor U3322 (N_3322,N_709,N_1555);
or U3323 (N_3323,N_646,N_1685);
xor U3324 (N_3324,N_1964,N_809);
and U3325 (N_3325,N_1501,N_86);
xnor U3326 (N_3326,N_392,N_309);
and U3327 (N_3327,N_429,N_588);
and U3328 (N_3328,N_920,N_1851);
or U3329 (N_3329,N_1437,N_592);
and U3330 (N_3330,N_1574,N_715);
or U3331 (N_3331,N_476,N_315);
and U3332 (N_3332,N_720,N_195);
and U3333 (N_3333,N_973,N_1330);
or U3334 (N_3334,N_174,N_772);
or U3335 (N_3335,N_1272,N_1853);
or U3336 (N_3336,N_1952,N_886);
or U3337 (N_3337,N_1944,N_1761);
nand U3338 (N_3338,N_266,N_1942);
nand U3339 (N_3339,N_1302,N_1702);
nand U3340 (N_3340,N_724,N_622);
nor U3341 (N_3341,N_936,N_1137);
and U3342 (N_3342,N_554,N_661);
or U3343 (N_3343,N_1985,N_476);
and U3344 (N_3344,N_710,N_1363);
or U3345 (N_3345,N_336,N_831);
and U3346 (N_3346,N_1529,N_409);
nand U3347 (N_3347,N_174,N_1907);
and U3348 (N_3348,N_580,N_1616);
or U3349 (N_3349,N_558,N_1545);
nand U3350 (N_3350,N_241,N_1086);
and U3351 (N_3351,N_1465,N_802);
nand U3352 (N_3352,N_715,N_339);
nand U3353 (N_3353,N_1141,N_1402);
nand U3354 (N_3354,N_1298,N_173);
nor U3355 (N_3355,N_943,N_1397);
and U3356 (N_3356,N_514,N_756);
and U3357 (N_3357,N_563,N_1747);
xnor U3358 (N_3358,N_1640,N_951);
nand U3359 (N_3359,N_1619,N_1729);
or U3360 (N_3360,N_1459,N_171);
or U3361 (N_3361,N_261,N_1900);
nand U3362 (N_3362,N_626,N_672);
nor U3363 (N_3363,N_1053,N_1946);
nor U3364 (N_3364,N_852,N_37);
nor U3365 (N_3365,N_1067,N_356);
xor U3366 (N_3366,N_39,N_1858);
nor U3367 (N_3367,N_797,N_1090);
xnor U3368 (N_3368,N_1515,N_574);
and U3369 (N_3369,N_552,N_1458);
nand U3370 (N_3370,N_1554,N_465);
xnor U3371 (N_3371,N_1600,N_59);
and U3372 (N_3372,N_1155,N_981);
or U3373 (N_3373,N_319,N_1665);
xnor U3374 (N_3374,N_302,N_1606);
or U3375 (N_3375,N_1095,N_399);
xor U3376 (N_3376,N_814,N_613);
xnor U3377 (N_3377,N_987,N_536);
nor U3378 (N_3378,N_168,N_945);
or U3379 (N_3379,N_420,N_1502);
or U3380 (N_3380,N_576,N_1371);
or U3381 (N_3381,N_1366,N_992);
nor U3382 (N_3382,N_1275,N_1904);
nand U3383 (N_3383,N_668,N_1250);
and U3384 (N_3384,N_119,N_1408);
nand U3385 (N_3385,N_1467,N_1657);
nand U3386 (N_3386,N_1700,N_1204);
or U3387 (N_3387,N_1664,N_1764);
or U3388 (N_3388,N_254,N_211);
nor U3389 (N_3389,N_1347,N_1242);
xnor U3390 (N_3390,N_1566,N_864);
or U3391 (N_3391,N_1794,N_1002);
nand U3392 (N_3392,N_1731,N_1451);
nand U3393 (N_3393,N_457,N_979);
nand U3394 (N_3394,N_1798,N_346);
nor U3395 (N_3395,N_831,N_1365);
nand U3396 (N_3396,N_817,N_1215);
nand U3397 (N_3397,N_1879,N_1236);
or U3398 (N_3398,N_260,N_528);
and U3399 (N_3399,N_725,N_78);
and U3400 (N_3400,N_1907,N_880);
and U3401 (N_3401,N_986,N_1615);
nor U3402 (N_3402,N_1774,N_871);
nor U3403 (N_3403,N_305,N_1937);
or U3404 (N_3404,N_1663,N_301);
xnor U3405 (N_3405,N_1482,N_1732);
nand U3406 (N_3406,N_267,N_855);
or U3407 (N_3407,N_1166,N_381);
xnor U3408 (N_3408,N_847,N_1970);
and U3409 (N_3409,N_715,N_1984);
xor U3410 (N_3410,N_797,N_377);
nand U3411 (N_3411,N_311,N_126);
or U3412 (N_3412,N_1242,N_1844);
nor U3413 (N_3413,N_1518,N_1003);
nand U3414 (N_3414,N_841,N_1673);
or U3415 (N_3415,N_103,N_343);
or U3416 (N_3416,N_1456,N_667);
and U3417 (N_3417,N_1435,N_630);
or U3418 (N_3418,N_1595,N_1425);
nor U3419 (N_3419,N_1353,N_574);
and U3420 (N_3420,N_904,N_1466);
xor U3421 (N_3421,N_336,N_484);
xnor U3422 (N_3422,N_989,N_731);
and U3423 (N_3423,N_1140,N_993);
and U3424 (N_3424,N_1647,N_1393);
xor U3425 (N_3425,N_634,N_790);
nand U3426 (N_3426,N_567,N_1269);
or U3427 (N_3427,N_214,N_1474);
and U3428 (N_3428,N_1243,N_709);
nor U3429 (N_3429,N_1248,N_1809);
xnor U3430 (N_3430,N_38,N_974);
or U3431 (N_3431,N_318,N_159);
nor U3432 (N_3432,N_723,N_989);
or U3433 (N_3433,N_454,N_1883);
or U3434 (N_3434,N_200,N_485);
and U3435 (N_3435,N_1593,N_1553);
or U3436 (N_3436,N_1415,N_911);
nand U3437 (N_3437,N_1366,N_329);
nor U3438 (N_3438,N_1610,N_194);
nand U3439 (N_3439,N_523,N_1887);
and U3440 (N_3440,N_1164,N_368);
or U3441 (N_3441,N_21,N_1530);
and U3442 (N_3442,N_1447,N_1792);
or U3443 (N_3443,N_675,N_1528);
nor U3444 (N_3444,N_646,N_882);
xnor U3445 (N_3445,N_883,N_1645);
nor U3446 (N_3446,N_1397,N_987);
or U3447 (N_3447,N_589,N_1591);
and U3448 (N_3448,N_1190,N_1867);
or U3449 (N_3449,N_1311,N_223);
nand U3450 (N_3450,N_1270,N_1819);
xnor U3451 (N_3451,N_1342,N_1973);
xnor U3452 (N_3452,N_1568,N_518);
nand U3453 (N_3453,N_370,N_1571);
and U3454 (N_3454,N_991,N_997);
or U3455 (N_3455,N_1943,N_1013);
nor U3456 (N_3456,N_350,N_1618);
nand U3457 (N_3457,N_1855,N_1159);
nand U3458 (N_3458,N_83,N_1417);
or U3459 (N_3459,N_512,N_890);
xnor U3460 (N_3460,N_1003,N_207);
nand U3461 (N_3461,N_783,N_1436);
xnor U3462 (N_3462,N_1040,N_1618);
nor U3463 (N_3463,N_1124,N_523);
nand U3464 (N_3464,N_1674,N_1832);
nor U3465 (N_3465,N_618,N_1316);
nand U3466 (N_3466,N_654,N_816);
nand U3467 (N_3467,N_952,N_782);
and U3468 (N_3468,N_1857,N_1107);
and U3469 (N_3469,N_1360,N_222);
and U3470 (N_3470,N_732,N_1451);
or U3471 (N_3471,N_1132,N_1201);
and U3472 (N_3472,N_626,N_1096);
xor U3473 (N_3473,N_1113,N_1760);
and U3474 (N_3474,N_1888,N_1398);
or U3475 (N_3475,N_1470,N_1575);
and U3476 (N_3476,N_1963,N_67);
and U3477 (N_3477,N_1339,N_1799);
or U3478 (N_3478,N_91,N_569);
nand U3479 (N_3479,N_1014,N_1677);
xnor U3480 (N_3480,N_1301,N_1641);
or U3481 (N_3481,N_1537,N_499);
and U3482 (N_3482,N_1715,N_1418);
nor U3483 (N_3483,N_436,N_1262);
nor U3484 (N_3484,N_1044,N_385);
xor U3485 (N_3485,N_1512,N_1572);
and U3486 (N_3486,N_1903,N_395);
xnor U3487 (N_3487,N_1824,N_1278);
or U3488 (N_3488,N_1244,N_1555);
nor U3489 (N_3489,N_677,N_703);
or U3490 (N_3490,N_1638,N_562);
xnor U3491 (N_3491,N_1064,N_1336);
nor U3492 (N_3492,N_278,N_529);
nand U3493 (N_3493,N_880,N_28);
nand U3494 (N_3494,N_1264,N_1426);
and U3495 (N_3495,N_427,N_1377);
and U3496 (N_3496,N_1938,N_1002);
and U3497 (N_3497,N_125,N_370);
nand U3498 (N_3498,N_1339,N_796);
and U3499 (N_3499,N_1052,N_984);
nand U3500 (N_3500,N_309,N_228);
xor U3501 (N_3501,N_1068,N_366);
xnor U3502 (N_3502,N_1016,N_525);
nand U3503 (N_3503,N_1183,N_1786);
xor U3504 (N_3504,N_773,N_881);
nand U3505 (N_3505,N_332,N_1294);
or U3506 (N_3506,N_944,N_186);
nor U3507 (N_3507,N_1224,N_1270);
or U3508 (N_3508,N_49,N_587);
nor U3509 (N_3509,N_1665,N_124);
nand U3510 (N_3510,N_593,N_23);
nand U3511 (N_3511,N_517,N_184);
nor U3512 (N_3512,N_1698,N_1123);
xnor U3513 (N_3513,N_1681,N_503);
nand U3514 (N_3514,N_371,N_643);
or U3515 (N_3515,N_919,N_1472);
nor U3516 (N_3516,N_101,N_1712);
nand U3517 (N_3517,N_1106,N_1257);
and U3518 (N_3518,N_598,N_1945);
and U3519 (N_3519,N_1047,N_502);
nor U3520 (N_3520,N_1886,N_1152);
or U3521 (N_3521,N_1829,N_739);
and U3522 (N_3522,N_791,N_292);
or U3523 (N_3523,N_1910,N_1699);
nand U3524 (N_3524,N_1143,N_927);
nor U3525 (N_3525,N_167,N_800);
nor U3526 (N_3526,N_310,N_1179);
or U3527 (N_3527,N_1956,N_89);
or U3528 (N_3528,N_1932,N_503);
and U3529 (N_3529,N_1499,N_1264);
nand U3530 (N_3530,N_1521,N_1402);
or U3531 (N_3531,N_1197,N_956);
and U3532 (N_3532,N_1698,N_59);
or U3533 (N_3533,N_1530,N_1710);
and U3534 (N_3534,N_80,N_1404);
nand U3535 (N_3535,N_1477,N_1608);
and U3536 (N_3536,N_717,N_1639);
nor U3537 (N_3537,N_259,N_936);
and U3538 (N_3538,N_1426,N_1168);
nand U3539 (N_3539,N_1450,N_738);
nor U3540 (N_3540,N_1839,N_896);
xor U3541 (N_3541,N_1511,N_24);
nand U3542 (N_3542,N_1593,N_846);
or U3543 (N_3543,N_1146,N_1403);
or U3544 (N_3544,N_1689,N_508);
and U3545 (N_3545,N_895,N_1786);
and U3546 (N_3546,N_132,N_434);
nor U3547 (N_3547,N_888,N_1984);
xor U3548 (N_3548,N_1159,N_1104);
xnor U3549 (N_3549,N_1811,N_515);
nand U3550 (N_3550,N_1910,N_918);
nor U3551 (N_3551,N_1625,N_635);
nor U3552 (N_3552,N_717,N_1777);
nor U3553 (N_3553,N_984,N_1061);
or U3554 (N_3554,N_986,N_967);
or U3555 (N_3555,N_700,N_55);
nand U3556 (N_3556,N_1262,N_797);
or U3557 (N_3557,N_1470,N_1423);
and U3558 (N_3558,N_1747,N_265);
nand U3559 (N_3559,N_125,N_37);
and U3560 (N_3560,N_1777,N_1826);
or U3561 (N_3561,N_1119,N_495);
nor U3562 (N_3562,N_1353,N_69);
nand U3563 (N_3563,N_1801,N_1268);
nor U3564 (N_3564,N_1953,N_664);
and U3565 (N_3565,N_1207,N_1397);
nor U3566 (N_3566,N_772,N_1409);
and U3567 (N_3567,N_336,N_944);
and U3568 (N_3568,N_597,N_1821);
nand U3569 (N_3569,N_1613,N_632);
nor U3570 (N_3570,N_1151,N_728);
nor U3571 (N_3571,N_1883,N_94);
and U3572 (N_3572,N_1643,N_42);
and U3573 (N_3573,N_1246,N_1568);
nor U3574 (N_3574,N_667,N_110);
nor U3575 (N_3575,N_1122,N_1712);
nor U3576 (N_3576,N_1612,N_1405);
and U3577 (N_3577,N_687,N_1699);
and U3578 (N_3578,N_1571,N_341);
nor U3579 (N_3579,N_701,N_733);
and U3580 (N_3580,N_1346,N_1942);
or U3581 (N_3581,N_1889,N_559);
nor U3582 (N_3582,N_1176,N_1026);
or U3583 (N_3583,N_1251,N_211);
nor U3584 (N_3584,N_627,N_846);
nor U3585 (N_3585,N_1230,N_591);
or U3586 (N_3586,N_557,N_1829);
nand U3587 (N_3587,N_1931,N_252);
nand U3588 (N_3588,N_953,N_629);
and U3589 (N_3589,N_1923,N_1791);
or U3590 (N_3590,N_749,N_330);
nand U3591 (N_3591,N_289,N_1320);
and U3592 (N_3592,N_1958,N_215);
or U3593 (N_3593,N_1750,N_1933);
nor U3594 (N_3594,N_789,N_9);
or U3595 (N_3595,N_1733,N_1206);
or U3596 (N_3596,N_1215,N_1406);
or U3597 (N_3597,N_215,N_1905);
nand U3598 (N_3598,N_422,N_1768);
nand U3599 (N_3599,N_1955,N_1559);
nor U3600 (N_3600,N_325,N_1995);
or U3601 (N_3601,N_1792,N_906);
nor U3602 (N_3602,N_1113,N_1074);
nand U3603 (N_3603,N_1547,N_803);
or U3604 (N_3604,N_517,N_1112);
nor U3605 (N_3605,N_108,N_814);
or U3606 (N_3606,N_1996,N_835);
and U3607 (N_3607,N_821,N_375);
or U3608 (N_3608,N_725,N_557);
and U3609 (N_3609,N_1200,N_1264);
or U3610 (N_3610,N_1431,N_339);
or U3611 (N_3611,N_1653,N_1675);
and U3612 (N_3612,N_500,N_1600);
xor U3613 (N_3613,N_696,N_432);
nand U3614 (N_3614,N_1872,N_1842);
and U3615 (N_3615,N_1545,N_894);
or U3616 (N_3616,N_694,N_903);
and U3617 (N_3617,N_886,N_407);
and U3618 (N_3618,N_1771,N_1239);
and U3619 (N_3619,N_1768,N_244);
nor U3620 (N_3620,N_1584,N_951);
xnor U3621 (N_3621,N_190,N_1341);
nand U3622 (N_3622,N_1324,N_1090);
and U3623 (N_3623,N_1424,N_220);
or U3624 (N_3624,N_327,N_1329);
nand U3625 (N_3625,N_729,N_161);
nor U3626 (N_3626,N_1278,N_932);
nor U3627 (N_3627,N_1563,N_40);
nor U3628 (N_3628,N_868,N_795);
nor U3629 (N_3629,N_1474,N_714);
nand U3630 (N_3630,N_1323,N_62);
or U3631 (N_3631,N_1191,N_1309);
or U3632 (N_3632,N_1570,N_98);
nor U3633 (N_3633,N_1343,N_1791);
nor U3634 (N_3634,N_1616,N_1770);
and U3635 (N_3635,N_1701,N_367);
nand U3636 (N_3636,N_46,N_1342);
xnor U3637 (N_3637,N_1497,N_1260);
xnor U3638 (N_3638,N_544,N_1309);
or U3639 (N_3639,N_493,N_1177);
nor U3640 (N_3640,N_57,N_23);
or U3641 (N_3641,N_1551,N_372);
nor U3642 (N_3642,N_561,N_1088);
nor U3643 (N_3643,N_121,N_1930);
nand U3644 (N_3644,N_1738,N_18);
nand U3645 (N_3645,N_1407,N_106);
nand U3646 (N_3646,N_983,N_919);
xnor U3647 (N_3647,N_558,N_643);
and U3648 (N_3648,N_611,N_831);
nor U3649 (N_3649,N_1649,N_532);
and U3650 (N_3650,N_594,N_955);
and U3651 (N_3651,N_868,N_195);
and U3652 (N_3652,N_1287,N_1221);
nand U3653 (N_3653,N_1503,N_315);
xnor U3654 (N_3654,N_544,N_881);
nand U3655 (N_3655,N_1084,N_622);
and U3656 (N_3656,N_1888,N_1610);
nand U3657 (N_3657,N_1017,N_766);
nand U3658 (N_3658,N_588,N_320);
and U3659 (N_3659,N_23,N_230);
xor U3660 (N_3660,N_486,N_522);
and U3661 (N_3661,N_455,N_1540);
xnor U3662 (N_3662,N_1872,N_36);
and U3663 (N_3663,N_1257,N_308);
or U3664 (N_3664,N_1837,N_0);
and U3665 (N_3665,N_325,N_313);
nor U3666 (N_3666,N_558,N_308);
nand U3667 (N_3667,N_318,N_302);
nand U3668 (N_3668,N_972,N_228);
nor U3669 (N_3669,N_544,N_1258);
or U3670 (N_3670,N_1726,N_1071);
and U3671 (N_3671,N_933,N_1343);
or U3672 (N_3672,N_1040,N_567);
and U3673 (N_3673,N_76,N_876);
nor U3674 (N_3674,N_573,N_1033);
and U3675 (N_3675,N_856,N_1804);
nand U3676 (N_3676,N_1535,N_1540);
and U3677 (N_3677,N_439,N_1543);
and U3678 (N_3678,N_130,N_435);
and U3679 (N_3679,N_1336,N_1465);
xor U3680 (N_3680,N_677,N_1230);
nor U3681 (N_3681,N_963,N_133);
nand U3682 (N_3682,N_125,N_404);
nor U3683 (N_3683,N_1462,N_1760);
nand U3684 (N_3684,N_1394,N_15);
nor U3685 (N_3685,N_1371,N_793);
nor U3686 (N_3686,N_326,N_343);
nor U3687 (N_3687,N_1396,N_178);
nand U3688 (N_3688,N_1403,N_343);
nor U3689 (N_3689,N_1057,N_168);
or U3690 (N_3690,N_1940,N_588);
or U3691 (N_3691,N_1284,N_623);
nand U3692 (N_3692,N_1609,N_1627);
xor U3693 (N_3693,N_1380,N_834);
or U3694 (N_3694,N_239,N_940);
or U3695 (N_3695,N_123,N_602);
nand U3696 (N_3696,N_985,N_1360);
or U3697 (N_3697,N_630,N_629);
nor U3698 (N_3698,N_1854,N_591);
nor U3699 (N_3699,N_1851,N_1638);
nor U3700 (N_3700,N_1867,N_1363);
and U3701 (N_3701,N_904,N_1600);
and U3702 (N_3702,N_1235,N_698);
xor U3703 (N_3703,N_85,N_782);
nand U3704 (N_3704,N_97,N_313);
nor U3705 (N_3705,N_1526,N_1669);
and U3706 (N_3706,N_1472,N_805);
or U3707 (N_3707,N_1848,N_1797);
or U3708 (N_3708,N_1234,N_140);
or U3709 (N_3709,N_1209,N_731);
xor U3710 (N_3710,N_147,N_1096);
nor U3711 (N_3711,N_488,N_1520);
and U3712 (N_3712,N_81,N_1614);
or U3713 (N_3713,N_1043,N_390);
and U3714 (N_3714,N_317,N_9);
xor U3715 (N_3715,N_643,N_615);
nor U3716 (N_3716,N_257,N_1801);
or U3717 (N_3717,N_227,N_363);
nor U3718 (N_3718,N_1175,N_400);
nand U3719 (N_3719,N_1733,N_403);
nor U3720 (N_3720,N_341,N_945);
and U3721 (N_3721,N_1997,N_717);
and U3722 (N_3722,N_1883,N_1454);
or U3723 (N_3723,N_296,N_1105);
and U3724 (N_3724,N_1459,N_1850);
nor U3725 (N_3725,N_255,N_65);
or U3726 (N_3726,N_1788,N_1515);
or U3727 (N_3727,N_1402,N_406);
and U3728 (N_3728,N_1226,N_847);
nor U3729 (N_3729,N_185,N_1324);
and U3730 (N_3730,N_1143,N_977);
and U3731 (N_3731,N_1153,N_819);
and U3732 (N_3732,N_87,N_1550);
or U3733 (N_3733,N_137,N_1529);
xor U3734 (N_3734,N_862,N_1979);
or U3735 (N_3735,N_1531,N_1916);
nor U3736 (N_3736,N_1819,N_47);
nor U3737 (N_3737,N_594,N_1242);
xnor U3738 (N_3738,N_470,N_1054);
and U3739 (N_3739,N_479,N_446);
nor U3740 (N_3740,N_209,N_1280);
and U3741 (N_3741,N_798,N_147);
or U3742 (N_3742,N_1830,N_1085);
nand U3743 (N_3743,N_171,N_1430);
xor U3744 (N_3744,N_692,N_604);
and U3745 (N_3745,N_1409,N_1498);
nor U3746 (N_3746,N_200,N_382);
nor U3747 (N_3747,N_1304,N_761);
and U3748 (N_3748,N_257,N_1577);
nand U3749 (N_3749,N_1523,N_1467);
and U3750 (N_3750,N_332,N_1784);
or U3751 (N_3751,N_1071,N_1143);
or U3752 (N_3752,N_842,N_180);
nor U3753 (N_3753,N_564,N_1914);
nand U3754 (N_3754,N_541,N_1464);
or U3755 (N_3755,N_1482,N_1207);
and U3756 (N_3756,N_1921,N_1644);
and U3757 (N_3757,N_1042,N_213);
and U3758 (N_3758,N_758,N_52);
nand U3759 (N_3759,N_1272,N_1093);
and U3760 (N_3760,N_1022,N_720);
or U3761 (N_3761,N_1710,N_253);
nor U3762 (N_3762,N_499,N_675);
nor U3763 (N_3763,N_145,N_1646);
or U3764 (N_3764,N_294,N_1165);
nor U3765 (N_3765,N_1199,N_982);
or U3766 (N_3766,N_1043,N_1081);
nor U3767 (N_3767,N_1748,N_1346);
xor U3768 (N_3768,N_850,N_469);
and U3769 (N_3769,N_74,N_369);
nand U3770 (N_3770,N_542,N_1168);
or U3771 (N_3771,N_1227,N_28);
nand U3772 (N_3772,N_1447,N_186);
nor U3773 (N_3773,N_891,N_1230);
and U3774 (N_3774,N_85,N_1290);
nor U3775 (N_3775,N_1122,N_926);
nor U3776 (N_3776,N_724,N_781);
nand U3777 (N_3777,N_1686,N_466);
or U3778 (N_3778,N_663,N_545);
nand U3779 (N_3779,N_887,N_387);
and U3780 (N_3780,N_1952,N_1208);
nor U3781 (N_3781,N_1515,N_1145);
nor U3782 (N_3782,N_1706,N_1064);
nand U3783 (N_3783,N_1665,N_41);
nor U3784 (N_3784,N_1267,N_751);
nor U3785 (N_3785,N_867,N_358);
or U3786 (N_3786,N_305,N_733);
nor U3787 (N_3787,N_1369,N_1441);
xnor U3788 (N_3788,N_338,N_1994);
and U3789 (N_3789,N_1817,N_1715);
and U3790 (N_3790,N_1671,N_1894);
nand U3791 (N_3791,N_1038,N_657);
nor U3792 (N_3792,N_58,N_494);
and U3793 (N_3793,N_221,N_1321);
or U3794 (N_3794,N_816,N_1208);
nor U3795 (N_3795,N_1665,N_517);
nor U3796 (N_3796,N_1610,N_1077);
nand U3797 (N_3797,N_258,N_154);
or U3798 (N_3798,N_623,N_856);
nor U3799 (N_3799,N_107,N_1317);
or U3800 (N_3800,N_1609,N_896);
xor U3801 (N_3801,N_1845,N_1842);
and U3802 (N_3802,N_579,N_562);
or U3803 (N_3803,N_1995,N_1634);
or U3804 (N_3804,N_979,N_612);
or U3805 (N_3805,N_382,N_1667);
or U3806 (N_3806,N_929,N_150);
xnor U3807 (N_3807,N_777,N_821);
xnor U3808 (N_3808,N_1489,N_1527);
nand U3809 (N_3809,N_1021,N_589);
nand U3810 (N_3810,N_132,N_1260);
nor U3811 (N_3811,N_204,N_761);
nand U3812 (N_3812,N_177,N_1415);
or U3813 (N_3813,N_481,N_992);
nor U3814 (N_3814,N_1473,N_863);
nor U3815 (N_3815,N_1256,N_852);
or U3816 (N_3816,N_1293,N_1073);
nor U3817 (N_3817,N_1205,N_162);
and U3818 (N_3818,N_1944,N_1641);
nand U3819 (N_3819,N_1519,N_962);
or U3820 (N_3820,N_1331,N_481);
or U3821 (N_3821,N_122,N_681);
nand U3822 (N_3822,N_190,N_1552);
xnor U3823 (N_3823,N_927,N_1462);
nand U3824 (N_3824,N_403,N_1177);
nor U3825 (N_3825,N_177,N_266);
or U3826 (N_3826,N_295,N_1726);
xnor U3827 (N_3827,N_1946,N_1089);
and U3828 (N_3828,N_852,N_1447);
nand U3829 (N_3829,N_622,N_1198);
or U3830 (N_3830,N_762,N_1969);
nor U3831 (N_3831,N_605,N_1783);
xor U3832 (N_3832,N_483,N_1131);
nor U3833 (N_3833,N_474,N_1563);
and U3834 (N_3834,N_930,N_628);
nor U3835 (N_3835,N_1579,N_553);
nor U3836 (N_3836,N_1245,N_1152);
nand U3837 (N_3837,N_1822,N_1313);
or U3838 (N_3838,N_30,N_1431);
nor U3839 (N_3839,N_761,N_645);
xnor U3840 (N_3840,N_1250,N_2);
xor U3841 (N_3841,N_1268,N_184);
nand U3842 (N_3842,N_138,N_12);
and U3843 (N_3843,N_256,N_919);
nand U3844 (N_3844,N_485,N_608);
nand U3845 (N_3845,N_235,N_53);
nor U3846 (N_3846,N_442,N_290);
nand U3847 (N_3847,N_752,N_581);
nor U3848 (N_3848,N_492,N_1432);
nand U3849 (N_3849,N_1850,N_1328);
or U3850 (N_3850,N_95,N_846);
and U3851 (N_3851,N_424,N_475);
and U3852 (N_3852,N_1402,N_41);
nor U3853 (N_3853,N_899,N_1711);
xnor U3854 (N_3854,N_1824,N_249);
or U3855 (N_3855,N_20,N_77);
nand U3856 (N_3856,N_1999,N_1705);
and U3857 (N_3857,N_700,N_1017);
and U3858 (N_3858,N_616,N_492);
or U3859 (N_3859,N_567,N_548);
nand U3860 (N_3860,N_1309,N_294);
and U3861 (N_3861,N_620,N_1063);
nor U3862 (N_3862,N_548,N_1680);
and U3863 (N_3863,N_1782,N_164);
or U3864 (N_3864,N_715,N_1703);
and U3865 (N_3865,N_431,N_361);
and U3866 (N_3866,N_1200,N_988);
and U3867 (N_3867,N_423,N_652);
nand U3868 (N_3868,N_95,N_1482);
nor U3869 (N_3869,N_1344,N_1920);
and U3870 (N_3870,N_170,N_1007);
or U3871 (N_3871,N_568,N_1313);
or U3872 (N_3872,N_1065,N_798);
and U3873 (N_3873,N_402,N_1626);
nor U3874 (N_3874,N_733,N_1152);
nor U3875 (N_3875,N_1740,N_782);
or U3876 (N_3876,N_1125,N_1235);
nor U3877 (N_3877,N_939,N_1069);
nand U3878 (N_3878,N_359,N_133);
nand U3879 (N_3879,N_843,N_1354);
or U3880 (N_3880,N_814,N_47);
or U3881 (N_3881,N_1302,N_821);
xor U3882 (N_3882,N_1256,N_317);
or U3883 (N_3883,N_32,N_355);
nor U3884 (N_3884,N_1832,N_528);
nor U3885 (N_3885,N_1210,N_903);
nand U3886 (N_3886,N_227,N_1407);
nand U3887 (N_3887,N_122,N_1883);
or U3888 (N_3888,N_1571,N_1007);
and U3889 (N_3889,N_1283,N_760);
nor U3890 (N_3890,N_1777,N_457);
and U3891 (N_3891,N_1725,N_1564);
and U3892 (N_3892,N_203,N_1976);
nor U3893 (N_3893,N_1233,N_1387);
nand U3894 (N_3894,N_1906,N_480);
or U3895 (N_3895,N_942,N_1874);
or U3896 (N_3896,N_465,N_1168);
nor U3897 (N_3897,N_986,N_1780);
or U3898 (N_3898,N_501,N_986);
xor U3899 (N_3899,N_725,N_496);
and U3900 (N_3900,N_1317,N_942);
or U3901 (N_3901,N_358,N_85);
or U3902 (N_3902,N_1814,N_833);
or U3903 (N_3903,N_1193,N_1880);
or U3904 (N_3904,N_588,N_1907);
nand U3905 (N_3905,N_1542,N_1523);
nand U3906 (N_3906,N_1326,N_1870);
xnor U3907 (N_3907,N_1212,N_156);
nand U3908 (N_3908,N_1591,N_1618);
or U3909 (N_3909,N_119,N_1184);
nand U3910 (N_3910,N_429,N_394);
and U3911 (N_3911,N_1085,N_1275);
or U3912 (N_3912,N_1809,N_1184);
or U3913 (N_3913,N_825,N_659);
and U3914 (N_3914,N_89,N_1823);
nand U3915 (N_3915,N_975,N_704);
and U3916 (N_3916,N_576,N_820);
nor U3917 (N_3917,N_149,N_923);
or U3918 (N_3918,N_134,N_990);
nand U3919 (N_3919,N_1710,N_302);
xor U3920 (N_3920,N_307,N_696);
or U3921 (N_3921,N_949,N_1186);
nand U3922 (N_3922,N_34,N_1874);
nor U3923 (N_3923,N_228,N_541);
or U3924 (N_3924,N_282,N_1616);
and U3925 (N_3925,N_1461,N_1718);
nor U3926 (N_3926,N_1835,N_364);
nand U3927 (N_3927,N_16,N_629);
or U3928 (N_3928,N_1502,N_1630);
or U3929 (N_3929,N_377,N_1503);
and U3930 (N_3930,N_187,N_363);
nand U3931 (N_3931,N_1775,N_1547);
or U3932 (N_3932,N_1323,N_527);
nand U3933 (N_3933,N_588,N_152);
or U3934 (N_3934,N_239,N_1892);
and U3935 (N_3935,N_1312,N_1809);
nand U3936 (N_3936,N_143,N_895);
nor U3937 (N_3937,N_732,N_1217);
or U3938 (N_3938,N_881,N_1278);
nand U3939 (N_3939,N_1329,N_687);
and U3940 (N_3940,N_1549,N_383);
nand U3941 (N_3941,N_220,N_1878);
or U3942 (N_3942,N_1405,N_499);
nor U3943 (N_3943,N_594,N_160);
xnor U3944 (N_3944,N_39,N_412);
and U3945 (N_3945,N_1804,N_751);
nor U3946 (N_3946,N_214,N_1144);
xor U3947 (N_3947,N_127,N_1646);
nand U3948 (N_3948,N_1051,N_1409);
and U3949 (N_3949,N_1937,N_116);
and U3950 (N_3950,N_861,N_1356);
nor U3951 (N_3951,N_895,N_571);
and U3952 (N_3952,N_1686,N_1086);
nand U3953 (N_3953,N_1332,N_731);
and U3954 (N_3954,N_1135,N_1112);
nor U3955 (N_3955,N_1099,N_1411);
and U3956 (N_3956,N_1574,N_499);
nand U3957 (N_3957,N_1535,N_602);
or U3958 (N_3958,N_414,N_1567);
or U3959 (N_3959,N_1660,N_1173);
nand U3960 (N_3960,N_1868,N_1871);
and U3961 (N_3961,N_462,N_1204);
or U3962 (N_3962,N_825,N_1332);
and U3963 (N_3963,N_662,N_1239);
or U3964 (N_3964,N_295,N_638);
nand U3965 (N_3965,N_1624,N_1838);
or U3966 (N_3966,N_1444,N_1697);
nand U3967 (N_3967,N_1601,N_1014);
nand U3968 (N_3968,N_1150,N_1156);
xnor U3969 (N_3969,N_1646,N_901);
nand U3970 (N_3970,N_691,N_423);
nor U3971 (N_3971,N_517,N_496);
and U3972 (N_3972,N_410,N_1732);
nand U3973 (N_3973,N_815,N_1438);
or U3974 (N_3974,N_1086,N_331);
nand U3975 (N_3975,N_800,N_1111);
and U3976 (N_3976,N_561,N_9);
nor U3977 (N_3977,N_435,N_509);
or U3978 (N_3978,N_348,N_143);
xor U3979 (N_3979,N_321,N_1172);
and U3980 (N_3980,N_835,N_723);
nor U3981 (N_3981,N_876,N_1158);
and U3982 (N_3982,N_762,N_1357);
nand U3983 (N_3983,N_375,N_1128);
nand U3984 (N_3984,N_1573,N_415);
and U3985 (N_3985,N_503,N_1026);
and U3986 (N_3986,N_218,N_334);
nand U3987 (N_3987,N_327,N_1992);
and U3988 (N_3988,N_768,N_723);
nand U3989 (N_3989,N_1725,N_843);
and U3990 (N_3990,N_1919,N_1631);
or U3991 (N_3991,N_1482,N_1781);
and U3992 (N_3992,N_1117,N_959);
nand U3993 (N_3993,N_405,N_1435);
nand U3994 (N_3994,N_1162,N_1397);
or U3995 (N_3995,N_761,N_1585);
nor U3996 (N_3996,N_1140,N_1491);
nand U3997 (N_3997,N_187,N_473);
nor U3998 (N_3998,N_1872,N_630);
nor U3999 (N_3999,N_1763,N_490);
nor U4000 (N_4000,N_3563,N_2469);
nand U4001 (N_4001,N_2180,N_3039);
nor U4002 (N_4002,N_2001,N_3539);
nor U4003 (N_4003,N_3217,N_3013);
and U4004 (N_4004,N_2101,N_3906);
nand U4005 (N_4005,N_3423,N_3114);
and U4006 (N_4006,N_3896,N_3600);
nand U4007 (N_4007,N_2157,N_3538);
nor U4008 (N_4008,N_3993,N_2024);
or U4009 (N_4009,N_2023,N_2031);
and U4010 (N_4010,N_2756,N_2422);
nor U4011 (N_4011,N_2902,N_3406);
nor U4012 (N_4012,N_3016,N_2100);
and U4013 (N_4013,N_3677,N_3527);
and U4014 (N_4014,N_2032,N_2194);
or U4015 (N_4015,N_2733,N_3089);
nor U4016 (N_4016,N_3831,N_2563);
nand U4017 (N_4017,N_2554,N_2729);
and U4018 (N_4018,N_2982,N_3657);
or U4019 (N_4019,N_3220,N_2235);
xnor U4020 (N_4020,N_3707,N_2213);
nand U4021 (N_4021,N_3366,N_2126);
nand U4022 (N_4022,N_2183,N_2285);
nand U4023 (N_4023,N_3582,N_3259);
and U4024 (N_4024,N_2717,N_2437);
and U4025 (N_4025,N_3065,N_3172);
and U4026 (N_4026,N_2116,N_2106);
and U4027 (N_4027,N_3303,N_2022);
or U4028 (N_4028,N_3273,N_3736);
and U4029 (N_4029,N_3353,N_3085);
or U4030 (N_4030,N_2340,N_2341);
or U4031 (N_4031,N_2476,N_3441);
nor U4032 (N_4032,N_2866,N_2491);
or U4033 (N_4033,N_2278,N_2042);
nand U4034 (N_4034,N_2887,N_2929);
and U4035 (N_4035,N_3115,N_2244);
nor U4036 (N_4036,N_2417,N_3876);
nand U4037 (N_4037,N_3669,N_3730);
and U4038 (N_4038,N_2710,N_2080);
xor U4039 (N_4039,N_2908,N_3358);
or U4040 (N_4040,N_2072,N_2938);
nor U4041 (N_4041,N_3087,N_2184);
xor U4042 (N_4042,N_2538,N_2452);
and U4043 (N_4043,N_2438,N_3910);
nor U4044 (N_4044,N_2348,N_2674);
or U4045 (N_4045,N_3569,N_3307);
and U4046 (N_4046,N_2609,N_3175);
and U4047 (N_4047,N_2245,N_2036);
nand U4048 (N_4048,N_3651,N_2696);
and U4049 (N_4049,N_2718,N_2127);
xnor U4050 (N_4050,N_3544,N_3478);
xnor U4051 (N_4051,N_3425,N_3477);
or U4052 (N_4052,N_2309,N_3103);
and U4053 (N_4053,N_3191,N_2344);
or U4054 (N_4054,N_2946,N_3480);
nand U4055 (N_4055,N_3891,N_2702);
or U4056 (N_4056,N_3324,N_3607);
nor U4057 (N_4057,N_2648,N_3095);
or U4058 (N_4058,N_2257,N_2201);
nand U4059 (N_4059,N_3380,N_2809);
or U4060 (N_4060,N_3225,N_3633);
xor U4061 (N_4061,N_2588,N_2470);
and U4062 (N_4062,N_3289,N_3858);
or U4063 (N_4063,N_2744,N_3928);
nand U4064 (N_4064,N_3755,N_2816);
or U4065 (N_4065,N_2271,N_3862);
or U4066 (N_4066,N_2955,N_3310);
nand U4067 (N_4067,N_3568,N_2292);
or U4068 (N_4068,N_3720,N_2658);
nor U4069 (N_4069,N_3552,N_2727);
nor U4070 (N_4070,N_2950,N_2583);
and U4071 (N_4071,N_2843,N_3258);
or U4072 (N_4072,N_3336,N_3378);
nor U4073 (N_4073,N_2377,N_2226);
and U4074 (N_4074,N_3968,N_2640);
or U4075 (N_4075,N_2220,N_3393);
and U4076 (N_4076,N_3705,N_3141);
nand U4077 (N_4077,N_3589,N_2364);
nor U4078 (N_4078,N_2992,N_2343);
and U4079 (N_4079,N_3464,N_2801);
nand U4080 (N_4080,N_3710,N_3841);
nand U4081 (N_4081,N_3404,N_2014);
nand U4082 (N_4082,N_2794,N_3124);
and U4083 (N_4083,N_2769,N_3835);
and U4084 (N_4084,N_2597,N_3966);
nand U4085 (N_4085,N_2082,N_2302);
or U4086 (N_4086,N_3543,N_2639);
nand U4087 (N_4087,N_3496,N_2954);
nand U4088 (N_4088,N_3032,N_3011);
nor U4089 (N_4089,N_2547,N_2517);
and U4090 (N_4090,N_2252,N_2686);
and U4091 (N_4091,N_3436,N_2709);
and U4092 (N_4092,N_2124,N_3239);
nor U4093 (N_4093,N_2839,N_3861);
xnor U4094 (N_4094,N_2990,N_3186);
nand U4095 (N_4095,N_2301,N_2649);
nand U4096 (N_4096,N_3675,N_3322);
or U4097 (N_4097,N_2111,N_3402);
nand U4098 (N_4098,N_2961,N_3774);
and U4099 (N_4099,N_2055,N_3793);
and U4100 (N_4100,N_2172,N_2638);
or U4101 (N_4101,N_3298,N_3714);
nor U4102 (N_4102,N_2948,N_2320);
or U4103 (N_4103,N_3929,N_3679);
and U4104 (N_4104,N_3510,N_2295);
and U4105 (N_4105,N_2490,N_2534);
nand U4106 (N_4106,N_2539,N_3961);
nand U4107 (N_4107,N_2618,N_2749);
and U4108 (N_4108,N_3129,N_2380);
nand U4109 (N_4109,N_3903,N_3266);
and U4110 (N_4110,N_3706,N_2813);
xnor U4111 (N_4111,N_2240,N_2643);
xor U4112 (N_4112,N_2305,N_2137);
xnor U4113 (N_4113,N_2266,N_2726);
nor U4114 (N_4114,N_2976,N_3960);
nand U4115 (N_4115,N_3078,N_3069);
or U4116 (N_4116,N_2317,N_3799);
and U4117 (N_4117,N_3357,N_3387);
and U4118 (N_4118,N_3160,N_2342);
or U4119 (N_4119,N_2028,N_3711);
nor U4120 (N_4120,N_2712,N_2013);
nor U4121 (N_4121,N_3019,N_3138);
and U4122 (N_4122,N_2963,N_3098);
nand U4123 (N_4123,N_3970,N_2551);
nand U4124 (N_4124,N_3434,N_2019);
or U4125 (N_4125,N_3269,N_3738);
or U4126 (N_4126,N_2384,N_2874);
nor U4127 (N_4127,N_2141,N_3549);
xor U4128 (N_4128,N_3853,N_3609);
nor U4129 (N_4129,N_2969,N_3665);
xnor U4130 (N_4130,N_2468,N_2943);
and U4131 (N_4131,N_3979,N_2251);
nand U4132 (N_4132,N_3066,N_3652);
nand U4133 (N_4133,N_3777,N_3666);
and U4134 (N_4134,N_3384,N_3830);
nand U4135 (N_4135,N_2993,N_3847);
or U4136 (N_4136,N_3163,N_2270);
and U4137 (N_4137,N_2409,N_2390);
and U4138 (N_4138,N_2817,N_2450);
nand U4139 (N_4139,N_2329,N_3060);
and U4140 (N_4140,N_2457,N_2569);
nor U4141 (N_4141,N_3494,N_2617);
or U4142 (N_4142,N_2176,N_3005);
nand U4143 (N_4143,N_2314,N_2647);
or U4144 (N_4144,N_3673,N_3629);
nand U4145 (N_4145,N_3224,N_2178);
or U4146 (N_4146,N_3886,N_2393);
nand U4147 (N_4147,N_2782,N_3797);
nand U4148 (N_4148,N_3389,N_3654);
nand U4149 (N_4149,N_2060,N_2766);
xor U4150 (N_4150,N_2406,N_3004);
or U4151 (N_4151,N_2949,N_2692);
or U4152 (N_4152,N_3828,N_3940);
nor U4153 (N_4153,N_3603,N_3430);
nand U4154 (N_4154,N_3709,N_2134);
and U4155 (N_4155,N_2510,N_2966);
nor U4156 (N_4156,N_3048,N_2246);
or U4157 (N_4157,N_3139,N_2935);
or U4158 (N_4158,N_2977,N_2304);
nand U4159 (N_4159,N_2502,N_3216);
nand U4160 (N_4160,N_3306,N_3758);
nand U4161 (N_4161,N_2919,N_2795);
nand U4162 (N_4162,N_2392,N_2722);
nand U4163 (N_4163,N_3344,N_2685);
xor U4164 (N_4164,N_2167,N_3596);
or U4165 (N_4165,N_2778,N_3703);
or U4166 (N_4166,N_2428,N_2802);
and U4167 (N_4167,N_3686,N_2549);
nor U4168 (N_4168,N_3647,N_3591);
and U4169 (N_4169,N_2870,N_3529);
nand U4170 (N_4170,N_2846,N_3504);
or U4171 (N_4171,N_3443,N_3056);
nand U4172 (N_4172,N_3040,N_3565);
and U4173 (N_4173,N_3002,N_2748);
nand U4174 (N_4174,N_3481,N_3299);
nor U4175 (N_4175,N_3786,N_2978);
nand U4176 (N_4176,N_2690,N_2807);
nand U4177 (N_4177,N_2300,N_3486);
xnor U4178 (N_4178,N_3165,N_2333);
xnor U4179 (N_4179,N_3640,N_3313);
nor U4180 (N_4180,N_3601,N_2256);
and U4181 (N_4181,N_3863,N_2303);
nor U4182 (N_4182,N_3128,N_2446);
nand U4183 (N_4183,N_3386,N_3467);
and U4184 (N_4184,N_2602,N_3099);
nor U4185 (N_4185,N_3685,N_2561);
or U4186 (N_4186,N_2282,N_3178);
nand U4187 (N_4187,N_2003,N_3028);
nand U4188 (N_4188,N_3233,N_2743);
nor U4189 (N_4189,N_2983,N_2808);
and U4190 (N_4190,N_3763,N_3489);
or U4191 (N_4191,N_3407,N_2630);
nor U4192 (N_4192,N_2560,N_3153);
nor U4193 (N_4193,N_2660,N_2361);
or U4194 (N_4194,N_3275,N_3608);
nor U4195 (N_4195,N_3899,N_3523);
and U4196 (N_4196,N_3716,N_2388);
xor U4197 (N_4197,N_3885,N_3688);
nor U4198 (N_4198,N_3694,N_3524);
and U4199 (N_4199,N_2725,N_3627);
nor U4200 (N_4200,N_2861,N_3576);
nor U4201 (N_4201,N_2037,N_3854);
nor U4202 (N_4202,N_2662,N_2833);
xnor U4203 (N_4203,N_2057,N_3789);
nand U4204 (N_4204,N_3164,N_3537);
or U4205 (N_4205,N_3426,N_3205);
or U4206 (N_4206,N_3147,N_3825);
nand U4207 (N_4207,N_2832,N_2796);
or U4208 (N_4208,N_3438,N_2994);
and U4209 (N_4209,N_3681,N_2845);
nand U4210 (N_4210,N_2960,N_2197);
nor U4211 (N_4211,N_3955,N_2723);
nand U4212 (N_4212,N_2664,N_2922);
nor U4213 (N_4213,N_2415,N_2511);
nand U4214 (N_4214,N_2558,N_3360);
and U4215 (N_4215,N_3248,N_3328);
xnor U4216 (N_4216,N_2144,N_2402);
and U4217 (N_4217,N_3012,N_2372);
nor U4218 (N_4218,N_2815,N_2604);
or U4219 (N_4219,N_3280,N_2035);
xor U4220 (N_4220,N_2093,N_3645);
nor U4221 (N_4221,N_3962,N_3382);
nand U4222 (N_4222,N_3924,N_2521);
nand U4223 (N_4223,N_2698,N_3689);
and U4224 (N_4224,N_2492,N_2087);
and U4225 (N_4225,N_3195,N_2541);
xor U4226 (N_4226,N_2207,N_2526);
and U4227 (N_4227,N_2218,N_3330);
nor U4228 (N_4228,N_2487,N_2947);
and U4229 (N_4229,N_2566,N_3356);
nand U4230 (N_4230,N_2427,N_3879);
nand U4231 (N_4231,N_3149,N_2442);
nor U4232 (N_4232,N_3327,N_3518);
and U4233 (N_4233,N_3047,N_3587);
or U4234 (N_4234,N_3733,N_2757);
nand U4235 (N_4235,N_2412,N_3517);
or U4236 (N_4236,N_2576,N_2916);
or U4237 (N_4237,N_3355,N_3123);
nand U4238 (N_4238,N_3638,N_2206);
or U4239 (N_4239,N_2186,N_2745);
nand U4240 (N_4240,N_2444,N_2128);
nor U4241 (N_4241,N_2483,N_3181);
nand U4242 (N_4242,N_3204,N_3131);
nand U4243 (N_4243,N_3169,N_2971);
or U4244 (N_4244,N_2524,N_3919);
nor U4245 (N_4245,N_2434,N_3192);
and U4246 (N_4246,N_2520,N_2362);
nor U4247 (N_4247,N_3431,N_2678);
and U4248 (N_4248,N_2932,N_3208);
and U4249 (N_4249,N_2423,N_3500);
or U4250 (N_4250,N_2544,N_3942);
or U4251 (N_4251,N_3001,N_3495);
nor U4252 (N_4252,N_3559,N_3490);
and U4253 (N_4253,N_3350,N_3871);
and U4254 (N_4254,N_3232,N_2234);
nand U4255 (N_4255,N_2884,N_2824);
and U4256 (N_4256,N_3251,N_3187);
nor U4257 (N_4257,N_3578,N_3454);
nand U4258 (N_4258,N_2871,N_3094);
xnor U4259 (N_4259,N_3945,N_3018);
nor U4260 (N_4260,N_3062,N_2570);
nand U4261 (N_4261,N_2294,N_3338);
and U4262 (N_4262,N_2738,N_2370);
and U4263 (N_4263,N_3833,N_3704);
or U4264 (N_4264,N_3548,N_2495);
or U4265 (N_4265,N_2852,N_3791);
or U4266 (N_4266,N_2407,N_3911);
and U4267 (N_4267,N_3038,N_3433);
nor U4268 (N_4268,N_3656,N_3915);
nor U4269 (N_4269,N_2831,N_3475);
xnor U4270 (N_4270,N_2182,N_2989);
or U4271 (N_4271,N_2202,N_3963);
and U4272 (N_4272,N_3832,N_3134);
and U4273 (N_4273,N_3663,N_3819);
or U4274 (N_4274,N_3551,N_2095);
nand U4275 (N_4275,N_2145,N_3405);
nor U4276 (N_4276,N_3713,N_3041);
or U4277 (N_4277,N_3492,N_3996);
xor U4278 (N_4278,N_2283,N_3947);
and U4279 (N_4279,N_3235,N_3764);
nand U4280 (N_4280,N_3905,N_2006);
or U4281 (N_4281,N_2460,N_2746);
or U4282 (N_4282,N_3695,N_3760);
nand U4283 (N_4283,N_3346,N_2885);
and U4284 (N_4284,N_2419,N_3190);
or U4285 (N_4285,N_2043,N_3938);
and U4286 (N_4286,N_2002,N_2222);
nor U4287 (N_4287,N_2138,N_3802);
nor U4288 (N_4288,N_2911,N_3820);
and U4289 (N_4289,N_3215,N_2613);
nor U4290 (N_4290,N_3868,N_2346);
nor U4291 (N_4291,N_2368,N_2061);
and U4292 (N_4292,N_2121,N_2680);
and U4293 (N_4293,N_3497,N_2559);
or U4294 (N_4294,N_3505,N_3068);
or U4295 (N_4295,N_3166,N_3347);
xor U4296 (N_4296,N_3721,N_2455);
nor U4297 (N_4297,N_3132,N_2077);
nand U4298 (N_4298,N_3840,N_3263);
and U4299 (N_4299,N_2791,N_3117);
xor U4300 (N_4300,N_3420,N_2985);
nand U4301 (N_4301,N_3156,N_2142);
and U4302 (N_4302,N_2907,N_3010);
nand U4303 (N_4303,N_3471,N_2532);
xor U4304 (N_4304,N_3717,N_2711);
and U4305 (N_4305,N_2161,N_2886);
nor U4306 (N_4306,N_2274,N_3560);
xor U4307 (N_4307,N_2820,N_2776);
nand U4308 (N_4308,N_2395,N_3463);
xnor U4309 (N_4309,N_3246,N_3250);
and U4310 (N_4310,N_3990,N_2737);
or U4311 (N_4311,N_2707,N_3823);
xor U4312 (N_4312,N_3566,N_2988);
and U4313 (N_4313,N_2158,N_2608);
nor U4314 (N_4314,N_2198,N_2253);
nor U4315 (N_4315,N_2531,N_2410);
or U4316 (N_4316,N_2731,N_3557);
nand U4317 (N_4317,N_3288,N_3749);
nand U4318 (N_4318,N_2265,N_3242);
and U4319 (N_4319,N_2533,N_3484);
nand U4320 (N_4320,N_3508,N_2355);
and U4321 (N_4321,N_3933,N_3301);
nand U4322 (N_4322,N_3267,N_3558);
nor U4323 (N_4323,N_3639,N_3992);
and U4324 (N_4324,N_2934,N_3877);
or U4325 (N_4325,N_2045,N_2385);
nor U4326 (N_4326,N_2620,N_3554);
and U4327 (N_4327,N_3768,N_2117);
and U4328 (N_4328,N_2728,N_2227);
nor U4329 (N_4329,N_2851,N_3584);
or U4330 (N_4330,N_2216,N_2318);
nand U4331 (N_4331,N_2633,N_3783);
and U4332 (N_4332,N_3340,N_3222);
or U4333 (N_4333,N_3697,N_3439);
nor U4334 (N_4334,N_2443,N_2196);
nand U4335 (N_4335,N_2430,N_2471);
and U4336 (N_4336,N_2814,N_2545);
nor U4337 (N_4337,N_3918,N_2572);
and U4338 (N_4338,N_2400,N_2478);
nor U4339 (N_4339,N_2840,N_2465);
nand U4340 (N_4340,N_2519,N_2688);
nor U4341 (N_4341,N_2426,N_2441);
nor U4342 (N_4342,N_3814,N_3110);
or U4343 (N_4343,N_2114,N_2634);
nor U4344 (N_4344,N_3650,N_2987);
or U4345 (N_4345,N_3621,N_2159);
and U4346 (N_4346,N_2091,N_3553);
nor U4347 (N_4347,N_2979,N_3021);
nand U4348 (N_4348,N_2927,N_2191);
or U4349 (N_4349,N_3779,N_3541);
and U4350 (N_4350,N_2498,N_2853);
or U4351 (N_4351,N_2958,N_2675);
nand U4352 (N_4352,N_3295,N_3145);
nand U4353 (N_4353,N_2310,N_2281);
nor U4354 (N_4354,N_3901,N_2068);
xor U4355 (N_4355,N_2264,N_2736);
or U4356 (N_4356,N_2695,N_2786);
nand U4357 (N_4357,N_2838,N_3482);
and U4358 (N_4358,N_3462,N_3312);
and U4359 (N_4359,N_2066,N_3874);
or U4360 (N_4360,N_2575,N_2593);
nand U4361 (N_4361,N_2965,N_3743);
xor U4362 (N_4362,N_3296,N_2030);
nor U4363 (N_4363,N_3029,N_2311);
and U4364 (N_4364,N_2973,N_2293);
and U4365 (N_4365,N_2512,N_3329);
nand U4366 (N_4366,N_2875,N_3790);
and U4367 (N_4367,N_3236,N_3447);
nor U4368 (N_4368,N_3408,N_3369);
nand U4369 (N_4369,N_3415,N_3105);
nor U4370 (N_4370,N_2398,N_3226);
and U4371 (N_4371,N_2288,N_3636);
nor U4372 (N_4372,N_3458,N_2872);
nor U4373 (N_4373,N_3411,N_3723);
and U4374 (N_4374,N_2075,N_2330);
or U4375 (N_4375,N_2162,N_3079);
nor U4376 (N_4376,N_3897,N_2548);
and U4377 (N_4377,N_2518,N_2243);
and U4378 (N_4378,N_3512,N_3308);
nor U4379 (N_4379,N_2254,N_2708);
nor U4380 (N_4380,N_2431,N_2826);
or U4381 (N_4381,N_2081,N_3150);
nand U4382 (N_4382,N_3281,N_2363);
and U4383 (N_4383,N_3741,N_2750);
or U4384 (N_4384,N_2650,N_3424);
nor U4385 (N_4385,N_3483,N_2867);
or U4386 (N_4386,N_3305,N_3152);
and U4387 (N_4387,N_2307,N_3852);
xnor U4388 (N_4388,N_2233,N_2386);
nand U4389 (N_4389,N_2981,N_2273);
or U4390 (N_4390,N_2332,N_2567);
nor U4391 (N_4391,N_2139,N_2912);
and U4392 (N_4392,N_3754,N_3249);
nand U4393 (N_4393,N_2464,N_3585);
nor U4394 (N_4394,N_2247,N_3488);
nor U4395 (N_4395,N_3572,N_3025);
nor U4396 (N_4396,N_3244,N_3212);
nand U4397 (N_4397,N_3573,N_2691);
nand U4398 (N_4398,N_2212,N_2753);
or U4399 (N_4399,N_3264,N_3412);
nand U4400 (N_4400,N_2759,N_2092);
and U4401 (N_4401,N_2669,N_2543);
xor U4402 (N_4402,N_3856,N_2258);
nand U4403 (N_4403,N_2018,N_3130);
and U4404 (N_4404,N_2882,N_3750);
or U4405 (N_4405,N_2078,N_2823);
or U4406 (N_4406,N_2337,N_2228);
or U4407 (N_4407,N_2530,N_3635);
nor U4408 (N_4408,N_3014,N_2936);
nand U4409 (N_4409,N_2975,N_3580);
nand U4410 (N_4410,N_3964,N_3290);
or U4411 (N_4411,N_3227,N_2525);
nor U4412 (N_4412,N_3932,N_2706);
nor U4413 (N_4413,N_2705,N_2998);
nor U4414 (N_4414,N_3804,N_2624);
nor U4415 (N_4415,N_3395,N_2047);
nor U4416 (N_4416,N_2174,N_3377);
or U4417 (N_4417,N_2574,N_3196);
and U4418 (N_4418,N_3096,N_3262);
nor U4419 (N_4419,N_2210,N_2356);
nor U4420 (N_4420,N_2834,N_2890);
or U4421 (N_4421,N_2466,N_2881);
nand U4422 (N_4422,N_3668,N_2177);
nor U4423 (N_4423,N_3926,N_3766);
or U4424 (N_4424,N_3487,N_3409);
nor U4425 (N_4425,N_2754,N_2094);
and U4426 (N_4426,N_2056,N_2339);
nand U4427 (N_4427,N_2836,N_3997);
and U4428 (N_4428,N_2523,N_2752);
xor U4429 (N_4429,N_2260,N_2486);
nor U4430 (N_4430,N_2917,N_2830);
nor U4431 (N_4431,N_2086,N_3354);
nor U4432 (N_4432,N_2170,N_3142);
nor U4433 (N_4433,N_3398,N_3618);
and U4434 (N_4434,N_3671,N_3373);
nor U4435 (N_4435,N_2798,N_3525);
nand U4436 (N_4436,N_3646,N_2335);
and U4437 (N_4437,N_3731,N_3370);
nor U4438 (N_4438,N_3034,N_2557);
and U4439 (N_4439,N_2399,N_2255);
nor U4440 (N_4440,N_2719,N_3534);
or U4441 (N_4441,N_2119,N_2528);
nand U4442 (N_4442,N_3737,N_2485);
xor U4443 (N_4443,N_2209,N_2897);
nand U4444 (N_4444,N_2587,N_3074);
or U4445 (N_4445,N_2589,N_3844);
and U4446 (N_4446,N_3140,N_2403);
and U4447 (N_4447,N_2005,N_2166);
and U4448 (N_4448,N_2803,N_2173);
and U4449 (N_4449,N_3634,N_2480);
nand U4450 (N_4450,N_3320,N_3837);
nor U4451 (N_4451,N_3214,N_3035);
and U4452 (N_4452,N_3416,N_3782);
nand U4453 (N_4453,N_3276,N_2734);
or U4454 (N_4454,N_3461,N_3507);
or U4455 (N_4455,N_3088,N_3279);
xor U4456 (N_4456,N_3291,N_3974);
nand U4457 (N_4457,N_3999,N_3352);
nand U4458 (N_4458,N_3351,N_2610);
nor U4459 (N_4459,N_2581,N_3403);
nor U4460 (N_4460,N_3630,N_3000);
nand U4461 (N_4461,N_3624,N_2923);
xor U4462 (N_4462,N_2107,N_2321);
nor U4463 (N_4463,N_2941,N_3958);
nor U4464 (N_4464,N_2432,N_2098);
nor U4465 (N_4465,N_2467,N_2232);
nor U4466 (N_4466,N_3889,N_2324);
nor U4467 (N_4467,N_2059,N_2396);
and U4468 (N_4468,N_3528,N_2862);
nand U4469 (N_4469,N_2793,N_3851);
or U4470 (N_4470,N_3946,N_3049);
or U4471 (N_4471,N_3729,N_2889);
and U4472 (N_4472,N_3031,N_3391);
or U4473 (N_4473,N_2672,N_2779);
or U4474 (N_4474,N_3473,N_3530);
and U4475 (N_4475,N_2892,N_2108);
and U4476 (N_4476,N_2050,N_3219);
and U4477 (N_4477,N_3927,N_3256);
and U4478 (N_4478,N_3812,N_3503);
or U4479 (N_4479,N_2312,N_3959);
xnor U4480 (N_4480,N_2268,N_3803);
and U4481 (N_4481,N_2704,N_3849);
nand U4482 (N_4482,N_3599,N_2125);
and U4483 (N_4483,N_3995,N_3780);
nor U4484 (N_4484,N_3452,N_2149);
or U4485 (N_4485,N_3364,N_3326);
or U4486 (N_4486,N_3188,N_2764);
nor U4487 (N_4487,N_3315,N_3054);
or U4488 (N_4488,N_2221,N_3293);
nor U4489 (N_4489,N_2347,N_3255);
and U4490 (N_4490,N_2799,N_3981);
nand U4491 (N_4491,N_3864,N_2016);
and U4492 (N_4492,N_2280,N_3894);
nor U4493 (N_4493,N_3977,N_3895);
xnor U4494 (N_4494,N_2806,N_3422);
or U4495 (N_4495,N_3146,N_3292);
and U4496 (N_4496,N_2942,N_2088);
and U4497 (N_4497,N_2160,N_3343);
nor U4498 (N_4498,N_3476,N_2187);
nand U4499 (N_4499,N_3309,N_2429);
and U4500 (N_4500,N_3171,N_3637);
nor U4501 (N_4501,N_3268,N_3641);
nand U4502 (N_4502,N_2375,N_3390);
nand U4503 (N_4503,N_2349,N_3333);
nor U4504 (N_4504,N_3816,N_3739);
nor U4505 (N_4505,N_2489,N_2225);
nor U4506 (N_4506,N_3363,N_2011);
and U4507 (N_4507,N_3339,N_3531);
xor U4508 (N_4508,N_3817,N_3796);
and U4509 (N_4509,N_3818,N_3365);
nand U4510 (N_4510,N_2109,N_3834);
or U4511 (N_4511,N_2358,N_3020);
nand U4512 (N_4512,N_2720,N_3440);
nor U4513 (N_4513,N_3643,N_2418);
or U4514 (N_4514,N_3311,N_2132);
nand U4515 (N_4515,N_2854,N_3335);
nor U4516 (N_4516,N_3965,N_3869);
nand U4517 (N_4517,N_3254,N_2325);
or U4518 (N_4518,N_3116,N_3880);
nand U4519 (N_4519,N_3113,N_3542);
nor U4520 (N_4520,N_2631,N_3051);
nor U4521 (N_4521,N_3923,N_3097);
nor U4522 (N_4522,N_3751,N_3300);
and U4523 (N_4523,N_2063,N_3881);
nand U4524 (N_4524,N_2249,N_3180);
nor U4525 (N_4525,N_2367,N_3987);
or U4526 (N_4526,N_2123,N_3571);
and U4527 (N_4527,N_2328,N_2996);
or U4528 (N_4528,N_2900,N_3459);
and U4529 (N_4529,N_3914,N_2627);
nor U4530 (N_4530,N_3472,N_2878);
and U4531 (N_4531,N_2474,N_3951);
nand U4532 (N_4532,N_2046,N_3792);
nor U4533 (N_4533,N_2967,N_3535);
nand U4534 (N_4534,N_3907,N_2496);
and U4535 (N_4535,N_2951,N_3316);
and U4536 (N_4536,N_2115,N_3590);
or U4537 (N_4537,N_2924,N_2103);
nor U4538 (N_4538,N_2805,N_3286);
or U4539 (N_4539,N_3392,N_2986);
nand U4540 (N_4540,N_2208,N_2546);
xnor U4541 (N_4541,N_3740,N_2904);
nor U4542 (N_4542,N_3174,N_3042);
nand U4543 (N_4543,N_3189,N_3957);
nor U4544 (N_4544,N_2898,N_3839);
or U4545 (N_4545,N_3183,N_3513);
nor U4546 (N_4546,N_2762,N_3860);
and U4547 (N_4547,N_3728,N_3661);
nand U4548 (N_4548,N_3297,N_3167);
nand U4549 (N_4549,N_3075,N_2424);
nor U4550 (N_4550,N_3939,N_3708);
nand U4551 (N_4551,N_3579,N_2394);
and U4552 (N_4552,N_3148,N_2147);
nand U4553 (N_4553,N_3597,N_2850);
and U4554 (N_4554,N_2069,N_3136);
or U4555 (N_4555,N_3765,N_2868);
nor U4556 (N_4556,N_2582,N_3781);
and U4557 (N_4557,N_2065,N_3325);
or U4558 (N_4558,N_3337,N_3734);
nand U4559 (N_4559,N_3623,N_2767);
and U4560 (N_4560,N_2224,N_3649);
nand U4561 (N_4561,N_3653,N_3023);
nand U4562 (N_4562,N_3100,N_2211);
xnor U4563 (N_4563,N_3692,N_2891);
nand U4564 (N_4564,N_2893,N_3719);
and U4565 (N_4565,N_3949,N_2326);
or U4566 (N_4566,N_3788,N_3253);
xor U4567 (N_4567,N_2239,N_3985);
nor U4568 (N_4568,N_2291,N_3798);
nand U4569 (N_4569,N_3127,N_3662);
or U4570 (N_4570,N_2636,N_2730);
nand U4571 (N_4571,N_2997,N_3161);
nand U4572 (N_4572,N_2503,N_3726);
and U4573 (N_4573,N_2642,N_3892);
and U4574 (N_4574,N_2945,N_2040);
and U4575 (N_4575,N_3043,N_3934);
nand U4576 (N_4576,N_2259,N_3349);
nand U4577 (N_4577,N_3449,N_2376);
or U4578 (N_4578,N_2579,N_3522);
or U4579 (N_4579,N_2621,N_3626);
or U4580 (N_4580,N_2628,N_2064);
nor U4581 (N_4581,N_2645,N_3223);
or U4582 (N_4582,N_2411,N_3260);
and U4583 (N_4583,N_2928,N_2999);
and U4584 (N_4584,N_3432,N_2858);
nand U4585 (N_4585,N_3606,N_3696);
nor U4586 (N_4586,N_2679,N_3270);
and U4587 (N_4587,N_3824,N_3093);
nor U4588 (N_4588,N_2821,N_2716);
nor U4589 (N_4589,N_2113,N_3509);
or U4590 (N_4590,N_2449,N_3064);
nand U4591 (N_4591,N_2535,N_3550);
nand U4592 (N_4592,N_2564,N_3052);
and U4593 (N_4593,N_3715,N_2837);
nand U4594 (N_4594,N_3271,N_2199);
nor U4595 (N_4595,N_2849,N_2508);
and U4596 (N_4596,N_3397,N_2668);
nand U4597 (N_4597,N_2404,N_3577);
or U4598 (N_4598,N_3973,N_3514);
nand U4599 (N_4599,N_2131,N_3602);
nand U4600 (N_4600,N_2482,N_3314);
or U4601 (N_4601,N_2556,N_3053);
or U4602 (N_4602,N_2171,N_3417);
or U4603 (N_4603,N_2181,N_2354);
and U4604 (N_4604,N_2694,N_2034);
or U4605 (N_4605,N_3194,N_2215);
nand U4606 (N_4606,N_3888,N_3284);
or U4607 (N_4607,N_3218,N_2027);
xor U4608 (N_4608,N_3515,N_3137);
and U4609 (N_4609,N_3120,N_3058);
xnor U4610 (N_4610,N_3943,N_2800);
nor U4611 (N_4611,N_2481,N_2378);
nand U4612 (N_4612,N_3265,N_2336);
nand U4613 (N_4613,N_2970,N_3375);
nor U4614 (N_4614,N_2479,N_2933);
nand U4615 (N_4615,N_3988,N_2536);
and U4616 (N_4616,N_2472,N_3331);
xnor U4617 (N_4617,N_3491,N_3843);
nor U4618 (N_4618,N_2164,N_3184);
nor U4619 (N_4619,N_3778,N_3611);
nand U4620 (N_4620,N_2964,N_3091);
and U4621 (N_4621,N_3536,N_3283);
or U4622 (N_4622,N_3969,N_2070);
and U4623 (N_4623,N_2373,N_3855);
nor U4624 (N_4624,N_2379,N_3108);
and U4625 (N_4625,N_3294,N_3177);
nor U4626 (N_4626,N_2864,N_2217);
or U4627 (N_4627,N_3445,N_2277);
and U4628 (N_4628,N_3024,N_3561);
or U4629 (N_4629,N_3272,N_3759);
nand U4630 (N_4630,N_3617,N_2635);
or U4631 (N_4631,N_2732,N_2527);
or U4632 (N_4632,N_3613,N_3619);
and U4633 (N_4633,N_2248,N_3682);
and U4634 (N_4634,N_2580,N_3935);
or U4635 (N_4635,N_3077,N_2687);
nand U4636 (N_4636,N_3506,N_3499);
and U4637 (N_4637,N_2319,N_2550);
and U4638 (N_4638,N_3727,N_2974);
and U4639 (N_4639,N_3015,N_2020);
nand U4640 (N_4640,N_2152,N_2083);
nand U4641 (N_4641,N_3371,N_2659);
nand U4642 (N_4642,N_2775,N_3151);
nand U4643 (N_4643,N_2740,N_2920);
nand U4644 (N_4644,N_3450,N_3479);
or U4645 (N_4645,N_3418,N_2345);
or U4646 (N_4646,N_2322,N_2577);
nand U4647 (N_4647,N_3362,N_3037);
nand U4648 (N_4648,N_3468,N_3867);
or U4649 (N_4649,N_2497,N_3735);
or U4650 (N_4650,N_2118,N_3193);
or U4651 (N_4651,N_3827,N_2873);
or U4652 (N_4652,N_3890,N_3941);
and U4653 (N_4653,N_2306,N_3615);
and U4654 (N_4654,N_3808,N_2895);
xor U4655 (N_4655,N_2596,N_3230);
or U4656 (N_4656,N_2350,N_2957);
nor U4657 (N_4657,N_3252,N_2021);
xnor U4658 (N_4658,N_2359,N_2972);
and U4659 (N_4659,N_3210,N_2382);
nand U4660 (N_4660,N_3502,N_3785);
or U4661 (N_4661,N_2741,N_2652);
nand U4662 (N_4662,N_3221,N_2625);
and U4663 (N_4663,N_3806,N_2458);
and U4664 (N_4664,N_3972,N_2366);
or U4665 (N_4665,N_3975,N_2190);
nor U4666 (N_4666,N_2699,N_2484);
and U4667 (N_4667,N_3421,N_2169);
and U4668 (N_4668,N_2788,N_2747);
and U4669 (N_4669,N_2085,N_3126);
and U4670 (N_4670,N_2953,N_2529);
nor U4671 (N_4671,N_2205,N_2189);
xor U4672 (N_4672,N_2073,N_3143);
or U4673 (N_4673,N_2237,N_2506);
nor U4674 (N_4674,N_2155,N_2456);
and U4675 (N_4675,N_2136,N_2540);
or U4676 (N_4676,N_3071,N_2937);
and U4677 (N_4677,N_3359,N_3826);
nor U4678 (N_4678,N_3683,N_2269);
nor U4679 (N_4679,N_2039,N_3546);
and U4680 (N_4680,N_2859,N_3702);
or U4681 (N_4681,N_2049,N_2453);
nand U4682 (N_4682,N_2493,N_2991);
and U4683 (N_4683,N_3956,N_3800);
nand U4684 (N_4684,N_2856,N_2338);
nor U4685 (N_4685,N_3243,N_3368);
nand U4686 (N_4686,N_2784,N_2007);
and U4687 (N_4687,N_3614,N_3865);
nor U4688 (N_4688,N_2369,N_3274);
nor U4689 (N_4689,N_2146,N_3693);
or U4690 (N_4690,N_3900,N_2276);
nor U4691 (N_4691,N_3429,N_3902);
nand U4692 (N_4692,N_2984,N_3470);
nand U4693 (N_4693,N_2835,N_3592);
or U4694 (N_4694,N_2905,N_3632);
nor U4695 (N_4695,N_2150,N_2903);
or U4696 (N_4696,N_2074,N_3446);
nor U4697 (N_4697,N_2657,N_2129);
nand U4698 (N_4698,N_3875,N_3564);
xor U4699 (N_4699,N_2461,N_3318);
nand U4700 (N_4700,N_2044,N_2598);
nand U4701 (N_4701,N_3971,N_2435);
nand U4702 (N_4702,N_3680,N_3700);
or U4703 (N_4703,N_2888,N_3342);
xor U4704 (N_4704,N_3588,N_2313);
or U4705 (N_4705,N_2646,N_3644);
and U4706 (N_4706,N_3676,N_3207);
or U4707 (N_4707,N_2869,N_3872);
xor U4708 (N_4708,N_3144,N_2681);
nand U4709 (N_4709,N_3104,N_3176);
nand U4710 (N_4710,N_3547,N_2773);
nor U4711 (N_4711,N_3757,N_3944);
nand U4712 (N_4712,N_3086,N_2287);
or U4713 (N_4713,N_3410,N_2792);
nand U4714 (N_4714,N_2565,N_2841);
or U4715 (N_4715,N_3684,N_3083);
or U4716 (N_4716,N_3050,N_2516);
and U4717 (N_4717,N_3701,N_2204);
or U4718 (N_4718,N_2571,N_2076);
xnor U4719 (N_4719,N_2894,N_3921);
nor U4720 (N_4720,N_3991,N_3036);
or U4721 (N_4721,N_2818,N_2316);
or U4722 (N_4722,N_3157,N_3642);
nand U4723 (N_4723,N_3348,N_2185);
and U4724 (N_4724,N_2876,N_2352);
nand U4725 (N_4725,N_2299,N_2944);
nand U4726 (N_4726,N_3444,N_2573);
nand U4727 (N_4727,N_3770,N_3427);
xor U4728 (N_4728,N_3511,N_3870);
or U4729 (N_4729,N_3321,N_2651);
xor U4730 (N_4730,N_3659,N_3385);
nor U4731 (N_4731,N_3809,N_3570);
xnor U4732 (N_4732,N_3989,N_3287);
nor U4733 (N_4733,N_3655,N_3383);
or U4734 (N_4734,N_3206,N_3076);
nand U4735 (N_4735,N_3775,N_3030);
or U4736 (N_4736,N_3485,N_2879);
nand U4737 (N_4737,N_2275,N_2272);
or U4738 (N_4738,N_3670,N_3229);
and U4739 (N_4739,N_2451,N_2143);
nor U4740 (N_4740,N_3761,N_2607);
or U4741 (N_4741,N_2626,N_3435);
or U4742 (N_4742,N_2462,N_3341);
and U4743 (N_4743,N_3784,N_2914);
and U4744 (N_4744,N_2188,N_2156);
or U4745 (N_4745,N_3983,N_2605);
or U4746 (N_4746,N_3762,N_2250);
and U4747 (N_4747,N_2896,N_3170);
xnor U4748 (N_4748,N_3691,N_2939);
or U4749 (N_4749,N_3811,N_2758);
nor U4750 (N_4750,N_2165,N_3866);
or U4751 (N_4751,N_3209,N_2447);
and U4752 (N_4752,N_3742,N_3197);
xnor U4753 (N_4753,N_3125,N_3323);
and U4754 (N_4754,N_3376,N_2553);
nand U4755 (N_4755,N_2600,N_3245);
and U4756 (N_4756,N_3712,N_2440);
or U4757 (N_4757,N_3724,N_3898);
and U4758 (N_4758,N_3567,N_2844);
nor U4759 (N_4759,N_2298,N_3154);
nand U4760 (N_4760,N_3203,N_3202);
and U4761 (N_4761,N_3893,N_3211);
nor U4762 (N_4762,N_2591,N_2012);
nor U4763 (N_4763,N_3748,N_2140);
and U4764 (N_4764,N_3231,N_2586);
or U4765 (N_4765,N_2777,N_3044);
nor U4766 (N_4766,N_2389,N_2684);
nand U4767 (N_4767,N_3556,N_3118);
nor U4768 (N_4768,N_2771,N_2331);
xor U4769 (N_4769,N_3631,N_3593);
and U4770 (N_4770,N_2238,N_3519);
xnor U4771 (N_4771,N_3771,N_2735);
or U4772 (N_4772,N_2656,N_2112);
nor U4773 (N_4773,N_2542,N_3007);
nor U4774 (N_4774,N_2925,N_3882);
or U4775 (N_4775,N_3747,N_2629);
and U4776 (N_4776,N_2822,N_3594);
nor U4777 (N_4777,N_2883,N_3625);
xor U4778 (N_4778,N_2595,N_2053);
nor U4779 (N_4779,N_2568,N_3850);
or U4780 (N_4780,N_3846,N_2405);
nor U4781 (N_4781,N_2819,N_3121);
nor U4782 (N_4782,N_2811,N_2847);
nand U4783 (N_4783,N_3612,N_3073);
and U4784 (N_4784,N_2670,N_2855);
or U4785 (N_4785,N_2284,N_2416);
nand U4786 (N_4786,N_3772,N_2425);
and U4787 (N_4787,N_2315,N_2787);
or U4788 (N_4788,N_3690,N_3912);
nor U4789 (N_4789,N_2097,N_2433);
nor U4790 (N_4790,N_2051,N_3008);
xor U4791 (N_4791,N_3769,N_2501);
or U4792 (N_4792,N_3842,N_2842);
nand U4793 (N_4793,N_2940,N_3278);
or U4794 (N_4794,N_3822,N_3428);
nand U4795 (N_4795,N_3345,N_2054);
nor U4796 (N_4796,N_3909,N_3419);
or U4797 (N_4797,N_2374,N_3238);
and U4798 (N_4798,N_2153,N_2009);
nor U4799 (N_4799,N_2214,N_2179);
nor U4800 (N_4800,N_3648,N_3493);
or U4801 (N_4801,N_3610,N_2488);
nor U4802 (N_4802,N_3756,N_3451);
nand U4803 (N_4803,N_3516,N_2713);
and U4804 (N_4804,N_2601,N_2089);
nor U4805 (N_4805,N_3658,N_2193);
or U4806 (N_4806,N_2448,N_3533);
or U4807 (N_4807,N_2365,N_3952);
nand U4808 (N_4808,N_3334,N_3474);
or U4809 (N_4809,N_3045,N_2096);
nand U4810 (N_4810,N_3583,N_2751);
nand U4811 (N_4811,N_2163,N_2203);
nand U4812 (N_4812,N_2671,N_2151);
nand U4813 (N_4813,N_2644,N_3119);
or U4814 (N_4814,N_2910,N_2327);
nor U4815 (N_4815,N_2594,N_2742);
xnor U4816 (N_4816,N_3857,N_2590);
nand U4817 (N_4817,N_2401,N_3698);
xor U4818 (N_4818,N_2262,N_2267);
xnor U4819 (N_4819,N_3057,N_2683);
nand U4820 (N_4820,N_3237,N_2084);
nor U4821 (N_4821,N_3936,N_2279);
or U4822 (N_4822,N_3437,N_2008);
nor U4823 (N_4823,N_2877,N_2555);
nand U4824 (N_4824,N_3848,N_2825);
and U4825 (N_4825,N_2952,N_2454);
xor U4826 (N_4826,N_2614,N_3017);
and U4827 (N_4827,N_3664,N_2290);
nor U4828 (N_4828,N_3061,N_3595);
nor U4829 (N_4829,N_2052,N_2192);
or U4830 (N_4830,N_2622,N_2682);
nand U4831 (N_4831,N_2915,N_3660);
or U4832 (N_4832,N_2901,N_2612);
nor U4833 (N_4833,N_3059,N_2038);
or U4834 (N_4834,N_2921,N_3448);
or U4835 (N_4835,N_2763,N_2099);
nor U4836 (N_4836,N_3813,N_3168);
and U4837 (N_4837,N_3465,N_2133);
or U4838 (N_4838,N_3986,N_3162);
xor U4839 (N_4839,N_3106,N_3285);
nand U4840 (N_4840,N_2459,N_3241);
and U4841 (N_4841,N_2663,N_3111);
nor U4842 (N_4842,N_2033,N_3767);
nand U4843 (N_4843,N_2017,N_3776);
and U4844 (N_4844,N_3752,N_2666);
nand U4845 (N_4845,N_2334,N_3112);
or U4846 (N_4846,N_3616,N_3374);
or U4847 (N_4847,N_2913,N_3586);
or U4848 (N_4848,N_3501,N_3821);
and U4849 (N_4849,N_2242,N_2959);
and U4850 (N_4850,N_2195,N_2926);
and U4851 (N_4851,N_3455,N_2804);
or U4852 (N_4852,N_3948,N_3033);
nor U4853 (N_4853,N_2286,N_3003);
or U4854 (N_4854,N_2880,N_3967);
or U4855 (N_4855,N_2774,N_2789);
nand U4856 (N_4856,N_2230,N_3829);
and U4857 (N_4857,N_3442,N_2863);
nand U4858 (N_4858,N_3372,N_2739);
or U4859 (N_4859,N_2829,N_2420);
nor U4860 (N_4860,N_3200,N_2421);
nor U4861 (N_4861,N_2296,N_3836);
xor U4862 (N_4862,N_3133,N_2000);
or U4863 (N_4863,N_3414,N_2135);
or U4864 (N_4864,N_3213,N_2026);
and U4865 (N_4865,N_2848,N_2623);
nor U4866 (N_4866,N_2785,N_3604);
xor U4867 (N_4867,N_3540,N_2562);
nand U4868 (N_4868,N_3917,N_3725);
nand U4869 (N_4869,N_2475,N_2689);
and U4870 (N_4870,N_3745,N_3520);
nor U4871 (N_4871,N_2673,N_3155);
and U4872 (N_4872,N_2110,N_3081);
xnor U4873 (N_4873,N_3521,N_3859);
nor U4874 (N_4874,N_2371,N_3277);
nor U4875 (N_4875,N_2079,N_3976);
nand U4876 (N_4876,N_3982,N_2724);
or U4877 (N_4877,N_2578,N_2148);
and U4878 (N_4878,N_2761,N_3009);
nand U4879 (N_4879,N_3887,N_3699);
and U4880 (N_4880,N_2391,N_3201);
xor U4881 (N_4881,N_3805,N_2102);
nand U4882 (N_4882,N_2105,N_3925);
and U4883 (N_4883,N_3498,N_2041);
nand U4884 (N_4884,N_2477,N_2058);
xor U4885 (N_4885,N_3080,N_2797);
or U4886 (N_4886,N_3883,N_3247);
and U4887 (N_4887,N_3466,N_3469);
nor U4888 (N_4888,N_2473,N_3878);
and U4889 (N_4889,N_2504,N_2537);
nor U4890 (N_4890,N_2584,N_2154);
or U4891 (N_4891,N_3937,N_3913);
nor U4892 (N_4892,N_2956,N_2514);
and U4893 (N_4893,N_3046,N_3667);
xor U4894 (N_4894,N_3575,N_3388);
nor U4895 (N_4895,N_3179,N_2665);
or U4896 (N_4896,N_3744,N_3379);
nor U4897 (N_4897,N_3581,N_2760);
and U4898 (N_4898,N_2827,N_2308);
nor U4899 (N_4899,N_3807,N_2071);
nor U4900 (N_4900,N_3332,N_2765);
xnor U4901 (N_4901,N_3678,N_3102);
and U4902 (N_4902,N_2812,N_2606);
and U4903 (N_4903,N_3457,N_2062);
nor U4904 (N_4904,N_2413,N_3732);
xor U4905 (N_4905,N_2509,N_3622);
or U4906 (N_4906,N_3545,N_2130);
or U4907 (N_4907,N_3773,N_3672);
and U4908 (N_4908,N_3787,N_3810);
nand U4909 (N_4909,N_2507,N_3361);
nor U4910 (N_4910,N_2463,N_2770);
and U4911 (N_4911,N_2585,N_3931);
nand U4912 (N_4912,N_3257,N_2918);
xnor U4913 (N_4913,N_2909,N_2494);
and U4914 (N_4914,N_2323,N_3978);
nand U4915 (N_4915,N_2241,N_3984);
nor U4916 (N_4916,N_2439,N_3953);
or U4917 (N_4917,N_2090,N_3101);
nor U4918 (N_4918,N_3801,N_2899);
xnor U4919 (N_4919,N_2263,N_2810);
nor U4920 (N_4920,N_3555,N_3950);
nand U4921 (N_4921,N_2025,N_3998);
nor U4922 (N_4922,N_2360,N_3401);
nor U4923 (N_4923,N_3107,N_2067);
or U4924 (N_4924,N_2029,N_3317);
or U4925 (N_4925,N_2522,N_3027);
or U4926 (N_4926,N_2236,N_3400);
and U4927 (N_4927,N_3173,N_3753);
and U4928 (N_4928,N_2615,N_3620);
and U4929 (N_4929,N_3908,N_3135);
nor U4930 (N_4930,N_2261,N_2104);
and U4931 (N_4931,N_2701,N_3261);
and U4932 (N_4932,N_3815,N_2783);
nor U4933 (N_4933,N_2980,N_2611);
or U4934 (N_4934,N_3980,N_3302);
nor U4935 (N_4935,N_3795,N_2168);
nor U4936 (N_4936,N_3598,N_2697);
and U4937 (N_4937,N_3240,N_3022);
and U4938 (N_4938,N_2616,N_3182);
and U4939 (N_4939,N_3109,N_3954);
nor U4940 (N_4940,N_3526,N_2175);
nor U4941 (N_4941,N_2289,N_2865);
or U4942 (N_4942,N_2414,N_2655);
xnor U4943 (N_4943,N_2667,N_3574);
and U4944 (N_4944,N_3234,N_2693);
nor U4945 (N_4945,N_3838,N_3628);
and U4946 (N_4946,N_2968,N_2004);
xnor U4947 (N_4947,N_2661,N_2599);
nor U4948 (N_4948,N_3198,N_2353);
or U4949 (N_4949,N_2603,N_2755);
or U4950 (N_4950,N_3396,N_2592);
nand U4951 (N_4951,N_3994,N_2408);
nor U4952 (N_4952,N_2930,N_2387);
nand U4953 (N_4953,N_3722,N_2397);
and U4954 (N_4954,N_3453,N_2231);
or U4955 (N_4955,N_2860,N_2122);
nor U4956 (N_4956,N_2931,N_2715);
nor U4957 (N_4957,N_2436,N_3067);
and U4958 (N_4958,N_3922,N_2962);
nor U4959 (N_4959,N_2010,N_3158);
nand U4960 (N_4960,N_3746,N_3920);
or U4961 (N_4961,N_3562,N_3394);
and U4962 (N_4962,N_2781,N_2445);
nand U4963 (N_4963,N_2351,N_2619);
xor U4964 (N_4964,N_2505,N_2383);
nor U4965 (N_4965,N_3122,N_2995);
xor U4966 (N_4966,N_3084,N_3063);
nand U4967 (N_4967,N_2700,N_3026);
nor U4968 (N_4968,N_3532,N_3916);
nand U4969 (N_4969,N_2515,N_2381);
or U4970 (N_4970,N_3930,N_3904);
and U4971 (N_4971,N_3367,N_3006);
or U4972 (N_4972,N_3282,N_3055);
or U4973 (N_4973,N_2513,N_3873);
xor U4974 (N_4974,N_2219,N_2768);
and U4975 (N_4975,N_2229,N_2906);
or U4976 (N_4976,N_3159,N_3718);
nor U4977 (N_4977,N_2048,N_3185);
nand U4978 (N_4978,N_3070,N_3456);
nor U4979 (N_4979,N_2714,N_3199);
xnor U4980 (N_4980,N_3605,N_2676);
nand U4981 (N_4981,N_2641,N_3413);
nor U4982 (N_4982,N_3381,N_2632);
and U4983 (N_4983,N_2703,N_3687);
and U4984 (N_4984,N_3304,N_2200);
and U4985 (N_4985,N_2637,N_3092);
and U4986 (N_4986,N_2499,N_2357);
nand U4987 (N_4987,N_3884,N_2790);
or U4988 (N_4988,N_2500,N_2297);
nor U4989 (N_4989,N_3319,N_3228);
xnor U4990 (N_4990,N_2772,N_2828);
or U4991 (N_4991,N_3794,N_2552);
xnor U4992 (N_4992,N_2223,N_3072);
nand U4993 (N_4993,N_3674,N_2654);
nor U4994 (N_4994,N_3082,N_2721);
nand U4995 (N_4995,N_3399,N_3460);
and U4996 (N_4996,N_2780,N_2653);
or U4997 (N_4997,N_3845,N_2857);
nor U4998 (N_4998,N_2677,N_2015);
xor U4999 (N_4999,N_2120,N_3090);
xor U5000 (N_5000,N_2468,N_3366);
nor U5001 (N_5001,N_2071,N_2513);
and U5002 (N_5002,N_3556,N_3422);
nor U5003 (N_5003,N_2356,N_2451);
xnor U5004 (N_5004,N_3833,N_3075);
nand U5005 (N_5005,N_3162,N_2539);
nor U5006 (N_5006,N_3001,N_3874);
or U5007 (N_5007,N_3026,N_2162);
nor U5008 (N_5008,N_2285,N_2798);
nand U5009 (N_5009,N_3942,N_3581);
nand U5010 (N_5010,N_3795,N_3955);
xnor U5011 (N_5011,N_3204,N_3452);
and U5012 (N_5012,N_3186,N_2960);
and U5013 (N_5013,N_2511,N_3534);
nand U5014 (N_5014,N_2353,N_2406);
and U5015 (N_5015,N_3502,N_2363);
nand U5016 (N_5016,N_3817,N_3195);
nor U5017 (N_5017,N_3895,N_2922);
or U5018 (N_5018,N_2649,N_3138);
or U5019 (N_5019,N_2901,N_3724);
and U5020 (N_5020,N_3522,N_2903);
xor U5021 (N_5021,N_3060,N_2861);
and U5022 (N_5022,N_2468,N_3553);
nand U5023 (N_5023,N_3643,N_3391);
xnor U5024 (N_5024,N_2569,N_3744);
nand U5025 (N_5025,N_2801,N_2253);
nor U5026 (N_5026,N_2028,N_2385);
or U5027 (N_5027,N_3594,N_3252);
nor U5028 (N_5028,N_2022,N_2239);
nor U5029 (N_5029,N_3056,N_3360);
nand U5030 (N_5030,N_2191,N_3360);
nor U5031 (N_5031,N_2150,N_2392);
or U5032 (N_5032,N_3936,N_3368);
or U5033 (N_5033,N_2202,N_3126);
nand U5034 (N_5034,N_2802,N_3774);
xnor U5035 (N_5035,N_2768,N_3408);
nor U5036 (N_5036,N_3673,N_2963);
and U5037 (N_5037,N_3895,N_2134);
nor U5038 (N_5038,N_3483,N_3602);
nor U5039 (N_5039,N_2828,N_3144);
nand U5040 (N_5040,N_2189,N_3721);
xnor U5041 (N_5041,N_3481,N_3242);
nor U5042 (N_5042,N_3629,N_2429);
or U5043 (N_5043,N_3513,N_3036);
nor U5044 (N_5044,N_3844,N_3781);
or U5045 (N_5045,N_2387,N_2655);
and U5046 (N_5046,N_3361,N_3341);
nor U5047 (N_5047,N_3080,N_2975);
nand U5048 (N_5048,N_2824,N_2216);
or U5049 (N_5049,N_3200,N_2771);
nand U5050 (N_5050,N_3018,N_2215);
xnor U5051 (N_5051,N_3201,N_2494);
nand U5052 (N_5052,N_3480,N_3311);
nor U5053 (N_5053,N_2529,N_2681);
xor U5054 (N_5054,N_3344,N_3016);
nand U5055 (N_5055,N_2445,N_3722);
nor U5056 (N_5056,N_3150,N_2947);
or U5057 (N_5057,N_3810,N_2370);
or U5058 (N_5058,N_3719,N_3455);
nor U5059 (N_5059,N_3714,N_2539);
nor U5060 (N_5060,N_3929,N_2437);
nor U5061 (N_5061,N_2537,N_2299);
nor U5062 (N_5062,N_2399,N_3114);
and U5063 (N_5063,N_2946,N_3331);
nor U5064 (N_5064,N_2106,N_2266);
or U5065 (N_5065,N_3917,N_2196);
nor U5066 (N_5066,N_3731,N_3683);
or U5067 (N_5067,N_3722,N_3875);
and U5068 (N_5068,N_3370,N_2269);
nor U5069 (N_5069,N_3835,N_3953);
and U5070 (N_5070,N_2391,N_3763);
and U5071 (N_5071,N_2738,N_2740);
and U5072 (N_5072,N_2457,N_3495);
and U5073 (N_5073,N_2547,N_2911);
and U5074 (N_5074,N_2374,N_3962);
and U5075 (N_5075,N_3308,N_3263);
nor U5076 (N_5076,N_2569,N_3400);
nand U5077 (N_5077,N_2148,N_3210);
nor U5078 (N_5078,N_2030,N_3989);
and U5079 (N_5079,N_2380,N_2070);
nor U5080 (N_5080,N_3107,N_2469);
and U5081 (N_5081,N_2279,N_3957);
and U5082 (N_5082,N_2317,N_3474);
nand U5083 (N_5083,N_3982,N_2388);
or U5084 (N_5084,N_3061,N_3309);
nand U5085 (N_5085,N_2955,N_3306);
and U5086 (N_5086,N_3780,N_3189);
xor U5087 (N_5087,N_2439,N_3938);
nand U5088 (N_5088,N_3063,N_3882);
or U5089 (N_5089,N_3302,N_2803);
and U5090 (N_5090,N_2040,N_3558);
and U5091 (N_5091,N_2726,N_3917);
and U5092 (N_5092,N_3101,N_3756);
and U5093 (N_5093,N_3555,N_2747);
and U5094 (N_5094,N_3863,N_3651);
nor U5095 (N_5095,N_2804,N_3690);
nor U5096 (N_5096,N_2466,N_3674);
nand U5097 (N_5097,N_3706,N_3544);
nor U5098 (N_5098,N_3556,N_2223);
or U5099 (N_5099,N_3806,N_2954);
and U5100 (N_5100,N_3317,N_3222);
nor U5101 (N_5101,N_3617,N_3562);
and U5102 (N_5102,N_2068,N_2792);
or U5103 (N_5103,N_3244,N_2017);
or U5104 (N_5104,N_2008,N_3758);
nand U5105 (N_5105,N_2170,N_3485);
and U5106 (N_5106,N_2266,N_3133);
or U5107 (N_5107,N_2236,N_2539);
nand U5108 (N_5108,N_3695,N_3045);
xor U5109 (N_5109,N_3070,N_3191);
or U5110 (N_5110,N_2240,N_2377);
xnor U5111 (N_5111,N_2559,N_3905);
nand U5112 (N_5112,N_3788,N_3573);
and U5113 (N_5113,N_3870,N_2892);
and U5114 (N_5114,N_3355,N_3958);
nand U5115 (N_5115,N_3025,N_3823);
nand U5116 (N_5116,N_2915,N_2312);
xnor U5117 (N_5117,N_2851,N_3286);
nor U5118 (N_5118,N_2010,N_3346);
nor U5119 (N_5119,N_2833,N_2731);
and U5120 (N_5120,N_3283,N_3600);
nand U5121 (N_5121,N_2623,N_2657);
or U5122 (N_5122,N_3183,N_2623);
nor U5123 (N_5123,N_2524,N_3665);
nor U5124 (N_5124,N_2479,N_2627);
nor U5125 (N_5125,N_2345,N_2412);
and U5126 (N_5126,N_3973,N_3652);
and U5127 (N_5127,N_2500,N_3502);
nand U5128 (N_5128,N_3510,N_2754);
nand U5129 (N_5129,N_2517,N_3127);
nand U5130 (N_5130,N_3340,N_2812);
or U5131 (N_5131,N_2145,N_2587);
xor U5132 (N_5132,N_2294,N_2597);
and U5133 (N_5133,N_2034,N_3426);
nand U5134 (N_5134,N_2938,N_2324);
xnor U5135 (N_5135,N_3912,N_2702);
nor U5136 (N_5136,N_2841,N_3487);
nand U5137 (N_5137,N_2640,N_2408);
or U5138 (N_5138,N_2025,N_2914);
and U5139 (N_5139,N_2901,N_2979);
xnor U5140 (N_5140,N_3776,N_3698);
xor U5141 (N_5141,N_2404,N_3430);
nand U5142 (N_5142,N_3546,N_3061);
nand U5143 (N_5143,N_3480,N_3539);
nor U5144 (N_5144,N_2852,N_3348);
and U5145 (N_5145,N_3114,N_3073);
nand U5146 (N_5146,N_3111,N_2552);
or U5147 (N_5147,N_3321,N_2336);
nor U5148 (N_5148,N_2436,N_2279);
nand U5149 (N_5149,N_3680,N_2840);
and U5150 (N_5150,N_3966,N_3618);
nor U5151 (N_5151,N_2796,N_3134);
nand U5152 (N_5152,N_2444,N_3240);
xnor U5153 (N_5153,N_2757,N_3216);
or U5154 (N_5154,N_2043,N_2118);
nor U5155 (N_5155,N_3513,N_3976);
nand U5156 (N_5156,N_3791,N_3602);
and U5157 (N_5157,N_2016,N_2785);
or U5158 (N_5158,N_2417,N_3145);
nor U5159 (N_5159,N_3191,N_2132);
or U5160 (N_5160,N_2319,N_3604);
or U5161 (N_5161,N_2737,N_2901);
or U5162 (N_5162,N_3576,N_3596);
and U5163 (N_5163,N_3017,N_3879);
nor U5164 (N_5164,N_3782,N_3916);
or U5165 (N_5165,N_2214,N_2980);
nor U5166 (N_5166,N_3592,N_2732);
or U5167 (N_5167,N_3789,N_2122);
and U5168 (N_5168,N_2767,N_3307);
nand U5169 (N_5169,N_3161,N_2111);
nor U5170 (N_5170,N_3995,N_2738);
and U5171 (N_5171,N_3815,N_2334);
and U5172 (N_5172,N_3025,N_3376);
or U5173 (N_5173,N_2315,N_2463);
or U5174 (N_5174,N_2832,N_2035);
nor U5175 (N_5175,N_3075,N_3561);
nor U5176 (N_5176,N_2165,N_3499);
or U5177 (N_5177,N_2282,N_2197);
nand U5178 (N_5178,N_3356,N_3456);
nand U5179 (N_5179,N_2140,N_3841);
nor U5180 (N_5180,N_3907,N_2592);
nor U5181 (N_5181,N_2943,N_2114);
nor U5182 (N_5182,N_2356,N_2103);
and U5183 (N_5183,N_2660,N_3795);
nand U5184 (N_5184,N_2539,N_2642);
or U5185 (N_5185,N_2919,N_2332);
nand U5186 (N_5186,N_3400,N_3203);
xor U5187 (N_5187,N_3688,N_3508);
nor U5188 (N_5188,N_3815,N_3125);
and U5189 (N_5189,N_2392,N_3346);
nand U5190 (N_5190,N_3680,N_3236);
and U5191 (N_5191,N_3689,N_2699);
nand U5192 (N_5192,N_3155,N_2701);
nand U5193 (N_5193,N_2651,N_3987);
xnor U5194 (N_5194,N_2641,N_2225);
and U5195 (N_5195,N_3926,N_3196);
nand U5196 (N_5196,N_2102,N_3114);
xnor U5197 (N_5197,N_2992,N_2381);
xor U5198 (N_5198,N_3223,N_2808);
nand U5199 (N_5199,N_2020,N_3807);
nand U5200 (N_5200,N_3545,N_3047);
or U5201 (N_5201,N_3712,N_2559);
and U5202 (N_5202,N_2941,N_3661);
and U5203 (N_5203,N_2174,N_2263);
and U5204 (N_5204,N_2592,N_2003);
nand U5205 (N_5205,N_3601,N_3396);
xor U5206 (N_5206,N_2500,N_2177);
nor U5207 (N_5207,N_2604,N_2837);
nand U5208 (N_5208,N_3242,N_2433);
nand U5209 (N_5209,N_2002,N_3658);
nand U5210 (N_5210,N_3134,N_3541);
nand U5211 (N_5211,N_3182,N_2697);
nor U5212 (N_5212,N_3025,N_3611);
and U5213 (N_5213,N_3305,N_3236);
and U5214 (N_5214,N_3712,N_3156);
or U5215 (N_5215,N_2070,N_3214);
xnor U5216 (N_5216,N_3666,N_3144);
and U5217 (N_5217,N_3365,N_2346);
xor U5218 (N_5218,N_3861,N_3174);
and U5219 (N_5219,N_2797,N_3217);
nor U5220 (N_5220,N_2699,N_3035);
nand U5221 (N_5221,N_3688,N_3004);
nand U5222 (N_5222,N_2862,N_2292);
and U5223 (N_5223,N_3170,N_2638);
nand U5224 (N_5224,N_3980,N_2338);
nand U5225 (N_5225,N_3344,N_2468);
and U5226 (N_5226,N_3568,N_2810);
nor U5227 (N_5227,N_2163,N_2741);
nand U5228 (N_5228,N_3033,N_3262);
nand U5229 (N_5229,N_2992,N_2964);
or U5230 (N_5230,N_2846,N_3849);
and U5231 (N_5231,N_3779,N_3653);
or U5232 (N_5232,N_2191,N_2623);
or U5233 (N_5233,N_2515,N_3647);
xor U5234 (N_5234,N_2449,N_2613);
xor U5235 (N_5235,N_3149,N_3406);
or U5236 (N_5236,N_2727,N_2751);
nand U5237 (N_5237,N_3592,N_3409);
and U5238 (N_5238,N_2229,N_3633);
nor U5239 (N_5239,N_3564,N_3871);
or U5240 (N_5240,N_2579,N_2994);
nor U5241 (N_5241,N_3578,N_3030);
nor U5242 (N_5242,N_2089,N_2494);
nor U5243 (N_5243,N_3771,N_2739);
and U5244 (N_5244,N_3862,N_2894);
nand U5245 (N_5245,N_2721,N_2463);
and U5246 (N_5246,N_2512,N_2936);
nand U5247 (N_5247,N_3309,N_3128);
or U5248 (N_5248,N_2148,N_3408);
and U5249 (N_5249,N_3627,N_2836);
or U5250 (N_5250,N_2638,N_3080);
xor U5251 (N_5251,N_3363,N_2164);
nor U5252 (N_5252,N_3808,N_3576);
nand U5253 (N_5253,N_3766,N_3273);
or U5254 (N_5254,N_2054,N_2351);
nand U5255 (N_5255,N_3537,N_3839);
nor U5256 (N_5256,N_3191,N_2514);
nor U5257 (N_5257,N_3086,N_3381);
xnor U5258 (N_5258,N_3104,N_3771);
nor U5259 (N_5259,N_2642,N_2989);
and U5260 (N_5260,N_2538,N_2949);
xor U5261 (N_5261,N_2835,N_2522);
nand U5262 (N_5262,N_2441,N_3835);
nand U5263 (N_5263,N_3001,N_2972);
or U5264 (N_5264,N_3651,N_3887);
and U5265 (N_5265,N_2804,N_3489);
and U5266 (N_5266,N_3307,N_2366);
or U5267 (N_5267,N_3910,N_2581);
nor U5268 (N_5268,N_2244,N_3964);
or U5269 (N_5269,N_3236,N_3287);
nand U5270 (N_5270,N_3326,N_2318);
nand U5271 (N_5271,N_2368,N_3843);
nand U5272 (N_5272,N_2749,N_2625);
and U5273 (N_5273,N_2641,N_3907);
or U5274 (N_5274,N_3665,N_3714);
xor U5275 (N_5275,N_3135,N_3847);
nand U5276 (N_5276,N_3766,N_2767);
xor U5277 (N_5277,N_3731,N_2057);
or U5278 (N_5278,N_2771,N_2985);
nand U5279 (N_5279,N_2975,N_3197);
and U5280 (N_5280,N_2610,N_3318);
xor U5281 (N_5281,N_3927,N_2278);
or U5282 (N_5282,N_2744,N_2105);
and U5283 (N_5283,N_3800,N_3588);
and U5284 (N_5284,N_3576,N_3372);
nor U5285 (N_5285,N_3804,N_3124);
and U5286 (N_5286,N_2061,N_2245);
and U5287 (N_5287,N_3602,N_3226);
or U5288 (N_5288,N_3299,N_2837);
or U5289 (N_5289,N_2375,N_2387);
nand U5290 (N_5290,N_2326,N_3355);
and U5291 (N_5291,N_2506,N_2508);
and U5292 (N_5292,N_2819,N_2900);
or U5293 (N_5293,N_3261,N_3084);
and U5294 (N_5294,N_3675,N_2085);
nor U5295 (N_5295,N_3571,N_3960);
nand U5296 (N_5296,N_2247,N_3592);
nand U5297 (N_5297,N_2662,N_2116);
nor U5298 (N_5298,N_3709,N_3390);
xor U5299 (N_5299,N_2570,N_2796);
nor U5300 (N_5300,N_3979,N_2105);
xnor U5301 (N_5301,N_3435,N_3505);
xnor U5302 (N_5302,N_2172,N_2476);
or U5303 (N_5303,N_3547,N_3108);
xnor U5304 (N_5304,N_3899,N_3806);
nor U5305 (N_5305,N_2811,N_3146);
nor U5306 (N_5306,N_2111,N_2138);
nand U5307 (N_5307,N_3798,N_2951);
xor U5308 (N_5308,N_3492,N_2602);
nor U5309 (N_5309,N_3362,N_2914);
or U5310 (N_5310,N_2420,N_2499);
or U5311 (N_5311,N_3979,N_3364);
nand U5312 (N_5312,N_3702,N_3818);
or U5313 (N_5313,N_3146,N_2008);
nor U5314 (N_5314,N_2621,N_2591);
nand U5315 (N_5315,N_2624,N_2053);
nor U5316 (N_5316,N_3998,N_3206);
or U5317 (N_5317,N_3089,N_2605);
nor U5318 (N_5318,N_2891,N_2120);
and U5319 (N_5319,N_2071,N_2922);
nor U5320 (N_5320,N_3912,N_2652);
nand U5321 (N_5321,N_3254,N_3910);
nor U5322 (N_5322,N_3457,N_3596);
nor U5323 (N_5323,N_3068,N_2496);
nor U5324 (N_5324,N_3433,N_2331);
nand U5325 (N_5325,N_3033,N_2648);
nand U5326 (N_5326,N_2637,N_2102);
nor U5327 (N_5327,N_2791,N_3510);
and U5328 (N_5328,N_3679,N_3367);
or U5329 (N_5329,N_2088,N_3044);
xnor U5330 (N_5330,N_2434,N_2948);
or U5331 (N_5331,N_2391,N_2956);
or U5332 (N_5332,N_2700,N_3628);
nand U5333 (N_5333,N_3289,N_3045);
or U5334 (N_5334,N_2862,N_2970);
nor U5335 (N_5335,N_3074,N_2907);
or U5336 (N_5336,N_3696,N_3033);
nor U5337 (N_5337,N_3387,N_2000);
nand U5338 (N_5338,N_2624,N_2806);
nor U5339 (N_5339,N_2663,N_3288);
nor U5340 (N_5340,N_3226,N_2601);
and U5341 (N_5341,N_3768,N_2847);
and U5342 (N_5342,N_3137,N_3862);
nand U5343 (N_5343,N_3175,N_2476);
nand U5344 (N_5344,N_2363,N_3049);
nor U5345 (N_5345,N_2468,N_2658);
or U5346 (N_5346,N_3817,N_2860);
and U5347 (N_5347,N_3228,N_2229);
nand U5348 (N_5348,N_2162,N_2662);
nor U5349 (N_5349,N_2832,N_3029);
xnor U5350 (N_5350,N_2784,N_3071);
xor U5351 (N_5351,N_3750,N_2020);
and U5352 (N_5352,N_3534,N_3638);
nand U5353 (N_5353,N_3093,N_2275);
and U5354 (N_5354,N_3329,N_2321);
nor U5355 (N_5355,N_2093,N_2383);
xnor U5356 (N_5356,N_2723,N_2931);
nand U5357 (N_5357,N_2659,N_3736);
or U5358 (N_5358,N_2929,N_3541);
nor U5359 (N_5359,N_3459,N_3091);
or U5360 (N_5360,N_3608,N_3566);
nand U5361 (N_5361,N_3831,N_3672);
and U5362 (N_5362,N_3122,N_2380);
nor U5363 (N_5363,N_2963,N_2052);
nor U5364 (N_5364,N_3877,N_3278);
or U5365 (N_5365,N_2791,N_3547);
and U5366 (N_5366,N_2652,N_3818);
nor U5367 (N_5367,N_3260,N_2753);
or U5368 (N_5368,N_3325,N_2791);
or U5369 (N_5369,N_2831,N_2185);
nor U5370 (N_5370,N_2499,N_3353);
xor U5371 (N_5371,N_2124,N_2215);
and U5372 (N_5372,N_2467,N_3751);
or U5373 (N_5373,N_3577,N_3045);
and U5374 (N_5374,N_2217,N_2150);
nor U5375 (N_5375,N_3346,N_3451);
xor U5376 (N_5376,N_2307,N_2829);
or U5377 (N_5377,N_2941,N_3762);
or U5378 (N_5378,N_2277,N_3514);
xnor U5379 (N_5379,N_2946,N_2754);
nor U5380 (N_5380,N_3243,N_3282);
or U5381 (N_5381,N_3852,N_2815);
and U5382 (N_5382,N_2657,N_3517);
nand U5383 (N_5383,N_3437,N_3398);
nor U5384 (N_5384,N_3927,N_2806);
nand U5385 (N_5385,N_3961,N_3637);
nor U5386 (N_5386,N_2674,N_3626);
and U5387 (N_5387,N_2570,N_2853);
or U5388 (N_5388,N_2762,N_3194);
nor U5389 (N_5389,N_3544,N_3253);
or U5390 (N_5390,N_2912,N_3208);
nand U5391 (N_5391,N_3611,N_2751);
nand U5392 (N_5392,N_3082,N_3648);
nor U5393 (N_5393,N_3026,N_3539);
nand U5394 (N_5394,N_3017,N_2171);
or U5395 (N_5395,N_2079,N_2363);
nor U5396 (N_5396,N_3511,N_3687);
and U5397 (N_5397,N_3634,N_2847);
xnor U5398 (N_5398,N_2370,N_3503);
xnor U5399 (N_5399,N_2054,N_2208);
and U5400 (N_5400,N_3437,N_2311);
or U5401 (N_5401,N_2455,N_3381);
nand U5402 (N_5402,N_2254,N_3522);
xor U5403 (N_5403,N_3480,N_2609);
nand U5404 (N_5404,N_3760,N_2668);
or U5405 (N_5405,N_2247,N_3203);
or U5406 (N_5406,N_3740,N_3515);
nor U5407 (N_5407,N_3161,N_3340);
nor U5408 (N_5408,N_2811,N_2243);
nand U5409 (N_5409,N_2707,N_3440);
nor U5410 (N_5410,N_2093,N_3071);
and U5411 (N_5411,N_3390,N_2411);
or U5412 (N_5412,N_3854,N_3712);
nor U5413 (N_5413,N_2849,N_2057);
nor U5414 (N_5414,N_2432,N_2829);
nor U5415 (N_5415,N_3528,N_2617);
nand U5416 (N_5416,N_2910,N_3559);
or U5417 (N_5417,N_3439,N_2523);
and U5418 (N_5418,N_3375,N_2248);
or U5419 (N_5419,N_2376,N_3994);
xor U5420 (N_5420,N_3833,N_3139);
or U5421 (N_5421,N_2110,N_2748);
nor U5422 (N_5422,N_2601,N_2867);
and U5423 (N_5423,N_2024,N_3047);
nor U5424 (N_5424,N_3810,N_2885);
nor U5425 (N_5425,N_2913,N_3452);
and U5426 (N_5426,N_3252,N_2135);
nand U5427 (N_5427,N_3152,N_2493);
and U5428 (N_5428,N_3362,N_2941);
nand U5429 (N_5429,N_3799,N_3422);
nand U5430 (N_5430,N_2503,N_2603);
or U5431 (N_5431,N_3528,N_3399);
or U5432 (N_5432,N_2887,N_2901);
nor U5433 (N_5433,N_2401,N_2122);
and U5434 (N_5434,N_3787,N_2917);
and U5435 (N_5435,N_2429,N_2134);
and U5436 (N_5436,N_3519,N_3380);
and U5437 (N_5437,N_3651,N_2300);
and U5438 (N_5438,N_3883,N_3968);
and U5439 (N_5439,N_3054,N_2637);
and U5440 (N_5440,N_3036,N_3584);
or U5441 (N_5441,N_2551,N_2627);
nor U5442 (N_5442,N_3513,N_2965);
nand U5443 (N_5443,N_3762,N_3875);
xor U5444 (N_5444,N_3403,N_3802);
nor U5445 (N_5445,N_3792,N_3798);
and U5446 (N_5446,N_3680,N_3382);
xnor U5447 (N_5447,N_3120,N_2836);
xnor U5448 (N_5448,N_2180,N_3009);
and U5449 (N_5449,N_3790,N_3740);
nand U5450 (N_5450,N_2651,N_3576);
nand U5451 (N_5451,N_2525,N_2460);
and U5452 (N_5452,N_3477,N_3003);
nor U5453 (N_5453,N_2714,N_3697);
nand U5454 (N_5454,N_2723,N_2255);
nor U5455 (N_5455,N_3488,N_2058);
nor U5456 (N_5456,N_3940,N_3480);
and U5457 (N_5457,N_2225,N_3172);
or U5458 (N_5458,N_2711,N_3454);
nor U5459 (N_5459,N_2159,N_3160);
nand U5460 (N_5460,N_3835,N_3241);
nor U5461 (N_5461,N_2652,N_2227);
xor U5462 (N_5462,N_3703,N_3620);
nor U5463 (N_5463,N_3025,N_2254);
nand U5464 (N_5464,N_2773,N_2575);
nand U5465 (N_5465,N_2979,N_3885);
xnor U5466 (N_5466,N_2415,N_3321);
and U5467 (N_5467,N_2476,N_2613);
or U5468 (N_5468,N_2567,N_3123);
nor U5469 (N_5469,N_3850,N_3683);
nor U5470 (N_5470,N_3236,N_3385);
nor U5471 (N_5471,N_3229,N_2936);
and U5472 (N_5472,N_2099,N_2862);
and U5473 (N_5473,N_2166,N_2290);
or U5474 (N_5474,N_3524,N_2384);
nand U5475 (N_5475,N_3599,N_3255);
xor U5476 (N_5476,N_2414,N_3541);
nor U5477 (N_5477,N_3510,N_2185);
nand U5478 (N_5478,N_3609,N_3759);
nor U5479 (N_5479,N_3892,N_3316);
or U5480 (N_5480,N_2342,N_2396);
xor U5481 (N_5481,N_3875,N_2858);
nor U5482 (N_5482,N_3127,N_3170);
and U5483 (N_5483,N_2452,N_3083);
and U5484 (N_5484,N_2137,N_3994);
nand U5485 (N_5485,N_3056,N_3895);
nand U5486 (N_5486,N_3719,N_3255);
or U5487 (N_5487,N_3462,N_3458);
nor U5488 (N_5488,N_3369,N_3235);
xor U5489 (N_5489,N_3595,N_3648);
nor U5490 (N_5490,N_2883,N_2512);
nor U5491 (N_5491,N_3041,N_2293);
nor U5492 (N_5492,N_2208,N_2499);
xnor U5493 (N_5493,N_2037,N_2115);
nand U5494 (N_5494,N_3059,N_3247);
nor U5495 (N_5495,N_3693,N_2193);
nand U5496 (N_5496,N_2450,N_2881);
nand U5497 (N_5497,N_2601,N_3241);
or U5498 (N_5498,N_3466,N_3172);
nand U5499 (N_5499,N_3433,N_3010);
nand U5500 (N_5500,N_2569,N_3344);
nor U5501 (N_5501,N_2163,N_2140);
nand U5502 (N_5502,N_3568,N_2967);
nor U5503 (N_5503,N_2585,N_3781);
or U5504 (N_5504,N_3465,N_3592);
nand U5505 (N_5505,N_3393,N_2376);
and U5506 (N_5506,N_3532,N_3457);
nor U5507 (N_5507,N_2193,N_2482);
or U5508 (N_5508,N_3193,N_2661);
nand U5509 (N_5509,N_2369,N_2292);
and U5510 (N_5510,N_2379,N_2813);
nor U5511 (N_5511,N_3087,N_3198);
nand U5512 (N_5512,N_2402,N_2453);
nor U5513 (N_5513,N_3918,N_2729);
nand U5514 (N_5514,N_3812,N_2893);
and U5515 (N_5515,N_2801,N_2791);
and U5516 (N_5516,N_2391,N_3644);
or U5517 (N_5517,N_3760,N_2349);
and U5518 (N_5518,N_2847,N_2774);
nand U5519 (N_5519,N_2408,N_3971);
nand U5520 (N_5520,N_2176,N_3057);
xor U5521 (N_5521,N_3732,N_2944);
nor U5522 (N_5522,N_2435,N_2952);
and U5523 (N_5523,N_3605,N_2864);
nor U5524 (N_5524,N_3136,N_3470);
nand U5525 (N_5525,N_3306,N_2748);
nand U5526 (N_5526,N_2435,N_2910);
nor U5527 (N_5527,N_2344,N_3396);
nand U5528 (N_5528,N_2071,N_2228);
nor U5529 (N_5529,N_3479,N_3087);
xnor U5530 (N_5530,N_3496,N_2083);
nand U5531 (N_5531,N_3767,N_3132);
nand U5532 (N_5532,N_3888,N_2804);
xor U5533 (N_5533,N_3827,N_2485);
and U5534 (N_5534,N_2532,N_2878);
nand U5535 (N_5535,N_2532,N_3542);
and U5536 (N_5536,N_2114,N_3106);
nand U5537 (N_5537,N_3268,N_2272);
xnor U5538 (N_5538,N_3157,N_3823);
nand U5539 (N_5539,N_2217,N_2570);
and U5540 (N_5540,N_2546,N_3485);
or U5541 (N_5541,N_3999,N_2437);
nor U5542 (N_5542,N_3223,N_2400);
or U5543 (N_5543,N_3863,N_2978);
nand U5544 (N_5544,N_3340,N_3512);
and U5545 (N_5545,N_2548,N_2465);
or U5546 (N_5546,N_3864,N_3433);
nand U5547 (N_5547,N_3697,N_2830);
or U5548 (N_5548,N_2114,N_3318);
nor U5549 (N_5549,N_2231,N_3052);
nand U5550 (N_5550,N_2808,N_2831);
nor U5551 (N_5551,N_3115,N_3815);
or U5552 (N_5552,N_3542,N_2706);
nor U5553 (N_5553,N_3682,N_3952);
xor U5554 (N_5554,N_3628,N_2851);
nor U5555 (N_5555,N_3512,N_3593);
nor U5556 (N_5556,N_3343,N_3751);
or U5557 (N_5557,N_3411,N_2629);
and U5558 (N_5558,N_2642,N_3771);
or U5559 (N_5559,N_2573,N_3153);
xor U5560 (N_5560,N_2433,N_2666);
nor U5561 (N_5561,N_3155,N_3842);
or U5562 (N_5562,N_2842,N_2665);
nand U5563 (N_5563,N_3516,N_2342);
nor U5564 (N_5564,N_3673,N_2131);
nor U5565 (N_5565,N_3670,N_3496);
nor U5566 (N_5566,N_3329,N_3922);
or U5567 (N_5567,N_2433,N_2356);
nand U5568 (N_5568,N_2246,N_2990);
nor U5569 (N_5569,N_3553,N_2353);
nand U5570 (N_5570,N_2731,N_2177);
xnor U5571 (N_5571,N_3519,N_2506);
or U5572 (N_5572,N_3359,N_3936);
or U5573 (N_5573,N_2754,N_2455);
nor U5574 (N_5574,N_2830,N_2714);
and U5575 (N_5575,N_3774,N_2066);
nor U5576 (N_5576,N_2538,N_2698);
and U5577 (N_5577,N_2874,N_3706);
or U5578 (N_5578,N_3012,N_2858);
and U5579 (N_5579,N_2718,N_2871);
or U5580 (N_5580,N_2386,N_2278);
xnor U5581 (N_5581,N_2047,N_3525);
and U5582 (N_5582,N_3856,N_2486);
nor U5583 (N_5583,N_3566,N_3239);
and U5584 (N_5584,N_2408,N_2296);
nand U5585 (N_5585,N_2434,N_3341);
nand U5586 (N_5586,N_2787,N_2027);
nand U5587 (N_5587,N_2384,N_2512);
or U5588 (N_5588,N_2414,N_2471);
and U5589 (N_5589,N_3741,N_2731);
or U5590 (N_5590,N_3268,N_2704);
nand U5591 (N_5591,N_3240,N_2020);
and U5592 (N_5592,N_3579,N_2204);
nor U5593 (N_5593,N_3373,N_3389);
nor U5594 (N_5594,N_3328,N_2222);
and U5595 (N_5595,N_2868,N_2201);
or U5596 (N_5596,N_2197,N_2134);
nand U5597 (N_5597,N_3026,N_3183);
and U5598 (N_5598,N_3178,N_3340);
and U5599 (N_5599,N_2774,N_2156);
and U5600 (N_5600,N_2309,N_3371);
and U5601 (N_5601,N_3065,N_3730);
xnor U5602 (N_5602,N_2479,N_3329);
nor U5603 (N_5603,N_3897,N_2034);
nand U5604 (N_5604,N_2075,N_2578);
and U5605 (N_5605,N_2991,N_3587);
nor U5606 (N_5606,N_2818,N_2932);
and U5607 (N_5607,N_2008,N_2920);
or U5608 (N_5608,N_2325,N_2818);
and U5609 (N_5609,N_2605,N_3673);
xnor U5610 (N_5610,N_3502,N_2089);
and U5611 (N_5611,N_2872,N_2143);
xnor U5612 (N_5612,N_3683,N_3820);
xor U5613 (N_5613,N_2341,N_2434);
or U5614 (N_5614,N_3553,N_3069);
nor U5615 (N_5615,N_3016,N_3884);
and U5616 (N_5616,N_2444,N_3404);
and U5617 (N_5617,N_2090,N_3124);
nand U5618 (N_5618,N_3803,N_2097);
or U5619 (N_5619,N_2153,N_2254);
or U5620 (N_5620,N_2146,N_2989);
xnor U5621 (N_5621,N_3660,N_2531);
or U5622 (N_5622,N_3190,N_3665);
and U5623 (N_5623,N_2686,N_3663);
nor U5624 (N_5624,N_2737,N_3664);
nor U5625 (N_5625,N_3044,N_2948);
xnor U5626 (N_5626,N_2595,N_3996);
or U5627 (N_5627,N_3268,N_3471);
nor U5628 (N_5628,N_2797,N_3028);
and U5629 (N_5629,N_3783,N_2016);
or U5630 (N_5630,N_2454,N_2304);
xor U5631 (N_5631,N_3027,N_3598);
xor U5632 (N_5632,N_3074,N_2060);
nor U5633 (N_5633,N_3436,N_3566);
or U5634 (N_5634,N_2834,N_2630);
nand U5635 (N_5635,N_3134,N_2850);
and U5636 (N_5636,N_2434,N_2345);
and U5637 (N_5637,N_2693,N_3406);
and U5638 (N_5638,N_2870,N_2214);
nor U5639 (N_5639,N_3609,N_2894);
or U5640 (N_5640,N_2233,N_2022);
xnor U5641 (N_5641,N_2504,N_3966);
and U5642 (N_5642,N_3117,N_2341);
or U5643 (N_5643,N_3695,N_2631);
nor U5644 (N_5644,N_2434,N_2230);
nand U5645 (N_5645,N_3289,N_2761);
and U5646 (N_5646,N_3161,N_3750);
or U5647 (N_5647,N_3266,N_2140);
nand U5648 (N_5648,N_2739,N_3778);
nand U5649 (N_5649,N_2356,N_2672);
and U5650 (N_5650,N_2689,N_2376);
nand U5651 (N_5651,N_2206,N_2408);
nor U5652 (N_5652,N_3502,N_2381);
nand U5653 (N_5653,N_3192,N_3726);
and U5654 (N_5654,N_2307,N_2482);
nor U5655 (N_5655,N_3584,N_3089);
nor U5656 (N_5656,N_2314,N_2799);
or U5657 (N_5657,N_3005,N_3467);
xor U5658 (N_5658,N_3654,N_3966);
or U5659 (N_5659,N_2076,N_2089);
nand U5660 (N_5660,N_3070,N_3885);
xnor U5661 (N_5661,N_3223,N_2387);
nor U5662 (N_5662,N_2349,N_2967);
nor U5663 (N_5663,N_3091,N_3151);
or U5664 (N_5664,N_2519,N_3551);
nand U5665 (N_5665,N_2269,N_2373);
or U5666 (N_5666,N_3002,N_3229);
nand U5667 (N_5667,N_2778,N_3764);
nand U5668 (N_5668,N_3250,N_2898);
nor U5669 (N_5669,N_3619,N_2366);
and U5670 (N_5670,N_3404,N_3058);
nand U5671 (N_5671,N_3908,N_2604);
or U5672 (N_5672,N_3188,N_2298);
or U5673 (N_5673,N_2714,N_2223);
and U5674 (N_5674,N_3813,N_3381);
or U5675 (N_5675,N_3867,N_3270);
or U5676 (N_5676,N_3351,N_2283);
or U5677 (N_5677,N_2101,N_3178);
or U5678 (N_5678,N_2661,N_3035);
and U5679 (N_5679,N_3616,N_3319);
nand U5680 (N_5680,N_3986,N_2574);
and U5681 (N_5681,N_2227,N_3523);
or U5682 (N_5682,N_3520,N_3012);
nor U5683 (N_5683,N_3068,N_3312);
or U5684 (N_5684,N_2968,N_3917);
and U5685 (N_5685,N_2015,N_2177);
or U5686 (N_5686,N_2119,N_2031);
or U5687 (N_5687,N_2673,N_2642);
nand U5688 (N_5688,N_2824,N_3763);
nand U5689 (N_5689,N_2714,N_3847);
xor U5690 (N_5690,N_3688,N_3765);
nor U5691 (N_5691,N_2070,N_3846);
xnor U5692 (N_5692,N_3846,N_3877);
or U5693 (N_5693,N_3190,N_3691);
or U5694 (N_5694,N_2428,N_2112);
and U5695 (N_5695,N_2908,N_3915);
nand U5696 (N_5696,N_2790,N_3185);
xnor U5697 (N_5697,N_3154,N_2134);
xor U5698 (N_5698,N_3433,N_3861);
or U5699 (N_5699,N_3986,N_2437);
nand U5700 (N_5700,N_3878,N_2917);
nor U5701 (N_5701,N_3094,N_2773);
nor U5702 (N_5702,N_3080,N_2483);
nand U5703 (N_5703,N_3252,N_2939);
nor U5704 (N_5704,N_3242,N_2565);
or U5705 (N_5705,N_2410,N_2092);
nor U5706 (N_5706,N_3437,N_3032);
nor U5707 (N_5707,N_3031,N_2172);
nand U5708 (N_5708,N_3696,N_3112);
nand U5709 (N_5709,N_3067,N_2255);
nand U5710 (N_5710,N_2764,N_2586);
nand U5711 (N_5711,N_3766,N_2135);
xnor U5712 (N_5712,N_2979,N_3263);
and U5713 (N_5713,N_3423,N_2413);
or U5714 (N_5714,N_2873,N_3446);
nand U5715 (N_5715,N_3056,N_2087);
and U5716 (N_5716,N_2580,N_2605);
xor U5717 (N_5717,N_2901,N_2076);
nand U5718 (N_5718,N_3165,N_3323);
nor U5719 (N_5719,N_2235,N_3393);
xor U5720 (N_5720,N_2024,N_3350);
and U5721 (N_5721,N_2652,N_2737);
or U5722 (N_5722,N_3697,N_3087);
nor U5723 (N_5723,N_3076,N_2113);
nor U5724 (N_5724,N_3523,N_2188);
and U5725 (N_5725,N_2209,N_2744);
nand U5726 (N_5726,N_2151,N_2135);
xnor U5727 (N_5727,N_3740,N_2047);
nand U5728 (N_5728,N_2805,N_2402);
nor U5729 (N_5729,N_3788,N_2788);
nor U5730 (N_5730,N_3110,N_3344);
nand U5731 (N_5731,N_3303,N_2349);
xnor U5732 (N_5732,N_2358,N_2819);
and U5733 (N_5733,N_2631,N_2816);
nand U5734 (N_5734,N_3265,N_2000);
or U5735 (N_5735,N_2587,N_3190);
or U5736 (N_5736,N_3038,N_2175);
nor U5737 (N_5737,N_3265,N_3544);
xnor U5738 (N_5738,N_2101,N_2718);
or U5739 (N_5739,N_2161,N_3166);
and U5740 (N_5740,N_2872,N_2515);
or U5741 (N_5741,N_3830,N_2152);
or U5742 (N_5742,N_2566,N_2458);
nand U5743 (N_5743,N_3494,N_3726);
nand U5744 (N_5744,N_2982,N_2105);
nand U5745 (N_5745,N_3575,N_2636);
nor U5746 (N_5746,N_2681,N_2625);
nor U5747 (N_5747,N_3562,N_2353);
or U5748 (N_5748,N_2112,N_3308);
or U5749 (N_5749,N_2383,N_2512);
or U5750 (N_5750,N_2140,N_3644);
and U5751 (N_5751,N_3615,N_3745);
nand U5752 (N_5752,N_2776,N_3511);
or U5753 (N_5753,N_2641,N_3996);
nand U5754 (N_5754,N_3687,N_2723);
nand U5755 (N_5755,N_2076,N_2575);
nor U5756 (N_5756,N_2385,N_3520);
or U5757 (N_5757,N_2144,N_3286);
or U5758 (N_5758,N_2048,N_3775);
nor U5759 (N_5759,N_2561,N_2535);
nand U5760 (N_5760,N_2067,N_3907);
or U5761 (N_5761,N_2735,N_2999);
or U5762 (N_5762,N_2721,N_3783);
or U5763 (N_5763,N_3256,N_2389);
or U5764 (N_5764,N_3215,N_3458);
nand U5765 (N_5765,N_2850,N_3076);
and U5766 (N_5766,N_2845,N_3626);
nand U5767 (N_5767,N_2449,N_3807);
nand U5768 (N_5768,N_3489,N_3200);
xor U5769 (N_5769,N_2761,N_2228);
nand U5770 (N_5770,N_2906,N_3344);
nor U5771 (N_5771,N_2128,N_2135);
nor U5772 (N_5772,N_2773,N_3131);
nor U5773 (N_5773,N_2104,N_3997);
nor U5774 (N_5774,N_3699,N_3119);
nand U5775 (N_5775,N_3950,N_2545);
nor U5776 (N_5776,N_3856,N_3052);
nor U5777 (N_5777,N_3732,N_3385);
xnor U5778 (N_5778,N_2443,N_2800);
nand U5779 (N_5779,N_2213,N_2265);
and U5780 (N_5780,N_3939,N_2957);
xor U5781 (N_5781,N_3782,N_3636);
or U5782 (N_5782,N_3073,N_2350);
and U5783 (N_5783,N_3462,N_3340);
or U5784 (N_5784,N_2043,N_3593);
nand U5785 (N_5785,N_2265,N_3149);
nand U5786 (N_5786,N_2870,N_3343);
or U5787 (N_5787,N_2528,N_3863);
xnor U5788 (N_5788,N_3015,N_2624);
nor U5789 (N_5789,N_2374,N_2675);
and U5790 (N_5790,N_3505,N_2196);
and U5791 (N_5791,N_2075,N_3834);
and U5792 (N_5792,N_3636,N_3793);
or U5793 (N_5793,N_2606,N_2274);
or U5794 (N_5794,N_3186,N_3413);
nand U5795 (N_5795,N_3911,N_3972);
and U5796 (N_5796,N_2958,N_2630);
nand U5797 (N_5797,N_3721,N_2647);
and U5798 (N_5798,N_3049,N_3632);
and U5799 (N_5799,N_2516,N_2710);
xor U5800 (N_5800,N_2112,N_3190);
nor U5801 (N_5801,N_2660,N_2632);
nand U5802 (N_5802,N_2449,N_2092);
nor U5803 (N_5803,N_3362,N_3794);
and U5804 (N_5804,N_2445,N_2667);
nand U5805 (N_5805,N_2487,N_2448);
or U5806 (N_5806,N_2973,N_3678);
nand U5807 (N_5807,N_2026,N_2876);
nand U5808 (N_5808,N_3340,N_2294);
or U5809 (N_5809,N_2979,N_3405);
xnor U5810 (N_5810,N_3842,N_2093);
nand U5811 (N_5811,N_3538,N_2446);
or U5812 (N_5812,N_3559,N_2496);
nor U5813 (N_5813,N_3717,N_3492);
nand U5814 (N_5814,N_2666,N_3329);
and U5815 (N_5815,N_3940,N_2313);
nand U5816 (N_5816,N_2270,N_2409);
nor U5817 (N_5817,N_3872,N_3520);
nor U5818 (N_5818,N_2428,N_2221);
nand U5819 (N_5819,N_3039,N_3587);
xor U5820 (N_5820,N_2161,N_2321);
or U5821 (N_5821,N_3250,N_2715);
nand U5822 (N_5822,N_2610,N_3655);
nand U5823 (N_5823,N_2227,N_3388);
nand U5824 (N_5824,N_3235,N_2084);
nor U5825 (N_5825,N_3597,N_3323);
nor U5826 (N_5826,N_3737,N_3662);
xnor U5827 (N_5827,N_3951,N_2097);
nor U5828 (N_5828,N_2743,N_2235);
and U5829 (N_5829,N_3453,N_3554);
or U5830 (N_5830,N_3272,N_2186);
nand U5831 (N_5831,N_3824,N_3176);
nor U5832 (N_5832,N_2087,N_2183);
and U5833 (N_5833,N_2537,N_2527);
nor U5834 (N_5834,N_3206,N_2075);
xnor U5835 (N_5835,N_2712,N_3150);
nor U5836 (N_5836,N_2002,N_3552);
nor U5837 (N_5837,N_2818,N_2544);
and U5838 (N_5838,N_2423,N_2241);
and U5839 (N_5839,N_3093,N_3332);
or U5840 (N_5840,N_2890,N_3031);
nor U5841 (N_5841,N_3172,N_2221);
nand U5842 (N_5842,N_2710,N_3065);
nor U5843 (N_5843,N_3056,N_3175);
nor U5844 (N_5844,N_3169,N_3520);
or U5845 (N_5845,N_3872,N_3252);
xor U5846 (N_5846,N_2991,N_2451);
or U5847 (N_5847,N_2516,N_2206);
or U5848 (N_5848,N_2107,N_3342);
or U5849 (N_5849,N_3582,N_2423);
and U5850 (N_5850,N_2298,N_3496);
and U5851 (N_5851,N_3014,N_2204);
or U5852 (N_5852,N_3350,N_3228);
and U5853 (N_5853,N_3405,N_3268);
nor U5854 (N_5854,N_3435,N_3194);
and U5855 (N_5855,N_2961,N_3722);
or U5856 (N_5856,N_3102,N_2354);
nor U5857 (N_5857,N_3427,N_3888);
nand U5858 (N_5858,N_3781,N_2385);
or U5859 (N_5859,N_2402,N_2482);
nand U5860 (N_5860,N_3509,N_2423);
nor U5861 (N_5861,N_3995,N_2598);
or U5862 (N_5862,N_2401,N_3341);
nor U5863 (N_5863,N_2361,N_3635);
and U5864 (N_5864,N_3317,N_2225);
or U5865 (N_5865,N_2218,N_2570);
and U5866 (N_5866,N_3301,N_2694);
nor U5867 (N_5867,N_2282,N_3059);
nor U5868 (N_5868,N_2274,N_2744);
xnor U5869 (N_5869,N_2869,N_3969);
and U5870 (N_5870,N_2035,N_2342);
nor U5871 (N_5871,N_2968,N_2238);
nand U5872 (N_5872,N_2690,N_3019);
xnor U5873 (N_5873,N_3683,N_2317);
nand U5874 (N_5874,N_2717,N_3419);
and U5875 (N_5875,N_2593,N_3325);
nand U5876 (N_5876,N_3865,N_3935);
or U5877 (N_5877,N_3901,N_2463);
nand U5878 (N_5878,N_3481,N_2932);
nand U5879 (N_5879,N_3653,N_3772);
nand U5880 (N_5880,N_3077,N_3134);
nand U5881 (N_5881,N_2287,N_2308);
nor U5882 (N_5882,N_3271,N_3795);
nand U5883 (N_5883,N_2579,N_2811);
xor U5884 (N_5884,N_2872,N_3542);
or U5885 (N_5885,N_2861,N_2235);
nand U5886 (N_5886,N_3151,N_3930);
or U5887 (N_5887,N_3480,N_2742);
xnor U5888 (N_5888,N_3526,N_2235);
and U5889 (N_5889,N_3345,N_2607);
nand U5890 (N_5890,N_3659,N_2076);
or U5891 (N_5891,N_2390,N_3581);
nor U5892 (N_5892,N_3515,N_3721);
nor U5893 (N_5893,N_3403,N_3905);
nand U5894 (N_5894,N_2643,N_3029);
and U5895 (N_5895,N_3411,N_3916);
nor U5896 (N_5896,N_3000,N_3504);
and U5897 (N_5897,N_2524,N_2273);
xor U5898 (N_5898,N_2096,N_2386);
nor U5899 (N_5899,N_3857,N_2676);
nor U5900 (N_5900,N_2586,N_2585);
or U5901 (N_5901,N_2506,N_2381);
xnor U5902 (N_5902,N_3705,N_2746);
nor U5903 (N_5903,N_3229,N_3619);
nor U5904 (N_5904,N_2336,N_3189);
and U5905 (N_5905,N_2307,N_2661);
nor U5906 (N_5906,N_3678,N_2718);
xnor U5907 (N_5907,N_3401,N_3017);
nand U5908 (N_5908,N_3551,N_2872);
nand U5909 (N_5909,N_3445,N_2922);
or U5910 (N_5910,N_3701,N_3212);
nand U5911 (N_5911,N_3329,N_3509);
or U5912 (N_5912,N_3491,N_3422);
or U5913 (N_5913,N_3232,N_3694);
nor U5914 (N_5914,N_2193,N_2078);
and U5915 (N_5915,N_3426,N_3799);
and U5916 (N_5916,N_3977,N_3486);
or U5917 (N_5917,N_3287,N_3964);
or U5918 (N_5918,N_3366,N_3714);
nor U5919 (N_5919,N_3298,N_3743);
and U5920 (N_5920,N_2528,N_3529);
nand U5921 (N_5921,N_3473,N_3546);
nor U5922 (N_5922,N_3653,N_2714);
or U5923 (N_5923,N_2415,N_3419);
xor U5924 (N_5924,N_3889,N_2484);
nand U5925 (N_5925,N_2203,N_3400);
and U5926 (N_5926,N_2460,N_2454);
nor U5927 (N_5927,N_2382,N_2393);
xnor U5928 (N_5928,N_2901,N_3266);
nand U5929 (N_5929,N_2032,N_2599);
nor U5930 (N_5930,N_3386,N_3391);
nand U5931 (N_5931,N_3014,N_2483);
or U5932 (N_5932,N_3563,N_2074);
nor U5933 (N_5933,N_2842,N_2341);
or U5934 (N_5934,N_3872,N_3174);
and U5935 (N_5935,N_2026,N_2185);
nor U5936 (N_5936,N_3340,N_3962);
xor U5937 (N_5937,N_3060,N_2072);
nor U5938 (N_5938,N_2831,N_3016);
nor U5939 (N_5939,N_2839,N_3848);
nor U5940 (N_5940,N_3746,N_3670);
nand U5941 (N_5941,N_2256,N_3983);
xnor U5942 (N_5942,N_2790,N_2918);
nand U5943 (N_5943,N_2106,N_2150);
and U5944 (N_5944,N_2502,N_3962);
or U5945 (N_5945,N_2231,N_2282);
or U5946 (N_5946,N_2336,N_3327);
and U5947 (N_5947,N_2833,N_3739);
or U5948 (N_5948,N_3443,N_2973);
nor U5949 (N_5949,N_2558,N_3595);
and U5950 (N_5950,N_2913,N_2674);
nor U5951 (N_5951,N_2023,N_3153);
nor U5952 (N_5952,N_3002,N_3221);
and U5953 (N_5953,N_3943,N_3451);
and U5954 (N_5954,N_2696,N_3626);
and U5955 (N_5955,N_3936,N_3301);
nor U5956 (N_5956,N_2943,N_3905);
nand U5957 (N_5957,N_2012,N_3901);
or U5958 (N_5958,N_2394,N_3343);
and U5959 (N_5959,N_2870,N_3360);
and U5960 (N_5960,N_3374,N_2405);
nand U5961 (N_5961,N_3307,N_3362);
and U5962 (N_5962,N_3761,N_2755);
nand U5963 (N_5963,N_2362,N_2991);
nor U5964 (N_5964,N_3050,N_3234);
and U5965 (N_5965,N_3913,N_3744);
and U5966 (N_5966,N_2300,N_2852);
and U5967 (N_5967,N_3657,N_2925);
and U5968 (N_5968,N_3444,N_3181);
or U5969 (N_5969,N_3945,N_2684);
nand U5970 (N_5970,N_2384,N_2672);
nor U5971 (N_5971,N_3502,N_2755);
or U5972 (N_5972,N_2546,N_3834);
nand U5973 (N_5973,N_2179,N_3542);
nor U5974 (N_5974,N_3372,N_3346);
xor U5975 (N_5975,N_3275,N_3479);
and U5976 (N_5976,N_2110,N_3891);
and U5977 (N_5977,N_3055,N_2670);
nand U5978 (N_5978,N_3885,N_2953);
nor U5979 (N_5979,N_2255,N_2430);
nor U5980 (N_5980,N_2634,N_3782);
or U5981 (N_5981,N_2668,N_2381);
or U5982 (N_5982,N_3523,N_2798);
nand U5983 (N_5983,N_3046,N_2790);
and U5984 (N_5984,N_2044,N_2112);
nor U5985 (N_5985,N_3588,N_3887);
and U5986 (N_5986,N_2127,N_2341);
nor U5987 (N_5987,N_2147,N_2023);
nor U5988 (N_5988,N_2876,N_3729);
or U5989 (N_5989,N_2910,N_3054);
and U5990 (N_5990,N_3840,N_3809);
or U5991 (N_5991,N_3447,N_2989);
or U5992 (N_5992,N_2841,N_3031);
or U5993 (N_5993,N_2715,N_2244);
and U5994 (N_5994,N_3375,N_2829);
and U5995 (N_5995,N_2953,N_2128);
nor U5996 (N_5996,N_2802,N_2976);
nand U5997 (N_5997,N_3721,N_2977);
and U5998 (N_5998,N_2071,N_2117);
xnor U5999 (N_5999,N_3823,N_2602);
and U6000 (N_6000,N_5860,N_5849);
and U6001 (N_6001,N_5581,N_5178);
nor U6002 (N_6002,N_4084,N_5437);
nor U6003 (N_6003,N_4006,N_4766);
nor U6004 (N_6004,N_4833,N_5946);
nand U6005 (N_6005,N_4765,N_4050);
or U6006 (N_6006,N_4018,N_4294);
and U6007 (N_6007,N_4751,N_5708);
nand U6008 (N_6008,N_4714,N_5229);
and U6009 (N_6009,N_4260,N_5249);
or U6010 (N_6010,N_5185,N_5538);
nand U6011 (N_6011,N_4355,N_4205);
or U6012 (N_6012,N_4853,N_4878);
and U6013 (N_6013,N_5638,N_4510);
and U6014 (N_6014,N_4204,N_5225);
nand U6015 (N_6015,N_4772,N_5092);
and U6016 (N_6016,N_4224,N_5498);
nand U6017 (N_6017,N_4841,N_5093);
nand U6018 (N_6018,N_4379,N_5692);
and U6019 (N_6019,N_5293,N_4791);
nor U6020 (N_6020,N_4614,N_4467);
nand U6021 (N_6021,N_4067,N_4960);
and U6022 (N_6022,N_5909,N_5806);
nand U6023 (N_6023,N_4316,N_5248);
and U6024 (N_6024,N_5877,N_5369);
nor U6025 (N_6025,N_5505,N_4807);
xor U6026 (N_6026,N_4547,N_4984);
nand U6027 (N_6027,N_4402,N_4832);
or U6028 (N_6028,N_4415,N_5868);
or U6029 (N_6029,N_4195,N_5556);
nor U6030 (N_6030,N_4210,N_5281);
or U6031 (N_6031,N_4054,N_5690);
or U6032 (N_6032,N_4673,N_4637);
nor U6033 (N_6033,N_4908,N_4008);
nand U6034 (N_6034,N_5375,N_4813);
and U6035 (N_6035,N_4460,N_4610);
and U6036 (N_6036,N_4362,N_4145);
nand U6037 (N_6037,N_4520,N_4571);
or U6038 (N_6038,N_5965,N_5425);
or U6039 (N_6039,N_4289,N_5964);
nor U6040 (N_6040,N_4444,N_5857);
nor U6041 (N_6041,N_4948,N_5183);
nand U6042 (N_6042,N_5450,N_5537);
or U6043 (N_6043,N_5606,N_5603);
nand U6044 (N_6044,N_5963,N_5753);
nand U6045 (N_6045,N_5101,N_4053);
and U6046 (N_6046,N_5641,N_4315);
xnor U6047 (N_6047,N_5910,N_5379);
and U6048 (N_6048,N_5940,N_4425);
or U6049 (N_6049,N_5215,N_5046);
nor U6050 (N_6050,N_5374,N_5322);
and U6051 (N_6051,N_5640,N_4662);
and U6052 (N_6052,N_4469,N_4836);
and U6053 (N_6053,N_4449,N_5770);
nor U6054 (N_6054,N_5604,N_5502);
xnor U6055 (N_6055,N_5053,N_4017);
and U6056 (N_6056,N_5095,N_4917);
nand U6057 (N_6057,N_4704,N_5162);
or U6058 (N_6058,N_4648,N_5722);
xor U6059 (N_6059,N_4870,N_4789);
xnor U6060 (N_6060,N_5099,N_5411);
nor U6061 (N_6061,N_4033,N_5831);
or U6062 (N_6062,N_4756,N_5930);
nand U6063 (N_6063,N_5810,N_4007);
or U6064 (N_6064,N_5888,N_5440);
nor U6065 (N_6065,N_4334,N_4919);
and U6066 (N_6066,N_5359,N_5491);
or U6067 (N_6067,N_4574,N_5022);
or U6068 (N_6068,N_4753,N_4335);
nand U6069 (N_6069,N_4345,N_5438);
nand U6070 (N_6070,N_5253,N_5230);
xnor U6071 (N_6071,N_5886,N_5625);
and U6072 (N_6072,N_5864,N_5325);
or U6073 (N_6073,N_5752,N_4521);
nand U6074 (N_6074,N_5371,N_5034);
nor U6075 (N_6075,N_5207,N_4578);
xnor U6076 (N_6076,N_4589,N_5203);
or U6077 (N_6077,N_5519,N_4906);
nand U6078 (N_6078,N_5482,N_5064);
nor U6079 (N_6079,N_4758,N_5144);
nor U6080 (N_6080,N_4428,N_4868);
and U6081 (N_6081,N_4617,N_4422);
or U6082 (N_6082,N_4681,N_4604);
or U6083 (N_6083,N_5647,N_5624);
or U6084 (N_6084,N_5589,N_4981);
xor U6085 (N_6085,N_4800,N_5004);
nor U6086 (N_6086,N_4650,N_5786);
nand U6087 (N_6087,N_5805,N_5989);
xor U6088 (N_6088,N_5789,N_5358);
or U6089 (N_6089,N_4044,N_5259);
or U6090 (N_6090,N_4546,N_5470);
nor U6091 (N_6091,N_5572,N_4944);
or U6092 (N_6092,N_4723,N_4667);
nand U6093 (N_6093,N_4707,N_5009);
nand U6094 (N_6094,N_4351,N_5191);
or U6095 (N_6095,N_4186,N_4646);
nand U6096 (N_6096,N_5173,N_4462);
nand U6097 (N_6097,N_5055,N_4200);
nor U6098 (N_6098,N_5585,N_5209);
or U6099 (N_6099,N_5509,N_4343);
or U6100 (N_6100,N_5315,N_4682);
and U6101 (N_6101,N_5829,N_5068);
and U6102 (N_6102,N_4923,N_5887);
nand U6103 (N_6103,N_4603,N_5146);
nor U6104 (N_6104,N_5620,N_5762);
nor U6105 (N_6105,N_4111,N_5199);
or U6106 (N_6106,N_4341,N_4702);
nand U6107 (N_6107,N_4471,N_4935);
xnor U6108 (N_6108,N_5266,N_5952);
and U6109 (N_6109,N_5891,N_5390);
nand U6110 (N_6110,N_4119,N_5736);
and U6111 (N_6111,N_5731,N_4697);
nor U6112 (N_6112,N_5244,N_5923);
nor U6113 (N_6113,N_4158,N_4430);
nor U6114 (N_6114,N_4312,N_5723);
and U6115 (N_6115,N_4222,N_4194);
xor U6116 (N_6116,N_5221,N_5196);
or U6117 (N_6117,N_4403,N_4463);
xor U6118 (N_6118,N_5555,N_4391);
and U6119 (N_6119,N_4573,N_4097);
nand U6120 (N_6120,N_5846,N_5847);
xor U6121 (N_6121,N_5681,N_4942);
xnor U6122 (N_6122,N_5597,N_4470);
and U6123 (N_6123,N_4846,N_4152);
and U6124 (N_6124,N_5160,N_4699);
and U6125 (N_6125,N_4827,N_5531);
or U6126 (N_6126,N_5205,N_4554);
nor U6127 (N_6127,N_5214,N_4619);
and U6128 (N_6128,N_4086,N_5894);
or U6129 (N_6129,N_4559,N_5635);
and U6130 (N_6130,N_4472,N_5168);
and U6131 (N_6131,N_4635,N_5982);
nand U6132 (N_6132,N_4142,N_5284);
or U6133 (N_6133,N_4065,N_4767);
xnor U6134 (N_6134,N_5151,N_5968);
nor U6135 (N_6135,N_4598,N_4980);
nor U6136 (N_6136,N_5458,N_5815);
and U6137 (N_6137,N_4639,N_4251);
nand U6138 (N_6138,N_5112,N_4239);
nand U6139 (N_6139,N_5003,N_5002);
nand U6140 (N_6140,N_5693,N_4214);
and U6141 (N_6141,N_5525,N_5302);
or U6142 (N_6142,N_5190,N_5659);
and U6143 (N_6143,N_4115,N_5686);
nand U6144 (N_6144,N_4911,N_4092);
nor U6145 (N_6145,N_4668,N_5251);
nor U6146 (N_6146,N_4277,N_4551);
and U6147 (N_6147,N_4404,N_4620);
nand U6148 (N_6148,N_4154,N_5993);
nor U6149 (N_6149,N_4708,N_4830);
and U6150 (N_6150,N_5258,N_4584);
and U6151 (N_6151,N_4144,N_5662);
nor U6152 (N_6152,N_4529,N_4882);
xor U6153 (N_6153,N_5582,N_4722);
or U6154 (N_6154,N_5828,N_5245);
and U6155 (N_6155,N_4419,N_4778);
nor U6156 (N_6156,N_4212,N_5726);
and U6157 (N_6157,N_4934,N_4601);
xor U6158 (N_6158,N_5674,N_5718);
nor U6159 (N_6159,N_4188,N_4450);
or U6160 (N_6160,N_4310,N_5404);
nor U6161 (N_6161,N_4004,N_5447);
and U6162 (N_6162,N_4622,N_4630);
or U6163 (N_6163,N_5468,N_5277);
nand U6164 (N_6164,N_5592,N_5439);
nor U6165 (N_6165,N_5433,N_5524);
or U6166 (N_6166,N_5759,N_5171);
nand U6167 (N_6167,N_5944,N_5755);
xor U6168 (N_6168,N_5774,N_5899);
or U6169 (N_6169,N_4649,N_5626);
xor U6170 (N_6170,N_5430,N_5552);
or U6171 (N_6171,N_5432,N_4728);
nand U6172 (N_6172,N_5106,N_4515);
xor U6173 (N_6173,N_5410,N_4609);
xnor U6174 (N_6174,N_5649,N_5901);
nor U6175 (N_6175,N_4180,N_4040);
nand U6176 (N_6176,N_4737,N_4393);
nor U6177 (N_6177,N_4417,N_4112);
nand U6178 (N_6178,N_5347,N_4982);
nand U6179 (N_6179,N_4406,N_4059);
xor U6180 (N_6180,N_5902,N_5826);
and U6181 (N_6181,N_4783,N_4692);
or U6182 (N_6182,N_4325,N_4150);
nor U6183 (N_6183,N_4465,N_5486);
nor U6184 (N_6184,N_5969,N_5085);
nand U6185 (N_6185,N_5932,N_4002);
nand U6186 (N_6186,N_5750,N_4411);
xor U6187 (N_6187,N_4856,N_4439);
or U6188 (N_6188,N_5271,N_4250);
and U6189 (N_6189,N_5282,N_5361);
nor U6190 (N_6190,N_4103,N_5445);
and U6191 (N_6191,N_4215,N_5181);
or U6192 (N_6192,N_4326,N_4922);
or U6193 (N_6193,N_5596,N_4275);
and U6194 (N_6194,N_5970,N_5599);
nand U6195 (N_6195,N_4716,N_5741);
or U6196 (N_6196,N_4322,N_4179);
and U6197 (N_6197,N_5986,N_5514);
nor U6198 (N_6198,N_5072,N_4485);
nor U6199 (N_6199,N_4132,N_4517);
nand U6200 (N_6200,N_5621,N_4745);
nand U6201 (N_6201,N_4433,N_4812);
or U6202 (N_6202,N_5320,N_4739);
and U6203 (N_6203,N_4400,N_5273);
nor U6204 (N_6204,N_5906,N_4500);
nand U6205 (N_6205,N_5286,N_4628);
nor U6206 (N_6206,N_4234,N_4509);
and U6207 (N_6207,N_5136,N_4558);
xor U6208 (N_6208,N_5922,N_4687);
nor U6209 (N_6209,N_5100,N_4370);
and U6210 (N_6210,N_4475,N_5794);
xnor U6211 (N_6211,N_4136,N_4997);
nand U6212 (N_6212,N_4424,N_4892);
nand U6213 (N_6213,N_4397,N_4976);
or U6214 (N_6214,N_4057,N_4265);
nor U6215 (N_6215,N_4255,N_5567);
nand U6216 (N_6216,N_4973,N_4837);
and U6217 (N_6217,N_5123,N_4503);
xnor U6218 (N_6218,N_5554,N_5078);
or U6219 (N_6219,N_4261,N_4652);
or U6220 (N_6220,N_4688,N_5462);
nor U6221 (N_6221,N_4993,N_4090);
or U6222 (N_6222,N_5813,N_4694);
nor U6223 (N_6223,N_4576,N_5878);
nand U6224 (N_6224,N_4641,N_4887);
and U6225 (N_6225,N_4700,N_5116);
nand U6226 (N_6226,N_5051,N_5811);
and U6227 (N_6227,N_4389,N_5962);
or U6228 (N_6228,N_5296,N_5623);
or U6229 (N_6229,N_5141,N_5569);
and U6230 (N_6230,N_5709,N_4690);
nor U6231 (N_6231,N_5330,N_5177);
and U6232 (N_6232,N_5147,N_5466);
and U6233 (N_6233,N_4219,N_4109);
or U6234 (N_6234,N_5074,N_4476);
or U6235 (N_6235,N_5052,N_4137);
xnor U6236 (N_6236,N_4254,N_4491);
or U6237 (N_6237,N_5619,N_5355);
or U6238 (N_6238,N_5639,N_5740);
nor U6239 (N_6239,N_5598,N_4534);
xnor U6240 (N_6240,N_5023,N_5010);
nand U6241 (N_6241,N_5685,N_4718);
or U6242 (N_6242,N_5668,N_5381);
xor U6243 (N_6243,N_5213,N_5073);
or U6244 (N_6244,N_4110,N_5084);
or U6245 (N_6245,N_4927,N_5063);
nand U6246 (N_6246,N_4918,N_4658);
nand U6247 (N_6247,N_4660,N_5795);
or U6248 (N_6248,N_4049,N_5754);
xor U6249 (N_6249,N_4062,N_5285);
or U6250 (N_6250,N_5992,N_4149);
or U6251 (N_6251,N_5176,N_4030);
and U6252 (N_6252,N_4867,N_5953);
and U6253 (N_6253,N_5911,N_4986);
nor U6254 (N_6254,N_4299,N_5070);
or U6255 (N_6255,N_5883,N_5687);
or U6256 (N_6256,N_5819,N_5274);
xnor U6257 (N_6257,N_5840,N_5839);
nor U6258 (N_6258,N_5479,N_4105);
or U6259 (N_6259,N_5204,N_5672);
nor U6260 (N_6260,N_4955,N_4327);
nor U6261 (N_6261,N_5545,N_5506);
xor U6262 (N_6262,N_5861,N_4169);
or U6263 (N_6263,N_4556,N_4123);
nor U6264 (N_6264,N_5384,N_4845);
and U6265 (N_6265,N_5169,N_4468);
nor U6266 (N_6266,N_5885,N_5903);
and U6267 (N_6267,N_4271,N_5825);
nor U6268 (N_6268,N_4615,N_4068);
nand U6269 (N_6269,N_5412,N_4645);
and U6270 (N_6270,N_5928,N_5108);
nand U6271 (N_6271,N_4877,N_5987);
nand U6272 (N_6272,N_5435,N_5316);
or U6273 (N_6273,N_4930,N_4596);
xor U6274 (N_6274,N_5027,N_4875);
nor U6275 (N_6275,N_5735,N_5793);
nor U6276 (N_6276,N_4020,N_4651);
nand U6277 (N_6277,N_5747,N_5790);
xor U6278 (N_6278,N_5311,N_4139);
and U6279 (N_6279,N_4037,N_5998);
and U6280 (N_6280,N_4931,N_5201);
nand U6281 (N_6281,N_4602,N_5362);
nor U6282 (N_6282,N_4323,N_4258);
nand U6283 (N_6283,N_5239,N_5796);
and U6284 (N_6284,N_4752,N_4907);
and U6285 (N_6285,N_5310,N_4954);
nor U6286 (N_6286,N_5919,N_5182);
and U6287 (N_6287,N_4599,N_4073);
nor U6288 (N_6288,N_5905,N_4296);
nand U6289 (N_6289,N_4512,N_5223);
and U6290 (N_6290,N_4587,N_5508);
and U6291 (N_6291,N_5131,N_5712);
and U6292 (N_6292,N_4039,N_4691);
or U6293 (N_6293,N_4496,N_5104);
and U6294 (N_6294,N_5044,N_4553);
nor U6295 (N_6295,N_4525,N_5247);
or U6296 (N_6296,N_5695,N_4542);
nor U6297 (N_6297,N_5563,N_5580);
or U6298 (N_6298,N_5113,N_5988);
or U6299 (N_6299,N_5079,N_5356);
nor U6300 (N_6300,N_5276,N_4297);
or U6301 (N_6301,N_5490,N_4543);
nand U6302 (N_6302,N_5038,N_4865);
nor U6303 (N_6303,N_4481,N_4001);
nand U6304 (N_6304,N_4191,N_5646);
nand U6305 (N_6305,N_5724,N_4202);
or U6306 (N_6306,N_5817,N_4815);
or U6307 (N_6307,N_5957,N_4307);
or U6308 (N_6308,N_5842,N_4611);
nor U6309 (N_6309,N_4101,N_5118);
and U6310 (N_6310,N_5518,N_5163);
and U6311 (N_6311,N_5283,N_4899);
and U6312 (N_6312,N_4834,N_4859);
nor U6313 (N_6313,N_5577,N_4431);
or U6314 (N_6314,N_4771,N_5391);
nand U6315 (N_6315,N_4134,N_4374);
nand U6316 (N_6316,N_4060,N_5855);
nor U6317 (N_6317,N_4285,N_5611);
nor U6318 (N_6318,N_4147,N_5780);
nor U6319 (N_6319,N_5977,N_5443);
nand U6320 (N_6320,N_4157,N_5226);
nor U6321 (N_6321,N_5727,N_4803);
nand U6322 (N_6322,N_4064,N_4042);
nor U6323 (N_6323,N_5497,N_4840);
and U6324 (N_6324,N_4790,N_4211);
nor U6325 (N_6325,N_4113,N_5816);
nor U6326 (N_6326,N_5985,N_4146);
nor U6327 (N_6327,N_5551,N_5870);
or U6328 (N_6328,N_4898,N_4757);
nand U6329 (N_6329,N_5526,N_4706);
or U6330 (N_6330,N_5880,N_5405);
nor U6331 (N_6331,N_5387,N_5363);
or U6332 (N_6332,N_5318,N_5544);
and U6333 (N_6333,N_5013,N_5973);
and U6334 (N_6334,N_5189,N_4367);
or U6335 (N_6335,N_4618,N_4066);
nor U6336 (N_6336,N_4924,N_4349);
and U6337 (N_6337,N_4184,N_5689);
and U6338 (N_6338,N_4929,N_4014);
and U6339 (N_6339,N_5610,N_5584);
xnor U6340 (N_6340,N_5395,N_5671);
nand U6341 (N_6341,N_5769,N_4028);
nand U6342 (N_6342,N_4860,N_5561);
or U6343 (N_6343,N_4987,N_5489);
or U6344 (N_6344,N_5801,N_4990);
nand U6345 (N_6345,N_5061,N_5557);
and U6346 (N_6346,N_4356,N_5820);
and U6347 (N_6347,N_4552,N_4290);
nand U6348 (N_6348,N_4544,N_5730);
nor U6349 (N_6349,N_5667,N_4979);
nor U6350 (N_6350,N_4394,N_4489);
or U6351 (N_6351,N_5488,N_4769);
xor U6352 (N_6352,N_5742,N_4705);
xnor U6353 (N_6353,N_5416,N_5393);
nand U6354 (N_6354,N_5081,N_4365);
xor U6355 (N_6355,N_4183,N_5351);
and U6356 (N_6356,N_4339,N_5788);
or U6357 (N_6357,N_4087,N_4616);
nor U6358 (N_6358,N_4644,N_5045);
nor U6359 (N_6359,N_4664,N_5339);
or U6360 (N_6360,N_4118,N_4484);
nor U6361 (N_6361,N_4088,N_5429);
nand U6362 (N_6362,N_4125,N_5423);
xor U6363 (N_6363,N_4161,N_4773);
nand U6364 (N_6364,N_5539,N_5630);
or U6365 (N_6365,N_5049,N_5926);
and U6366 (N_6366,N_4385,N_5991);
and U6367 (N_6367,N_5814,N_4114);
nand U6368 (N_6368,N_4155,N_4328);
nor U6369 (N_6369,N_5756,N_4392);
xor U6370 (N_6370,N_5837,N_4715);
xnor U6371 (N_6371,N_5420,N_4776);
or U6372 (N_6372,N_5924,N_5260);
nor U6373 (N_6373,N_5622,N_5958);
nor U6374 (N_6374,N_4881,N_5083);
nor U6375 (N_6375,N_4130,N_4932);
or U6376 (N_6376,N_5377,N_4458);
xnor U6377 (N_6377,N_5553,N_5135);
and U6378 (N_6378,N_5366,N_5874);
nor U6379 (N_6379,N_5008,N_5783);
xor U6380 (N_6380,N_4770,N_5757);
and U6381 (N_6381,N_5507,N_4089);
or U6382 (N_6382,N_5001,N_4540);
and U6383 (N_6383,N_5441,N_4902);
and U6384 (N_6384,N_4647,N_5396);
and U6385 (N_6385,N_5843,N_4124);
and U6386 (N_6386,N_5132,N_5800);
or U6387 (N_6387,N_4075,N_4304);
nand U6388 (N_6388,N_4683,N_4654);
and U6389 (N_6389,N_4093,N_4903);
nor U6390 (N_6390,N_5663,N_5609);
nand U6391 (N_6391,N_4872,N_4741);
and U6392 (N_6392,N_5595,N_5124);
and U6393 (N_6393,N_5210,N_5453);
xnor U6394 (N_6394,N_5402,N_4880);
or U6395 (N_6395,N_4848,N_4809);
and U6396 (N_6396,N_5446,N_5863);
or U6397 (N_6397,N_5219,N_4711);
nor U6398 (N_6398,N_4989,N_5541);
or U6399 (N_6399,N_5459,N_4457);
or U6400 (N_6400,N_4177,N_4873);
nor U6401 (N_6401,N_4350,N_4170);
nand U6402 (N_6402,N_5702,N_4826);
and U6403 (N_6403,N_4505,N_5494);
nand U6404 (N_6404,N_5900,N_5130);
nor U6405 (N_6405,N_4223,N_5385);
and U6406 (N_6406,N_5020,N_4975);
and U6407 (N_6407,N_4861,N_4862);
and U6408 (N_6408,N_4781,N_4288);
nor U6409 (N_6409,N_5768,N_5066);
and U6410 (N_6410,N_4527,N_5576);
nor U6411 (N_6411,N_5711,N_4443);
and U6412 (N_6412,N_4311,N_4912);
xnor U6413 (N_6413,N_4538,N_5252);
nor U6414 (N_6414,N_4131,N_5613);
or U6415 (N_6415,N_5612,N_4532);
or U6416 (N_6416,N_4495,N_4324);
or U6417 (N_6417,N_5651,N_5559);
nor U6418 (N_6418,N_5743,N_5654);
nor U6419 (N_6419,N_4977,N_5372);
and U6420 (N_6420,N_4732,N_5866);
or U6421 (N_6421,N_4201,N_4780);
or U6422 (N_6422,N_5884,N_5583);
and U6423 (N_6423,N_4423,N_5238);
nor U6424 (N_6424,N_4336,N_4079);
or U6425 (N_6425,N_4670,N_5587);
xor U6426 (N_6426,N_4675,N_5862);
nand U6427 (N_6427,N_5487,N_5103);
or U6428 (N_6428,N_4523,N_5547);
or U6429 (N_6429,N_4442,N_5501);
nand U6430 (N_6430,N_4747,N_4025);
nand U6431 (N_6431,N_5275,N_4626);
nand U6432 (N_6432,N_5047,N_4381);
or U6433 (N_6433,N_4844,N_4590);
nor U6434 (N_6434,N_4869,N_4096);
nor U6435 (N_6435,N_4566,N_5392);
nand U6436 (N_6436,N_5570,N_4560);
nand U6437 (N_6437,N_5335,N_4189);
nand U6438 (N_6438,N_4164,N_5424);
xnor U6439 (N_6439,N_5499,N_4185);
nand U6440 (N_6440,N_5272,N_5014);
and U6441 (N_6441,N_5707,N_5267);
or U6442 (N_6442,N_5254,N_4669);
xor U6443 (N_6443,N_4712,N_5029);
nand U6444 (N_6444,N_5543,N_4678);
and U6445 (N_6445,N_4182,N_4709);
nand U6446 (N_6446,N_5032,N_4220);
and U6447 (N_6447,N_5975,N_5972);
and U6448 (N_6448,N_5463,N_5836);
nor U6449 (N_6449,N_4689,N_5720);
and U6450 (N_6450,N_4666,N_5120);
nor U6451 (N_6451,N_4302,N_5798);
xnor U6452 (N_6452,N_5737,N_5172);
or U6453 (N_6453,N_4308,N_5808);
nor U6454 (N_6454,N_4719,N_5342);
and U6455 (N_6455,N_4052,N_4221);
and U6456 (N_6456,N_5180,N_4998);
and U6457 (N_6457,N_4029,N_5297);
and U6458 (N_6458,N_4418,N_4801);
and U6459 (N_6459,N_4421,N_4725);
or U6460 (N_6460,N_4570,N_5725);
or U6461 (N_6461,N_4199,N_5920);
nor U6462 (N_6462,N_4102,N_5781);
and U6463 (N_6463,N_5011,N_5715);
xnor U6464 (N_6464,N_4634,N_4744);
nor U6465 (N_6465,N_4390,N_5607);
nor U6466 (N_6466,N_4274,N_5154);
nor U6467 (N_6467,N_4083,N_4493);
nand U6468 (N_6468,N_4380,N_5608);
xnor U6469 (N_6469,N_4550,N_5195);
xnor U6470 (N_6470,N_4376,N_4347);
or U6471 (N_6471,N_5234,N_5354);
or U6472 (N_6472,N_4300,N_5564);
nor U6473 (N_6473,N_4508,N_4730);
xor U6474 (N_6474,N_4821,N_5575);
nor U6475 (N_6475,N_5775,N_4337);
or U6476 (N_6476,N_5389,N_4386);
xor U6477 (N_6477,N_4436,N_5939);
nand U6478 (N_6478,N_5650,N_4579);
nand U6479 (N_6479,N_4591,N_5767);
nor U6480 (N_6480,N_4023,N_5881);
and U6481 (N_6481,N_5948,N_4755);
nand U6482 (N_6482,N_4676,N_4933);
xnor U6483 (N_6483,N_5005,N_5763);
or U6484 (N_6484,N_4779,N_5328);
and U6485 (N_6485,N_5661,N_4192);
and U6486 (N_6486,N_5307,N_4298);
and U6487 (N_6487,N_5548,N_4607);
nor U6488 (N_6488,N_5476,N_5807);
and U6489 (N_6489,N_5309,N_5017);
or U6490 (N_6490,N_5628,N_4401);
nor U6491 (N_6491,N_4937,N_4748);
and U6492 (N_6492,N_5691,N_4226);
xor U6493 (N_6493,N_4344,N_4248);
nand U6494 (N_6494,N_4502,N_5949);
and U6495 (N_6495,N_4010,N_4514);
nand U6496 (N_6496,N_5455,N_5186);
nand U6497 (N_6497,N_5758,N_4893);
or U6498 (N_6498,N_4531,N_4750);
or U6499 (N_6499,N_4346,N_4287);
nor U6500 (N_6500,N_5999,N_4266);
nand U6501 (N_6501,N_5778,N_4270);
nand U6502 (N_6502,N_4372,N_4116);
nand U6503 (N_6503,N_4160,N_5174);
or U6504 (N_6504,N_4557,N_5317);
nand U6505 (N_6505,N_4498,N_4043);
nand U6506 (N_6506,N_4247,N_5015);
nand U6507 (N_6507,N_4541,N_5858);
nor U6508 (N_6508,N_5150,N_5121);
nand U6509 (N_6509,N_4129,N_5835);
and U6510 (N_6510,N_4572,N_5333);
nor U6511 (N_6511,N_4005,N_4378);
xnor U6512 (N_6512,N_5632,N_5086);
or U6513 (N_6513,N_4340,N_5026);
nor U6514 (N_6514,N_5571,N_5352);
or U6515 (N_6515,N_5175,N_5105);
nand U6516 (N_6516,N_5019,N_5699);
or U6517 (N_6517,N_4108,N_4282);
xnor U6518 (N_6518,N_5530,N_4964);
nand U6519 (N_6519,N_4738,N_4580);
and U6520 (N_6520,N_5528,N_5337);
or U6521 (N_6521,N_5591,N_5114);
xnor U6522 (N_6522,N_4454,N_4594);
nor U6523 (N_6523,N_4916,N_4009);
and U6524 (N_6524,N_4874,N_4713);
or U6525 (N_6525,N_4742,N_4313);
or U6526 (N_6526,N_4069,N_5098);
nor U6527 (N_6527,N_4141,N_5306);
nor U6528 (N_6528,N_4293,N_4583);
nand U6529 (N_6529,N_4885,N_5682);
nor U6530 (N_6530,N_5102,N_4342);
nand U6531 (N_6531,N_4360,N_4838);
nor U6532 (N_6532,N_4561,N_5208);
nor U6533 (N_6533,N_5305,N_5263);
xor U6534 (N_6534,N_4884,N_4585);
or U6535 (N_6535,N_4720,N_4904);
or U6536 (N_6536,N_5071,N_5560);
nand U6537 (N_6537,N_4015,N_5128);
xnor U6538 (N_6538,N_4363,N_5024);
or U6539 (N_6539,N_5367,N_5745);
xor U6540 (N_6540,N_4268,N_5890);
nand U6541 (N_6541,N_5133,N_5644);
or U6542 (N_6542,N_4640,N_4166);
nand U6543 (N_6543,N_5586,N_5278);
xnor U6544 (N_6544,N_4051,N_5428);
and U6545 (N_6545,N_5167,N_4076);
and U6546 (N_6546,N_4095,N_5043);
nor U6547 (N_6547,N_4581,N_4913);
and U6548 (N_6548,N_5594,N_4317);
nor U6549 (N_6549,N_4963,N_5579);
or U6550 (N_6550,N_4264,N_5791);
nor U6551 (N_6551,N_5115,N_5976);
nand U6552 (N_6552,N_4410,N_5035);
and U6553 (N_6553,N_5631,N_5166);
and U6554 (N_6554,N_5733,N_4278);
nand U6555 (N_6555,N_4227,N_5918);
and U6556 (N_6556,N_5824,N_4486);
or U6557 (N_6557,N_5527,N_4717);
nor U6558 (N_6558,N_4788,N_4420);
xor U6559 (N_6559,N_4000,N_5534);
and U6560 (N_6560,N_4127,N_4985);
and U6561 (N_6561,N_5578,N_4920);
nand U6562 (N_6562,N_4782,N_4575);
nand U6563 (N_6563,N_5967,N_5818);
nand U6564 (N_6564,N_4022,N_5895);
nor U6565 (N_6565,N_5850,N_4273);
or U6566 (N_6566,N_5960,N_4721);
or U6567 (N_6567,N_5218,N_5652);
and U6568 (N_6568,N_4999,N_5848);
nand U6569 (N_6569,N_4126,N_5772);
or U6570 (N_6570,N_5748,N_5666);
nor U6571 (N_6571,N_4408,N_4643);
or U6572 (N_6572,N_4905,N_5670);
nand U6573 (N_6573,N_5966,N_4513);
nor U6574 (N_6574,N_4252,N_5399);
nor U6575 (N_6575,N_5016,N_5738);
nor U6576 (N_6576,N_4162,N_5995);
or U6577 (N_6577,N_4971,N_4041);
xor U6578 (N_6578,N_5542,N_5036);
nor U6579 (N_6579,N_5897,N_5521);
and U6580 (N_6580,N_5056,N_5787);
and U6581 (N_6581,N_4464,N_5904);
and U6582 (N_6582,N_4504,N_5469);
or U6583 (N_6583,N_5942,N_4321);
nor U6584 (N_6584,N_5675,N_5996);
nand U6585 (N_6585,N_5323,N_5294);
or U6586 (N_6586,N_5984,N_4446);
and U6587 (N_6587,N_4764,N_5407);
or U6588 (N_6588,N_4729,N_5184);
nor U6589 (N_6589,N_5345,N_4740);
and U6590 (N_6590,N_4197,N_4608);
nor U6591 (N_6591,N_4843,N_4600);
and U6592 (N_6592,N_5865,N_4249);
nand U6593 (N_6593,N_4679,N_4193);
and U6594 (N_6594,N_4850,N_5478);
nand U6595 (N_6595,N_5771,N_4961);
xnor U6596 (N_6596,N_5503,N_5627);
and U6597 (N_6597,N_5943,N_5935);
and U6598 (N_6598,N_4056,N_4939);
or U6599 (N_6599,N_4019,N_4435);
xor U6600 (N_6600,N_4229,N_4359);
nand U6601 (N_6601,N_4217,N_5125);
nor U6602 (N_6602,N_4698,N_5134);
and U6603 (N_6603,N_4733,N_4516);
nand U6604 (N_6604,N_5232,N_4256);
or U6605 (N_6605,N_4358,N_5464);
and U6606 (N_6606,N_4562,N_4104);
or U6607 (N_6607,N_5804,N_5080);
and U6608 (N_6608,N_5892,N_5107);
or U6609 (N_6609,N_4026,N_4777);
nor U6610 (N_6610,N_5504,N_4627);
xnor U6611 (N_6611,N_5030,N_5713);
xnor U6612 (N_6612,N_5669,N_4685);
nand U6613 (N_6613,N_5934,N_5341);
and U6614 (N_6614,N_4657,N_5406);
nand U6615 (N_6615,N_4743,N_5295);
nor U6616 (N_6616,N_5496,N_5202);
or U6617 (N_6617,N_5802,N_4962);
nand U6618 (N_6618,N_4459,N_5088);
xnor U6619 (N_6619,N_5188,N_4956);
nand U6620 (N_6620,N_4795,N_5368);
nor U6621 (N_6621,N_5684,N_5574);
or U6622 (N_6622,N_4235,N_4448);
or U6623 (N_6623,N_5974,N_4368);
or U6624 (N_6624,N_5451,N_5653);
and U6625 (N_6625,N_5921,N_4291);
nand U6626 (N_6626,N_5481,N_5600);
nor U6627 (N_6627,N_5536,N_4967);
nand U6628 (N_6628,N_4507,N_4888);
and U6629 (N_6629,N_4936,N_4653);
and U6630 (N_6630,N_5091,N_5290);
nor U6631 (N_6631,N_5761,N_5028);
and U6632 (N_6632,N_5779,N_5535);
nor U6633 (N_6633,N_4451,N_5090);
nand U6634 (N_6634,N_5637,N_4974);
nand U6635 (N_6635,N_4330,N_4382);
nand U6636 (N_6636,N_5021,N_4817);
nor U6637 (N_6637,N_4992,N_5197);
and U6638 (N_6638,N_5844,N_5336);
or U6639 (N_6639,N_5456,N_4949);
or U6640 (N_6640,N_5159,N_4526);
nor U6641 (N_6641,N_5289,N_5673);
nor U6642 (N_6642,N_5364,N_5980);
xnor U6643 (N_6643,N_4384,N_5058);
nor U6644 (N_6644,N_4950,N_5688);
nand U6645 (N_6645,N_4405,N_5110);
nand U6646 (N_6646,N_5614,N_5853);
nand U6647 (N_6647,N_4851,N_5550);
nor U6648 (N_6648,N_5397,N_5994);
nor U6649 (N_6649,N_5799,N_4965);
nand U6650 (N_6650,N_4168,N_4122);
or U6651 (N_6651,N_5217,N_5845);
nand U6652 (N_6652,N_4361,N_5927);
xor U6653 (N_6653,N_4941,N_4638);
and U6654 (N_6654,N_5658,N_4441);
nand U6655 (N_6655,N_4632,N_5751);
nand U6656 (N_6656,N_5057,N_4246);
or U6657 (N_6657,N_4677,N_5040);
nand U6658 (N_6658,N_4128,N_4055);
nand U6659 (N_6659,N_4357,N_5418);
nand U6660 (N_6660,N_4735,N_5326);
and U6661 (N_6661,N_4206,N_4536);
xor U6662 (N_6662,N_5075,N_4595);
nor U6663 (N_6663,N_5299,N_5383);
and U6664 (N_6664,N_4633,N_5231);
and U6665 (N_6665,N_5558,N_4240);
and U6666 (N_6666,N_4805,N_4479);
or U6667 (N_6667,N_5566,N_5329);
nand U6668 (N_6668,N_4100,N_5950);
nor U6669 (N_6669,N_4338,N_4890);
or U6670 (N_6670,N_5054,N_5913);
nand U6671 (N_6671,N_4236,N_5593);
and U6672 (N_6672,N_4921,N_4172);
nand U6673 (N_6673,N_5956,N_4629);
or U6674 (N_6674,N_5403,N_5137);
nand U6675 (N_6675,N_4565,N_4301);
and U6676 (N_6676,N_5288,N_5097);
and U6677 (N_6677,N_4085,N_4659);
nand U6678 (N_6678,N_4333,N_4926);
xnor U6679 (N_6679,N_4663,N_4857);
and U6680 (N_6680,N_5041,N_4331);
nor U6681 (N_6681,N_4613,N_5873);
nand U6682 (N_6682,N_5492,N_5048);
nor U6683 (N_6683,N_4684,N_5262);
nand U6684 (N_6684,N_5812,N_4569);
nor U6685 (N_6685,N_5517,N_5785);
nor U6686 (N_6686,N_5126,N_5744);
nor U6687 (N_6687,N_5703,N_4117);
nand U6688 (N_6688,N_4511,N_4314);
nor U6689 (N_6689,N_5415,N_4106);
nand U6690 (N_6690,N_5340,N_5250);
and U6691 (N_6691,N_5933,N_4031);
and U6692 (N_6692,N_4928,N_4427);
and U6693 (N_6693,N_4563,N_5655);
nor U6694 (N_6694,N_4187,N_4148);
or U6695 (N_6695,N_4259,N_4074);
xor U6696 (N_6696,N_5270,N_5292);
nand U6697 (N_6697,N_5457,N_5382);
nor U6698 (N_6698,N_4655,N_5461);
nor U6699 (N_6699,N_5938,N_5198);
and U6700 (N_6700,N_4332,N_4852);
or U6701 (N_6701,N_5350,N_4822);
or U6702 (N_6702,N_5549,N_5155);
or U6703 (N_6703,N_4243,N_5493);
nor U6704 (N_6704,N_4178,N_4453);
xor U6705 (N_6705,N_4366,N_4951);
nor U6706 (N_6706,N_5419,N_5660);
nand U6707 (N_6707,N_4024,N_5694);
xnor U6708 (N_6708,N_4281,N_4606);
nor U6709 (N_6709,N_4013,N_4286);
or U6710 (N_6710,N_4364,N_4946);
nor U6711 (N_6711,N_4806,N_4456);
nor U6712 (N_6712,N_5343,N_4354);
nand U6713 (N_6713,N_4377,N_5475);
and U6714 (N_6714,N_4808,N_4957);
nor U6715 (N_6715,N_5512,N_5264);
nor U6716 (N_6716,N_4703,N_4231);
and U6717 (N_6717,N_5792,N_5227);
nor U6718 (N_6718,N_4165,N_5917);
and U6719 (N_6719,N_4522,N_4909);
and U6720 (N_6720,N_5480,N_5766);
and U6721 (N_6721,N_4399,N_5119);
or U6722 (N_6722,N_4070,N_5832);
xor U6723 (N_6723,N_4480,N_5319);
and U6724 (N_6724,N_5914,N_4876);
xnor U6725 (N_6725,N_4107,N_4292);
nor U6726 (N_6726,N_4034,N_4478);
xor U6727 (N_6727,N_5427,N_4021);
and U6728 (N_6728,N_5148,N_5076);
nor U6729 (N_6729,N_4492,N_4855);
nor U6730 (N_6730,N_5300,N_5228);
and U6731 (N_6731,N_5700,N_5436);
xor U6732 (N_6732,N_4003,N_5852);
or U6733 (N_6733,N_5431,N_5562);
and U6734 (N_6734,N_5007,N_4894);
and U6735 (N_6735,N_5158,N_5386);
or U6736 (N_6736,N_4373,N_5602);
or U6737 (N_6737,N_4810,N_5233);
and U6738 (N_6738,N_4225,N_4306);
xor U6739 (N_6739,N_4094,N_5656);
nand U6740 (N_6740,N_4133,N_5876);
xor U6741 (N_6741,N_4895,N_5413);
or U6742 (N_6742,N_5338,N_4048);
nor U6743 (N_6743,N_5414,N_5471);
nor U6744 (N_6744,N_4012,N_5908);
nand U6745 (N_6745,N_5981,N_5616);
and U6746 (N_6746,N_4891,N_4533);
and U6747 (N_6747,N_4455,N_4253);
nor U6748 (N_6748,N_4879,N_5732);
nor U6749 (N_6749,N_4952,N_5678);
and U6750 (N_6750,N_5241,N_4804);
or U6751 (N_6751,N_5077,N_5129);
nand U6752 (N_6752,N_4245,N_4263);
and U6753 (N_6753,N_4494,N_5997);
nand U6754 (N_6754,N_4605,N_4409);
xor U6755 (N_6755,N_5216,N_4383);
or U6756 (N_6756,N_5573,N_4318);
xnor U6757 (N_6757,N_4539,N_5452);
nor U6758 (N_6758,N_5483,N_4959);
nor U6759 (N_6759,N_5243,N_5312);
xnor U6760 (N_6760,N_4996,N_5360);
nand U6761 (N_6761,N_4968,N_5401);
nor U6762 (N_6762,N_5268,N_5344);
nor U6763 (N_6763,N_4889,N_5510);
or U6764 (N_6764,N_5679,N_4586);
or U6765 (N_6765,N_5615,N_5879);
nand U6766 (N_6766,N_4710,N_5353);
nand U6767 (N_6767,N_5645,N_4661);
nor U6768 (N_6768,N_5050,N_4058);
nand U6769 (N_6769,N_4284,N_4763);
and U6770 (N_6770,N_5222,N_4151);
nor U6771 (N_6771,N_4695,N_5827);
nand U6772 (N_6772,N_5065,N_4624);
nor U6773 (N_6773,N_4482,N_4045);
nor U6774 (N_6774,N_5279,N_4190);
nand U6775 (N_6775,N_4966,N_5334);
nand U6776 (N_6776,N_5729,N_4693);
nand U6777 (N_6777,N_4680,N_4320);
and U6778 (N_6778,N_5139,N_4623);
and U6779 (N_6779,N_5696,N_5206);
nand U6780 (N_6780,N_4099,N_5301);
nand U6781 (N_6781,N_5220,N_5164);
and U6782 (N_6782,N_4656,N_5683);
xnor U6783 (N_6783,N_4295,N_4672);
nand U6784 (N_6784,N_4797,N_5760);
nand U6785 (N_6785,N_4519,N_5303);
or U6786 (N_6786,N_5532,N_5648);
or U6787 (N_6787,N_5376,N_5031);
and U6788 (N_6788,N_4835,N_4438);
nor U6789 (N_6789,N_4731,N_5448);
or U6790 (N_6790,N_5854,N_4272);
and U6791 (N_6791,N_5346,N_5511);
or U6792 (N_6792,N_4413,N_5821);
nor U6793 (N_6793,N_4818,N_4545);
nor U6794 (N_6794,N_5916,N_4994);
and U6795 (N_6795,N_4820,N_5465);
or U6796 (N_6796,N_5951,N_4866);
nor U6797 (N_6797,N_4784,N_5449);
xor U6798 (N_6798,N_4167,N_5867);
nand U6799 (N_6799,N_5145,N_5947);
or U6800 (N_6800,N_4988,N_5959);
nor U6801 (N_6801,N_4537,N_4785);
or U6802 (N_6802,N_4631,N_4824);
xor U6803 (N_6803,N_4388,N_5236);
or U6804 (N_6804,N_5871,N_4228);
or U6805 (N_6805,N_5192,N_4665);
and U6806 (N_6806,N_4276,N_5565);
and U6807 (N_6807,N_5701,N_5896);
and U6808 (N_6808,N_5069,N_4466);
and U6809 (N_6809,N_5111,N_4279);
xor U6810 (N_6810,N_5314,N_5000);
nor U6811 (N_6811,N_4871,N_5882);
or U6812 (N_6812,N_4814,N_4671);
and U6813 (N_6813,N_5931,N_4958);
nor U6814 (N_6814,N_5717,N_4241);
xor U6815 (N_6815,N_4970,N_4071);
nand U6816 (N_6816,N_4196,N_5127);
or U6817 (N_6817,N_4794,N_5983);
or U6818 (N_6818,N_4371,N_4636);
xnor U6819 (N_6819,N_4143,N_5117);
xor U6820 (N_6820,N_4768,N_5705);
or U6821 (N_6821,N_5954,N_5636);
and U6822 (N_6822,N_4839,N_4230);
and U6823 (N_6823,N_5851,N_4078);
and U6824 (N_6824,N_5618,N_4972);
nand U6825 (N_6825,N_4063,N_4138);
and U6826 (N_6826,N_4762,N_5941);
nand U6827 (N_6827,N_4208,N_5764);
nand U6828 (N_6828,N_4303,N_4940);
and U6829 (N_6829,N_5211,N_5212);
xor U6830 (N_6830,N_5349,N_4798);
and U6831 (N_6831,N_5422,N_5721);
or U6832 (N_6832,N_4269,N_5287);
nor U6833 (N_6833,N_5157,N_4518);
or U6834 (N_6834,N_5875,N_4398);
nor U6835 (N_6835,N_5109,N_4216);
or U6836 (N_6836,N_4432,N_4232);
or U6837 (N_6837,N_4915,N_4793);
or U6838 (N_6838,N_5348,N_5809);
and U6839 (N_6839,N_4412,N_5716);
or U6840 (N_6840,N_5039,N_4163);
nand U6841 (N_6841,N_5417,N_5697);
nand U6842 (N_6842,N_4396,N_4452);
or U6843 (N_6843,N_5830,N_5513);
nor U6844 (N_6844,N_5140,N_4945);
or U6845 (N_6845,N_4257,N_5859);
or U6846 (N_6846,N_5937,N_5929);
and U6847 (N_6847,N_5676,N_4036);
or U6848 (N_6848,N_4233,N_4642);
or U6849 (N_6849,N_4176,N_4597);
nor U6850 (N_6850,N_4407,N_4238);
nor U6851 (N_6851,N_5776,N_4749);
and U6852 (N_6852,N_4437,N_5194);
nand U6853 (N_6853,N_5484,N_5324);
or U6854 (N_6854,N_4900,N_5142);
nor U6855 (N_6855,N_5601,N_4461);
and U6856 (N_6856,N_4395,N_5629);
or U6857 (N_6857,N_5664,N_5605);
nand U6858 (N_6858,N_4592,N_4121);
nand U6859 (N_6859,N_5936,N_5138);
nand U6860 (N_6860,N_5149,N_4901);
nor U6861 (N_6861,N_4736,N_4686);
xor U6862 (N_6862,N_5714,N_4568);
and U6863 (N_6863,N_5680,N_4329);
and U6864 (N_6864,N_4847,N_4829);
nand U6865 (N_6865,N_4886,N_5634);
nand U6866 (N_6866,N_4925,N_5643);
or U6867 (N_6867,N_4811,N_4244);
nand U6868 (N_6868,N_4207,N_5907);
and U6869 (N_6869,N_5633,N_5060);
nand U6870 (N_6870,N_5308,N_4305);
and U6871 (N_6871,N_5945,N_4816);
or U6872 (N_6872,N_5257,N_4375);
nor U6873 (N_6873,N_4548,N_5472);
nand U6874 (N_6874,N_5434,N_4174);
nor U6875 (N_6875,N_5313,N_5321);
nand U6876 (N_6876,N_5485,N_4761);
nor U6877 (N_6877,N_5380,N_4506);
nand U6878 (N_6878,N_4046,N_4625);
nor U6879 (N_6879,N_5665,N_5096);
nand U6880 (N_6880,N_4696,N_4734);
nor U6881 (N_6881,N_5529,N_5327);
nand U6882 (N_6882,N_5193,N_4528);
and U6883 (N_6883,N_5087,N_4429);
or U6884 (N_6884,N_4072,N_5094);
xnor U6885 (N_6885,N_5915,N_5777);
and U6886 (N_6886,N_4549,N_4447);
or U6887 (N_6887,N_5224,N_5460);
nor U6888 (N_6888,N_4796,N_5421);
nor U6889 (N_6889,N_4819,N_5161);
nor U6890 (N_6890,N_5500,N_4978);
nand U6891 (N_6891,N_5971,N_4943);
or U6892 (N_6892,N_5523,N_5365);
or U6893 (N_6893,N_4473,N_4218);
nor U6894 (N_6894,N_5834,N_4501);
nand U6895 (N_6895,N_5869,N_4746);
or U6896 (N_6896,N_5473,N_4490);
or U6897 (N_6897,N_5797,N_4564);
or U6898 (N_6898,N_5394,N_5370);
nor U6899 (N_6899,N_5200,N_4792);
or U6900 (N_6900,N_5782,N_4038);
nand U6901 (N_6901,N_5856,N_4140);
and U6902 (N_6902,N_5833,N_5706);
or U6903 (N_6903,N_5784,N_4499);
nor U6904 (N_6904,N_4047,N_5255);
or U6905 (N_6905,N_5773,N_4674);
nor U6906 (N_6906,N_5454,N_5898);
or U6907 (N_6907,N_5265,N_5979);
nand U6908 (N_6908,N_5409,N_4883);
or U6909 (N_6909,N_5590,N_4799);
nor U6910 (N_6910,N_5067,N_4416);
nand U6911 (N_6911,N_5520,N_4262);
and U6912 (N_6912,N_5388,N_5822);
or U6913 (N_6913,N_5746,N_5256);
and U6914 (N_6914,N_5153,N_5739);
nand U6915 (N_6915,N_4858,N_4153);
xor U6916 (N_6916,N_5269,N_5331);
or U6917 (N_6917,N_5533,N_4369);
and U6918 (N_6918,N_5240,N_4524);
and U6919 (N_6919,N_4011,N_5400);
nor U6920 (N_6920,N_5235,N_5516);
nor U6921 (N_6921,N_4953,N_4488);
or U6922 (N_6922,N_4969,N_4701);
nand U6923 (N_6923,N_4445,N_5617);
nand U6924 (N_6924,N_4267,N_4825);
nand U6925 (N_6925,N_4352,N_4995);
nand U6926 (N_6926,N_4135,N_4091);
or U6927 (N_6927,N_4727,N_5710);
or U6928 (N_6928,N_4348,N_5237);
nor U6929 (N_6929,N_5728,N_5749);
and U6930 (N_6930,N_5037,N_4483);
nor U6931 (N_6931,N_5568,N_4910);
xor U6932 (N_6932,N_4530,N_4181);
nand U6933 (N_6933,N_4035,N_4914);
and U6934 (N_6934,N_4854,N_4612);
nand U6935 (N_6935,N_4061,N_4175);
and U6936 (N_6936,N_5025,N_4171);
nand U6937 (N_6937,N_5978,N_4309);
and U6938 (N_6938,N_5378,N_5657);
xnor U6939 (N_6939,N_4849,N_5872);
or U6940 (N_6940,N_4582,N_5089);
or U6941 (N_6941,N_5152,N_5122);
and U6942 (N_6942,N_5889,N_4947);
or U6943 (N_6943,N_5823,N_5242);
and U6944 (N_6944,N_4173,N_5495);
nand U6945 (N_6945,N_4726,N_4016);
and U6946 (N_6946,N_4213,N_4387);
nor U6947 (N_6947,N_4159,N_4209);
nand U6948 (N_6948,N_5803,N_5156);
or U6949 (N_6949,N_5838,N_5719);
or U6950 (N_6950,N_5467,N_5261);
or U6951 (N_6951,N_4802,N_5546);
nand U6952 (N_6952,N_4724,N_5642);
nor U6953 (N_6953,N_4353,N_5515);
nor U6954 (N_6954,N_5298,N_4760);
nor U6955 (N_6955,N_4567,N_4198);
nand U6956 (N_6956,N_4080,N_5474);
and U6957 (N_6957,N_4938,N_5925);
or U6958 (N_6958,N_5012,N_4487);
nor U6959 (N_6959,N_5704,N_4077);
nor U6960 (N_6960,N_5042,N_4120);
and U6961 (N_6961,N_4203,N_4831);
nand U6962 (N_6962,N_4588,N_4098);
nor U6963 (N_6963,N_5426,N_4864);
or U6964 (N_6964,N_5540,N_5179);
nor U6965 (N_6965,N_5059,N_5912);
nand U6966 (N_6966,N_4593,N_5588);
and U6967 (N_6967,N_4434,N_4082);
and U6968 (N_6968,N_4991,N_5291);
or U6969 (N_6969,N_4828,N_4474);
nor U6970 (N_6970,N_4426,N_5442);
nor U6971 (N_6971,N_5990,N_4983);
xor U6972 (N_6972,N_4081,N_4787);
or U6973 (N_6973,N_5398,N_5961);
and U6974 (N_6974,N_5522,N_5165);
nand U6975 (N_6975,N_5170,N_4775);
or U6976 (N_6976,N_4497,N_4842);
nor U6977 (N_6977,N_5677,N_4754);
or U6978 (N_6978,N_5062,N_5143);
and U6979 (N_6979,N_4237,N_4621);
nor U6980 (N_6980,N_4759,N_5477);
and U6981 (N_6981,N_4280,N_4027);
or U6982 (N_6982,N_5006,N_5304);
and U6983 (N_6983,N_4897,N_4535);
or U6984 (N_6984,N_5841,N_5444);
or U6985 (N_6985,N_4896,N_5698);
or U6986 (N_6986,N_4283,N_5408);
nand U6987 (N_6987,N_4440,N_5765);
or U6988 (N_6988,N_5357,N_4823);
or U6989 (N_6989,N_4774,N_4555);
or U6990 (N_6990,N_4414,N_4477);
nand U6991 (N_6991,N_5246,N_5373);
nand U6992 (N_6992,N_5187,N_5893);
or U6993 (N_6993,N_4863,N_5734);
nand U6994 (N_6994,N_4242,N_4032);
nor U6995 (N_6995,N_4786,N_5082);
nor U6996 (N_6996,N_5018,N_5332);
or U6997 (N_6997,N_4577,N_5955);
and U6998 (N_6998,N_5280,N_4156);
xor U6999 (N_6999,N_5033,N_4319);
nand U7000 (N_7000,N_4442,N_4441);
and U7001 (N_7001,N_4176,N_4663);
nand U7002 (N_7002,N_5876,N_5938);
xor U7003 (N_7003,N_5598,N_4211);
and U7004 (N_7004,N_5756,N_4168);
nand U7005 (N_7005,N_5108,N_4490);
nor U7006 (N_7006,N_4130,N_5912);
or U7007 (N_7007,N_5612,N_5961);
nand U7008 (N_7008,N_4694,N_5570);
and U7009 (N_7009,N_4813,N_4431);
and U7010 (N_7010,N_5560,N_5323);
and U7011 (N_7011,N_5159,N_4158);
xnor U7012 (N_7012,N_5802,N_4290);
nor U7013 (N_7013,N_4840,N_5293);
or U7014 (N_7014,N_4491,N_4860);
or U7015 (N_7015,N_4473,N_4897);
nor U7016 (N_7016,N_4420,N_5369);
nor U7017 (N_7017,N_5886,N_4637);
nand U7018 (N_7018,N_5156,N_5678);
nand U7019 (N_7019,N_4955,N_5160);
nand U7020 (N_7020,N_4019,N_5064);
and U7021 (N_7021,N_5095,N_4677);
and U7022 (N_7022,N_4108,N_4508);
nor U7023 (N_7023,N_4845,N_5298);
nand U7024 (N_7024,N_4766,N_4662);
nor U7025 (N_7025,N_5688,N_4140);
nor U7026 (N_7026,N_4975,N_5097);
or U7027 (N_7027,N_5985,N_4445);
xor U7028 (N_7028,N_4282,N_4816);
or U7029 (N_7029,N_4340,N_4446);
nand U7030 (N_7030,N_5638,N_4965);
nand U7031 (N_7031,N_5682,N_4656);
nor U7032 (N_7032,N_4405,N_4839);
or U7033 (N_7033,N_5521,N_4551);
or U7034 (N_7034,N_4286,N_5121);
nand U7035 (N_7035,N_5875,N_4327);
nor U7036 (N_7036,N_5409,N_5253);
or U7037 (N_7037,N_4738,N_5008);
or U7038 (N_7038,N_4150,N_4355);
nand U7039 (N_7039,N_5716,N_5653);
nor U7040 (N_7040,N_4600,N_4102);
xnor U7041 (N_7041,N_4557,N_5916);
nand U7042 (N_7042,N_4483,N_4195);
nand U7043 (N_7043,N_5929,N_4945);
nor U7044 (N_7044,N_5849,N_4761);
nor U7045 (N_7045,N_4265,N_4130);
and U7046 (N_7046,N_4752,N_5693);
nor U7047 (N_7047,N_4298,N_5429);
nand U7048 (N_7048,N_4392,N_4619);
or U7049 (N_7049,N_4568,N_4151);
nor U7050 (N_7050,N_5049,N_5339);
or U7051 (N_7051,N_5358,N_4732);
nor U7052 (N_7052,N_4775,N_4466);
nor U7053 (N_7053,N_5083,N_5033);
or U7054 (N_7054,N_5188,N_5962);
and U7055 (N_7055,N_4140,N_5580);
nand U7056 (N_7056,N_5555,N_4580);
and U7057 (N_7057,N_4430,N_5154);
or U7058 (N_7058,N_4418,N_4678);
and U7059 (N_7059,N_4775,N_5902);
and U7060 (N_7060,N_4576,N_5781);
nor U7061 (N_7061,N_5485,N_4837);
nor U7062 (N_7062,N_4955,N_5166);
or U7063 (N_7063,N_5269,N_4982);
xnor U7064 (N_7064,N_4113,N_5499);
nor U7065 (N_7065,N_4583,N_4167);
or U7066 (N_7066,N_5617,N_5932);
nor U7067 (N_7067,N_4360,N_4897);
nand U7068 (N_7068,N_4858,N_4238);
nand U7069 (N_7069,N_5091,N_5183);
nor U7070 (N_7070,N_4406,N_5982);
xnor U7071 (N_7071,N_4949,N_5860);
nor U7072 (N_7072,N_5137,N_5110);
and U7073 (N_7073,N_4718,N_5641);
or U7074 (N_7074,N_4146,N_5281);
nand U7075 (N_7075,N_5532,N_4344);
nand U7076 (N_7076,N_4481,N_5265);
nor U7077 (N_7077,N_5327,N_5230);
nand U7078 (N_7078,N_4514,N_5509);
or U7079 (N_7079,N_5347,N_5570);
or U7080 (N_7080,N_4733,N_5177);
nand U7081 (N_7081,N_5699,N_4340);
nand U7082 (N_7082,N_4918,N_4499);
or U7083 (N_7083,N_4596,N_5330);
and U7084 (N_7084,N_4216,N_4380);
nand U7085 (N_7085,N_4005,N_5332);
and U7086 (N_7086,N_5179,N_4491);
xor U7087 (N_7087,N_4466,N_5888);
and U7088 (N_7088,N_5076,N_5006);
and U7089 (N_7089,N_5268,N_4009);
nand U7090 (N_7090,N_4270,N_4716);
nor U7091 (N_7091,N_5411,N_4522);
or U7092 (N_7092,N_4437,N_4865);
nand U7093 (N_7093,N_5408,N_4860);
or U7094 (N_7094,N_5653,N_4838);
nand U7095 (N_7095,N_4213,N_4551);
or U7096 (N_7096,N_4027,N_4278);
and U7097 (N_7097,N_5771,N_4189);
and U7098 (N_7098,N_4357,N_4422);
nand U7099 (N_7099,N_5888,N_4115);
or U7100 (N_7100,N_4253,N_5650);
or U7101 (N_7101,N_5368,N_5349);
nor U7102 (N_7102,N_4768,N_5606);
nand U7103 (N_7103,N_5974,N_4312);
or U7104 (N_7104,N_5117,N_4631);
nand U7105 (N_7105,N_4785,N_4944);
and U7106 (N_7106,N_5880,N_4865);
nor U7107 (N_7107,N_4924,N_4781);
or U7108 (N_7108,N_5083,N_5437);
and U7109 (N_7109,N_4822,N_4981);
nand U7110 (N_7110,N_4995,N_4294);
and U7111 (N_7111,N_4822,N_5830);
or U7112 (N_7112,N_5441,N_5991);
or U7113 (N_7113,N_4796,N_5146);
nor U7114 (N_7114,N_4493,N_5993);
or U7115 (N_7115,N_4736,N_5045);
or U7116 (N_7116,N_5528,N_4510);
nor U7117 (N_7117,N_5340,N_5473);
nand U7118 (N_7118,N_5424,N_5407);
nor U7119 (N_7119,N_4269,N_4968);
nor U7120 (N_7120,N_5577,N_4727);
and U7121 (N_7121,N_4318,N_4618);
or U7122 (N_7122,N_5680,N_5717);
nor U7123 (N_7123,N_5603,N_4778);
or U7124 (N_7124,N_4557,N_4106);
and U7125 (N_7125,N_5824,N_5216);
and U7126 (N_7126,N_5475,N_4753);
nand U7127 (N_7127,N_4905,N_4024);
and U7128 (N_7128,N_5300,N_5996);
or U7129 (N_7129,N_5191,N_5559);
xor U7130 (N_7130,N_5369,N_5421);
nor U7131 (N_7131,N_5007,N_4810);
nor U7132 (N_7132,N_5698,N_5422);
and U7133 (N_7133,N_5273,N_5606);
and U7134 (N_7134,N_5130,N_4818);
and U7135 (N_7135,N_4768,N_5700);
xnor U7136 (N_7136,N_5824,N_5779);
nand U7137 (N_7137,N_5177,N_4192);
nand U7138 (N_7138,N_5680,N_5642);
nor U7139 (N_7139,N_5324,N_5365);
nor U7140 (N_7140,N_5290,N_5112);
and U7141 (N_7141,N_5030,N_5903);
nand U7142 (N_7142,N_4163,N_5997);
nand U7143 (N_7143,N_5399,N_4037);
and U7144 (N_7144,N_5785,N_5023);
nand U7145 (N_7145,N_5042,N_4229);
nor U7146 (N_7146,N_5151,N_5063);
and U7147 (N_7147,N_4727,N_5333);
xor U7148 (N_7148,N_5414,N_5985);
and U7149 (N_7149,N_4471,N_5146);
nor U7150 (N_7150,N_5244,N_4343);
xor U7151 (N_7151,N_4421,N_4269);
nand U7152 (N_7152,N_4283,N_5897);
or U7153 (N_7153,N_5749,N_4986);
nand U7154 (N_7154,N_4796,N_5723);
nand U7155 (N_7155,N_5359,N_5363);
or U7156 (N_7156,N_4223,N_4005);
nand U7157 (N_7157,N_4481,N_4402);
or U7158 (N_7158,N_4734,N_5624);
nand U7159 (N_7159,N_4788,N_5700);
or U7160 (N_7160,N_4923,N_5247);
nand U7161 (N_7161,N_5434,N_4410);
or U7162 (N_7162,N_4276,N_5062);
and U7163 (N_7163,N_5467,N_4277);
or U7164 (N_7164,N_4625,N_5094);
and U7165 (N_7165,N_5053,N_5058);
nand U7166 (N_7166,N_4303,N_4027);
nand U7167 (N_7167,N_4963,N_4592);
xor U7168 (N_7168,N_5753,N_4767);
nor U7169 (N_7169,N_5914,N_4977);
xnor U7170 (N_7170,N_4361,N_5072);
nor U7171 (N_7171,N_5628,N_4382);
nor U7172 (N_7172,N_5781,N_4617);
or U7173 (N_7173,N_4278,N_4962);
nor U7174 (N_7174,N_4736,N_5735);
and U7175 (N_7175,N_4640,N_5947);
or U7176 (N_7176,N_4635,N_5390);
or U7177 (N_7177,N_5721,N_4154);
or U7178 (N_7178,N_5812,N_4520);
and U7179 (N_7179,N_4540,N_5625);
and U7180 (N_7180,N_5995,N_4427);
nor U7181 (N_7181,N_5259,N_4123);
xor U7182 (N_7182,N_5180,N_5137);
and U7183 (N_7183,N_5952,N_4685);
nand U7184 (N_7184,N_5154,N_5456);
nand U7185 (N_7185,N_4505,N_5647);
and U7186 (N_7186,N_5041,N_5478);
nor U7187 (N_7187,N_4631,N_5525);
or U7188 (N_7188,N_4154,N_5346);
nand U7189 (N_7189,N_5893,N_4198);
nand U7190 (N_7190,N_4328,N_4582);
nor U7191 (N_7191,N_4780,N_5456);
or U7192 (N_7192,N_4331,N_4563);
or U7193 (N_7193,N_4357,N_5717);
nor U7194 (N_7194,N_5704,N_4015);
nand U7195 (N_7195,N_4864,N_4620);
nor U7196 (N_7196,N_4934,N_4692);
and U7197 (N_7197,N_4414,N_4248);
nand U7198 (N_7198,N_4160,N_4919);
and U7199 (N_7199,N_4954,N_5096);
or U7200 (N_7200,N_4661,N_5979);
and U7201 (N_7201,N_5272,N_4129);
nand U7202 (N_7202,N_5772,N_4303);
nand U7203 (N_7203,N_4389,N_5713);
or U7204 (N_7204,N_4894,N_5956);
and U7205 (N_7205,N_5605,N_5653);
and U7206 (N_7206,N_5181,N_5824);
and U7207 (N_7207,N_4023,N_4330);
or U7208 (N_7208,N_5185,N_5193);
nor U7209 (N_7209,N_4305,N_4858);
xor U7210 (N_7210,N_4291,N_4327);
or U7211 (N_7211,N_4693,N_5437);
or U7212 (N_7212,N_5598,N_4987);
xor U7213 (N_7213,N_5991,N_4883);
or U7214 (N_7214,N_4256,N_4391);
nand U7215 (N_7215,N_5841,N_4678);
or U7216 (N_7216,N_5663,N_5606);
nor U7217 (N_7217,N_4860,N_5006);
nand U7218 (N_7218,N_5645,N_5509);
and U7219 (N_7219,N_5332,N_5319);
nand U7220 (N_7220,N_5649,N_4998);
xnor U7221 (N_7221,N_5945,N_5246);
nor U7222 (N_7222,N_4472,N_5852);
or U7223 (N_7223,N_4818,N_5289);
nand U7224 (N_7224,N_5398,N_4231);
nor U7225 (N_7225,N_4499,N_5030);
nand U7226 (N_7226,N_4668,N_4773);
nor U7227 (N_7227,N_4796,N_4959);
and U7228 (N_7228,N_5259,N_4782);
or U7229 (N_7229,N_5332,N_4554);
nand U7230 (N_7230,N_5081,N_4590);
or U7231 (N_7231,N_4663,N_4490);
or U7232 (N_7232,N_4135,N_4841);
and U7233 (N_7233,N_4162,N_5053);
nand U7234 (N_7234,N_5372,N_5455);
nand U7235 (N_7235,N_5771,N_5369);
and U7236 (N_7236,N_5388,N_4556);
nor U7237 (N_7237,N_5383,N_5104);
or U7238 (N_7238,N_4410,N_5987);
or U7239 (N_7239,N_5967,N_5701);
or U7240 (N_7240,N_4960,N_5478);
nand U7241 (N_7241,N_4162,N_4640);
nand U7242 (N_7242,N_4162,N_4051);
or U7243 (N_7243,N_4291,N_4685);
or U7244 (N_7244,N_5901,N_4455);
and U7245 (N_7245,N_4991,N_4796);
nand U7246 (N_7246,N_5721,N_5598);
nand U7247 (N_7247,N_5415,N_5851);
or U7248 (N_7248,N_4470,N_5544);
or U7249 (N_7249,N_5192,N_4684);
and U7250 (N_7250,N_4042,N_5788);
nand U7251 (N_7251,N_4204,N_5298);
and U7252 (N_7252,N_5732,N_4972);
nand U7253 (N_7253,N_5786,N_4300);
or U7254 (N_7254,N_4887,N_5079);
and U7255 (N_7255,N_4171,N_5897);
and U7256 (N_7256,N_4092,N_5944);
and U7257 (N_7257,N_5685,N_5041);
or U7258 (N_7258,N_4337,N_5885);
nand U7259 (N_7259,N_4416,N_4678);
xnor U7260 (N_7260,N_4155,N_4260);
or U7261 (N_7261,N_5985,N_5120);
and U7262 (N_7262,N_5242,N_5373);
or U7263 (N_7263,N_4054,N_4466);
or U7264 (N_7264,N_4828,N_4640);
or U7265 (N_7265,N_4271,N_5870);
xor U7266 (N_7266,N_4712,N_5013);
nor U7267 (N_7267,N_5852,N_5869);
nor U7268 (N_7268,N_4005,N_5645);
and U7269 (N_7269,N_5311,N_5643);
nor U7270 (N_7270,N_4085,N_4806);
nor U7271 (N_7271,N_5064,N_5488);
and U7272 (N_7272,N_5947,N_4928);
nand U7273 (N_7273,N_4555,N_4749);
or U7274 (N_7274,N_5802,N_5787);
or U7275 (N_7275,N_4838,N_5030);
and U7276 (N_7276,N_4248,N_4666);
xnor U7277 (N_7277,N_5580,N_4757);
or U7278 (N_7278,N_4888,N_4618);
and U7279 (N_7279,N_5275,N_5097);
and U7280 (N_7280,N_4925,N_4734);
or U7281 (N_7281,N_5187,N_4914);
nand U7282 (N_7282,N_5644,N_5729);
or U7283 (N_7283,N_4345,N_4206);
nor U7284 (N_7284,N_4069,N_4536);
nor U7285 (N_7285,N_5911,N_5812);
xnor U7286 (N_7286,N_5569,N_4852);
and U7287 (N_7287,N_5292,N_5869);
and U7288 (N_7288,N_4476,N_5529);
nand U7289 (N_7289,N_4918,N_5864);
or U7290 (N_7290,N_5916,N_4621);
xor U7291 (N_7291,N_4218,N_4506);
nand U7292 (N_7292,N_4734,N_4675);
and U7293 (N_7293,N_4985,N_4196);
or U7294 (N_7294,N_4102,N_5152);
or U7295 (N_7295,N_5429,N_5441);
or U7296 (N_7296,N_5054,N_5251);
nand U7297 (N_7297,N_4194,N_4284);
nor U7298 (N_7298,N_4654,N_5636);
nand U7299 (N_7299,N_5771,N_5201);
xnor U7300 (N_7300,N_5696,N_4138);
and U7301 (N_7301,N_5871,N_5532);
nor U7302 (N_7302,N_5326,N_4561);
or U7303 (N_7303,N_5027,N_4904);
nor U7304 (N_7304,N_4690,N_4631);
or U7305 (N_7305,N_5605,N_4828);
xor U7306 (N_7306,N_5033,N_4426);
nand U7307 (N_7307,N_5785,N_5584);
nor U7308 (N_7308,N_4192,N_5729);
nand U7309 (N_7309,N_4727,N_5668);
nor U7310 (N_7310,N_5628,N_5647);
or U7311 (N_7311,N_5065,N_5001);
nand U7312 (N_7312,N_5752,N_4514);
and U7313 (N_7313,N_5309,N_5077);
and U7314 (N_7314,N_4448,N_4854);
nor U7315 (N_7315,N_4253,N_5965);
nand U7316 (N_7316,N_5412,N_5636);
nand U7317 (N_7317,N_4233,N_5168);
or U7318 (N_7318,N_5259,N_5517);
nor U7319 (N_7319,N_4935,N_5475);
or U7320 (N_7320,N_5430,N_4164);
xnor U7321 (N_7321,N_5441,N_5355);
or U7322 (N_7322,N_4758,N_4056);
and U7323 (N_7323,N_5957,N_5289);
and U7324 (N_7324,N_4538,N_5905);
nand U7325 (N_7325,N_5222,N_5256);
nor U7326 (N_7326,N_5290,N_4770);
or U7327 (N_7327,N_5893,N_5307);
xor U7328 (N_7328,N_5036,N_4092);
or U7329 (N_7329,N_4097,N_4469);
or U7330 (N_7330,N_5792,N_4668);
or U7331 (N_7331,N_4013,N_4505);
and U7332 (N_7332,N_5563,N_4951);
and U7333 (N_7333,N_4464,N_4663);
or U7334 (N_7334,N_4188,N_5604);
nor U7335 (N_7335,N_4619,N_5509);
and U7336 (N_7336,N_4930,N_4072);
and U7337 (N_7337,N_5074,N_4099);
or U7338 (N_7338,N_5351,N_5029);
nor U7339 (N_7339,N_5172,N_5365);
or U7340 (N_7340,N_5042,N_4441);
and U7341 (N_7341,N_5587,N_5235);
and U7342 (N_7342,N_5065,N_5761);
nand U7343 (N_7343,N_4019,N_4088);
or U7344 (N_7344,N_5267,N_5787);
or U7345 (N_7345,N_5657,N_4197);
and U7346 (N_7346,N_5830,N_5721);
or U7347 (N_7347,N_5238,N_4707);
nand U7348 (N_7348,N_4129,N_5130);
nand U7349 (N_7349,N_5802,N_4493);
and U7350 (N_7350,N_5125,N_4859);
or U7351 (N_7351,N_4281,N_5332);
nand U7352 (N_7352,N_5188,N_5643);
or U7353 (N_7353,N_4802,N_4256);
and U7354 (N_7354,N_5034,N_5520);
or U7355 (N_7355,N_4624,N_5986);
nor U7356 (N_7356,N_5619,N_5539);
and U7357 (N_7357,N_4033,N_4524);
nand U7358 (N_7358,N_4795,N_4916);
and U7359 (N_7359,N_5603,N_5234);
nor U7360 (N_7360,N_4130,N_5503);
and U7361 (N_7361,N_4677,N_4927);
and U7362 (N_7362,N_5470,N_5305);
nor U7363 (N_7363,N_5095,N_5604);
nand U7364 (N_7364,N_5854,N_4479);
and U7365 (N_7365,N_5243,N_4310);
nand U7366 (N_7366,N_4581,N_4796);
nor U7367 (N_7367,N_4935,N_4567);
or U7368 (N_7368,N_4430,N_4099);
nand U7369 (N_7369,N_5957,N_4088);
or U7370 (N_7370,N_5832,N_5743);
and U7371 (N_7371,N_5025,N_4494);
nand U7372 (N_7372,N_4471,N_4987);
or U7373 (N_7373,N_4384,N_5815);
or U7374 (N_7374,N_5656,N_5015);
or U7375 (N_7375,N_4392,N_5612);
and U7376 (N_7376,N_5555,N_5527);
or U7377 (N_7377,N_4919,N_4052);
and U7378 (N_7378,N_4642,N_4164);
or U7379 (N_7379,N_4598,N_4346);
nand U7380 (N_7380,N_5319,N_4596);
nor U7381 (N_7381,N_4024,N_5898);
or U7382 (N_7382,N_4169,N_5108);
and U7383 (N_7383,N_4332,N_4892);
and U7384 (N_7384,N_5999,N_5297);
nand U7385 (N_7385,N_5630,N_5315);
nor U7386 (N_7386,N_4590,N_5712);
or U7387 (N_7387,N_5656,N_4699);
nand U7388 (N_7388,N_4877,N_4449);
xnor U7389 (N_7389,N_4574,N_4705);
nor U7390 (N_7390,N_5476,N_4051);
nor U7391 (N_7391,N_4566,N_4925);
and U7392 (N_7392,N_5613,N_4017);
nor U7393 (N_7393,N_5685,N_4025);
and U7394 (N_7394,N_4541,N_4493);
and U7395 (N_7395,N_4393,N_4537);
nand U7396 (N_7396,N_4668,N_4099);
or U7397 (N_7397,N_5420,N_4653);
xnor U7398 (N_7398,N_5891,N_5322);
or U7399 (N_7399,N_4542,N_4367);
and U7400 (N_7400,N_4460,N_4760);
xnor U7401 (N_7401,N_5976,N_5273);
and U7402 (N_7402,N_5023,N_4165);
or U7403 (N_7403,N_5123,N_5067);
and U7404 (N_7404,N_5230,N_4005);
nand U7405 (N_7405,N_5771,N_5526);
or U7406 (N_7406,N_4730,N_5436);
xnor U7407 (N_7407,N_4281,N_5814);
nor U7408 (N_7408,N_5941,N_5523);
nor U7409 (N_7409,N_5307,N_4146);
and U7410 (N_7410,N_5946,N_4345);
and U7411 (N_7411,N_5886,N_5729);
xnor U7412 (N_7412,N_5185,N_4554);
or U7413 (N_7413,N_4769,N_5165);
xor U7414 (N_7414,N_5438,N_5244);
nor U7415 (N_7415,N_5012,N_5029);
nor U7416 (N_7416,N_4805,N_5892);
and U7417 (N_7417,N_5464,N_4335);
or U7418 (N_7418,N_5340,N_5440);
or U7419 (N_7419,N_5307,N_5246);
xor U7420 (N_7420,N_4175,N_5653);
and U7421 (N_7421,N_5419,N_4256);
xnor U7422 (N_7422,N_5945,N_5093);
and U7423 (N_7423,N_5080,N_4116);
or U7424 (N_7424,N_5835,N_4249);
nor U7425 (N_7425,N_5026,N_5273);
or U7426 (N_7426,N_4345,N_5930);
and U7427 (N_7427,N_4369,N_5168);
or U7428 (N_7428,N_5743,N_4694);
nor U7429 (N_7429,N_5876,N_5994);
or U7430 (N_7430,N_5386,N_5363);
nor U7431 (N_7431,N_5686,N_4203);
nand U7432 (N_7432,N_5851,N_5536);
or U7433 (N_7433,N_5715,N_5019);
or U7434 (N_7434,N_4480,N_4888);
nor U7435 (N_7435,N_5399,N_5664);
xor U7436 (N_7436,N_5710,N_5332);
and U7437 (N_7437,N_4994,N_4196);
nor U7438 (N_7438,N_5006,N_4241);
or U7439 (N_7439,N_4070,N_4290);
and U7440 (N_7440,N_4675,N_4288);
nor U7441 (N_7441,N_4748,N_4598);
nor U7442 (N_7442,N_4091,N_5181);
nor U7443 (N_7443,N_5117,N_4167);
nor U7444 (N_7444,N_5763,N_4006);
nor U7445 (N_7445,N_4586,N_4170);
nor U7446 (N_7446,N_4758,N_5638);
xnor U7447 (N_7447,N_4614,N_4175);
nand U7448 (N_7448,N_5154,N_4729);
nand U7449 (N_7449,N_4090,N_5462);
and U7450 (N_7450,N_5917,N_5549);
nand U7451 (N_7451,N_5395,N_5564);
and U7452 (N_7452,N_5909,N_5718);
or U7453 (N_7453,N_4482,N_4503);
or U7454 (N_7454,N_5214,N_5539);
and U7455 (N_7455,N_5170,N_5360);
xor U7456 (N_7456,N_4789,N_5203);
or U7457 (N_7457,N_4689,N_5471);
and U7458 (N_7458,N_5662,N_4605);
and U7459 (N_7459,N_4283,N_4540);
nand U7460 (N_7460,N_4006,N_4718);
nor U7461 (N_7461,N_5427,N_5931);
nand U7462 (N_7462,N_5223,N_4110);
and U7463 (N_7463,N_5521,N_5817);
nand U7464 (N_7464,N_5200,N_5364);
and U7465 (N_7465,N_5573,N_4793);
or U7466 (N_7466,N_5743,N_4426);
nor U7467 (N_7467,N_5846,N_4865);
nor U7468 (N_7468,N_5378,N_5706);
and U7469 (N_7469,N_5573,N_4788);
and U7470 (N_7470,N_4824,N_5046);
and U7471 (N_7471,N_4933,N_5430);
and U7472 (N_7472,N_5195,N_4830);
nor U7473 (N_7473,N_4390,N_4185);
nor U7474 (N_7474,N_4899,N_4276);
or U7475 (N_7475,N_4332,N_5442);
or U7476 (N_7476,N_5072,N_5772);
nor U7477 (N_7477,N_4561,N_5837);
and U7478 (N_7478,N_4536,N_4209);
nand U7479 (N_7479,N_4968,N_5961);
nor U7480 (N_7480,N_4275,N_5886);
nand U7481 (N_7481,N_4889,N_4208);
nor U7482 (N_7482,N_4398,N_4305);
and U7483 (N_7483,N_5538,N_5681);
and U7484 (N_7484,N_5891,N_5066);
or U7485 (N_7485,N_5159,N_4093);
nand U7486 (N_7486,N_4850,N_5086);
xor U7487 (N_7487,N_4168,N_5543);
or U7488 (N_7488,N_4278,N_5723);
xnor U7489 (N_7489,N_4680,N_5393);
and U7490 (N_7490,N_4957,N_4209);
xnor U7491 (N_7491,N_5311,N_4324);
or U7492 (N_7492,N_5779,N_5569);
or U7493 (N_7493,N_5772,N_5824);
or U7494 (N_7494,N_4103,N_4437);
nor U7495 (N_7495,N_4539,N_4987);
nand U7496 (N_7496,N_4444,N_5296);
nor U7497 (N_7497,N_4093,N_4052);
or U7498 (N_7498,N_4658,N_4596);
and U7499 (N_7499,N_5715,N_4571);
and U7500 (N_7500,N_4494,N_5463);
nand U7501 (N_7501,N_5278,N_4523);
and U7502 (N_7502,N_4769,N_5205);
or U7503 (N_7503,N_5691,N_4120);
or U7504 (N_7504,N_4732,N_5631);
and U7505 (N_7505,N_5690,N_5541);
and U7506 (N_7506,N_4662,N_4509);
or U7507 (N_7507,N_4971,N_5921);
or U7508 (N_7508,N_5270,N_5079);
nand U7509 (N_7509,N_4917,N_5607);
or U7510 (N_7510,N_5500,N_5621);
nor U7511 (N_7511,N_5790,N_4275);
nor U7512 (N_7512,N_5700,N_4099);
nand U7513 (N_7513,N_4149,N_5137);
or U7514 (N_7514,N_5876,N_5144);
nand U7515 (N_7515,N_4588,N_5330);
xor U7516 (N_7516,N_5159,N_4413);
nor U7517 (N_7517,N_5331,N_4852);
nand U7518 (N_7518,N_5785,N_4727);
nor U7519 (N_7519,N_5778,N_4069);
nand U7520 (N_7520,N_5965,N_4774);
xor U7521 (N_7521,N_4826,N_4452);
nor U7522 (N_7522,N_4127,N_5533);
nor U7523 (N_7523,N_4991,N_4107);
nand U7524 (N_7524,N_5469,N_5942);
or U7525 (N_7525,N_4436,N_4397);
or U7526 (N_7526,N_4306,N_4780);
or U7527 (N_7527,N_5354,N_4896);
nor U7528 (N_7528,N_5824,N_4774);
nor U7529 (N_7529,N_5708,N_4466);
nand U7530 (N_7530,N_5525,N_4400);
nor U7531 (N_7531,N_5387,N_5709);
or U7532 (N_7532,N_4909,N_4565);
nor U7533 (N_7533,N_5115,N_5958);
xnor U7534 (N_7534,N_4073,N_4433);
xnor U7535 (N_7535,N_4090,N_5651);
nand U7536 (N_7536,N_4021,N_4498);
nor U7537 (N_7537,N_5127,N_5518);
nor U7538 (N_7538,N_4643,N_4054);
nand U7539 (N_7539,N_5079,N_4902);
nor U7540 (N_7540,N_4797,N_4418);
nand U7541 (N_7541,N_5471,N_5904);
nor U7542 (N_7542,N_4303,N_4054);
nand U7543 (N_7543,N_4696,N_4962);
nor U7544 (N_7544,N_5126,N_5942);
nand U7545 (N_7545,N_4976,N_4370);
or U7546 (N_7546,N_5882,N_5978);
xor U7547 (N_7547,N_5740,N_4818);
and U7548 (N_7548,N_4775,N_4427);
and U7549 (N_7549,N_5647,N_4791);
or U7550 (N_7550,N_5694,N_4300);
nand U7551 (N_7551,N_4061,N_4943);
nand U7552 (N_7552,N_4468,N_4865);
and U7553 (N_7553,N_4991,N_4224);
nand U7554 (N_7554,N_4567,N_5747);
and U7555 (N_7555,N_4464,N_4393);
nor U7556 (N_7556,N_4962,N_4939);
nand U7557 (N_7557,N_5165,N_5387);
nand U7558 (N_7558,N_4786,N_4145);
and U7559 (N_7559,N_4975,N_5480);
or U7560 (N_7560,N_5107,N_4149);
or U7561 (N_7561,N_5371,N_5530);
nor U7562 (N_7562,N_4506,N_5442);
nand U7563 (N_7563,N_4896,N_5431);
nor U7564 (N_7564,N_5764,N_5938);
or U7565 (N_7565,N_4285,N_4493);
and U7566 (N_7566,N_5398,N_5521);
nor U7567 (N_7567,N_5340,N_4554);
nand U7568 (N_7568,N_4759,N_5636);
nand U7569 (N_7569,N_5536,N_5133);
nand U7570 (N_7570,N_5480,N_5924);
nor U7571 (N_7571,N_4115,N_4196);
nor U7572 (N_7572,N_5862,N_5889);
nand U7573 (N_7573,N_4885,N_4767);
nand U7574 (N_7574,N_4378,N_4039);
or U7575 (N_7575,N_5778,N_4162);
or U7576 (N_7576,N_4440,N_5839);
nand U7577 (N_7577,N_5765,N_4607);
and U7578 (N_7578,N_4758,N_5425);
or U7579 (N_7579,N_4438,N_5070);
or U7580 (N_7580,N_5834,N_4012);
and U7581 (N_7581,N_5900,N_4128);
xnor U7582 (N_7582,N_5369,N_4500);
and U7583 (N_7583,N_5812,N_5636);
or U7584 (N_7584,N_5358,N_5666);
xor U7585 (N_7585,N_5879,N_5721);
nand U7586 (N_7586,N_5369,N_4432);
or U7587 (N_7587,N_4057,N_4845);
nand U7588 (N_7588,N_4962,N_5754);
or U7589 (N_7589,N_4631,N_4121);
xnor U7590 (N_7590,N_4638,N_5231);
or U7591 (N_7591,N_4977,N_4469);
or U7592 (N_7592,N_5925,N_5568);
nor U7593 (N_7593,N_5858,N_4750);
or U7594 (N_7594,N_5139,N_5240);
and U7595 (N_7595,N_5263,N_5501);
nor U7596 (N_7596,N_4927,N_5606);
nor U7597 (N_7597,N_4123,N_4169);
or U7598 (N_7598,N_5986,N_5921);
or U7599 (N_7599,N_4688,N_4708);
and U7600 (N_7600,N_4148,N_4835);
and U7601 (N_7601,N_4650,N_5753);
nand U7602 (N_7602,N_4031,N_5907);
nor U7603 (N_7603,N_5125,N_4033);
and U7604 (N_7604,N_4872,N_4624);
or U7605 (N_7605,N_4735,N_4652);
xor U7606 (N_7606,N_5300,N_4541);
nand U7607 (N_7607,N_5685,N_5348);
nand U7608 (N_7608,N_5582,N_5266);
nand U7609 (N_7609,N_5265,N_5101);
or U7610 (N_7610,N_5088,N_5428);
or U7611 (N_7611,N_4351,N_5969);
nor U7612 (N_7612,N_5676,N_4424);
and U7613 (N_7613,N_5453,N_4072);
and U7614 (N_7614,N_4793,N_5954);
nand U7615 (N_7615,N_4319,N_5207);
and U7616 (N_7616,N_5347,N_4914);
nand U7617 (N_7617,N_5319,N_5764);
or U7618 (N_7618,N_4432,N_4684);
xnor U7619 (N_7619,N_5055,N_4897);
nand U7620 (N_7620,N_5060,N_4617);
and U7621 (N_7621,N_4740,N_4060);
or U7622 (N_7622,N_5097,N_5062);
nand U7623 (N_7623,N_5778,N_5463);
nor U7624 (N_7624,N_4862,N_5936);
or U7625 (N_7625,N_5356,N_4456);
nand U7626 (N_7626,N_5905,N_5507);
and U7627 (N_7627,N_5921,N_4658);
xor U7628 (N_7628,N_5538,N_4485);
or U7629 (N_7629,N_4120,N_5443);
nand U7630 (N_7630,N_4922,N_4059);
nor U7631 (N_7631,N_4198,N_5589);
xor U7632 (N_7632,N_4391,N_5390);
xnor U7633 (N_7633,N_4660,N_5805);
nor U7634 (N_7634,N_5474,N_4133);
or U7635 (N_7635,N_5055,N_5200);
and U7636 (N_7636,N_4064,N_5253);
nand U7637 (N_7637,N_5689,N_4932);
nor U7638 (N_7638,N_4363,N_5081);
nor U7639 (N_7639,N_5640,N_5224);
and U7640 (N_7640,N_4409,N_5827);
nand U7641 (N_7641,N_5794,N_5442);
and U7642 (N_7642,N_4477,N_5931);
nand U7643 (N_7643,N_5550,N_5587);
nor U7644 (N_7644,N_4503,N_5256);
nand U7645 (N_7645,N_5910,N_5640);
or U7646 (N_7646,N_4412,N_4662);
and U7647 (N_7647,N_5009,N_4511);
and U7648 (N_7648,N_5131,N_4413);
nor U7649 (N_7649,N_4604,N_5233);
nor U7650 (N_7650,N_4780,N_5453);
and U7651 (N_7651,N_5164,N_4504);
or U7652 (N_7652,N_5397,N_5346);
and U7653 (N_7653,N_5358,N_5525);
nor U7654 (N_7654,N_5661,N_4992);
nand U7655 (N_7655,N_5756,N_4418);
and U7656 (N_7656,N_4846,N_4839);
or U7657 (N_7657,N_4474,N_4808);
or U7658 (N_7658,N_4537,N_4374);
or U7659 (N_7659,N_5554,N_5946);
xnor U7660 (N_7660,N_5154,N_5860);
nor U7661 (N_7661,N_4772,N_4225);
nor U7662 (N_7662,N_5042,N_4567);
or U7663 (N_7663,N_5957,N_4835);
nand U7664 (N_7664,N_5791,N_4343);
nor U7665 (N_7665,N_4965,N_5647);
nor U7666 (N_7666,N_5497,N_4821);
xor U7667 (N_7667,N_4615,N_5953);
or U7668 (N_7668,N_5576,N_5104);
or U7669 (N_7669,N_4928,N_5014);
nand U7670 (N_7670,N_4104,N_5976);
and U7671 (N_7671,N_4053,N_4980);
and U7672 (N_7672,N_4364,N_4529);
or U7673 (N_7673,N_4941,N_4756);
nor U7674 (N_7674,N_5669,N_5271);
nor U7675 (N_7675,N_5610,N_4960);
and U7676 (N_7676,N_5972,N_4881);
nand U7677 (N_7677,N_5371,N_5978);
xnor U7678 (N_7678,N_5315,N_4546);
and U7679 (N_7679,N_5258,N_5743);
nor U7680 (N_7680,N_5638,N_5842);
or U7681 (N_7681,N_5454,N_5550);
or U7682 (N_7682,N_4266,N_5373);
nor U7683 (N_7683,N_4575,N_4774);
or U7684 (N_7684,N_5598,N_5930);
xnor U7685 (N_7685,N_5514,N_4288);
or U7686 (N_7686,N_4465,N_4322);
xor U7687 (N_7687,N_5776,N_5478);
or U7688 (N_7688,N_4913,N_5856);
and U7689 (N_7689,N_5636,N_5834);
or U7690 (N_7690,N_4078,N_4093);
xnor U7691 (N_7691,N_5077,N_5484);
or U7692 (N_7692,N_5685,N_5865);
xnor U7693 (N_7693,N_5198,N_4621);
or U7694 (N_7694,N_4644,N_5840);
nor U7695 (N_7695,N_4205,N_5459);
and U7696 (N_7696,N_4679,N_5325);
and U7697 (N_7697,N_4106,N_5850);
or U7698 (N_7698,N_4619,N_4966);
or U7699 (N_7699,N_4512,N_5389);
and U7700 (N_7700,N_4296,N_4365);
nand U7701 (N_7701,N_4058,N_5608);
xnor U7702 (N_7702,N_4795,N_4945);
nor U7703 (N_7703,N_4003,N_5584);
or U7704 (N_7704,N_4046,N_5915);
nor U7705 (N_7705,N_4615,N_5355);
and U7706 (N_7706,N_4957,N_5640);
and U7707 (N_7707,N_5658,N_5579);
nand U7708 (N_7708,N_5852,N_5870);
or U7709 (N_7709,N_4644,N_4592);
xnor U7710 (N_7710,N_5880,N_4678);
nand U7711 (N_7711,N_5639,N_4313);
and U7712 (N_7712,N_5332,N_5835);
nand U7713 (N_7713,N_4052,N_4382);
and U7714 (N_7714,N_5397,N_5041);
or U7715 (N_7715,N_5979,N_4960);
nand U7716 (N_7716,N_5464,N_4692);
or U7717 (N_7717,N_4227,N_4363);
nand U7718 (N_7718,N_5973,N_5012);
and U7719 (N_7719,N_5300,N_5375);
xor U7720 (N_7720,N_4652,N_4129);
nand U7721 (N_7721,N_4919,N_4485);
or U7722 (N_7722,N_5251,N_5589);
or U7723 (N_7723,N_4122,N_4667);
nor U7724 (N_7724,N_5404,N_5186);
or U7725 (N_7725,N_4730,N_5011);
and U7726 (N_7726,N_4545,N_5385);
or U7727 (N_7727,N_5425,N_5559);
nor U7728 (N_7728,N_5375,N_4729);
or U7729 (N_7729,N_4833,N_5492);
and U7730 (N_7730,N_4688,N_5190);
nand U7731 (N_7731,N_4175,N_4260);
nor U7732 (N_7732,N_5320,N_4565);
and U7733 (N_7733,N_4538,N_5989);
nand U7734 (N_7734,N_5302,N_4188);
nand U7735 (N_7735,N_4941,N_4595);
nor U7736 (N_7736,N_4894,N_4381);
nor U7737 (N_7737,N_5752,N_4072);
nor U7738 (N_7738,N_4463,N_5224);
and U7739 (N_7739,N_5265,N_5912);
nor U7740 (N_7740,N_4631,N_4083);
nor U7741 (N_7741,N_5188,N_4395);
nor U7742 (N_7742,N_5387,N_5400);
and U7743 (N_7743,N_4006,N_5260);
nand U7744 (N_7744,N_5557,N_5746);
nand U7745 (N_7745,N_4837,N_5870);
nor U7746 (N_7746,N_5881,N_4310);
xor U7747 (N_7747,N_4388,N_5571);
and U7748 (N_7748,N_4063,N_4917);
nor U7749 (N_7749,N_5465,N_4283);
and U7750 (N_7750,N_4743,N_5745);
nand U7751 (N_7751,N_5261,N_4938);
and U7752 (N_7752,N_5137,N_4079);
or U7753 (N_7753,N_5166,N_5368);
nor U7754 (N_7754,N_5165,N_5661);
or U7755 (N_7755,N_4078,N_4972);
and U7756 (N_7756,N_5779,N_4651);
and U7757 (N_7757,N_5997,N_4740);
and U7758 (N_7758,N_5744,N_5651);
and U7759 (N_7759,N_5720,N_5923);
xor U7760 (N_7760,N_5829,N_4633);
nor U7761 (N_7761,N_4304,N_5134);
xor U7762 (N_7762,N_4329,N_5408);
and U7763 (N_7763,N_5618,N_5651);
nand U7764 (N_7764,N_4295,N_4463);
nand U7765 (N_7765,N_4717,N_5371);
nand U7766 (N_7766,N_4507,N_4954);
nor U7767 (N_7767,N_5702,N_5235);
nand U7768 (N_7768,N_4725,N_5702);
xnor U7769 (N_7769,N_5005,N_4387);
and U7770 (N_7770,N_5863,N_5993);
nor U7771 (N_7771,N_5140,N_4096);
and U7772 (N_7772,N_4898,N_5945);
and U7773 (N_7773,N_5655,N_4164);
and U7774 (N_7774,N_4101,N_4988);
or U7775 (N_7775,N_5421,N_5374);
nor U7776 (N_7776,N_5318,N_4038);
and U7777 (N_7777,N_5556,N_5623);
or U7778 (N_7778,N_5260,N_4224);
nor U7779 (N_7779,N_4623,N_4206);
nand U7780 (N_7780,N_4773,N_4407);
xor U7781 (N_7781,N_4232,N_4163);
nor U7782 (N_7782,N_4794,N_5106);
nor U7783 (N_7783,N_5460,N_4615);
xor U7784 (N_7784,N_4213,N_4764);
xnor U7785 (N_7785,N_5926,N_4978);
xnor U7786 (N_7786,N_5554,N_4032);
nand U7787 (N_7787,N_5591,N_5862);
nor U7788 (N_7788,N_4658,N_5170);
nor U7789 (N_7789,N_4532,N_5401);
nor U7790 (N_7790,N_5759,N_5647);
nor U7791 (N_7791,N_5458,N_4443);
nand U7792 (N_7792,N_4601,N_5395);
nor U7793 (N_7793,N_5179,N_5561);
or U7794 (N_7794,N_5333,N_5055);
nand U7795 (N_7795,N_4726,N_4663);
or U7796 (N_7796,N_5642,N_4934);
and U7797 (N_7797,N_4087,N_4762);
and U7798 (N_7798,N_4553,N_5127);
nor U7799 (N_7799,N_4455,N_5664);
or U7800 (N_7800,N_4553,N_5069);
nand U7801 (N_7801,N_4199,N_5740);
and U7802 (N_7802,N_5489,N_5260);
nor U7803 (N_7803,N_4289,N_5148);
nand U7804 (N_7804,N_4861,N_4977);
nor U7805 (N_7805,N_5820,N_4413);
or U7806 (N_7806,N_5529,N_5601);
and U7807 (N_7807,N_5161,N_4035);
nand U7808 (N_7808,N_4879,N_5032);
and U7809 (N_7809,N_5233,N_4846);
or U7810 (N_7810,N_5782,N_5204);
nand U7811 (N_7811,N_5640,N_5087);
nor U7812 (N_7812,N_5690,N_4104);
or U7813 (N_7813,N_5760,N_4415);
nor U7814 (N_7814,N_4229,N_5895);
and U7815 (N_7815,N_5414,N_4470);
nor U7816 (N_7816,N_5698,N_5305);
xnor U7817 (N_7817,N_4919,N_4622);
or U7818 (N_7818,N_5822,N_4233);
nor U7819 (N_7819,N_4329,N_5963);
nor U7820 (N_7820,N_4440,N_5957);
nor U7821 (N_7821,N_5376,N_5064);
and U7822 (N_7822,N_4474,N_5431);
or U7823 (N_7823,N_4566,N_4898);
or U7824 (N_7824,N_5561,N_5316);
or U7825 (N_7825,N_4082,N_5792);
and U7826 (N_7826,N_4365,N_5165);
and U7827 (N_7827,N_4752,N_4398);
and U7828 (N_7828,N_5810,N_4545);
or U7829 (N_7829,N_4502,N_5421);
or U7830 (N_7830,N_4153,N_5987);
nand U7831 (N_7831,N_5757,N_5601);
or U7832 (N_7832,N_5379,N_4609);
nand U7833 (N_7833,N_5367,N_5483);
or U7834 (N_7834,N_4479,N_4988);
or U7835 (N_7835,N_4090,N_5285);
or U7836 (N_7836,N_5008,N_4751);
nor U7837 (N_7837,N_5501,N_5329);
nand U7838 (N_7838,N_4961,N_5835);
nor U7839 (N_7839,N_5317,N_5471);
nor U7840 (N_7840,N_5201,N_4943);
nand U7841 (N_7841,N_4327,N_5843);
xnor U7842 (N_7842,N_4322,N_5101);
xor U7843 (N_7843,N_5927,N_4859);
nor U7844 (N_7844,N_4983,N_5920);
and U7845 (N_7845,N_5346,N_5951);
nor U7846 (N_7846,N_5271,N_4462);
nand U7847 (N_7847,N_5721,N_4886);
nor U7848 (N_7848,N_5286,N_4850);
xor U7849 (N_7849,N_4476,N_4153);
or U7850 (N_7850,N_5152,N_4345);
or U7851 (N_7851,N_4085,N_5472);
or U7852 (N_7852,N_5153,N_5657);
and U7853 (N_7853,N_4441,N_5307);
nand U7854 (N_7854,N_5066,N_5666);
nand U7855 (N_7855,N_4884,N_4247);
nand U7856 (N_7856,N_4242,N_4094);
xnor U7857 (N_7857,N_4277,N_4990);
nand U7858 (N_7858,N_4606,N_5256);
or U7859 (N_7859,N_4558,N_4330);
xor U7860 (N_7860,N_5924,N_5178);
nand U7861 (N_7861,N_5953,N_4355);
xnor U7862 (N_7862,N_4917,N_5465);
and U7863 (N_7863,N_4366,N_4246);
or U7864 (N_7864,N_5877,N_4050);
xor U7865 (N_7865,N_5692,N_5696);
or U7866 (N_7866,N_5945,N_5171);
nand U7867 (N_7867,N_5430,N_4470);
or U7868 (N_7868,N_4242,N_4305);
or U7869 (N_7869,N_5390,N_5726);
and U7870 (N_7870,N_4892,N_4318);
xnor U7871 (N_7871,N_5168,N_4039);
nor U7872 (N_7872,N_4604,N_4178);
or U7873 (N_7873,N_5678,N_4775);
nand U7874 (N_7874,N_5242,N_4598);
or U7875 (N_7875,N_5729,N_5236);
and U7876 (N_7876,N_5776,N_4314);
and U7877 (N_7877,N_5314,N_5465);
and U7878 (N_7878,N_4002,N_4532);
or U7879 (N_7879,N_5487,N_5848);
nand U7880 (N_7880,N_4936,N_4846);
and U7881 (N_7881,N_4959,N_4384);
and U7882 (N_7882,N_5771,N_5339);
nor U7883 (N_7883,N_4203,N_5103);
nand U7884 (N_7884,N_5182,N_5205);
and U7885 (N_7885,N_4200,N_4355);
nand U7886 (N_7886,N_5714,N_5496);
and U7887 (N_7887,N_5807,N_5816);
nor U7888 (N_7888,N_5949,N_4786);
nor U7889 (N_7889,N_5981,N_5914);
or U7890 (N_7890,N_5278,N_5479);
nor U7891 (N_7891,N_5153,N_5338);
and U7892 (N_7892,N_5240,N_5150);
xnor U7893 (N_7893,N_4712,N_5310);
or U7894 (N_7894,N_4898,N_4071);
or U7895 (N_7895,N_4184,N_4805);
and U7896 (N_7896,N_4385,N_5732);
nand U7897 (N_7897,N_5635,N_5005);
xnor U7898 (N_7898,N_5601,N_5871);
nor U7899 (N_7899,N_5679,N_4753);
and U7900 (N_7900,N_5363,N_5723);
or U7901 (N_7901,N_4978,N_5594);
or U7902 (N_7902,N_4675,N_5209);
nand U7903 (N_7903,N_4737,N_5141);
or U7904 (N_7904,N_4573,N_4496);
and U7905 (N_7905,N_4216,N_5687);
or U7906 (N_7906,N_5930,N_4446);
nor U7907 (N_7907,N_5122,N_5760);
nor U7908 (N_7908,N_5445,N_5305);
nor U7909 (N_7909,N_5734,N_5101);
nand U7910 (N_7910,N_5271,N_4427);
and U7911 (N_7911,N_4265,N_5034);
nor U7912 (N_7912,N_4310,N_5808);
or U7913 (N_7913,N_5997,N_5239);
or U7914 (N_7914,N_5912,N_5154);
nand U7915 (N_7915,N_4443,N_5566);
nand U7916 (N_7916,N_5373,N_4256);
nand U7917 (N_7917,N_4423,N_4140);
or U7918 (N_7918,N_5195,N_5099);
and U7919 (N_7919,N_4544,N_4092);
or U7920 (N_7920,N_5570,N_5288);
and U7921 (N_7921,N_5110,N_5399);
or U7922 (N_7922,N_4970,N_4043);
or U7923 (N_7923,N_5263,N_4891);
nand U7924 (N_7924,N_5879,N_5746);
and U7925 (N_7925,N_5547,N_4781);
nor U7926 (N_7926,N_4135,N_4124);
and U7927 (N_7927,N_4378,N_4644);
nand U7928 (N_7928,N_4430,N_5516);
and U7929 (N_7929,N_4742,N_5709);
nor U7930 (N_7930,N_4650,N_4502);
xor U7931 (N_7931,N_5152,N_4036);
nor U7932 (N_7932,N_5824,N_4861);
and U7933 (N_7933,N_4870,N_5731);
nor U7934 (N_7934,N_4045,N_4224);
nand U7935 (N_7935,N_5879,N_4465);
nor U7936 (N_7936,N_4351,N_4323);
nor U7937 (N_7937,N_4472,N_5703);
xor U7938 (N_7938,N_5918,N_5196);
nand U7939 (N_7939,N_5033,N_5936);
and U7940 (N_7940,N_4752,N_5195);
or U7941 (N_7941,N_5093,N_5623);
nor U7942 (N_7942,N_5161,N_4327);
nor U7943 (N_7943,N_4812,N_5922);
nor U7944 (N_7944,N_4931,N_5764);
and U7945 (N_7945,N_5323,N_5949);
nand U7946 (N_7946,N_5104,N_4528);
and U7947 (N_7947,N_5195,N_5358);
nand U7948 (N_7948,N_5950,N_4718);
or U7949 (N_7949,N_4732,N_4366);
nand U7950 (N_7950,N_5886,N_5335);
or U7951 (N_7951,N_4028,N_4345);
nor U7952 (N_7952,N_5466,N_5111);
xnor U7953 (N_7953,N_5840,N_5018);
or U7954 (N_7954,N_4220,N_5462);
nor U7955 (N_7955,N_5671,N_5562);
and U7956 (N_7956,N_4065,N_4667);
and U7957 (N_7957,N_4067,N_5495);
nor U7958 (N_7958,N_4128,N_5289);
or U7959 (N_7959,N_5384,N_4580);
or U7960 (N_7960,N_4237,N_4985);
and U7961 (N_7961,N_5854,N_5253);
nor U7962 (N_7962,N_5677,N_4736);
or U7963 (N_7963,N_5977,N_5457);
xor U7964 (N_7964,N_5766,N_4027);
nand U7965 (N_7965,N_5278,N_4910);
nor U7966 (N_7966,N_4993,N_5818);
or U7967 (N_7967,N_5757,N_4994);
or U7968 (N_7968,N_5281,N_5337);
and U7969 (N_7969,N_5887,N_5557);
nand U7970 (N_7970,N_4572,N_4693);
nand U7971 (N_7971,N_4402,N_4915);
nand U7972 (N_7972,N_4565,N_5584);
and U7973 (N_7973,N_4563,N_4250);
or U7974 (N_7974,N_5477,N_4445);
and U7975 (N_7975,N_5180,N_4252);
nor U7976 (N_7976,N_5342,N_4756);
or U7977 (N_7977,N_4823,N_4799);
and U7978 (N_7978,N_5239,N_4033);
nand U7979 (N_7979,N_4408,N_5085);
nand U7980 (N_7980,N_5356,N_4706);
nor U7981 (N_7981,N_5903,N_5134);
xor U7982 (N_7982,N_4196,N_5797);
xor U7983 (N_7983,N_4769,N_5752);
or U7984 (N_7984,N_4557,N_5789);
nor U7985 (N_7985,N_4731,N_4571);
xnor U7986 (N_7986,N_5155,N_4129);
and U7987 (N_7987,N_4477,N_4166);
nand U7988 (N_7988,N_4091,N_4185);
nand U7989 (N_7989,N_4317,N_5160);
and U7990 (N_7990,N_4329,N_4373);
xor U7991 (N_7991,N_5286,N_4093);
nand U7992 (N_7992,N_4953,N_5354);
and U7993 (N_7993,N_5129,N_4577);
nand U7994 (N_7994,N_5879,N_4553);
and U7995 (N_7995,N_5122,N_5653);
nor U7996 (N_7996,N_5724,N_4462);
and U7997 (N_7997,N_5240,N_4415);
xor U7998 (N_7998,N_5819,N_5732);
or U7999 (N_7999,N_4919,N_4705);
nand U8000 (N_8000,N_6147,N_7031);
nor U8001 (N_8001,N_7873,N_7215);
nand U8002 (N_8002,N_7808,N_6264);
or U8003 (N_8003,N_6241,N_7434);
and U8004 (N_8004,N_6851,N_7381);
nor U8005 (N_8005,N_6565,N_6761);
and U8006 (N_8006,N_6848,N_6063);
nor U8007 (N_8007,N_7401,N_7298);
or U8008 (N_8008,N_7986,N_7322);
xor U8009 (N_8009,N_6963,N_6987);
nand U8010 (N_8010,N_6204,N_6925);
and U8011 (N_8011,N_7084,N_6237);
and U8012 (N_8012,N_6605,N_6990);
or U8013 (N_8013,N_7558,N_6879);
nor U8014 (N_8014,N_6575,N_6858);
and U8015 (N_8015,N_7019,N_7767);
or U8016 (N_8016,N_6236,N_7646);
and U8017 (N_8017,N_7069,N_7457);
nor U8018 (N_8018,N_7036,N_6257);
or U8019 (N_8019,N_6459,N_7086);
nor U8020 (N_8020,N_6277,N_6569);
nor U8021 (N_8021,N_6956,N_7487);
xnor U8022 (N_8022,N_7200,N_6056);
nor U8023 (N_8023,N_6768,N_6642);
or U8024 (N_8024,N_7929,N_7095);
xor U8025 (N_8025,N_6300,N_7917);
nor U8026 (N_8026,N_7476,N_6545);
or U8027 (N_8027,N_6746,N_7816);
nor U8028 (N_8028,N_7000,N_7516);
or U8029 (N_8029,N_6296,N_7283);
nor U8030 (N_8030,N_6738,N_6188);
or U8031 (N_8031,N_7587,N_6415);
nor U8032 (N_8032,N_6064,N_7602);
or U8033 (N_8033,N_6551,N_6590);
nor U8034 (N_8034,N_6330,N_7217);
xnor U8035 (N_8035,N_6492,N_7009);
nand U8036 (N_8036,N_7969,N_7409);
nor U8037 (N_8037,N_7778,N_7752);
and U8038 (N_8038,N_6409,N_6627);
and U8039 (N_8039,N_7187,N_7888);
and U8040 (N_8040,N_6539,N_7053);
nor U8041 (N_8041,N_7327,N_7363);
and U8042 (N_8042,N_7337,N_7334);
nor U8043 (N_8043,N_6600,N_7681);
nor U8044 (N_8044,N_7208,N_6484);
nor U8045 (N_8045,N_6587,N_7670);
nor U8046 (N_8046,N_7464,N_6391);
nor U8047 (N_8047,N_7291,N_6903);
or U8048 (N_8048,N_7403,N_7627);
nor U8049 (N_8049,N_7512,N_7912);
or U8050 (N_8050,N_7211,N_7539);
nand U8051 (N_8051,N_6230,N_6473);
and U8052 (N_8052,N_7206,N_6747);
nand U8053 (N_8053,N_6502,N_7796);
and U8054 (N_8054,N_7465,N_7210);
nor U8055 (N_8055,N_7102,N_7046);
and U8056 (N_8056,N_6643,N_7357);
nor U8057 (N_8057,N_6304,N_6465);
nor U8058 (N_8058,N_7252,N_7544);
xor U8059 (N_8059,N_7203,N_6468);
nor U8060 (N_8060,N_7571,N_7493);
and U8061 (N_8061,N_6035,N_6291);
nand U8062 (N_8062,N_6080,N_6788);
and U8063 (N_8063,N_6434,N_6198);
xor U8064 (N_8064,N_6666,N_6352);
xnor U8065 (N_8065,N_7529,N_6295);
and U8066 (N_8066,N_7010,N_7073);
nand U8067 (N_8067,N_6260,N_7345);
nand U8068 (N_8068,N_6714,N_7109);
nand U8069 (N_8069,N_7205,N_7887);
or U8070 (N_8070,N_6262,N_7309);
nor U8071 (N_8071,N_6057,N_6427);
and U8072 (N_8072,N_7197,N_6730);
xnor U8073 (N_8073,N_6027,N_6396);
xor U8074 (N_8074,N_7083,N_6022);
xor U8075 (N_8075,N_6458,N_6496);
and U8076 (N_8076,N_6856,N_6753);
nand U8077 (N_8077,N_6322,N_7908);
and U8078 (N_8078,N_6633,N_6685);
xnor U8079 (N_8079,N_7249,N_7076);
xor U8080 (N_8080,N_7899,N_6461);
or U8081 (N_8081,N_6735,N_7325);
nor U8082 (N_8082,N_6374,N_6514);
nand U8083 (N_8083,N_7407,N_6001);
or U8084 (N_8084,N_7154,N_6966);
nand U8085 (N_8085,N_7007,N_7843);
nor U8086 (N_8086,N_6896,N_7624);
or U8087 (N_8087,N_6214,N_7896);
and U8088 (N_8088,N_7270,N_7675);
and U8089 (N_8089,N_6683,N_7127);
nor U8090 (N_8090,N_6517,N_6721);
and U8091 (N_8091,N_6478,N_7994);
and U8092 (N_8092,N_6348,N_7295);
or U8093 (N_8093,N_6748,N_6782);
and U8094 (N_8094,N_6696,N_6549);
or U8095 (N_8095,N_7920,N_6594);
nor U8096 (N_8096,N_7718,N_7108);
or U8097 (N_8097,N_7674,N_6499);
nand U8098 (N_8098,N_6049,N_7094);
and U8099 (N_8099,N_7881,N_6139);
or U8100 (N_8100,N_6812,N_7915);
xor U8101 (N_8101,N_6155,N_7429);
nor U8102 (N_8102,N_6258,N_6687);
and U8103 (N_8103,N_6135,N_6610);
and U8104 (N_8104,N_7745,N_6331);
and U8105 (N_8105,N_7134,N_6061);
or U8106 (N_8106,N_6817,N_6611);
nor U8107 (N_8107,N_6711,N_6612);
or U8108 (N_8108,N_7408,N_6273);
nand U8109 (N_8109,N_6649,N_6926);
or U8110 (N_8110,N_7157,N_6112);
nor U8111 (N_8111,N_7836,N_6104);
and U8112 (N_8112,N_7034,N_6560);
and U8113 (N_8113,N_7607,N_6238);
xnor U8114 (N_8114,N_7188,N_6037);
nand U8115 (N_8115,N_7444,N_7064);
nor U8116 (N_8116,N_6816,N_7097);
and U8117 (N_8117,N_6981,N_7030);
or U8118 (N_8118,N_7405,N_7780);
nand U8119 (N_8119,N_6213,N_7932);
nand U8120 (N_8120,N_7443,N_7527);
or U8121 (N_8121,N_7015,N_7425);
and U8122 (N_8122,N_7501,N_7140);
and U8123 (N_8123,N_7642,N_6700);
or U8124 (N_8124,N_6176,N_7844);
and U8125 (N_8125,N_6286,N_6640);
xnor U8126 (N_8126,N_7988,N_6799);
and U8127 (N_8127,N_7124,N_7392);
or U8128 (N_8128,N_6441,N_6708);
nand U8129 (N_8129,N_7411,N_7850);
and U8130 (N_8130,N_6947,N_6327);
nand U8131 (N_8131,N_7286,N_7535);
and U8132 (N_8132,N_7546,N_6092);
and U8133 (N_8133,N_6486,N_7940);
xor U8134 (N_8134,N_7687,N_6538);
nand U8135 (N_8135,N_7554,N_6664);
or U8136 (N_8136,N_6900,N_6979);
nor U8137 (N_8137,N_7742,N_6224);
nor U8138 (N_8138,N_7166,N_6574);
nor U8139 (N_8139,N_7107,N_7694);
nor U8140 (N_8140,N_6046,N_7671);
or U8141 (N_8141,N_6173,N_7077);
nor U8142 (N_8142,N_6862,N_7002);
or U8143 (N_8143,N_6247,N_7864);
nor U8144 (N_8144,N_7787,N_6680);
or U8145 (N_8145,N_7641,N_6452);
and U8146 (N_8146,N_6393,N_7279);
xnor U8147 (N_8147,N_7978,N_6240);
and U8148 (N_8148,N_6703,N_7532);
or U8149 (N_8149,N_6618,N_6002);
nand U8150 (N_8150,N_7598,N_7042);
or U8151 (N_8151,N_6929,N_7592);
nand U8152 (N_8152,N_7852,N_6191);
nand U8153 (N_8153,N_7093,N_7989);
xor U8154 (N_8154,N_6078,N_6119);
nor U8155 (N_8155,N_6655,N_6811);
and U8156 (N_8156,N_7751,N_6839);
and U8157 (N_8157,N_6794,N_6469);
xor U8158 (N_8158,N_6462,N_6637);
nand U8159 (N_8159,N_6945,N_6973);
or U8160 (N_8160,N_6242,N_6184);
nor U8161 (N_8161,N_7763,N_6202);
and U8162 (N_8162,N_6248,N_7739);
nor U8163 (N_8163,N_7660,N_7474);
nor U8164 (N_8164,N_6233,N_6067);
and U8165 (N_8165,N_7824,N_7563);
or U8166 (N_8166,N_7186,N_6471);
and U8167 (N_8167,N_6940,N_6361);
nand U8168 (N_8168,N_7927,N_6624);
and U8169 (N_8169,N_6239,N_7386);
nand U8170 (N_8170,N_7891,N_7182);
nor U8171 (N_8171,N_6091,N_6228);
or U8172 (N_8172,N_7422,N_6373);
nand U8173 (N_8173,N_6846,N_7013);
and U8174 (N_8174,N_7623,N_6040);
nand U8175 (N_8175,N_7479,N_7936);
xnor U8176 (N_8176,N_6036,N_6394);
nor U8177 (N_8177,N_7370,N_6166);
or U8178 (N_8178,N_7551,N_6494);
or U8179 (N_8179,N_6745,N_7894);
and U8180 (N_8180,N_6132,N_7358);
and U8181 (N_8181,N_7471,N_6907);
nor U8182 (N_8182,N_7014,N_7880);
nor U8183 (N_8183,N_6977,N_7058);
and U8184 (N_8184,N_7290,N_6775);
xor U8185 (N_8185,N_6466,N_6579);
xnor U8186 (N_8186,N_6426,N_7236);
nor U8187 (N_8187,N_7938,N_6250);
and U8188 (N_8188,N_7181,N_6029);
or U8189 (N_8189,N_6842,N_7770);
nand U8190 (N_8190,N_7885,N_6321);
nor U8191 (N_8191,N_7667,N_7918);
nand U8192 (N_8192,N_6491,N_6408);
and U8193 (N_8193,N_6283,N_6095);
nand U8194 (N_8194,N_6975,N_7586);
nand U8195 (N_8195,N_7606,N_6523);
xnor U8196 (N_8196,N_7721,N_7673);
or U8197 (N_8197,N_7662,N_7934);
xnor U8198 (N_8198,N_6834,N_6720);
nand U8199 (N_8199,N_6149,N_6728);
nor U8200 (N_8200,N_6167,N_6397);
nor U8201 (N_8201,N_6103,N_6252);
or U8202 (N_8202,N_6395,N_7819);
xor U8203 (N_8203,N_7343,N_6456);
xor U8204 (N_8204,N_7706,N_7065);
and U8205 (N_8205,N_6174,N_6784);
or U8206 (N_8206,N_7815,N_6678);
nand U8207 (N_8207,N_7113,N_7783);
xor U8208 (N_8208,N_6561,N_7608);
xnor U8209 (N_8209,N_7591,N_6619);
and U8210 (N_8210,N_6912,N_6559);
nand U8211 (N_8211,N_6644,N_6853);
nor U8212 (N_8212,N_7132,N_6333);
and U8213 (N_8213,N_7521,N_7016);
and U8214 (N_8214,N_6133,N_7189);
and U8215 (N_8215,N_7398,N_7074);
nor U8216 (N_8216,N_7690,N_7241);
and U8217 (N_8217,N_7812,N_6197);
nand U8218 (N_8218,N_7404,N_7332);
and U8219 (N_8219,N_6392,N_6163);
nor U8220 (N_8220,N_7461,N_7294);
nor U8221 (N_8221,N_7483,N_6553);
nand U8222 (N_8222,N_6054,N_6875);
and U8223 (N_8223,N_6079,N_7976);
xnor U8224 (N_8224,N_7289,N_7027);
nand U8225 (N_8225,N_7958,N_7017);
or U8226 (N_8226,N_7305,N_7903);
and U8227 (N_8227,N_6910,N_6855);
nand U8228 (N_8228,N_7696,N_7230);
nor U8229 (N_8229,N_6860,N_7484);
nand U8230 (N_8230,N_7922,N_7272);
xor U8231 (N_8231,N_6004,N_7513);
nor U8232 (N_8232,N_6183,N_6449);
nor U8233 (N_8233,N_7703,N_7428);
nor U8234 (N_8234,N_7541,N_7259);
nand U8235 (N_8235,N_6108,N_6222);
nor U8236 (N_8236,N_7734,N_7306);
nor U8237 (N_8237,N_6866,N_6109);
and U8238 (N_8238,N_7697,N_6513);
xor U8239 (N_8239,N_7238,N_6769);
nand U8240 (N_8240,N_7713,N_7910);
and U8241 (N_8241,N_6765,N_6121);
or U8242 (N_8242,N_7818,N_7245);
nand U8243 (N_8243,N_7583,N_7119);
xor U8244 (N_8244,N_7080,N_6127);
xor U8245 (N_8245,N_6725,N_6805);
and U8246 (N_8246,N_7090,N_7098);
nand U8247 (N_8247,N_6152,N_7364);
or U8248 (N_8248,N_7665,N_7717);
xnor U8249 (N_8249,N_6882,N_6620);
nor U8250 (N_8250,N_7420,N_6086);
nor U8251 (N_8251,N_7835,N_7982);
nor U8252 (N_8252,N_7360,N_6013);
nand U8253 (N_8253,N_6504,N_7302);
nor U8254 (N_8254,N_6350,N_7079);
nand U8255 (N_8255,N_6182,N_7255);
xor U8256 (N_8256,N_6457,N_7509);
or U8257 (N_8257,N_6942,N_6845);
and U8258 (N_8258,N_7384,N_6582);
nand U8259 (N_8259,N_7515,N_7728);
and U8260 (N_8260,N_7693,N_6636);
or U8261 (N_8261,N_6081,N_7239);
nand U8262 (N_8262,N_6810,N_7247);
nor U8263 (N_8263,N_7737,N_7643);
or U8264 (N_8264,N_7112,N_7389);
or U8265 (N_8265,N_6442,N_6278);
nor U8266 (N_8266,N_6573,N_6930);
nor U8267 (N_8267,N_6244,N_6557);
nor U8268 (N_8268,N_7339,N_6325);
and U8269 (N_8269,N_6501,N_7326);
nor U8270 (N_8270,N_7913,N_7158);
xor U8271 (N_8271,N_7235,N_7984);
or U8272 (N_8272,N_7024,N_7234);
nor U8273 (N_8273,N_7757,N_7178);
xnor U8274 (N_8274,N_6251,N_7176);
nand U8275 (N_8275,N_7765,N_6967);
xnor U8276 (N_8276,N_7820,N_6776);
xnor U8277 (N_8277,N_7756,N_7975);
nor U8278 (N_8278,N_7284,N_7822);
nand U8279 (N_8279,N_7710,N_6915);
nand U8280 (N_8280,N_6012,N_7271);
or U8281 (N_8281,N_7865,N_6195);
nor U8282 (N_8282,N_6177,N_7099);
or U8283 (N_8283,N_6229,N_6976);
nor U8284 (N_8284,N_7350,N_6707);
or U8285 (N_8285,N_7658,N_6863);
xnor U8286 (N_8286,N_7365,N_7695);
nor U8287 (N_8287,N_6740,N_7388);
and U8288 (N_8288,N_6764,N_7463);
nor U8289 (N_8289,N_6285,N_7705);
or U8290 (N_8290,N_7897,N_7629);
and U8291 (N_8291,N_7831,N_7803);
and U8292 (N_8292,N_6245,N_6343);
or U8293 (N_8293,N_6652,N_6570);
xnor U8294 (N_8294,N_6632,N_7638);
nand U8295 (N_8295,N_6943,N_7653);
and U8296 (N_8296,N_7995,N_6450);
and U8297 (N_8297,N_6511,N_6781);
nand U8298 (N_8298,N_7611,N_7048);
nand U8299 (N_8299,N_6181,N_6010);
xor U8300 (N_8300,N_7089,N_7147);
nand U8301 (N_8301,N_7714,N_6686);
or U8302 (N_8302,N_7761,N_7258);
or U8303 (N_8303,N_6448,N_7898);
or U8304 (N_8304,N_6309,N_6998);
nand U8305 (N_8305,N_6367,N_6463);
nand U8306 (N_8306,N_6984,N_7806);
and U8307 (N_8307,N_7814,N_7735);
nor U8308 (N_8308,N_6822,N_7315);
nor U8309 (N_8309,N_7135,N_6288);
or U8310 (N_8310,N_6881,N_6113);
nor U8311 (N_8311,N_7626,N_6274);
and U8312 (N_8312,N_6071,N_7954);
nor U8313 (N_8313,N_7771,N_6602);
nand U8314 (N_8314,N_6340,N_6718);
and U8315 (N_8315,N_7799,N_6335);
and U8316 (N_8316,N_7273,N_6803);
or U8317 (N_8317,N_6980,N_7688);
and U8318 (N_8318,N_6047,N_7453);
and U8319 (N_8319,N_6031,N_6089);
or U8320 (N_8320,N_7870,N_7834);
xnor U8321 (N_8321,N_6008,N_7860);
nor U8322 (N_8322,N_7123,N_7753);
nand U8323 (N_8323,N_7467,N_6555);
nor U8324 (N_8324,N_7828,N_7595);
nor U8325 (N_8325,N_6952,N_6556);
nor U8326 (N_8326,N_6464,N_6151);
xor U8327 (N_8327,N_7825,N_6532);
and U8328 (N_8328,N_7656,N_7227);
nand U8329 (N_8329,N_6783,N_6982);
nor U8330 (N_8330,N_7222,N_6599);
and U8331 (N_8331,N_6922,N_6682);
xnor U8332 (N_8332,N_7506,N_6698);
or U8333 (N_8333,N_7435,N_6874);
nor U8334 (N_8334,N_6411,N_6887);
nor U8335 (N_8335,N_6835,N_6261);
and U8336 (N_8336,N_7576,N_6017);
or U8337 (N_8337,N_7689,N_7307);
nor U8338 (N_8338,N_6535,N_7029);
and U8339 (N_8339,N_7297,N_7971);
xor U8340 (N_8340,N_6604,N_7025);
and U8341 (N_8341,N_7341,N_7256);
xnor U8342 (N_8342,N_7666,N_7191);
nor U8343 (N_8343,N_7415,N_6186);
nand U8344 (N_8344,N_6986,N_7857);
or U8345 (N_8345,N_6840,N_7708);
nor U8346 (N_8346,N_6737,N_7723);
or U8347 (N_8347,N_7281,N_7138);
or U8348 (N_8348,N_7946,N_7055);
and U8349 (N_8349,N_6097,N_6613);
and U8350 (N_8350,N_7021,N_7747);
nor U8351 (N_8351,N_7131,N_7679);
nand U8352 (N_8352,N_7565,N_7151);
or U8353 (N_8353,N_7573,N_7331);
nand U8354 (N_8354,N_6412,N_7202);
and U8355 (N_8355,N_6398,N_6476);
nor U8356 (N_8356,N_7352,N_6428);
nand U8357 (N_8357,N_7242,N_6650);
or U8358 (N_8358,N_6914,N_7199);
nand U8359 (N_8359,N_7848,N_6847);
nor U8360 (N_8360,N_7101,N_7701);
or U8361 (N_8361,N_7669,N_6774);
or U8362 (N_8362,N_6493,N_6052);
nor U8363 (N_8363,N_6364,N_6212);
nand U8364 (N_8364,N_7488,N_7762);
nand U8365 (N_8365,N_7416,N_7071);
or U8366 (N_8366,N_7589,N_6219);
and U8367 (N_8367,N_7059,N_7584);
and U8368 (N_8368,N_7702,N_7051);
xnor U8369 (N_8369,N_6315,N_7862);
or U8370 (N_8370,N_7351,N_6292);
xnor U8371 (N_8371,N_7125,N_6886);
and U8372 (N_8372,N_6438,N_6281);
nor U8373 (N_8373,N_7141,N_7128);
and U8374 (N_8374,N_6075,N_6231);
nand U8375 (N_8375,N_6094,N_7323);
or U8376 (N_8376,N_7035,N_6485);
or U8377 (N_8377,N_7433,N_6578);
nand U8378 (N_8378,N_7028,N_7872);
xor U8379 (N_8379,N_7011,N_6892);
or U8380 (N_8380,N_6148,N_7939);
nand U8381 (N_8381,N_6924,N_6607);
or U8382 (N_8382,N_7460,N_6430);
and U8383 (N_8383,N_7970,N_6477);
nor U8384 (N_8384,N_6772,N_6105);
nand U8385 (N_8385,N_7937,N_6934);
nand U8386 (N_8386,N_7263,N_7481);
nand U8387 (N_8387,N_6994,N_6821);
and U8388 (N_8388,N_7324,N_6324);
nor U8389 (N_8389,N_7562,N_7746);
and U8390 (N_8390,N_6701,N_7981);
or U8391 (N_8391,N_6960,N_6388);
or U8392 (N_8392,N_7489,N_6505);
xnor U8393 (N_8393,N_6736,N_6669);
nand U8394 (N_8394,N_7786,N_6741);
nor U8395 (N_8395,N_6066,N_6993);
and U8396 (N_8396,N_6813,N_6717);
nand U8397 (N_8397,N_7963,N_7725);
and U8398 (N_8398,N_6358,N_6142);
nand U8399 (N_8399,N_7413,N_6332);
nor U8400 (N_8400,N_6927,N_6280);
and U8401 (N_8401,N_6831,N_7261);
and U8402 (N_8402,N_7537,N_6826);
and U8403 (N_8403,N_7711,N_6709);
or U8404 (N_8404,N_7630,N_7867);
and U8405 (N_8405,N_7317,N_6524);
nand U8406 (N_8406,N_6823,N_7397);
and U8407 (N_8407,N_6082,N_7190);
nand U8408 (N_8408,N_7795,N_6498);
or U8409 (N_8409,N_7900,N_7180);
nor U8410 (N_8410,N_7251,N_7846);
or U8411 (N_8411,N_6677,N_7472);
nor U8412 (N_8412,N_6317,N_7882);
nand U8413 (N_8413,N_6419,N_6662);
or U8414 (N_8414,N_6235,N_6098);
nand U8415 (N_8415,N_6106,N_6454);
or U8416 (N_8416,N_6387,N_6546);
or U8417 (N_8417,N_6420,N_7229);
or U8418 (N_8418,N_7901,N_7316);
or U8419 (N_8419,N_6588,N_7220);
or U8420 (N_8420,N_7743,N_7605);
nor U8421 (N_8421,N_7293,N_6654);
and U8422 (N_8422,N_7144,N_7427);
or U8423 (N_8423,N_6804,N_7277);
or U8424 (N_8424,N_6995,N_7810);
or U8425 (N_8425,N_7044,N_7373);
and U8426 (N_8426,N_7333,N_6948);
nand U8427 (N_8427,N_7394,N_6221);
xor U8428 (N_8428,N_7678,N_6827);
nor U8429 (N_8429,N_7574,N_6232);
or U8430 (N_8430,N_6180,N_7254);
nor U8431 (N_8431,N_6403,N_7047);
and U8432 (N_8432,N_7792,N_6647);
or U8433 (N_8433,N_6667,N_7052);
xor U8434 (N_8434,N_6410,N_6297);
nand U8435 (N_8435,N_7149,N_6985);
nand U8436 (N_8436,N_7632,N_7153);
nand U8437 (N_8437,N_6316,N_6625);
nor U8438 (N_8438,N_7740,N_7957);
nand U8439 (N_8439,N_7192,N_7798);
or U8440 (N_8440,N_7423,N_7164);
nand U8441 (N_8441,N_6483,N_6656);
nor U8442 (N_8442,N_6134,N_6023);
nand U8443 (N_8443,N_6787,N_7750);
nor U8444 (N_8444,N_6699,N_7517);
nor U8445 (N_8445,N_7490,N_7715);
and U8446 (N_8446,N_6865,N_6124);
nand U8447 (N_8447,N_6989,N_7772);
and U8448 (N_8448,N_6145,N_7684);
nor U8449 (N_8449,N_7797,N_7387);
nand U8450 (N_8450,N_7223,N_7347);
and U8451 (N_8451,N_6190,N_6716);
or U8452 (N_8452,N_6530,N_7372);
or U8453 (N_8453,N_7979,N_6136);
xor U8454 (N_8454,N_7237,N_7300);
nor U8455 (N_8455,N_7935,N_7508);
nand U8456 (N_8456,N_7943,N_6543);
nand U8457 (N_8457,N_7906,N_6158);
or U8458 (N_8458,N_6868,N_6085);
xor U8459 (N_8459,N_6672,N_7956);
nand U8460 (N_8460,N_7198,N_7161);
nor U8461 (N_8461,N_7185,N_6595);
or U8462 (N_8462,N_6983,N_6414);
and U8463 (N_8463,N_6193,N_6904);
or U8464 (N_8464,N_6641,N_6634);
or U8465 (N_8465,N_7499,N_7441);
or U8466 (N_8466,N_6824,N_6857);
nand U8467 (N_8467,N_7038,N_7832);
or U8468 (N_8468,N_6888,N_7103);
or U8469 (N_8469,N_6674,N_7749);
nor U8470 (N_8470,N_7773,N_6506);
nor U8471 (N_8471,N_7581,N_6440);
nand U8472 (N_8472,N_7032,N_7207);
nand U8473 (N_8473,N_7748,N_7661);
nand U8474 (N_8474,N_7686,N_7118);
or U8475 (N_8475,N_7983,N_7121);
or U8476 (N_8476,N_7023,N_7580);
and U8477 (N_8477,N_7950,N_7879);
nor U8478 (N_8478,N_6390,N_6313);
nor U8479 (N_8479,N_7367,N_7195);
nand U8480 (N_8480,N_7063,N_6120);
xnor U8481 (N_8481,N_6931,N_6731);
nand U8482 (N_8482,N_6178,N_6129);
xnor U8483 (N_8483,N_6162,N_6968);
nand U8484 (N_8484,N_6921,N_6377);
or U8485 (N_8485,N_6692,N_7480);
and U8486 (N_8486,N_6110,N_6844);
xor U8487 (N_8487,N_7654,N_7619);
nor U8488 (N_8488,N_6808,N_6205);
nand U8489 (N_8489,N_6270,N_7839);
or U8490 (N_8490,N_7775,N_7240);
and U8491 (N_8491,N_6932,N_6349);
or U8492 (N_8492,N_7949,N_7018);
nor U8493 (N_8493,N_6342,N_6734);
nand U8494 (N_8494,N_6389,N_7170);
or U8495 (N_8495,N_7082,N_7497);
nor U8496 (N_8496,N_6521,N_7547);
and U8497 (N_8497,N_6760,N_7171);
or U8498 (N_8498,N_6616,N_6864);
xor U8499 (N_8499,N_6779,N_7104);
or U8500 (N_8500,N_7486,N_6225);
nor U8501 (N_8501,N_6744,N_7226);
nor U8502 (N_8502,N_6552,N_6101);
and U8503 (N_8503,N_6160,N_7346);
and U8504 (N_8504,N_7612,N_6360);
and U8505 (N_8505,N_6531,N_7145);
xnor U8506 (N_8506,N_7572,N_6381);
or U8507 (N_8507,N_7603,N_7916);
or U8508 (N_8508,N_6339,N_7827);
nor U8509 (N_8509,N_6567,N_7155);
nand U8510 (N_8510,N_7526,N_6362);
and U8511 (N_8511,N_7650,N_6347);
or U8512 (N_8512,N_7907,N_7883);
or U8513 (N_8513,N_7553,N_6336);
nor U8514 (N_8514,N_6444,N_6488);
nor U8515 (N_8515,N_6596,N_6218);
and U8516 (N_8516,N_7944,N_7847);
nor U8517 (N_8517,N_6346,N_6131);
nor U8518 (N_8518,N_6577,N_6453);
or U8519 (N_8519,N_6639,N_7964);
xor U8520 (N_8520,N_7699,N_7732);
and U8521 (N_8521,N_6704,N_6021);
or U8522 (N_8522,N_6818,N_7837);
or U8523 (N_8523,N_7451,N_6833);
or U8524 (N_8524,N_6526,N_7356);
or U8525 (N_8525,N_7418,N_6424);
xnor U8526 (N_8526,N_6055,N_7459);
and U8527 (N_8527,N_7162,N_7437);
or U8528 (N_8528,N_6282,N_7233);
xor U8529 (N_8529,N_7033,N_7342);
or U8530 (N_8530,N_6534,N_6111);
nand U8531 (N_8531,N_7201,N_7376);
or U8532 (N_8532,N_7269,N_7628);
and U8533 (N_8533,N_6179,N_6038);
nor U8534 (N_8534,N_7303,N_7928);
nor U8535 (N_8535,N_6263,N_7842);
and U8536 (N_8536,N_6581,N_7942);
or U8537 (N_8537,N_7858,N_6006);
nor U8538 (N_8538,N_7566,N_7456);
nand U8539 (N_8539,N_6069,N_6433);
and U8540 (N_8540,N_6015,N_6118);
xnor U8541 (N_8541,N_6814,N_6626);
or U8542 (N_8542,N_7353,N_6726);
or U8543 (N_8543,N_6460,N_6154);
nand U8544 (N_8544,N_7878,N_7005);
nand U8545 (N_8545,N_6077,N_6815);
nand U8546 (N_8546,N_6905,N_6843);
nor U8547 (N_8547,N_6568,N_7774);
nand U8548 (N_8548,N_7478,N_6946);
or U8549 (N_8549,N_7120,N_6099);
nor U8550 (N_8550,N_6503,N_7945);
or U8551 (N_8551,N_7193,N_6899);
or U8552 (N_8552,N_6482,N_6034);
or U8553 (N_8553,N_6369,N_6096);
nor U8554 (N_8554,N_6593,N_6871);
nor U8555 (N_8555,N_6786,N_7175);
nand U8556 (N_8556,N_7722,N_7784);
nand U8557 (N_8557,N_7727,N_6954);
or U8558 (N_8558,N_6719,N_6025);
and U8559 (N_8559,N_6289,N_7601);
or U8560 (N_8560,N_6246,N_6691);
xnor U8561 (N_8561,N_6512,N_7941);
xnor U8562 (N_8562,N_7301,N_6234);
nand U8563 (N_8563,N_7452,N_7543);
nand U8564 (N_8564,N_6294,N_6060);
nand U8565 (N_8565,N_7440,N_7545);
or U8566 (N_8566,N_6432,N_7729);
nor U8567 (N_8567,N_6515,N_7368);
nor U8568 (N_8568,N_6771,N_7213);
and U8569 (N_8569,N_6615,N_6849);
or U8570 (N_8570,N_6991,N_7664);
nor U8571 (N_8571,N_6777,N_6750);
nand U8572 (N_8572,N_7996,N_7760);
and U8573 (N_8573,N_7039,N_7886);
and U8574 (N_8574,N_6638,N_7336);
nor U8575 (N_8575,N_7482,N_7779);
or U8576 (N_8576,N_6150,N_7785);
or U8577 (N_8577,N_6970,N_6284);
nor U8578 (N_8578,N_7766,N_6757);
nand U8579 (N_8579,N_6712,N_7133);
and U8580 (N_8580,N_6423,N_6992);
and U8581 (N_8581,N_7111,N_6259);
or U8582 (N_8582,N_6019,N_7863);
and U8583 (N_8583,N_7947,N_6911);
or U8584 (N_8584,N_7304,N_7594);
nor U8585 (N_8585,N_6789,N_7895);
nand U8586 (N_8586,N_6563,N_7851);
xnor U8587 (N_8587,N_6366,N_7621);
nand U8588 (N_8588,N_7244,N_6386);
or U8589 (N_8589,N_7436,N_7550);
xnor U8590 (N_8590,N_7789,N_7282);
nand U8591 (N_8591,N_6876,N_6908);
or U8592 (N_8592,N_6418,N_6093);
nand U8593 (N_8593,N_7495,N_7142);
and U8594 (N_8594,N_7136,N_7794);
or U8595 (N_8595,N_7800,N_7477);
or U8596 (N_8596,N_6068,N_6445);
nand U8597 (N_8597,N_6436,N_6533);
and U8598 (N_8598,N_7159,N_7519);
and U8599 (N_8599,N_6308,N_6306);
nand U8600 (N_8600,N_6651,N_6944);
nand U8601 (N_8601,N_6210,N_7531);
or U8602 (N_8602,N_7406,N_6016);
xor U8603 (N_8603,N_6072,N_7380);
and U8604 (N_8604,N_6630,N_7359);
nor U8605 (N_8605,N_7597,N_6107);
nand U8606 (N_8606,N_6661,N_7412);
and U8607 (N_8607,N_6268,N_7620);
and U8608 (N_8608,N_7496,N_7354);
nand U8609 (N_8609,N_6227,N_6164);
or U8610 (N_8610,N_6800,N_7174);
nand U8611 (N_8611,N_6852,N_6913);
or U8612 (N_8612,N_6614,N_7966);
or U8613 (N_8613,N_6076,N_7876);
nand U8614 (N_8614,N_6583,N_7559);
nor U8615 (N_8615,N_6326,N_7657);
or U8616 (N_8616,N_6175,N_7972);
or U8617 (N_8617,N_7712,N_7068);
nand U8618 (N_8618,N_7361,N_6657);
or U8619 (N_8619,N_7385,N_7542);
or U8620 (N_8620,N_7676,N_7348);
or U8621 (N_8621,N_7578,N_6895);
nor U8622 (N_8622,N_7314,N_7977);
and U8623 (N_8623,N_6256,N_6759);
nor U8624 (N_8624,N_6951,N_7755);
nand U8625 (N_8625,N_7006,N_6825);
and U8626 (N_8626,N_6850,N_7383);
and U8627 (N_8627,N_6891,N_7518);
nor U8628 (N_8628,N_7020,N_7769);
or U8629 (N_8629,N_6901,N_7275);
nor U8630 (N_8630,N_6937,N_6589);
nand U8631 (N_8631,N_7146,N_7570);
and U8632 (N_8632,N_6949,N_6962);
nor U8633 (N_8633,N_7776,N_7395);
and U8634 (N_8634,N_7582,N_7668);
nand U8635 (N_8635,N_7968,N_6401);
nand U8636 (N_8636,N_7634,N_7871);
or U8637 (N_8637,N_7417,N_6688);
or U8638 (N_8638,N_7869,N_7329);
nor U8639 (N_8639,N_7805,N_7040);
or U8640 (N_8640,N_7951,N_6659);
and U8641 (N_8641,N_6007,N_6749);
and U8642 (N_8642,N_7043,N_6706);
and U8643 (N_8643,N_6663,N_7439);
xnor U8644 (N_8644,N_6507,N_7232);
nor U8645 (N_8645,N_6045,N_7177);
nor U8646 (N_8646,N_7163,N_7262);
nand U8647 (N_8647,N_7652,N_6050);
or U8648 (N_8648,N_7631,N_7682);
or U8649 (N_8649,N_7698,N_7868);
nor U8650 (N_8650,N_7070,N_6558);
nor U8651 (N_8651,N_7530,N_7788);
and U8652 (N_8652,N_6014,N_6048);
or U8653 (N_8653,N_6715,N_6074);
or U8654 (N_8654,N_6115,N_6705);
and U8655 (N_8655,N_7991,N_6935);
and U8656 (N_8656,N_6658,N_6443);
nor U8657 (N_8657,N_6653,N_6955);
or U8658 (N_8658,N_6837,N_7100);
or U8659 (N_8659,N_7168,N_6431);
and U8660 (N_8660,N_7374,N_6571);
and U8661 (N_8661,N_6520,N_7057);
or U8662 (N_8662,N_7672,N_7644);
or U8663 (N_8663,N_6318,N_6540);
or U8664 (N_8664,N_7117,N_6157);
nand U8665 (N_8665,N_6413,N_6287);
xor U8666 (N_8666,N_6971,N_6126);
nor U8667 (N_8667,N_7625,N_6201);
nor U8668 (N_8668,N_6353,N_6713);
and U8669 (N_8669,N_6902,N_7455);
nand U8670 (N_8670,N_6550,N_6695);
nand U8671 (N_8671,N_6670,N_6928);
nand U8672 (N_8672,N_6729,N_7260);
nor U8673 (N_8673,N_7861,N_7266);
nor U8674 (N_8674,N_7533,N_6479);
nor U8675 (N_8675,N_6576,N_6838);
nor U8676 (N_8676,N_7585,N_6312);
nor U8677 (N_8677,N_7635,N_7782);
nand U8678 (N_8678,N_7905,N_6059);
and U8679 (N_8679,N_7485,N_7338);
xnor U8680 (N_8680,N_6676,N_7997);
and U8681 (N_8681,N_6733,N_7833);
nand U8682 (N_8682,N_7224,N_7926);
or U8683 (N_8683,N_6368,N_7552);
nor U8684 (N_8684,N_6724,N_6628);
or U8685 (N_8685,N_7904,N_6088);
nand U8686 (N_8686,N_6878,N_6623);
xor U8687 (N_8687,N_6603,N_6694);
nor U8688 (N_8688,N_6030,N_7507);
and U8689 (N_8689,N_6344,N_6102);
or U8690 (N_8690,N_6003,N_7320);
and U8691 (N_8691,N_6226,N_6953);
and U8692 (N_8692,N_6541,N_7877);
nor U8693 (N_8693,N_6311,N_6884);
and U8694 (N_8694,N_6301,N_7148);
xnor U8695 (N_8695,N_7012,N_6939);
nand U8696 (N_8696,N_7257,N_6684);
nand U8697 (N_8697,N_6580,N_7296);
and U8698 (N_8698,N_7618,N_6140);
nor U8699 (N_8699,N_6972,N_7736);
xnor U8700 (N_8700,N_7974,N_7599);
nand U8701 (N_8701,N_6544,N_7319);
nand U8702 (N_8702,N_7617,N_6299);
nor U8703 (N_8703,N_7391,N_7577);
xnor U8704 (N_8704,N_6536,N_6372);
nor U8705 (N_8705,N_7369,N_6159);
nor U8706 (N_8706,N_7003,N_6751);
nor U8707 (N_8707,N_7821,N_7998);
or U8708 (N_8708,N_7209,N_6497);
nor U8709 (N_8709,N_7114,N_7045);
or U8710 (N_8710,N_7285,N_6548);
nor U8711 (N_8711,N_7924,N_7081);
nand U8712 (N_8712,N_6254,N_7129);
and U8713 (N_8713,N_6307,N_7724);
and U8714 (N_8714,N_6770,N_6447);
nand U8715 (N_8715,N_7575,N_7764);
nor U8716 (N_8716,N_7616,N_7008);
or U8717 (N_8717,N_6123,N_7680);
and U8718 (N_8718,N_7328,N_7639);
nor U8719 (N_8719,N_7402,N_6671);
nor U8720 (N_8720,N_7438,N_6756);
and U8721 (N_8721,N_6384,N_7349);
and U8722 (N_8722,N_6791,N_6345);
or U8723 (N_8723,N_6528,N_6762);
and U8724 (N_8724,N_6217,N_6957);
and U8725 (N_8725,N_7651,N_6870);
nor U8726 (N_8726,N_7731,N_6156);
xnor U8727 (N_8727,N_6796,N_6354);
nor U8728 (N_8728,N_6042,N_7143);
nand U8729 (N_8729,N_6885,N_7066);
and U8730 (N_8730,N_7091,N_7037);
or U8731 (N_8731,N_7568,N_6645);
and U8732 (N_8732,N_6936,N_6116);
nor U8733 (N_8733,N_6065,N_6032);
xor U8734 (N_8734,N_7709,N_6303);
or U8735 (N_8735,N_7999,N_7524);
nand U8736 (N_8736,N_6200,N_7067);
nor U8737 (N_8737,N_6889,N_7733);
nand U8738 (N_8738,N_7993,N_7758);
xnor U8739 (N_8739,N_6591,N_6893);
or U8740 (N_8740,N_7054,N_7449);
and U8741 (N_8741,N_7875,N_6601);
nand U8742 (N_8742,N_6480,N_7930);
or U8743 (N_8743,N_6938,N_7511);
or U8744 (N_8744,N_7830,N_6755);
nor U8745 (N_8745,N_6137,N_7473);
or U8746 (N_8746,N_7985,N_6293);
xnor U8747 (N_8747,N_7399,N_6338);
or U8748 (N_8748,N_7194,N_6689);
nand U8749 (N_8749,N_7022,N_7311);
or U8750 (N_8750,N_6161,N_7169);
xnor U8751 (N_8751,N_6185,N_6171);
nand U8752 (N_8752,N_7225,N_6400);
or U8753 (N_8753,N_6832,N_6279);
or U8754 (N_8754,N_7919,N_7889);
and U8755 (N_8755,N_7633,N_7801);
nor U8756 (N_8756,N_7777,N_7962);
nand U8757 (N_8757,N_6629,N_6806);
nand U8758 (N_8758,N_6519,N_7952);
nand U8759 (N_8759,N_7948,N_7596);
and U8760 (N_8760,N_6690,N_6216);
nand U8761 (N_8761,N_6051,N_7292);
and U8762 (N_8762,N_6192,N_6621);
nor U8763 (N_8763,N_6170,N_6836);
nand U8764 (N_8764,N_7312,N_7636);
and U8765 (N_8765,N_6801,N_6527);
and U8766 (N_8766,N_6778,N_6062);
and U8767 (N_8767,N_6780,N_7866);
and U8768 (N_8768,N_6489,N_7965);
xnor U8769 (N_8769,N_6090,N_7072);
or U8770 (N_8770,N_7525,N_6363);
and U8771 (N_8771,N_6407,N_7953);
xnor U8772 (N_8772,N_6518,N_6117);
nand U8773 (N_8773,N_7845,N_6351);
and U8774 (N_8774,N_7466,N_7462);
and U8775 (N_8775,N_7231,N_6635);
nand U8776 (N_8776,N_6495,N_7555);
and U8777 (N_8777,N_7564,N_7126);
nand U8778 (N_8778,N_7165,N_7152);
and U8779 (N_8779,N_7228,N_7278);
or U8780 (N_8780,N_6084,N_6319);
xnor U8781 (N_8781,N_6965,N_7909);
or U8782 (N_8782,N_7390,N_7719);
nand U8783 (N_8783,N_6024,N_7265);
and U8784 (N_8784,N_7468,N_6668);
nand U8785 (N_8785,N_7060,N_7960);
and U8786 (N_8786,N_7967,N_6203);
or U8787 (N_8787,N_7744,N_6172);
nor U8788 (N_8788,N_6382,N_6693);
nand U8789 (N_8789,N_7092,N_7609);
or U8790 (N_8790,N_6996,N_6341);
nor U8791 (N_8791,N_6189,N_7829);
and U8792 (N_8792,N_7130,N_7085);
xor U8793 (N_8793,N_6883,N_7534);
nor U8794 (N_8794,N_6861,N_7593);
xor U8795 (N_8795,N_6920,N_7902);
nor U8796 (N_8796,N_7419,N_7826);
xor U8797 (N_8797,N_7366,N_7448);
nand U8798 (N_8798,N_7004,N_7378);
and U8799 (N_8799,N_7400,N_6011);
and U8800 (N_8800,N_6405,N_6125);
xnor U8801 (N_8801,N_7414,N_6795);
nand U8802 (N_8802,N_7854,N_7540);
nor U8803 (N_8803,N_6743,N_6959);
or U8804 (N_8804,N_6375,N_7500);
nand U8805 (N_8805,N_6114,N_6380);
or U8806 (N_8806,N_6923,N_6673);
or U8807 (N_8807,N_6510,N_6269);
or U8808 (N_8808,N_7716,N_7610);
nand U8809 (N_8809,N_7538,N_6421);
and U8810 (N_8810,N_7557,N_7931);
xor U8811 (N_8811,N_7649,N_6169);
or U8812 (N_8812,N_7856,N_6697);
nand U8813 (N_8813,N_7110,N_6820);
and U8814 (N_8814,N_7726,N_6675);
and U8815 (N_8815,N_7990,N_6005);
nand U8816 (N_8816,N_7933,N_7614);
nor U8817 (N_8817,N_7704,N_7150);
nand U8818 (N_8818,N_6646,N_6044);
and U8819 (N_8819,N_7137,N_7214);
nand U8820 (N_8820,N_7212,N_6841);
xnor U8821 (N_8821,N_6334,N_6566);
or U8822 (N_8822,N_6429,N_6723);
xnor U8823 (N_8823,N_6370,N_6437);
and U8824 (N_8824,N_6710,N_7288);
and U8825 (N_8825,N_6215,N_6809);
or U8826 (N_8826,N_7561,N_7410);
or U8827 (N_8827,N_6455,N_7707);
and U8828 (N_8828,N_6958,N_7645);
nand U8829 (N_8829,N_6073,N_7893);
nand U8830 (N_8830,N_7992,N_6969);
xor U8831 (N_8831,N_6829,N_7371);
nor U8832 (N_8832,N_7424,N_7335);
nand U8833 (N_8833,N_7741,N_6585);
xor U8834 (N_8834,N_6964,N_6337);
and U8835 (N_8835,N_7884,N_7973);
and U8836 (N_8836,N_7310,N_6867);
nand U8837 (N_8837,N_7925,N_6754);
xnor U8838 (N_8838,N_6302,N_6660);
nand U8839 (N_8839,N_6830,N_6209);
and U8840 (N_8840,N_6357,N_6978);
or U8841 (N_8841,N_6586,N_6622);
or U8842 (N_8842,N_6043,N_7075);
and U8843 (N_8843,N_6467,N_7026);
and U8844 (N_8844,N_7355,N_6516);
and U8845 (N_8845,N_7637,N_7167);
and U8846 (N_8846,N_7362,N_6028);
nor U8847 (N_8847,N_7590,N_6379);
nand U8848 (N_8848,N_6508,N_7791);
and U8849 (N_8849,N_6828,N_6275);
and U8850 (N_8850,N_6742,N_6041);
and U8851 (N_8851,N_7196,N_7313);
nand U8852 (N_8852,N_7655,N_7446);
or U8853 (N_8853,N_6727,N_6211);
nor U8854 (N_8854,N_7049,N_7961);
nor U8855 (N_8855,N_6802,N_7056);
nand U8856 (N_8856,N_6206,N_7730);
or U8857 (N_8857,N_7802,N_6562);
nor U8858 (N_8858,N_6792,N_7793);
nor U8859 (N_8859,N_6439,N_7505);
or U8860 (N_8860,N_6087,N_7430);
nand U8861 (N_8861,N_7308,N_6877);
or U8862 (N_8862,N_7344,N_7683);
nor U8863 (N_8863,N_7921,N_7393);
nor U8864 (N_8864,N_7523,N_7781);
nand U8865 (N_8865,N_6916,N_6807);
nor U8866 (N_8866,N_6785,N_6265);
and U8867 (N_8867,N_6490,N_7160);
and U8868 (N_8868,N_7442,N_7379);
or U8869 (N_8869,N_7340,N_6933);
or U8870 (N_8870,N_6529,N_7280);
and U8871 (N_8871,N_7569,N_6165);
xnor U8872 (N_8872,N_7179,N_7243);
nor U8873 (N_8873,N_6554,N_6194);
nor U8874 (N_8874,N_7299,N_7849);
and U8875 (N_8875,N_6143,N_6475);
nor U8876 (N_8876,N_6854,N_7528);
or U8877 (N_8877,N_7622,N_7088);
nor U8878 (N_8878,N_6220,N_6542);
nor U8879 (N_8879,N_7116,N_6609);
nand U8880 (N_8880,N_7183,N_6472);
or U8881 (N_8881,N_7426,N_6416);
and U8882 (N_8882,N_7809,N_6974);
and U8883 (N_8883,N_6572,N_6406);
or U8884 (N_8884,N_6053,N_6584);
nand U8885 (N_8885,N_7959,N_6355);
nand U8886 (N_8886,N_7720,N_6272);
nor U8887 (N_8887,N_6819,N_6702);
nand U8888 (N_8888,N_7807,N_6187);
and U8889 (N_8889,N_6168,N_7685);
nor U8890 (N_8890,N_7105,N_7458);
nor U8891 (N_8891,N_7890,N_6058);
and U8892 (N_8892,N_7549,N_6547);
and U8893 (N_8893,N_7874,N_6305);
or U8894 (N_8894,N_7447,N_6276);
xnor U8895 (N_8895,N_6009,N_7504);
xnor U8896 (N_8896,N_7218,N_7855);
and U8897 (N_8897,N_7804,N_7604);
or U8898 (N_8898,N_6153,N_7246);
or U8899 (N_8899,N_6999,N_6329);
nand U8900 (N_8900,N_7494,N_7838);
or U8901 (N_8901,N_7450,N_6890);
and U8902 (N_8902,N_6767,N_6752);
nor U8903 (N_8903,N_6665,N_7738);
or U8904 (N_8904,N_6383,N_7475);
nor U8905 (N_8905,N_7648,N_6417);
or U8906 (N_8906,N_7790,N_7659);
and U8907 (N_8907,N_6267,N_7087);
nor U8908 (N_8908,N_6070,N_7454);
or U8909 (N_8909,N_7677,N_6404);
nand U8910 (N_8910,N_7514,N_6310);
nor U8911 (N_8911,N_6681,N_6146);
nand U8912 (N_8912,N_7823,N_7817);
nor U8913 (N_8913,N_6988,N_6470);
nand U8914 (N_8914,N_7536,N_6608);
nand U8915 (N_8915,N_7139,N_6020);
and U8916 (N_8916,N_7078,N_6873);
nand U8917 (N_8917,N_6997,N_7001);
or U8918 (N_8918,N_7375,N_7579);
nor U8919 (N_8919,N_7267,N_6950);
or U8920 (N_8920,N_7522,N_6128);
and U8921 (N_8921,N_6243,N_7264);
or U8922 (N_8922,N_7274,N_7853);
nor U8923 (N_8923,N_7615,N_6422);
and U8924 (N_8924,N_6435,N_6592);
and U8925 (N_8925,N_7813,N_7287);
or U8926 (N_8926,N_6207,N_7062);
or U8927 (N_8927,N_6141,N_6402);
nor U8928 (N_8928,N_6793,N_7914);
and U8929 (N_8929,N_7172,N_6290);
xnor U8930 (N_8930,N_7377,N_6323);
or U8931 (N_8931,N_7892,N_6425);
or U8932 (N_8932,N_7911,N_6648);
nand U8933 (N_8933,N_6763,N_6000);
xnor U8934 (N_8934,N_7691,N_6298);
nand U8935 (N_8935,N_6564,N_6790);
or U8936 (N_8936,N_7841,N_7470);
and U8937 (N_8937,N_6722,N_6487);
or U8938 (N_8938,N_6018,N_6144);
and U8939 (N_8939,N_6872,N_6365);
and U8940 (N_8940,N_7759,N_7556);
or U8941 (N_8941,N_6773,N_6894);
nand U8942 (N_8942,N_7754,N_7647);
nand U8943 (N_8943,N_6941,N_7156);
or U8944 (N_8944,N_7330,N_6033);
nor U8945 (N_8945,N_6797,N_6758);
nand U8946 (N_8946,N_6917,N_7498);
and U8947 (N_8947,N_7811,N_7445);
xnor U8948 (N_8948,N_7276,N_6919);
nand U8949 (N_8949,N_7096,N_6869);
and U8950 (N_8950,N_6378,N_7253);
or U8951 (N_8951,N_6138,N_6909);
nor U8952 (N_8952,N_6606,N_7061);
nand U8953 (N_8953,N_7520,N_6376);
nand U8954 (N_8954,N_6314,N_7431);
nand U8955 (N_8955,N_6385,N_6597);
nand U8956 (N_8956,N_7663,N_6039);
nor U8957 (N_8957,N_7250,N_7548);
and U8958 (N_8958,N_7248,N_6961);
and U8959 (N_8959,N_7469,N_7041);
nand U8960 (N_8960,N_6371,N_7421);
nand U8961 (N_8961,N_6208,N_6249);
nor U8962 (N_8962,N_7115,N_6897);
nor U8963 (N_8963,N_6446,N_6359);
nor U8964 (N_8964,N_7184,N_7980);
and U8965 (N_8965,N_6500,N_6732);
nand U8966 (N_8966,N_6537,N_7692);
nor U8967 (N_8967,N_6223,N_6271);
and U8968 (N_8968,N_6253,N_7382);
xnor U8969 (N_8969,N_6196,N_7492);
and U8970 (N_8970,N_7432,N_7859);
xor U8971 (N_8971,N_7221,N_6509);
nand U8972 (N_8972,N_6399,N_6522);
nand U8973 (N_8973,N_6130,N_7588);
or U8974 (N_8974,N_6100,N_7955);
nand U8975 (N_8975,N_6083,N_6631);
or U8976 (N_8976,N_7502,N_7491);
nand U8977 (N_8977,N_7106,N_6679);
and U8978 (N_8978,N_6525,N_7216);
nand U8979 (N_8979,N_6918,N_6798);
nor U8980 (N_8980,N_6898,N_6906);
and U8981 (N_8981,N_7600,N_7768);
nor U8982 (N_8982,N_7987,N_6255);
nor U8983 (N_8983,N_7640,N_7204);
nor U8984 (N_8984,N_6859,N_7560);
nand U8985 (N_8985,N_7268,N_6739);
or U8986 (N_8986,N_7613,N_7567);
or U8987 (N_8987,N_7219,N_7923);
or U8988 (N_8988,N_6320,N_6199);
and U8989 (N_8989,N_6617,N_7321);
nand U8990 (N_8990,N_7050,N_7840);
or U8991 (N_8991,N_6356,N_6481);
nor U8992 (N_8992,N_7700,N_6598);
and U8993 (N_8993,N_6880,N_6026);
nor U8994 (N_8994,N_6451,N_6266);
nor U8995 (N_8995,N_6766,N_6474);
or U8996 (N_8996,N_7510,N_7396);
nor U8997 (N_8997,N_7173,N_7503);
nand U8998 (N_8998,N_7122,N_7318);
and U8999 (N_8999,N_6328,N_6122);
nor U9000 (N_9000,N_7842,N_7911);
xnor U9001 (N_9001,N_7729,N_7845);
or U9002 (N_9002,N_7281,N_7299);
or U9003 (N_9003,N_6905,N_7230);
or U9004 (N_9004,N_7462,N_7734);
and U9005 (N_9005,N_7903,N_6434);
nor U9006 (N_9006,N_6610,N_7635);
nor U9007 (N_9007,N_6708,N_7042);
nand U9008 (N_9008,N_6509,N_6211);
nor U9009 (N_9009,N_6664,N_7834);
nand U9010 (N_9010,N_6285,N_6066);
nand U9011 (N_9011,N_6740,N_6968);
and U9012 (N_9012,N_7757,N_7791);
or U9013 (N_9013,N_7648,N_6129);
and U9014 (N_9014,N_6185,N_6966);
nand U9015 (N_9015,N_7046,N_6810);
or U9016 (N_9016,N_6930,N_6407);
or U9017 (N_9017,N_7236,N_6050);
nor U9018 (N_9018,N_7544,N_7587);
nor U9019 (N_9019,N_7861,N_7011);
xnor U9020 (N_9020,N_6843,N_6682);
or U9021 (N_9021,N_6787,N_7264);
nand U9022 (N_9022,N_6907,N_7879);
xnor U9023 (N_9023,N_6124,N_6972);
nand U9024 (N_9024,N_6359,N_6183);
and U9025 (N_9025,N_7889,N_6357);
nor U9026 (N_9026,N_6502,N_6612);
and U9027 (N_9027,N_7164,N_7331);
nor U9028 (N_9028,N_6625,N_6902);
and U9029 (N_9029,N_7091,N_7426);
nand U9030 (N_9030,N_7735,N_7454);
nor U9031 (N_9031,N_6776,N_6041);
nor U9032 (N_9032,N_7950,N_6550);
and U9033 (N_9033,N_7252,N_7499);
nor U9034 (N_9034,N_7261,N_6820);
and U9035 (N_9035,N_6971,N_6853);
or U9036 (N_9036,N_6334,N_7856);
nand U9037 (N_9037,N_7421,N_7338);
and U9038 (N_9038,N_6419,N_6225);
nand U9039 (N_9039,N_7263,N_7212);
and U9040 (N_9040,N_6265,N_7141);
nand U9041 (N_9041,N_7088,N_6751);
nor U9042 (N_9042,N_7712,N_6140);
nor U9043 (N_9043,N_7088,N_7452);
nor U9044 (N_9044,N_7569,N_6553);
or U9045 (N_9045,N_6976,N_7995);
nand U9046 (N_9046,N_6608,N_7020);
nor U9047 (N_9047,N_6304,N_6518);
nor U9048 (N_9048,N_6904,N_6726);
xor U9049 (N_9049,N_6101,N_6311);
or U9050 (N_9050,N_7880,N_6232);
and U9051 (N_9051,N_7839,N_6022);
and U9052 (N_9052,N_6734,N_7372);
and U9053 (N_9053,N_7534,N_7326);
or U9054 (N_9054,N_7719,N_7825);
or U9055 (N_9055,N_7635,N_6601);
nand U9056 (N_9056,N_6316,N_6577);
or U9057 (N_9057,N_7513,N_7939);
or U9058 (N_9058,N_6731,N_6275);
or U9059 (N_9059,N_6848,N_6794);
and U9060 (N_9060,N_6620,N_6277);
and U9061 (N_9061,N_6427,N_6843);
nor U9062 (N_9062,N_6929,N_6736);
nand U9063 (N_9063,N_6484,N_6540);
nor U9064 (N_9064,N_6732,N_6070);
or U9065 (N_9065,N_6153,N_6246);
and U9066 (N_9066,N_7138,N_6320);
and U9067 (N_9067,N_6901,N_7842);
nor U9068 (N_9068,N_6944,N_6879);
nand U9069 (N_9069,N_7173,N_6785);
and U9070 (N_9070,N_7991,N_6439);
or U9071 (N_9071,N_6995,N_7669);
nand U9072 (N_9072,N_7712,N_7370);
or U9073 (N_9073,N_7834,N_6186);
nor U9074 (N_9074,N_7264,N_6521);
or U9075 (N_9075,N_7650,N_6414);
nor U9076 (N_9076,N_7014,N_6611);
nand U9077 (N_9077,N_6992,N_6148);
and U9078 (N_9078,N_6222,N_6361);
nand U9079 (N_9079,N_7222,N_7602);
and U9080 (N_9080,N_7467,N_7103);
nand U9081 (N_9081,N_7555,N_6026);
nor U9082 (N_9082,N_6222,N_6132);
or U9083 (N_9083,N_7373,N_6748);
or U9084 (N_9084,N_6696,N_7194);
nand U9085 (N_9085,N_6846,N_7570);
nand U9086 (N_9086,N_6963,N_7144);
and U9087 (N_9087,N_6310,N_6078);
nand U9088 (N_9088,N_6757,N_7931);
or U9089 (N_9089,N_7705,N_6738);
and U9090 (N_9090,N_7559,N_6353);
or U9091 (N_9091,N_7536,N_7811);
or U9092 (N_9092,N_6931,N_6074);
and U9093 (N_9093,N_7308,N_6458);
and U9094 (N_9094,N_7989,N_7470);
nor U9095 (N_9095,N_6331,N_6014);
or U9096 (N_9096,N_7474,N_7909);
or U9097 (N_9097,N_7853,N_7510);
nor U9098 (N_9098,N_7804,N_6176);
nor U9099 (N_9099,N_7886,N_7129);
nand U9100 (N_9100,N_7731,N_6517);
nor U9101 (N_9101,N_7143,N_6011);
and U9102 (N_9102,N_6738,N_6424);
xor U9103 (N_9103,N_6520,N_6313);
nor U9104 (N_9104,N_6479,N_6978);
nand U9105 (N_9105,N_7113,N_6574);
and U9106 (N_9106,N_6033,N_6242);
or U9107 (N_9107,N_7158,N_6075);
xnor U9108 (N_9108,N_6761,N_7312);
nand U9109 (N_9109,N_6450,N_6714);
nand U9110 (N_9110,N_7662,N_7003);
xnor U9111 (N_9111,N_6478,N_7036);
nor U9112 (N_9112,N_6199,N_7140);
or U9113 (N_9113,N_7621,N_7618);
xnor U9114 (N_9114,N_6743,N_7802);
nor U9115 (N_9115,N_7075,N_6741);
and U9116 (N_9116,N_6579,N_7687);
nor U9117 (N_9117,N_6335,N_6387);
or U9118 (N_9118,N_7013,N_6180);
nor U9119 (N_9119,N_6277,N_7794);
or U9120 (N_9120,N_7589,N_7415);
or U9121 (N_9121,N_7463,N_6411);
or U9122 (N_9122,N_7127,N_7347);
nand U9123 (N_9123,N_6645,N_7871);
xnor U9124 (N_9124,N_7003,N_7854);
and U9125 (N_9125,N_7605,N_7695);
nor U9126 (N_9126,N_7881,N_7829);
and U9127 (N_9127,N_7190,N_7753);
or U9128 (N_9128,N_6090,N_6102);
or U9129 (N_9129,N_7794,N_7445);
and U9130 (N_9130,N_6316,N_6707);
and U9131 (N_9131,N_6873,N_7863);
or U9132 (N_9132,N_6904,N_6851);
nand U9133 (N_9133,N_6330,N_7116);
xnor U9134 (N_9134,N_7163,N_7790);
or U9135 (N_9135,N_6409,N_6607);
nor U9136 (N_9136,N_7644,N_6474);
xor U9137 (N_9137,N_6605,N_7650);
nand U9138 (N_9138,N_6687,N_7322);
nand U9139 (N_9139,N_6760,N_6456);
xor U9140 (N_9140,N_7979,N_7108);
nor U9141 (N_9141,N_6181,N_7934);
and U9142 (N_9142,N_6152,N_6697);
nor U9143 (N_9143,N_7803,N_7518);
or U9144 (N_9144,N_7187,N_6218);
or U9145 (N_9145,N_7128,N_6024);
nor U9146 (N_9146,N_7814,N_7959);
nand U9147 (N_9147,N_6625,N_7381);
or U9148 (N_9148,N_6935,N_7565);
or U9149 (N_9149,N_7145,N_6077);
nor U9150 (N_9150,N_7139,N_6321);
xor U9151 (N_9151,N_7956,N_6607);
nand U9152 (N_9152,N_6183,N_7860);
xor U9153 (N_9153,N_7126,N_6911);
nand U9154 (N_9154,N_7445,N_7974);
and U9155 (N_9155,N_7063,N_7844);
xor U9156 (N_9156,N_6451,N_7928);
xor U9157 (N_9157,N_7736,N_7397);
and U9158 (N_9158,N_6935,N_6012);
nor U9159 (N_9159,N_6796,N_7956);
nor U9160 (N_9160,N_6340,N_6553);
and U9161 (N_9161,N_6960,N_6584);
and U9162 (N_9162,N_7944,N_6234);
xor U9163 (N_9163,N_6696,N_6087);
nand U9164 (N_9164,N_6096,N_7351);
or U9165 (N_9165,N_6874,N_6848);
nor U9166 (N_9166,N_7072,N_6501);
nand U9167 (N_9167,N_6315,N_7148);
nand U9168 (N_9168,N_7951,N_7720);
or U9169 (N_9169,N_6077,N_7649);
nand U9170 (N_9170,N_6947,N_7548);
or U9171 (N_9171,N_6806,N_6728);
or U9172 (N_9172,N_6093,N_6277);
and U9173 (N_9173,N_6143,N_6478);
nor U9174 (N_9174,N_6180,N_7339);
nor U9175 (N_9175,N_7241,N_6773);
nand U9176 (N_9176,N_6399,N_6104);
and U9177 (N_9177,N_6455,N_6137);
nand U9178 (N_9178,N_7272,N_7061);
or U9179 (N_9179,N_6570,N_6630);
nor U9180 (N_9180,N_6710,N_7428);
xor U9181 (N_9181,N_6000,N_7856);
or U9182 (N_9182,N_6634,N_7660);
nor U9183 (N_9183,N_7758,N_7902);
nor U9184 (N_9184,N_7909,N_6931);
nand U9185 (N_9185,N_7728,N_6508);
or U9186 (N_9186,N_6524,N_7609);
and U9187 (N_9187,N_7679,N_6321);
nand U9188 (N_9188,N_6230,N_7794);
and U9189 (N_9189,N_6407,N_7339);
xor U9190 (N_9190,N_7244,N_7735);
or U9191 (N_9191,N_6643,N_6194);
and U9192 (N_9192,N_6279,N_6127);
nand U9193 (N_9193,N_7585,N_6393);
or U9194 (N_9194,N_6534,N_6265);
or U9195 (N_9195,N_6906,N_6740);
xnor U9196 (N_9196,N_7189,N_7263);
nand U9197 (N_9197,N_6040,N_7023);
or U9198 (N_9198,N_6473,N_6059);
and U9199 (N_9199,N_6677,N_7075);
and U9200 (N_9200,N_6355,N_7767);
nand U9201 (N_9201,N_7813,N_7414);
or U9202 (N_9202,N_6645,N_6316);
or U9203 (N_9203,N_7614,N_6538);
xor U9204 (N_9204,N_6120,N_7184);
and U9205 (N_9205,N_7765,N_6628);
nor U9206 (N_9206,N_6898,N_7548);
nor U9207 (N_9207,N_7082,N_6613);
or U9208 (N_9208,N_7053,N_6249);
or U9209 (N_9209,N_6732,N_7551);
and U9210 (N_9210,N_6158,N_6313);
or U9211 (N_9211,N_6160,N_6820);
or U9212 (N_9212,N_6838,N_6519);
or U9213 (N_9213,N_7078,N_6819);
or U9214 (N_9214,N_7311,N_6206);
xor U9215 (N_9215,N_6717,N_7432);
nand U9216 (N_9216,N_6485,N_7444);
xnor U9217 (N_9217,N_6654,N_6119);
nor U9218 (N_9218,N_6682,N_7352);
and U9219 (N_9219,N_7134,N_7234);
or U9220 (N_9220,N_7300,N_6662);
and U9221 (N_9221,N_7144,N_7685);
nand U9222 (N_9222,N_7391,N_6995);
nand U9223 (N_9223,N_7113,N_6694);
nor U9224 (N_9224,N_6387,N_6591);
nor U9225 (N_9225,N_7699,N_7501);
and U9226 (N_9226,N_7450,N_6491);
nand U9227 (N_9227,N_7677,N_7305);
nand U9228 (N_9228,N_7524,N_7980);
nand U9229 (N_9229,N_7416,N_6307);
xor U9230 (N_9230,N_7074,N_6344);
nand U9231 (N_9231,N_6128,N_7687);
nand U9232 (N_9232,N_6621,N_7203);
and U9233 (N_9233,N_6724,N_6959);
nor U9234 (N_9234,N_6176,N_6894);
nand U9235 (N_9235,N_7340,N_6869);
and U9236 (N_9236,N_6588,N_7140);
nand U9237 (N_9237,N_6168,N_6725);
xor U9238 (N_9238,N_7814,N_6245);
nor U9239 (N_9239,N_7345,N_7898);
or U9240 (N_9240,N_6780,N_6154);
xnor U9241 (N_9241,N_6727,N_7613);
and U9242 (N_9242,N_7385,N_7584);
or U9243 (N_9243,N_6099,N_6609);
or U9244 (N_9244,N_6935,N_6001);
xor U9245 (N_9245,N_6027,N_6314);
and U9246 (N_9246,N_7478,N_7185);
or U9247 (N_9247,N_7410,N_7317);
or U9248 (N_9248,N_7488,N_6971);
nand U9249 (N_9249,N_7286,N_6505);
or U9250 (N_9250,N_7787,N_6756);
nor U9251 (N_9251,N_6080,N_7769);
nand U9252 (N_9252,N_6757,N_6669);
or U9253 (N_9253,N_6103,N_6529);
nand U9254 (N_9254,N_7591,N_7835);
nor U9255 (N_9255,N_7122,N_7530);
nor U9256 (N_9256,N_6121,N_7215);
nor U9257 (N_9257,N_6238,N_7226);
nor U9258 (N_9258,N_6264,N_7368);
nand U9259 (N_9259,N_7638,N_7800);
or U9260 (N_9260,N_6111,N_7886);
and U9261 (N_9261,N_7611,N_7213);
nand U9262 (N_9262,N_6535,N_7298);
nor U9263 (N_9263,N_7977,N_6908);
nor U9264 (N_9264,N_6350,N_7020);
and U9265 (N_9265,N_7937,N_7627);
nand U9266 (N_9266,N_6167,N_6703);
or U9267 (N_9267,N_7716,N_6441);
and U9268 (N_9268,N_6086,N_7670);
nand U9269 (N_9269,N_6840,N_7881);
and U9270 (N_9270,N_6614,N_7095);
xnor U9271 (N_9271,N_7487,N_7626);
and U9272 (N_9272,N_6761,N_6244);
or U9273 (N_9273,N_6231,N_7781);
or U9274 (N_9274,N_6034,N_6092);
and U9275 (N_9275,N_6036,N_7452);
or U9276 (N_9276,N_7790,N_7241);
or U9277 (N_9277,N_7220,N_6138);
and U9278 (N_9278,N_6786,N_6144);
or U9279 (N_9279,N_7459,N_6628);
and U9280 (N_9280,N_7837,N_6413);
nor U9281 (N_9281,N_6229,N_7657);
and U9282 (N_9282,N_6700,N_6221);
nand U9283 (N_9283,N_7443,N_7539);
and U9284 (N_9284,N_7965,N_6383);
or U9285 (N_9285,N_7634,N_7887);
or U9286 (N_9286,N_6859,N_7461);
nor U9287 (N_9287,N_6725,N_6572);
xor U9288 (N_9288,N_7681,N_7307);
nand U9289 (N_9289,N_6823,N_7059);
nor U9290 (N_9290,N_7377,N_6684);
and U9291 (N_9291,N_6355,N_6136);
or U9292 (N_9292,N_6970,N_7017);
and U9293 (N_9293,N_6231,N_6798);
nor U9294 (N_9294,N_7359,N_7945);
nor U9295 (N_9295,N_7264,N_6320);
and U9296 (N_9296,N_7047,N_7954);
or U9297 (N_9297,N_7682,N_7132);
or U9298 (N_9298,N_7020,N_7168);
or U9299 (N_9299,N_7209,N_7608);
xnor U9300 (N_9300,N_7370,N_6783);
nor U9301 (N_9301,N_7067,N_6561);
and U9302 (N_9302,N_6341,N_7146);
nor U9303 (N_9303,N_7466,N_6508);
or U9304 (N_9304,N_6492,N_7961);
nand U9305 (N_9305,N_6730,N_6779);
nand U9306 (N_9306,N_7054,N_7326);
or U9307 (N_9307,N_6833,N_6692);
nand U9308 (N_9308,N_6440,N_7671);
nor U9309 (N_9309,N_7732,N_7447);
or U9310 (N_9310,N_7017,N_7303);
nand U9311 (N_9311,N_6324,N_7000);
and U9312 (N_9312,N_7237,N_7184);
xnor U9313 (N_9313,N_7859,N_6367);
or U9314 (N_9314,N_7952,N_7787);
nor U9315 (N_9315,N_6358,N_7700);
or U9316 (N_9316,N_6397,N_7574);
or U9317 (N_9317,N_6067,N_6672);
or U9318 (N_9318,N_6360,N_7974);
nand U9319 (N_9319,N_6414,N_6916);
nor U9320 (N_9320,N_6660,N_7891);
and U9321 (N_9321,N_6261,N_7303);
xnor U9322 (N_9322,N_6920,N_6438);
or U9323 (N_9323,N_7158,N_6029);
xnor U9324 (N_9324,N_6206,N_7786);
or U9325 (N_9325,N_6722,N_7170);
nand U9326 (N_9326,N_6390,N_7502);
or U9327 (N_9327,N_6287,N_6317);
or U9328 (N_9328,N_6286,N_6701);
or U9329 (N_9329,N_7448,N_6253);
nand U9330 (N_9330,N_7547,N_7884);
nand U9331 (N_9331,N_7801,N_6400);
nor U9332 (N_9332,N_6261,N_7378);
nor U9333 (N_9333,N_7759,N_7570);
or U9334 (N_9334,N_7188,N_6155);
and U9335 (N_9335,N_6513,N_7044);
or U9336 (N_9336,N_6574,N_6584);
nand U9337 (N_9337,N_7120,N_7650);
or U9338 (N_9338,N_7887,N_7039);
nor U9339 (N_9339,N_6501,N_6543);
nor U9340 (N_9340,N_6470,N_7255);
xor U9341 (N_9341,N_6188,N_6889);
or U9342 (N_9342,N_6563,N_7984);
nand U9343 (N_9343,N_7258,N_6494);
xor U9344 (N_9344,N_6387,N_7107);
xnor U9345 (N_9345,N_7840,N_7943);
xor U9346 (N_9346,N_6178,N_7979);
nor U9347 (N_9347,N_6594,N_7173);
and U9348 (N_9348,N_7872,N_7929);
or U9349 (N_9349,N_6640,N_7963);
nand U9350 (N_9350,N_6589,N_7012);
nand U9351 (N_9351,N_7362,N_6332);
or U9352 (N_9352,N_6076,N_6697);
nor U9353 (N_9353,N_6716,N_7331);
or U9354 (N_9354,N_6748,N_6669);
and U9355 (N_9355,N_6981,N_6282);
and U9356 (N_9356,N_6610,N_7926);
and U9357 (N_9357,N_7741,N_7864);
and U9358 (N_9358,N_6144,N_6865);
and U9359 (N_9359,N_6969,N_6459);
and U9360 (N_9360,N_6129,N_7703);
and U9361 (N_9361,N_7042,N_7306);
and U9362 (N_9362,N_7541,N_7048);
nor U9363 (N_9363,N_6610,N_7395);
and U9364 (N_9364,N_6735,N_7309);
or U9365 (N_9365,N_6843,N_7541);
and U9366 (N_9366,N_6040,N_6922);
and U9367 (N_9367,N_7012,N_7523);
nor U9368 (N_9368,N_7289,N_6970);
or U9369 (N_9369,N_6977,N_6874);
xor U9370 (N_9370,N_6883,N_7036);
and U9371 (N_9371,N_7924,N_7893);
and U9372 (N_9372,N_7846,N_6515);
and U9373 (N_9373,N_7185,N_7280);
nand U9374 (N_9374,N_6966,N_7293);
and U9375 (N_9375,N_6845,N_7183);
nand U9376 (N_9376,N_7018,N_6383);
xor U9377 (N_9377,N_7223,N_7055);
or U9378 (N_9378,N_7138,N_7001);
and U9379 (N_9379,N_7169,N_6043);
and U9380 (N_9380,N_6594,N_6085);
and U9381 (N_9381,N_6943,N_7031);
and U9382 (N_9382,N_6359,N_7072);
nor U9383 (N_9383,N_7171,N_6550);
and U9384 (N_9384,N_7245,N_6857);
or U9385 (N_9385,N_7379,N_6444);
nor U9386 (N_9386,N_7916,N_6795);
nor U9387 (N_9387,N_6180,N_6108);
xnor U9388 (N_9388,N_6762,N_7373);
nand U9389 (N_9389,N_6627,N_6070);
nand U9390 (N_9390,N_6381,N_7105);
nor U9391 (N_9391,N_6496,N_6363);
nor U9392 (N_9392,N_7941,N_6170);
or U9393 (N_9393,N_7565,N_7647);
nand U9394 (N_9394,N_6397,N_6562);
nor U9395 (N_9395,N_6920,N_6894);
and U9396 (N_9396,N_6913,N_6803);
nand U9397 (N_9397,N_6017,N_7781);
and U9398 (N_9398,N_7935,N_7040);
nor U9399 (N_9399,N_6595,N_6929);
xor U9400 (N_9400,N_7450,N_7207);
and U9401 (N_9401,N_7833,N_7509);
or U9402 (N_9402,N_7891,N_6795);
nor U9403 (N_9403,N_6378,N_7206);
and U9404 (N_9404,N_6764,N_7940);
nor U9405 (N_9405,N_6684,N_7250);
nand U9406 (N_9406,N_6354,N_6174);
nor U9407 (N_9407,N_7420,N_7987);
nand U9408 (N_9408,N_7450,N_7862);
or U9409 (N_9409,N_6376,N_7819);
nor U9410 (N_9410,N_6511,N_7980);
nand U9411 (N_9411,N_7363,N_6585);
nand U9412 (N_9412,N_6146,N_7404);
nor U9413 (N_9413,N_7563,N_6026);
nand U9414 (N_9414,N_7507,N_7539);
and U9415 (N_9415,N_7567,N_6046);
xnor U9416 (N_9416,N_7496,N_7886);
nand U9417 (N_9417,N_7012,N_6243);
nand U9418 (N_9418,N_6615,N_6116);
and U9419 (N_9419,N_7772,N_7281);
xor U9420 (N_9420,N_7752,N_7538);
nor U9421 (N_9421,N_7711,N_6496);
nand U9422 (N_9422,N_7668,N_7078);
xnor U9423 (N_9423,N_7442,N_6631);
or U9424 (N_9424,N_7940,N_6046);
and U9425 (N_9425,N_6144,N_7385);
nor U9426 (N_9426,N_7977,N_7601);
or U9427 (N_9427,N_7635,N_6163);
nor U9428 (N_9428,N_6250,N_7375);
nor U9429 (N_9429,N_6240,N_6656);
or U9430 (N_9430,N_6253,N_7670);
nand U9431 (N_9431,N_6372,N_6661);
or U9432 (N_9432,N_7159,N_7027);
nor U9433 (N_9433,N_6810,N_6847);
nor U9434 (N_9434,N_6200,N_6015);
xor U9435 (N_9435,N_6686,N_7151);
and U9436 (N_9436,N_6128,N_6938);
nand U9437 (N_9437,N_6905,N_7059);
or U9438 (N_9438,N_7387,N_6499);
or U9439 (N_9439,N_6006,N_7560);
xor U9440 (N_9440,N_6154,N_7946);
nand U9441 (N_9441,N_7433,N_7909);
and U9442 (N_9442,N_6472,N_7650);
xnor U9443 (N_9443,N_6370,N_6265);
nor U9444 (N_9444,N_7513,N_7382);
or U9445 (N_9445,N_6934,N_6537);
and U9446 (N_9446,N_6999,N_6683);
or U9447 (N_9447,N_7984,N_6637);
nand U9448 (N_9448,N_7771,N_7194);
nand U9449 (N_9449,N_7865,N_6089);
nand U9450 (N_9450,N_7231,N_7553);
nor U9451 (N_9451,N_7118,N_6294);
or U9452 (N_9452,N_7104,N_7811);
nor U9453 (N_9453,N_6784,N_7506);
nand U9454 (N_9454,N_7918,N_7313);
or U9455 (N_9455,N_6436,N_6665);
nand U9456 (N_9456,N_7047,N_7244);
nand U9457 (N_9457,N_7479,N_7613);
nor U9458 (N_9458,N_6648,N_7776);
and U9459 (N_9459,N_6008,N_6435);
and U9460 (N_9460,N_7879,N_6081);
xnor U9461 (N_9461,N_7320,N_6346);
nand U9462 (N_9462,N_6385,N_7415);
nand U9463 (N_9463,N_7705,N_6992);
xor U9464 (N_9464,N_7147,N_7328);
nor U9465 (N_9465,N_7463,N_7422);
xnor U9466 (N_9466,N_6786,N_7277);
and U9467 (N_9467,N_7040,N_6313);
nor U9468 (N_9468,N_7973,N_6864);
nand U9469 (N_9469,N_7509,N_7424);
nand U9470 (N_9470,N_6793,N_7954);
nor U9471 (N_9471,N_7123,N_6036);
xnor U9472 (N_9472,N_6480,N_7365);
xor U9473 (N_9473,N_6221,N_7121);
xor U9474 (N_9474,N_7387,N_6307);
or U9475 (N_9475,N_6066,N_7923);
or U9476 (N_9476,N_6385,N_6995);
and U9477 (N_9477,N_6721,N_6758);
or U9478 (N_9478,N_6340,N_7038);
nor U9479 (N_9479,N_7915,N_6751);
and U9480 (N_9480,N_7933,N_6780);
nand U9481 (N_9481,N_7855,N_7045);
nor U9482 (N_9482,N_7152,N_6000);
and U9483 (N_9483,N_7542,N_6155);
or U9484 (N_9484,N_7470,N_7858);
nor U9485 (N_9485,N_6229,N_7332);
nand U9486 (N_9486,N_6373,N_7180);
and U9487 (N_9487,N_7464,N_6698);
nor U9488 (N_9488,N_6354,N_6359);
or U9489 (N_9489,N_6060,N_6845);
nand U9490 (N_9490,N_7818,N_7674);
nand U9491 (N_9491,N_6434,N_7127);
xnor U9492 (N_9492,N_6811,N_7036);
and U9493 (N_9493,N_6870,N_6454);
and U9494 (N_9494,N_6095,N_7761);
xor U9495 (N_9495,N_7576,N_6604);
nor U9496 (N_9496,N_7304,N_6187);
nor U9497 (N_9497,N_7999,N_6138);
nor U9498 (N_9498,N_6706,N_7622);
or U9499 (N_9499,N_7358,N_7574);
nor U9500 (N_9500,N_6953,N_6530);
nand U9501 (N_9501,N_7118,N_6438);
nor U9502 (N_9502,N_6092,N_6698);
or U9503 (N_9503,N_7094,N_7347);
nand U9504 (N_9504,N_6158,N_6299);
and U9505 (N_9505,N_7952,N_6927);
nand U9506 (N_9506,N_7637,N_7799);
nand U9507 (N_9507,N_6456,N_7614);
nand U9508 (N_9508,N_7043,N_7099);
xnor U9509 (N_9509,N_6324,N_7021);
or U9510 (N_9510,N_7581,N_7045);
nor U9511 (N_9511,N_7610,N_6768);
and U9512 (N_9512,N_7885,N_6748);
nand U9513 (N_9513,N_7473,N_6771);
nand U9514 (N_9514,N_7760,N_7133);
nor U9515 (N_9515,N_7631,N_6640);
or U9516 (N_9516,N_6132,N_7649);
or U9517 (N_9517,N_6741,N_6935);
nor U9518 (N_9518,N_6775,N_6255);
nand U9519 (N_9519,N_7305,N_6317);
or U9520 (N_9520,N_7677,N_6624);
or U9521 (N_9521,N_7409,N_7151);
or U9522 (N_9522,N_6899,N_6511);
nand U9523 (N_9523,N_7990,N_7578);
nand U9524 (N_9524,N_6389,N_7956);
or U9525 (N_9525,N_7348,N_6758);
and U9526 (N_9526,N_7386,N_6609);
xor U9527 (N_9527,N_6852,N_6822);
or U9528 (N_9528,N_7018,N_6582);
nand U9529 (N_9529,N_6975,N_7190);
nand U9530 (N_9530,N_7935,N_6176);
and U9531 (N_9531,N_6284,N_6526);
or U9532 (N_9532,N_7433,N_7629);
nor U9533 (N_9533,N_6288,N_6523);
nor U9534 (N_9534,N_6483,N_6209);
and U9535 (N_9535,N_6477,N_6499);
nand U9536 (N_9536,N_6944,N_7232);
xnor U9537 (N_9537,N_7120,N_6881);
nand U9538 (N_9538,N_7400,N_6596);
xnor U9539 (N_9539,N_7400,N_6832);
and U9540 (N_9540,N_6847,N_6912);
or U9541 (N_9541,N_7736,N_6583);
nand U9542 (N_9542,N_6751,N_6371);
and U9543 (N_9543,N_7933,N_7897);
xnor U9544 (N_9544,N_6984,N_7821);
nand U9545 (N_9545,N_7722,N_7348);
nand U9546 (N_9546,N_7281,N_6753);
nor U9547 (N_9547,N_7454,N_7448);
nand U9548 (N_9548,N_6661,N_6086);
nand U9549 (N_9549,N_6527,N_7374);
and U9550 (N_9550,N_6457,N_7426);
or U9551 (N_9551,N_7678,N_7192);
nand U9552 (N_9552,N_7024,N_6080);
nand U9553 (N_9553,N_6259,N_6156);
nor U9554 (N_9554,N_7806,N_6118);
and U9555 (N_9555,N_7469,N_6337);
nor U9556 (N_9556,N_7158,N_7950);
and U9557 (N_9557,N_7154,N_6102);
nor U9558 (N_9558,N_7376,N_7919);
nand U9559 (N_9559,N_7341,N_7514);
or U9560 (N_9560,N_6332,N_7550);
or U9561 (N_9561,N_6397,N_6933);
nor U9562 (N_9562,N_6487,N_6086);
and U9563 (N_9563,N_6231,N_7977);
or U9564 (N_9564,N_6422,N_7791);
nor U9565 (N_9565,N_6852,N_7581);
and U9566 (N_9566,N_6660,N_7195);
or U9567 (N_9567,N_7147,N_7996);
or U9568 (N_9568,N_7304,N_7945);
nand U9569 (N_9569,N_6810,N_7354);
and U9570 (N_9570,N_7254,N_7185);
or U9571 (N_9571,N_7051,N_7812);
nand U9572 (N_9572,N_6556,N_6510);
or U9573 (N_9573,N_7355,N_6016);
nor U9574 (N_9574,N_6127,N_6400);
xor U9575 (N_9575,N_7137,N_6054);
nor U9576 (N_9576,N_7005,N_7397);
nand U9577 (N_9577,N_7106,N_7405);
xnor U9578 (N_9578,N_6559,N_6538);
and U9579 (N_9579,N_7985,N_6977);
or U9580 (N_9580,N_6932,N_6414);
and U9581 (N_9581,N_6704,N_6511);
nor U9582 (N_9582,N_6169,N_6077);
and U9583 (N_9583,N_6957,N_6214);
xor U9584 (N_9584,N_7648,N_6263);
or U9585 (N_9585,N_7143,N_6051);
xor U9586 (N_9586,N_7013,N_7731);
nand U9587 (N_9587,N_6491,N_7351);
nor U9588 (N_9588,N_7419,N_6540);
xor U9589 (N_9589,N_6285,N_6353);
and U9590 (N_9590,N_6113,N_7824);
nand U9591 (N_9591,N_7378,N_6007);
or U9592 (N_9592,N_6361,N_6144);
or U9593 (N_9593,N_6538,N_7632);
and U9594 (N_9594,N_7753,N_7521);
xnor U9595 (N_9595,N_6882,N_7829);
and U9596 (N_9596,N_6799,N_7146);
xnor U9597 (N_9597,N_7416,N_7060);
xnor U9598 (N_9598,N_7164,N_6652);
nor U9599 (N_9599,N_7850,N_7704);
nor U9600 (N_9600,N_7813,N_7120);
or U9601 (N_9601,N_7984,N_6383);
nand U9602 (N_9602,N_7114,N_6275);
nand U9603 (N_9603,N_7428,N_7972);
or U9604 (N_9604,N_7270,N_6126);
and U9605 (N_9605,N_6761,N_7769);
and U9606 (N_9606,N_6855,N_6597);
or U9607 (N_9607,N_6267,N_6444);
nor U9608 (N_9608,N_7685,N_6329);
nor U9609 (N_9609,N_7817,N_6204);
nor U9610 (N_9610,N_7081,N_7188);
or U9611 (N_9611,N_6432,N_7094);
nand U9612 (N_9612,N_6191,N_7082);
nand U9613 (N_9613,N_7988,N_7195);
and U9614 (N_9614,N_7517,N_7427);
nand U9615 (N_9615,N_6201,N_6774);
or U9616 (N_9616,N_6144,N_7724);
nand U9617 (N_9617,N_7651,N_7534);
nand U9618 (N_9618,N_7691,N_7181);
xnor U9619 (N_9619,N_6843,N_7607);
and U9620 (N_9620,N_6491,N_7129);
xor U9621 (N_9621,N_6649,N_6907);
nand U9622 (N_9622,N_7000,N_6982);
nand U9623 (N_9623,N_6154,N_6208);
nand U9624 (N_9624,N_6218,N_6627);
xnor U9625 (N_9625,N_6923,N_7565);
nand U9626 (N_9626,N_6608,N_6955);
or U9627 (N_9627,N_7528,N_7838);
and U9628 (N_9628,N_6515,N_7833);
or U9629 (N_9629,N_6776,N_6979);
nand U9630 (N_9630,N_6683,N_6019);
and U9631 (N_9631,N_6679,N_7107);
and U9632 (N_9632,N_6233,N_6172);
and U9633 (N_9633,N_7829,N_6608);
and U9634 (N_9634,N_7080,N_7990);
and U9635 (N_9635,N_7335,N_7625);
and U9636 (N_9636,N_6054,N_6058);
nor U9637 (N_9637,N_7665,N_6507);
nor U9638 (N_9638,N_7439,N_6250);
nand U9639 (N_9639,N_6722,N_7122);
xor U9640 (N_9640,N_7267,N_7561);
nor U9641 (N_9641,N_7246,N_7478);
nor U9642 (N_9642,N_6162,N_6791);
and U9643 (N_9643,N_6989,N_6393);
nand U9644 (N_9644,N_6618,N_6120);
nand U9645 (N_9645,N_6251,N_6971);
nand U9646 (N_9646,N_6411,N_7621);
and U9647 (N_9647,N_6274,N_7758);
and U9648 (N_9648,N_6523,N_7458);
and U9649 (N_9649,N_6865,N_7659);
nor U9650 (N_9650,N_6702,N_6138);
nand U9651 (N_9651,N_6582,N_7314);
nand U9652 (N_9652,N_7132,N_6609);
xor U9653 (N_9653,N_7848,N_6659);
or U9654 (N_9654,N_7613,N_6492);
xor U9655 (N_9655,N_7014,N_6403);
nand U9656 (N_9656,N_6937,N_7235);
nor U9657 (N_9657,N_6205,N_6697);
and U9658 (N_9658,N_7029,N_6547);
and U9659 (N_9659,N_6369,N_6612);
nor U9660 (N_9660,N_7512,N_7446);
or U9661 (N_9661,N_7155,N_7596);
nor U9662 (N_9662,N_7076,N_7131);
xnor U9663 (N_9663,N_7247,N_6757);
nand U9664 (N_9664,N_7831,N_6065);
nand U9665 (N_9665,N_7915,N_7657);
nor U9666 (N_9666,N_6735,N_7685);
or U9667 (N_9667,N_7148,N_7659);
nor U9668 (N_9668,N_7227,N_6026);
nand U9669 (N_9669,N_6147,N_7494);
nor U9670 (N_9670,N_7199,N_7674);
nor U9671 (N_9671,N_6617,N_6997);
or U9672 (N_9672,N_7722,N_7277);
and U9673 (N_9673,N_6542,N_6342);
or U9674 (N_9674,N_6193,N_7299);
and U9675 (N_9675,N_7982,N_6635);
and U9676 (N_9676,N_7119,N_7329);
or U9677 (N_9677,N_6326,N_6145);
or U9678 (N_9678,N_7732,N_7412);
or U9679 (N_9679,N_7899,N_6701);
or U9680 (N_9680,N_7573,N_6601);
nand U9681 (N_9681,N_6042,N_6937);
xnor U9682 (N_9682,N_6391,N_6358);
and U9683 (N_9683,N_6615,N_7412);
and U9684 (N_9684,N_7589,N_7551);
nand U9685 (N_9685,N_7193,N_7455);
nor U9686 (N_9686,N_6755,N_6962);
nor U9687 (N_9687,N_7787,N_7414);
xnor U9688 (N_9688,N_6011,N_7187);
nand U9689 (N_9689,N_7229,N_7736);
xnor U9690 (N_9690,N_7791,N_6677);
xor U9691 (N_9691,N_7489,N_6125);
nand U9692 (N_9692,N_6361,N_6263);
or U9693 (N_9693,N_6348,N_7300);
and U9694 (N_9694,N_7460,N_7084);
nand U9695 (N_9695,N_6017,N_6385);
or U9696 (N_9696,N_7132,N_7082);
nand U9697 (N_9697,N_6807,N_6343);
xnor U9698 (N_9698,N_6381,N_6045);
xnor U9699 (N_9699,N_7657,N_6118);
and U9700 (N_9700,N_6868,N_6308);
or U9701 (N_9701,N_7875,N_7061);
or U9702 (N_9702,N_6303,N_7190);
nand U9703 (N_9703,N_6464,N_7096);
nand U9704 (N_9704,N_6482,N_7548);
nor U9705 (N_9705,N_6061,N_7141);
nor U9706 (N_9706,N_7052,N_7530);
nand U9707 (N_9707,N_7021,N_7587);
and U9708 (N_9708,N_7088,N_6030);
or U9709 (N_9709,N_6921,N_7902);
xnor U9710 (N_9710,N_7578,N_7379);
xnor U9711 (N_9711,N_7572,N_7743);
or U9712 (N_9712,N_7635,N_7495);
or U9713 (N_9713,N_6507,N_7847);
or U9714 (N_9714,N_7199,N_7451);
nand U9715 (N_9715,N_6475,N_6491);
xor U9716 (N_9716,N_6462,N_7536);
and U9717 (N_9717,N_6113,N_7188);
nor U9718 (N_9718,N_6990,N_6306);
or U9719 (N_9719,N_6108,N_6729);
or U9720 (N_9720,N_7057,N_6658);
nor U9721 (N_9721,N_7082,N_6474);
nand U9722 (N_9722,N_7204,N_6032);
nor U9723 (N_9723,N_6574,N_7022);
nand U9724 (N_9724,N_7128,N_7355);
xor U9725 (N_9725,N_6236,N_6555);
and U9726 (N_9726,N_7947,N_7706);
or U9727 (N_9727,N_6824,N_7283);
and U9728 (N_9728,N_7741,N_6590);
nor U9729 (N_9729,N_6623,N_6698);
nand U9730 (N_9730,N_6976,N_7667);
nand U9731 (N_9731,N_7457,N_7504);
nor U9732 (N_9732,N_7763,N_7383);
nor U9733 (N_9733,N_7709,N_7162);
nand U9734 (N_9734,N_6204,N_6087);
nor U9735 (N_9735,N_7813,N_6106);
nand U9736 (N_9736,N_6179,N_6003);
or U9737 (N_9737,N_6069,N_7610);
and U9738 (N_9738,N_7463,N_6396);
or U9739 (N_9739,N_6775,N_7653);
nor U9740 (N_9740,N_6818,N_7937);
nand U9741 (N_9741,N_7170,N_6065);
nor U9742 (N_9742,N_6334,N_6519);
nand U9743 (N_9743,N_6250,N_6737);
or U9744 (N_9744,N_7778,N_6636);
or U9745 (N_9745,N_7172,N_6871);
nand U9746 (N_9746,N_6402,N_6252);
or U9747 (N_9747,N_7011,N_6220);
nor U9748 (N_9748,N_7797,N_6485);
nor U9749 (N_9749,N_6746,N_6440);
and U9750 (N_9750,N_6043,N_6889);
or U9751 (N_9751,N_7013,N_7281);
or U9752 (N_9752,N_7483,N_6678);
or U9753 (N_9753,N_7601,N_7433);
nor U9754 (N_9754,N_7187,N_7870);
nand U9755 (N_9755,N_7843,N_7432);
nand U9756 (N_9756,N_6879,N_7740);
nor U9757 (N_9757,N_6060,N_6113);
or U9758 (N_9758,N_6071,N_6913);
and U9759 (N_9759,N_7979,N_6668);
nor U9760 (N_9760,N_7863,N_6669);
nand U9761 (N_9761,N_7550,N_7356);
and U9762 (N_9762,N_6753,N_6504);
nor U9763 (N_9763,N_6348,N_7774);
or U9764 (N_9764,N_6777,N_7323);
and U9765 (N_9765,N_6178,N_6524);
nor U9766 (N_9766,N_7336,N_7659);
and U9767 (N_9767,N_7548,N_6062);
and U9768 (N_9768,N_7201,N_6464);
xnor U9769 (N_9769,N_7925,N_6799);
nor U9770 (N_9770,N_7570,N_7953);
nand U9771 (N_9771,N_6264,N_6070);
nand U9772 (N_9772,N_7751,N_7805);
and U9773 (N_9773,N_6960,N_6390);
nor U9774 (N_9774,N_6432,N_7654);
or U9775 (N_9775,N_6665,N_7193);
and U9776 (N_9776,N_6664,N_6154);
nand U9777 (N_9777,N_7061,N_7726);
and U9778 (N_9778,N_7172,N_7460);
or U9779 (N_9779,N_7260,N_7399);
or U9780 (N_9780,N_6838,N_6622);
and U9781 (N_9781,N_6525,N_6513);
nand U9782 (N_9782,N_7579,N_7502);
and U9783 (N_9783,N_7583,N_6454);
and U9784 (N_9784,N_6462,N_6640);
and U9785 (N_9785,N_6411,N_7110);
xnor U9786 (N_9786,N_7549,N_7383);
nand U9787 (N_9787,N_7483,N_7437);
nor U9788 (N_9788,N_7953,N_7324);
nand U9789 (N_9789,N_6515,N_7170);
and U9790 (N_9790,N_7395,N_7513);
or U9791 (N_9791,N_6886,N_7119);
or U9792 (N_9792,N_6085,N_7206);
or U9793 (N_9793,N_6828,N_7200);
or U9794 (N_9794,N_7734,N_6484);
or U9795 (N_9795,N_7157,N_6360);
nor U9796 (N_9796,N_7479,N_7335);
xnor U9797 (N_9797,N_6780,N_6912);
and U9798 (N_9798,N_7254,N_6231);
nor U9799 (N_9799,N_7577,N_7001);
or U9800 (N_9800,N_7138,N_6336);
nor U9801 (N_9801,N_6161,N_6457);
and U9802 (N_9802,N_6195,N_7241);
or U9803 (N_9803,N_7758,N_6636);
nor U9804 (N_9804,N_6330,N_7315);
nor U9805 (N_9805,N_7529,N_7687);
nand U9806 (N_9806,N_6901,N_7144);
or U9807 (N_9807,N_6443,N_6914);
nand U9808 (N_9808,N_6452,N_6561);
or U9809 (N_9809,N_6587,N_7453);
nor U9810 (N_9810,N_6013,N_6168);
nor U9811 (N_9811,N_7000,N_6658);
nand U9812 (N_9812,N_7150,N_7070);
nor U9813 (N_9813,N_7115,N_6134);
and U9814 (N_9814,N_6438,N_7853);
or U9815 (N_9815,N_6987,N_7545);
and U9816 (N_9816,N_6940,N_7831);
and U9817 (N_9817,N_7397,N_6789);
or U9818 (N_9818,N_7712,N_6208);
and U9819 (N_9819,N_6548,N_6422);
and U9820 (N_9820,N_6442,N_7063);
and U9821 (N_9821,N_7067,N_6629);
nand U9822 (N_9822,N_6344,N_7824);
and U9823 (N_9823,N_7273,N_7539);
or U9824 (N_9824,N_6232,N_7832);
nand U9825 (N_9825,N_7797,N_6176);
or U9826 (N_9826,N_7714,N_6275);
nand U9827 (N_9827,N_7519,N_7358);
and U9828 (N_9828,N_7598,N_6807);
xnor U9829 (N_9829,N_7144,N_7228);
or U9830 (N_9830,N_7887,N_7743);
nor U9831 (N_9831,N_6446,N_7783);
or U9832 (N_9832,N_7169,N_6216);
nand U9833 (N_9833,N_7307,N_6925);
nand U9834 (N_9834,N_7355,N_6221);
nand U9835 (N_9835,N_7843,N_6332);
nand U9836 (N_9836,N_6272,N_6488);
and U9837 (N_9837,N_7123,N_6843);
and U9838 (N_9838,N_7240,N_7582);
nand U9839 (N_9839,N_7598,N_6154);
or U9840 (N_9840,N_6290,N_7058);
nand U9841 (N_9841,N_6780,N_6490);
or U9842 (N_9842,N_6921,N_7595);
nand U9843 (N_9843,N_7673,N_6846);
nand U9844 (N_9844,N_7177,N_6592);
and U9845 (N_9845,N_7971,N_6292);
nand U9846 (N_9846,N_7591,N_6157);
nand U9847 (N_9847,N_6339,N_6382);
or U9848 (N_9848,N_6154,N_6760);
xor U9849 (N_9849,N_7691,N_7462);
or U9850 (N_9850,N_6207,N_7653);
and U9851 (N_9851,N_7302,N_7922);
and U9852 (N_9852,N_7968,N_7263);
nor U9853 (N_9853,N_7630,N_6571);
xnor U9854 (N_9854,N_7757,N_7945);
nand U9855 (N_9855,N_7659,N_7698);
or U9856 (N_9856,N_6950,N_7894);
nand U9857 (N_9857,N_6794,N_6176);
nand U9858 (N_9858,N_6141,N_6293);
xnor U9859 (N_9859,N_7146,N_6417);
and U9860 (N_9860,N_7123,N_6174);
nor U9861 (N_9861,N_6428,N_7066);
or U9862 (N_9862,N_6938,N_7504);
or U9863 (N_9863,N_7200,N_7136);
nor U9864 (N_9864,N_6425,N_7617);
and U9865 (N_9865,N_7726,N_6542);
nor U9866 (N_9866,N_7261,N_7897);
or U9867 (N_9867,N_6589,N_6122);
and U9868 (N_9868,N_7879,N_7077);
or U9869 (N_9869,N_6464,N_7939);
and U9870 (N_9870,N_6472,N_6903);
xnor U9871 (N_9871,N_6609,N_6134);
and U9872 (N_9872,N_7249,N_6671);
nor U9873 (N_9873,N_6886,N_7773);
nor U9874 (N_9874,N_7481,N_7694);
and U9875 (N_9875,N_6294,N_7944);
or U9876 (N_9876,N_7467,N_7548);
or U9877 (N_9877,N_7957,N_7758);
or U9878 (N_9878,N_7937,N_7727);
nor U9879 (N_9879,N_6850,N_7794);
or U9880 (N_9880,N_6855,N_6192);
and U9881 (N_9881,N_6112,N_7656);
nor U9882 (N_9882,N_6521,N_7984);
or U9883 (N_9883,N_6214,N_6832);
or U9884 (N_9884,N_6444,N_7271);
and U9885 (N_9885,N_7349,N_7631);
or U9886 (N_9886,N_6681,N_6764);
or U9887 (N_9887,N_6880,N_7458);
and U9888 (N_9888,N_6404,N_7730);
or U9889 (N_9889,N_7124,N_7724);
or U9890 (N_9890,N_7909,N_7664);
and U9891 (N_9891,N_6235,N_6885);
nand U9892 (N_9892,N_7099,N_7893);
and U9893 (N_9893,N_6597,N_6314);
or U9894 (N_9894,N_6952,N_7142);
and U9895 (N_9895,N_7622,N_6994);
and U9896 (N_9896,N_6726,N_6961);
nand U9897 (N_9897,N_6787,N_6847);
or U9898 (N_9898,N_6304,N_6505);
xor U9899 (N_9899,N_6353,N_7859);
and U9900 (N_9900,N_6937,N_7694);
nor U9901 (N_9901,N_6938,N_7513);
xor U9902 (N_9902,N_6214,N_6312);
or U9903 (N_9903,N_7810,N_6614);
or U9904 (N_9904,N_6835,N_7697);
xor U9905 (N_9905,N_7247,N_6783);
nand U9906 (N_9906,N_6293,N_7949);
nor U9907 (N_9907,N_6429,N_6461);
and U9908 (N_9908,N_7569,N_6834);
nand U9909 (N_9909,N_7783,N_7347);
and U9910 (N_9910,N_7489,N_7057);
or U9911 (N_9911,N_7415,N_7380);
and U9912 (N_9912,N_6572,N_6421);
or U9913 (N_9913,N_7948,N_7599);
nor U9914 (N_9914,N_6928,N_7309);
or U9915 (N_9915,N_7394,N_7227);
nor U9916 (N_9916,N_7158,N_6721);
or U9917 (N_9917,N_7511,N_6492);
xnor U9918 (N_9918,N_7976,N_6841);
and U9919 (N_9919,N_6433,N_6365);
and U9920 (N_9920,N_6051,N_7268);
or U9921 (N_9921,N_6876,N_7701);
and U9922 (N_9922,N_6554,N_7511);
xnor U9923 (N_9923,N_6978,N_7169);
xor U9924 (N_9924,N_7321,N_7796);
xnor U9925 (N_9925,N_7709,N_7250);
and U9926 (N_9926,N_7858,N_6028);
or U9927 (N_9927,N_7070,N_6710);
or U9928 (N_9928,N_7901,N_7947);
or U9929 (N_9929,N_7385,N_7921);
and U9930 (N_9930,N_6502,N_6031);
nor U9931 (N_9931,N_6787,N_6100);
and U9932 (N_9932,N_7776,N_6996);
nand U9933 (N_9933,N_6713,N_7020);
or U9934 (N_9934,N_6217,N_7982);
and U9935 (N_9935,N_7205,N_7948);
or U9936 (N_9936,N_7740,N_6487);
and U9937 (N_9937,N_7314,N_6266);
and U9938 (N_9938,N_7905,N_6444);
nand U9939 (N_9939,N_6801,N_7433);
nor U9940 (N_9940,N_7833,N_7745);
nor U9941 (N_9941,N_6020,N_7833);
nand U9942 (N_9942,N_7207,N_6903);
nand U9943 (N_9943,N_7247,N_7881);
nor U9944 (N_9944,N_6885,N_6518);
nand U9945 (N_9945,N_7214,N_6748);
nand U9946 (N_9946,N_7536,N_7030);
nand U9947 (N_9947,N_7302,N_7887);
xnor U9948 (N_9948,N_7106,N_7988);
nand U9949 (N_9949,N_6974,N_6586);
or U9950 (N_9950,N_6025,N_7401);
and U9951 (N_9951,N_6661,N_6472);
nor U9952 (N_9952,N_7071,N_6983);
nor U9953 (N_9953,N_6311,N_7952);
or U9954 (N_9954,N_6554,N_7832);
nor U9955 (N_9955,N_6861,N_6123);
or U9956 (N_9956,N_6893,N_6574);
or U9957 (N_9957,N_6842,N_7935);
nor U9958 (N_9958,N_7429,N_7856);
nor U9959 (N_9959,N_7347,N_7961);
or U9960 (N_9960,N_7281,N_7778);
nand U9961 (N_9961,N_6310,N_7763);
nor U9962 (N_9962,N_6683,N_7881);
xnor U9963 (N_9963,N_7227,N_7160);
nor U9964 (N_9964,N_7774,N_7921);
and U9965 (N_9965,N_7348,N_6414);
nor U9966 (N_9966,N_6912,N_6781);
and U9967 (N_9967,N_6190,N_7824);
nand U9968 (N_9968,N_6430,N_7962);
and U9969 (N_9969,N_7175,N_7456);
or U9970 (N_9970,N_7485,N_6483);
nor U9971 (N_9971,N_6179,N_6600);
or U9972 (N_9972,N_7432,N_6200);
xnor U9973 (N_9973,N_7799,N_7896);
nor U9974 (N_9974,N_6458,N_7104);
and U9975 (N_9975,N_7975,N_7844);
xnor U9976 (N_9976,N_7975,N_7458);
or U9977 (N_9977,N_7651,N_6368);
and U9978 (N_9978,N_7040,N_7660);
and U9979 (N_9979,N_6913,N_6539);
nand U9980 (N_9980,N_6889,N_7038);
nand U9981 (N_9981,N_7172,N_6943);
and U9982 (N_9982,N_6278,N_6042);
nor U9983 (N_9983,N_6780,N_6491);
and U9984 (N_9984,N_7294,N_6790);
and U9985 (N_9985,N_7087,N_6452);
or U9986 (N_9986,N_7242,N_7566);
nand U9987 (N_9987,N_7100,N_6750);
or U9988 (N_9988,N_6452,N_7948);
or U9989 (N_9989,N_7899,N_6188);
and U9990 (N_9990,N_6598,N_6499);
and U9991 (N_9991,N_6918,N_6838);
or U9992 (N_9992,N_7349,N_6597);
and U9993 (N_9993,N_6650,N_6997);
nor U9994 (N_9994,N_6047,N_7716);
nand U9995 (N_9995,N_7016,N_7210);
and U9996 (N_9996,N_7380,N_6605);
nor U9997 (N_9997,N_6319,N_7158);
nor U9998 (N_9998,N_7498,N_7061);
or U9999 (N_9999,N_7580,N_7834);
or U10000 (N_10000,N_8182,N_9172);
and U10001 (N_10001,N_8797,N_8954);
nand U10002 (N_10002,N_8903,N_8846);
nor U10003 (N_10003,N_9686,N_9466);
xor U10004 (N_10004,N_9939,N_9186);
or U10005 (N_10005,N_8329,N_9909);
or U10006 (N_10006,N_9456,N_8408);
and U10007 (N_10007,N_8990,N_9424);
and U10008 (N_10008,N_9638,N_8998);
xor U10009 (N_10009,N_9825,N_9930);
or U10010 (N_10010,N_8298,N_8442);
or U10011 (N_10011,N_8682,N_9067);
xor U10012 (N_10012,N_9816,N_8301);
nor U10013 (N_10013,N_9232,N_9159);
and U10014 (N_10014,N_8997,N_9734);
nand U10015 (N_10015,N_8170,N_8135);
and U10016 (N_10016,N_9913,N_9807);
nor U10017 (N_10017,N_8089,N_9286);
or U10018 (N_10018,N_8392,N_8029);
nor U10019 (N_10019,N_9020,N_9918);
nor U10020 (N_10020,N_9979,N_8163);
nand U10021 (N_10021,N_9268,N_9205);
nand U10022 (N_10022,N_8852,N_8529);
xnor U10023 (N_10023,N_9303,N_8400);
or U10024 (N_10024,N_9900,N_9077);
and U10025 (N_10025,N_9097,N_8021);
nor U10026 (N_10026,N_8932,N_9530);
xor U10027 (N_10027,N_8896,N_9472);
and U10028 (N_10028,N_8981,N_8890);
or U10029 (N_10029,N_8321,N_9084);
and U10030 (N_10030,N_8055,N_8638);
and U10031 (N_10031,N_8702,N_9748);
nor U10032 (N_10032,N_9753,N_8547);
nand U10033 (N_10033,N_8088,N_9532);
nor U10034 (N_10034,N_8022,N_9922);
nand U10035 (N_10035,N_8763,N_8709);
and U10036 (N_10036,N_9203,N_9740);
or U10037 (N_10037,N_8935,N_8827);
nand U10038 (N_10038,N_9414,N_9502);
nand U10039 (N_10039,N_8794,N_8753);
xor U10040 (N_10040,N_9174,N_8479);
nor U10041 (N_10041,N_9980,N_8663);
nor U10042 (N_10042,N_8995,N_9643);
or U10043 (N_10043,N_9299,N_9945);
nand U10044 (N_10044,N_8750,N_8677);
nand U10045 (N_10045,N_9648,N_9024);
or U10046 (N_10046,N_8785,N_8410);
xnor U10047 (N_10047,N_9861,N_8936);
or U10048 (N_10048,N_9711,N_8715);
or U10049 (N_10049,N_9361,N_8601);
or U10050 (N_10050,N_8081,N_8421);
or U10051 (N_10051,N_9607,N_9765);
or U10052 (N_10052,N_9782,N_8095);
nand U10053 (N_10053,N_8978,N_8538);
nand U10054 (N_10054,N_8251,N_9082);
nand U10055 (N_10055,N_9291,N_8793);
or U10056 (N_10056,N_8107,N_9309);
nand U10057 (N_10057,N_9636,N_9368);
nand U10058 (N_10058,N_9046,N_9381);
or U10059 (N_10059,N_9070,N_9546);
nor U10060 (N_10060,N_8098,N_9273);
or U10061 (N_10061,N_9146,N_9064);
or U10062 (N_10062,N_9253,N_8411);
or U10063 (N_10063,N_9427,N_8803);
nor U10064 (N_10064,N_9104,N_9801);
or U10065 (N_10065,N_9495,N_9614);
or U10066 (N_10066,N_8657,N_9944);
or U10067 (N_10067,N_9572,N_8207);
and U10068 (N_10068,N_9738,N_8085);
and U10069 (N_10069,N_8099,N_9359);
and U10070 (N_10070,N_9221,N_9783);
and U10071 (N_10071,N_9013,N_8204);
and U10072 (N_10072,N_8431,N_8539);
nand U10073 (N_10073,N_8805,N_9177);
xnor U10074 (N_10074,N_8623,N_9010);
nand U10075 (N_10075,N_8439,N_9600);
or U10076 (N_10076,N_8059,N_8983);
and U10077 (N_10077,N_8551,N_9540);
or U10078 (N_10078,N_8327,N_9371);
nor U10079 (N_10079,N_9586,N_9398);
nor U10080 (N_10080,N_9343,N_8955);
and U10081 (N_10081,N_8028,N_9356);
or U10082 (N_10082,N_9248,N_8687);
and U10083 (N_10083,N_9580,N_9790);
or U10084 (N_10084,N_9876,N_9470);
nand U10085 (N_10085,N_8473,N_9292);
xor U10086 (N_10086,N_8842,N_8171);
xnor U10087 (N_10087,N_8974,N_8643);
nand U10088 (N_10088,N_8299,N_9829);
or U10089 (N_10089,N_9053,N_8986);
or U10090 (N_10090,N_8331,N_8549);
nor U10091 (N_10091,N_8553,N_9797);
nor U10092 (N_10092,N_8150,N_9948);
nor U10093 (N_10093,N_8712,N_8596);
nand U10094 (N_10094,N_9805,N_9851);
and U10095 (N_10095,N_9644,N_9435);
and U10096 (N_10096,N_9812,N_9353);
or U10097 (N_10097,N_8821,N_8219);
nor U10098 (N_10098,N_9731,N_9525);
or U10099 (N_10099,N_9276,N_9283);
or U10100 (N_10100,N_8044,N_8660);
nor U10101 (N_10101,N_9231,N_9187);
nand U10102 (N_10102,N_8911,N_9244);
nor U10103 (N_10103,N_8308,N_9976);
nor U10104 (N_10104,N_9620,N_9327);
and U10105 (N_10105,N_8880,N_9406);
or U10106 (N_10106,N_8245,N_8965);
nor U10107 (N_10107,N_9729,N_9601);
nand U10108 (N_10108,N_9934,N_9306);
and U10109 (N_10109,N_8372,N_9415);
or U10110 (N_10110,N_8295,N_9854);
nand U10111 (N_10111,N_8428,N_9955);
and U10112 (N_10112,N_9950,N_8909);
or U10113 (N_10113,N_9687,N_9412);
nand U10114 (N_10114,N_9637,N_9723);
nor U10115 (N_10115,N_9668,N_9933);
nand U10116 (N_10116,N_8336,N_8783);
nor U10117 (N_10117,N_8406,N_8719);
nor U10118 (N_10118,N_8187,N_8949);
and U10119 (N_10119,N_8233,N_9565);
nor U10120 (N_10120,N_9655,N_8654);
nor U10121 (N_10121,N_9049,N_8923);
nor U10122 (N_10122,N_8658,N_8863);
or U10123 (N_10123,N_8288,N_9337);
and U10124 (N_10124,N_8686,N_8563);
or U10125 (N_10125,N_8109,N_8378);
and U10126 (N_10126,N_8748,N_9213);
and U10127 (N_10127,N_9258,N_8090);
nor U10128 (N_10128,N_8031,N_8250);
and U10129 (N_10129,N_8418,N_9217);
or U10130 (N_10130,N_8145,N_8355);
and U10131 (N_10131,N_8987,N_9094);
and U10132 (N_10132,N_8362,N_8625);
xor U10133 (N_10133,N_8840,N_9521);
and U10134 (N_10134,N_9014,N_9015);
nor U10135 (N_10135,N_8594,N_9233);
and U10136 (N_10136,N_9664,N_8968);
or U10137 (N_10137,N_9092,N_9660);
nor U10138 (N_10138,N_9150,N_9452);
nand U10139 (N_10139,N_8620,N_8943);
nor U10140 (N_10140,N_9863,N_9430);
xnor U10141 (N_10141,N_8404,N_8312);
and U10142 (N_10142,N_9761,N_8272);
or U10143 (N_10143,N_8086,N_8721);
and U10144 (N_10144,N_8957,N_9019);
nand U10145 (N_10145,N_9606,N_8169);
nand U10146 (N_10146,N_8665,N_9338);
nor U10147 (N_10147,N_8064,N_9308);
xnor U10148 (N_10148,N_9228,N_9744);
or U10149 (N_10149,N_8074,N_9163);
and U10150 (N_10150,N_8789,N_9514);
nor U10151 (N_10151,N_9847,N_9647);
and U10152 (N_10152,N_9075,N_8609);
and U10153 (N_10153,N_9208,N_9106);
or U10154 (N_10154,N_8886,N_8699);
nor U10155 (N_10155,N_9493,N_8722);
nand U10156 (N_10156,N_9635,N_9946);
and U10157 (N_10157,N_9333,N_9973);
nor U10158 (N_10158,N_8924,N_9551);
nor U10159 (N_10159,N_9195,N_8056);
and U10160 (N_10160,N_8144,N_8477);
or U10161 (N_10161,N_9113,N_8693);
xor U10162 (N_10162,N_8588,N_8158);
and U10163 (N_10163,N_9017,N_8931);
nor U10164 (N_10164,N_8466,N_9853);
nor U10165 (N_10165,N_8894,N_9780);
or U10166 (N_10166,N_9619,N_8007);
nor U10167 (N_10167,N_8166,N_9622);
and U10168 (N_10168,N_8275,N_8116);
nor U10169 (N_10169,N_8337,N_9775);
nor U10170 (N_10170,N_8037,N_8615);
and U10171 (N_10171,N_9193,N_9912);
nand U10172 (N_10172,N_9088,N_8223);
xnor U10173 (N_10173,N_9073,N_9440);
nand U10174 (N_10174,N_8613,N_9055);
and U10175 (N_10175,N_9408,N_8820);
and U10176 (N_10176,N_8427,N_9690);
nand U10177 (N_10177,N_9788,N_9531);
nor U10178 (N_10178,N_9705,N_8208);
nand U10179 (N_10179,N_9178,N_9140);
nor U10180 (N_10180,N_9870,N_9869);
and U10181 (N_10181,N_9182,N_9988);
or U10182 (N_10182,N_8456,N_9066);
and U10183 (N_10183,N_9260,N_9237);
and U10184 (N_10184,N_9842,N_9448);
and U10185 (N_10185,N_9348,N_9943);
and U10186 (N_10186,N_8485,N_9667);
xnor U10187 (N_10187,N_9995,N_8206);
nand U10188 (N_10188,N_9840,N_9692);
nor U10189 (N_10189,N_8776,N_9862);
and U10190 (N_10190,N_8213,N_9428);
and U10191 (N_10191,N_8703,N_9839);
nand U10192 (N_10192,N_8707,N_8122);
nor U10193 (N_10193,N_9553,N_8384);
and U10194 (N_10194,N_9868,N_9384);
nor U10195 (N_10195,N_8281,N_8590);
or U10196 (N_10196,N_8478,N_9305);
or U10197 (N_10197,N_9194,N_9036);
and U10198 (N_10198,N_9784,N_8258);
nand U10199 (N_10199,N_8919,N_8459);
nand U10200 (N_10200,N_8772,N_9087);
nor U10201 (N_10201,N_8354,N_9158);
and U10202 (N_10202,N_9416,N_9204);
nand U10203 (N_10203,N_8097,N_9672);
or U10204 (N_10204,N_8867,N_9541);
and U10205 (N_10205,N_9144,N_8118);
nor U10206 (N_10206,N_9575,N_9557);
nand U10207 (N_10207,N_8440,N_8697);
nor U10208 (N_10208,N_9977,N_9091);
nand U10209 (N_10209,N_8576,N_8670);
nand U10210 (N_10210,N_9986,N_9624);
or U10211 (N_10211,N_8254,N_8773);
nor U10212 (N_10212,N_9791,N_8447);
nor U10213 (N_10213,N_9068,N_9754);
nand U10214 (N_10214,N_8189,N_8950);
and U10215 (N_10215,N_8389,N_9763);
nor U10216 (N_10216,N_9069,N_8471);
or U10217 (N_10217,N_8711,N_9599);
nand U10218 (N_10218,N_9042,N_9227);
or U10219 (N_10219,N_9215,N_8181);
nand U10220 (N_10220,N_8045,N_8357);
xor U10221 (N_10221,N_8527,N_9008);
nand U10222 (N_10222,N_9402,N_9369);
nand U10223 (N_10223,N_8521,N_9028);
nor U10224 (N_10224,N_8662,N_8878);
nor U10225 (N_10225,N_8133,N_8268);
nor U10226 (N_10226,N_9375,N_8157);
nand U10227 (N_10227,N_8291,N_9363);
and U10228 (N_10228,N_9974,N_8649);
nor U10229 (N_10229,N_9706,N_8519);
nand U10230 (N_10230,N_8744,N_9379);
and U10231 (N_10231,N_9503,N_9992);
nand U10232 (N_10232,N_9282,N_8586);
and U10233 (N_10233,N_8103,N_9483);
nor U10234 (N_10234,N_9724,N_8173);
or U10235 (N_10235,N_8869,N_9374);
nand U10236 (N_10236,N_8339,N_9315);
and U10237 (N_10237,N_8335,N_9824);
and U10238 (N_10238,N_8795,N_9143);
and U10239 (N_10239,N_8946,N_8778);
nand U10240 (N_10240,N_9603,N_8104);
xnor U10241 (N_10241,N_9190,N_9076);
or U10242 (N_10242,N_8490,N_8496);
nor U10243 (N_10243,N_8835,N_9991);
or U10244 (N_10244,N_9778,N_9544);
nand U10245 (N_10245,N_8728,N_8328);
nor U10246 (N_10246,N_8141,N_9582);
or U10247 (N_10247,N_8603,N_9935);
nand U10248 (N_10248,N_9639,N_9828);
or U10249 (N_10249,N_8115,N_8832);
and U10250 (N_10250,N_8984,N_9405);
or U10251 (N_10251,N_8102,N_8239);
and U10252 (N_10252,N_8787,N_9394);
or U10253 (N_10253,N_9490,N_9718);
and U10254 (N_10254,N_8651,N_9859);
or U10255 (N_10255,N_9044,N_8433);
and U10256 (N_10256,N_9279,N_8648);
and U10257 (N_10257,N_9662,N_8422);
or U10258 (N_10258,N_8489,N_9362);
nand U10259 (N_10259,N_9684,N_8664);
nor U10260 (N_10260,N_8426,N_9832);
nand U10261 (N_10261,N_8515,N_8026);
or U10262 (N_10262,N_8856,N_8353);
nand U10263 (N_10263,N_9674,N_9968);
nand U10264 (N_10264,N_9081,N_9366);
nor U10265 (N_10265,N_9629,N_8151);
or U10266 (N_10266,N_9399,N_8540);
and U10267 (N_10267,N_8520,N_8641);
nor U10268 (N_10268,N_8083,N_9025);
xnor U10269 (N_10269,N_9243,N_8667);
or U10270 (N_10270,N_9903,N_9189);
nor U10271 (N_10271,N_9899,N_8154);
xnor U10272 (N_10272,N_8800,N_8417);
nor U10273 (N_10273,N_8153,N_9485);
and U10274 (N_10274,N_8374,N_9730);
or U10275 (N_10275,N_8070,N_8132);
nand U10276 (N_10276,N_8148,N_9888);
nor U10277 (N_10277,N_8242,N_8191);
and U10278 (N_10278,N_8380,N_8830);
or U10279 (N_10279,N_9443,N_9925);
nand U10280 (N_10280,N_9200,N_9133);
or U10281 (N_10281,N_8991,N_9093);
and U10282 (N_10282,N_9160,N_9479);
nor U10283 (N_10283,N_9026,N_9891);
or U10284 (N_10284,N_9835,N_8444);
and U10285 (N_10285,N_8348,N_8416);
nand U10286 (N_10286,N_8967,N_9486);
nor U10287 (N_10287,N_8390,N_9115);
nand U10288 (N_10288,N_8514,N_9849);
nor U10289 (N_10289,N_9071,N_8105);
nor U10290 (N_10290,N_8409,N_8303);
xor U10291 (N_10291,N_9746,N_8460);
or U10292 (N_10292,N_8541,N_9852);
and U10293 (N_10293,N_8033,N_8745);
or U10294 (N_10294,N_9978,N_9242);
xor U10295 (N_10295,N_9167,N_8685);
nor U10296 (N_10296,N_8391,N_9915);
nor U10297 (N_10297,N_9882,N_8696);
nand U10298 (N_10298,N_9206,N_9155);
nand U10299 (N_10299,N_9442,N_9289);
and U10300 (N_10300,N_8084,N_8761);
nand U10301 (N_10301,N_9739,N_9389);
nand U10302 (N_10302,N_9665,N_9858);
xnor U10303 (N_10303,N_9449,N_9278);
nor U10304 (N_10304,N_8196,N_9340);
nor U10305 (N_10305,N_8113,N_8435);
nand U10306 (N_10306,N_8854,N_9994);
nor U10307 (N_10307,N_9128,N_9728);
nor U10308 (N_10308,N_8899,N_9760);
nand U10309 (N_10309,N_9577,N_9130);
or U10310 (N_10310,N_9651,N_9578);
and U10311 (N_10311,N_9675,N_9523);
nand U10312 (N_10312,N_8111,N_9387);
xor U10313 (N_10313,N_9464,N_8221);
or U10314 (N_10314,N_9170,N_9681);
xnor U10315 (N_10315,N_9112,N_8143);
and U10316 (N_10316,N_8286,N_8972);
nor U10317 (N_10317,N_9583,N_8680);
or U10318 (N_10318,N_8513,N_8566);
nand U10319 (N_10319,N_8383,N_8762);
nand U10320 (N_10320,N_8629,N_8733);
and U10321 (N_10321,N_9608,N_8398);
nor U10322 (N_10322,N_8718,N_9513);
nor U10323 (N_10323,N_8264,N_8175);
nand U10324 (N_10324,N_9520,N_9218);
nor U10325 (N_10325,N_9391,N_8066);
or U10326 (N_10326,N_8689,N_9390);
or U10327 (N_10327,N_8244,N_8347);
and U10328 (N_10328,N_9589,N_8970);
nand U10329 (N_10329,N_8727,N_9111);
nor U10330 (N_10330,N_8945,N_9236);
and U10331 (N_10331,N_8973,N_8907);
nand U10332 (N_10332,N_9080,N_9039);
xor U10333 (N_10333,N_9936,N_8533);
and U10334 (N_10334,N_8005,N_8860);
nor U10335 (N_10335,N_8545,N_9222);
nor U10336 (N_10336,N_8237,N_9972);
nor U10337 (N_10337,N_8634,N_8216);
nand U10338 (N_10338,N_8558,N_9984);
or U10339 (N_10339,N_9197,N_8598);
or U10340 (N_10340,N_9998,N_9779);
nor U10341 (N_10341,N_9697,N_9357);
xor U10342 (N_10342,N_8669,N_9074);
nand U10343 (N_10343,N_8332,N_8290);
or U10344 (N_10344,N_9207,N_9680);
nor U10345 (N_10345,N_9814,N_9180);
nor U10346 (N_10346,N_9538,N_9453);
nand U10347 (N_10347,N_8307,N_9226);
nor U10348 (N_10348,N_8504,N_8914);
or U10349 (N_10349,N_9669,N_8072);
nor U10350 (N_10350,N_8094,N_8544);
or U10351 (N_10351,N_8593,N_9507);
or U10352 (N_10352,N_9400,N_9060);
nand U10353 (N_10353,N_8063,N_9191);
nor U10354 (N_10354,N_9096,N_8351);
and U10355 (N_10355,N_8069,N_9319);
and U10356 (N_10356,N_9336,N_8925);
nor U10357 (N_10357,N_8626,N_9331);
nand U10358 (N_10358,N_8215,N_9127);
xnor U10359 (N_10359,N_9896,N_9764);
nor U10360 (N_10360,N_8430,N_8947);
xor U10361 (N_10361,N_8396,N_9623);
nor U10362 (N_10362,N_8225,N_9506);
nand U10363 (N_10363,N_8386,N_9002);
and U10364 (N_10364,N_9012,N_8554);
and U10365 (N_10365,N_8349,N_8371);
nor U10366 (N_10366,N_8448,N_8786);
nor U10367 (N_10367,N_9777,N_9004);
and U10368 (N_10368,N_9615,N_9649);
xnor U10369 (N_10369,N_8823,N_9677);
nand U10370 (N_10370,N_8532,N_8735);
or U10371 (N_10371,N_8898,N_9947);
nor U10372 (N_10372,N_9659,N_9285);
nand U10373 (N_10373,N_8849,N_8159);
or U10374 (N_10374,N_8587,N_9886);
nand U10375 (N_10375,N_8388,N_9838);
nand U10376 (N_10376,N_8270,N_8882);
nand U10377 (N_10377,N_9241,N_8222);
nor U10378 (N_10378,N_8742,N_8611);
nand U10379 (N_10379,N_8263,N_9314);
or U10380 (N_10380,N_9156,N_9249);
nor U10381 (N_10381,N_8877,N_8700);
xor U10382 (N_10382,N_9528,N_8614);
and U10383 (N_10383,N_9120,N_8049);
xnor U10384 (N_10384,N_8333,N_9820);
nor U10385 (N_10385,N_9883,N_8659);
and U10386 (N_10386,N_8012,N_9566);
nor U10387 (N_10387,N_8020,N_9999);
and U10388 (N_10388,N_9604,N_9196);
and U10389 (N_10389,N_8988,N_8969);
xnor U10390 (N_10390,N_9942,N_9656);
or U10391 (N_10391,N_8937,N_8042);
nor U10392 (N_10392,N_9247,N_9893);
nor U10393 (N_10393,N_8412,N_8673);
or U10394 (N_10394,N_9833,N_9574);
nor U10395 (N_10395,N_9003,N_9632);
nand U10396 (N_10396,N_8872,N_8829);
or U10397 (N_10397,N_8199,N_8458);
nand U10398 (N_10398,N_9109,N_8160);
nor U10399 (N_10399,N_8437,N_9489);
nand U10400 (N_10400,N_8304,N_8688);
nor U10401 (N_10401,N_8363,N_9393);
and U10402 (N_10402,N_9785,N_9845);
or U10403 (N_10403,N_8075,N_8246);
nand U10404 (N_10404,N_8161,N_8220);
xnor U10405 (N_10405,N_8274,N_9041);
and U10406 (N_10406,N_9420,N_8054);
and U10407 (N_10407,N_8790,N_8273);
nor U10408 (N_10408,N_8096,N_8377);
nand U10409 (N_10409,N_8804,N_8676);
or U10410 (N_10410,N_8198,N_8732);
and U10411 (N_10411,N_8452,N_9750);
and U10412 (N_10412,N_9919,N_9457);
nor U10413 (N_10413,N_8106,N_8505);
xnor U10414 (N_10414,N_8197,N_8350);
or U10415 (N_10415,N_8912,N_8725);
nand U10416 (N_10416,N_9515,N_8356);
or U10417 (N_10417,N_8176,N_8100);
nor U10418 (N_10418,N_8482,N_8313);
nand U10419 (N_10419,N_9179,N_9202);
nor U10420 (N_10420,N_8399,N_9749);
nand U10421 (N_10421,N_9100,N_9445);
or U10422 (N_10422,N_9524,N_8807);
or U10423 (N_10423,N_9560,N_9238);
nor U10424 (N_10424,N_8018,N_9719);
nor U10425 (N_10425,N_8730,N_8340);
nor U10426 (N_10426,N_9272,N_8009);
nor U10427 (N_10427,N_9545,N_9373);
and U10428 (N_10428,N_9009,N_9928);
xnor U10429 (N_10429,N_8468,N_8325);
nand U10430 (N_10430,N_9808,N_8491);
or U10431 (N_10431,N_9108,N_8777);
and U10432 (N_10432,N_8210,N_8724);
and U10433 (N_10433,N_9924,N_9168);
or U10434 (N_10434,N_8833,N_8977);
xnor U10435 (N_10435,N_9223,N_8155);
nor U10436 (N_10436,N_8708,N_8124);
nand U10437 (N_10437,N_8602,N_9118);
and U10438 (N_10438,N_8261,N_9011);
and U10439 (N_10439,N_8368,N_9981);
and U10440 (N_10440,N_9229,N_8650);
xnor U10441 (N_10441,N_8238,N_9031);
nor U10442 (N_10442,N_9481,N_9762);
nor U10443 (N_10443,N_9881,N_8087);
nand U10444 (N_10444,N_9822,N_9795);
xnor U10445 (N_10445,N_9539,N_8755);
nand U10446 (N_10446,N_8559,N_8865);
and U10447 (N_10447,N_9467,N_8508);
and U10448 (N_10448,N_8480,N_8975);
xor U10449 (N_10449,N_8605,N_8597);
nor U10450 (N_10450,N_8324,N_9770);
or U10451 (N_10451,N_9561,N_9358);
nand U10452 (N_10452,N_9230,N_9700);
or U10453 (N_10453,N_8910,N_9685);
nand U10454 (N_10454,N_9841,N_9458);
nor U10455 (N_10455,N_9509,N_9512);
nand U10456 (N_10456,N_9628,N_8874);
nor U10457 (N_10457,N_9296,N_9444);
and U10458 (N_10458,N_8231,N_9147);
or U10459 (N_10459,N_9409,N_9609);
and U10460 (N_10460,N_8771,N_9431);
nand U10461 (N_10461,N_9103,N_8030);
nor U10462 (N_10462,N_8736,N_9755);
xor U10463 (N_10463,N_8780,N_9261);
nand U10464 (N_10464,N_8423,N_9846);
nor U10465 (N_10465,N_8592,N_8524);
or U10466 (N_10466,N_9275,N_8958);
or U10467 (N_10467,N_8917,N_8526);
nor U10468 (N_10468,N_9184,N_8445);
xor U10469 (N_10469,N_8938,N_9792);
or U10470 (N_10470,N_9799,N_8200);
nand U10471 (N_10471,N_9617,N_8057);
nand U10472 (N_10472,N_8203,N_9904);
and U10473 (N_10473,N_9114,N_9879);
and U10474 (N_10474,N_9821,N_8413);
nor U10475 (N_10475,N_9054,N_9969);
nand U10476 (N_10476,N_9721,N_8152);
nand U10477 (N_10477,N_9450,N_8060);
xnor U10478 (N_10478,N_9872,N_9421);
nor U10479 (N_10479,N_8516,N_9311);
xnor U10480 (N_10480,N_8738,N_9475);
nor U10481 (N_10481,N_9745,N_9953);
nor U10482 (N_10482,N_9809,N_8610);
nand U10483 (N_10483,N_9256,N_8739);
nor U10484 (N_10484,N_9352,N_8073);
or U10485 (N_10485,N_9699,N_9559);
or U10486 (N_10486,N_9908,N_8193);
xnor U10487 (N_10487,N_8309,N_9878);
and U10488 (N_10488,N_9220,N_8616);
or U10489 (N_10489,N_8067,N_8752);
xnor U10490 (N_10490,N_9712,N_8214);
nor U10491 (N_10491,N_8209,N_9201);
nor U10492 (N_10492,N_8338,N_9982);
xor U10493 (N_10493,N_8844,N_9511);
or U10494 (N_10494,N_8117,N_8741);
and U10495 (N_10495,N_9488,N_9110);
nor U10496 (N_10496,N_8916,N_9594);
nand U10497 (N_10497,N_8234,N_8259);
or U10498 (N_10498,N_9403,N_8017);
or U10499 (N_10499,N_9864,N_8265);
and U10500 (N_10500,N_9722,N_8746);
xor U10501 (N_10501,N_8692,N_8006);
or U10502 (N_10502,N_8565,N_8817);
and U10503 (N_10503,N_8655,N_8901);
nor U10504 (N_10504,N_9552,N_8282);
and U10505 (N_10505,N_8573,N_9902);
nor U10506 (N_10506,N_9429,N_8717);
and U10507 (N_10507,N_8497,N_8897);
nor U10508 (N_10508,N_9786,N_8751);
nor U10509 (N_10509,N_8985,N_8394);
and U10510 (N_10510,N_8893,N_9126);
or U10511 (N_10511,N_8656,N_9473);
nor U10512 (N_10512,N_8205,N_9326);
xnor U10513 (N_10513,N_8358,N_8498);
or U10514 (N_10514,N_9673,N_9704);
nor U10515 (N_10515,N_8360,N_9625);
or U10516 (N_10516,N_9985,N_8499);
or U10517 (N_10517,N_8600,N_9463);
nand U10518 (N_10518,N_9715,N_9122);
or U10519 (N_10519,N_8622,N_8522);
or U10520 (N_10520,N_8369,N_8334);
nor U10521 (N_10521,N_9288,N_8366);
nand U10522 (N_10522,N_9504,N_8875);
or U10523 (N_10523,N_9713,N_8393);
xor U10524 (N_10524,N_8365,N_8822);
or U10525 (N_10525,N_9519,N_8053);
nand U10526 (N_10526,N_8624,N_9342);
or U10527 (N_10527,N_9702,N_8443);
nor U10528 (N_10528,N_8474,N_9696);
nand U10529 (N_10529,N_8904,N_9107);
or U10530 (N_10530,N_9162,N_8962);
nor U10531 (N_10531,N_8632,N_9378);
xnor U10532 (N_10532,N_8379,N_8232);
or U10533 (N_10533,N_9693,N_8749);
nand U10534 (N_10534,N_8010,N_8774);
nor U10535 (N_10535,N_8517,N_8889);
xnor U10536 (N_10536,N_9302,N_8228);
nor U10537 (N_10537,N_8402,N_8112);
and U10538 (N_10538,N_9446,N_9173);
nand U10539 (N_10539,N_9252,N_8462);
nand U10540 (N_10540,N_8837,N_8420);
or U10541 (N_10541,N_9817,N_9733);
nand U10542 (N_10542,N_8041,N_8454);
and U10543 (N_10543,N_8419,N_9266);
and U10544 (N_10544,N_9796,N_9246);
or U10545 (N_10545,N_9666,N_9294);
or U10546 (N_10546,N_8582,N_9078);
nor U10547 (N_10547,N_9937,N_8511);
or U10548 (N_10548,N_8283,N_9396);
and U10549 (N_10549,N_9695,N_9587);
nand U10550 (N_10550,N_8802,N_9726);
and U10551 (N_10551,N_9332,N_9460);
xnor U10552 (N_10552,N_8472,N_8811);
and U10553 (N_10553,N_8486,N_9496);
xnor U10554 (N_10554,N_8341,N_9047);
or U10555 (N_10555,N_9921,N_9757);
nand U10556 (N_10556,N_8078,N_9166);
and U10557 (N_10557,N_9548,N_9905);
nand U10558 (N_10558,N_8212,N_8782);
and U10559 (N_10559,N_9307,N_8449);
xnor U10560 (N_10560,N_8186,N_9768);
and U10561 (N_10561,N_9304,N_8760);
or U10562 (N_10562,N_9585,N_9516);
or U10563 (N_10563,N_8885,N_9810);
xnor U10564 (N_10564,N_8976,N_8289);
nor U10565 (N_10565,N_8884,N_8825);
and U10566 (N_10566,N_9491,N_9875);
and U10567 (N_10567,N_8813,N_9018);
and U10568 (N_10568,N_9259,N_8960);
nand U10569 (N_10569,N_9301,N_9958);
or U10570 (N_10570,N_8311,N_9694);
xor U10571 (N_10571,N_8121,N_9347);
nor U10572 (N_10572,N_8604,N_9322);
nor U10573 (N_10573,N_8071,N_8343);
nand U10574 (N_10574,N_9059,N_8126);
xnor U10575 (N_10575,N_8627,N_9434);
nand U10576 (N_10576,N_9037,N_8034);
or U10577 (N_10577,N_9679,N_9929);
or U10578 (N_10578,N_9441,N_8346);
nand U10579 (N_10579,N_9683,N_9906);
nor U10580 (N_10580,N_9235,N_8562);
nand U10581 (N_10581,N_9410,N_8192);
or U10582 (N_10582,N_8509,N_8000);
nor U10583 (N_10583,N_9926,N_9265);
and U10584 (N_10584,N_8831,N_8180);
xnor U10585 (N_10585,N_9250,N_8941);
nor U10586 (N_10586,N_8229,N_9927);
or U10587 (N_10587,N_8306,N_8174);
or U10588 (N_10588,N_9335,N_9670);
and U10589 (N_10589,N_8630,N_8577);
nor U10590 (N_10590,N_9766,N_8952);
nor U10591 (N_10591,N_9183,N_9756);
nor U10592 (N_10592,N_9759,N_9576);
or U10593 (N_10593,N_9914,N_9613);
nor U10594 (N_10594,N_8564,N_8873);
or U10595 (N_10595,N_8570,N_8025);
nor U10596 (N_10596,N_9284,N_9297);
nand U10597 (N_10597,N_8202,N_8591);
nor U10598 (N_10598,N_9295,N_8194);
and U10599 (N_10599,N_8999,N_8747);
or U10600 (N_10600,N_9316,N_8754);
or U10601 (N_10601,N_8939,N_9661);
nand U10602 (N_10602,N_8149,N_8572);
xor U10603 (N_10603,N_9997,N_9892);
nor U10604 (N_10604,N_9800,N_8463);
nor U10605 (N_10605,N_8930,N_9372);
nor U10606 (N_10606,N_8201,N_9567);
or U10607 (N_10607,N_8027,N_9119);
and U10608 (N_10608,N_8706,N_9462);
and U10609 (N_10609,N_9318,N_9482);
nor U10610 (N_10610,N_8345,N_8248);
nand U10611 (N_10611,N_8858,N_9526);
nor U10612 (N_10612,N_9798,N_9264);
or U10613 (N_10613,N_8179,N_9058);
nand U10614 (N_10614,N_8940,N_9225);
or U10615 (N_10615,N_8920,N_9967);
nor U10616 (N_10616,N_8227,N_9964);
nand U10617 (N_10617,N_9451,N_8876);
and U10618 (N_10618,N_9772,N_8168);
and U10619 (N_10619,N_9618,N_9072);
xnor U10620 (N_10620,N_9439,N_8134);
or U10621 (N_10621,N_9176,N_8068);
nor U10622 (N_10622,N_9157,N_9602);
or U10623 (N_10623,N_8895,N_8461);
nand U10624 (N_10624,N_8989,N_8080);
nand U10625 (N_10625,N_9099,N_8195);
or U10626 (N_10626,N_9364,N_9465);
nor U10627 (N_10627,N_8183,N_8791);
and U10628 (N_10628,N_9423,N_9469);
or U10629 (N_10629,N_9654,N_8531);
or U10630 (N_10630,N_9471,N_9323);
xor U10631 (N_10631,N_8507,N_9267);
nand U10632 (N_10632,N_8645,N_9224);
nor U10633 (N_10633,N_9138,N_9563);
nor U10634 (N_10634,N_9823,N_9413);
nand U10635 (N_10635,N_9941,N_9543);
and U10636 (N_10636,N_8518,N_9181);
nor U10637 (N_10637,N_8450,N_9045);
or U10638 (N_10638,N_9689,N_8266);
nand U10639 (N_10639,N_8555,N_8801);
nand U10640 (N_10640,N_8704,N_9940);
nand U10641 (N_10641,N_9642,N_8296);
or U10642 (N_10642,N_9508,N_8048);
nor U10643 (N_10643,N_8501,N_9787);
xnor U10644 (N_10644,N_9626,N_9932);
nor U10645 (N_10645,N_9987,N_8775);
nor U10646 (N_10646,N_8484,N_8077);
nand U10647 (N_10647,N_9534,N_8211);
and U10648 (N_10648,N_9630,N_8188);
or U10649 (N_10649,N_9437,N_9293);
and U10650 (N_10650,N_8185,N_8902);
nor U10651 (N_10651,N_8726,N_8996);
or U10652 (N_10652,N_8277,N_9123);
nor U10653 (N_10653,N_8888,N_9963);
and U10654 (N_10654,N_9344,N_9831);
nand U10655 (N_10655,N_8796,N_9171);
nand U10656 (N_10656,N_8698,N_8293);
nor U10657 (N_10657,N_9380,N_8280);
and U10658 (N_10658,N_8589,N_8317);
or U10659 (N_10659,N_9461,N_8535);
or U10660 (N_10660,N_9145,N_8612);
nor U10661 (N_10661,N_8578,N_8167);
nand U10662 (N_10662,N_8959,N_8879);
and U10663 (N_10663,N_8451,N_8848);
nand U10664 (N_10664,N_8644,N_8140);
and U10665 (N_10665,N_8502,N_9844);
nand U10666 (N_10666,N_9793,N_8734);
nor U10667 (N_10667,N_8361,N_8137);
xnor U10668 (N_10668,N_8424,N_9569);
nor U10669 (N_10669,N_8184,N_9474);
nor U10670 (N_10670,N_9533,N_9383);
nor U10671 (N_10671,N_8672,N_9907);
or U10672 (N_10672,N_8495,N_9751);
nand U10673 (N_10673,N_9737,N_9634);
nor U10674 (N_10674,N_9447,N_8666);
xnor U10675 (N_10675,N_8723,N_8494);
and U10676 (N_10676,N_8128,N_9501);
and U10677 (N_10677,N_9860,N_9627);
and U10678 (N_10678,N_9573,N_9382);
nor U10679 (N_10679,N_8381,N_9678);
nor U10680 (N_10680,N_8536,N_8757);
and U10681 (N_10681,N_8839,N_8798);
nor U10682 (N_10682,N_9641,N_8364);
xor U10683 (N_10683,N_8561,N_8767);
nand U10684 (N_10684,N_8305,N_9240);
nand U10685 (N_10685,N_8963,N_9653);
nand U10686 (N_10686,N_8883,N_8713);
and U10687 (N_10687,N_9494,N_9487);
nor U10688 (N_10688,N_9499,N_9717);
or U10689 (N_10689,N_9529,N_9300);
nor U10690 (N_10690,N_9165,N_9007);
and U10691 (N_10691,N_8262,N_9510);
nand U10692 (N_10692,N_8695,N_8701);
and U10693 (N_10693,N_8836,N_9781);
nor U10694 (N_10694,N_8768,N_8429);
and U10695 (N_10695,N_9280,N_9454);
or U10696 (N_10696,N_9149,N_8226);
xor U10697 (N_10697,N_8806,N_8934);
nand U10698 (N_10698,N_9736,N_9735);
or U10699 (N_10699,N_8892,N_8323);
nor U10700 (N_10700,N_8847,N_9522);
nor U10701 (N_10701,N_9804,N_9057);
nand U10702 (N_10702,N_8870,N_9098);
nor U10703 (N_10703,N_9478,N_8344);
and U10704 (N_10704,N_8314,N_9836);
nor U10705 (N_10705,N_9554,N_9547);
and U10706 (N_10706,N_8756,N_8230);
nand U10707 (N_10707,N_8640,N_9610);
nor U10708 (N_10708,N_9774,N_9043);
and U10709 (N_10709,N_8476,N_9830);
nor U10710 (N_10710,N_8500,N_8003);
xor U10711 (N_10711,N_8457,N_9897);
or U10712 (N_10712,N_8120,N_9579);
nand U10713 (N_10713,N_8926,N_9034);
and U10714 (N_10714,N_9274,N_9281);
nand U10715 (N_10715,N_8980,N_8928);
xor U10716 (N_10716,N_8058,N_9219);
and U10717 (N_10717,N_9758,N_9954);
nand U10718 (N_10718,N_9920,N_8011);
nand U10719 (N_10719,N_8146,N_8933);
or U10720 (N_10720,N_8862,N_9773);
nor U10721 (N_10721,N_8190,N_8887);
or U10722 (N_10722,N_8868,N_9148);
and U10723 (N_10723,N_8267,N_9650);
and U10724 (N_10724,N_9083,N_9355);
nand U10725 (N_10725,N_8130,N_8764);
nor U10726 (N_10726,N_9588,N_9251);
nor U10727 (N_10727,N_9971,N_9211);
and U10728 (N_10728,N_8956,N_9199);
nand U10729 (N_10729,N_9124,N_9826);
nand U10730 (N_10730,N_8310,N_8560);
nand U10731 (N_10731,N_8271,N_9269);
nor U10732 (N_10732,N_9827,N_9334);
and U10733 (N_10733,N_8172,N_8326);
or U10734 (N_10734,N_8617,N_8674);
and U10735 (N_10735,N_8779,N_8784);
nor U10736 (N_10736,N_8278,N_8859);
or U10737 (N_10737,N_8818,N_9255);
and U10738 (N_10738,N_8082,N_8915);
or U10739 (N_10739,N_8729,N_9271);
or U10740 (N_10740,N_9117,N_9698);
and U10741 (N_10741,N_8382,N_8671);
nand U10742 (N_10742,N_8043,N_9153);
nand U10743 (N_10743,N_9542,N_8781);
and U10744 (N_10744,N_8062,N_8855);
or U10745 (N_10745,N_9709,N_9033);
nor U10746 (N_10746,N_9965,N_9850);
nand U10747 (N_10747,N_8464,N_9433);
and U10748 (N_10748,N_9404,N_8694);
and U10749 (N_10749,N_8285,N_9917);
nor U10750 (N_10750,N_8008,N_8114);
or U10751 (N_10751,N_9767,N_8255);
and U10752 (N_10752,N_8136,N_8425);
nand U10753 (N_10753,N_9418,N_8528);
nor U10754 (N_10754,N_9714,N_8013);
and U10755 (N_10755,N_9422,N_9931);
nand U10756 (N_10756,N_8581,N_8236);
and U10757 (N_10757,N_9298,N_9263);
xnor U10758 (N_10758,N_8683,N_8032);
nand U10759 (N_10759,N_9027,N_8759);
nor U10760 (N_10760,N_8469,N_9131);
nand U10761 (N_10761,N_8982,N_9345);
nand U10762 (N_10762,N_8812,N_8036);
or U10763 (N_10763,N_9564,N_8864);
or U10764 (N_10764,N_9254,N_9970);
xnor U10765 (N_10765,N_9132,N_9819);
and U10766 (N_10766,N_9951,N_8397);
and U10767 (N_10767,N_9125,N_8001);
nor U10768 (N_10768,N_9234,N_9803);
and U10769 (N_10769,N_8110,N_8853);
and U10770 (N_10770,N_9593,N_9164);
nor U10771 (N_10771,N_8580,N_8716);
nand U10772 (N_10772,N_8953,N_8493);
xor U10773 (N_10773,N_9386,N_9455);
and U10774 (N_10774,N_9349,N_8373);
and U10775 (N_10775,N_9392,N_9874);
or U10776 (N_10776,N_8300,N_8621);
nor U10777 (N_10777,N_8523,N_8619);
and U10778 (N_10778,N_8550,N_8217);
or U10779 (N_10779,N_8537,N_8287);
or U10780 (N_10780,N_8342,N_9346);
nor U10781 (N_10781,N_9732,N_8574);
and U10782 (N_10782,N_8359,N_9535);
or U10783 (N_10783,N_9152,N_8569);
nor U10784 (N_10784,N_8123,N_9239);
xor U10785 (N_10785,N_8971,N_9596);
xnor U10786 (N_10786,N_8297,N_9657);
nor U10787 (N_10787,N_8138,N_9834);
nand U10788 (N_10788,N_8690,N_9848);
nor U10789 (N_10789,N_9742,N_9425);
xnor U10790 (N_10790,N_8828,N_8636);
or U10791 (N_10791,N_9727,N_9116);
nand U10792 (N_10792,N_8260,N_9707);
nor U10793 (N_10793,N_8395,N_9571);
nor U10794 (N_10794,N_8076,N_8178);
nand U10795 (N_10795,N_8092,N_8376);
nor U10796 (N_10796,N_9837,N_9631);
and U10797 (N_10797,N_9350,N_9584);
or U10798 (N_10798,N_8256,N_8900);
or U10799 (N_10799,N_8618,N_9426);
xor U10800 (N_10800,N_8441,N_9161);
and U10801 (N_10801,N_9376,N_9771);
or U10802 (N_10802,N_8014,N_8465);
nor U10803 (N_10803,N_8816,N_8415);
nor U10804 (N_10804,N_9050,N_8024);
and U10805 (N_10805,N_9815,N_9873);
nand U10806 (N_10806,N_8320,N_9048);
and U10807 (N_10807,N_9354,N_8047);
nand U10808 (N_10808,N_9813,N_8668);
nand U10809 (N_10809,N_9102,N_8678);
and U10810 (N_10810,N_8269,N_8675);
and U10811 (N_10811,N_8681,N_8948);
xnor U10812 (N_10812,N_8714,N_9001);
or U10813 (N_10813,N_8814,N_8039);
or U10814 (N_10814,N_8162,N_9313);
nor U10815 (N_10815,N_8483,N_8557);
nand U10816 (N_10816,N_9789,N_8119);
nor U10817 (N_10817,N_8607,N_9101);
and U10818 (N_10818,N_8131,N_8921);
nand U10819 (N_10819,N_9056,N_8841);
nor U10820 (N_10820,N_8548,N_9794);
xor U10821 (N_10821,N_9136,N_9989);
nand U10822 (N_10822,N_9811,N_8405);
and U10823 (N_10823,N_8731,N_8608);
and U10824 (N_10824,N_9029,N_9135);
nand U10825 (N_10825,N_8276,N_8407);
nor U10826 (N_10826,N_8628,N_9000);
nor U10827 (N_10827,N_9960,N_9419);
or U10828 (N_10828,N_9497,N_9975);
and U10829 (N_10829,N_9432,N_9351);
nand U10830 (N_10830,N_8646,N_9095);
or U10831 (N_10831,N_8652,N_8571);
nor U10832 (N_10832,N_8108,N_8467);
nor U10833 (N_10833,N_9377,N_9818);
nand U10834 (N_10834,N_8575,N_9198);
nor U10835 (N_10835,N_9663,N_8165);
nand U10836 (N_10836,N_8235,N_9949);
nor U10837 (N_10837,N_8401,N_8679);
xnor U10838 (N_10838,N_9006,N_8845);
or U10839 (N_10839,N_9562,N_9210);
and U10840 (N_10840,N_8595,N_8319);
nor U10841 (N_10841,N_8653,N_9016);
nand U10842 (N_10842,N_8446,N_9129);
xnor U10843 (N_10843,N_8101,N_9324);
or U10844 (N_10844,N_8302,N_9498);
and U10845 (N_10845,N_9671,N_9857);
xnor U10846 (N_10846,N_8147,N_9438);
and U10847 (N_10847,N_8913,N_8815);
and U10848 (N_10848,N_8534,N_9505);
nor U10849 (N_10849,N_9966,N_8927);
nand U10850 (N_10850,N_8918,N_9216);
nand U10851 (N_10851,N_9407,N_9468);
xor U10852 (N_10852,N_8253,N_9032);
or U10853 (N_10853,N_8164,N_8556);
nor U10854 (N_10854,N_9752,N_8488);
xnor U10855 (N_10855,N_8455,N_9492);
xnor U10856 (N_10856,N_8294,N_9401);
xor U10857 (N_10857,N_8546,N_9262);
xnor U10858 (N_10858,N_9085,N_9865);
nor U10859 (N_10859,N_8512,N_8315);
and U10860 (N_10860,N_8470,N_8808);
nor U10861 (N_10861,N_9367,N_9898);
and U10862 (N_10862,N_9983,N_8881);
nor U10863 (N_10863,N_9633,N_9121);
and U10864 (N_10864,N_9703,N_8929);
or U10865 (N_10865,N_8740,N_9151);
and U10866 (N_10866,N_9590,N_9741);
nor U10867 (N_10867,N_9592,N_9021);
and U10868 (N_10868,N_9209,N_9646);
xor U10869 (N_10869,N_9856,N_9035);
nand U10870 (N_10870,N_8002,N_8375);
or U10871 (N_10871,N_8810,N_8637);
nor U10872 (N_10872,N_8633,N_8257);
and U10873 (N_10873,N_8438,N_8871);
nand U10874 (N_10874,N_8705,N_9598);
nand U10875 (N_10875,N_8951,N_8322);
xor U10876 (N_10876,N_8770,N_8050);
and U10877 (N_10877,N_9154,N_9993);
xor U10878 (N_10878,N_8543,N_9038);
nand U10879 (N_10879,N_9611,N_8436);
nor U10880 (N_10880,N_8857,N_8584);
nor U10881 (N_10881,N_8606,N_8583);
or U10882 (N_10882,N_8769,N_9329);
nor U10883 (N_10883,N_9105,N_8922);
or U10884 (N_10884,N_9537,N_9890);
nand U10885 (N_10885,N_9959,N_8905);
and U10886 (N_10886,N_9640,N_9597);
nor U10887 (N_10887,N_8506,N_8525);
nand U10888 (N_10888,N_9802,N_8792);
nand U10889 (N_10889,N_9086,N_9555);
nand U10890 (N_10890,N_8819,N_9581);
nand U10891 (N_10891,N_8125,N_8906);
and U10892 (N_10892,N_9691,N_9330);
nor U10893 (N_10893,N_8579,N_9616);
or U10894 (N_10894,N_8966,N_9459);
xnor U10895 (N_10895,N_9395,N_8758);
or U10896 (N_10896,N_9388,N_9962);
or U10897 (N_10897,N_8639,N_8481);
nand U10898 (N_10898,N_8961,N_9568);
xor U10899 (N_10899,N_8035,N_9961);
or U10900 (N_10900,N_8492,N_9645);
or U10901 (N_10901,N_9370,N_9867);
nor U10902 (N_10902,N_9517,N_9957);
nand U10903 (N_10903,N_9134,N_8318);
or U10904 (N_10904,N_8599,N_8635);
and U10905 (N_10905,N_8079,N_8994);
xor U10906 (N_10906,N_8838,N_8434);
nor U10907 (N_10907,N_8799,N_9720);
nor U10908 (N_10908,N_9901,N_8908);
and U10909 (N_10909,N_9137,N_9889);
nand U10910 (N_10910,N_8891,N_9317);
and U10911 (N_10911,N_9621,N_9290);
nor U10912 (N_10912,N_9895,N_9871);
nor U10913 (N_10913,N_9527,N_9040);
or U10914 (N_10914,N_9339,N_8487);
xnor U10915 (N_10915,N_8023,N_8684);
nand U10916 (N_10916,N_9365,N_9325);
nor U10917 (N_10917,N_9312,N_9476);
and U10918 (N_10918,N_9417,N_8851);
or U10919 (N_10919,N_9411,N_8475);
nand U10920 (N_10920,N_8850,N_8052);
and U10921 (N_10921,N_8065,N_9436);
nand U10922 (N_10922,N_9676,N_9843);
or U10923 (N_10923,N_9556,N_9022);
nand U10924 (N_10924,N_8292,N_9052);
nand U10925 (N_10925,N_9484,N_9477);
nor U10926 (N_10926,N_9570,N_9558);
nor U10927 (N_10927,N_9956,N_9938);
nor U10928 (N_10928,N_9360,N_9652);
or U10929 (N_10929,N_9688,N_8743);
nand U10930 (N_10930,N_9923,N_9910);
or U10931 (N_10931,N_9030,N_8552);
nand U10932 (N_10932,N_9855,N_8432);
or U10933 (N_10933,N_9062,N_8061);
xor U10934 (N_10934,N_9536,N_8284);
or U10935 (N_10935,N_8944,N_9701);
nand U10936 (N_10936,N_8093,N_9328);
nand U10937 (N_10937,N_9257,N_8710);
and U10938 (N_10938,N_9090,N_8352);
and U10939 (N_10939,N_9591,N_8247);
nand U10940 (N_10940,N_8385,N_9175);
xor U10941 (N_10941,N_8177,N_9023);
nor U10942 (N_10942,N_9776,N_8585);
nor U10943 (N_10943,N_8243,N_8737);
nor U10944 (N_10944,N_9320,N_8766);
or U10945 (N_10945,N_8142,N_8503);
or U10946 (N_10946,N_9310,N_8661);
or U10947 (N_10947,N_8403,N_8240);
nor U10948 (N_10948,N_9916,N_9612);
and U10949 (N_10949,N_8542,N_8414);
xnor U10950 (N_10950,N_8156,N_9079);
xnor U10951 (N_10951,N_8249,N_8316);
or U10952 (N_10952,N_8330,N_9397);
and U10953 (N_10953,N_9911,N_8992);
or U10954 (N_10954,N_9658,N_8866);
or U10955 (N_10955,N_8387,N_8016);
nand U10956 (N_10956,N_8861,N_8809);
nand U10957 (N_10957,N_9287,N_8019);
or U10958 (N_10958,N_9894,N_9212);
or U10959 (N_10959,N_8765,N_9065);
and U10960 (N_10960,N_9605,N_8843);
and U10961 (N_10961,N_9880,N_8979);
or U10962 (N_10962,N_8964,N_9185);
nand U10963 (N_10963,N_8642,N_8568);
xor U10964 (N_10964,N_8691,N_8510);
nand U10965 (N_10965,N_9063,N_8824);
or U10966 (N_10966,N_9996,N_8530);
and U10967 (N_10967,N_9245,N_8826);
nand U10968 (N_10968,N_9747,N_9595);
nand U10969 (N_10969,N_9710,N_9051);
and U10970 (N_10970,N_9708,N_9769);
nor U10971 (N_10971,N_8453,N_9549);
or U10972 (N_10972,N_9005,N_9192);
or U10973 (N_10973,N_8129,N_9550);
and U10974 (N_10974,N_9884,N_8139);
or U10975 (N_10975,N_9270,N_8040);
or U10976 (N_10976,N_8241,N_9188);
or U10977 (N_10977,N_9141,N_9682);
nor U10978 (N_10978,N_8367,N_8720);
nand U10979 (N_10979,N_8370,N_8004);
and U10980 (N_10980,N_8942,N_9169);
nor U10981 (N_10981,N_9990,N_8015);
or U10982 (N_10982,N_8224,N_9866);
and U10983 (N_10983,N_9139,N_8091);
nand U10984 (N_10984,N_9061,N_9877);
nor U10985 (N_10985,N_9806,N_9518);
or U10986 (N_10986,N_9952,N_9743);
nand U10987 (N_10987,N_8631,N_9887);
nand U10988 (N_10988,N_8993,N_9142);
xor U10989 (N_10989,N_9385,N_9089);
nand U10990 (N_10990,N_9341,N_9500);
and U10991 (N_10991,N_8647,N_9716);
or U10992 (N_10992,N_8051,N_8834);
and U10993 (N_10993,N_9480,N_8252);
nor U10994 (N_10994,N_8046,N_8038);
nor U10995 (N_10995,N_9321,N_8567);
or U10996 (N_10996,N_9214,N_8127);
nor U10997 (N_10997,N_9277,N_8218);
and U10998 (N_10998,N_9885,N_8788);
and U10999 (N_10999,N_8279,N_9725);
nor U11000 (N_11000,N_8598,N_8896);
nor U11001 (N_11001,N_9351,N_9849);
nand U11002 (N_11002,N_8715,N_9355);
xnor U11003 (N_11003,N_8548,N_8831);
nor U11004 (N_11004,N_9996,N_9654);
and U11005 (N_11005,N_9912,N_9849);
or U11006 (N_11006,N_8001,N_8669);
and U11007 (N_11007,N_9056,N_8813);
nor U11008 (N_11008,N_8061,N_8015);
or U11009 (N_11009,N_8006,N_9771);
nor U11010 (N_11010,N_8368,N_8785);
or U11011 (N_11011,N_8749,N_9298);
nand U11012 (N_11012,N_8963,N_8687);
nor U11013 (N_11013,N_8877,N_9673);
nor U11014 (N_11014,N_8375,N_9377);
and U11015 (N_11015,N_9881,N_9671);
or U11016 (N_11016,N_8413,N_8184);
or U11017 (N_11017,N_8472,N_9415);
nor U11018 (N_11018,N_8574,N_8183);
xnor U11019 (N_11019,N_9213,N_9652);
xnor U11020 (N_11020,N_9530,N_8508);
or U11021 (N_11021,N_9790,N_9571);
nor U11022 (N_11022,N_8547,N_9282);
nor U11023 (N_11023,N_9233,N_8761);
nor U11024 (N_11024,N_9082,N_8948);
nand U11025 (N_11025,N_8842,N_8835);
or U11026 (N_11026,N_9474,N_8010);
nand U11027 (N_11027,N_9606,N_9554);
nor U11028 (N_11028,N_8201,N_9642);
and U11029 (N_11029,N_9045,N_8418);
nand U11030 (N_11030,N_9751,N_9017);
and U11031 (N_11031,N_8068,N_8774);
nand U11032 (N_11032,N_9357,N_8861);
or U11033 (N_11033,N_8700,N_8020);
xnor U11034 (N_11034,N_9248,N_9590);
and U11035 (N_11035,N_9267,N_8904);
and U11036 (N_11036,N_8313,N_8859);
nand U11037 (N_11037,N_9841,N_8719);
or U11038 (N_11038,N_9664,N_9762);
nand U11039 (N_11039,N_9374,N_8993);
xnor U11040 (N_11040,N_9466,N_8751);
or U11041 (N_11041,N_9136,N_8648);
xnor U11042 (N_11042,N_9993,N_8758);
xnor U11043 (N_11043,N_9441,N_9423);
nand U11044 (N_11044,N_8327,N_9676);
or U11045 (N_11045,N_8091,N_9761);
or U11046 (N_11046,N_9585,N_9077);
and U11047 (N_11047,N_8428,N_8497);
nand U11048 (N_11048,N_9149,N_8965);
or U11049 (N_11049,N_9729,N_9809);
or U11050 (N_11050,N_9863,N_9317);
and U11051 (N_11051,N_8946,N_9606);
and U11052 (N_11052,N_8904,N_8201);
nand U11053 (N_11053,N_8583,N_8320);
nand U11054 (N_11054,N_9017,N_9407);
xor U11055 (N_11055,N_9887,N_9872);
or U11056 (N_11056,N_9444,N_9599);
nand U11057 (N_11057,N_8381,N_8264);
nor U11058 (N_11058,N_8726,N_9914);
or U11059 (N_11059,N_9199,N_9316);
or U11060 (N_11060,N_9875,N_8039);
or U11061 (N_11061,N_8223,N_8652);
nor U11062 (N_11062,N_8566,N_8555);
or U11063 (N_11063,N_8250,N_9181);
nand U11064 (N_11064,N_9252,N_9483);
and U11065 (N_11065,N_9515,N_8559);
and U11066 (N_11066,N_9391,N_9718);
nor U11067 (N_11067,N_9985,N_8686);
nand U11068 (N_11068,N_9035,N_8009);
or U11069 (N_11069,N_9953,N_9570);
nor U11070 (N_11070,N_9926,N_8541);
and U11071 (N_11071,N_9765,N_9048);
and U11072 (N_11072,N_9557,N_8242);
nor U11073 (N_11073,N_8215,N_9184);
nand U11074 (N_11074,N_8440,N_8425);
nand U11075 (N_11075,N_9563,N_8172);
nor U11076 (N_11076,N_8540,N_8179);
or U11077 (N_11077,N_8535,N_8903);
nand U11078 (N_11078,N_9812,N_9697);
nand U11079 (N_11079,N_8773,N_8420);
or U11080 (N_11080,N_8468,N_8429);
or U11081 (N_11081,N_9574,N_8357);
and U11082 (N_11082,N_8345,N_8617);
or U11083 (N_11083,N_8408,N_8208);
nand U11084 (N_11084,N_8020,N_9962);
or U11085 (N_11085,N_9161,N_9140);
nor U11086 (N_11086,N_8410,N_8082);
nor U11087 (N_11087,N_9866,N_9104);
or U11088 (N_11088,N_8520,N_9425);
nand U11089 (N_11089,N_8545,N_9639);
xor U11090 (N_11090,N_9883,N_9606);
nor U11091 (N_11091,N_8073,N_9930);
or U11092 (N_11092,N_9599,N_8481);
nor U11093 (N_11093,N_9694,N_8674);
nand U11094 (N_11094,N_8056,N_9922);
nor U11095 (N_11095,N_8828,N_9249);
nor U11096 (N_11096,N_9605,N_8504);
and U11097 (N_11097,N_8687,N_9109);
and U11098 (N_11098,N_8274,N_9037);
nor U11099 (N_11099,N_8898,N_8752);
or U11100 (N_11100,N_9479,N_8694);
nand U11101 (N_11101,N_9768,N_8097);
and U11102 (N_11102,N_8986,N_9017);
or U11103 (N_11103,N_8656,N_9843);
or U11104 (N_11104,N_9388,N_8624);
xor U11105 (N_11105,N_9794,N_8454);
nand U11106 (N_11106,N_9550,N_9445);
nor U11107 (N_11107,N_9691,N_9253);
nor U11108 (N_11108,N_9952,N_9162);
or U11109 (N_11109,N_8864,N_8103);
nand U11110 (N_11110,N_8519,N_9147);
nand U11111 (N_11111,N_9368,N_8626);
nand U11112 (N_11112,N_9617,N_8461);
nor U11113 (N_11113,N_9324,N_8205);
nor U11114 (N_11114,N_9304,N_8928);
and U11115 (N_11115,N_9212,N_9611);
and U11116 (N_11116,N_9093,N_9817);
and U11117 (N_11117,N_9777,N_8903);
nand U11118 (N_11118,N_8850,N_8398);
nor U11119 (N_11119,N_9736,N_8626);
or U11120 (N_11120,N_9211,N_8597);
nor U11121 (N_11121,N_8855,N_8985);
or U11122 (N_11122,N_8856,N_9026);
and U11123 (N_11123,N_8007,N_8543);
and U11124 (N_11124,N_9958,N_8295);
nand U11125 (N_11125,N_8828,N_8387);
and U11126 (N_11126,N_8812,N_8976);
or U11127 (N_11127,N_9052,N_8289);
nand U11128 (N_11128,N_9025,N_9671);
or U11129 (N_11129,N_8997,N_8521);
and U11130 (N_11130,N_8317,N_9537);
xnor U11131 (N_11131,N_9217,N_8860);
and U11132 (N_11132,N_8097,N_8596);
and U11133 (N_11133,N_8345,N_9570);
and U11134 (N_11134,N_9964,N_8900);
and U11135 (N_11135,N_8271,N_8241);
nor U11136 (N_11136,N_9446,N_8956);
and U11137 (N_11137,N_8479,N_8222);
nor U11138 (N_11138,N_9518,N_8144);
nor U11139 (N_11139,N_8337,N_9934);
xnor U11140 (N_11140,N_9941,N_9015);
nand U11141 (N_11141,N_8147,N_8829);
nand U11142 (N_11142,N_8974,N_9987);
and U11143 (N_11143,N_9961,N_8824);
xnor U11144 (N_11144,N_8610,N_9470);
nand U11145 (N_11145,N_9853,N_9997);
or U11146 (N_11146,N_9859,N_8116);
and U11147 (N_11147,N_9624,N_9609);
nand U11148 (N_11148,N_9093,N_9746);
and U11149 (N_11149,N_8593,N_9381);
xnor U11150 (N_11150,N_8362,N_8135);
nand U11151 (N_11151,N_9710,N_8059);
and U11152 (N_11152,N_8358,N_9701);
nand U11153 (N_11153,N_8447,N_9421);
and U11154 (N_11154,N_8919,N_8330);
or U11155 (N_11155,N_9778,N_8175);
or U11156 (N_11156,N_8385,N_8773);
nand U11157 (N_11157,N_8256,N_9805);
and U11158 (N_11158,N_8780,N_9849);
or U11159 (N_11159,N_9227,N_9931);
nand U11160 (N_11160,N_8059,N_9462);
xor U11161 (N_11161,N_8261,N_9147);
or U11162 (N_11162,N_8912,N_8860);
nand U11163 (N_11163,N_9694,N_9530);
xor U11164 (N_11164,N_8598,N_8358);
and U11165 (N_11165,N_8102,N_9220);
and U11166 (N_11166,N_9850,N_8713);
nor U11167 (N_11167,N_8945,N_9854);
xor U11168 (N_11168,N_9730,N_9997);
nand U11169 (N_11169,N_8819,N_9803);
or U11170 (N_11170,N_9974,N_9420);
or U11171 (N_11171,N_8095,N_9202);
xor U11172 (N_11172,N_9763,N_9935);
nor U11173 (N_11173,N_9964,N_9564);
and U11174 (N_11174,N_8241,N_8801);
or U11175 (N_11175,N_9398,N_8052);
nor U11176 (N_11176,N_9591,N_8387);
nor U11177 (N_11177,N_9438,N_8528);
nand U11178 (N_11178,N_9712,N_9575);
and U11179 (N_11179,N_9051,N_8027);
nor U11180 (N_11180,N_9458,N_8688);
nand U11181 (N_11181,N_8435,N_8527);
or U11182 (N_11182,N_8858,N_8886);
nand U11183 (N_11183,N_9250,N_9766);
nand U11184 (N_11184,N_8132,N_9555);
nor U11185 (N_11185,N_8601,N_9891);
or U11186 (N_11186,N_8610,N_9964);
nor U11187 (N_11187,N_9498,N_8802);
nand U11188 (N_11188,N_8758,N_9624);
xor U11189 (N_11189,N_8571,N_9657);
and U11190 (N_11190,N_9446,N_8561);
nand U11191 (N_11191,N_8468,N_9431);
nand U11192 (N_11192,N_9391,N_8380);
or U11193 (N_11193,N_8723,N_9155);
nand U11194 (N_11194,N_8770,N_9904);
and U11195 (N_11195,N_9975,N_8169);
xor U11196 (N_11196,N_9300,N_9122);
and U11197 (N_11197,N_9474,N_8820);
nor U11198 (N_11198,N_9727,N_8789);
and U11199 (N_11199,N_9243,N_9291);
nand U11200 (N_11200,N_8625,N_8783);
and U11201 (N_11201,N_9631,N_8751);
and U11202 (N_11202,N_9874,N_8413);
xor U11203 (N_11203,N_9444,N_8920);
and U11204 (N_11204,N_8909,N_9874);
xor U11205 (N_11205,N_8696,N_9270);
nor U11206 (N_11206,N_9018,N_8030);
nand U11207 (N_11207,N_9496,N_8606);
nand U11208 (N_11208,N_8719,N_9654);
or U11209 (N_11209,N_8182,N_9392);
nor U11210 (N_11210,N_9190,N_9514);
or U11211 (N_11211,N_9989,N_9896);
nand U11212 (N_11212,N_9745,N_8647);
or U11213 (N_11213,N_9256,N_9813);
nand U11214 (N_11214,N_8373,N_8928);
and U11215 (N_11215,N_9833,N_8047);
and U11216 (N_11216,N_9223,N_9632);
nand U11217 (N_11217,N_8744,N_9410);
or U11218 (N_11218,N_8449,N_9823);
nand U11219 (N_11219,N_8150,N_9317);
nor U11220 (N_11220,N_8017,N_9991);
nand U11221 (N_11221,N_8372,N_9551);
xor U11222 (N_11222,N_9209,N_8386);
nor U11223 (N_11223,N_9379,N_9319);
nand U11224 (N_11224,N_8757,N_9178);
nand U11225 (N_11225,N_9608,N_9857);
and U11226 (N_11226,N_9371,N_9749);
nor U11227 (N_11227,N_9468,N_8297);
xnor U11228 (N_11228,N_8332,N_9775);
and U11229 (N_11229,N_9097,N_8512);
nor U11230 (N_11230,N_8205,N_8979);
and U11231 (N_11231,N_9134,N_9797);
or U11232 (N_11232,N_9501,N_8097);
xnor U11233 (N_11233,N_8886,N_8014);
and U11234 (N_11234,N_9482,N_8775);
or U11235 (N_11235,N_8772,N_9339);
nand U11236 (N_11236,N_9126,N_8865);
or U11237 (N_11237,N_9469,N_8311);
nand U11238 (N_11238,N_9733,N_9334);
nor U11239 (N_11239,N_9425,N_8855);
and U11240 (N_11240,N_8875,N_8465);
or U11241 (N_11241,N_8016,N_9836);
or U11242 (N_11242,N_9791,N_8617);
nand U11243 (N_11243,N_8654,N_8203);
and U11244 (N_11244,N_9355,N_9181);
nand U11245 (N_11245,N_9657,N_8674);
nor U11246 (N_11246,N_9940,N_9095);
xnor U11247 (N_11247,N_8794,N_9371);
nand U11248 (N_11248,N_8837,N_8017);
or U11249 (N_11249,N_8430,N_9355);
xnor U11250 (N_11250,N_9597,N_8484);
xnor U11251 (N_11251,N_9472,N_8295);
xor U11252 (N_11252,N_9271,N_8635);
and U11253 (N_11253,N_8885,N_9077);
or U11254 (N_11254,N_9258,N_9357);
and U11255 (N_11255,N_8384,N_9338);
and U11256 (N_11256,N_9860,N_9674);
nand U11257 (N_11257,N_8049,N_9900);
xor U11258 (N_11258,N_9292,N_8391);
or U11259 (N_11259,N_9871,N_9167);
nand U11260 (N_11260,N_8367,N_8590);
or U11261 (N_11261,N_9550,N_9456);
and U11262 (N_11262,N_8683,N_8161);
nor U11263 (N_11263,N_9195,N_9338);
and U11264 (N_11264,N_9187,N_8243);
or U11265 (N_11265,N_9363,N_8185);
nand U11266 (N_11266,N_9479,N_8534);
or U11267 (N_11267,N_9955,N_8624);
or U11268 (N_11268,N_9792,N_8860);
nor U11269 (N_11269,N_9282,N_9560);
xor U11270 (N_11270,N_9379,N_9745);
or U11271 (N_11271,N_8424,N_8595);
or U11272 (N_11272,N_9642,N_8815);
nor U11273 (N_11273,N_8880,N_8484);
nor U11274 (N_11274,N_9853,N_8266);
nor U11275 (N_11275,N_8600,N_8223);
nor U11276 (N_11276,N_8385,N_8506);
or U11277 (N_11277,N_8436,N_9514);
nand U11278 (N_11278,N_9328,N_9329);
xnor U11279 (N_11279,N_8362,N_8109);
and U11280 (N_11280,N_9737,N_9074);
nor U11281 (N_11281,N_9483,N_9717);
nand U11282 (N_11282,N_8454,N_9925);
nand U11283 (N_11283,N_9192,N_9877);
nor U11284 (N_11284,N_9854,N_8201);
nand U11285 (N_11285,N_8231,N_8302);
nor U11286 (N_11286,N_8068,N_8335);
or U11287 (N_11287,N_9316,N_9348);
nor U11288 (N_11288,N_8621,N_8608);
xnor U11289 (N_11289,N_8647,N_8411);
nor U11290 (N_11290,N_8397,N_9367);
or U11291 (N_11291,N_8747,N_9335);
nand U11292 (N_11292,N_8674,N_8587);
and U11293 (N_11293,N_8948,N_8126);
nor U11294 (N_11294,N_9525,N_8415);
or U11295 (N_11295,N_9671,N_9728);
nand U11296 (N_11296,N_9505,N_9239);
or U11297 (N_11297,N_9966,N_9008);
or U11298 (N_11298,N_8128,N_9906);
nand U11299 (N_11299,N_9735,N_8136);
nor U11300 (N_11300,N_9934,N_8993);
nor U11301 (N_11301,N_8492,N_9560);
nand U11302 (N_11302,N_8964,N_8200);
and U11303 (N_11303,N_8758,N_9226);
nor U11304 (N_11304,N_9064,N_9596);
or U11305 (N_11305,N_9134,N_9525);
nor U11306 (N_11306,N_9780,N_8691);
nor U11307 (N_11307,N_9176,N_8137);
xnor U11308 (N_11308,N_9974,N_9538);
nand U11309 (N_11309,N_9185,N_9949);
or U11310 (N_11310,N_8788,N_9453);
and U11311 (N_11311,N_9471,N_8306);
nor U11312 (N_11312,N_8030,N_8649);
nor U11313 (N_11313,N_8113,N_8777);
or U11314 (N_11314,N_9308,N_8763);
xnor U11315 (N_11315,N_9575,N_9959);
and U11316 (N_11316,N_9878,N_9475);
nor U11317 (N_11317,N_8043,N_8706);
nor U11318 (N_11318,N_9618,N_8600);
and U11319 (N_11319,N_9848,N_8134);
nand U11320 (N_11320,N_9548,N_8586);
or U11321 (N_11321,N_9971,N_8548);
or U11322 (N_11322,N_8086,N_8672);
nor U11323 (N_11323,N_9410,N_8080);
nand U11324 (N_11324,N_9050,N_8373);
or U11325 (N_11325,N_8959,N_9716);
nor U11326 (N_11326,N_9454,N_9018);
or U11327 (N_11327,N_8728,N_8379);
xor U11328 (N_11328,N_8514,N_8160);
nor U11329 (N_11329,N_8113,N_8078);
nand U11330 (N_11330,N_9343,N_9801);
and U11331 (N_11331,N_8902,N_8392);
or U11332 (N_11332,N_9471,N_8159);
nor U11333 (N_11333,N_9860,N_9863);
and U11334 (N_11334,N_8497,N_8427);
nand U11335 (N_11335,N_8020,N_9145);
or U11336 (N_11336,N_8980,N_8186);
nand U11337 (N_11337,N_8810,N_9891);
and U11338 (N_11338,N_9643,N_9578);
or U11339 (N_11339,N_9408,N_8558);
or U11340 (N_11340,N_8425,N_9461);
nor U11341 (N_11341,N_8949,N_8602);
nand U11342 (N_11342,N_8141,N_8550);
or U11343 (N_11343,N_8538,N_8063);
and U11344 (N_11344,N_9820,N_9501);
xor U11345 (N_11345,N_9241,N_9439);
and U11346 (N_11346,N_9326,N_9748);
nand U11347 (N_11347,N_9790,N_9877);
xnor U11348 (N_11348,N_8472,N_8744);
or U11349 (N_11349,N_8877,N_9628);
or U11350 (N_11350,N_8634,N_9632);
nor U11351 (N_11351,N_9348,N_8114);
or U11352 (N_11352,N_9731,N_9564);
nand U11353 (N_11353,N_9747,N_8032);
nor U11354 (N_11354,N_9464,N_9545);
and U11355 (N_11355,N_8186,N_9873);
nand U11356 (N_11356,N_8897,N_9243);
nand U11357 (N_11357,N_9903,N_8588);
or U11358 (N_11358,N_8324,N_8212);
and U11359 (N_11359,N_9921,N_9275);
nand U11360 (N_11360,N_8905,N_9016);
or U11361 (N_11361,N_8244,N_9083);
and U11362 (N_11362,N_8136,N_9792);
nor U11363 (N_11363,N_9015,N_9598);
or U11364 (N_11364,N_8311,N_8534);
xor U11365 (N_11365,N_9968,N_8699);
and U11366 (N_11366,N_9732,N_8611);
and U11367 (N_11367,N_8852,N_9313);
or U11368 (N_11368,N_9077,N_9001);
nor U11369 (N_11369,N_8474,N_9225);
and U11370 (N_11370,N_9495,N_8526);
nand U11371 (N_11371,N_8632,N_8090);
xnor U11372 (N_11372,N_9480,N_8355);
nor U11373 (N_11373,N_8920,N_9331);
and U11374 (N_11374,N_9478,N_9142);
and U11375 (N_11375,N_9416,N_9593);
and U11376 (N_11376,N_9699,N_8507);
nand U11377 (N_11377,N_9352,N_9264);
nand U11378 (N_11378,N_9546,N_9183);
or U11379 (N_11379,N_9500,N_9790);
nor U11380 (N_11380,N_8109,N_9664);
and U11381 (N_11381,N_9119,N_8346);
nand U11382 (N_11382,N_9468,N_9678);
and U11383 (N_11383,N_8884,N_8398);
nand U11384 (N_11384,N_9752,N_9847);
and U11385 (N_11385,N_8831,N_8072);
or U11386 (N_11386,N_8785,N_8112);
or U11387 (N_11387,N_8037,N_8600);
nand U11388 (N_11388,N_9126,N_8439);
nor U11389 (N_11389,N_8311,N_9982);
nor U11390 (N_11390,N_8224,N_9747);
and U11391 (N_11391,N_9156,N_8258);
and U11392 (N_11392,N_9210,N_8759);
or U11393 (N_11393,N_8217,N_8282);
nand U11394 (N_11394,N_9260,N_9158);
or U11395 (N_11395,N_8966,N_9986);
or U11396 (N_11396,N_8779,N_8438);
or U11397 (N_11397,N_8936,N_8883);
and U11398 (N_11398,N_9224,N_8034);
and U11399 (N_11399,N_8644,N_9204);
or U11400 (N_11400,N_8316,N_9776);
nand U11401 (N_11401,N_8016,N_8928);
or U11402 (N_11402,N_8232,N_9340);
nor U11403 (N_11403,N_9987,N_9543);
nor U11404 (N_11404,N_8177,N_9719);
xor U11405 (N_11405,N_8610,N_9692);
nor U11406 (N_11406,N_8955,N_9258);
xnor U11407 (N_11407,N_9436,N_8004);
and U11408 (N_11408,N_8100,N_9614);
nor U11409 (N_11409,N_8931,N_8948);
and U11410 (N_11410,N_9170,N_8969);
nor U11411 (N_11411,N_9213,N_9469);
nor U11412 (N_11412,N_9115,N_8798);
nor U11413 (N_11413,N_8510,N_8757);
or U11414 (N_11414,N_9982,N_9750);
and U11415 (N_11415,N_8386,N_8776);
or U11416 (N_11416,N_8859,N_9626);
nand U11417 (N_11417,N_9820,N_8098);
and U11418 (N_11418,N_9665,N_9782);
nand U11419 (N_11419,N_8752,N_8785);
nor U11420 (N_11420,N_8754,N_8703);
and U11421 (N_11421,N_8966,N_9457);
nor U11422 (N_11422,N_8156,N_9406);
and U11423 (N_11423,N_8680,N_8159);
and U11424 (N_11424,N_8605,N_8158);
nor U11425 (N_11425,N_8428,N_9089);
nor U11426 (N_11426,N_9687,N_9748);
nand U11427 (N_11427,N_9157,N_8750);
xnor U11428 (N_11428,N_9333,N_9002);
or U11429 (N_11429,N_9008,N_8223);
nor U11430 (N_11430,N_9118,N_9656);
nand U11431 (N_11431,N_9646,N_8460);
nand U11432 (N_11432,N_9463,N_8847);
nor U11433 (N_11433,N_9080,N_8783);
or U11434 (N_11434,N_8483,N_8452);
or U11435 (N_11435,N_8205,N_8675);
and U11436 (N_11436,N_9566,N_9473);
nor U11437 (N_11437,N_8263,N_8534);
nand U11438 (N_11438,N_8347,N_9615);
nand U11439 (N_11439,N_9413,N_9078);
xnor U11440 (N_11440,N_8765,N_8852);
and U11441 (N_11441,N_8376,N_9624);
nand U11442 (N_11442,N_8693,N_9542);
nand U11443 (N_11443,N_8560,N_9335);
and U11444 (N_11444,N_9272,N_8353);
nand U11445 (N_11445,N_8395,N_8140);
nor U11446 (N_11446,N_9140,N_8176);
nor U11447 (N_11447,N_8968,N_8410);
nand U11448 (N_11448,N_8897,N_8636);
and U11449 (N_11449,N_8864,N_9555);
or U11450 (N_11450,N_8808,N_8122);
nand U11451 (N_11451,N_8792,N_8941);
and U11452 (N_11452,N_9669,N_9254);
nor U11453 (N_11453,N_9826,N_9890);
xor U11454 (N_11454,N_8675,N_9639);
nand U11455 (N_11455,N_9520,N_9554);
and U11456 (N_11456,N_8157,N_8108);
and U11457 (N_11457,N_8957,N_8007);
nand U11458 (N_11458,N_8762,N_8057);
xor U11459 (N_11459,N_9625,N_9339);
xor U11460 (N_11460,N_8453,N_9777);
and U11461 (N_11461,N_9904,N_8536);
nand U11462 (N_11462,N_8155,N_9294);
or U11463 (N_11463,N_8209,N_9745);
xnor U11464 (N_11464,N_9155,N_9217);
xor U11465 (N_11465,N_9681,N_8386);
or U11466 (N_11466,N_9594,N_9670);
nor U11467 (N_11467,N_9568,N_9913);
and U11468 (N_11468,N_8971,N_9326);
xnor U11469 (N_11469,N_9003,N_9276);
or U11470 (N_11470,N_8837,N_9268);
nand U11471 (N_11471,N_9088,N_9103);
and U11472 (N_11472,N_9525,N_8675);
and U11473 (N_11473,N_8367,N_9250);
nor U11474 (N_11474,N_9424,N_9869);
nor U11475 (N_11475,N_9862,N_8097);
nand U11476 (N_11476,N_9659,N_9937);
nand U11477 (N_11477,N_8417,N_8168);
xor U11478 (N_11478,N_8686,N_8702);
xor U11479 (N_11479,N_8512,N_8798);
or U11480 (N_11480,N_9778,N_9844);
xor U11481 (N_11481,N_9161,N_9825);
nand U11482 (N_11482,N_8776,N_9789);
and U11483 (N_11483,N_8875,N_8482);
nor U11484 (N_11484,N_9196,N_9876);
nor U11485 (N_11485,N_8109,N_8341);
nand U11486 (N_11486,N_9211,N_8742);
or U11487 (N_11487,N_9830,N_8084);
or U11488 (N_11488,N_9016,N_9754);
and U11489 (N_11489,N_8487,N_8770);
and U11490 (N_11490,N_9993,N_9719);
and U11491 (N_11491,N_9046,N_8445);
or U11492 (N_11492,N_8789,N_9333);
nor U11493 (N_11493,N_8128,N_8226);
nor U11494 (N_11494,N_8601,N_9326);
or U11495 (N_11495,N_8208,N_9045);
nor U11496 (N_11496,N_9339,N_8964);
or U11497 (N_11497,N_8352,N_9061);
nand U11498 (N_11498,N_8813,N_8525);
nor U11499 (N_11499,N_9276,N_9165);
nor U11500 (N_11500,N_8764,N_8865);
and U11501 (N_11501,N_9337,N_8943);
and U11502 (N_11502,N_8163,N_9944);
or U11503 (N_11503,N_9840,N_9649);
nand U11504 (N_11504,N_9478,N_9679);
and U11505 (N_11505,N_9713,N_8422);
and U11506 (N_11506,N_9191,N_9514);
or U11507 (N_11507,N_8293,N_8817);
and U11508 (N_11508,N_9815,N_8107);
nor U11509 (N_11509,N_9214,N_8525);
nor U11510 (N_11510,N_8946,N_9785);
or U11511 (N_11511,N_9645,N_9120);
nor U11512 (N_11512,N_8631,N_8221);
nor U11513 (N_11513,N_9616,N_8226);
nand U11514 (N_11514,N_8494,N_9794);
nor U11515 (N_11515,N_9578,N_8245);
nand U11516 (N_11516,N_9808,N_9699);
nand U11517 (N_11517,N_9488,N_8218);
and U11518 (N_11518,N_9773,N_9763);
nor U11519 (N_11519,N_9458,N_8243);
nand U11520 (N_11520,N_8734,N_8978);
nor U11521 (N_11521,N_9848,N_8326);
xnor U11522 (N_11522,N_8122,N_9631);
nand U11523 (N_11523,N_8239,N_9816);
nor U11524 (N_11524,N_8051,N_8959);
xnor U11525 (N_11525,N_8481,N_8633);
and U11526 (N_11526,N_9689,N_8992);
nor U11527 (N_11527,N_9792,N_8344);
nor U11528 (N_11528,N_9468,N_9679);
nor U11529 (N_11529,N_9060,N_9924);
and U11530 (N_11530,N_8520,N_8689);
or U11531 (N_11531,N_8107,N_8638);
nand U11532 (N_11532,N_9688,N_8195);
xor U11533 (N_11533,N_9279,N_8665);
and U11534 (N_11534,N_8630,N_9114);
nand U11535 (N_11535,N_8145,N_8603);
and U11536 (N_11536,N_8828,N_8287);
or U11537 (N_11537,N_8244,N_8499);
and U11538 (N_11538,N_9625,N_8203);
and U11539 (N_11539,N_9541,N_8611);
nand U11540 (N_11540,N_9200,N_9671);
nor U11541 (N_11541,N_9087,N_9686);
and U11542 (N_11542,N_8779,N_8287);
nand U11543 (N_11543,N_9126,N_8365);
nor U11544 (N_11544,N_9131,N_9603);
nand U11545 (N_11545,N_8977,N_9050);
or U11546 (N_11546,N_8367,N_8994);
nand U11547 (N_11547,N_8812,N_9845);
nor U11548 (N_11548,N_9681,N_9727);
or U11549 (N_11549,N_9460,N_8540);
nor U11550 (N_11550,N_9433,N_8639);
nor U11551 (N_11551,N_8194,N_8285);
and U11552 (N_11552,N_8861,N_8611);
nor U11553 (N_11553,N_8294,N_8259);
or U11554 (N_11554,N_9269,N_9659);
or U11555 (N_11555,N_9665,N_9803);
or U11556 (N_11556,N_8619,N_8682);
xnor U11557 (N_11557,N_9100,N_8547);
and U11558 (N_11558,N_8235,N_8136);
nand U11559 (N_11559,N_9024,N_8513);
nor U11560 (N_11560,N_8571,N_9334);
and U11561 (N_11561,N_8838,N_9058);
nor U11562 (N_11562,N_9772,N_8632);
or U11563 (N_11563,N_9339,N_9508);
nand U11564 (N_11564,N_8609,N_8830);
and U11565 (N_11565,N_9322,N_9581);
or U11566 (N_11566,N_9050,N_8597);
nor U11567 (N_11567,N_8862,N_8159);
and U11568 (N_11568,N_9853,N_9828);
and U11569 (N_11569,N_8822,N_9080);
and U11570 (N_11570,N_9266,N_9006);
nand U11571 (N_11571,N_9762,N_9552);
nor U11572 (N_11572,N_9985,N_9142);
and U11573 (N_11573,N_8141,N_8549);
nand U11574 (N_11574,N_9149,N_9336);
or U11575 (N_11575,N_8185,N_9733);
nor U11576 (N_11576,N_8561,N_9484);
nor U11577 (N_11577,N_8019,N_8304);
nor U11578 (N_11578,N_8444,N_9599);
nor U11579 (N_11579,N_9021,N_8890);
or U11580 (N_11580,N_9394,N_9847);
nand U11581 (N_11581,N_9774,N_8255);
nor U11582 (N_11582,N_9131,N_8182);
and U11583 (N_11583,N_8413,N_8066);
nand U11584 (N_11584,N_8823,N_9127);
nand U11585 (N_11585,N_8661,N_8775);
nand U11586 (N_11586,N_8122,N_9094);
nor U11587 (N_11587,N_8726,N_9189);
nor U11588 (N_11588,N_9714,N_9488);
nor U11589 (N_11589,N_8298,N_9439);
and U11590 (N_11590,N_9751,N_8703);
nor U11591 (N_11591,N_9440,N_8858);
nor U11592 (N_11592,N_8245,N_8700);
or U11593 (N_11593,N_9065,N_9459);
nor U11594 (N_11594,N_9257,N_8756);
and U11595 (N_11595,N_9142,N_8580);
nor U11596 (N_11596,N_8621,N_8894);
nand U11597 (N_11597,N_8028,N_9212);
or U11598 (N_11598,N_9125,N_8850);
and U11599 (N_11599,N_8150,N_9057);
and U11600 (N_11600,N_8565,N_8900);
xor U11601 (N_11601,N_9545,N_9640);
nor U11602 (N_11602,N_8657,N_8246);
nor U11603 (N_11603,N_8671,N_8377);
xnor U11604 (N_11604,N_9321,N_9839);
xnor U11605 (N_11605,N_8785,N_8195);
or U11606 (N_11606,N_9949,N_8139);
xor U11607 (N_11607,N_9270,N_8024);
nand U11608 (N_11608,N_9101,N_8112);
nand U11609 (N_11609,N_8300,N_9725);
nor U11610 (N_11610,N_8479,N_9458);
or U11611 (N_11611,N_9767,N_9286);
and U11612 (N_11612,N_8558,N_8120);
and U11613 (N_11613,N_8912,N_9937);
nand U11614 (N_11614,N_9281,N_8269);
nand U11615 (N_11615,N_8652,N_9118);
nor U11616 (N_11616,N_8644,N_8971);
nor U11617 (N_11617,N_8278,N_9682);
and U11618 (N_11618,N_9417,N_8186);
or U11619 (N_11619,N_8419,N_9426);
nor U11620 (N_11620,N_8497,N_8695);
nor U11621 (N_11621,N_9901,N_9688);
and U11622 (N_11622,N_9567,N_8561);
or U11623 (N_11623,N_8025,N_9807);
nand U11624 (N_11624,N_8651,N_9006);
xnor U11625 (N_11625,N_9494,N_9047);
nor U11626 (N_11626,N_9751,N_8426);
nand U11627 (N_11627,N_9975,N_9743);
nor U11628 (N_11628,N_8822,N_9415);
nor U11629 (N_11629,N_8932,N_9090);
or U11630 (N_11630,N_8424,N_9696);
nor U11631 (N_11631,N_8592,N_9665);
nor U11632 (N_11632,N_9672,N_8311);
or U11633 (N_11633,N_9499,N_9879);
nor U11634 (N_11634,N_9274,N_8446);
xnor U11635 (N_11635,N_9741,N_8769);
or U11636 (N_11636,N_8489,N_9451);
or U11637 (N_11637,N_9694,N_8349);
or U11638 (N_11638,N_8387,N_8138);
nand U11639 (N_11639,N_9644,N_8684);
xor U11640 (N_11640,N_9084,N_8269);
nand U11641 (N_11641,N_8176,N_8820);
or U11642 (N_11642,N_9297,N_8558);
nor U11643 (N_11643,N_8958,N_8708);
nand U11644 (N_11644,N_9869,N_8563);
or U11645 (N_11645,N_9683,N_8571);
or U11646 (N_11646,N_9268,N_9906);
nor U11647 (N_11647,N_9610,N_9722);
and U11648 (N_11648,N_9663,N_8050);
nor U11649 (N_11649,N_8255,N_9305);
nand U11650 (N_11650,N_9261,N_9817);
nor U11651 (N_11651,N_8967,N_8635);
or U11652 (N_11652,N_9051,N_9792);
or U11653 (N_11653,N_8690,N_9164);
xnor U11654 (N_11654,N_8433,N_8384);
nor U11655 (N_11655,N_8834,N_8354);
nor U11656 (N_11656,N_9484,N_9004);
and U11657 (N_11657,N_8364,N_8807);
nand U11658 (N_11658,N_9615,N_9863);
nor U11659 (N_11659,N_9880,N_8796);
xor U11660 (N_11660,N_9562,N_9872);
xnor U11661 (N_11661,N_8448,N_8292);
nor U11662 (N_11662,N_8081,N_9020);
and U11663 (N_11663,N_8132,N_9164);
or U11664 (N_11664,N_8979,N_9913);
nor U11665 (N_11665,N_8383,N_9441);
nor U11666 (N_11666,N_9521,N_8237);
or U11667 (N_11667,N_9231,N_9384);
nor U11668 (N_11668,N_9351,N_8061);
or U11669 (N_11669,N_8229,N_8074);
nand U11670 (N_11670,N_8720,N_8795);
nand U11671 (N_11671,N_8333,N_8760);
nand U11672 (N_11672,N_8190,N_9772);
nand U11673 (N_11673,N_9435,N_9634);
xnor U11674 (N_11674,N_8534,N_8539);
nand U11675 (N_11675,N_9590,N_9833);
and U11676 (N_11676,N_8487,N_8799);
nand U11677 (N_11677,N_8552,N_8625);
or U11678 (N_11678,N_8396,N_8283);
or U11679 (N_11679,N_9207,N_9766);
nand U11680 (N_11680,N_8462,N_8328);
nor U11681 (N_11681,N_9666,N_9153);
or U11682 (N_11682,N_8427,N_8690);
and U11683 (N_11683,N_9914,N_8831);
and U11684 (N_11684,N_9889,N_8197);
or U11685 (N_11685,N_8072,N_8849);
nand U11686 (N_11686,N_9594,N_9798);
nand U11687 (N_11687,N_8408,N_8685);
nand U11688 (N_11688,N_9744,N_9838);
or U11689 (N_11689,N_8504,N_8332);
nand U11690 (N_11690,N_9483,N_9507);
and U11691 (N_11691,N_9063,N_9266);
xnor U11692 (N_11692,N_8176,N_8036);
nor U11693 (N_11693,N_8141,N_9107);
or U11694 (N_11694,N_8606,N_9879);
or U11695 (N_11695,N_8027,N_9642);
or U11696 (N_11696,N_9638,N_8928);
or U11697 (N_11697,N_8963,N_9214);
nor U11698 (N_11698,N_9558,N_9229);
and U11699 (N_11699,N_9393,N_9103);
xor U11700 (N_11700,N_9119,N_9993);
nor U11701 (N_11701,N_9538,N_9135);
and U11702 (N_11702,N_9074,N_9282);
and U11703 (N_11703,N_8641,N_8533);
xor U11704 (N_11704,N_9999,N_9883);
xnor U11705 (N_11705,N_8906,N_9978);
nor U11706 (N_11706,N_9043,N_8516);
or U11707 (N_11707,N_8311,N_9424);
nor U11708 (N_11708,N_9525,N_9169);
xnor U11709 (N_11709,N_9422,N_9083);
and U11710 (N_11710,N_9742,N_9344);
nand U11711 (N_11711,N_9802,N_9481);
nand U11712 (N_11712,N_9759,N_8942);
nor U11713 (N_11713,N_9997,N_9048);
nand U11714 (N_11714,N_8648,N_8454);
nand U11715 (N_11715,N_8569,N_8179);
nor U11716 (N_11716,N_8239,N_8673);
xor U11717 (N_11717,N_8973,N_9191);
and U11718 (N_11718,N_8382,N_8832);
and U11719 (N_11719,N_9163,N_8137);
xor U11720 (N_11720,N_8166,N_9487);
xnor U11721 (N_11721,N_9539,N_9514);
or U11722 (N_11722,N_8578,N_8426);
or U11723 (N_11723,N_8675,N_8078);
and U11724 (N_11724,N_9429,N_9822);
and U11725 (N_11725,N_8847,N_9501);
nand U11726 (N_11726,N_9756,N_8673);
nor U11727 (N_11727,N_8908,N_8266);
nor U11728 (N_11728,N_9970,N_9682);
or U11729 (N_11729,N_9067,N_8400);
or U11730 (N_11730,N_9284,N_8883);
nand U11731 (N_11731,N_8081,N_9136);
nand U11732 (N_11732,N_9366,N_9498);
or U11733 (N_11733,N_8617,N_8579);
or U11734 (N_11734,N_9773,N_9750);
or U11735 (N_11735,N_8364,N_9518);
nand U11736 (N_11736,N_8894,N_9253);
nor U11737 (N_11737,N_9729,N_9119);
and U11738 (N_11738,N_8532,N_8946);
or U11739 (N_11739,N_8627,N_9598);
or U11740 (N_11740,N_9924,N_9167);
and U11741 (N_11741,N_9608,N_9521);
nor U11742 (N_11742,N_8791,N_9582);
nand U11743 (N_11743,N_8855,N_9586);
and U11744 (N_11744,N_8676,N_8867);
and U11745 (N_11745,N_9655,N_9848);
or U11746 (N_11746,N_9974,N_9568);
or U11747 (N_11747,N_9960,N_8586);
nand U11748 (N_11748,N_8802,N_9978);
xnor U11749 (N_11749,N_8670,N_8426);
nor U11750 (N_11750,N_9674,N_9166);
nor U11751 (N_11751,N_8149,N_8323);
xnor U11752 (N_11752,N_9176,N_9087);
nand U11753 (N_11753,N_8880,N_9421);
xor U11754 (N_11754,N_9893,N_8696);
nor U11755 (N_11755,N_8530,N_9925);
nand U11756 (N_11756,N_8206,N_8939);
nor U11757 (N_11757,N_9279,N_8185);
or U11758 (N_11758,N_9159,N_8622);
or U11759 (N_11759,N_9977,N_9380);
nor U11760 (N_11760,N_9490,N_8245);
nor U11761 (N_11761,N_9317,N_8684);
or U11762 (N_11762,N_8206,N_9810);
nor U11763 (N_11763,N_8469,N_8021);
and U11764 (N_11764,N_9382,N_8585);
or U11765 (N_11765,N_8671,N_9522);
nor U11766 (N_11766,N_8096,N_9877);
nand U11767 (N_11767,N_9888,N_9483);
nand U11768 (N_11768,N_8876,N_8086);
and U11769 (N_11769,N_9016,N_9007);
nor U11770 (N_11770,N_8144,N_8894);
and U11771 (N_11771,N_9240,N_8019);
nor U11772 (N_11772,N_9772,N_9765);
xnor U11773 (N_11773,N_8784,N_9457);
nor U11774 (N_11774,N_9994,N_8444);
or U11775 (N_11775,N_9289,N_9496);
nor U11776 (N_11776,N_9160,N_8631);
nand U11777 (N_11777,N_8471,N_9368);
or U11778 (N_11778,N_9549,N_9374);
nand U11779 (N_11779,N_9271,N_8293);
nor U11780 (N_11780,N_8797,N_8852);
nor U11781 (N_11781,N_9854,N_9202);
or U11782 (N_11782,N_8734,N_8862);
or U11783 (N_11783,N_9558,N_9409);
and U11784 (N_11784,N_8548,N_9695);
or U11785 (N_11785,N_8693,N_8080);
or U11786 (N_11786,N_8685,N_9100);
and U11787 (N_11787,N_9321,N_9483);
nand U11788 (N_11788,N_8686,N_9488);
or U11789 (N_11789,N_9396,N_9913);
xnor U11790 (N_11790,N_8713,N_9710);
and U11791 (N_11791,N_9801,N_8598);
nand U11792 (N_11792,N_9779,N_9864);
or U11793 (N_11793,N_8494,N_9992);
xnor U11794 (N_11794,N_9549,N_9545);
or U11795 (N_11795,N_8657,N_9629);
or U11796 (N_11796,N_8804,N_8343);
and U11797 (N_11797,N_9606,N_9970);
or U11798 (N_11798,N_8649,N_8680);
and U11799 (N_11799,N_8620,N_9927);
or U11800 (N_11800,N_8306,N_8783);
or U11801 (N_11801,N_8215,N_8115);
nor U11802 (N_11802,N_8977,N_8707);
nor U11803 (N_11803,N_8269,N_9658);
and U11804 (N_11804,N_8198,N_9776);
nand U11805 (N_11805,N_8434,N_9713);
nor U11806 (N_11806,N_9324,N_8646);
xnor U11807 (N_11807,N_9818,N_8026);
and U11808 (N_11808,N_9190,N_9136);
nand U11809 (N_11809,N_8331,N_8213);
nand U11810 (N_11810,N_9193,N_9343);
or U11811 (N_11811,N_9353,N_8988);
or U11812 (N_11812,N_8126,N_9017);
and U11813 (N_11813,N_9016,N_8397);
nand U11814 (N_11814,N_9927,N_9180);
nor U11815 (N_11815,N_8518,N_9017);
or U11816 (N_11816,N_8374,N_8403);
and U11817 (N_11817,N_9899,N_9816);
and U11818 (N_11818,N_8165,N_9194);
or U11819 (N_11819,N_9202,N_8063);
and U11820 (N_11820,N_9366,N_8572);
and U11821 (N_11821,N_9407,N_8073);
nor U11822 (N_11822,N_9788,N_9005);
or U11823 (N_11823,N_8781,N_8185);
or U11824 (N_11824,N_9185,N_9328);
nand U11825 (N_11825,N_8291,N_8666);
and U11826 (N_11826,N_9135,N_8375);
xor U11827 (N_11827,N_9799,N_8150);
xnor U11828 (N_11828,N_9924,N_8307);
and U11829 (N_11829,N_9443,N_8653);
and U11830 (N_11830,N_9405,N_8989);
or U11831 (N_11831,N_8164,N_8706);
nor U11832 (N_11832,N_8925,N_8687);
nor U11833 (N_11833,N_9725,N_8510);
nor U11834 (N_11834,N_8320,N_9576);
and U11835 (N_11835,N_8976,N_8231);
or U11836 (N_11836,N_9199,N_9872);
nor U11837 (N_11837,N_8085,N_9828);
and U11838 (N_11838,N_8762,N_8962);
xor U11839 (N_11839,N_8131,N_9809);
or U11840 (N_11840,N_9892,N_9835);
nor U11841 (N_11841,N_9647,N_9229);
and U11842 (N_11842,N_9697,N_9824);
or U11843 (N_11843,N_9006,N_9662);
or U11844 (N_11844,N_9340,N_9636);
or U11845 (N_11845,N_9601,N_9335);
nor U11846 (N_11846,N_8167,N_8375);
nand U11847 (N_11847,N_8958,N_8848);
nor U11848 (N_11848,N_9332,N_9500);
and U11849 (N_11849,N_9983,N_8334);
or U11850 (N_11850,N_9333,N_8116);
nand U11851 (N_11851,N_9526,N_9099);
nand U11852 (N_11852,N_9602,N_9402);
or U11853 (N_11853,N_8364,N_8479);
and U11854 (N_11854,N_9222,N_9185);
xor U11855 (N_11855,N_8145,N_8202);
nor U11856 (N_11856,N_9522,N_9660);
xnor U11857 (N_11857,N_8616,N_9266);
or U11858 (N_11858,N_8919,N_9382);
and U11859 (N_11859,N_8978,N_9409);
or U11860 (N_11860,N_9354,N_9699);
or U11861 (N_11861,N_9791,N_8084);
nand U11862 (N_11862,N_9644,N_8922);
nor U11863 (N_11863,N_8789,N_8322);
or U11864 (N_11864,N_9160,N_8125);
and U11865 (N_11865,N_9111,N_8685);
or U11866 (N_11866,N_8166,N_8984);
nor U11867 (N_11867,N_8423,N_8936);
and U11868 (N_11868,N_8048,N_9355);
nor U11869 (N_11869,N_8510,N_9303);
nor U11870 (N_11870,N_8893,N_8898);
nand U11871 (N_11871,N_8906,N_9278);
and U11872 (N_11872,N_8150,N_9238);
and U11873 (N_11873,N_8842,N_8775);
xor U11874 (N_11874,N_9784,N_9147);
or U11875 (N_11875,N_9149,N_8794);
nand U11876 (N_11876,N_8277,N_8253);
and U11877 (N_11877,N_8464,N_9989);
and U11878 (N_11878,N_9889,N_9658);
and U11879 (N_11879,N_9347,N_9912);
nor U11880 (N_11880,N_9833,N_8494);
or U11881 (N_11881,N_8495,N_8180);
and U11882 (N_11882,N_8772,N_9462);
nor U11883 (N_11883,N_9734,N_9766);
nand U11884 (N_11884,N_9487,N_9935);
or U11885 (N_11885,N_8594,N_8931);
or U11886 (N_11886,N_9828,N_9579);
nor U11887 (N_11887,N_8732,N_9396);
nor U11888 (N_11888,N_9751,N_8499);
or U11889 (N_11889,N_9725,N_9181);
xnor U11890 (N_11890,N_8830,N_9727);
nand U11891 (N_11891,N_9417,N_9028);
or U11892 (N_11892,N_9112,N_8168);
or U11893 (N_11893,N_8068,N_8951);
or U11894 (N_11894,N_9937,N_8349);
nor U11895 (N_11895,N_8936,N_9881);
nand U11896 (N_11896,N_8191,N_9557);
xor U11897 (N_11897,N_9884,N_8232);
xor U11898 (N_11898,N_8138,N_9130);
nand U11899 (N_11899,N_9713,N_9104);
nand U11900 (N_11900,N_9178,N_9844);
nor U11901 (N_11901,N_8197,N_9895);
or U11902 (N_11902,N_8815,N_8728);
and U11903 (N_11903,N_9190,N_9267);
and U11904 (N_11904,N_8078,N_9666);
nand U11905 (N_11905,N_8536,N_9027);
nand U11906 (N_11906,N_8554,N_8749);
and U11907 (N_11907,N_8707,N_8831);
nor U11908 (N_11908,N_8318,N_8141);
or U11909 (N_11909,N_9331,N_8640);
nor U11910 (N_11910,N_8118,N_9712);
nand U11911 (N_11911,N_9648,N_9092);
and U11912 (N_11912,N_8776,N_8208);
nand U11913 (N_11913,N_9160,N_8011);
and U11914 (N_11914,N_8408,N_8433);
nor U11915 (N_11915,N_9482,N_9396);
nand U11916 (N_11916,N_8040,N_9385);
xnor U11917 (N_11917,N_8709,N_9529);
or U11918 (N_11918,N_9878,N_9592);
and U11919 (N_11919,N_9472,N_8465);
or U11920 (N_11920,N_8360,N_9377);
nand U11921 (N_11921,N_8201,N_9575);
nand U11922 (N_11922,N_9353,N_9956);
nand U11923 (N_11923,N_9239,N_8243);
or U11924 (N_11924,N_8445,N_8249);
xor U11925 (N_11925,N_8059,N_8439);
nor U11926 (N_11926,N_8858,N_9438);
nand U11927 (N_11927,N_8813,N_8247);
xor U11928 (N_11928,N_8756,N_8268);
xor U11929 (N_11929,N_8312,N_8112);
or U11930 (N_11930,N_9099,N_9478);
or U11931 (N_11931,N_9077,N_8751);
xnor U11932 (N_11932,N_9818,N_9661);
and U11933 (N_11933,N_9246,N_9940);
nand U11934 (N_11934,N_9024,N_8283);
or U11935 (N_11935,N_9936,N_9273);
nor U11936 (N_11936,N_9062,N_9953);
nand U11937 (N_11937,N_9179,N_9747);
and U11938 (N_11938,N_9017,N_8331);
or U11939 (N_11939,N_9488,N_8351);
nor U11940 (N_11940,N_9956,N_9957);
nand U11941 (N_11941,N_8198,N_9228);
nor U11942 (N_11942,N_9718,N_8623);
nor U11943 (N_11943,N_9641,N_9044);
and U11944 (N_11944,N_8687,N_9537);
and U11945 (N_11945,N_8815,N_9032);
and U11946 (N_11946,N_9887,N_8634);
xor U11947 (N_11947,N_9725,N_9559);
nand U11948 (N_11948,N_8912,N_8204);
nor U11949 (N_11949,N_8762,N_9061);
or U11950 (N_11950,N_9972,N_9324);
and U11951 (N_11951,N_8045,N_9863);
nand U11952 (N_11952,N_8919,N_8316);
nor U11953 (N_11953,N_8770,N_8386);
or U11954 (N_11954,N_8510,N_9545);
nor U11955 (N_11955,N_8597,N_8363);
or U11956 (N_11956,N_8242,N_8009);
nor U11957 (N_11957,N_9695,N_9867);
nand U11958 (N_11958,N_8760,N_9337);
nand U11959 (N_11959,N_9223,N_9121);
nor U11960 (N_11960,N_8451,N_8467);
xnor U11961 (N_11961,N_8115,N_9079);
nor U11962 (N_11962,N_9566,N_9832);
nand U11963 (N_11963,N_8697,N_8222);
nor U11964 (N_11964,N_9211,N_9340);
nor U11965 (N_11965,N_9406,N_8084);
and U11966 (N_11966,N_8001,N_9604);
nand U11967 (N_11967,N_8008,N_9971);
nand U11968 (N_11968,N_9190,N_9597);
nor U11969 (N_11969,N_8116,N_9816);
nor U11970 (N_11970,N_9817,N_8775);
nor U11971 (N_11971,N_9890,N_9124);
nor U11972 (N_11972,N_8124,N_8078);
nor U11973 (N_11973,N_9274,N_8019);
and U11974 (N_11974,N_9489,N_8757);
and U11975 (N_11975,N_8267,N_9814);
nor U11976 (N_11976,N_8755,N_8284);
nor U11977 (N_11977,N_9859,N_8511);
and U11978 (N_11978,N_8341,N_8523);
nand U11979 (N_11979,N_8262,N_8680);
and U11980 (N_11980,N_9857,N_9325);
or U11981 (N_11981,N_9196,N_8783);
nor U11982 (N_11982,N_8867,N_9064);
nand U11983 (N_11983,N_8428,N_8684);
and U11984 (N_11984,N_9691,N_8373);
nor U11985 (N_11985,N_8989,N_9482);
nor U11986 (N_11986,N_8711,N_9199);
nor U11987 (N_11987,N_8649,N_9731);
xnor U11988 (N_11988,N_8217,N_9403);
and U11989 (N_11989,N_8017,N_9810);
or U11990 (N_11990,N_8504,N_9287);
or U11991 (N_11991,N_8983,N_9485);
nor U11992 (N_11992,N_8596,N_9726);
or U11993 (N_11993,N_9529,N_9080);
nand U11994 (N_11994,N_8337,N_8883);
xnor U11995 (N_11995,N_8550,N_8091);
or U11996 (N_11996,N_9754,N_9054);
nand U11997 (N_11997,N_8150,N_8201);
or U11998 (N_11998,N_9659,N_8122);
nand U11999 (N_11999,N_9714,N_8815);
or U12000 (N_12000,N_10276,N_10042);
nor U12001 (N_12001,N_11758,N_11224);
nor U12002 (N_12002,N_11153,N_11111);
and U12003 (N_12003,N_11609,N_10333);
nand U12004 (N_12004,N_10208,N_11946);
and U12005 (N_12005,N_11030,N_10409);
nor U12006 (N_12006,N_10257,N_11721);
or U12007 (N_12007,N_10590,N_10559);
and U12008 (N_12008,N_11966,N_10800);
and U12009 (N_12009,N_11212,N_11831);
nor U12010 (N_12010,N_11062,N_10776);
nor U12011 (N_12011,N_10361,N_11216);
and U12012 (N_12012,N_10269,N_10150);
or U12013 (N_12013,N_11565,N_10859);
nand U12014 (N_12014,N_10445,N_11431);
xor U12015 (N_12015,N_10071,N_11045);
and U12016 (N_12016,N_10373,N_11717);
nor U12017 (N_12017,N_10787,N_11108);
or U12018 (N_12018,N_10526,N_11747);
or U12019 (N_12019,N_11652,N_11907);
and U12020 (N_12020,N_10006,N_11147);
and U12021 (N_12021,N_11607,N_10053);
nand U12022 (N_12022,N_11630,N_11067);
or U12023 (N_12023,N_10392,N_10791);
nand U12024 (N_12024,N_11398,N_11736);
nor U12025 (N_12025,N_11188,N_10539);
nor U12026 (N_12026,N_10789,N_10075);
nand U12027 (N_12027,N_10946,N_11750);
nand U12028 (N_12028,N_10380,N_11463);
nand U12029 (N_12029,N_11848,N_10721);
nor U12030 (N_12030,N_11491,N_10144);
and U12031 (N_12031,N_11932,N_10556);
nand U12032 (N_12032,N_11438,N_10083);
and U12033 (N_12033,N_11873,N_10616);
and U12034 (N_12034,N_11315,N_11994);
and U12035 (N_12035,N_11625,N_11540);
and U12036 (N_12036,N_11584,N_10436);
or U12037 (N_12037,N_10295,N_11432);
or U12038 (N_12038,N_10716,N_10076);
xnor U12039 (N_12039,N_11175,N_10466);
nor U12040 (N_12040,N_10981,N_10775);
nand U12041 (N_12041,N_10762,N_10290);
xor U12042 (N_12042,N_10665,N_11031);
and U12043 (N_12043,N_10266,N_10822);
and U12044 (N_12044,N_11751,N_11354);
or U12045 (N_12045,N_11569,N_11744);
nand U12046 (N_12046,N_10655,N_11768);
xor U12047 (N_12047,N_10989,N_11096);
or U12048 (N_12048,N_10210,N_10214);
nand U12049 (N_12049,N_10914,N_11702);
xnor U12050 (N_12050,N_10272,N_10154);
or U12051 (N_12051,N_10085,N_11316);
or U12052 (N_12052,N_11012,N_11197);
nor U12053 (N_12053,N_10934,N_11020);
or U12054 (N_12054,N_10522,N_11528);
xor U12055 (N_12055,N_11566,N_10799);
xor U12056 (N_12056,N_10956,N_11228);
nor U12057 (N_12057,N_10782,N_11856);
and U12058 (N_12058,N_11833,N_11749);
xnor U12059 (N_12059,N_11169,N_11809);
and U12060 (N_12060,N_10704,N_11213);
nand U12061 (N_12061,N_11631,N_11259);
or U12062 (N_12062,N_10843,N_10564);
nand U12063 (N_12063,N_10215,N_11962);
and U12064 (N_12064,N_11104,N_10766);
and U12065 (N_12065,N_11040,N_10813);
nand U12066 (N_12066,N_10286,N_11454);
or U12067 (N_12067,N_11414,N_11507);
nand U12068 (N_12068,N_11332,N_11254);
or U12069 (N_12069,N_11824,N_11255);
nor U12070 (N_12070,N_11514,N_11065);
and U12071 (N_12071,N_10719,N_10759);
nand U12072 (N_12072,N_10217,N_10474);
nor U12073 (N_12073,N_11193,N_11064);
or U12074 (N_12074,N_11992,N_10429);
nor U12075 (N_12075,N_11982,N_11035);
xor U12076 (N_12076,N_11655,N_11286);
nor U12077 (N_12077,N_11754,N_10932);
nor U12078 (N_12078,N_10430,N_11157);
nor U12079 (N_12079,N_11861,N_10434);
or U12080 (N_12080,N_11371,N_11384);
and U12081 (N_12081,N_10901,N_10519);
or U12082 (N_12082,N_10896,N_10585);
or U12083 (N_12083,N_10143,N_11564);
and U12084 (N_12084,N_10457,N_10335);
nor U12085 (N_12085,N_10754,N_10236);
nand U12086 (N_12086,N_11386,N_10726);
nor U12087 (N_12087,N_11123,N_11364);
or U12088 (N_12088,N_11196,N_10199);
nor U12089 (N_12089,N_11801,N_10611);
and U12090 (N_12090,N_10820,N_11502);
or U12091 (N_12091,N_10012,N_10640);
and U12092 (N_12092,N_10666,N_10057);
nand U12093 (N_12093,N_10991,N_10378);
and U12094 (N_12094,N_11931,N_10988);
or U12095 (N_12095,N_11874,N_10234);
or U12096 (N_12096,N_11636,N_10173);
nor U12097 (N_12097,N_10493,N_11855);
nor U12098 (N_12098,N_10853,N_11958);
xor U12099 (N_12099,N_10770,N_10740);
nor U12100 (N_12100,N_11303,N_11843);
nor U12101 (N_12101,N_10366,N_10596);
and U12102 (N_12102,N_11296,N_11428);
and U12103 (N_12103,N_10259,N_10542);
nor U12104 (N_12104,N_10984,N_10861);
nand U12105 (N_12105,N_10900,N_10305);
nor U12106 (N_12106,N_10648,N_11603);
nor U12107 (N_12107,N_11529,N_10043);
and U12108 (N_12108,N_10692,N_11248);
nor U12109 (N_12109,N_10803,N_11974);
and U12110 (N_12110,N_10937,N_11764);
and U12111 (N_12111,N_11077,N_11021);
nand U12112 (N_12112,N_10252,N_11671);
nor U12113 (N_12113,N_11722,N_11408);
xor U12114 (N_12114,N_10685,N_11234);
or U12115 (N_12115,N_10352,N_10709);
and U12116 (N_12116,N_10348,N_10182);
or U12117 (N_12117,N_11489,N_11544);
and U12118 (N_12118,N_11681,N_11849);
and U12119 (N_12119,N_11588,N_11929);
nand U12120 (N_12120,N_11484,N_11927);
nand U12121 (N_12121,N_10203,N_11322);
and U12122 (N_12122,N_10487,N_10880);
nand U12123 (N_12123,N_10131,N_10662);
and U12124 (N_12124,N_10906,N_10218);
and U12125 (N_12125,N_11699,N_10541);
nand U12126 (N_12126,N_10889,N_10595);
nor U12127 (N_12127,N_11079,N_10239);
and U12128 (N_12128,N_10110,N_10245);
nor U12129 (N_12129,N_11301,N_11028);
and U12130 (N_12130,N_10060,N_10494);
and U12131 (N_12131,N_10465,N_10367);
or U12132 (N_12132,N_10400,N_11290);
nor U12133 (N_12133,N_11445,N_11081);
and U12134 (N_12134,N_10138,N_10983);
nor U12135 (N_12135,N_11710,N_11146);
nand U12136 (N_12136,N_10582,N_11916);
and U12137 (N_12137,N_11601,N_11942);
xor U12138 (N_12138,N_10146,N_10788);
or U12139 (N_12139,N_10231,N_10694);
xnor U12140 (N_12140,N_11888,N_10960);
nor U12141 (N_12141,N_11014,N_11378);
and U12142 (N_12142,N_11898,N_10032);
nor U12143 (N_12143,N_10273,N_11466);
nor U12144 (N_12144,N_11732,N_10279);
xor U12145 (N_12145,N_11583,N_11957);
or U12146 (N_12146,N_10314,N_11359);
or U12147 (N_12147,N_11651,N_11106);
and U12148 (N_12148,N_11708,N_11906);
or U12149 (N_12149,N_10503,N_11127);
and U12150 (N_12150,N_11353,N_10477);
and U12151 (N_12151,N_11349,N_10261);
nand U12152 (N_12152,N_11317,N_10927);
xnor U12153 (N_12153,N_11665,N_10003);
nand U12154 (N_12154,N_11662,N_10402);
nand U12155 (N_12155,N_11572,N_11447);
nand U12156 (N_12156,N_10454,N_11415);
nand U12157 (N_12157,N_11339,N_10793);
and U12158 (N_12158,N_10962,N_11404);
xor U12159 (N_12159,N_11046,N_11239);
nor U12160 (N_12160,N_10077,N_10625);
and U12161 (N_12161,N_10224,N_11120);
or U12162 (N_12162,N_10451,N_10472);
or U12163 (N_12163,N_10354,N_11490);
nand U12164 (N_12164,N_11069,N_10656);
and U12165 (N_12165,N_11939,N_10478);
or U12166 (N_12166,N_11073,N_11458);
nand U12167 (N_12167,N_10365,N_10289);
nor U12168 (N_12168,N_11811,N_10317);
or U12169 (N_12169,N_10773,N_10769);
and U12170 (N_12170,N_11177,N_10415);
or U12171 (N_12171,N_10175,N_10055);
nor U12172 (N_12172,N_11306,N_10115);
nand U12173 (N_12173,N_10159,N_11117);
or U12174 (N_12174,N_11219,N_10836);
nor U12175 (N_12175,N_10578,N_11760);
nand U12176 (N_12176,N_11766,N_10284);
and U12177 (N_12177,N_11853,N_11495);
nand U12178 (N_12178,N_10007,N_11869);
nand U12179 (N_12179,N_11273,N_11941);
and U12180 (N_12180,N_11791,N_11739);
nor U12181 (N_12181,N_10809,N_10216);
nand U12182 (N_12182,N_10690,N_10184);
and U12183 (N_12183,N_10912,N_11728);
or U12184 (N_12184,N_10802,N_11820);
and U12185 (N_12185,N_10262,N_10686);
and U12186 (N_12186,N_11264,N_10019);
nand U12187 (N_12187,N_11094,N_10976);
xor U12188 (N_12188,N_10768,N_11761);
nor U12189 (N_12189,N_11167,N_10928);
nand U12190 (N_12190,N_10490,N_11468);
nor U12191 (N_12191,N_11084,N_11598);
or U12192 (N_12192,N_11538,N_11176);
xor U12193 (N_12193,N_11150,N_11510);
nor U12194 (N_12194,N_11712,N_10369);
or U12195 (N_12195,N_11960,N_11052);
nand U12196 (N_12196,N_11166,N_11901);
nand U12197 (N_12197,N_10291,N_11780);
and U12198 (N_12198,N_10479,N_11344);
and U12199 (N_12199,N_10950,N_10021);
nand U12200 (N_12200,N_10411,N_10117);
nand U12201 (N_12201,N_11406,N_11852);
or U12202 (N_12202,N_11646,N_10260);
and U12203 (N_12203,N_10185,N_10078);
nand U12204 (N_12204,N_10650,N_10223);
or U12205 (N_12205,N_10090,N_10840);
nand U12206 (N_12206,N_10674,N_11629);
and U12207 (N_12207,N_10486,N_10283);
and U12208 (N_12208,N_10767,N_11740);
and U12209 (N_12209,N_10221,N_10095);
or U12210 (N_12210,N_11661,N_10842);
nand U12211 (N_12211,N_10838,N_11334);
xor U12212 (N_12212,N_10974,N_11218);
nand U12213 (N_12213,N_10913,N_10362);
nand U12214 (N_12214,N_11304,N_10013);
xor U12215 (N_12215,N_10325,N_11782);
nand U12216 (N_12216,N_11112,N_10328);
nand U12217 (N_12217,N_11101,N_11793);
nor U12218 (N_12218,N_11837,N_11003);
or U12219 (N_12219,N_11433,N_11834);
nor U12220 (N_12220,N_11361,N_10041);
or U12221 (N_12221,N_10387,N_10644);
and U12222 (N_12222,N_11987,N_10610);
and U12223 (N_12223,N_10498,N_10638);
or U12224 (N_12224,N_10763,N_11309);
or U12225 (N_12225,N_11692,N_11242);
nand U12226 (N_12226,N_11473,N_10841);
nor U12227 (N_12227,N_11327,N_10020);
or U12228 (N_12228,N_10620,N_11562);
nor U12229 (N_12229,N_10693,N_10751);
or U12230 (N_12230,N_10732,N_10601);
or U12231 (N_12231,N_10160,N_10702);
xor U12232 (N_12232,N_10292,N_11493);
or U12233 (N_12233,N_10275,N_11482);
or U12234 (N_12234,N_11536,N_10464);
nor U12235 (N_12235,N_11614,N_10147);
or U12236 (N_12236,N_11924,N_10460);
and U12237 (N_12237,N_10222,N_10165);
nand U12238 (N_12238,N_11311,N_11779);
nor U12239 (N_12239,N_10848,N_11642);
nand U12240 (N_12240,N_10864,N_10895);
nor U12241 (N_12241,N_10296,N_10897);
and U12242 (N_12242,N_10183,N_11753);
or U12243 (N_12243,N_11733,N_11241);
or U12244 (N_12244,N_11783,N_10850);
nor U12245 (N_12245,N_10112,N_10379);
nor U12246 (N_12246,N_10845,N_11523);
nor U12247 (N_12247,N_11172,N_10384);
nand U12248 (N_12248,N_10450,N_11318);
nor U12249 (N_12249,N_11345,N_11295);
nor U12250 (N_12250,N_10546,N_11302);
nor U12251 (N_12251,N_11757,N_11815);
or U12252 (N_12252,N_10197,N_10660);
or U12253 (N_12253,N_10811,N_10715);
nand U12254 (N_12254,N_10098,N_10758);
and U12255 (N_12255,N_11517,N_11719);
nand U12256 (N_12256,N_11862,N_11501);
or U12257 (N_12257,N_10080,N_11223);
and U12258 (N_12258,N_11356,N_10152);
and U12259 (N_12259,N_11525,N_11180);
nor U12260 (N_12260,N_11455,N_10229);
and U12261 (N_12261,N_10672,N_11503);
nor U12262 (N_12262,N_10018,N_11822);
nand U12263 (N_12263,N_10826,N_11679);
or U12264 (N_12264,N_10534,N_10764);
nand U12265 (N_12265,N_11478,N_11179);
nand U12266 (N_12266,N_11397,N_10485);
or U12267 (N_12267,N_10200,N_10922);
nor U12268 (N_12268,N_10047,N_10461);
xor U12269 (N_12269,N_11706,N_10658);
or U12270 (N_12270,N_11784,N_10920);
nor U12271 (N_12271,N_11969,N_10393);
or U12272 (N_12272,N_11578,N_10860);
or U12273 (N_12273,N_11881,N_10476);
nand U12274 (N_12274,N_10600,N_11152);
or U12275 (N_12275,N_11441,N_11628);
nand U12276 (N_12276,N_11026,N_10285);
and U12277 (N_12277,N_11838,N_10254);
xnor U12278 (N_12278,N_10492,N_10313);
or U12279 (N_12279,N_10647,N_11477);
and U12280 (N_12280,N_11400,N_10324);
nand U12281 (N_12281,N_11451,N_10207);
nand U12282 (N_12282,N_11618,N_10684);
xnor U12283 (N_12283,N_11896,N_11854);
or U12284 (N_12284,N_10894,N_11649);
and U12285 (N_12285,N_10968,N_11335);
nand U12286 (N_12286,N_11707,N_11570);
or U12287 (N_12287,N_10780,N_11277);
or U12288 (N_12288,N_10375,N_10915);
or U12289 (N_12289,N_10433,N_11430);
or U12290 (N_12290,N_10998,N_11648);
and U12291 (N_12291,N_10548,N_10323);
nor U12292 (N_12292,N_10688,N_10502);
nor U12293 (N_12293,N_10263,N_10888);
nor U12294 (N_12294,N_11922,N_11110);
and U12295 (N_12295,N_10488,N_11682);
and U12296 (N_12296,N_10550,N_11936);
nor U12297 (N_12297,N_10796,N_11637);
nand U12298 (N_12298,N_11990,N_11421);
or U12299 (N_12299,N_11413,N_10441);
nand U12300 (N_12300,N_11006,N_11229);
and U12301 (N_12301,N_11289,N_10587);
nand U12302 (N_12302,N_11043,N_10343);
nor U12303 (N_12303,N_10404,N_11158);
nor U12304 (N_12304,N_10288,N_10986);
nor U12305 (N_12305,N_11975,N_10442);
nor U12306 (N_12306,N_10421,N_11324);
or U12307 (N_12307,N_10753,N_11579);
or U12308 (N_12308,N_11352,N_11799);
or U12309 (N_12309,N_11456,N_10281);
xnor U12310 (N_12310,N_11920,N_10881);
nand U12311 (N_12311,N_11847,N_10171);
and U12312 (N_12312,N_10680,N_10985);
or U12313 (N_12313,N_11943,N_10372);
nand U12314 (N_12314,N_10642,N_10280);
or U12315 (N_12315,N_10667,N_10801);
and U12316 (N_12316,N_10708,N_10654);
xnor U12317 (N_12317,N_10696,N_10355);
nand U12318 (N_12318,N_11586,N_10576);
or U12319 (N_12319,N_11806,N_11004);
nand U12320 (N_12320,N_10449,N_11659);
nand U12321 (N_12321,N_10997,N_10815);
or U12322 (N_12322,N_11392,N_10471);
or U12323 (N_12323,N_10537,N_11705);
xnor U12324 (N_12324,N_11965,N_10760);
and U12325 (N_12325,N_11981,N_11553);
and U12326 (N_12326,N_10456,N_10311);
or U12327 (N_12327,N_11836,N_10856);
nor U12328 (N_12328,N_10562,N_11530);
xnor U12329 (N_12329,N_11971,N_11870);
xor U12330 (N_12330,N_11019,N_10874);
and U12331 (N_12331,N_11961,N_10785);
xnor U12332 (N_12332,N_11996,N_10959);
nand U12333 (N_12333,N_11919,N_10581);
nand U12334 (N_12334,N_11238,N_11686);
nand U12335 (N_12335,N_10855,N_11554);
and U12336 (N_12336,N_10570,N_10942);
or U12337 (N_12337,N_10887,N_10423);
nor U12338 (N_12338,N_10196,N_11235);
and U12339 (N_12339,N_11312,N_11159);
or U12340 (N_12340,N_11674,N_11623);
nand U12341 (N_12341,N_10011,N_11243);
nand U12342 (N_12342,N_11527,N_11333);
nand U12343 (N_12343,N_11812,N_11908);
xnor U12344 (N_12344,N_11305,N_10613);
and U12345 (N_12345,N_11660,N_10302);
and U12346 (N_12346,N_10882,N_11376);
and U12347 (N_12347,N_11367,N_10586);
and U12348 (N_12348,N_11912,N_10381);
or U12349 (N_12349,N_10432,N_11670);
nand U12350 (N_12350,N_11860,N_11231);
nand U12351 (N_12351,N_10700,N_11198);
nor U12352 (N_12352,N_11685,N_11174);
and U12353 (N_12353,N_11443,N_11276);
or U12354 (N_12354,N_10268,N_10253);
nor U12355 (N_12355,N_11145,N_10706);
nor U12356 (N_12356,N_11545,N_10885);
nor U12357 (N_12357,N_11464,N_11844);
nor U12358 (N_12358,N_11913,N_11829);
or U12359 (N_12359,N_10063,N_11805);
xor U12360 (N_12360,N_11055,N_11369);
xnor U12361 (N_12361,N_11083,N_10963);
or U12362 (N_12362,N_10635,N_10250);
nand U12363 (N_12363,N_10405,N_11797);
nor U12364 (N_12364,N_10385,N_11561);
or U12365 (N_12365,N_11313,N_10446);
xnor U12366 (N_12366,N_10058,N_10247);
nand U12367 (N_12367,N_11446,N_11675);
nor U12368 (N_12368,N_11270,N_10149);
or U12369 (N_12369,N_11730,N_11267);
nor U12370 (N_12370,N_11085,N_10641);
nor U12371 (N_12371,N_10204,N_10037);
and U12372 (N_12372,N_10004,N_11669);
nand U12373 (N_12373,N_10459,N_10308);
and U12374 (N_12374,N_10558,N_11186);
and U12375 (N_12375,N_11115,N_11887);
nor U12376 (N_12376,N_10926,N_10500);
and U12377 (N_12377,N_10825,N_10024);
or U12378 (N_12378,N_11729,N_11752);
nor U12379 (N_12379,N_11391,N_10228);
nor U12380 (N_12380,N_10322,N_11155);
or U12381 (N_12381,N_11192,N_11709);
nor U12382 (N_12382,N_10816,N_10341);
or U12383 (N_12383,N_11057,N_10359);
or U12384 (N_12384,N_11059,N_10748);
nor U12385 (N_12385,N_10427,N_10108);
nor U12386 (N_12386,N_10046,N_10969);
and U12387 (N_12387,N_10121,N_11534);
nand U12388 (N_12388,N_10639,N_10230);
nand U12389 (N_12389,N_10072,N_10863);
nand U12390 (N_12390,N_10109,N_10784);
nor U12391 (N_12391,N_10818,N_10734);
nand U12392 (N_12392,N_10332,N_10670);
and U12393 (N_12393,N_11785,N_10101);
and U12394 (N_12394,N_10572,N_11892);
and U12395 (N_12395,N_11066,N_10844);
nor U12396 (N_12396,N_10870,N_10049);
and U12397 (N_12397,N_10722,N_11471);
nand U12398 (N_12398,N_10307,N_10972);
or U12399 (N_12399,N_10482,N_11556);
xor U12400 (N_12400,N_10971,N_10039);
xnor U12401 (N_12401,N_11880,N_10087);
nor U12402 (N_12402,N_10795,N_11160);
and U12403 (N_12403,N_11735,N_11162);
nor U12404 (N_12404,N_10326,N_10164);
and U12405 (N_12405,N_11156,N_11411);
or U12406 (N_12406,N_11549,N_11459);
and U12407 (N_12407,N_11496,N_10623);
nor U12408 (N_12408,N_10491,N_10176);
nor U12409 (N_12409,N_10104,N_11380);
and U12410 (N_12410,N_10201,N_10752);
nand U12411 (N_12411,N_11299,N_11154);
or U12412 (N_12412,N_11134,N_10256);
or U12413 (N_12413,N_10933,N_11351);
xnor U12414 (N_12414,N_10967,N_11465);
or U12415 (N_12415,N_10678,N_10306);
nor U12416 (N_12416,N_11602,N_11426);
or U12417 (N_12417,N_10489,N_11038);
or U12418 (N_12418,N_10652,N_10594);
nand U12419 (N_12419,N_11830,N_11615);
or U12420 (N_12420,N_11571,N_11483);
or U12421 (N_12421,N_11656,N_10808);
or U12422 (N_12422,N_11900,N_10814);
nand U12423 (N_12423,N_11668,N_10851);
nand U12424 (N_12424,N_11436,N_10082);
and U12425 (N_12425,N_11608,N_11078);
or U12426 (N_12426,N_10089,N_11488);
xor U12427 (N_12427,N_11976,N_10418);
nor U12428 (N_12428,N_11362,N_11437);
and U12429 (N_12429,N_10606,N_11593);
nand U12430 (N_12430,N_10637,N_10810);
nor U12431 (N_12431,N_10403,N_10137);
and U12432 (N_12432,N_11616,N_10170);
or U12433 (N_12433,N_11845,N_11015);
nor U12434 (N_12434,N_11688,N_10270);
nand U12435 (N_12435,N_10941,N_11310);
or U12436 (N_12436,N_10691,N_10805);
xnor U12437 (N_12437,N_11944,N_10151);
or U12438 (N_12438,N_11734,N_10347);
nand U12439 (N_12439,N_10727,N_10918);
nor U12440 (N_12440,N_10961,N_10633);
nand U12441 (N_12441,N_10346,N_10733);
nor U12442 (N_12442,N_10629,N_11048);
and U12443 (N_12443,N_10824,N_11533);
or U12444 (N_12444,N_10134,N_11050);
or U12445 (N_12445,N_11060,N_10663);
xor U12446 (N_12446,N_11864,N_11989);
or U12447 (N_12447,N_11245,N_11505);
xnor U12448 (N_12448,N_11221,N_11082);
and U12449 (N_12449,N_10599,N_10036);
or U12450 (N_12450,N_10829,N_10038);
nand U12451 (N_12451,N_11605,N_10909);
nand U12452 (N_12452,N_10917,N_11405);
nor U12453 (N_12453,N_10025,N_10697);
nand U12454 (N_12454,N_11125,N_10779);
or U12455 (N_12455,N_11010,N_10987);
nor U12456 (N_12456,N_11988,N_10687);
nand U12457 (N_12457,N_11140,N_11725);
or U12458 (N_12458,N_10597,N_11442);
nand U12459 (N_12459,N_10589,N_10675);
or U12460 (N_12460,N_11576,N_10426);
or U12461 (N_12461,N_10931,N_11143);
or U12462 (N_12462,N_10939,N_11798);
nand U12463 (N_12463,N_10031,N_11808);
or U12464 (N_12464,N_10008,N_11298);
nor U12465 (N_12465,N_11210,N_10579);
nor U12466 (N_12466,N_10837,N_10073);
and U12467 (N_12467,N_10107,N_11423);
xnor U12468 (N_12468,N_11567,N_11170);
and U12469 (N_12469,N_11449,N_10249);
nand U12470 (N_12470,N_10166,N_11416);
or U12471 (N_12471,N_11051,N_10093);
or U12472 (N_12472,N_11998,N_10806);
or U12473 (N_12473,N_10303,N_11786);
or U12474 (N_12474,N_10051,N_11563);
or U12475 (N_12475,N_10545,N_11804);
or U12476 (N_12476,N_11858,N_10088);
xor U12477 (N_12477,N_11025,N_11979);
xnor U12478 (N_12478,N_11915,N_10749);
or U12479 (N_12479,N_10265,N_10653);
nand U12480 (N_12480,N_10035,N_10181);
or U12481 (N_12481,N_11418,N_10676);
nor U12482 (N_12482,N_11841,N_11279);
or U12483 (N_12483,N_10617,N_11291);
or U12484 (N_12484,N_10739,N_11063);
and U12485 (N_12485,N_10938,N_11149);
nand U12486 (N_12486,N_10607,N_11183);
or U12487 (N_12487,N_11676,N_10227);
and U12488 (N_12488,N_10626,N_10778);
and U12489 (N_12489,N_10287,N_10743);
nor U12490 (N_12490,N_11895,N_11129);
or U12491 (N_12491,N_10513,N_11839);
xnor U12492 (N_12492,N_10511,N_10267);
or U12493 (N_12493,N_10009,N_11287);
nand U12494 (N_12494,N_11202,N_10849);
or U12495 (N_12495,N_10156,N_11644);
nand U12496 (N_12496,N_10294,N_11813);
and U12497 (N_12497,N_11448,N_10532);
nor U12498 (N_12498,N_10977,N_11516);
nand U12499 (N_12499,N_10846,N_10563);
nand U12500 (N_12500,N_10907,N_11535);
nand U12501 (N_12501,N_10420,N_11027);
nand U12502 (N_12502,N_11788,N_11995);
and U12503 (N_12503,N_11089,N_10714);
and U12504 (N_12504,N_10929,N_10530);
xnor U12505 (N_12505,N_10455,N_11100);
or U12506 (N_12506,N_10293,N_11165);
nand U12507 (N_12507,N_11878,N_10394);
nor U12508 (N_12508,N_11080,N_11000);
or U12509 (N_12509,N_10958,N_11551);
or U12510 (N_12510,N_11591,N_10718);
nor U12511 (N_12511,N_10005,N_11486);
or U12512 (N_12512,N_11945,N_11582);
nand U12513 (N_12513,N_10193,N_11091);
nand U12514 (N_12514,N_10756,N_10774);
nor U12515 (N_12515,N_10299,N_11696);
or U12516 (N_12516,N_11225,N_11952);
nor U12517 (N_12517,N_10924,N_10321);
nand U12518 (N_12518,N_10908,N_11790);
and U12519 (N_12519,N_10624,N_10439);
nand U12520 (N_12520,N_10462,N_10139);
and U12521 (N_12521,N_11200,N_11105);
xor U12522 (N_12522,N_11548,N_11550);
xor U12523 (N_12523,N_11792,N_10627);
nand U12524 (N_12524,N_10310,N_10129);
or U12525 (N_12525,N_10334,N_11875);
nand U12526 (N_12526,N_11597,N_11340);
or U12527 (N_12527,N_11250,N_11453);
nand U12528 (N_12528,N_11742,N_10565);
nor U12529 (N_12529,N_10167,N_11789);
nor U12530 (N_12530,N_10886,N_10561);
or U12531 (N_12531,N_11698,N_11918);
nand U12532 (N_12532,N_11963,N_10664);
nand U12533 (N_12533,N_10738,N_11775);
nor U12534 (N_12534,N_11113,N_10980);
xor U12535 (N_12535,N_11741,N_11726);
nor U12536 (N_12536,N_10584,N_11182);
and U12537 (N_12537,N_11949,N_10410);
or U12538 (N_12538,N_11810,N_10575);
or U12539 (N_12539,N_10437,N_10475);
and U12540 (N_12540,N_10979,N_11444);
or U12541 (N_12541,N_10710,N_10349);
or U12542 (N_12542,N_11622,N_11930);
nor U12543 (N_12543,N_10225,N_10240);
or U12544 (N_12544,N_11624,N_11552);
xor U12545 (N_12545,N_11058,N_10484);
or U12546 (N_12546,N_11541,N_10344);
and U12547 (N_12547,N_11914,N_10940);
nor U12548 (N_12548,N_11321,N_10271);
nor U12549 (N_12549,N_10495,N_11269);
or U12550 (N_12550,N_10079,N_11181);
xor U12551 (N_12551,N_10543,N_10698);
nor U12552 (N_12552,N_11278,N_10833);
and U12553 (N_12553,N_10921,N_11330);
nand U12554 (N_12554,N_10871,N_10797);
or U12555 (N_12555,N_10383,N_10557);
nor U12556 (N_12556,N_11365,N_11275);
or U12557 (N_12557,N_11638,N_10902);
xnor U12558 (N_12558,N_10136,N_11476);
and U12559 (N_12559,N_11704,N_11697);
and U12560 (N_12560,N_10884,N_10552);
or U12561 (N_12561,N_10242,N_10591);
nor U12562 (N_12562,N_11587,N_10246);
nand U12563 (N_12563,N_10496,N_10614);
or U12564 (N_12564,N_10056,N_11388);
nand U12565 (N_12565,N_11107,N_11539);
or U12566 (N_12566,N_10412,N_11594);
or U12567 (N_12567,N_10248,N_11122);
and U12568 (N_12568,N_10761,N_10538);
or U12569 (N_12569,N_10391,N_10040);
nor U12570 (N_12570,N_10188,N_10671);
xnor U12571 (N_12571,N_10114,N_10211);
nand U12572 (N_12572,N_11236,N_10202);
nand U12573 (N_12573,N_11738,N_11131);
nor U12574 (N_12574,N_11577,N_11244);
or U12575 (N_12575,N_11542,N_11214);
nand U12576 (N_12576,N_11955,N_10017);
or U12577 (N_12577,N_11821,N_10453);
and U12578 (N_12578,N_11977,N_11497);
or U12579 (N_12579,N_11184,N_10054);
nor U12580 (N_12580,N_10179,N_10052);
nand U12581 (N_12581,N_11825,N_10443);
xnor U12582 (N_12582,N_10919,N_10592);
nor U12583 (N_12583,N_10251,N_11208);
or U12584 (N_12584,N_10377,N_11385);
nand U12585 (N_12585,N_11161,N_10309);
nand U12586 (N_12586,N_11294,N_11138);
and U12587 (N_12587,N_10520,N_10551);
nor U12588 (N_12588,N_10068,N_10948);
nor U12589 (N_12589,N_11509,N_10677);
nor U12590 (N_12590,N_11191,N_11226);
nand U12591 (N_12591,N_11039,N_11033);
or U12592 (N_12592,N_11581,N_11935);
nand U12593 (N_12593,N_10126,N_10645);
nor U12594 (N_12594,N_11846,N_11522);
nand U12595 (N_12595,N_11425,N_10990);
nand U12596 (N_12596,N_10413,N_10830);
and U12597 (N_12597,N_11897,N_10745);
nor U12598 (N_12598,N_10244,N_11366);
or U12599 (N_12599,N_11247,N_10125);
and U12600 (N_12600,N_11827,N_11018);
and U12601 (N_12601,N_10717,N_10936);
and U12602 (N_12602,N_10096,N_11396);
or U12603 (N_12603,N_11300,N_10529);
nor U12604 (N_12604,N_11993,N_11720);
and U12605 (N_12605,N_10957,N_11911);
and U12606 (N_12606,N_11617,N_11375);
and U12607 (N_12607,N_11133,N_11504);
or U12608 (N_12608,N_11393,N_11954);
nand U12609 (N_12609,N_11889,N_11419);
or U12610 (N_12610,N_10277,N_11016);
and U12611 (N_12611,N_10944,N_11337);
or U12612 (N_12612,N_10390,N_11690);
nor U12613 (N_12613,N_11654,N_10371);
nor U12614 (N_12614,N_11061,N_11042);
nand U12615 (N_12615,N_11222,N_11047);
nor U12616 (N_12616,N_10514,N_10866);
or U12617 (N_12617,N_10904,N_10463);
xor U12618 (N_12618,N_10945,N_11755);
and U12619 (N_12619,N_10424,N_11088);
or U12620 (N_12620,N_10910,N_11613);
nand U12621 (N_12621,N_10893,N_10525);
and U12622 (N_12622,N_11716,N_10646);
or U12623 (N_12623,N_10081,N_11109);
and U12624 (N_12624,N_10583,N_11620);
or U12625 (N_12625,N_10206,N_11677);
nor U12626 (N_12626,N_11580,N_10831);
nor U12627 (N_12627,N_10001,N_11684);
or U12628 (N_12628,N_11691,N_10506);
and U12629 (N_12629,N_10059,N_10631);
nand U12630 (N_12630,N_11360,N_10536);
or U12631 (N_12631,N_11148,N_11802);
xnor U12632 (N_12632,N_11009,N_10527);
nor U12633 (N_12633,N_10515,N_11401);
nand U12634 (N_12634,N_10705,N_10747);
or U12635 (N_12635,N_10045,N_11403);
or U12636 (N_12636,N_10723,N_11817);
xnor U12637 (N_12637,N_11633,N_10386);
or U12638 (N_12638,N_11023,N_11189);
xor U12639 (N_12639,N_10140,N_10389);
nand U12640 (N_12640,N_11410,N_11054);
or U12641 (N_12641,N_11460,N_10169);
nor U12642 (N_12642,N_11209,N_10069);
or U12643 (N_12643,N_10161,N_11859);
and U12644 (N_12644,N_10636,N_10661);
nor U12645 (N_12645,N_11980,N_10103);
or U12646 (N_12646,N_10376,N_10858);
xor U12647 (N_12647,N_11288,N_10955);
xnor U12648 (N_12648,N_10345,N_10966);
or U12649 (N_12649,N_10823,N_10241);
xnor U12650 (N_12650,N_10615,N_11872);
or U12651 (N_12651,N_10571,N_10304);
nand U12652 (N_12652,N_10757,N_11293);
nand U12653 (N_12653,N_11102,N_10873);
nand U12654 (N_12654,N_10419,N_11338);
and U12655 (N_12655,N_11767,N_10892);
nor U12656 (N_12656,N_11097,N_11467);
nor U12657 (N_12657,N_10923,N_10540);
or U12658 (N_12658,N_10807,N_10812);
or U12659 (N_12659,N_11185,N_10876);
or U12660 (N_12660,N_11232,N_11984);
nand U12661 (N_12661,N_11521,N_10111);
or U12662 (N_12662,N_11252,N_10930);
xnor U12663 (N_12663,N_10100,N_10622);
and U12664 (N_12664,N_11883,N_10396);
nor U12665 (N_12665,N_10226,N_10243);
nand U12666 (N_12666,N_10220,N_10605);
nor U12667 (N_12667,N_10123,N_10407);
nor U12668 (N_12668,N_10862,N_11070);
and U12669 (N_12669,N_11095,N_11325);
nand U12670 (N_12670,N_11227,N_11121);
and U12671 (N_12671,N_11257,N_11475);
and U12672 (N_12672,N_11559,N_10517);
nor U12673 (N_12673,N_10238,N_10724);
or U12674 (N_12674,N_11440,N_10995);
nand U12675 (N_12675,N_11842,N_11387);
xor U12676 (N_12676,N_10116,N_11867);
nor U12677 (N_12677,N_11612,N_10350);
and U12678 (N_12678,N_11787,N_11141);
nand U12679 (N_12679,N_10781,N_10531);
or U12680 (N_12680,N_10106,N_11991);
and U12681 (N_12681,N_10879,N_10499);
and U12682 (N_12682,N_11765,N_11972);
nor U12683 (N_12683,N_11068,N_10192);
or U12684 (N_12684,N_10553,N_11693);
nand U12685 (N_12685,N_11499,N_10194);
or U12686 (N_12686,N_10133,N_11814);
or U12687 (N_12687,N_10356,N_11029);
or U12688 (N_12688,N_11053,N_10190);
nor U12689 (N_12689,N_10408,N_11868);
and U12690 (N_12690,N_10431,N_10993);
nand U12691 (N_12691,N_10360,N_10728);
and U12692 (N_12692,N_10010,N_11713);
or U12693 (N_12693,N_11126,N_10094);
xnor U12694 (N_12694,N_11923,N_10504);
and U12695 (N_12695,N_10682,N_11985);
nor U12696 (N_12696,N_11635,N_11090);
and U12697 (N_12697,N_10868,N_11515);
nor U12698 (N_12698,N_11292,N_10994);
and U12699 (N_12699,N_11714,N_11424);
nor U12700 (N_12700,N_10746,N_11590);
and U12701 (N_12701,N_11034,N_11978);
or U12702 (N_12702,N_11763,N_10975);
nand U12703 (N_12703,N_11341,N_10331);
and U12704 (N_12704,N_10162,N_10951);
nor U12705 (N_12705,N_10973,N_11168);
xnor U12706 (N_12706,N_10297,N_10555);
and U12707 (N_12707,N_10015,N_11164);
nand U12708 (N_12708,N_11778,N_11274);
xor U12709 (N_12709,N_11639,N_11557);
and U12710 (N_12710,N_10554,N_10163);
nor U12711 (N_12711,N_10683,N_11007);
and U12712 (N_12712,N_10736,N_11745);
and U12713 (N_12713,N_11494,N_11619);
nor U12714 (N_12714,N_11715,N_11573);
nand U12715 (N_12715,N_11701,N_11137);
nand U12716 (N_12716,N_10120,N_11871);
nand U12717 (N_12717,N_11604,N_10237);
and U12718 (N_12718,N_10388,N_10947);
xnor U12719 (N_12719,N_11024,N_11256);
or U12720 (N_12720,N_10452,N_11819);
or U12721 (N_12721,N_10839,N_11513);
nor U12722 (N_12722,N_11389,N_10730);
nor U12723 (N_12723,N_11217,N_11925);
xnor U12724 (N_12724,N_11748,N_10772);
nand U12725 (N_12725,N_11498,N_11653);
and U12726 (N_12726,N_10318,N_10357);
nor U12727 (N_12727,N_10438,N_10065);
nor U12728 (N_12728,N_11877,N_11934);
nor U12729 (N_12729,N_10911,N_10679);
or U12730 (N_12730,N_11461,N_11355);
and U12731 (N_12731,N_10735,N_10703);
nand U12732 (N_12732,N_11072,N_11342);
and U12733 (N_12733,N_11395,N_11611);
xor U12734 (N_12734,N_10014,N_10062);
nor U12735 (N_12735,N_11882,N_10336);
nor U12736 (N_12736,N_10510,N_10030);
and U12737 (N_12737,N_10135,N_11230);
nor U12738 (N_12738,N_11071,N_10209);
or U12739 (N_12739,N_10783,N_10066);
nand U12740 (N_12740,N_10609,N_11114);
and U12741 (N_12741,N_10189,N_11201);
xor U12742 (N_12742,N_11253,N_10821);
and U12743 (N_12743,N_11546,N_10965);
or U12744 (N_12744,N_11771,N_11124);
xor U12745 (N_12745,N_10621,N_10699);
nor U12746 (N_12746,N_11532,N_11171);
or U12747 (N_12747,N_11592,N_11574);
nand U12748 (N_12748,N_11328,N_10523);
nand U12749 (N_12749,N_10854,N_11323);
or U12750 (N_12750,N_10668,N_10187);
nand U12751 (N_12751,N_11937,N_10061);
and U12752 (N_12752,N_11435,N_10835);
or U12753 (N_12753,N_10342,N_10435);
nor U12754 (N_12754,N_11240,N_10026);
nand U12755 (N_12755,N_11627,N_10469);
and U12756 (N_12756,N_10765,N_11032);
and U12757 (N_12757,N_10741,N_11011);
or U12758 (N_12758,N_10422,N_10869);
xor U12759 (N_12759,N_10467,N_11876);
or U12760 (N_12760,N_11119,N_10000);
and U12761 (N_12761,N_11087,N_10533);
xor U12762 (N_12762,N_10016,N_11596);
and U12763 (N_12763,N_11260,N_10852);
or U12764 (N_12764,N_11973,N_11518);
nand U12765 (N_12765,N_10777,N_10695);
nor U12766 (N_12766,N_10832,N_11850);
xnor U12767 (N_12767,N_11420,N_11022);
nand U12768 (N_12768,N_10729,N_10002);
nor U12769 (N_12769,N_11381,N_11508);
nor U12770 (N_12770,N_11481,N_10128);
nor U12771 (N_12771,N_10028,N_10573);
or U12772 (N_12772,N_11694,N_11429);
and U12773 (N_12773,N_11928,N_10480);
nor U12774 (N_12774,N_10034,N_11723);
or U12775 (N_12775,N_11469,N_11777);
nor U12776 (N_12776,N_11673,N_11951);
or U12777 (N_12777,N_11905,N_11645);
nand U12778 (N_12778,N_10044,N_10050);
and U12779 (N_12779,N_10593,N_11926);
and U12780 (N_12780,N_11886,N_10255);
nor U12781 (N_12781,N_10521,N_10483);
nand U12782 (N_12782,N_11086,N_10560);
and U12783 (N_12783,N_10235,N_10612);
xnor U12784 (N_12784,N_10580,N_11543);
nor U12785 (N_12785,N_10458,N_10659);
and U12786 (N_12786,N_10118,N_11103);
and U12787 (N_12787,N_10711,N_10070);
or U12788 (N_12788,N_11178,N_10157);
xor U12789 (N_12789,N_11412,N_10312);
nand U12790 (N_12790,N_10132,N_10899);
and U12791 (N_12791,N_11272,N_11664);
nand U12792 (N_12792,N_10731,N_10569);
nor U12793 (N_12793,N_10440,N_11678);
and U12794 (N_12794,N_11135,N_11358);
nor U12795 (N_12795,N_10022,N_11357);
and U12796 (N_12796,N_11001,N_10481);
nand U12797 (N_12797,N_11796,N_11005);
nand U12798 (N_12798,N_10744,N_11832);
nand U12799 (N_12799,N_10353,N_10319);
nor U12800 (N_12800,N_11520,N_11347);
nor U12801 (N_12801,N_10566,N_10651);
and U12802 (N_12802,N_11575,N_11118);
and U12803 (N_12803,N_11139,N_11207);
nor U12804 (N_12804,N_11485,N_10996);
and U12805 (N_12805,N_11314,N_11261);
and U12806 (N_12806,N_10544,N_10416);
and U12807 (N_12807,N_10395,N_10232);
or U12808 (N_12808,N_10577,N_11997);
or U12809 (N_12809,N_11640,N_10794);
nand U12810 (N_12810,N_11851,N_10872);
nor U12811 (N_12811,N_11450,N_10628);
nor U12812 (N_12812,N_10713,N_10337);
nand U12813 (N_12813,N_11144,N_11866);
nand U12814 (N_12814,N_11263,N_11373);
and U12815 (N_12815,N_11409,N_11890);
nand U12816 (N_12816,N_11606,N_11422);
nand U12817 (N_12817,N_10351,N_11319);
or U12818 (N_12818,N_11370,N_11377);
nor U12819 (N_12819,N_10447,N_11884);
and U12820 (N_12820,N_11285,N_10604);
nor U12821 (N_12821,N_11840,N_11800);
and U12822 (N_12822,N_11372,N_10508);
xnor U12823 (N_12823,N_10444,N_11938);
and U12824 (N_12824,N_10278,N_10374);
or U12825 (N_12825,N_11695,N_11835);
nor U12826 (N_12826,N_10535,N_11281);
and U12827 (N_12827,N_10632,N_10316);
or U12828 (N_12828,N_11940,N_11163);
nor U12829 (N_12829,N_11857,N_11632);
or U12830 (N_12830,N_11909,N_11658);
or U12831 (N_12831,N_11056,N_10358);
or U12832 (N_12832,N_10720,N_11641);
nand U12833 (N_12833,N_11199,N_11948);
and U12834 (N_12834,N_11439,N_10195);
and U12835 (N_12835,N_11331,N_11910);
and U12836 (N_12836,N_11970,N_11382);
nor U12837 (N_12837,N_11128,N_11595);
xor U12838 (N_12838,N_11487,N_10382);
or U12839 (N_12839,N_10949,N_11634);
and U12840 (N_12840,N_10999,N_10124);
xnor U12841 (N_12841,N_11266,N_11233);
nand U12842 (N_12842,N_10033,N_10619);
or U12843 (N_12843,N_11151,N_10890);
and U12844 (N_12844,N_11899,N_11950);
and U12845 (N_12845,N_11271,N_10401);
and U12846 (N_12846,N_10634,N_10274);
or U12847 (N_12847,N_11268,N_10099);
nor U12848 (N_12848,N_11399,N_10608);
and U12849 (N_12849,N_10834,N_11036);
nand U12850 (N_12850,N_11251,N_11903);
xor U12851 (N_12851,N_11434,N_10468);
nor U12852 (N_12852,N_11049,N_11647);
or U12853 (N_12853,N_10867,N_11986);
and U12854 (N_12854,N_10771,N_11457);
nor U12855 (N_12855,N_10127,N_10320);
nor U12856 (N_12856,N_10315,N_10023);
nor U12857 (N_12857,N_11511,N_10282);
xnor U12858 (N_12858,N_11600,N_11308);
nor U12859 (N_12859,N_11657,N_10064);
nand U12860 (N_12860,N_11672,N_11703);
or U12861 (N_12861,N_10086,N_11130);
and U12862 (N_12862,N_11480,N_11326);
or U12863 (N_12863,N_11902,N_10512);
xnor U12864 (N_12864,N_10470,N_11683);
or U12865 (N_12865,N_10643,N_10417);
xnor U12866 (N_12866,N_11531,N_11759);
nand U12867 (N_12867,N_11724,N_10574);
xor U12868 (N_12868,N_11320,N_10516);
nor U12869 (N_12869,N_10172,N_11585);
nor U12870 (N_12870,N_10865,N_11462);
xor U12871 (N_12871,N_11781,N_11967);
nor U12872 (N_12872,N_11307,N_10817);
xnor U12873 (N_12873,N_10798,N_10105);
and U12874 (N_12874,N_11700,N_11650);
xnor U12875 (N_12875,N_11921,N_11075);
nand U12876 (N_12876,N_11999,N_11008);
nand U12877 (N_12877,N_10174,N_10233);
nor U12878 (N_12878,N_11013,N_11711);
or U12879 (N_12879,N_11626,N_10505);
xor U12880 (N_12880,N_10953,N_11891);
nand U12881 (N_12881,N_11610,N_10725);
nor U12882 (N_12882,N_11743,N_11205);
and U12883 (N_12883,N_11194,N_10084);
or U12884 (N_12884,N_11379,N_11826);
and U12885 (N_12885,N_10122,N_10742);
xor U12886 (N_12886,N_11680,N_10180);
nor U12887 (N_12887,N_11863,N_11718);
and U12888 (N_12888,N_10130,N_11667);
nor U12889 (N_12889,N_10370,N_10649);
nor U12890 (N_12890,N_11099,N_11731);
or U12891 (N_12891,N_10707,N_10935);
nor U12892 (N_12892,N_11537,N_10964);
nand U12893 (N_12893,N_11237,N_11280);
nor U12894 (N_12894,N_11329,N_10145);
and U12895 (N_12895,N_11374,N_10524);
nand U12896 (N_12896,N_11098,N_11017);
nor U12897 (N_12897,N_10518,N_10158);
nand U12898 (N_12898,N_10448,N_10528);
nor U12899 (N_12899,N_10364,N_11555);
and U12900 (N_12900,N_11968,N_11558);
and U12901 (N_12901,N_10258,N_10790);
and U12902 (N_12902,N_11220,N_10689);
and U12903 (N_12903,N_10509,N_10792);
or U12904 (N_12904,N_10501,N_11472);
nor U12905 (N_12905,N_11187,N_10712);
and U12906 (N_12906,N_10298,N_11190);
or U12907 (N_12907,N_10507,N_11076);
xnor U12908 (N_12908,N_11402,N_11663);
nand U12909 (N_12909,N_10943,N_11041);
and U12910 (N_12910,N_11383,N_11093);
nor U12911 (N_12911,N_11136,N_11265);
and U12912 (N_12912,N_10177,N_10219);
nand U12913 (N_12913,N_10602,N_11727);
nand U12914 (N_12914,N_11044,N_11795);
or U12915 (N_12915,N_10178,N_10978);
nor U12916 (N_12916,N_11506,N_10588);
or U12917 (N_12917,N_11893,N_10198);
and U12918 (N_12918,N_10847,N_11470);
and U12919 (N_12919,N_10428,N_11348);
nor U12920 (N_12920,N_11599,N_10828);
or U12921 (N_12921,N_10155,N_10168);
and U12922 (N_12922,N_10701,N_11947);
nor U12923 (N_12923,N_11492,N_10091);
and U12924 (N_12924,N_10191,N_11959);
nand U12925 (N_12925,N_11666,N_11512);
or U12926 (N_12926,N_10074,N_11737);
nor U12927 (N_12927,N_10891,N_10329);
xnor U12928 (N_12928,N_11524,N_11282);
and U12929 (N_12929,N_10819,N_11343);
nor U12930 (N_12930,N_10878,N_10330);
nand U12931 (N_12931,N_10092,N_10300);
nand U12932 (N_12932,N_11002,N_11132);
and U12933 (N_12933,N_10603,N_11621);
nor U12934 (N_12934,N_10804,N_10827);
nor U12935 (N_12935,N_10925,N_11933);
nand U12936 (N_12936,N_11474,N_11816);
or U12937 (N_12937,N_11865,N_11519);
nand U12938 (N_12938,N_11589,N_10212);
or U12939 (N_12939,N_11828,N_11823);
nor U12940 (N_12940,N_10669,N_11643);
nand U12941 (N_12941,N_11203,N_10681);
or U12942 (N_12942,N_11452,N_10916);
and U12943 (N_12943,N_11770,N_11262);
nor U12944 (N_12944,N_11195,N_10213);
or U12945 (N_12945,N_11879,N_10567);
nand U12946 (N_12946,N_10473,N_10414);
or U12947 (N_12947,N_11956,N_10338);
nor U12948 (N_12948,N_10630,N_10368);
or U12949 (N_12949,N_10898,N_11560);
xor U12950 (N_12950,N_10970,N_10097);
nor U12951 (N_12951,N_11547,N_11894);
and U12952 (N_12952,N_10737,N_11350);
or U12953 (N_12953,N_11173,N_10029);
nand U12954 (N_12954,N_11204,N_11885);
nand U12955 (N_12955,N_10153,N_11776);
and U12956 (N_12956,N_11142,N_11568);
nor U12957 (N_12957,N_11803,N_11206);
or U12958 (N_12958,N_10618,N_10992);
xnor U12959 (N_12959,N_11689,N_11773);
xor U12960 (N_12960,N_10142,N_10327);
and U12961 (N_12961,N_10141,N_10119);
and U12962 (N_12962,N_11390,N_10954);
and U12963 (N_12963,N_10905,N_11246);
and U12964 (N_12964,N_10339,N_11211);
xnor U12965 (N_12965,N_11283,N_11479);
nand U12966 (N_12966,N_10903,N_11116);
nor U12967 (N_12967,N_10982,N_11904);
nor U12968 (N_12968,N_10497,N_11917);
and U12969 (N_12969,N_11336,N_11526);
and U12970 (N_12970,N_11092,N_11794);
nor U12971 (N_12971,N_10205,N_10875);
and U12972 (N_12972,N_11427,N_10301);
nor U12973 (N_12973,N_10406,N_11346);
or U12974 (N_12974,N_10102,N_11687);
nand U12975 (N_12975,N_10568,N_10397);
or U12976 (N_12976,N_11249,N_11368);
nand U12977 (N_12977,N_10549,N_11774);
nor U12978 (N_12978,N_10547,N_10398);
xnor U12979 (N_12979,N_10673,N_11772);
xnor U12980 (N_12980,N_11407,N_10425);
and U12981 (N_12981,N_11807,N_11037);
or U12982 (N_12982,N_11297,N_10340);
and U12983 (N_12983,N_10113,N_11500);
nand U12984 (N_12984,N_10186,N_11983);
nand U12985 (N_12985,N_11394,N_10857);
and U12986 (N_12986,N_10148,N_11215);
and U12987 (N_12987,N_10877,N_11074);
or U12988 (N_12988,N_11762,N_10755);
nor U12989 (N_12989,N_10264,N_10067);
and U12990 (N_12990,N_11417,N_10048);
nand U12991 (N_12991,N_11284,N_11964);
nor U12992 (N_12992,N_10657,N_10883);
and U12993 (N_12993,N_11756,N_11818);
or U12994 (N_12994,N_11769,N_11363);
nor U12995 (N_12995,N_10952,N_10399);
or U12996 (N_12996,N_10598,N_10027);
nor U12997 (N_12997,N_10750,N_10363);
or U12998 (N_12998,N_11953,N_11258);
nand U12999 (N_12999,N_11746,N_10786);
xor U13000 (N_13000,N_11573,N_10569);
nor U13001 (N_13001,N_11856,N_10571);
nand U13002 (N_13002,N_10876,N_10415);
or U13003 (N_13003,N_11068,N_11217);
or U13004 (N_13004,N_10745,N_11344);
or U13005 (N_13005,N_11917,N_11934);
nor U13006 (N_13006,N_10887,N_11762);
nor U13007 (N_13007,N_11894,N_11035);
nand U13008 (N_13008,N_11233,N_11799);
or U13009 (N_13009,N_10136,N_10128);
and U13010 (N_13010,N_10885,N_11948);
or U13011 (N_13011,N_10191,N_10738);
and U13012 (N_13012,N_10895,N_11798);
nor U13013 (N_13013,N_11750,N_11093);
or U13014 (N_13014,N_11882,N_10130);
or U13015 (N_13015,N_10202,N_10396);
nand U13016 (N_13016,N_10886,N_10443);
nor U13017 (N_13017,N_11069,N_10977);
or U13018 (N_13018,N_10849,N_11145);
nand U13019 (N_13019,N_11360,N_11744);
and U13020 (N_13020,N_11328,N_10630);
nand U13021 (N_13021,N_10793,N_10818);
xnor U13022 (N_13022,N_10903,N_11013);
nand U13023 (N_13023,N_11172,N_10666);
and U13024 (N_13024,N_11415,N_11718);
nor U13025 (N_13025,N_10941,N_10794);
or U13026 (N_13026,N_11493,N_10870);
nand U13027 (N_13027,N_10750,N_11088);
nand U13028 (N_13028,N_10827,N_10103);
nor U13029 (N_13029,N_11811,N_11461);
and U13030 (N_13030,N_11001,N_11223);
nor U13031 (N_13031,N_11051,N_10103);
xor U13032 (N_13032,N_10430,N_10065);
nand U13033 (N_13033,N_11701,N_10976);
or U13034 (N_13034,N_10582,N_10882);
and U13035 (N_13035,N_10144,N_10632);
nor U13036 (N_13036,N_11861,N_11877);
nor U13037 (N_13037,N_10612,N_10207);
nand U13038 (N_13038,N_11508,N_10642);
and U13039 (N_13039,N_11494,N_10390);
xnor U13040 (N_13040,N_10594,N_10855);
or U13041 (N_13041,N_10888,N_11548);
or U13042 (N_13042,N_11818,N_10141);
xor U13043 (N_13043,N_11986,N_11457);
nand U13044 (N_13044,N_10890,N_11558);
xor U13045 (N_13045,N_11145,N_11044);
or U13046 (N_13046,N_11152,N_11744);
nor U13047 (N_13047,N_10363,N_10580);
nor U13048 (N_13048,N_10733,N_11868);
nor U13049 (N_13049,N_11590,N_11050);
or U13050 (N_13050,N_11113,N_10359);
or U13051 (N_13051,N_11762,N_10842);
nand U13052 (N_13052,N_10181,N_11357);
nand U13053 (N_13053,N_11007,N_11440);
nor U13054 (N_13054,N_10164,N_10586);
nor U13055 (N_13055,N_11497,N_11527);
nand U13056 (N_13056,N_10680,N_10070);
and U13057 (N_13057,N_10710,N_11236);
nor U13058 (N_13058,N_11313,N_10789);
nand U13059 (N_13059,N_11872,N_11414);
nand U13060 (N_13060,N_11708,N_10097);
nor U13061 (N_13061,N_10403,N_11339);
nand U13062 (N_13062,N_11678,N_11264);
or U13063 (N_13063,N_11324,N_10377);
and U13064 (N_13064,N_11266,N_11026);
nor U13065 (N_13065,N_10482,N_11972);
and U13066 (N_13066,N_10736,N_11802);
and U13067 (N_13067,N_11539,N_11692);
and U13068 (N_13068,N_11454,N_10533);
nor U13069 (N_13069,N_11726,N_11026);
nor U13070 (N_13070,N_10934,N_11119);
nor U13071 (N_13071,N_11947,N_10313);
and U13072 (N_13072,N_11547,N_10024);
nor U13073 (N_13073,N_10077,N_10948);
xnor U13074 (N_13074,N_11724,N_10514);
nor U13075 (N_13075,N_11600,N_11984);
or U13076 (N_13076,N_10718,N_11894);
and U13077 (N_13077,N_10873,N_11504);
xor U13078 (N_13078,N_10115,N_11253);
and U13079 (N_13079,N_11814,N_11362);
and U13080 (N_13080,N_11593,N_10033);
or U13081 (N_13081,N_11586,N_10135);
nand U13082 (N_13082,N_11080,N_11638);
nor U13083 (N_13083,N_11880,N_10668);
nor U13084 (N_13084,N_11756,N_10647);
nand U13085 (N_13085,N_11208,N_10781);
xnor U13086 (N_13086,N_10136,N_11347);
or U13087 (N_13087,N_10120,N_11236);
or U13088 (N_13088,N_11536,N_11502);
nand U13089 (N_13089,N_11803,N_11285);
or U13090 (N_13090,N_11784,N_10449);
nand U13091 (N_13091,N_11444,N_11116);
nor U13092 (N_13092,N_11306,N_10490);
and U13093 (N_13093,N_10280,N_10301);
nand U13094 (N_13094,N_11300,N_10770);
and U13095 (N_13095,N_10095,N_10209);
nor U13096 (N_13096,N_10422,N_10064);
or U13097 (N_13097,N_11761,N_11121);
and U13098 (N_13098,N_10685,N_10560);
and U13099 (N_13099,N_10766,N_11910);
nor U13100 (N_13100,N_11801,N_10557);
or U13101 (N_13101,N_11865,N_10580);
and U13102 (N_13102,N_10089,N_10783);
nand U13103 (N_13103,N_10662,N_10176);
nor U13104 (N_13104,N_11291,N_10773);
xor U13105 (N_13105,N_10861,N_10712);
or U13106 (N_13106,N_10256,N_11850);
nor U13107 (N_13107,N_11442,N_11843);
or U13108 (N_13108,N_11823,N_11088);
and U13109 (N_13109,N_11518,N_11746);
and U13110 (N_13110,N_11641,N_11185);
or U13111 (N_13111,N_11932,N_11618);
nand U13112 (N_13112,N_10106,N_11053);
and U13113 (N_13113,N_11788,N_11778);
nor U13114 (N_13114,N_11246,N_11074);
nand U13115 (N_13115,N_10334,N_10649);
nor U13116 (N_13116,N_10486,N_10649);
nor U13117 (N_13117,N_10798,N_11557);
and U13118 (N_13118,N_10411,N_10018);
nor U13119 (N_13119,N_11435,N_10723);
and U13120 (N_13120,N_10669,N_10556);
nor U13121 (N_13121,N_11526,N_10870);
and U13122 (N_13122,N_11602,N_10217);
nor U13123 (N_13123,N_10908,N_11518);
nor U13124 (N_13124,N_11230,N_10753);
or U13125 (N_13125,N_11120,N_11780);
nand U13126 (N_13126,N_10532,N_10398);
nand U13127 (N_13127,N_10749,N_10849);
nand U13128 (N_13128,N_10286,N_11364);
or U13129 (N_13129,N_11107,N_11693);
nand U13130 (N_13130,N_11022,N_11104);
nand U13131 (N_13131,N_11322,N_11225);
nand U13132 (N_13132,N_11496,N_10903);
or U13133 (N_13133,N_10406,N_11290);
or U13134 (N_13134,N_11271,N_10482);
nor U13135 (N_13135,N_10813,N_11667);
and U13136 (N_13136,N_10893,N_10829);
or U13137 (N_13137,N_10007,N_11104);
xnor U13138 (N_13138,N_11505,N_10294);
and U13139 (N_13139,N_11757,N_10204);
xor U13140 (N_13140,N_11393,N_11362);
nor U13141 (N_13141,N_11308,N_11548);
and U13142 (N_13142,N_11290,N_11114);
or U13143 (N_13143,N_11063,N_11659);
nand U13144 (N_13144,N_10928,N_11974);
xor U13145 (N_13145,N_10197,N_10086);
nand U13146 (N_13146,N_11892,N_11314);
nand U13147 (N_13147,N_11701,N_10202);
nor U13148 (N_13148,N_10541,N_11274);
and U13149 (N_13149,N_11056,N_10859);
or U13150 (N_13150,N_10140,N_10006);
and U13151 (N_13151,N_10505,N_11164);
and U13152 (N_13152,N_11050,N_10365);
nor U13153 (N_13153,N_10487,N_10982);
or U13154 (N_13154,N_10487,N_11622);
xnor U13155 (N_13155,N_11127,N_10878);
or U13156 (N_13156,N_10263,N_11785);
nand U13157 (N_13157,N_10599,N_11513);
and U13158 (N_13158,N_10667,N_10232);
nor U13159 (N_13159,N_10730,N_11477);
nor U13160 (N_13160,N_11424,N_11259);
nand U13161 (N_13161,N_11142,N_11543);
and U13162 (N_13162,N_11572,N_10360);
xor U13163 (N_13163,N_11487,N_10791);
or U13164 (N_13164,N_10495,N_10234);
nor U13165 (N_13165,N_11537,N_11410);
nor U13166 (N_13166,N_10870,N_10431);
nand U13167 (N_13167,N_10364,N_10764);
or U13168 (N_13168,N_11779,N_10154);
or U13169 (N_13169,N_10553,N_11193);
nand U13170 (N_13170,N_10159,N_10525);
nand U13171 (N_13171,N_11506,N_11107);
nand U13172 (N_13172,N_11884,N_10154);
and U13173 (N_13173,N_10727,N_10447);
xnor U13174 (N_13174,N_11698,N_10220);
or U13175 (N_13175,N_11116,N_10881);
and U13176 (N_13176,N_10416,N_10172);
or U13177 (N_13177,N_10453,N_11654);
or U13178 (N_13178,N_10084,N_10945);
nor U13179 (N_13179,N_11464,N_10464);
nor U13180 (N_13180,N_11766,N_10848);
or U13181 (N_13181,N_10323,N_10626);
or U13182 (N_13182,N_10602,N_10697);
or U13183 (N_13183,N_10445,N_11773);
nor U13184 (N_13184,N_10948,N_11110);
xnor U13185 (N_13185,N_10642,N_11084);
or U13186 (N_13186,N_10386,N_10663);
or U13187 (N_13187,N_10225,N_11291);
nor U13188 (N_13188,N_11172,N_11889);
and U13189 (N_13189,N_10974,N_11777);
nand U13190 (N_13190,N_10094,N_10167);
and U13191 (N_13191,N_10946,N_10042);
nor U13192 (N_13192,N_10349,N_10480);
and U13193 (N_13193,N_10276,N_11581);
nor U13194 (N_13194,N_11898,N_10447);
nand U13195 (N_13195,N_10283,N_10742);
or U13196 (N_13196,N_11711,N_11664);
and U13197 (N_13197,N_10028,N_11256);
or U13198 (N_13198,N_11636,N_11022);
or U13199 (N_13199,N_10498,N_10311);
nor U13200 (N_13200,N_10117,N_10170);
xnor U13201 (N_13201,N_11747,N_10287);
nor U13202 (N_13202,N_11741,N_10634);
or U13203 (N_13203,N_11130,N_10554);
nor U13204 (N_13204,N_10754,N_10410);
or U13205 (N_13205,N_10454,N_10687);
or U13206 (N_13206,N_11888,N_10073);
nor U13207 (N_13207,N_10943,N_11642);
and U13208 (N_13208,N_10123,N_11874);
nor U13209 (N_13209,N_11732,N_11096);
and U13210 (N_13210,N_11979,N_10852);
and U13211 (N_13211,N_10029,N_10368);
nand U13212 (N_13212,N_10491,N_10702);
xnor U13213 (N_13213,N_11632,N_10937);
nand U13214 (N_13214,N_11607,N_11365);
nand U13215 (N_13215,N_10618,N_11764);
nand U13216 (N_13216,N_11349,N_10417);
and U13217 (N_13217,N_11583,N_10776);
nor U13218 (N_13218,N_11971,N_11391);
or U13219 (N_13219,N_11712,N_10718);
nand U13220 (N_13220,N_11516,N_11803);
nand U13221 (N_13221,N_10752,N_10643);
or U13222 (N_13222,N_10354,N_10758);
nor U13223 (N_13223,N_11472,N_11097);
nor U13224 (N_13224,N_10980,N_11938);
nand U13225 (N_13225,N_10451,N_10580);
nand U13226 (N_13226,N_10000,N_11243);
nand U13227 (N_13227,N_10347,N_11998);
nor U13228 (N_13228,N_10383,N_10229);
nor U13229 (N_13229,N_10118,N_10970);
nand U13230 (N_13230,N_10987,N_10888);
and U13231 (N_13231,N_10078,N_11964);
nor U13232 (N_13232,N_10351,N_10551);
nand U13233 (N_13233,N_11893,N_10776);
nand U13234 (N_13234,N_11403,N_11484);
and U13235 (N_13235,N_11363,N_10185);
nor U13236 (N_13236,N_10079,N_10947);
or U13237 (N_13237,N_11516,N_11672);
or U13238 (N_13238,N_10524,N_10153);
nand U13239 (N_13239,N_11539,N_10362);
xnor U13240 (N_13240,N_11467,N_11706);
and U13241 (N_13241,N_10602,N_11289);
nor U13242 (N_13242,N_10444,N_11293);
nand U13243 (N_13243,N_11119,N_11352);
nand U13244 (N_13244,N_11617,N_11924);
or U13245 (N_13245,N_11542,N_11310);
xor U13246 (N_13246,N_10081,N_10578);
nand U13247 (N_13247,N_10670,N_11388);
xnor U13248 (N_13248,N_10740,N_10738);
nand U13249 (N_13249,N_11809,N_11623);
nand U13250 (N_13250,N_11280,N_11434);
nand U13251 (N_13251,N_11116,N_11152);
and U13252 (N_13252,N_10252,N_11586);
nor U13253 (N_13253,N_11309,N_11893);
nor U13254 (N_13254,N_10496,N_10904);
or U13255 (N_13255,N_11672,N_11137);
and U13256 (N_13256,N_11539,N_11468);
or U13257 (N_13257,N_10616,N_10558);
nand U13258 (N_13258,N_11088,N_11557);
nand U13259 (N_13259,N_10387,N_11399);
or U13260 (N_13260,N_11267,N_10751);
nand U13261 (N_13261,N_10725,N_11015);
and U13262 (N_13262,N_10580,N_10071);
nand U13263 (N_13263,N_10414,N_10026);
or U13264 (N_13264,N_10996,N_10744);
or U13265 (N_13265,N_11392,N_10094);
nand U13266 (N_13266,N_11906,N_10882);
xor U13267 (N_13267,N_10209,N_10316);
xnor U13268 (N_13268,N_10669,N_10331);
xor U13269 (N_13269,N_11243,N_11374);
nor U13270 (N_13270,N_11651,N_10512);
nor U13271 (N_13271,N_11521,N_10282);
and U13272 (N_13272,N_10222,N_10423);
or U13273 (N_13273,N_10337,N_11871);
or U13274 (N_13274,N_10502,N_10034);
or U13275 (N_13275,N_11592,N_11824);
xnor U13276 (N_13276,N_10534,N_11601);
and U13277 (N_13277,N_10682,N_11068);
and U13278 (N_13278,N_11986,N_10730);
xor U13279 (N_13279,N_11525,N_10609);
nand U13280 (N_13280,N_10633,N_11589);
nor U13281 (N_13281,N_11913,N_10551);
nor U13282 (N_13282,N_11273,N_10806);
nand U13283 (N_13283,N_11783,N_10938);
nand U13284 (N_13284,N_11197,N_11380);
nand U13285 (N_13285,N_11155,N_11813);
and U13286 (N_13286,N_10149,N_10808);
and U13287 (N_13287,N_11820,N_10568);
nand U13288 (N_13288,N_10883,N_11147);
nor U13289 (N_13289,N_11332,N_11397);
nand U13290 (N_13290,N_11759,N_10268);
nand U13291 (N_13291,N_11345,N_11091);
nand U13292 (N_13292,N_11440,N_11078);
nor U13293 (N_13293,N_11977,N_10143);
or U13294 (N_13294,N_11744,N_11707);
or U13295 (N_13295,N_10947,N_10295);
xnor U13296 (N_13296,N_10382,N_11053);
nor U13297 (N_13297,N_10257,N_10477);
and U13298 (N_13298,N_10126,N_10284);
nor U13299 (N_13299,N_11225,N_11058);
nand U13300 (N_13300,N_11099,N_10989);
or U13301 (N_13301,N_11212,N_10455);
nand U13302 (N_13302,N_11028,N_10838);
and U13303 (N_13303,N_10767,N_11675);
and U13304 (N_13304,N_10971,N_11211);
nor U13305 (N_13305,N_10701,N_11589);
nor U13306 (N_13306,N_11699,N_10401);
and U13307 (N_13307,N_10376,N_10726);
nand U13308 (N_13308,N_10348,N_11289);
or U13309 (N_13309,N_11629,N_10639);
nor U13310 (N_13310,N_11224,N_11898);
nor U13311 (N_13311,N_11688,N_10527);
nand U13312 (N_13312,N_10936,N_11936);
or U13313 (N_13313,N_10824,N_11926);
nor U13314 (N_13314,N_10025,N_11980);
nand U13315 (N_13315,N_11416,N_11163);
and U13316 (N_13316,N_10107,N_10372);
nand U13317 (N_13317,N_10765,N_11329);
nor U13318 (N_13318,N_10460,N_11690);
nor U13319 (N_13319,N_11447,N_11424);
xor U13320 (N_13320,N_10839,N_11003);
and U13321 (N_13321,N_11116,N_11280);
and U13322 (N_13322,N_10288,N_11915);
or U13323 (N_13323,N_10821,N_10289);
or U13324 (N_13324,N_10898,N_10986);
and U13325 (N_13325,N_11552,N_11939);
nand U13326 (N_13326,N_11921,N_11140);
nand U13327 (N_13327,N_11610,N_11351);
and U13328 (N_13328,N_10679,N_11511);
nor U13329 (N_13329,N_11369,N_11695);
nand U13330 (N_13330,N_10993,N_10983);
nor U13331 (N_13331,N_10670,N_10567);
or U13332 (N_13332,N_11291,N_10768);
nand U13333 (N_13333,N_11873,N_11584);
and U13334 (N_13334,N_10882,N_11793);
nor U13335 (N_13335,N_11912,N_10001);
nand U13336 (N_13336,N_10293,N_11703);
and U13337 (N_13337,N_11399,N_10610);
or U13338 (N_13338,N_10733,N_10653);
nand U13339 (N_13339,N_10669,N_11639);
nand U13340 (N_13340,N_10646,N_11620);
and U13341 (N_13341,N_11017,N_11202);
nor U13342 (N_13342,N_10907,N_10635);
and U13343 (N_13343,N_10074,N_10582);
xnor U13344 (N_13344,N_11055,N_10350);
xor U13345 (N_13345,N_10363,N_11239);
or U13346 (N_13346,N_10830,N_10756);
xor U13347 (N_13347,N_11658,N_11332);
and U13348 (N_13348,N_10511,N_10116);
nand U13349 (N_13349,N_10971,N_11454);
or U13350 (N_13350,N_10851,N_10962);
and U13351 (N_13351,N_10284,N_11712);
nand U13352 (N_13352,N_11366,N_11874);
or U13353 (N_13353,N_11118,N_10359);
nor U13354 (N_13354,N_10268,N_10462);
or U13355 (N_13355,N_10712,N_11576);
nand U13356 (N_13356,N_10332,N_11915);
nand U13357 (N_13357,N_11598,N_10499);
or U13358 (N_13358,N_11137,N_11099);
nand U13359 (N_13359,N_10304,N_11943);
nand U13360 (N_13360,N_10573,N_10464);
or U13361 (N_13361,N_10880,N_10958);
or U13362 (N_13362,N_10608,N_11696);
or U13363 (N_13363,N_10473,N_10462);
nor U13364 (N_13364,N_10695,N_10205);
nor U13365 (N_13365,N_10594,N_11753);
and U13366 (N_13366,N_11979,N_10891);
nor U13367 (N_13367,N_11060,N_11468);
or U13368 (N_13368,N_11564,N_10810);
and U13369 (N_13369,N_10519,N_10707);
nand U13370 (N_13370,N_10433,N_11225);
or U13371 (N_13371,N_11514,N_11012);
nand U13372 (N_13372,N_11549,N_10706);
xor U13373 (N_13373,N_10321,N_11905);
nand U13374 (N_13374,N_10386,N_10081);
and U13375 (N_13375,N_10900,N_11086);
nand U13376 (N_13376,N_11058,N_10112);
nor U13377 (N_13377,N_11353,N_10584);
or U13378 (N_13378,N_10789,N_11297);
xnor U13379 (N_13379,N_11100,N_11336);
or U13380 (N_13380,N_10926,N_10661);
and U13381 (N_13381,N_11761,N_10848);
nor U13382 (N_13382,N_10877,N_11660);
nor U13383 (N_13383,N_10106,N_11072);
nand U13384 (N_13384,N_11954,N_11456);
or U13385 (N_13385,N_10954,N_10653);
or U13386 (N_13386,N_11634,N_10678);
or U13387 (N_13387,N_10433,N_11877);
or U13388 (N_13388,N_10713,N_11556);
or U13389 (N_13389,N_10057,N_10333);
nor U13390 (N_13390,N_11951,N_10166);
xor U13391 (N_13391,N_11963,N_11587);
or U13392 (N_13392,N_11959,N_10679);
or U13393 (N_13393,N_10724,N_11836);
and U13394 (N_13394,N_10138,N_10982);
and U13395 (N_13395,N_11205,N_11929);
nand U13396 (N_13396,N_11100,N_10844);
and U13397 (N_13397,N_11503,N_11906);
or U13398 (N_13398,N_10131,N_11945);
or U13399 (N_13399,N_10870,N_11084);
nor U13400 (N_13400,N_10254,N_11496);
nor U13401 (N_13401,N_10571,N_11264);
and U13402 (N_13402,N_11894,N_10172);
nand U13403 (N_13403,N_11182,N_11856);
xor U13404 (N_13404,N_10634,N_11685);
or U13405 (N_13405,N_11116,N_10328);
nor U13406 (N_13406,N_11094,N_11072);
nand U13407 (N_13407,N_10527,N_11593);
xnor U13408 (N_13408,N_11711,N_11108);
nor U13409 (N_13409,N_10088,N_11379);
nand U13410 (N_13410,N_10238,N_10380);
nand U13411 (N_13411,N_11639,N_11070);
nor U13412 (N_13412,N_10706,N_10899);
xor U13413 (N_13413,N_11251,N_11878);
nor U13414 (N_13414,N_10247,N_10399);
xor U13415 (N_13415,N_11843,N_11481);
and U13416 (N_13416,N_11355,N_10552);
nand U13417 (N_13417,N_10646,N_11226);
and U13418 (N_13418,N_11221,N_10063);
nor U13419 (N_13419,N_10418,N_11865);
and U13420 (N_13420,N_11399,N_11824);
and U13421 (N_13421,N_11536,N_11591);
xor U13422 (N_13422,N_10022,N_10954);
and U13423 (N_13423,N_10271,N_10170);
and U13424 (N_13424,N_10593,N_11241);
or U13425 (N_13425,N_10021,N_11430);
xnor U13426 (N_13426,N_10132,N_11820);
or U13427 (N_13427,N_10867,N_10238);
or U13428 (N_13428,N_10143,N_11054);
and U13429 (N_13429,N_11683,N_11742);
xnor U13430 (N_13430,N_10819,N_11784);
nand U13431 (N_13431,N_11134,N_10424);
and U13432 (N_13432,N_11922,N_10766);
nand U13433 (N_13433,N_10365,N_11918);
nand U13434 (N_13434,N_10065,N_10633);
xor U13435 (N_13435,N_11895,N_10520);
nand U13436 (N_13436,N_10123,N_10457);
and U13437 (N_13437,N_11043,N_11456);
nor U13438 (N_13438,N_11353,N_11706);
and U13439 (N_13439,N_11441,N_11588);
and U13440 (N_13440,N_10545,N_11073);
and U13441 (N_13441,N_10150,N_10599);
or U13442 (N_13442,N_10592,N_10889);
or U13443 (N_13443,N_10841,N_11811);
or U13444 (N_13444,N_11591,N_11631);
and U13445 (N_13445,N_10634,N_11568);
or U13446 (N_13446,N_11604,N_11276);
nor U13447 (N_13447,N_11344,N_10189);
and U13448 (N_13448,N_10929,N_10582);
xor U13449 (N_13449,N_10218,N_10200);
nand U13450 (N_13450,N_11964,N_10134);
nor U13451 (N_13451,N_11903,N_10752);
xnor U13452 (N_13452,N_10039,N_10075);
or U13453 (N_13453,N_10976,N_10447);
and U13454 (N_13454,N_11916,N_11547);
xnor U13455 (N_13455,N_11243,N_11490);
nor U13456 (N_13456,N_11980,N_10806);
nor U13457 (N_13457,N_11867,N_10349);
and U13458 (N_13458,N_11904,N_11031);
or U13459 (N_13459,N_10291,N_11525);
nand U13460 (N_13460,N_10590,N_11838);
nor U13461 (N_13461,N_11852,N_10578);
nand U13462 (N_13462,N_11177,N_11415);
xnor U13463 (N_13463,N_10446,N_10375);
and U13464 (N_13464,N_10325,N_11893);
and U13465 (N_13465,N_10906,N_11900);
and U13466 (N_13466,N_10884,N_10633);
or U13467 (N_13467,N_11668,N_10247);
and U13468 (N_13468,N_10992,N_10315);
nand U13469 (N_13469,N_11030,N_10615);
nor U13470 (N_13470,N_10523,N_10248);
and U13471 (N_13471,N_11787,N_10870);
and U13472 (N_13472,N_11243,N_10399);
xnor U13473 (N_13473,N_11165,N_10468);
or U13474 (N_13474,N_10126,N_11292);
or U13475 (N_13475,N_11075,N_10485);
xor U13476 (N_13476,N_10859,N_10527);
and U13477 (N_13477,N_11563,N_10109);
nor U13478 (N_13478,N_11262,N_10788);
and U13479 (N_13479,N_11097,N_11349);
nor U13480 (N_13480,N_10087,N_11623);
or U13481 (N_13481,N_11847,N_11955);
or U13482 (N_13482,N_11264,N_11436);
nand U13483 (N_13483,N_10626,N_10692);
nand U13484 (N_13484,N_11216,N_10136);
and U13485 (N_13485,N_11211,N_11199);
and U13486 (N_13486,N_10527,N_11616);
nand U13487 (N_13487,N_10447,N_11359);
and U13488 (N_13488,N_10359,N_11779);
or U13489 (N_13489,N_11301,N_11428);
nor U13490 (N_13490,N_11652,N_10040);
nand U13491 (N_13491,N_11139,N_10456);
nor U13492 (N_13492,N_10735,N_11370);
nand U13493 (N_13493,N_10289,N_10847);
nor U13494 (N_13494,N_11472,N_11054);
xnor U13495 (N_13495,N_11313,N_10292);
and U13496 (N_13496,N_10709,N_10908);
nand U13497 (N_13497,N_11526,N_10515);
nand U13498 (N_13498,N_10214,N_10701);
nand U13499 (N_13499,N_11052,N_10149);
or U13500 (N_13500,N_11514,N_10406);
nor U13501 (N_13501,N_10518,N_11434);
or U13502 (N_13502,N_10713,N_11083);
or U13503 (N_13503,N_11031,N_11995);
or U13504 (N_13504,N_11092,N_10324);
nor U13505 (N_13505,N_11769,N_10875);
nand U13506 (N_13506,N_10027,N_10876);
or U13507 (N_13507,N_11660,N_10032);
xor U13508 (N_13508,N_11662,N_11474);
or U13509 (N_13509,N_10139,N_10757);
nor U13510 (N_13510,N_11764,N_10961);
or U13511 (N_13511,N_10988,N_11912);
nand U13512 (N_13512,N_11514,N_10236);
and U13513 (N_13513,N_11403,N_11160);
nor U13514 (N_13514,N_10548,N_10466);
nand U13515 (N_13515,N_11784,N_10702);
nand U13516 (N_13516,N_10167,N_11919);
xnor U13517 (N_13517,N_11898,N_10121);
and U13518 (N_13518,N_10394,N_11648);
nor U13519 (N_13519,N_11347,N_11109);
and U13520 (N_13520,N_11895,N_11788);
or U13521 (N_13521,N_11786,N_11736);
xor U13522 (N_13522,N_10205,N_11529);
nand U13523 (N_13523,N_10716,N_10750);
xor U13524 (N_13524,N_10382,N_11879);
and U13525 (N_13525,N_11392,N_10182);
and U13526 (N_13526,N_11565,N_10486);
and U13527 (N_13527,N_10693,N_11737);
xnor U13528 (N_13528,N_10421,N_11511);
or U13529 (N_13529,N_11015,N_11603);
nor U13530 (N_13530,N_10887,N_10360);
and U13531 (N_13531,N_10448,N_11395);
nand U13532 (N_13532,N_10056,N_10720);
nand U13533 (N_13533,N_11059,N_11608);
and U13534 (N_13534,N_10160,N_10958);
xor U13535 (N_13535,N_11363,N_11229);
or U13536 (N_13536,N_11962,N_11380);
nor U13537 (N_13537,N_10962,N_11525);
and U13538 (N_13538,N_11081,N_11664);
and U13539 (N_13539,N_10094,N_10218);
nor U13540 (N_13540,N_11875,N_11628);
and U13541 (N_13541,N_11276,N_10906);
or U13542 (N_13542,N_10101,N_11292);
nand U13543 (N_13543,N_10880,N_11831);
and U13544 (N_13544,N_11777,N_10531);
nand U13545 (N_13545,N_11608,N_10679);
nand U13546 (N_13546,N_11273,N_11149);
and U13547 (N_13547,N_11640,N_11520);
or U13548 (N_13548,N_10996,N_10324);
nor U13549 (N_13549,N_11962,N_11474);
xnor U13550 (N_13550,N_10404,N_10034);
or U13551 (N_13551,N_10640,N_10054);
and U13552 (N_13552,N_10175,N_11238);
or U13553 (N_13553,N_10950,N_10437);
and U13554 (N_13554,N_10860,N_10759);
nand U13555 (N_13555,N_11617,N_10101);
and U13556 (N_13556,N_10970,N_10841);
and U13557 (N_13557,N_10077,N_10593);
and U13558 (N_13558,N_10869,N_11860);
nor U13559 (N_13559,N_10176,N_10407);
nor U13560 (N_13560,N_11544,N_11716);
nor U13561 (N_13561,N_10269,N_11909);
nor U13562 (N_13562,N_11895,N_10591);
or U13563 (N_13563,N_10023,N_11782);
nand U13564 (N_13564,N_10322,N_11815);
nand U13565 (N_13565,N_11814,N_10240);
and U13566 (N_13566,N_11776,N_11283);
nor U13567 (N_13567,N_11450,N_11380);
nor U13568 (N_13568,N_10627,N_10875);
nor U13569 (N_13569,N_11355,N_10510);
nor U13570 (N_13570,N_10371,N_10358);
or U13571 (N_13571,N_10050,N_10840);
xnor U13572 (N_13572,N_10231,N_10944);
xor U13573 (N_13573,N_10298,N_11130);
or U13574 (N_13574,N_11635,N_10441);
or U13575 (N_13575,N_10126,N_10417);
nand U13576 (N_13576,N_10470,N_10568);
and U13577 (N_13577,N_11789,N_11876);
nor U13578 (N_13578,N_10226,N_10060);
nand U13579 (N_13579,N_10819,N_11799);
xnor U13580 (N_13580,N_11486,N_11262);
and U13581 (N_13581,N_10925,N_11311);
nor U13582 (N_13582,N_10730,N_10001);
or U13583 (N_13583,N_11691,N_11178);
xor U13584 (N_13584,N_10609,N_11471);
or U13585 (N_13585,N_10196,N_11085);
nand U13586 (N_13586,N_11299,N_11522);
nor U13587 (N_13587,N_11434,N_11413);
and U13588 (N_13588,N_10498,N_11947);
nor U13589 (N_13589,N_11953,N_11886);
xor U13590 (N_13590,N_11167,N_10279);
nor U13591 (N_13591,N_10735,N_11726);
nand U13592 (N_13592,N_11947,N_10243);
or U13593 (N_13593,N_11528,N_11335);
nor U13594 (N_13594,N_10910,N_11865);
or U13595 (N_13595,N_11042,N_10501);
nor U13596 (N_13596,N_11456,N_11911);
nand U13597 (N_13597,N_10558,N_10483);
and U13598 (N_13598,N_11662,N_10022);
and U13599 (N_13599,N_11525,N_11660);
or U13600 (N_13600,N_10396,N_11064);
xnor U13601 (N_13601,N_10912,N_10270);
or U13602 (N_13602,N_11665,N_11155);
nor U13603 (N_13603,N_10699,N_11483);
nand U13604 (N_13604,N_10610,N_10843);
xnor U13605 (N_13605,N_11894,N_10900);
and U13606 (N_13606,N_11399,N_10216);
and U13607 (N_13607,N_11523,N_10512);
or U13608 (N_13608,N_11469,N_11095);
nor U13609 (N_13609,N_11729,N_11833);
nand U13610 (N_13610,N_11817,N_10247);
nor U13611 (N_13611,N_10810,N_10886);
nor U13612 (N_13612,N_10889,N_11514);
nor U13613 (N_13613,N_11869,N_11916);
xnor U13614 (N_13614,N_11792,N_10873);
xor U13615 (N_13615,N_10096,N_11813);
and U13616 (N_13616,N_10790,N_11403);
and U13617 (N_13617,N_10584,N_10843);
nand U13618 (N_13618,N_11893,N_10371);
or U13619 (N_13619,N_11820,N_10840);
xor U13620 (N_13620,N_11495,N_11003);
xnor U13621 (N_13621,N_11538,N_10504);
nand U13622 (N_13622,N_11355,N_10562);
nand U13623 (N_13623,N_11447,N_10879);
or U13624 (N_13624,N_11333,N_11648);
and U13625 (N_13625,N_10415,N_11866);
or U13626 (N_13626,N_11443,N_11231);
or U13627 (N_13627,N_10185,N_10917);
nand U13628 (N_13628,N_11070,N_11289);
and U13629 (N_13629,N_11198,N_10898);
nor U13630 (N_13630,N_10452,N_10216);
nor U13631 (N_13631,N_10488,N_10425);
or U13632 (N_13632,N_10983,N_10933);
or U13633 (N_13633,N_10439,N_10387);
nand U13634 (N_13634,N_11419,N_10698);
and U13635 (N_13635,N_11709,N_10281);
nand U13636 (N_13636,N_11412,N_11059);
nand U13637 (N_13637,N_11505,N_10389);
and U13638 (N_13638,N_10593,N_11368);
and U13639 (N_13639,N_11338,N_11275);
and U13640 (N_13640,N_11357,N_11817);
nand U13641 (N_13641,N_11071,N_10085);
and U13642 (N_13642,N_11496,N_10348);
nand U13643 (N_13643,N_10192,N_10848);
xor U13644 (N_13644,N_10303,N_11608);
nand U13645 (N_13645,N_11036,N_10589);
xnor U13646 (N_13646,N_11572,N_10315);
and U13647 (N_13647,N_11075,N_10295);
or U13648 (N_13648,N_11259,N_10501);
and U13649 (N_13649,N_11933,N_10356);
and U13650 (N_13650,N_10020,N_10871);
and U13651 (N_13651,N_10422,N_11905);
or U13652 (N_13652,N_10128,N_10160);
and U13653 (N_13653,N_11219,N_10601);
nand U13654 (N_13654,N_10130,N_11028);
and U13655 (N_13655,N_11497,N_10283);
and U13656 (N_13656,N_10845,N_10571);
and U13657 (N_13657,N_11064,N_11311);
and U13658 (N_13658,N_11809,N_11140);
or U13659 (N_13659,N_11811,N_10167);
or U13660 (N_13660,N_11263,N_11421);
and U13661 (N_13661,N_11542,N_11533);
and U13662 (N_13662,N_11554,N_11547);
nor U13663 (N_13663,N_11064,N_10220);
or U13664 (N_13664,N_10275,N_10451);
xor U13665 (N_13665,N_10152,N_10031);
nor U13666 (N_13666,N_10714,N_11856);
nand U13667 (N_13667,N_11589,N_11319);
nor U13668 (N_13668,N_11838,N_10526);
xnor U13669 (N_13669,N_10899,N_11583);
and U13670 (N_13670,N_11853,N_11046);
or U13671 (N_13671,N_11281,N_10360);
nand U13672 (N_13672,N_11208,N_11420);
and U13673 (N_13673,N_10765,N_11338);
nand U13674 (N_13674,N_10004,N_10698);
and U13675 (N_13675,N_10797,N_10920);
and U13676 (N_13676,N_11824,N_10009);
nand U13677 (N_13677,N_10691,N_10024);
nand U13678 (N_13678,N_10676,N_11092);
nor U13679 (N_13679,N_10808,N_11061);
nand U13680 (N_13680,N_10010,N_11366);
or U13681 (N_13681,N_10465,N_11665);
nor U13682 (N_13682,N_10691,N_10233);
nand U13683 (N_13683,N_11330,N_11541);
nand U13684 (N_13684,N_11731,N_10280);
nor U13685 (N_13685,N_11361,N_10024);
nand U13686 (N_13686,N_10664,N_10976);
xnor U13687 (N_13687,N_11193,N_10720);
nand U13688 (N_13688,N_10388,N_11165);
nand U13689 (N_13689,N_11867,N_11743);
xor U13690 (N_13690,N_10150,N_10127);
nor U13691 (N_13691,N_11635,N_11978);
or U13692 (N_13692,N_11221,N_11653);
nor U13693 (N_13693,N_10087,N_10188);
nor U13694 (N_13694,N_10126,N_11580);
or U13695 (N_13695,N_11523,N_10251);
and U13696 (N_13696,N_11081,N_10275);
and U13697 (N_13697,N_10510,N_11762);
nor U13698 (N_13698,N_10309,N_10002);
nor U13699 (N_13699,N_10281,N_11741);
nand U13700 (N_13700,N_11741,N_11718);
nor U13701 (N_13701,N_11917,N_11009);
xor U13702 (N_13702,N_10504,N_11869);
nor U13703 (N_13703,N_11017,N_10718);
nand U13704 (N_13704,N_10170,N_10588);
nand U13705 (N_13705,N_10761,N_10525);
or U13706 (N_13706,N_10959,N_10339);
nand U13707 (N_13707,N_11159,N_10944);
and U13708 (N_13708,N_10861,N_10123);
nor U13709 (N_13709,N_10801,N_10804);
or U13710 (N_13710,N_10332,N_10686);
nor U13711 (N_13711,N_11029,N_11643);
nand U13712 (N_13712,N_10190,N_11647);
nor U13713 (N_13713,N_10989,N_11868);
nand U13714 (N_13714,N_10727,N_10790);
nand U13715 (N_13715,N_11687,N_11580);
xor U13716 (N_13716,N_10595,N_10343);
or U13717 (N_13717,N_11217,N_11401);
and U13718 (N_13718,N_11744,N_10165);
or U13719 (N_13719,N_10848,N_11310);
and U13720 (N_13720,N_10344,N_11391);
nor U13721 (N_13721,N_11108,N_11045);
nor U13722 (N_13722,N_11195,N_11526);
nand U13723 (N_13723,N_11044,N_11017);
nor U13724 (N_13724,N_11996,N_11464);
nand U13725 (N_13725,N_10346,N_11465);
nand U13726 (N_13726,N_11617,N_10442);
or U13727 (N_13727,N_10088,N_11673);
xor U13728 (N_13728,N_10280,N_11612);
nand U13729 (N_13729,N_11900,N_11651);
and U13730 (N_13730,N_10614,N_11360);
nand U13731 (N_13731,N_11834,N_10691);
xor U13732 (N_13732,N_11172,N_10595);
or U13733 (N_13733,N_11905,N_11285);
nand U13734 (N_13734,N_10144,N_11049);
xor U13735 (N_13735,N_10182,N_10128);
or U13736 (N_13736,N_11516,N_10826);
xnor U13737 (N_13737,N_11377,N_10582);
or U13738 (N_13738,N_11692,N_10360);
nor U13739 (N_13739,N_10076,N_10193);
and U13740 (N_13740,N_10607,N_10370);
nand U13741 (N_13741,N_11947,N_11023);
nor U13742 (N_13742,N_11134,N_10402);
xnor U13743 (N_13743,N_11255,N_10935);
or U13744 (N_13744,N_11854,N_10367);
or U13745 (N_13745,N_10054,N_11869);
xor U13746 (N_13746,N_10697,N_11279);
or U13747 (N_13747,N_11010,N_10269);
or U13748 (N_13748,N_10042,N_10639);
nor U13749 (N_13749,N_10540,N_11721);
or U13750 (N_13750,N_10709,N_10898);
and U13751 (N_13751,N_10687,N_11930);
and U13752 (N_13752,N_11342,N_11194);
and U13753 (N_13753,N_10799,N_10278);
and U13754 (N_13754,N_11259,N_10910);
nor U13755 (N_13755,N_11887,N_10538);
nand U13756 (N_13756,N_10001,N_11409);
or U13757 (N_13757,N_11110,N_10217);
and U13758 (N_13758,N_10730,N_11951);
or U13759 (N_13759,N_10106,N_11181);
and U13760 (N_13760,N_10143,N_10524);
and U13761 (N_13761,N_11702,N_11638);
and U13762 (N_13762,N_10091,N_10570);
nor U13763 (N_13763,N_11883,N_11337);
or U13764 (N_13764,N_10843,N_10777);
and U13765 (N_13765,N_10904,N_11980);
and U13766 (N_13766,N_11983,N_10026);
and U13767 (N_13767,N_11175,N_10616);
nor U13768 (N_13768,N_10019,N_10726);
nand U13769 (N_13769,N_11447,N_10390);
nor U13770 (N_13770,N_10828,N_10025);
xnor U13771 (N_13771,N_11410,N_10162);
and U13772 (N_13772,N_11462,N_11364);
or U13773 (N_13773,N_11755,N_10809);
or U13774 (N_13774,N_11872,N_10227);
xnor U13775 (N_13775,N_10269,N_10476);
and U13776 (N_13776,N_10499,N_11428);
nor U13777 (N_13777,N_11810,N_10901);
nand U13778 (N_13778,N_11594,N_10849);
and U13779 (N_13779,N_11997,N_11128);
nor U13780 (N_13780,N_10452,N_10418);
or U13781 (N_13781,N_10140,N_11174);
xnor U13782 (N_13782,N_10889,N_10820);
nand U13783 (N_13783,N_10518,N_10276);
and U13784 (N_13784,N_11404,N_10301);
nand U13785 (N_13785,N_10865,N_10009);
nand U13786 (N_13786,N_10652,N_11458);
and U13787 (N_13787,N_11752,N_11867);
and U13788 (N_13788,N_10285,N_11162);
or U13789 (N_13789,N_10890,N_10929);
and U13790 (N_13790,N_11280,N_10906);
and U13791 (N_13791,N_11339,N_11922);
nand U13792 (N_13792,N_10186,N_10907);
or U13793 (N_13793,N_10237,N_10053);
or U13794 (N_13794,N_10656,N_11246);
nand U13795 (N_13795,N_11642,N_11674);
nor U13796 (N_13796,N_10278,N_11867);
and U13797 (N_13797,N_11394,N_10400);
or U13798 (N_13798,N_11813,N_10458);
nor U13799 (N_13799,N_10484,N_10363);
and U13800 (N_13800,N_11675,N_11962);
or U13801 (N_13801,N_10997,N_11076);
xor U13802 (N_13802,N_11022,N_10796);
and U13803 (N_13803,N_11448,N_10667);
nor U13804 (N_13804,N_11581,N_11866);
or U13805 (N_13805,N_11449,N_10264);
and U13806 (N_13806,N_11904,N_10052);
and U13807 (N_13807,N_11645,N_10692);
nand U13808 (N_13808,N_11508,N_11527);
or U13809 (N_13809,N_11402,N_11822);
or U13810 (N_13810,N_10312,N_10546);
nor U13811 (N_13811,N_10824,N_10309);
nor U13812 (N_13812,N_11876,N_11742);
or U13813 (N_13813,N_10985,N_10454);
nand U13814 (N_13814,N_11543,N_11252);
nor U13815 (N_13815,N_10693,N_11160);
and U13816 (N_13816,N_10207,N_11737);
and U13817 (N_13817,N_11559,N_11822);
xnor U13818 (N_13818,N_11270,N_11948);
nand U13819 (N_13819,N_11408,N_11183);
or U13820 (N_13820,N_11373,N_11103);
or U13821 (N_13821,N_10164,N_10084);
or U13822 (N_13822,N_10584,N_10023);
and U13823 (N_13823,N_11166,N_11842);
nor U13824 (N_13824,N_11880,N_11567);
nand U13825 (N_13825,N_10451,N_10492);
or U13826 (N_13826,N_10395,N_10334);
or U13827 (N_13827,N_10892,N_10209);
nor U13828 (N_13828,N_10854,N_11878);
nor U13829 (N_13829,N_10578,N_11058);
nor U13830 (N_13830,N_10985,N_10961);
xnor U13831 (N_13831,N_10400,N_10283);
nand U13832 (N_13832,N_11000,N_10166);
nor U13833 (N_13833,N_11270,N_11218);
or U13834 (N_13834,N_11280,N_10346);
and U13835 (N_13835,N_10708,N_10534);
or U13836 (N_13836,N_11391,N_10520);
or U13837 (N_13837,N_10907,N_10240);
xnor U13838 (N_13838,N_11248,N_10813);
or U13839 (N_13839,N_10004,N_11107);
or U13840 (N_13840,N_11783,N_10410);
and U13841 (N_13841,N_10772,N_10649);
nor U13842 (N_13842,N_10276,N_10911);
or U13843 (N_13843,N_11313,N_10888);
nand U13844 (N_13844,N_10333,N_11674);
or U13845 (N_13845,N_10532,N_10521);
xnor U13846 (N_13846,N_10081,N_10748);
nor U13847 (N_13847,N_11206,N_10897);
or U13848 (N_13848,N_11107,N_11185);
nor U13849 (N_13849,N_11078,N_10755);
or U13850 (N_13850,N_11327,N_11115);
nor U13851 (N_13851,N_11701,N_11042);
nand U13852 (N_13852,N_11000,N_11625);
nor U13853 (N_13853,N_11009,N_11705);
and U13854 (N_13854,N_11528,N_11006);
or U13855 (N_13855,N_10232,N_10755);
and U13856 (N_13856,N_10835,N_10241);
or U13857 (N_13857,N_11784,N_11550);
nand U13858 (N_13858,N_10246,N_11734);
nand U13859 (N_13859,N_11351,N_10056);
nand U13860 (N_13860,N_11853,N_10292);
nand U13861 (N_13861,N_10003,N_11933);
or U13862 (N_13862,N_11256,N_10759);
nor U13863 (N_13863,N_10692,N_11268);
or U13864 (N_13864,N_10204,N_10114);
nand U13865 (N_13865,N_11154,N_11999);
nand U13866 (N_13866,N_11476,N_10384);
and U13867 (N_13867,N_11130,N_11763);
nand U13868 (N_13868,N_11061,N_11035);
nor U13869 (N_13869,N_11190,N_11134);
or U13870 (N_13870,N_11049,N_11208);
and U13871 (N_13871,N_10229,N_11987);
nand U13872 (N_13872,N_10687,N_11822);
and U13873 (N_13873,N_11986,N_11045);
or U13874 (N_13874,N_11782,N_11787);
nor U13875 (N_13875,N_10904,N_11263);
xnor U13876 (N_13876,N_11544,N_10491);
and U13877 (N_13877,N_11715,N_11013);
or U13878 (N_13878,N_11861,N_11798);
nor U13879 (N_13879,N_11865,N_10729);
nand U13880 (N_13880,N_10274,N_11132);
or U13881 (N_13881,N_10174,N_11139);
xor U13882 (N_13882,N_10680,N_11470);
nand U13883 (N_13883,N_11503,N_10502);
nand U13884 (N_13884,N_11684,N_10184);
or U13885 (N_13885,N_11730,N_10937);
or U13886 (N_13886,N_11651,N_10278);
nand U13887 (N_13887,N_11401,N_10101);
or U13888 (N_13888,N_10253,N_10126);
xnor U13889 (N_13889,N_11918,N_10684);
and U13890 (N_13890,N_10866,N_10359);
and U13891 (N_13891,N_10155,N_11561);
or U13892 (N_13892,N_10373,N_10713);
or U13893 (N_13893,N_11795,N_10845);
xnor U13894 (N_13894,N_10491,N_11217);
or U13895 (N_13895,N_11282,N_11946);
nor U13896 (N_13896,N_11589,N_11725);
or U13897 (N_13897,N_11818,N_10439);
nor U13898 (N_13898,N_10436,N_11609);
xor U13899 (N_13899,N_10132,N_11117);
or U13900 (N_13900,N_11763,N_10653);
nand U13901 (N_13901,N_11287,N_11572);
and U13902 (N_13902,N_11560,N_11942);
or U13903 (N_13903,N_10716,N_10536);
nand U13904 (N_13904,N_11243,N_10807);
nand U13905 (N_13905,N_11155,N_11480);
nor U13906 (N_13906,N_10494,N_10031);
nand U13907 (N_13907,N_11453,N_11862);
nor U13908 (N_13908,N_11634,N_11724);
or U13909 (N_13909,N_11973,N_10804);
or U13910 (N_13910,N_10068,N_10579);
and U13911 (N_13911,N_10223,N_11237);
nor U13912 (N_13912,N_10596,N_11808);
nor U13913 (N_13913,N_11000,N_10306);
nor U13914 (N_13914,N_10301,N_10527);
nor U13915 (N_13915,N_11640,N_10534);
or U13916 (N_13916,N_11495,N_10776);
nor U13917 (N_13917,N_11774,N_10708);
xor U13918 (N_13918,N_11833,N_11764);
and U13919 (N_13919,N_11781,N_10387);
nor U13920 (N_13920,N_10792,N_11315);
nor U13921 (N_13921,N_10860,N_11577);
and U13922 (N_13922,N_10456,N_10273);
nand U13923 (N_13923,N_10876,N_11481);
nor U13924 (N_13924,N_11570,N_11975);
nand U13925 (N_13925,N_11136,N_11780);
and U13926 (N_13926,N_10713,N_10049);
nor U13927 (N_13927,N_11437,N_10630);
nand U13928 (N_13928,N_11526,N_10004);
nor U13929 (N_13929,N_10722,N_10962);
and U13930 (N_13930,N_10473,N_11600);
nor U13931 (N_13931,N_11242,N_11138);
nor U13932 (N_13932,N_10095,N_10281);
nor U13933 (N_13933,N_11645,N_11567);
nand U13934 (N_13934,N_11215,N_10176);
nor U13935 (N_13935,N_11885,N_11809);
and U13936 (N_13936,N_11826,N_11201);
nor U13937 (N_13937,N_11499,N_10890);
nor U13938 (N_13938,N_10529,N_11116);
or U13939 (N_13939,N_10145,N_10431);
or U13940 (N_13940,N_10132,N_10726);
nand U13941 (N_13941,N_10047,N_10184);
or U13942 (N_13942,N_10619,N_10039);
xor U13943 (N_13943,N_10074,N_11201);
nor U13944 (N_13944,N_11547,N_10583);
and U13945 (N_13945,N_10908,N_11382);
or U13946 (N_13946,N_11506,N_10621);
and U13947 (N_13947,N_11779,N_10106);
and U13948 (N_13948,N_10768,N_11796);
or U13949 (N_13949,N_10916,N_11495);
and U13950 (N_13950,N_11578,N_10270);
or U13951 (N_13951,N_11824,N_11556);
or U13952 (N_13952,N_10797,N_11348);
nand U13953 (N_13953,N_11007,N_10137);
or U13954 (N_13954,N_10235,N_11470);
and U13955 (N_13955,N_10114,N_10236);
nor U13956 (N_13956,N_11099,N_11322);
or U13957 (N_13957,N_11729,N_10557);
xor U13958 (N_13958,N_11849,N_10616);
nand U13959 (N_13959,N_11422,N_11073);
and U13960 (N_13960,N_10145,N_10011);
nor U13961 (N_13961,N_10741,N_10391);
nand U13962 (N_13962,N_10792,N_11905);
nand U13963 (N_13963,N_10193,N_11796);
nand U13964 (N_13964,N_11361,N_11686);
nor U13965 (N_13965,N_10820,N_10551);
and U13966 (N_13966,N_11295,N_11734);
nor U13967 (N_13967,N_10864,N_11712);
and U13968 (N_13968,N_10261,N_10114);
xor U13969 (N_13969,N_10038,N_10128);
nand U13970 (N_13970,N_10853,N_11834);
and U13971 (N_13971,N_10591,N_11584);
nand U13972 (N_13972,N_11303,N_10785);
nand U13973 (N_13973,N_10001,N_11283);
nor U13974 (N_13974,N_11817,N_11095);
nand U13975 (N_13975,N_11826,N_10293);
and U13976 (N_13976,N_11076,N_10179);
and U13977 (N_13977,N_11210,N_10523);
xnor U13978 (N_13978,N_10435,N_11713);
or U13979 (N_13979,N_10388,N_10757);
and U13980 (N_13980,N_11579,N_10886);
or U13981 (N_13981,N_11923,N_11252);
nand U13982 (N_13982,N_11973,N_10369);
xnor U13983 (N_13983,N_11249,N_10733);
nand U13984 (N_13984,N_11926,N_10618);
and U13985 (N_13985,N_11773,N_10225);
or U13986 (N_13986,N_11413,N_11315);
or U13987 (N_13987,N_11411,N_10520);
nor U13988 (N_13988,N_10611,N_11198);
and U13989 (N_13989,N_10231,N_11158);
or U13990 (N_13990,N_11053,N_11589);
nor U13991 (N_13991,N_10750,N_11231);
nor U13992 (N_13992,N_11792,N_11727);
xor U13993 (N_13993,N_10036,N_10441);
or U13994 (N_13994,N_10558,N_10235);
and U13995 (N_13995,N_10256,N_11128);
nor U13996 (N_13996,N_10486,N_11592);
nor U13997 (N_13997,N_11654,N_10639);
and U13998 (N_13998,N_11562,N_10690);
nor U13999 (N_13999,N_11651,N_11028);
and U14000 (N_14000,N_12854,N_12131);
nor U14001 (N_14001,N_13138,N_12066);
nand U14002 (N_14002,N_12267,N_13079);
and U14003 (N_14003,N_12242,N_12705);
or U14004 (N_14004,N_12792,N_12771);
or U14005 (N_14005,N_13664,N_13496);
or U14006 (N_14006,N_12880,N_12037);
or U14007 (N_14007,N_12064,N_12121);
xnor U14008 (N_14008,N_12348,N_13192);
or U14009 (N_14009,N_12904,N_12025);
xnor U14010 (N_14010,N_13893,N_12747);
or U14011 (N_14011,N_13176,N_12832);
and U14012 (N_14012,N_13584,N_12351);
nand U14013 (N_14013,N_13678,N_13730);
xnor U14014 (N_14014,N_13284,N_13766);
or U14015 (N_14015,N_12198,N_12767);
xnor U14016 (N_14016,N_13306,N_13157);
and U14017 (N_14017,N_12799,N_13348);
and U14018 (N_14018,N_12769,N_13513);
and U14019 (N_14019,N_13511,N_12754);
nand U14020 (N_14020,N_12777,N_12236);
nor U14021 (N_14021,N_12925,N_12055);
and U14022 (N_14022,N_12495,N_13864);
nand U14023 (N_14023,N_12726,N_12975);
nor U14024 (N_14024,N_13517,N_13793);
or U14025 (N_14025,N_12424,N_12192);
and U14026 (N_14026,N_12572,N_13007);
nand U14027 (N_14027,N_12344,N_13525);
and U14028 (N_14028,N_13540,N_12720);
xor U14029 (N_14029,N_12251,N_12165);
and U14030 (N_14030,N_12691,N_13474);
or U14031 (N_14031,N_12229,N_12846);
nor U14032 (N_14032,N_12523,N_13961);
nand U14033 (N_14033,N_13419,N_12127);
and U14034 (N_14034,N_12544,N_12914);
and U14035 (N_14035,N_12103,N_13287);
nor U14036 (N_14036,N_13870,N_13498);
or U14037 (N_14037,N_13813,N_13705);
nand U14038 (N_14038,N_13376,N_12171);
and U14039 (N_14039,N_13951,N_13797);
and U14040 (N_14040,N_13018,N_12535);
or U14041 (N_14041,N_12428,N_12871);
and U14042 (N_14042,N_13676,N_12390);
nor U14043 (N_14043,N_12094,N_13193);
nor U14044 (N_14044,N_12524,N_12658);
nand U14045 (N_14045,N_12281,N_13729);
nand U14046 (N_14046,N_12892,N_12901);
and U14047 (N_14047,N_12470,N_13072);
and U14048 (N_14048,N_13994,N_12737);
nand U14049 (N_14049,N_12326,N_13697);
and U14050 (N_14050,N_13005,N_13716);
nor U14051 (N_14051,N_13572,N_12261);
nor U14052 (N_14052,N_13317,N_12757);
and U14053 (N_14053,N_13950,N_13330);
and U14054 (N_14054,N_13954,N_13497);
nand U14055 (N_14055,N_12764,N_12178);
nor U14056 (N_14056,N_12987,N_12485);
and U14057 (N_14057,N_12160,N_13354);
nor U14058 (N_14058,N_12296,N_13033);
nor U14059 (N_14059,N_12237,N_12943);
and U14060 (N_14060,N_12598,N_12505);
and U14061 (N_14061,N_12034,N_12033);
nand U14062 (N_14062,N_13050,N_13506);
nand U14063 (N_14063,N_12245,N_12835);
nand U14064 (N_14064,N_13314,N_13381);
nor U14065 (N_14065,N_12389,N_12923);
and U14066 (N_14066,N_13680,N_13651);
nand U14067 (N_14067,N_12665,N_12933);
xnor U14068 (N_14068,N_13089,N_13170);
and U14069 (N_14069,N_13985,N_13605);
nand U14070 (N_14070,N_13930,N_12097);
nand U14071 (N_14071,N_13597,N_12842);
or U14072 (N_14072,N_12466,N_12784);
or U14073 (N_14073,N_12280,N_12942);
nand U14074 (N_14074,N_12869,N_13989);
nor U14075 (N_14075,N_13336,N_12013);
or U14076 (N_14076,N_12785,N_12147);
xnor U14077 (N_14077,N_12973,N_12526);
and U14078 (N_14078,N_12611,N_12681);
nor U14079 (N_14079,N_13475,N_12527);
nor U14080 (N_14080,N_13649,N_12413);
and U14081 (N_14081,N_12459,N_12856);
nor U14082 (N_14082,N_13819,N_13960);
nor U14083 (N_14083,N_13370,N_12490);
nor U14084 (N_14084,N_13812,N_12041);
and U14085 (N_14085,N_12643,N_13167);
nor U14086 (N_14086,N_12656,N_12994);
and U14087 (N_14087,N_13241,N_13899);
nor U14088 (N_14088,N_13095,N_12995);
nand U14089 (N_14089,N_12950,N_12944);
nor U14090 (N_14090,N_13181,N_12986);
nor U14091 (N_14091,N_13739,N_13409);
or U14092 (N_14092,N_13932,N_12885);
and U14093 (N_14093,N_13924,N_12346);
nand U14094 (N_14094,N_13149,N_12060);
nand U14095 (N_14095,N_12126,N_12024);
and U14096 (N_14096,N_12782,N_13830);
or U14097 (N_14097,N_13201,N_13783);
or U14098 (N_14098,N_13957,N_13096);
xor U14099 (N_14099,N_13345,N_12517);
nor U14100 (N_14100,N_13353,N_12168);
xnor U14101 (N_14101,N_13159,N_12708);
or U14102 (N_14102,N_13359,N_12800);
xnor U14103 (N_14103,N_13788,N_12735);
and U14104 (N_14104,N_12197,N_13818);
and U14105 (N_14105,N_12822,N_12476);
or U14106 (N_14106,N_12167,N_13078);
or U14107 (N_14107,N_13615,N_12555);
or U14108 (N_14108,N_12032,N_13626);
and U14109 (N_14109,N_13856,N_12303);
or U14110 (N_14110,N_13097,N_12831);
and U14111 (N_14111,N_13016,N_12633);
xnor U14112 (N_14112,N_12608,N_13561);
nand U14113 (N_14113,N_12453,N_12403);
nor U14114 (N_14114,N_12189,N_13493);
and U14115 (N_14115,N_12780,N_13903);
nand U14116 (N_14116,N_13443,N_12534);
nor U14117 (N_14117,N_13223,N_13148);
or U14118 (N_14118,N_12623,N_13748);
and U14119 (N_14119,N_13792,N_12439);
nand U14120 (N_14120,N_13334,N_12583);
xnor U14121 (N_14121,N_12588,N_12253);
nand U14122 (N_14122,N_13227,N_12514);
or U14123 (N_14123,N_13865,N_13177);
nor U14124 (N_14124,N_13717,N_12661);
nor U14125 (N_14125,N_13900,N_13846);
nor U14126 (N_14126,N_12020,N_13583);
xor U14127 (N_14127,N_13635,N_12778);
and U14128 (N_14128,N_12293,N_12689);
and U14129 (N_14129,N_12112,N_12352);
and U14130 (N_14130,N_13612,N_13065);
and U14131 (N_14131,N_12420,N_12104);
nand U14132 (N_14132,N_12776,N_12905);
nor U14133 (N_14133,N_12012,N_12163);
nand U14134 (N_14134,N_12325,N_12741);
and U14135 (N_14135,N_13160,N_13703);
xnor U14136 (N_14136,N_13294,N_13146);
nor U14137 (N_14137,N_12088,N_13367);
and U14138 (N_14138,N_12157,N_13083);
nor U14139 (N_14139,N_13617,N_13544);
nor U14140 (N_14140,N_12089,N_13045);
and U14141 (N_14141,N_12049,N_13198);
nor U14142 (N_14142,N_13553,N_13028);
or U14143 (N_14143,N_12815,N_12759);
nor U14144 (N_14144,N_13648,N_13161);
and U14145 (N_14145,N_12414,N_12796);
or U14146 (N_14146,N_13022,N_12028);
nand U14147 (N_14147,N_12742,N_13868);
nor U14148 (N_14148,N_13976,N_13530);
nand U14149 (N_14149,N_12627,N_12095);
and U14150 (N_14150,N_12044,N_12662);
nor U14151 (N_14151,N_13945,N_12177);
nand U14152 (N_14152,N_12216,N_12998);
nor U14153 (N_14153,N_12145,N_13158);
and U14154 (N_14154,N_12515,N_12356);
or U14155 (N_14155,N_13189,N_12123);
xor U14156 (N_14156,N_13608,N_13963);
or U14157 (N_14157,N_12212,N_12011);
and U14158 (N_14158,N_13744,N_12309);
nor U14159 (N_14159,N_13549,N_12913);
and U14160 (N_14160,N_13838,N_12077);
and U14161 (N_14161,N_13833,N_12209);
nand U14162 (N_14162,N_12482,N_12614);
or U14163 (N_14163,N_13636,N_13623);
xnor U14164 (N_14164,N_13757,N_13915);
and U14165 (N_14165,N_12391,N_13829);
or U14166 (N_14166,N_13331,N_13880);
and U14167 (N_14167,N_12781,N_12573);
nor U14168 (N_14168,N_13273,N_12117);
and U14169 (N_14169,N_12317,N_12884);
and U14170 (N_14170,N_13172,N_13629);
nand U14171 (N_14171,N_13631,N_12556);
nor U14172 (N_14172,N_13811,N_12124);
nor U14173 (N_14173,N_12429,N_13275);
xnor U14174 (N_14174,N_13430,N_13416);
and U14175 (N_14175,N_12340,N_12738);
nor U14176 (N_14176,N_12158,N_13587);
nor U14177 (N_14177,N_13768,N_13923);
nor U14178 (N_14178,N_12492,N_12829);
nand U14179 (N_14179,N_12603,N_12070);
xor U14180 (N_14180,N_12230,N_12632);
nor U14181 (N_14181,N_12536,N_13239);
xor U14182 (N_14182,N_13199,N_12574);
xor U14183 (N_14183,N_12408,N_13683);
or U14184 (N_14184,N_12957,N_13858);
and U14185 (N_14185,N_12175,N_13059);
nand U14186 (N_14186,N_13745,N_13029);
or U14187 (N_14187,N_13031,N_12920);
nor U14188 (N_14188,N_12810,N_12146);
or U14189 (N_14189,N_12875,N_13175);
nand U14190 (N_14190,N_13279,N_12220);
nor U14191 (N_14191,N_12503,N_12062);
and U14192 (N_14192,N_13413,N_12305);
nor U14193 (N_14193,N_13861,N_13098);
nand U14194 (N_14194,N_12706,N_13435);
nor U14195 (N_14195,N_13290,N_13424);
nor U14196 (N_14196,N_13538,N_12074);
xor U14197 (N_14197,N_12581,N_12010);
and U14198 (N_14198,N_12543,N_13968);
nor U14199 (N_14199,N_13845,N_12926);
nand U14200 (N_14200,N_12442,N_12551);
or U14201 (N_14201,N_12073,N_12313);
nor U14202 (N_14202,N_13388,N_13966);
nor U14203 (N_14203,N_13944,N_12257);
or U14204 (N_14204,N_12762,N_13338);
or U14205 (N_14205,N_12377,N_13836);
xnor U14206 (N_14206,N_13194,N_12756);
nand U14207 (N_14207,N_13820,N_13489);
nand U14208 (N_14208,N_12007,N_13316);
nor U14209 (N_14209,N_13659,N_13088);
nor U14210 (N_14210,N_13313,N_12208);
nand U14211 (N_14211,N_13934,N_13478);
nand U14212 (N_14212,N_13032,N_13888);
nand U14213 (N_14213,N_12223,N_13979);
nand U14214 (N_14214,N_13180,N_12031);
or U14215 (N_14215,N_12723,N_13809);
or U14216 (N_14216,N_13991,N_13816);
nor U14217 (N_14217,N_13779,N_12366);
or U14218 (N_14218,N_13499,N_13441);
and U14219 (N_14219,N_12525,N_13277);
or U14220 (N_14220,N_13070,N_13922);
and U14221 (N_14221,N_12941,N_12059);
or U14222 (N_14222,N_13296,N_12151);
xor U14223 (N_14223,N_12663,N_13415);
nor U14224 (N_14224,N_13222,N_13125);
or U14225 (N_14225,N_12432,N_12761);
or U14226 (N_14226,N_13668,N_12278);
nand U14227 (N_14227,N_13375,N_12787);
xor U14228 (N_14228,N_12248,N_12501);
and U14229 (N_14229,N_12620,N_13295);
and U14230 (N_14230,N_13360,N_12879);
nor U14231 (N_14231,N_12672,N_12903);
or U14232 (N_14232,N_12310,N_12636);
nand U14233 (N_14233,N_12746,N_12946);
nand U14234 (N_14234,N_12697,N_13103);
nor U14235 (N_14235,N_13548,N_12287);
nand U14236 (N_14236,N_12530,N_12316);
or U14237 (N_14237,N_12695,N_12322);
nor U14238 (N_14238,N_12051,N_12203);
nor U14239 (N_14239,N_13974,N_12873);
and U14240 (N_14240,N_13719,N_12646);
nand U14241 (N_14241,N_13644,N_12824);
nand U14242 (N_14242,N_12793,N_13105);
or U14243 (N_14243,N_13469,N_13611);
nand U14244 (N_14244,N_12054,N_13408);
or U14245 (N_14245,N_12692,N_12181);
nor U14246 (N_14246,N_13806,N_12292);
and U14247 (N_14247,N_12794,N_12014);
and U14248 (N_14248,N_13853,N_13586);
nand U14249 (N_14249,N_12455,N_13828);
or U14250 (N_14250,N_12850,N_12898);
nor U14251 (N_14251,N_12407,N_13689);
nor U14252 (N_14252,N_13575,N_13737);
xnor U14253 (N_14253,N_13965,N_13881);
nor U14254 (N_14254,N_12069,N_13302);
or U14255 (N_14255,N_13731,N_12685);
or U14256 (N_14256,N_13885,N_12065);
or U14257 (N_14257,N_13904,N_13318);
and U14258 (N_14258,N_13132,N_13602);
nor U14259 (N_14259,N_12385,N_12789);
nand U14260 (N_14260,N_12022,N_13162);
or U14261 (N_14261,N_13339,N_12865);
xor U14262 (N_14262,N_12225,N_13634);
or U14263 (N_14263,N_12677,N_13406);
xor U14264 (N_14264,N_13484,N_12409);
and U14265 (N_14265,N_12629,N_12830);
or U14266 (N_14266,N_13344,N_13726);
nor U14267 (N_14267,N_13400,N_13077);
or U14268 (N_14268,N_12868,N_13929);
or U14269 (N_14269,N_12595,N_13321);
or U14270 (N_14270,N_13568,N_12451);
or U14271 (N_14271,N_12259,N_13749);
nor U14272 (N_14272,N_12110,N_12788);
nand U14273 (N_14273,N_13195,N_12508);
nor U14274 (N_14274,N_12397,N_12797);
or U14275 (N_14275,N_13799,N_13291);
and U14276 (N_14276,N_12048,N_13850);
nor U14277 (N_14277,N_13849,N_13461);
and U14278 (N_14278,N_12231,N_13217);
nor U14279 (N_14279,N_13735,N_12299);
or U14280 (N_14280,N_12119,N_12773);
nand U14281 (N_14281,N_13448,N_13479);
nand U14282 (N_14282,N_12335,N_12376);
nand U14283 (N_14283,N_12491,N_13606);
nor U14284 (N_14284,N_13431,N_13384);
and U14285 (N_14285,N_13686,N_13271);
or U14286 (N_14286,N_12058,N_12954);
nor U14287 (N_14287,N_13688,N_12602);
nor U14288 (N_14288,N_13564,N_13008);
and U14289 (N_14289,N_12339,N_12255);
or U14290 (N_14290,N_12642,N_13335);
and U14291 (N_14291,N_13472,N_12355);
xor U14292 (N_14292,N_13734,N_13677);
or U14293 (N_14293,N_12113,N_12249);
and U14294 (N_14294,N_13718,N_13949);
xor U14295 (N_14295,N_12162,N_12795);
nor U14296 (N_14296,N_12431,N_13233);
and U14297 (N_14297,N_13589,N_13998);
and U14298 (N_14298,N_13337,N_12380);
nand U14299 (N_14299,N_12387,N_12384);
nand U14300 (N_14300,N_13075,N_13604);
nand U14301 (N_14301,N_13245,N_13808);
xor U14302 (N_14302,N_12132,N_12516);
or U14303 (N_14303,N_13569,N_13129);
nand U14304 (N_14304,N_13449,N_13463);
nor U14305 (N_14305,N_12246,N_12184);
xnor U14306 (N_14306,N_13450,N_13789);
xor U14307 (N_14307,N_13933,N_12053);
and U14308 (N_14308,N_13796,N_12215);
or U14309 (N_14309,N_12654,N_13100);
and U14310 (N_14310,N_12959,N_12276);
or U14311 (N_14311,N_13882,N_12497);
nand U14312 (N_14312,N_12772,N_12176);
or U14313 (N_14313,N_12307,N_13377);
nor U14314 (N_14314,N_12269,N_12506);
and U14315 (N_14315,N_13468,N_12130);
and U14316 (N_14316,N_13872,N_13001);
and U14317 (N_14317,N_12331,N_13996);
or U14318 (N_14318,N_13143,N_13600);
nor U14319 (N_14319,N_13283,N_12847);
nor U14320 (N_14320,N_13365,N_12895);
nor U14321 (N_14321,N_12199,N_13320);
nor U14322 (N_14322,N_13758,N_12838);
nor U14323 (N_14323,N_13082,N_13130);
nor U14324 (N_14324,N_12840,N_13014);
nand U14325 (N_14325,N_12454,N_12148);
nand U14326 (N_14326,N_12382,N_13666);
nand U14327 (N_14327,N_12233,N_13117);
nor U14328 (N_14328,N_12486,N_13554);
or U14329 (N_14329,N_13019,N_13692);
xnor U14330 (N_14330,N_12101,N_12365);
nor U14331 (N_14331,N_12955,N_13988);
and U14332 (N_14332,N_12042,N_12989);
and U14333 (N_14333,N_13978,N_13128);
nor U14334 (N_14334,N_13622,N_12930);
nand U14335 (N_14335,N_12166,N_13570);
or U14336 (N_14336,N_12985,N_12240);
nand U14337 (N_14337,N_12019,N_13567);
nand U14338 (N_14338,N_12128,N_13107);
xnor U14339 (N_14339,N_12308,N_12043);
nand U14340 (N_14340,N_13364,N_13049);
xnor U14341 (N_14341,N_12479,N_13535);
nand U14342 (N_14342,N_13073,N_12717);
nor U14343 (N_14343,N_12279,N_13753);
nand U14344 (N_14344,N_13613,N_12702);
xor U14345 (N_14345,N_13781,N_12564);
and U14346 (N_14346,N_12180,N_12449);
nor U14347 (N_14347,N_13959,N_12272);
nor U14348 (N_14348,N_13147,N_12922);
nor U14349 (N_14349,N_13169,N_13303);
nand U14350 (N_14350,N_13026,N_13462);
xnor U14351 (N_14351,N_13311,N_13706);
or U14352 (N_14352,N_12715,N_12939);
nor U14353 (N_14353,N_12561,N_12586);
nand U14354 (N_14354,N_12820,N_12217);
or U14355 (N_14355,N_13814,N_13747);
or U14356 (N_14356,N_13975,N_12529);
or U14357 (N_14357,N_13051,N_13145);
nand U14358 (N_14358,N_13024,N_13759);
nand U14359 (N_14359,N_12988,N_13660);
or U14360 (N_14360,N_12463,N_13682);
or U14361 (N_14361,N_13052,N_13111);
and U14362 (N_14362,N_13545,N_13067);
or U14363 (N_14363,N_13352,N_12333);
nand U14364 (N_14364,N_12056,N_13732);
or U14365 (N_14365,N_12039,N_13843);
nor U14366 (N_14366,N_12819,N_13973);
or U14367 (N_14367,N_13141,N_12990);
nand U14368 (N_14368,N_12578,N_13531);
nor U14369 (N_14369,N_13183,N_12256);
nand U14370 (N_14370,N_13254,N_13574);
nor U14371 (N_14371,N_13981,N_12727);
or U14372 (N_14372,N_12133,N_12657);
and U14373 (N_14373,N_12202,N_12412);
xor U14374 (N_14374,N_12520,N_13557);
and U14375 (N_14375,N_13543,N_12461);
nand U14376 (N_14376,N_13702,N_12935);
nand U14377 (N_14377,N_13451,N_13514);
nor U14378 (N_14378,N_12640,N_13984);
or U14379 (N_14379,N_12716,N_13310);
nand U14380 (N_14380,N_13956,N_12383);
nor U14381 (N_14381,N_13837,N_12774);
and U14382 (N_14382,N_12206,N_12760);
nand U14383 (N_14383,N_12183,N_13048);
or U14384 (N_14384,N_13342,N_12190);
or U14385 (N_14385,N_12948,N_12770);
xor U14386 (N_14386,N_12908,N_13216);
nand U14387 (N_14387,N_12226,N_13656);
and U14388 (N_14388,N_12559,N_13109);
and U14389 (N_14389,N_12631,N_13857);
and U14390 (N_14390,N_12634,N_12619);
nand U14391 (N_14391,N_13278,N_13698);
or U14392 (N_14392,N_13601,N_12801);
or U14393 (N_14393,N_12809,N_12533);
nand U14394 (N_14394,N_13438,N_13456);
nand U14395 (N_14395,N_13150,N_13684);
nor U14396 (N_14396,N_12857,N_12582);
nor U14397 (N_14397,N_12956,N_13420);
and U14398 (N_14398,N_12813,N_13151);
xnor U14399 (N_14399,N_12638,N_13204);
or U14400 (N_14400,N_13750,N_13723);
or U14401 (N_14401,N_13270,N_12932);
nor U14402 (N_14402,N_12046,N_13361);
nand U14403 (N_14403,N_13867,N_13269);
xnor U14404 (N_14404,N_12244,N_12899);
or U14405 (N_14405,N_13405,N_13209);
and U14406 (N_14406,N_12243,N_12870);
nor U14407 (N_14407,N_13707,N_12188);
nor U14408 (N_14408,N_13765,N_13369);
xor U14409 (N_14409,N_13790,N_13712);
nor U14410 (N_14410,N_13139,N_13063);
nor U14411 (N_14411,N_13910,N_13559);
xnor U14412 (N_14412,N_13418,N_13196);
and U14413 (N_14413,N_12675,N_13154);
or U14414 (N_14414,N_13522,N_12567);
nand U14415 (N_14415,N_12684,N_13743);
or U14416 (N_14416,N_13560,N_13023);
or U14417 (N_14417,N_13693,N_12645);
nand U14418 (N_14418,N_12260,N_12404);
or U14419 (N_14419,N_13822,N_12156);
nand U14420 (N_14420,N_13440,N_13094);
or U14421 (N_14421,N_12550,N_13464);
and U14422 (N_14422,N_13764,N_12538);
or U14423 (N_14423,N_13447,N_13581);
nand U14424 (N_14424,N_13142,N_12068);
and U14425 (N_14425,N_13926,N_12021);
nand U14426 (N_14426,N_12469,N_13661);
or U14427 (N_14427,N_13392,N_13774);
xnor U14428 (N_14428,N_13382,N_12500);
or U14429 (N_14429,N_12775,N_12722);
nand U14430 (N_14430,N_12896,N_13010);
nand U14431 (N_14431,N_13439,N_12766);
or U14432 (N_14432,N_12537,N_13533);
and U14433 (N_14433,N_12982,N_12395);
nor U14434 (N_14434,N_13547,N_12791);
and U14435 (N_14435,N_12086,N_13741);
and U14436 (N_14436,N_13034,N_12639);
and U14437 (N_14437,N_13911,N_12977);
and U14438 (N_14438,N_12858,N_12332);
or U14439 (N_14439,N_12600,N_12265);
or U14440 (N_14440,N_13071,N_13432);
and U14441 (N_14441,N_13665,N_12144);
nor U14442 (N_14442,N_12076,N_12916);
or U14443 (N_14443,N_13247,N_12386);
nor U14444 (N_14444,N_12001,N_12152);
xnor U14445 (N_14445,N_13841,N_13672);
or U14446 (N_14446,N_13437,N_12668);
and U14447 (N_14447,N_12328,N_12698);
nor U14448 (N_14448,N_13596,N_13847);
nor U14449 (N_14449,N_13285,N_12258);
and U14450 (N_14450,N_12493,N_12063);
xor U14451 (N_14451,N_12354,N_12368);
nand U14452 (N_14452,N_12411,N_12301);
or U14453 (N_14453,N_12509,N_13243);
nand U14454 (N_14454,N_12465,N_12828);
nand U14455 (N_14455,N_12604,N_13115);
xor U14456 (N_14456,N_13645,N_13068);
or U14457 (N_14457,N_12890,N_13452);
and U14458 (N_14458,N_13887,N_13218);
and U14459 (N_14459,N_13436,N_12931);
nor U14460 (N_14460,N_13304,N_12000);
and U14461 (N_14461,N_13326,N_12458);
and U14462 (N_14462,N_13041,N_12378);
and U14463 (N_14463,N_13947,N_12125);
nor U14464 (N_14464,N_13952,N_13925);
or U14465 (N_14465,N_12751,N_12297);
nor U14466 (N_14466,N_13658,N_13894);
nor U14467 (N_14467,N_13357,N_12511);
or U14468 (N_14468,N_13886,N_13112);
or U14469 (N_14469,N_12098,N_12628);
nand U14470 (N_14470,N_12472,N_13308);
nand U14471 (N_14471,N_13179,N_12510);
or U14472 (N_14472,N_12252,N_13240);
nor U14473 (N_14473,N_12513,N_13460);
xor U14474 (N_14474,N_13453,N_13268);
and U14475 (N_14475,N_12863,N_13579);
or U14476 (N_14476,N_13417,N_12753);
nand U14477 (N_14477,N_12081,N_12343);
or U14478 (N_14478,N_13999,N_12610);
or U14479 (N_14479,N_12023,N_12005);
nand U14480 (N_14480,N_13491,N_12921);
and U14481 (N_14481,N_12962,N_12521);
nor U14482 (N_14482,N_12438,N_12363);
and U14483 (N_14483,N_13862,N_13770);
xnor U14484 (N_14484,N_13633,N_12498);
xor U14485 (N_14485,N_13669,N_12907);
nand U14486 (N_14486,N_12575,N_12882);
nor U14487 (N_14487,N_12700,N_12504);
and U14488 (N_14488,N_12548,N_13831);
and U14489 (N_14489,N_12765,N_12427);
and U14490 (N_14490,N_12591,N_13044);
nor U14491 (N_14491,N_12002,N_13340);
and U14492 (N_14492,N_12143,N_12690);
nor U14493 (N_14493,N_13883,N_13372);
and U14494 (N_14494,N_12910,N_12963);
xnor U14495 (N_14495,N_12671,N_12290);
and U14496 (N_14496,N_12649,N_12361);
nor U14497 (N_14497,N_13099,N_12972);
or U14498 (N_14498,N_13657,N_13652);
nand U14499 (N_14499,N_12029,N_12277);
and U14500 (N_14500,N_13709,N_12845);
or U14501 (N_14501,N_12379,N_12150);
or U14502 (N_14502,N_12546,N_13740);
nor U14503 (N_14503,N_13912,N_12558);
or U14504 (N_14504,N_13704,N_13775);
nand U14505 (N_14505,N_12234,N_12418);
nand U14506 (N_14506,N_12839,N_12008);
or U14507 (N_14507,N_13523,N_13234);
nand U14508 (N_14508,N_13992,N_12441);
nand U14509 (N_14509,N_13394,N_12360);
nand U14510 (N_14510,N_12139,N_13242);
or U14511 (N_14511,N_13558,N_12109);
and U14512 (N_14512,N_13835,N_12239);
and U14513 (N_14513,N_13208,N_12483);
and U14514 (N_14514,N_12666,N_12283);
xnor U14515 (N_14515,N_12596,N_13200);
xnor U14516 (N_14516,N_12833,N_12349);
and U14517 (N_14517,N_13492,N_12855);
nand U14518 (N_14518,N_12878,N_12860);
nand U14519 (N_14519,N_13896,N_12512);
xnor U14520 (N_14520,N_12653,N_13066);
nand U14521 (N_14521,N_12035,N_13153);
nor U14522 (N_14522,N_12318,N_13329);
and U14523 (N_14523,N_12211,N_12618);
nor U14524 (N_14524,N_13650,N_13509);
nor U14525 (N_14525,N_12091,N_13038);
nand U14526 (N_14526,N_12375,N_13914);
or U14527 (N_14527,N_13319,N_12435);
xnor U14528 (N_14528,N_12090,N_12194);
nand U14529 (N_14529,N_13173,N_12732);
or U14530 (N_14530,N_12474,N_12545);
or U14531 (N_14531,N_13715,N_12704);
nor U14532 (N_14532,N_13685,N_13537);
and U14533 (N_14533,N_13264,N_13126);
nor U14534 (N_14534,N_13632,N_12319);
and U14535 (N_14535,N_12853,N_13391);
or U14536 (N_14536,N_12866,N_13322);
xnor U14537 (N_14537,N_12997,N_12410);
nand U14538 (N_14538,N_13913,N_13387);
xnor U14539 (N_14539,N_12302,N_13058);
or U14540 (N_14540,N_12464,N_13446);
nand U14541 (N_14541,N_13238,N_13800);
nand U14542 (N_14542,N_13997,N_12017);
and U14543 (N_14543,N_13309,N_13210);
and U14544 (N_14544,N_13501,N_13039);
or U14545 (N_14545,N_13795,N_13905);
or U14546 (N_14546,N_13398,N_12731);
nor U14547 (N_14547,N_13724,N_13494);
and U14548 (N_14548,N_12953,N_12739);
nand U14549 (N_14549,N_12802,N_12467);
xnor U14550 (N_14550,N_13378,N_12607);
nor U14551 (N_14551,N_13733,N_13445);
nor U14552 (N_14552,N_12709,N_12321);
and U14553 (N_14553,N_12422,N_13211);
and U14554 (N_14554,N_12547,N_13002);
nand U14555 (N_14555,N_12961,N_13580);
nand U14556 (N_14556,N_13347,N_13694);
and U14557 (N_14557,N_13519,N_13742);
nor U14558 (N_14558,N_13490,N_12481);
and U14559 (N_14559,N_13798,N_12593);
xor U14560 (N_14560,N_13476,N_13371);
or U14561 (N_14561,N_12009,N_13889);
and U14562 (N_14562,N_12122,N_13054);
xnor U14563 (N_14563,N_12334,N_12811);
and U14564 (N_14564,N_13520,N_13871);
nand U14565 (N_14565,N_12003,N_13423);
nand U14566 (N_14566,N_13108,N_12915);
xnor U14567 (N_14567,N_13137,N_13346);
or U14568 (N_14568,N_12447,N_12338);
nor U14569 (N_14569,N_13422,N_13232);
and U14570 (N_14570,N_13654,N_13231);
or U14571 (N_14571,N_12728,N_13972);
and U14572 (N_14572,N_13266,N_12312);
xnor U14573 (N_14573,N_13892,N_12185);
nand U14574 (N_14574,N_12528,N_13226);
or U14575 (N_14575,N_12952,N_12398);
nand U14576 (N_14576,N_13860,N_12625);
or U14577 (N_14577,N_13552,N_13197);
xnor U14578 (N_14578,N_12291,N_13970);
and U14579 (N_14579,N_12193,N_12118);
and U14580 (N_14580,N_12195,N_13401);
nand U14581 (N_14581,N_12266,N_12655);
nand U14582 (N_14582,N_13516,N_12949);
or U14583 (N_14583,N_12693,N_13842);
nand U14584 (N_14584,N_12883,N_13228);
or U14585 (N_14585,N_12696,N_13875);
nor U14586 (N_14586,N_13118,N_13315);
nand U14587 (N_14587,N_13582,N_12745);
nand U14588 (N_14588,N_13555,N_13508);
nor U14589 (N_14589,N_12577,N_12947);
nand U14590 (N_14590,N_13297,N_12200);
nor U14591 (N_14591,N_13121,N_12889);
or U14592 (N_14592,N_12480,N_13958);
and U14593 (N_14593,N_13168,N_13935);
and U14594 (N_14594,N_13465,N_13986);
and U14595 (N_14595,N_13598,N_12342);
nand U14596 (N_14596,N_13133,N_12918);
nand U14597 (N_14597,N_12494,N_13414);
nand U14598 (N_14598,N_13752,N_13395);
nand U14599 (N_14599,N_13257,N_13573);
nor U14600 (N_14600,N_13165,N_13466);
and U14601 (N_14601,N_13086,N_12075);
nor U14602 (N_14602,N_12964,N_12659);
nor U14603 (N_14603,N_13866,N_12238);
nand U14604 (N_14604,N_12664,N_13119);
and U14605 (N_14605,N_13990,N_12273);
nor U14606 (N_14606,N_12394,N_12680);
or U14607 (N_14607,N_13021,N_13186);
nand U14608 (N_14608,N_12440,N_13455);
nor U14609 (N_14609,N_13220,N_12864);
nand U14610 (N_14610,N_13203,N_12734);
nor U14611 (N_14611,N_12740,N_13485);
xor U14612 (N_14612,N_12660,N_12247);
or U14613 (N_14613,N_13879,N_13953);
nand U14614 (N_14614,N_13515,N_12803);
xor U14615 (N_14615,N_12979,N_13349);
or U14616 (N_14616,N_13917,N_12980);
nor U14617 (N_14617,N_12609,N_12733);
nor U14618 (N_14618,N_13873,N_13943);
nand U14619 (N_14619,N_12817,N_12562);
and U14620 (N_14620,N_12900,N_13471);
or U14621 (N_14621,N_13607,N_13069);
and U14622 (N_14622,N_12730,N_13874);
or U14623 (N_14623,N_13013,N_12324);
nor U14624 (N_14624,N_12288,N_13164);
nand U14625 (N_14625,N_12207,N_13628);
nor U14626 (N_14626,N_13721,N_13794);
or U14627 (N_14627,N_12306,N_12976);
or U14628 (N_14628,N_13043,N_13341);
nand U14629 (N_14629,N_13120,N_12067);
or U14630 (N_14630,N_13012,N_13618);
or U14631 (N_14631,N_12093,N_13738);
nand U14632 (N_14632,N_12539,N_13093);
and U14633 (N_14633,N_13614,N_12204);
nand U14634 (N_14634,N_12912,N_13259);
nor U14635 (N_14635,N_12841,N_13834);
nor U14636 (N_14636,N_13504,N_13131);
nand U14637 (N_14637,N_12592,N_13603);
and U14638 (N_14638,N_13638,N_12456);
nor U14639 (N_14639,N_13332,N_12057);
nor U14640 (N_14640,N_12004,N_12417);
or U14641 (N_14641,N_13003,N_12140);
nor U14642 (N_14642,N_13076,N_13720);
or U14643 (N_14643,N_12106,N_13276);
nand U14644 (N_14644,N_13403,N_12676);
nor U14645 (N_14645,N_13116,N_13529);
or U14646 (N_14646,N_13769,N_13594);
and U14647 (N_14647,N_13102,N_13546);
nor U14648 (N_14648,N_13434,N_12298);
or U14649 (N_14649,N_13062,N_12674);
xor U14650 (N_14650,N_13385,N_13207);
and U14651 (N_14651,N_13713,N_13967);
or U14652 (N_14652,N_13675,N_12170);
nand U14653 (N_14653,N_12262,N_13328);
and U14654 (N_14654,N_12872,N_13256);
and U14655 (N_14655,N_12960,N_13937);
or U14656 (N_14656,N_12566,N_13566);
nor U14657 (N_14657,N_13487,N_12647);
nor U14658 (N_14658,N_13363,N_12228);
nand U14659 (N_14659,N_13655,N_12396);
nand U14660 (N_14660,N_12748,N_13939);
nor U14661 (N_14661,N_12852,N_12701);
nand U14662 (N_14662,N_12568,N_12268);
nor U14663 (N_14663,N_12392,N_13585);
nor U14664 (N_14664,N_12285,N_12750);
nor U14665 (N_14665,N_12475,N_12902);
nor U14666 (N_14666,N_12129,N_12108);
nand U14667 (N_14667,N_13215,N_12393);
xor U14668 (N_14668,N_12254,N_13620);
nand U14669 (N_14669,N_12703,N_13980);
nand U14670 (N_14670,N_13263,N_13246);
nor U14671 (N_14671,N_13576,N_12711);
nor U14672 (N_14672,N_13772,N_13433);
nand U14673 (N_14673,N_13237,N_13884);
nand U14674 (N_14674,N_13562,N_12488);
nand U14675 (N_14675,N_12372,N_12201);
or U14676 (N_14676,N_13667,N_12958);
nand U14677 (N_14677,N_13642,N_12560);
xor U14678 (N_14678,N_12981,N_13187);
and U14679 (N_14679,N_12423,N_12937);
nor U14680 (N_14680,N_12359,N_13085);
xor U14681 (N_14681,N_13791,N_13827);
nor U14682 (N_14682,N_12499,N_12874);
xor U14683 (N_14683,N_12137,N_12082);
nand U14684 (N_14684,N_12218,N_13495);
or U14685 (N_14685,N_13902,N_12214);
nor U14686 (N_14686,N_13470,N_13272);
nor U14687 (N_14687,N_13127,N_13824);
xor U14688 (N_14688,N_13258,N_12174);
and U14689 (N_14689,N_13897,N_12554);
nand U14690 (N_14690,N_13020,N_12585);
nor U14691 (N_14691,N_12861,N_12936);
and U14692 (N_14692,N_13876,N_12083);
nor U14693 (N_14693,N_13687,N_13056);
nand U14694 (N_14694,N_12909,N_12191);
xor U14695 (N_14695,N_12138,N_12489);
or U14696 (N_14696,N_12725,N_13110);
nor U14697 (N_14697,N_13477,N_13253);
nand U14698 (N_14698,N_13760,N_12182);
xor U14699 (N_14699,N_12616,N_13616);
nand U14700 (N_14700,N_12818,N_12169);
or U14701 (N_14701,N_13941,N_12434);
or U14702 (N_14702,N_13286,N_13969);
nand U14703 (N_14703,N_13877,N_13380);
nor U14704 (N_14704,N_12315,N_13389);
xor U14705 (N_14705,N_13852,N_12341);
nand U14706 (N_14706,N_12768,N_12388);
nor U14707 (N_14707,N_12807,N_13163);
and U14708 (N_14708,N_12477,N_13407);
nand U14709 (N_14709,N_13591,N_12263);
or U14710 (N_14710,N_13588,N_13323);
nor U14711 (N_14711,N_13803,N_13249);
nor U14712 (N_14712,N_13289,N_12992);
or U14713 (N_14713,N_12134,N_13025);
or U14714 (N_14714,N_13305,N_13293);
nor U14715 (N_14715,N_12808,N_13411);
nor U14716 (N_14716,N_12615,N_12084);
and U14717 (N_14717,N_13662,N_12891);
nor U14718 (N_14718,N_12460,N_13244);
nand U14719 (N_14719,N_12471,N_13483);
nor U14720 (N_14720,N_13442,N_12849);
xnor U14721 (N_14721,N_12016,N_13184);
nand U14722 (N_14722,N_12507,N_13927);
nand U14723 (N_14723,N_13444,N_12589);
or U14724 (N_14724,N_12522,N_13521);
xnor U14725 (N_14725,N_13909,N_12650);
nor U14726 (N_14726,N_13637,N_13274);
nand U14727 (N_14727,N_12061,N_12402);
nand U14728 (N_14728,N_12862,N_13936);
or U14729 (N_14729,N_12844,N_12786);
and U14730 (N_14730,N_12314,N_13639);
nor U14731 (N_14731,N_13851,N_12219);
or U14732 (N_14732,N_12232,N_12473);
and U14733 (N_14733,N_13235,N_12928);
nand U14734 (N_14734,N_13810,N_13373);
nor U14735 (N_14735,N_13236,N_12951);
or U14736 (N_14736,N_12116,N_12336);
nand U14737 (N_14737,N_13754,N_13280);
nand U14738 (N_14738,N_13505,N_12940);
nor U14739 (N_14739,N_13593,N_13512);
or U14740 (N_14740,N_13004,N_12938);
nor U14741 (N_14741,N_12330,N_13938);
nor U14742 (N_14742,N_13036,N_12679);
nor U14743 (N_14743,N_13262,N_12092);
nand U14744 (N_14744,N_12984,N_13890);
or U14745 (N_14745,N_13728,N_13224);
nor U14746 (N_14746,N_12018,N_13482);
and U14747 (N_14747,N_12637,N_12644);
or U14748 (N_14748,N_13844,N_12087);
nor U14749 (N_14749,N_12848,N_12719);
nor U14750 (N_14750,N_12271,N_13532);
nand U14751 (N_14751,N_12295,N_13817);
nor U14752 (N_14752,N_12250,N_12927);
nor U14753 (N_14753,N_12173,N_13832);
nand U14754 (N_14754,N_13312,N_13815);
nand U14755 (N_14755,N_13534,N_12805);
xnor U14756 (N_14756,N_13011,N_13480);
nor U14757 (N_14757,N_12945,N_12078);
nor U14758 (N_14758,N_12906,N_13551);
nand U14759 (N_14759,N_13777,N_13190);
nand U14760 (N_14760,N_12729,N_13178);
nand U14761 (N_14761,N_12448,N_12478);
or U14762 (N_14762,N_13805,N_13895);
nand U14763 (N_14763,N_12282,N_12999);
nor U14764 (N_14764,N_13299,N_12599);
and U14765 (N_14765,N_13124,N_12821);
and U14766 (N_14766,N_13114,N_13599);
nand U14767 (N_14767,N_13691,N_13854);
or U14768 (N_14768,N_13397,N_13901);
or U14769 (N_14769,N_12161,N_13000);
xnor U14770 (N_14770,N_12264,N_13518);
and U14771 (N_14771,N_12135,N_12040);
or U14772 (N_14772,N_13009,N_13592);
xor U14773 (N_14773,N_12758,N_12172);
nand U14774 (N_14774,N_13987,N_12405);
and U14775 (N_14775,N_13404,N_12590);
or U14776 (N_14776,N_12678,N_12641);
nor U14777 (N_14777,N_12584,N_12496);
nor U14778 (N_14778,N_13630,N_13977);
nand U14779 (N_14779,N_13571,N_13106);
or U14780 (N_14780,N_13122,N_12834);
nor U14781 (N_14781,N_13964,N_13060);
nor U14782 (N_14782,N_12816,N_13412);
nand U14783 (N_14783,N_12362,N_13425);
and U14784 (N_14784,N_13113,N_13057);
or U14785 (N_14785,N_12996,N_12694);
nand U14786 (N_14786,N_13653,N_13042);
xor U14787 (N_14787,N_12450,N_13307);
and U14788 (N_14788,N_13467,N_13647);
or U14789 (N_14789,N_12099,N_12686);
or U14790 (N_14790,N_12155,N_13459);
nand U14791 (N_14791,N_13502,N_12688);
or U14792 (N_14792,N_13017,N_12399);
xnor U14793 (N_14793,N_12519,N_12886);
nand U14794 (N_14794,N_13393,N_13955);
xor U14795 (N_14795,N_12721,N_12851);
nor U14796 (N_14796,N_12345,N_13982);
nor U14797 (N_14797,N_12430,N_13174);
nor U14798 (N_14798,N_12580,N_12827);
nand U14799 (N_14799,N_13486,N_12426);
or U14800 (N_14800,N_13940,N_13962);
nand U14801 (N_14801,N_13428,N_13214);
nand U14802 (N_14802,N_13248,N_13080);
nand U14803 (N_14803,N_13090,N_13681);
and U14804 (N_14804,N_12783,N_12983);
and U14805 (N_14805,N_12210,N_13251);
xnor U14806 (N_14806,N_13971,N_13092);
and U14807 (N_14807,N_12993,N_12710);
nor U14808 (N_14808,N_12120,N_12736);
or U14809 (N_14809,N_12141,N_12045);
nor U14810 (N_14810,N_13776,N_13383);
or U14811 (N_14811,N_13536,N_13565);
and U14812 (N_14812,N_12823,N_13061);
or U14813 (N_14813,N_13379,N_12888);
and U14814 (N_14814,N_12867,N_12576);
nand U14815 (N_14815,N_13261,N_13621);
nand U14816 (N_14816,N_12337,N_13916);
or U14817 (N_14817,N_13301,N_13763);
nor U14818 (N_14818,N_12713,N_13087);
and U14819 (N_14819,N_13427,N_12924);
and U14820 (N_14820,N_12699,N_13690);
or U14821 (N_14821,N_12683,N_13784);
and U14822 (N_14822,N_13807,N_13942);
nor U14823 (N_14823,N_13983,N_12531);
nor U14824 (N_14824,N_13255,N_13786);
nor U14825 (N_14825,N_12179,N_13577);
xor U14826 (N_14826,N_12542,N_13578);
nor U14827 (N_14827,N_13140,N_12224);
or U14828 (N_14828,N_12401,N_13212);
and U14829 (N_14829,N_13185,N_12353);
or U14830 (N_14830,N_13767,N_12552);
and U14831 (N_14831,N_13804,N_12241);
or U14832 (N_14832,N_12613,N_13358);
nand U14833 (N_14833,N_12294,N_12015);
nor U14834 (N_14834,N_13995,N_13027);
nor U14835 (N_14835,N_12859,N_12502);
xor U14836 (N_14836,N_13627,N_13053);
and U14837 (N_14837,N_13823,N_12036);
nand U14838 (N_14838,N_12601,N_12357);
or U14839 (N_14839,N_12425,N_13761);
nand U14840 (N_14840,N_13035,N_12102);
xnor U14841 (N_14841,N_12755,N_13205);
or U14842 (N_14842,N_13030,N_13037);
and U14843 (N_14843,N_13646,N_12443);
nor U14844 (N_14844,N_13663,N_12114);
or U14845 (N_14845,N_12347,N_12071);
nor U14846 (N_14846,N_13458,N_12630);
or U14847 (N_14847,N_13134,N_12487);
nand U14848 (N_14848,N_12806,N_12436);
or U14849 (N_14849,N_12779,N_13055);
or U14850 (N_14850,N_13206,N_13640);
nand U14851 (N_14851,N_13643,N_12557);
or U14852 (N_14852,N_12804,N_13454);
or U14853 (N_14853,N_13155,N_13221);
or U14854 (N_14854,N_12648,N_12714);
and U14855 (N_14855,N_12669,N_13481);
xnor U14856 (N_14856,N_12374,N_13182);
or U14857 (N_14857,N_13500,N_12622);
nor U14858 (N_14858,N_13671,N_12159);
xnor U14859 (N_14859,N_12164,N_13773);
and U14860 (N_14860,N_12919,N_13152);
xnor U14861 (N_14861,N_12187,N_12416);
or U14862 (N_14862,N_13736,N_13429);
nand U14863 (N_14863,N_12718,N_12897);
nor U14864 (N_14864,N_12100,N_13641);
nor U14865 (N_14865,N_12894,N_13333);
nor U14866 (N_14866,N_12826,N_12457);
and U14867 (N_14867,N_12626,N_12350);
nand U14868 (N_14868,N_12052,N_13590);
or U14869 (N_14869,N_13386,N_13402);
and U14870 (N_14870,N_13993,N_13840);
xnor U14871 (N_14871,N_12367,N_13046);
nor U14872 (N_14872,N_12370,N_12876);
nor U14873 (N_14873,N_13679,N_12752);
and U14874 (N_14874,N_13488,N_13906);
or U14875 (N_14875,N_13219,N_12462);
nor U14876 (N_14876,N_12227,N_12111);
xnor U14877 (N_14877,N_13563,N_12594);
and U14878 (N_14878,N_12437,N_13229);
nand U14879 (N_14879,N_13366,N_13526);
nand U14880 (N_14880,N_13542,N_13281);
or U14881 (N_14881,N_13267,N_12991);
or U14882 (N_14882,N_12814,N_12687);
nor U14883 (N_14883,N_13918,N_13368);
or U14884 (N_14884,N_13390,N_13746);
nor U14885 (N_14885,N_12651,N_12154);
nor U14886 (N_14886,N_12038,N_13695);
and U14887 (N_14887,N_13821,N_13780);
and U14888 (N_14888,N_12274,N_12917);
nand U14889 (N_14889,N_13878,N_12877);
nand U14890 (N_14890,N_12468,N_13006);
nor U14891 (N_14891,N_13144,N_12825);
and U14892 (N_14892,N_13674,N_12978);
nor U14893 (N_14893,N_13710,N_12030);
and U14894 (N_14894,N_13528,N_12235);
or U14895 (N_14895,N_12186,N_12652);
and U14896 (N_14896,N_13699,N_12540);
nor U14897 (N_14897,N_12222,N_12970);
or U14898 (N_14898,N_13324,N_13751);
nor U14899 (N_14899,N_12763,N_12284);
xor U14900 (N_14900,N_13782,N_12749);
and U14901 (N_14901,N_13421,N_12969);
nand U14902 (N_14902,N_13550,N_12579);
and U14903 (N_14903,N_13202,N_13931);
nor U14904 (N_14904,N_12080,N_12587);
nor U14905 (N_14905,N_13839,N_13171);
and U14906 (N_14906,N_13188,N_12381);
nor U14907 (N_14907,N_13946,N_13040);
or U14908 (N_14908,N_13785,N_12635);
nand U14909 (N_14909,N_13300,N_12971);
nor U14910 (N_14910,N_12929,N_12597);
xnor U14911 (N_14911,N_12286,N_12006);
and U14912 (N_14912,N_13081,N_12532);
nand U14913 (N_14913,N_13252,N_12105);
nand U14914 (N_14914,N_13399,N_13524);
nor U14915 (N_14915,N_13362,N_13541);
and U14916 (N_14916,N_12881,N_12452);
nor U14917 (N_14917,N_12724,N_13771);
nand U14918 (N_14918,N_12446,N_13701);
or U14919 (N_14919,N_13595,N_12670);
or U14920 (N_14920,N_12221,N_13919);
nand U14921 (N_14921,N_13104,N_13426);
and U14922 (N_14922,N_12743,N_12744);
nand U14923 (N_14923,N_12373,N_12115);
or U14924 (N_14924,N_13624,N_13230);
and U14925 (N_14925,N_12569,N_13225);
nor U14926 (N_14926,N_12136,N_12707);
nor U14927 (N_14927,N_13265,N_13350);
nor U14928 (N_14928,N_13325,N_12327);
nor U14929 (N_14929,N_12605,N_12079);
and U14930 (N_14930,N_13825,N_12606);
nor U14931 (N_14931,N_12887,N_13670);
xnor U14932 (N_14932,N_13503,N_12270);
nand U14933 (N_14933,N_13787,N_12541);
nand U14934 (N_14934,N_13727,N_13527);
or U14935 (N_14935,N_13711,N_13848);
and U14936 (N_14936,N_12484,N_12565);
or U14937 (N_14937,N_13282,N_12149);
and U14938 (N_14938,N_13074,N_13457);
nand U14939 (N_14939,N_13064,N_13755);
nor U14940 (N_14940,N_12419,N_12444);
nand U14941 (N_14941,N_13539,N_12966);
nor U14942 (N_14942,N_13625,N_12790);
or U14943 (N_14943,N_13250,N_12320);
and U14944 (N_14944,N_13135,N_12712);
nand U14945 (N_14945,N_12518,N_12974);
or U14946 (N_14946,N_12300,N_13725);
and U14947 (N_14947,N_12549,N_13374);
and U14948 (N_14948,N_13351,N_12213);
xor U14949 (N_14949,N_13756,N_12400);
and U14950 (N_14950,N_13123,N_13288);
and U14951 (N_14951,N_12289,N_12911);
nand U14952 (N_14952,N_12553,N_13869);
nor U14953 (N_14953,N_12682,N_13473);
and U14954 (N_14954,N_13355,N_13556);
or U14955 (N_14955,N_13801,N_13898);
and U14956 (N_14956,N_12934,N_12196);
and U14957 (N_14957,N_13260,N_12406);
nor U14958 (N_14958,N_12205,N_13863);
nand U14959 (N_14959,N_12893,N_12433);
and U14960 (N_14960,N_12445,N_12275);
or U14961 (N_14961,N_12798,N_13609);
nand U14962 (N_14962,N_12323,N_13213);
and U14963 (N_14963,N_13166,N_12624);
or U14964 (N_14964,N_13327,N_12617);
nor U14965 (N_14965,N_13619,N_13778);
and U14966 (N_14966,N_12085,N_12570);
and U14967 (N_14967,N_13156,N_13700);
nand U14968 (N_14968,N_12358,N_12836);
nor U14969 (N_14969,N_13891,N_12107);
nor U14970 (N_14970,N_13047,N_12027);
and U14971 (N_14971,N_12329,N_13298);
or U14972 (N_14972,N_13510,N_13855);
and U14973 (N_14973,N_13714,N_12843);
nand U14974 (N_14974,N_13920,N_12364);
or U14975 (N_14975,N_12369,N_13908);
xor U14976 (N_14976,N_13696,N_13292);
nor U14977 (N_14977,N_12812,N_13410);
or U14978 (N_14978,N_13948,N_13802);
and U14979 (N_14979,N_12142,N_12371);
or U14980 (N_14980,N_12612,N_13708);
or U14981 (N_14981,N_13610,N_13907);
or U14982 (N_14982,N_13356,N_13928);
nor U14983 (N_14983,N_13396,N_13859);
or U14984 (N_14984,N_12837,N_12026);
or U14985 (N_14985,N_12667,N_12153);
and U14986 (N_14986,N_12673,N_13921);
nand U14987 (N_14987,N_12050,N_12965);
nor U14988 (N_14988,N_12415,N_12571);
nand U14989 (N_14989,N_13015,N_12563);
nor U14990 (N_14990,N_13136,N_13826);
or U14991 (N_14991,N_13762,N_13722);
nand U14992 (N_14992,N_13507,N_13101);
and U14993 (N_14993,N_12096,N_13091);
nand U14994 (N_14994,N_13673,N_12304);
nand U14995 (N_14995,N_12047,N_12072);
nand U14996 (N_14996,N_13343,N_13084);
nand U14997 (N_14997,N_12967,N_12621);
xor U14998 (N_14998,N_12311,N_13191);
and U14999 (N_14999,N_12968,N_12421);
or U15000 (N_15000,N_13787,N_13659);
and U15001 (N_15001,N_12650,N_12188);
nand U15002 (N_15002,N_13701,N_12974);
nand U15003 (N_15003,N_13597,N_12801);
or U15004 (N_15004,N_13815,N_12456);
and U15005 (N_15005,N_12878,N_13791);
or U15006 (N_15006,N_12192,N_13171);
nand U15007 (N_15007,N_13195,N_13003);
and U15008 (N_15008,N_12056,N_12938);
and U15009 (N_15009,N_13945,N_12216);
nand U15010 (N_15010,N_13049,N_12049);
and U15011 (N_15011,N_12437,N_13677);
nor U15012 (N_15012,N_13724,N_12757);
xnor U15013 (N_15013,N_13814,N_13840);
nand U15014 (N_15014,N_12971,N_12578);
xor U15015 (N_15015,N_13238,N_13272);
nor U15016 (N_15016,N_12644,N_12614);
or U15017 (N_15017,N_13883,N_13056);
or U15018 (N_15018,N_13154,N_12595);
nor U15019 (N_15019,N_13755,N_13093);
and U15020 (N_15020,N_13909,N_12690);
nor U15021 (N_15021,N_13078,N_12053);
xor U15022 (N_15022,N_13503,N_13886);
nor U15023 (N_15023,N_12747,N_13451);
or U15024 (N_15024,N_13718,N_13330);
or U15025 (N_15025,N_13074,N_13372);
nor U15026 (N_15026,N_13002,N_12683);
xor U15027 (N_15027,N_12706,N_13710);
nor U15028 (N_15028,N_13942,N_12506);
nand U15029 (N_15029,N_12295,N_12507);
and U15030 (N_15030,N_13888,N_13968);
nand U15031 (N_15031,N_13927,N_13912);
nand U15032 (N_15032,N_13239,N_13826);
and U15033 (N_15033,N_13012,N_12745);
and U15034 (N_15034,N_13876,N_13760);
and U15035 (N_15035,N_13688,N_12879);
and U15036 (N_15036,N_13966,N_12095);
xnor U15037 (N_15037,N_13387,N_12579);
and U15038 (N_15038,N_13437,N_12096);
nor U15039 (N_15039,N_12962,N_12205);
and U15040 (N_15040,N_13811,N_12855);
and U15041 (N_15041,N_12897,N_13652);
nor U15042 (N_15042,N_12390,N_12444);
or U15043 (N_15043,N_13548,N_12909);
or U15044 (N_15044,N_13739,N_12444);
nor U15045 (N_15045,N_13283,N_13385);
and U15046 (N_15046,N_13490,N_13211);
or U15047 (N_15047,N_13574,N_13836);
and U15048 (N_15048,N_12438,N_13321);
or U15049 (N_15049,N_13594,N_13789);
nor U15050 (N_15050,N_13996,N_12343);
xor U15051 (N_15051,N_13231,N_12792);
and U15052 (N_15052,N_12639,N_13117);
and U15053 (N_15053,N_13324,N_13011);
or U15054 (N_15054,N_13525,N_12219);
nand U15055 (N_15055,N_12972,N_12007);
nand U15056 (N_15056,N_13276,N_13376);
nor U15057 (N_15057,N_13982,N_12004);
nand U15058 (N_15058,N_13504,N_13045);
and U15059 (N_15059,N_12992,N_13955);
and U15060 (N_15060,N_13655,N_13573);
and U15061 (N_15061,N_12147,N_13169);
or U15062 (N_15062,N_12082,N_12926);
and U15063 (N_15063,N_12029,N_13083);
nor U15064 (N_15064,N_13605,N_13476);
nor U15065 (N_15065,N_12926,N_12245);
and U15066 (N_15066,N_13837,N_12360);
xor U15067 (N_15067,N_13468,N_12505);
nor U15068 (N_15068,N_13753,N_12687);
or U15069 (N_15069,N_12266,N_13452);
and U15070 (N_15070,N_12419,N_12489);
nor U15071 (N_15071,N_13114,N_13505);
nor U15072 (N_15072,N_13214,N_13895);
xnor U15073 (N_15073,N_13476,N_12498);
nor U15074 (N_15074,N_13437,N_13168);
xor U15075 (N_15075,N_13408,N_13567);
or U15076 (N_15076,N_13507,N_13437);
xnor U15077 (N_15077,N_13525,N_13364);
nand U15078 (N_15078,N_13262,N_13161);
nand U15079 (N_15079,N_12726,N_12277);
xnor U15080 (N_15080,N_12357,N_12717);
xnor U15081 (N_15081,N_12767,N_12511);
or U15082 (N_15082,N_13759,N_13380);
or U15083 (N_15083,N_13266,N_13254);
nand U15084 (N_15084,N_12058,N_12525);
and U15085 (N_15085,N_12370,N_12661);
nor U15086 (N_15086,N_12136,N_12553);
and U15087 (N_15087,N_12459,N_12314);
or U15088 (N_15088,N_13019,N_13287);
and U15089 (N_15089,N_12812,N_13045);
nand U15090 (N_15090,N_12973,N_13269);
nand U15091 (N_15091,N_12322,N_12224);
or U15092 (N_15092,N_13955,N_13370);
xor U15093 (N_15093,N_12779,N_12767);
or U15094 (N_15094,N_12146,N_12357);
or U15095 (N_15095,N_13966,N_13043);
nor U15096 (N_15096,N_12928,N_13548);
xnor U15097 (N_15097,N_12999,N_12420);
or U15098 (N_15098,N_13593,N_12609);
or U15099 (N_15099,N_12372,N_12159);
nor U15100 (N_15100,N_13057,N_12773);
nand U15101 (N_15101,N_13755,N_12478);
nand U15102 (N_15102,N_12341,N_13049);
or U15103 (N_15103,N_12118,N_13518);
and U15104 (N_15104,N_13809,N_13950);
and U15105 (N_15105,N_13792,N_12328);
or U15106 (N_15106,N_12803,N_13002);
or U15107 (N_15107,N_13401,N_13040);
xnor U15108 (N_15108,N_13277,N_13519);
nand U15109 (N_15109,N_13648,N_12519);
xor U15110 (N_15110,N_12219,N_12845);
nand U15111 (N_15111,N_13542,N_13427);
and U15112 (N_15112,N_13011,N_13131);
nor U15113 (N_15113,N_12007,N_12644);
nor U15114 (N_15114,N_13335,N_12355);
or U15115 (N_15115,N_13242,N_12529);
or U15116 (N_15116,N_13755,N_13138);
nand U15117 (N_15117,N_12994,N_12688);
nand U15118 (N_15118,N_12317,N_12624);
nand U15119 (N_15119,N_13577,N_13509);
nor U15120 (N_15120,N_13545,N_13994);
or U15121 (N_15121,N_13240,N_12360);
nand U15122 (N_15122,N_12831,N_12559);
nand U15123 (N_15123,N_12516,N_12439);
nand U15124 (N_15124,N_13067,N_13237);
or U15125 (N_15125,N_12533,N_13127);
or U15126 (N_15126,N_12832,N_13683);
nor U15127 (N_15127,N_12437,N_12186);
nand U15128 (N_15128,N_12139,N_12644);
or U15129 (N_15129,N_13799,N_13789);
nor U15130 (N_15130,N_12431,N_12081);
or U15131 (N_15131,N_13930,N_12211);
and U15132 (N_15132,N_12089,N_13620);
xor U15133 (N_15133,N_12230,N_12052);
nor U15134 (N_15134,N_13303,N_12872);
nand U15135 (N_15135,N_12229,N_13892);
nand U15136 (N_15136,N_12417,N_13160);
or U15137 (N_15137,N_13116,N_13222);
and U15138 (N_15138,N_12285,N_12691);
nand U15139 (N_15139,N_12024,N_13489);
nand U15140 (N_15140,N_12011,N_13175);
or U15141 (N_15141,N_12404,N_12277);
or U15142 (N_15142,N_13887,N_12855);
nand U15143 (N_15143,N_12245,N_13587);
or U15144 (N_15144,N_12897,N_12004);
and U15145 (N_15145,N_12953,N_13475);
and U15146 (N_15146,N_12245,N_12811);
or U15147 (N_15147,N_13036,N_12412);
nand U15148 (N_15148,N_12232,N_13507);
xnor U15149 (N_15149,N_13616,N_12118);
xnor U15150 (N_15150,N_12945,N_12632);
xnor U15151 (N_15151,N_13688,N_13083);
nand U15152 (N_15152,N_13380,N_12626);
or U15153 (N_15153,N_12913,N_12480);
nand U15154 (N_15154,N_12225,N_13369);
nand U15155 (N_15155,N_12682,N_12352);
nor U15156 (N_15156,N_13438,N_12865);
or U15157 (N_15157,N_13992,N_12668);
nor U15158 (N_15158,N_13865,N_12382);
nand U15159 (N_15159,N_12957,N_13341);
nand U15160 (N_15160,N_13106,N_12803);
nor U15161 (N_15161,N_12464,N_12415);
and U15162 (N_15162,N_12129,N_13476);
or U15163 (N_15163,N_12839,N_12189);
and U15164 (N_15164,N_12474,N_12561);
nor U15165 (N_15165,N_13019,N_12692);
xor U15166 (N_15166,N_13557,N_12684);
nor U15167 (N_15167,N_12839,N_12091);
nand U15168 (N_15168,N_13469,N_12686);
xnor U15169 (N_15169,N_13116,N_13142);
and U15170 (N_15170,N_12463,N_13343);
and U15171 (N_15171,N_13191,N_13166);
and U15172 (N_15172,N_13179,N_13843);
and U15173 (N_15173,N_13226,N_12663);
nand U15174 (N_15174,N_12567,N_13083);
nand U15175 (N_15175,N_12736,N_13917);
nand U15176 (N_15176,N_13773,N_12908);
or U15177 (N_15177,N_13489,N_12565);
and U15178 (N_15178,N_13243,N_12792);
and U15179 (N_15179,N_12190,N_12753);
nor U15180 (N_15180,N_12934,N_13642);
nand U15181 (N_15181,N_12517,N_12378);
nand U15182 (N_15182,N_13488,N_12066);
nor U15183 (N_15183,N_13820,N_12288);
or U15184 (N_15184,N_12576,N_13547);
nor U15185 (N_15185,N_13997,N_12505);
or U15186 (N_15186,N_12143,N_12649);
nand U15187 (N_15187,N_12356,N_13795);
and U15188 (N_15188,N_13742,N_13149);
or U15189 (N_15189,N_13794,N_13780);
nor U15190 (N_15190,N_12216,N_12165);
or U15191 (N_15191,N_12709,N_12382);
or U15192 (N_15192,N_13545,N_12825);
nor U15193 (N_15193,N_13558,N_12566);
nand U15194 (N_15194,N_12468,N_13840);
nand U15195 (N_15195,N_13887,N_12516);
and U15196 (N_15196,N_12735,N_12284);
or U15197 (N_15197,N_12645,N_12340);
nor U15198 (N_15198,N_13890,N_12764);
nor U15199 (N_15199,N_13192,N_13970);
nand U15200 (N_15200,N_13136,N_13523);
and U15201 (N_15201,N_13966,N_12989);
nand U15202 (N_15202,N_12931,N_13577);
nor U15203 (N_15203,N_13624,N_13298);
nor U15204 (N_15204,N_12739,N_13195);
nor U15205 (N_15205,N_13345,N_12810);
nand U15206 (N_15206,N_13218,N_13968);
nand U15207 (N_15207,N_12440,N_13704);
or U15208 (N_15208,N_12016,N_12456);
or U15209 (N_15209,N_12233,N_12919);
or U15210 (N_15210,N_12283,N_12931);
xnor U15211 (N_15211,N_12041,N_12214);
nand U15212 (N_15212,N_12788,N_13404);
xnor U15213 (N_15213,N_12120,N_13678);
or U15214 (N_15214,N_13868,N_12847);
nor U15215 (N_15215,N_12252,N_13863);
and U15216 (N_15216,N_12037,N_12986);
nand U15217 (N_15217,N_12597,N_13818);
nor U15218 (N_15218,N_13636,N_12872);
or U15219 (N_15219,N_12561,N_12851);
or U15220 (N_15220,N_13470,N_12955);
or U15221 (N_15221,N_13382,N_13302);
nand U15222 (N_15222,N_12599,N_12100);
nor U15223 (N_15223,N_12972,N_12321);
or U15224 (N_15224,N_13094,N_13635);
and U15225 (N_15225,N_12927,N_13132);
nand U15226 (N_15226,N_12451,N_12832);
nor U15227 (N_15227,N_12226,N_12905);
and U15228 (N_15228,N_13402,N_12661);
nor U15229 (N_15229,N_13287,N_13348);
or U15230 (N_15230,N_13616,N_13681);
nand U15231 (N_15231,N_12000,N_12083);
nor U15232 (N_15232,N_12049,N_12030);
or U15233 (N_15233,N_12046,N_13044);
or U15234 (N_15234,N_13716,N_13020);
nor U15235 (N_15235,N_13884,N_13712);
xor U15236 (N_15236,N_12863,N_12777);
nand U15237 (N_15237,N_13096,N_13337);
nor U15238 (N_15238,N_13669,N_13378);
nand U15239 (N_15239,N_12869,N_12659);
nand U15240 (N_15240,N_12763,N_13850);
xnor U15241 (N_15241,N_12623,N_12092);
nand U15242 (N_15242,N_12743,N_12741);
nand U15243 (N_15243,N_12234,N_13489);
xor U15244 (N_15244,N_13506,N_13568);
and U15245 (N_15245,N_13545,N_12718);
and U15246 (N_15246,N_13489,N_12308);
nand U15247 (N_15247,N_12793,N_12512);
xnor U15248 (N_15248,N_13614,N_12442);
and U15249 (N_15249,N_13499,N_12024);
nand U15250 (N_15250,N_13174,N_12653);
xor U15251 (N_15251,N_13686,N_12410);
xnor U15252 (N_15252,N_13097,N_13878);
and U15253 (N_15253,N_13492,N_13990);
nand U15254 (N_15254,N_12867,N_12887);
or U15255 (N_15255,N_13407,N_12375);
nand U15256 (N_15256,N_13105,N_12512);
nor U15257 (N_15257,N_13304,N_13182);
xor U15258 (N_15258,N_13424,N_12269);
nand U15259 (N_15259,N_13469,N_12055);
or U15260 (N_15260,N_13964,N_13632);
xor U15261 (N_15261,N_12451,N_12101);
nand U15262 (N_15262,N_13234,N_12274);
and U15263 (N_15263,N_12584,N_12019);
nor U15264 (N_15264,N_12164,N_13808);
nor U15265 (N_15265,N_13427,N_12740);
or U15266 (N_15266,N_12674,N_12883);
nor U15267 (N_15267,N_13944,N_12865);
nand U15268 (N_15268,N_12161,N_12119);
and U15269 (N_15269,N_13813,N_12530);
or U15270 (N_15270,N_12841,N_13785);
xnor U15271 (N_15271,N_12630,N_12453);
or U15272 (N_15272,N_12744,N_13020);
xor U15273 (N_15273,N_13332,N_13521);
nor U15274 (N_15274,N_13753,N_13443);
nand U15275 (N_15275,N_13217,N_13617);
and U15276 (N_15276,N_13757,N_12023);
xor U15277 (N_15277,N_13988,N_13953);
nand U15278 (N_15278,N_13581,N_13324);
nor U15279 (N_15279,N_13221,N_13444);
nor U15280 (N_15280,N_13992,N_13383);
and U15281 (N_15281,N_13152,N_13229);
xnor U15282 (N_15282,N_12894,N_12343);
and U15283 (N_15283,N_12074,N_12631);
xnor U15284 (N_15284,N_13454,N_13473);
nor U15285 (N_15285,N_13066,N_12947);
and U15286 (N_15286,N_12070,N_13192);
nand U15287 (N_15287,N_12261,N_13996);
nor U15288 (N_15288,N_12940,N_13659);
xor U15289 (N_15289,N_12611,N_13102);
or U15290 (N_15290,N_13707,N_13794);
and U15291 (N_15291,N_12165,N_12862);
nor U15292 (N_15292,N_13454,N_13546);
xor U15293 (N_15293,N_12901,N_13990);
and U15294 (N_15294,N_13793,N_12012);
and U15295 (N_15295,N_12756,N_13323);
or U15296 (N_15296,N_13882,N_12868);
nor U15297 (N_15297,N_13053,N_12622);
or U15298 (N_15298,N_13669,N_13946);
nor U15299 (N_15299,N_13708,N_13571);
nor U15300 (N_15300,N_13400,N_13571);
or U15301 (N_15301,N_12962,N_12447);
nor U15302 (N_15302,N_13246,N_12157);
nand U15303 (N_15303,N_12717,N_13687);
or U15304 (N_15304,N_13792,N_13152);
xor U15305 (N_15305,N_12993,N_12423);
and U15306 (N_15306,N_13041,N_13767);
nand U15307 (N_15307,N_12506,N_12733);
nand U15308 (N_15308,N_12155,N_13100);
xor U15309 (N_15309,N_13603,N_13042);
or U15310 (N_15310,N_13633,N_12786);
nand U15311 (N_15311,N_13494,N_12881);
or U15312 (N_15312,N_12050,N_13043);
nand U15313 (N_15313,N_13342,N_12693);
and U15314 (N_15314,N_12158,N_13014);
xnor U15315 (N_15315,N_13176,N_13679);
and U15316 (N_15316,N_12157,N_12905);
and U15317 (N_15317,N_13182,N_12077);
and U15318 (N_15318,N_13352,N_13970);
or U15319 (N_15319,N_13987,N_13739);
and U15320 (N_15320,N_13039,N_13545);
and U15321 (N_15321,N_12996,N_12745);
nor U15322 (N_15322,N_12446,N_13095);
nor U15323 (N_15323,N_12162,N_12675);
nand U15324 (N_15324,N_12553,N_13339);
nand U15325 (N_15325,N_12317,N_12075);
nor U15326 (N_15326,N_12967,N_13560);
nand U15327 (N_15327,N_13487,N_12791);
and U15328 (N_15328,N_13580,N_12662);
and U15329 (N_15329,N_12644,N_12124);
nor U15330 (N_15330,N_12984,N_13487);
nor U15331 (N_15331,N_12571,N_13972);
or U15332 (N_15332,N_12673,N_12882);
and U15333 (N_15333,N_13467,N_13650);
nand U15334 (N_15334,N_13318,N_13319);
nand U15335 (N_15335,N_13501,N_13779);
and U15336 (N_15336,N_12465,N_13764);
nand U15337 (N_15337,N_13783,N_12611);
nor U15338 (N_15338,N_12561,N_12845);
or U15339 (N_15339,N_12213,N_13524);
nand U15340 (N_15340,N_12598,N_12247);
or U15341 (N_15341,N_12309,N_12727);
nand U15342 (N_15342,N_13662,N_13250);
nor U15343 (N_15343,N_13581,N_13085);
or U15344 (N_15344,N_13962,N_13475);
nor U15345 (N_15345,N_12639,N_12735);
xnor U15346 (N_15346,N_13992,N_12909);
and U15347 (N_15347,N_12571,N_13567);
and U15348 (N_15348,N_12116,N_13265);
or U15349 (N_15349,N_12825,N_12691);
or U15350 (N_15350,N_12256,N_13349);
or U15351 (N_15351,N_13654,N_13772);
nor U15352 (N_15352,N_12767,N_12732);
and U15353 (N_15353,N_13097,N_13914);
nor U15354 (N_15354,N_13521,N_13063);
and U15355 (N_15355,N_13390,N_13106);
nand U15356 (N_15356,N_13982,N_13351);
and U15357 (N_15357,N_13729,N_12544);
or U15358 (N_15358,N_12702,N_12501);
nand U15359 (N_15359,N_13732,N_12375);
nor U15360 (N_15360,N_13237,N_13582);
or U15361 (N_15361,N_12002,N_13592);
nand U15362 (N_15362,N_12665,N_13599);
or U15363 (N_15363,N_13463,N_12314);
and U15364 (N_15364,N_12271,N_12266);
nor U15365 (N_15365,N_13811,N_12309);
nand U15366 (N_15366,N_13052,N_12129);
or U15367 (N_15367,N_13101,N_13040);
nand U15368 (N_15368,N_12834,N_13208);
and U15369 (N_15369,N_12059,N_12513);
or U15370 (N_15370,N_12606,N_12058);
or U15371 (N_15371,N_12688,N_13291);
nor U15372 (N_15372,N_13384,N_13946);
nand U15373 (N_15373,N_13605,N_13761);
or U15374 (N_15374,N_13007,N_13305);
xor U15375 (N_15375,N_12924,N_13444);
nand U15376 (N_15376,N_13968,N_13219);
or U15377 (N_15377,N_13014,N_12613);
and U15378 (N_15378,N_12913,N_13738);
nand U15379 (N_15379,N_12496,N_13015);
and U15380 (N_15380,N_13015,N_13572);
nand U15381 (N_15381,N_12868,N_12858);
xor U15382 (N_15382,N_13764,N_13401);
or U15383 (N_15383,N_13372,N_13815);
or U15384 (N_15384,N_12638,N_12831);
nor U15385 (N_15385,N_13447,N_12863);
xor U15386 (N_15386,N_12470,N_12108);
xor U15387 (N_15387,N_13446,N_12822);
nor U15388 (N_15388,N_13559,N_12951);
or U15389 (N_15389,N_12118,N_13857);
xor U15390 (N_15390,N_13207,N_13286);
or U15391 (N_15391,N_12243,N_13878);
nor U15392 (N_15392,N_12716,N_12292);
nand U15393 (N_15393,N_13490,N_13507);
xor U15394 (N_15394,N_12098,N_12589);
nor U15395 (N_15395,N_12144,N_12804);
xnor U15396 (N_15396,N_12466,N_13901);
nor U15397 (N_15397,N_12226,N_13335);
nand U15398 (N_15398,N_12782,N_12615);
nor U15399 (N_15399,N_13825,N_13662);
nand U15400 (N_15400,N_13196,N_13347);
or U15401 (N_15401,N_13339,N_13585);
or U15402 (N_15402,N_12135,N_13538);
nand U15403 (N_15403,N_13133,N_12471);
nor U15404 (N_15404,N_13924,N_13705);
nor U15405 (N_15405,N_13256,N_13575);
nand U15406 (N_15406,N_13909,N_13728);
xor U15407 (N_15407,N_12202,N_13424);
nand U15408 (N_15408,N_12820,N_12160);
or U15409 (N_15409,N_13826,N_13186);
or U15410 (N_15410,N_13478,N_12416);
xor U15411 (N_15411,N_13961,N_12751);
nor U15412 (N_15412,N_13435,N_12534);
and U15413 (N_15413,N_12989,N_13050);
and U15414 (N_15414,N_13215,N_13256);
or U15415 (N_15415,N_13401,N_12286);
and U15416 (N_15416,N_12676,N_13138);
nand U15417 (N_15417,N_12141,N_13892);
or U15418 (N_15418,N_13675,N_12204);
nand U15419 (N_15419,N_13992,N_13847);
nand U15420 (N_15420,N_12379,N_13389);
and U15421 (N_15421,N_12178,N_12413);
and U15422 (N_15422,N_12197,N_12020);
nand U15423 (N_15423,N_13917,N_13906);
or U15424 (N_15424,N_12099,N_12550);
or U15425 (N_15425,N_13074,N_13249);
nand U15426 (N_15426,N_12384,N_13797);
and U15427 (N_15427,N_13727,N_12418);
nand U15428 (N_15428,N_13692,N_12524);
xnor U15429 (N_15429,N_12153,N_12189);
or U15430 (N_15430,N_13798,N_13575);
xnor U15431 (N_15431,N_12375,N_13651);
nand U15432 (N_15432,N_13900,N_13548);
nor U15433 (N_15433,N_13797,N_13415);
and U15434 (N_15434,N_13806,N_12209);
nor U15435 (N_15435,N_13402,N_13508);
or U15436 (N_15436,N_13408,N_12458);
or U15437 (N_15437,N_12878,N_12616);
or U15438 (N_15438,N_12432,N_13766);
nand U15439 (N_15439,N_13260,N_13544);
nand U15440 (N_15440,N_12792,N_13701);
or U15441 (N_15441,N_13125,N_13803);
and U15442 (N_15442,N_12672,N_12565);
and U15443 (N_15443,N_13171,N_12822);
nor U15444 (N_15444,N_12740,N_13300);
and U15445 (N_15445,N_13026,N_13876);
xnor U15446 (N_15446,N_12426,N_13399);
or U15447 (N_15447,N_12111,N_13778);
nor U15448 (N_15448,N_13276,N_12502);
or U15449 (N_15449,N_12932,N_13094);
xor U15450 (N_15450,N_12869,N_12106);
xnor U15451 (N_15451,N_12833,N_13695);
or U15452 (N_15452,N_13552,N_13493);
or U15453 (N_15453,N_13124,N_12238);
nor U15454 (N_15454,N_13565,N_13781);
or U15455 (N_15455,N_13398,N_13304);
xnor U15456 (N_15456,N_12022,N_12309);
or U15457 (N_15457,N_12970,N_12769);
and U15458 (N_15458,N_13034,N_13916);
and U15459 (N_15459,N_13783,N_12943);
and U15460 (N_15460,N_13265,N_12424);
and U15461 (N_15461,N_12086,N_13504);
xnor U15462 (N_15462,N_13736,N_13640);
or U15463 (N_15463,N_13480,N_13726);
nor U15464 (N_15464,N_13429,N_12672);
xnor U15465 (N_15465,N_12847,N_13610);
or U15466 (N_15466,N_13197,N_12160);
and U15467 (N_15467,N_12834,N_12039);
and U15468 (N_15468,N_12484,N_12949);
nand U15469 (N_15469,N_13880,N_13143);
and U15470 (N_15470,N_12805,N_12122);
xnor U15471 (N_15471,N_12199,N_12065);
nand U15472 (N_15472,N_13194,N_12581);
and U15473 (N_15473,N_12512,N_13440);
nor U15474 (N_15474,N_12746,N_13015);
nand U15475 (N_15475,N_13396,N_13450);
nor U15476 (N_15476,N_13613,N_13067);
nand U15477 (N_15477,N_13638,N_12110);
and U15478 (N_15478,N_12134,N_12414);
or U15479 (N_15479,N_12763,N_12752);
and U15480 (N_15480,N_12527,N_12769);
nand U15481 (N_15481,N_13962,N_12206);
or U15482 (N_15482,N_12129,N_13586);
or U15483 (N_15483,N_13229,N_13635);
nand U15484 (N_15484,N_13511,N_12920);
or U15485 (N_15485,N_13124,N_12579);
nand U15486 (N_15486,N_12103,N_12929);
nand U15487 (N_15487,N_12143,N_12226);
nor U15488 (N_15488,N_12610,N_12727);
nand U15489 (N_15489,N_12279,N_12913);
nor U15490 (N_15490,N_13862,N_13061);
or U15491 (N_15491,N_12136,N_12175);
or U15492 (N_15492,N_13886,N_12571);
nor U15493 (N_15493,N_12296,N_13183);
xnor U15494 (N_15494,N_12823,N_13917);
nand U15495 (N_15495,N_12966,N_13709);
xor U15496 (N_15496,N_13102,N_12220);
nor U15497 (N_15497,N_13846,N_13737);
or U15498 (N_15498,N_13401,N_13571);
and U15499 (N_15499,N_12337,N_13552);
nor U15500 (N_15500,N_13806,N_12787);
nor U15501 (N_15501,N_13360,N_12304);
nor U15502 (N_15502,N_13582,N_12949);
xnor U15503 (N_15503,N_12047,N_13006);
and U15504 (N_15504,N_13187,N_12359);
nor U15505 (N_15505,N_12497,N_12819);
and U15506 (N_15506,N_12299,N_12414);
or U15507 (N_15507,N_12019,N_13299);
and U15508 (N_15508,N_13544,N_12851);
or U15509 (N_15509,N_12131,N_12872);
nand U15510 (N_15510,N_13545,N_13085);
nor U15511 (N_15511,N_12738,N_13912);
or U15512 (N_15512,N_12533,N_13450);
or U15513 (N_15513,N_13747,N_13232);
and U15514 (N_15514,N_13188,N_13268);
or U15515 (N_15515,N_13062,N_12351);
and U15516 (N_15516,N_13854,N_13335);
and U15517 (N_15517,N_12150,N_13803);
nand U15518 (N_15518,N_12701,N_13046);
nor U15519 (N_15519,N_13381,N_13065);
nand U15520 (N_15520,N_12850,N_13840);
nand U15521 (N_15521,N_12910,N_12667);
nor U15522 (N_15522,N_12757,N_12963);
and U15523 (N_15523,N_12178,N_13546);
nand U15524 (N_15524,N_12931,N_13458);
nand U15525 (N_15525,N_13142,N_13851);
and U15526 (N_15526,N_12732,N_12918);
nand U15527 (N_15527,N_13148,N_13663);
and U15528 (N_15528,N_13613,N_12398);
and U15529 (N_15529,N_12297,N_13246);
and U15530 (N_15530,N_13564,N_12176);
nor U15531 (N_15531,N_12858,N_12253);
nor U15532 (N_15532,N_13345,N_13353);
nand U15533 (N_15533,N_13338,N_12458);
or U15534 (N_15534,N_13086,N_13514);
nand U15535 (N_15535,N_12213,N_12081);
nand U15536 (N_15536,N_13857,N_13445);
or U15537 (N_15537,N_12593,N_12868);
and U15538 (N_15538,N_12968,N_13622);
and U15539 (N_15539,N_13358,N_13879);
nand U15540 (N_15540,N_12180,N_12074);
nor U15541 (N_15541,N_12549,N_13460);
nor U15542 (N_15542,N_13810,N_12649);
nor U15543 (N_15543,N_13510,N_13905);
nor U15544 (N_15544,N_12022,N_13409);
or U15545 (N_15545,N_13274,N_13907);
or U15546 (N_15546,N_12447,N_13565);
nor U15547 (N_15547,N_13766,N_12619);
and U15548 (N_15548,N_13924,N_12687);
or U15549 (N_15549,N_13802,N_12495);
or U15550 (N_15550,N_13909,N_12708);
and U15551 (N_15551,N_12266,N_12133);
or U15552 (N_15552,N_13959,N_13271);
and U15553 (N_15553,N_12060,N_12722);
nor U15554 (N_15554,N_12528,N_13954);
and U15555 (N_15555,N_13455,N_12772);
and U15556 (N_15556,N_13018,N_13483);
and U15557 (N_15557,N_12615,N_13576);
and U15558 (N_15558,N_12172,N_12999);
nand U15559 (N_15559,N_13807,N_13435);
nand U15560 (N_15560,N_12216,N_12637);
nand U15561 (N_15561,N_12979,N_13735);
nor U15562 (N_15562,N_12395,N_13870);
and U15563 (N_15563,N_12704,N_13307);
nand U15564 (N_15564,N_12785,N_13775);
or U15565 (N_15565,N_13506,N_13676);
nand U15566 (N_15566,N_13136,N_12272);
and U15567 (N_15567,N_13825,N_12535);
nand U15568 (N_15568,N_12430,N_12113);
nor U15569 (N_15569,N_12889,N_12006);
xnor U15570 (N_15570,N_13614,N_12337);
and U15571 (N_15571,N_12873,N_13573);
nand U15572 (N_15572,N_12899,N_13974);
and U15573 (N_15573,N_13860,N_13057);
nand U15574 (N_15574,N_12021,N_12556);
or U15575 (N_15575,N_13851,N_12430);
or U15576 (N_15576,N_12307,N_13149);
or U15577 (N_15577,N_13479,N_13925);
nor U15578 (N_15578,N_12084,N_13575);
or U15579 (N_15579,N_12333,N_12855);
nor U15580 (N_15580,N_13030,N_12914);
and U15581 (N_15581,N_12640,N_13245);
or U15582 (N_15582,N_12587,N_13299);
nor U15583 (N_15583,N_12618,N_13464);
xnor U15584 (N_15584,N_12704,N_12844);
nand U15585 (N_15585,N_13338,N_13322);
and U15586 (N_15586,N_13145,N_12510);
nand U15587 (N_15587,N_13952,N_12295);
nor U15588 (N_15588,N_12166,N_13434);
nor U15589 (N_15589,N_12219,N_13059);
or U15590 (N_15590,N_13149,N_13599);
nand U15591 (N_15591,N_12642,N_12938);
and U15592 (N_15592,N_12302,N_12205);
nor U15593 (N_15593,N_13070,N_12108);
and U15594 (N_15594,N_13693,N_12901);
nand U15595 (N_15595,N_12992,N_13756);
and U15596 (N_15596,N_13968,N_13092);
and U15597 (N_15597,N_13078,N_13269);
nor U15598 (N_15598,N_12238,N_13224);
nand U15599 (N_15599,N_12432,N_12108);
and U15600 (N_15600,N_12728,N_13797);
and U15601 (N_15601,N_13250,N_13941);
and U15602 (N_15602,N_12559,N_12302);
nand U15603 (N_15603,N_13411,N_13845);
nor U15604 (N_15604,N_13752,N_13385);
xnor U15605 (N_15605,N_13264,N_12589);
and U15606 (N_15606,N_13351,N_12988);
or U15607 (N_15607,N_12254,N_13143);
or U15608 (N_15608,N_13699,N_13773);
nand U15609 (N_15609,N_12088,N_13848);
and U15610 (N_15610,N_12108,N_12270);
and U15611 (N_15611,N_13888,N_13448);
and U15612 (N_15612,N_12814,N_13932);
nor U15613 (N_15613,N_13573,N_12063);
nor U15614 (N_15614,N_12588,N_12597);
xnor U15615 (N_15615,N_12513,N_12809);
nand U15616 (N_15616,N_12918,N_12778);
xnor U15617 (N_15617,N_12538,N_12047);
or U15618 (N_15618,N_13459,N_13634);
nor U15619 (N_15619,N_13436,N_12391);
and U15620 (N_15620,N_13579,N_13451);
and U15621 (N_15621,N_13788,N_13115);
or U15622 (N_15622,N_13562,N_12211);
or U15623 (N_15623,N_13971,N_12634);
and U15624 (N_15624,N_12420,N_13250);
xor U15625 (N_15625,N_13796,N_12612);
or U15626 (N_15626,N_12470,N_13853);
or U15627 (N_15627,N_12184,N_12240);
or U15628 (N_15628,N_13891,N_13624);
or U15629 (N_15629,N_13758,N_12763);
nand U15630 (N_15630,N_13054,N_12207);
nor U15631 (N_15631,N_12035,N_12375);
and U15632 (N_15632,N_13192,N_12049);
nor U15633 (N_15633,N_12507,N_12503);
or U15634 (N_15634,N_12929,N_12873);
xor U15635 (N_15635,N_12054,N_12435);
or U15636 (N_15636,N_12463,N_13384);
and U15637 (N_15637,N_12060,N_12480);
or U15638 (N_15638,N_13396,N_13694);
and U15639 (N_15639,N_13947,N_13121);
and U15640 (N_15640,N_13069,N_12220);
nor U15641 (N_15641,N_13993,N_12149);
nand U15642 (N_15642,N_12365,N_13100);
and U15643 (N_15643,N_13261,N_13598);
nor U15644 (N_15644,N_13454,N_13790);
nor U15645 (N_15645,N_12361,N_12691);
nor U15646 (N_15646,N_13315,N_13556);
nand U15647 (N_15647,N_13149,N_13452);
xnor U15648 (N_15648,N_12366,N_12318);
nor U15649 (N_15649,N_12074,N_13363);
xnor U15650 (N_15650,N_13422,N_13115);
and U15651 (N_15651,N_12883,N_12007);
or U15652 (N_15652,N_13418,N_12851);
xor U15653 (N_15653,N_12778,N_12196);
or U15654 (N_15654,N_12022,N_13658);
xnor U15655 (N_15655,N_12274,N_12081);
or U15656 (N_15656,N_13858,N_12428);
or U15657 (N_15657,N_12713,N_13763);
or U15658 (N_15658,N_13562,N_12521);
or U15659 (N_15659,N_13600,N_12214);
nand U15660 (N_15660,N_13759,N_13279);
and U15661 (N_15661,N_12537,N_12067);
nor U15662 (N_15662,N_13340,N_13726);
nand U15663 (N_15663,N_13337,N_13585);
or U15664 (N_15664,N_12230,N_13544);
nand U15665 (N_15665,N_13031,N_12824);
and U15666 (N_15666,N_12273,N_13472);
nor U15667 (N_15667,N_13996,N_13123);
nand U15668 (N_15668,N_13680,N_12304);
nand U15669 (N_15669,N_13411,N_12617);
and U15670 (N_15670,N_13146,N_12426);
nand U15671 (N_15671,N_12838,N_12404);
xor U15672 (N_15672,N_13985,N_13296);
nand U15673 (N_15673,N_13795,N_13229);
or U15674 (N_15674,N_12444,N_12654);
nor U15675 (N_15675,N_13179,N_12275);
and U15676 (N_15676,N_12914,N_13810);
nor U15677 (N_15677,N_13724,N_13854);
or U15678 (N_15678,N_12827,N_12717);
nand U15679 (N_15679,N_12061,N_13507);
and U15680 (N_15680,N_12448,N_13259);
nand U15681 (N_15681,N_12746,N_12120);
nor U15682 (N_15682,N_12221,N_13466);
nand U15683 (N_15683,N_12432,N_12588);
nor U15684 (N_15684,N_13206,N_13098);
and U15685 (N_15685,N_12074,N_12719);
and U15686 (N_15686,N_13562,N_13823);
or U15687 (N_15687,N_12974,N_13635);
nand U15688 (N_15688,N_13720,N_12406);
nor U15689 (N_15689,N_13257,N_12728);
and U15690 (N_15690,N_12206,N_12127);
or U15691 (N_15691,N_12689,N_13025);
and U15692 (N_15692,N_12314,N_12680);
or U15693 (N_15693,N_12603,N_12261);
and U15694 (N_15694,N_13604,N_13053);
nor U15695 (N_15695,N_12786,N_12110);
nor U15696 (N_15696,N_12227,N_12627);
nand U15697 (N_15697,N_13387,N_12578);
or U15698 (N_15698,N_13377,N_12431);
nor U15699 (N_15699,N_13949,N_12226);
nand U15700 (N_15700,N_12629,N_13409);
nor U15701 (N_15701,N_12498,N_12943);
nor U15702 (N_15702,N_12993,N_13819);
and U15703 (N_15703,N_12044,N_13217);
xor U15704 (N_15704,N_13653,N_12562);
and U15705 (N_15705,N_12385,N_12868);
nor U15706 (N_15706,N_12557,N_12363);
and U15707 (N_15707,N_13961,N_12356);
xnor U15708 (N_15708,N_13892,N_12504);
nor U15709 (N_15709,N_12465,N_12232);
and U15710 (N_15710,N_13535,N_12920);
and U15711 (N_15711,N_13560,N_12162);
nor U15712 (N_15712,N_13930,N_12375);
or U15713 (N_15713,N_13916,N_12749);
xnor U15714 (N_15714,N_13453,N_12083);
or U15715 (N_15715,N_13792,N_13061);
or U15716 (N_15716,N_12856,N_13879);
or U15717 (N_15717,N_12678,N_12780);
and U15718 (N_15718,N_12697,N_12297);
and U15719 (N_15719,N_12125,N_13398);
nand U15720 (N_15720,N_12293,N_13481);
nand U15721 (N_15721,N_13996,N_12104);
nand U15722 (N_15722,N_13201,N_13016);
and U15723 (N_15723,N_12055,N_12320);
nor U15724 (N_15724,N_13684,N_13214);
nor U15725 (N_15725,N_12821,N_13149);
and U15726 (N_15726,N_12626,N_13817);
nor U15727 (N_15727,N_13860,N_12042);
xnor U15728 (N_15728,N_13747,N_13807);
nand U15729 (N_15729,N_13245,N_13070);
nor U15730 (N_15730,N_12717,N_13043);
xor U15731 (N_15731,N_12961,N_12372);
and U15732 (N_15732,N_13855,N_13693);
xor U15733 (N_15733,N_13245,N_12532);
nand U15734 (N_15734,N_13047,N_13662);
and U15735 (N_15735,N_13205,N_12162);
nor U15736 (N_15736,N_13686,N_13144);
nand U15737 (N_15737,N_12230,N_12463);
nand U15738 (N_15738,N_13371,N_13589);
nor U15739 (N_15739,N_13079,N_12618);
nand U15740 (N_15740,N_13618,N_12238);
and U15741 (N_15741,N_13271,N_12313);
and U15742 (N_15742,N_12602,N_13332);
xor U15743 (N_15743,N_12811,N_12520);
nand U15744 (N_15744,N_12725,N_13242);
xor U15745 (N_15745,N_12532,N_12515);
xor U15746 (N_15746,N_12370,N_13284);
and U15747 (N_15747,N_12347,N_12492);
nand U15748 (N_15748,N_12144,N_12686);
and U15749 (N_15749,N_13519,N_12734);
and U15750 (N_15750,N_13416,N_13694);
nand U15751 (N_15751,N_13694,N_12544);
nand U15752 (N_15752,N_12661,N_13092);
nor U15753 (N_15753,N_12130,N_12853);
and U15754 (N_15754,N_13767,N_12320);
nor U15755 (N_15755,N_13680,N_12515);
nor U15756 (N_15756,N_12286,N_13121);
and U15757 (N_15757,N_13449,N_13037);
or U15758 (N_15758,N_13331,N_12446);
or U15759 (N_15759,N_13437,N_13167);
and U15760 (N_15760,N_12835,N_13488);
nor U15761 (N_15761,N_13280,N_12104);
nand U15762 (N_15762,N_12717,N_12214);
nand U15763 (N_15763,N_12864,N_12265);
nand U15764 (N_15764,N_13692,N_13740);
nand U15765 (N_15765,N_13432,N_12001);
nand U15766 (N_15766,N_12012,N_12969);
nor U15767 (N_15767,N_12890,N_12114);
and U15768 (N_15768,N_12459,N_12927);
and U15769 (N_15769,N_12014,N_12119);
nand U15770 (N_15770,N_13526,N_12672);
xnor U15771 (N_15771,N_12846,N_13978);
nand U15772 (N_15772,N_13939,N_12354);
nand U15773 (N_15773,N_12118,N_12673);
and U15774 (N_15774,N_13025,N_13425);
xnor U15775 (N_15775,N_13493,N_12593);
nor U15776 (N_15776,N_12182,N_13673);
xnor U15777 (N_15777,N_13673,N_13098);
and U15778 (N_15778,N_12024,N_13186);
and U15779 (N_15779,N_12929,N_12498);
nand U15780 (N_15780,N_12529,N_13360);
nor U15781 (N_15781,N_13949,N_13070);
and U15782 (N_15782,N_12026,N_13904);
nand U15783 (N_15783,N_13539,N_13093);
nand U15784 (N_15784,N_12128,N_13218);
nor U15785 (N_15785,N_13414,N_12831);
and U15786 (N_15786,N_13379,N_13088);
and U15787 (N_15787,N_12827,N_13721);
nor U15788 (N_15788,N_12364,N_12643);
nor U15789 (N_15789,N_12808,N_12290);
xnor U15790 (N_15790,N_13168,N_13617);
nand U15791 (N_15791,N_12691,N_13075);
nor U15792 (N_15792,N_12784,N_12855);
xor U15793 (N_15793,N_12838,N_12052);
nor U15794 (N_15794,N_13999,N_13892);
nor U15795 (N_15795,N_13627,N_13389);
xor U15796 (N_15796,N_12448,N_13417);
xor U15797 (N_15797,N_13922,N_13543);
xor U15798 (N_15798,N_13912,N_13766);
xor U15799 (N_15799,N_12351,N_13839);
nor U15800 (N_15800,N_12581,N_13872);
xor U15801 (N_15801,N_13259,N_13628);
and U15802 (N_15802,N_13796,N_13660);
and U15803 (N_15803,N_13612,N_12874);
and U15804 (N_15804,N_12905,N_12362);
or U15805 (N_15805,N_13831,N_12892);
or U15806 (N_15806,N_13469,N_13737);
xnor U15807 (N_15807,N_12130,N_12180);
or U15808 (N_15808,N_13646,N_12495);
nor U15809 (N_15809,N_13491,N_13220);
nand U15810 (N_15810,N_12863,N_13139);
or U15811 (N_15811,N_13206,N_12972);
xnor U15812 (N_15812,N_13096,N_13014);
or U15813 (N_15813,N_12234,N_13262);
xor U15814 (N_15814,N_12313,N_13296);
or U15815 (N_15815,N_12843,N_12419);
and U15816 (N_15816,N_12790,N_12504);
nand U15817 (N_15817,N_12355,N_12740);
or U15818 (N_15818,N_13096,N_13010);
nor U15819 (N_15819,N_12465,N_13931);
or U15820 (N_15820,N_13239,N_12757);
nand U15821 (N_15821,N_13555,N_12328);
and U15822 (N_15822,N_13912,N_12367);
and U15823 (N_15823,N_12615,N_12929);
xnor U15824 (N_15824,N_12069,N_12624);
nand U15825 (N_15825,N_12764,N_12127);
nor U15826 (N_15826,N_13762,N_13328);
or U15827 (N_15827,N_13808,N_13238);
nor U15828 (N_15828,N_12459,N_13520);
and U15829 (N_15829,N_13516,N_12556);
and U15830 (N_15830,N_13642,N_12811);
nor U15831 (N_15831,N_12850,N_13417);
nand U15832 (N_15832,N_12362,N_13305);
nand U15833 (N_15833,N_12978,N_12508);
and U15834 (N_15834,N_13818,N_12281);
and U15835 (N_15835,N_13283,N_12001);
nor U15836 (N_15836,N_12689,N_13266);
or U15837 (N_15837,N_12569,N_12375);
and U15838 (N_15838,N_13051,N_12863);
and U15839 (N_15839,N_13952,N_12928);
xnor U15840 (N_15840,N_13002,N_12320);
or U15841 (N_15841,N_13663,N_13046);
or U15842 (N_15842,N_12433,N_13744);
and U15843 (N_15843,N_13954,N_13408);
nor U15844 (N_15844,N_12771,N_12648);
and U15845 (N_15845,N_12610,N_13765);
and U15846 (N_15846,N_12799,N_13375);
or U15847 (N_15847,N_13319,N_13989);
xnor U15848 (N_15848,N_13139,N_13866);
xor U15849 (N_15849,N_13354,N_13324);
nand U15850 (N_15850,N_13999,N_13028);
or U15851 (N_15851,N_12912,N_13013);
and U15852 (N_15852,N_12950,N_12356);
nand U15853 (N_15853,N_13835,N_13587);
nand U15854 (N_15854,N_12119,N_13288);
or U15855 (N_15855,N_13041,N_12630);
or U15856 (N_15856,N_12857,N_13284);
nor U15857 (N_15857,N_12935,N_13704);
xor U15858 (N_15858,N_12449,N_13431);
or U15859 (N_15859,N_12635,N_12800);
and U15860 (N_15860,N_12571,N_12915);
and U15861 (N_15861,N_12817,N_13360);
and U15862 (N_15862,N_13671,N_12597);
or U15863 (N_15863,N_13215,N_13163);
nor U15864 (N_15864,N_13107,N_13986);
nor U15865 (N_15865,N_13391,N_12285);
nor U15866 (N_15866,N_13879,N_12321);
or U15867 (N_15867,N_12314,N_13161);
nand U15868 (N_15868,N_13548,N_12834);
and U15869 (N_15869,N_13627,N_13538);
nor U15870 (N_15870,N_12694,N_12541);
nor U15871 (N_15871,N_13748,N_12232);
and U15872 (N_15872,N_13190,N_12084);
or U15873 (N_15873,N_12107,N_13508);
nor U15874 (N_15874,N_13925,N_12022);
nand U15875 (N_15875,N_12092,N_12302);
nor U15876 (N_15876,N_12414,N_13078);
nand U15877 (N_15877,N_12340,N_13725);
or U15878 (N_15878,N_13621,N_12112);
nor U15879 (N_15879,N_12081,N_12659);
and U15880 (N_15880,N_12935,N_12860);
and U15881 (N_15881,N_13201,N_12535);
and U15882 (N_15882,N_13415,N_13322);
and U15883 (N_15883,N_12100,N_13072);
nor U15884 (N_15884,N_13351,N_12479);
or U15885 (N_15885,N_13057,N_13647);
xor U15886 (N_15886,N_13907,N_12215);
nand U15887 (N_15887,N_12147,N_13018);
nand U15888 (N_15888,N_13389,N_12527);
nand U15889 (N_15889,N_12673,N_12871);
and U15890 (N_15890,N_12489,N_12620);
xnor U15891 (N_15891,N_12437,N_13919);
nand U15892 (N_15892,N_13684,N_13529);
and U15893 (N_15893,N_13578,N_13388);
or U15894 (N_15894,N_13992,N_13067);
and U15895 (N_15895,N_13958,N_13136);
nand U15896 (N_15896,N_13740,N_12232);
nor U15897 (N_15897,N_12015,N_12782);
nor U15898 (N_15898,N_13520,N_12853);
and U15899 (N_15899,N_12114,N_12281);
nand U15900 (N_15900,N_12090,N_13561);
nor U15901 (N_15901,N_12466,N_12794);
nor U15902 (N_15902,N_12770,N_13550);
nor U15903 (N_15903,N_12857,N_12314);
or U15904 (N_15904,N_12759,N_13535);
or U15905 (N_15905,N_12705,N_13533);
or U15906 (N_15906,N_13261,N_12652);
and U15907 (N_15907,N_12126,N_13316);
nand U15908 (N_15908,N_13977,N_12731);
nor U15909 (N_15909,N_13962,N_13784);
nand U15910 (N_15910,N_12871,N_12843);
or U15911 (N_15911,N_13309,N_13765);
and U15912 (N_15912,N_13471,N_12331);
nor U15913 (N_15913,N_12491,N_12341);
nor U15914 (N_15914,N_12838,N_13825);
xnor U15915 (N_15915,N_13419,N_12197);
and U15916 (N_15916,N_12510,N_13976);
and U15917 (N_15917,N_13808,N_13837);
nor U15918 (N_15918,N_12390,N_13385);
and U15919 (N_15919,N_13278,N_13213);
nor U15920 (N_15920,N_12433,N_13407);
nand U15921 (N_15921,N_12693,N_12191);
or U15922 (N_15922,N_12472,N_12921);
nand U15923 (N_15923,N_13201,N_12372);
nand U15924 (N_15924,N_12542,N_13889);
nand U15925 (N_15925,N_12361,N_12220);
and U15926 (N_15926,N_12633,N_12798);
or U15927 (N_15927,N_13542,N_13125);
nor U15928 (N_15928,N_12728,N_13785);
and U15929 (N_15929,N_12166,N_13199);
nand U15930 (N_15930,N_12781,N_12413);
or U15931 (N_15931,N_13921,N_12963);
nor U15932 (N_15932,N_12450,N_12400);
nand U15933 (N_15933,N_13157,N_12148);
or U15934 (N_15934,N_13052,N_12946);
xor U15935 (N_15935,N_13289,N_13380);
nand U15936 (N_15936,N_12240,N_12504);
and U15937 (N_15937,N_12352,N_13085);
or U15938 (N_15938,N_12410,N_12851);
nor U15939 (N_15939,N_13573,N_13083);
and U15940 (N_15940,N_12659,N_13221);
nor U15941 (N_15941,N_12843,N_13936);
nand U15942 (N_15942,N_12603,N_13610);
or U15943 (N_15943,N_12464,N_13641);
nand U15944 (N_15944,N_12364,N_13833);
or U15945 (N_15945,N_12936,N_13137);
and U15946 (N_15946,N_13510,N_12592);
nand U15947 (N_15947,N_13850,N_13300);
and U15948 (N_15948,N_12727,N_13768);
or U15949 (N_15949,N_13335,N_12951);
nand U15950 (N_15950,N_13855,N_13883);
nor U15951 (N_15951,N_13714,N_12298);
nand U15952 (N_15952,N_12430,N_13496);
nor U15953 (N_15953,N_13050,N_13722);
nor U15954 (N_15954,N_12629,N_12041);
and U15955 (N_15955,N_13930,N_13439);
or U15956 (N_15956,N_13762,N_13121);
or U15957 (N_15957,N_13544,N_12482);
nor U15958 (N_15958,N_12936,N_13686);
nor U15959 (N_15959,N_13685,N_13171);
and U15960 (N_15960,N_13835,N_13446);
and U15961 (N_15961,N_13386,N_12266);
xnor U15962 (N_15962,N_13647,N_12332);
xnor U15963 (N_15963,N_13173,N_13165);
nor U15964 (N_15964,N_12952,N_13022);
and U15965 (N_15965,N_12735,N_13647);
or U15966 (N_15966,N_13705,N_13779);
and U15967 (N_15967,N_12998,N_12612);
nor U15968 (N_15968,N_12201,N_13887);
or U15969 (N_15969,N_12946,N_12026);
nor U15970 (N_15970,N_13289,N_13483);
nor U15971 (N_15971,N_12700,N_13705);
or U15972 (N_15972,N_13017,N_12898);
xor U15973 (N_15973,N_13927,N_12602);
nor U15974 (N_15974,N_12389,N_13441);
nand U15975 (N_15975,N_12942,N_12695);
xor U15976 (N_15976,N_13398,N_13020);
and U15977 (N_15977,N_12417,N_13902);
nand U15978 (N_15978,N_13375,N_12019);
or U15979 (N_15979,N_12776,N_12389);
nor U15980 (N_15980,N_13193,N_13878);
nand U15981 (N_15981,N_13443,N_12473);
nor U15982 (N_15982,N_12608,N_12349);
nand U15983 (N_15983,N_12254,N_12854);
nand U15984 (N_15984,N_13432,N_13187);
or U15985 (N_15985,N_13633,N_12631);
and U15986 (N_15986,N_13133,N_13923);
nand U15987 (N_15987,N_12701,N_13714);
and U15988 (N_15988,N_12562,N_13069);
nor U15989 (N_15989,N_13922,N_12178);
nand U15990 (N_15990,N_13273,N_13290);
nor U15991 (N_15991,N_13543,N_12469);
xnor U15992 (N_15992,N_13310,N_13939);
nor U15993 (N_15993,N_12730,N_12339);
nand U15994 (N_15994,N_13091,N_13205);
or U15995 (N_15995,N_13900,N_12455);
nor U15996 (N_15996,N_13003,N_12671);
nor U15997 (N_15997,N_13324,N_12469);
or U15998 (N_15998,N_13634,N_13501);
xnor U15999 (N_15999,N_12636,N_13561);
nand U16000 (N_16000,N_14951,N_15296);
nor U16001 (N_16001,N_14509,N_14867);
nand U16002 (N_16002,N_14684,N_15874);
and U16003 (N_16003,N_14146,N_14644);
nor U16004 (N_16004,N_15125,N_14419);
nor U16005 (N_16005,N_15828,N_14504);
and U16006 (N_16006,N_14099,N_15587);
or U16007 (N_16007,N_14877,N_14861);
nand U16008 (N_16008,N_15080,N_14941);
nor U16009 (N_16009,N_15973,N_14107);
xnor U16010 (N_16010,N_15856,N_14091);
and U16011 (N_16011,N_15982,N_15954);
nand U16012 (N_16012,N_14387,N_15060);
nand U16013 (N_16013,N_15319,N_15946);
or U16014 (N_16014,N_15482,N_14349);
nor U16015 (N_16015,N_14222,N_14487);
nor U16016 (N_16016,N_14437,N_15112);
nor U16017 (N_16017,N_14599,N_14448);
xor U16018 (N_16018,N_15656,N_14417);
nand U16019 (N_16019,N_15998,N_14161);
nand U16020 (N_16020,N_15870,N_14042);
or U16021 (N_16021,N_15198,N_14870);
or U16022 (N_16022,N_14351,N_15688);
or U16023 (N_16023,N_14709,N_14949);
nand U16024 (N_16024,N_15417,N_14239);
and U16025 (N_16025,N_14163,N_14992);
nor U16026 (N_16026,N_14835,N_15880);
nor U16027 (N_16027,N_15333,N_14059);
or U16028 (N_16028,N_15097,N_15464);
nor U16029 (N_16029,N_14589,N_14791);
xor U16030 (N_16030,N_14399,N_15472);
nor U16031 (N_16031,N_14762,N_14392);
or U16032 (N_16032,N_15021,N_15837);
nor U16033 (N_16033,N_14343,N_14982);
nor U16034 (N_16034,N_14680,N_14070);
xnor U16035 (N_16035,N_14544,N_15193);
nand U16036 (N_16036,N_14041,N_15813);
nand U16037 (N_16037,N_15226,N_14449);
or U16038 (N_16038,N_15903,N_14014);
xnor U16039 (N_16039,N_15768,N_15832);
nand U16040 (N_16040,N_15011,N_15612);
or U16041 (N_16041,N_14893,N_14501);
and U16042 (N_16042,N_15326,N_14192);
xor U16043 (N_16043,N_14388,N_14431);
or U16044 (N_16044,N_15222,N_15732);
nand U16045 (N_16045,N_14434,N_15788);
xor U16046 (N_16046,N_15879,N_14816);
nor U16047 (N_16047,N_14965,N_15552);
nand U16048 (N_16048,N_15944,N_15019);
xnor U16049 (N_16049,N_15001,N_14275);
or U16050 (N_16050,N_15098,N_14821);
nand U16051 (N_16051,N_14984,N_14196);
or U16052 (N_16052,N_14190,N_15167);
or U16053 (N_16053,N_14715,N_14324);
nand U16054 (N_16054,N_14790,N_15206);
or U16055 (N_16055,N_15943,N_14697);
or U16056 (N_16056,N_14944,N_15983);
and U16057 (N_16057,N_15245,N_15002);
xnor U16058 (N_16058,N_15966,N_15711);
xor U16059 (N_16059,N_15137,N_15811);
nand U16060 (N_16060,N_14083,N_15975);
and U16061 (N_16061,N_14360,N_14722);
nor U16062 (N_16062,N_15479,N_14495);
nand U16063 (N_16063,N_14172,N_14649);
and U16064 (N_16064,N_14040,N_15241);
nand U16065 (N_16065,N_14223,N_15093);
and U16066 (N_16066,N_14592,N_14761);
nor U16067 (N_16067,N_15704,N_15558);
and U16068 (N_16068,N_15530,N_15260);
and U16069 (N_16069,N_14545,N_14229);
nand U16070 (N_16070,N_14553,N_15175);
nand U16071 (N_16071,N_14466,N_15580);
and U16072 (N_16072,N_15276,N_15505);
nor U16073 (N_16073,N_14962,N_15481);
nor U16074 (N_16074,N_14654,N_14114);
or U16075 (N_16075,N_14998,N_14297);
xor U16076 (N_16076,N_14942,N_15706);
or U16077 (N_16077,N_14159,N_14887);
or U16078 (N_16078,N_14116,N_14754);
nand U16079 (N_16079,N_15030,N_15070);
or U16080 (N_16080,N_14674,N_15212);
or U16081 (N_16081,N_14374,N_14533);
and U16082 (N_16082,N_14935,N_14338);
or U16083 (N_16083,N_15191,N_14988);
nand U16084 (N_16084,N_15473,N_14915);
xor U16085 (N_16085,N_15765,N_15275);
nand U16086 (N_16086,N_15540,N_15246);
nand U16087 (N_16087,N_14145,N_14376);
nor U16088 (N_16088,N_15985,N_15224);
nor U16089 (N_16089,N_15781,N_14102);
or U16090 (N_16090,N_14327,N_14752);
and U16091 (N_16091,N_15757,N_15715);
or U16092 (N_16092,N_15795,N_15027);
or U16093 (N_16093,N_14357,N_15763);
xor U16094 (N_16094,N_15234,N_14566);
nor U16095 (N_16095,N_15786,N_15075);
or U16096 (N_16096,N_14314,N_15589);
and U16097 (N_16097,N_14142,N_14403);
or U16098 (N_16098,N_14595,N_15869);
and U16099 (N_16099,N_15186,N_14226);
and U16100 (N_16100,N_14587,N_14727);
nor U16101 (N_16101,N_15452,N_14945);
or U16102 (N_16102,N_14299,N_15357);
or U16103 (N_16103,N_14272,N_14414);
or U16104 (N_16104,N_15350,N_14305);
or U16105 (N_16105,N_15769,N_14350);
nand U16106 (N_16106,N_15114,N_14927);
nand U16107 (N_16107,N_15690,N_15082);
xor U16108 (N_16108,N_14095,N_15913);
or U16109 (N_16109,N_14999,N_15121);
nor U16110 (N_16110,N_14515,N_14796);
nor U16111 (N_16111,N_15861,N_15057);
nand U16112 (N_16112,N_15359,N_14651);
and U16113 (N_16113,N_15631,N_15753);
nor U16114 (N_16114,N_15285,N_14681);
or U16115 (N_16115,N_15852,N_14892);
and U16116 (N_16116,N_14691,N_15407);
and U16117 (N_16117,N_14078,N_14108);
nor U16118 (N_16118,N_14735,N_15513);
nor U16119 (N_16119,N_15272,N_15981);
or U16120 (N_16120,N_15734,N_14720);
xnor U16121 (N_16121,N_15658,N_15192);
nand U16122 (N_16122,N_14373,N_15637);
and U16123 (N_16123,N_15923,N_14631);
nor U16124 (N_16124,N_14391,N_15709);
or U16125 (N_16125,N_15375,N_14215);
or U16126 (N_16126,N_15997,N_14265);
nand U16127 (N_16127,N_15814,N_14841);
xnor U16128 (N_16128,N_14243,N_14492);
or U16129 (N_16129,N_15664,N_15238);
nand U16130 (N_16130,N_14885,N_15782);
nor U16131 (N_16131,N_15267,N_15091);
nor U16132 (N_16132,N_14217,N_15079);
nand U16133 (N_16133,N_15504,N_15979);
or U16134 (N_16134,N_14189,N_14436);
nand U16135 (N_16135,N_15610,N_14795);
nand U16136 (N_16136,N_15428,N_14639);
or U16137 (N_16137,N_15697,N_15099);
or U16138 (N_16138,N_15563,N_14986);
nor U16139 (N_16139,N_14187,N_14817);
or U16140 (N_16140,N_14706,N_14894);
or U16141 (N_16141,N_14415,N_15162);
or U16142 (N_16142,N_15169,N_14692);
or U16143 (N_16143,N_15687,N_14936);
xnor U16144 (N_16144,N_14136,N_14932);
nand U16145 (N_16145,N_15933,N_14689);
nor U16146 (N_16146,N_15032,N_14728);
or U16147 (N_16147,N_14925,N_15957);
nand U16148 (N_16148,N_15144,N_14057);
nand U16149 (N_16149,N_14268,N_14862);
or U16150 (N_16150,N_14626,N_14581);
nor U16151 (N_16151,N_14276,N_15755);
nand U16152 (N_16152,N_15300,N_15083);
nand U16153 (N_16153,N_15659,N_15559);
or U16154 (N_16154,N_14247,N_14315);
nor U16155 (N_16155,N_14552,N_14288);
and U16156 (N_16156,N_15767,N_14777);
nor U16157 (N_16157,N_14718,N_15055);
or U16158 (N_16158,N_15003,N_14298);
nand U16159 (N_16159,N_15416,N_15415);
or U16160 (N_16160,N_15301,N_14921);
and U16161 (N_16161,N_14560,N_14645);
and U16162 (N_16162,N_15387,N_15088);
or U16163 (N_16163,N_14179,N_15063);
or U16164 (N_16164,N_15199,N_14522);
or U16165 (N_16165,N_15705,N_15834);
xnor U16166 (N_16166,N_15372,N_14123);
nor U16167 (N_16167,N_15293,N_14402);
nand U16168 (N_16168,N_15466,N_15672);
nand U16169 (N_16169,N_15833,N_15851);
nor U16170 (N_16170,N_15108,N_15758);
nand U16171 (N_16171,N_15178,N_15335);
and U16172 (N_16172,N_15130,N_14975);
nand U16173 (N_16173,N_15243,N_15330);
or U16174 (N_16174,N_14696,N_14055);
nor U16175 (N_16175,N_15527,N_15255);
or U16176 (N_16176,N_15392,N_14044);
xnor U16177 (N_16177,N_15752,N_14046);
nand U16178 (N_16178,N_14331,N_14489);
or U16179 (N_16179,N_14130,N_14705);
nand U16180 (N_16180,N_14908,N_14667);
and U16181 (N_16181,N_15277,N_15219);
nor U16182 (N_16182,N_15320,N_14236);
nor U16183 (N_16183,N_14439,N_15528);
or U16184 (N_16184,N_15262,N_14904);
nor U16185 (N_16185,N_15645,N_14588);
and U16186 (N_16186,N_15666,N_15179);
nor U16187 (N_16187,N_15622,N_15430);
xnor U16188 (N_16188,N_14913,N_14269);
and U16189 (N_16189,N_15521,N_14928);
or U16190 (N_16190,N_14097,N_14620);
or U16191 (N_16191,N_15154,N_14124);
or U16192 (N_16192,N_14428,N_14424);
or U16193 (N_16193,N_15056,N_14005);
nand U16194 (N_16194,N_15052,N_15764);
or U16195 (N_16195,N_15196,N_14548);
nand U16196 (N_16196,N_15756,N_14623);
nand U16197 (N_16197,N_15737,N_15936);
nor U16198 (N_16198,N_14201,N_15433);
or U16199 (N_16199,N_15013,N_15595);
and U16200 (N_16200,N_15994,N_15693);
nand U16201 (N_16201,N_15691,N_15218);
and U16202 (N_16202,N_15050,N_15887);
nand U16203 (N_16203,N_15584,N_15515);
or U16204 (N_16204,N_14410,N_14191);
and U16205 (N_16205,N_14611,N_14122);
nand U16206 (N_16206,N_14979,N_14568);
or U16207 (N_16207,N_14693,N_14937);
and U16208 (N_16208,N_15292,N_14829);
and U16209 (N_16209,N_15860,N_15022);
and U16210 (N_16210,N_15567,N_15976);
or U16211 (N_16211,N_14567,N_14039);
and U16212 (N_16212,N_15878,N_14084);
xnor U16213 (N_16213,N_15233,N_14868);
nor U16214 (N_16214,N_15723,N_15081);
nor U16215 (N_16215,N_14408,N_14759);
nor U16216 (N_16216,N_14372,N_15522);
nor U16217 (N_16217,N_15462,N_15486);
nor U16218 (N_16218,N_15639,N_15247);
nand U16219 (N_16219,N_14633,N_14764);
nor U16220 (N_16220,N_15331,N_14612);
nand U16221 (N_16221,N_15534,N_14686);
nor U16222 (N_16222,N_14524,N_14105);
or U16223 (N_16223,N_14300,N_14571);
or U16224 (N_16224,N_15801,N_14469);
nor U16225 (N_16225,N_14855,N_14966);
nand U16226 (N_16226,N_14255,N_14820);
or U16227 (N_16227,N_15015,N_15653);
or U16228 (N_16228,N_14637,N_15404);
or U16229 (N_16229,N_14648,N_14144);
or U16230 (N_16230,N_14362,N_14241);
or U16231 (N_16231,N_15498,N_15256);
nand U16232 (N_16232,N_15037,N_15143);
or U16233 (N_16233,N_15731,N_15648);
nand U16234 (N_16234,N_14446,N_14429);
or U16235 (N_16235,N_14530,N_14094);
nor U16236 (N_16236,N_14453,N_15745);
or U16237 (N_16237,N_15394,N_15902);
nand U16238 (N_16238,N_14394,N_15471);
nand U16239 (N_16239,N_15306,N_14657);
and U16240 (N_16240,N_15549,N_15204);
nor U16241 (N_16241,N_14580,N_14760);
nor U16242 (N_16242,N_14412,N_14157);
nor U16243 (N_16243,N_15924,N_15626);
and U16244 (N_16244,N_14682,N_15971);
xor U16245 (N_16245,N_15122,N_14493);
xor U16246 (N_16246,N_15872,N_15545);
nand U16247 (N_16247,N_14987,N_15237);
nor U16248 (N_16248,N_14656,N_15646);
nor U16249 (N_16249,N_14807,N_14874);
and U16250 (N_16250,N_14200,N_14563);
nor U16251 (N_16251,N_14433,N_14521);
nand U16252 (N_16252,N_15673,N_15823);
or U16253 (N_16253,N_14475,N_15474);
nor U16254 (N_16254,N_14038,N_14404);
nor U16255 (N_16255,N_14801,N_15842);
nand U16256 (N_16256,N_14658,N_15604);
nand U16257 (N_16257,N_15980,N_14371);
nand U16258 (N_16258,N_15850,N_15820);
nor U16259 (N_16259,N_14216,N_15215);
nor U16260 (N_16260,N_15889,N_14342);
nor U16261 (N_16261,N_15235,N_15332);
nand U16262 (N_16262,N_14134,N_14677);
nor U16263 (N_16263,N_15628,N_15992);
xnor U16264 (N_16264,N_15607,N_14505);
and U16265 (N_16265,N_15524,N_15111);
and U16266 (N_16266,N_14220,N_14248);
nor U16267 (N_16267,N_15602,N_14880);
and U16268 (N_16268,N_15354,N_14073);
nor U16269 (N_16269,N_14930,N_15347);
nor U16270 (N_16270,N_15286,N_15397);
nand U16271 (N_16271,N_15592,N_15597);
nor U16272 (N_16272,N_14920,N_14481);
or U16273 (N_16273,N_15195,N_14670);
and U16274 (N_16274,N_15507,N_15855);
and U16275 (N_16275,N_14398,N_14729);
or U16276 (N_16276,N_15438,N_14018);
or U16277 (N_16277,N_14012,N_14939);
or U16278 (N_16278,N_15366,N_15085);
nor U16279 (N_16279,N_14529,N_14717);
and U16280 (N_16280,N_15259,N_15271);
nand U16281 (N_16281,N_14721,N_14339);
nor U16282 (N_16282,N_15411,N_15819);
and U16283 (N_16283,N_15974,N_15023);
nand U16284 (N_16284,N_15362,N_15046);
nor U16285 (N_16285,N_15551,N_14701);
nand U16286 (N_16286,N_15644,N_14284);
or U16287 (N_16287,N_14176,N_14174);
and U16288 (N_16288,N_14775,N_15240);
or U16289 (N_16289,N_15211,N_15594);
nor U16290 (N_16290,N_14502,N_15965);
nand U16291 (N_16291,N_15383,N_15729);
nor U16292 (N_16292,N_15989,N_15173);
xor U16293 (N_16293,N_15773,N_14411);
nand U16294 (N_16294,N_15952,N_14698);
xnor U16295 (N_16295,N_15155,N_14778);
nand U16296 (N_16296,N_15996,N_14496);
and U16297 (N_16297,N_15270,N_15437);
nand U16298 (N_16298,N_14451,N_15217);
and U16299 (N_16299,N_14053,N_14918);
and U16300 (N_16300,N_14112,N_15053);
or U16301 (N_16301,N_15294,N_14167);
nand U16302 (N_16302,N_15264,N_15562);
and U16303 (N_16303,N_14212,N_14066);
or U16304 (N_16304,N_15156,N_14900);
and U16305 (N_16305,N_14557,N_14271);
nor U16306 (N_16306,N_14379,N_14249);
xor U16307 (N_16307,N_14559,N_15713);
nor U16308 (N_16308,N_14508,N_14789);
and U16309 (N_16309,N_14295,N_15868);
and U16310 (N_16310,N_14177,N_14856);
nand U16311 (N_16311,N_15410,N_14614);
or U16312 (N_16312,N_15386,N_15113);
nand U16313 (N_16313,N_15864,N_14234);
and U16314 (N_16314,N_14723,N_14804);
and U16315 (N_16315,N_15477,N_14185);
nand U16316 (N_16316,N_14832,N_15789);
or U16317 (N_16317,N_15058,N_15857);
nor U16318 (N_16318,N_14008,N_14209);
nand U16319 (N_16319,N_14699,N_14384);
or U16320 (N_16320,N_14093,N_14825);
or U16321 (N_16321,N_14903,N_15905);
and U16322 (N_16322,N_14155,N_14554);
nor U16323 (N_16323,N_14938,N_14990);
nor U16324 (N_16324,N_14213,N_14895);
nor U16325 (N_16325,N_14369,N_15461);
and U16326 (N_16326,N_14527,N_14964);
xor U16327 (N_16327,N_15345,N_15726);
nand U16328 (N_16328,N_15883,N_15812);
nor U16329 (N_16329,N_15546,N_15636);
nor U16330 (N_16330,N_14126,N_15858);
nor U16331 (N_16331,N_15741,N_15184);
and U16332 (N_16332,N_14457,N_14098);
nand U16333 (N_16333,N_14258,N_15710);
and U16334 (N_16334,N_15496,N_15408);
or U16335 (N_16335,N_14011,N_15554);
nor U16336 (N_16336,N_15051,N_15048);
or U16337 (N_16337,N_14273,N_15574);
or U16338 (N_16338,N_15614,N_15341);
and U16339 (N_16339,N_14477,N_14814);
and U16340 (N_16340,N_14584,N_14075);
or U16341 (N_16341,N_15748,N_15624);
or U16342 (N_16342,N_14793,N_14772);
xor U16343 (N_16343,N_14875,N_15892);
and U16344 (N_16344,N_15373,N_14025);
nor U16345 (N_16345,N_15134,N_15401);
xor U16346 (N_16346,N_15389,N_15844);
and U16347 (N_16347,N_14923,N_14463);
nor U16348 (N_16348,N_15356,N_15999);
and U16349 (N_16349,N_14266,N_14837);
and U16350 (N_16350,N_14341,N_14556);
and U16351 (N_16351,N_14438,N_14077);
or U16352 (N_16352,N_14732,N_14911);
nor U16353 (N_16353,N_14251,N_14238);
and U16354 (N_16354,N_14652,N_15958);
nand U16355 (N_16355,N_14850,N_14943);
nand U16356 (N_16356,N_15824,N_14204);
or U16357 (N_16357,N_14321,N_14395);
or U16358 (N_16358,N_14983,N_14052);
or U16359 (N_16359,N_14643,N_15579);
nor U16360 (N_16360,N_14051,N_14323);
nor U16361 (N_16361,N_14100,N_14565);
nand U16362 (N_16362,N_14886,N_14954);
nor U16363 (N_16363,N_14293,N_15603);
and U16364 (N_16364,N_15995,N_15570);
or U16365 (N_16365,N_14488,N_15086);
or U16366 (N_16366,N_15251,N_15714);
nand U16367 (N_16367,N_14193,N_14037);
nor U16368 (N_16368,N_14061,N_14365);
or U16369 (N_16369,N_14002,N_14573);
or U16370 (N_16370,N_14017,N_14188);
and U16371 (N_16371,N_15336,N_15109);
nand U16372 (N_16372,N_14719,N_15329);
xnor U16373 (N_16373,N_15412,N_15470);
or U16374 (N_16374,N_14186,N_14104);
nor U16375 (N_16375,N_14838,N_14842);
and U16376 (N_16376,N_14541,N_15266);
or U16377 (N_16377,N_14879,N_15573);
or U16378 (N_16378,N_14198,N_14304);
and U16379 (N_16379,N_14967,N_15564);
nor U16380 (N_16380,N_15059,N_14004);
nor U16381 (N_16381,N_14278,N_14844);
or U16382 (N_16382,N_15848,N_15586);
and U16383 (N_16383,N_14259,N_15572);
or U16384 (N_16384,N_15951,N_15232);
or U16385 (N_16385,N_15516,N_15681);
or U16386 (N_16386,N_14767,N_15065);
nor U16387 (N_16387,N_15476,N_15956);
xor U16388 (N_16388,N_15725,N_15601);
or U16389 (N_16389,N_14497,N_15761);
nand U16390 (N_16390,N_15771,N_14934);
nand U16391 (N_16391,N_14958,N_15103);
nor U16392 (N_16392,N_15728,N_15377);
or U16393 (N_16393,N_14596,N_14301);
or U16394 (N_16394,N_14542,N_14029);
nand U16395 (N_16395,N_14598,N_14166);
or U16396 (N_16396,N_15719,N_14907);
nor U16397 (N_16397,N_14929,N_15535);
and U16398 (N_16398,N_15147,N_15176);
or U16399 (N_16399,N_14427,N_15938);
xor U16400 (N_16400,N_14853,N_15442);
nor U16401 (N_16401,N_14182,N_14716);
nand U16402 (N_16402,N_15617,N_15378);
and U16403 (N_16403,N_15261,N_15164);
or U16404 (N_16404,N_15871,N_15340);
or U16405 (N_16405,N_15017,N_15928);
nor U16406 (N_16406,N_14473,N_14738);
nand U16407 (N_16407,N_15279,N_14847);
or U16408 (N_16408,N_15792,N_14450);
nand U16409 (N_16409,N_14725,N_15608);
nand U16410 (N_16410,N_15785,N_14758);
nand U16411 (N_16411,N_14663,N_15702);
nor U16412 (N_16412,N_14978,N_15606);
or U16413 (N_16413,N_14036,N_14027);
nand U16414 (N_16414,N_14555,N_15396);
nand U16415 (N_16415,N_14630,N_15542);
nor U16416 (N_16416,N_15308,N_15619);
and U16417 (N_16417,N_14460,N_15585);
nand U16418 (N_16418,N_15543,N_15544);
nand U16419 (N_16419,N_14603,N_15930);
nor U16420 (N_16420,N_15039,N_14865);
xnor U16421 (N_16421,N_14413,N_14836);
nor U16422 (N_16422,N_15128,N_15455);
and U16423 (N_16423,N_14957,N_15148);
xnor U16424 (N_16424,N_15077,N_14462);
nor U16425 (N_16425,N_15927,N_15071);
or U16426 (N_16426,N_15126,N_14579);
or U16427 (N_16427,N_15388,N_15738);
or U16428 (N_16428,N_14367,N_15506);
nand U16429 (N_16429,N_15853,N_14308);
nand U16430 (N_16430,N_14065,N_15096);
nand U16431 (N_16431,N_15135,N_14531);
nand U16432 (N_16432,N_15827,N_15242);
or U16433 (N_16433,N_14609,N_15216);
and U16434 (N_16434,N_14526,N_15133);
or U16435 (N_16435,N_14876,N_15364);
nand U16436 (N_16436,N_14447,N_15815);
or U16437 (N_16437,N_14562,N_15718);
and U16438 (N_16438,N_15456,N_14549);
and U16439 (N_16439,N_15682,N_14525);
or U16440 (N_16440,N_14386,N_15818);
xnor U16441 (N_16441,N_14898,N_15207);
nor U16442 (N_16442,N_14237,N_15403);
or U16443 (N_16443,N_15406,N_14006);
and U16444 (N_16444,N_14171,N_14787);
xor U16445 (N_16445,N_15074,N_14685);
xor U16446 (N_16446,N_14669,N_15399);
nand U16447 (N_16447,N_15797,N_14523);
nor U16448 (N_16448,N_15613,N_15280);
nor U16449 (N_16449,N_15634,N_14089);
nor U16450 (N_16450,N_15054,N_15104);
nor U16451 (N_16451,N_14478,N_14605);
or U16452 (N_16452,N_14292,N_14583);
nor U16453 (N_16453,N_14889,N_14302);
nand U16454 (N_16454,N_15171,N_14843);
or U16455 (N_16455,N_14062,N_15635);
or U16456 (N_16456,N_14955,N_15281);
nand U16457 (N_16457,N_15724,N_14390);
nor U16458 (N_16458,N_14981,N_14613);
or U16459 (N_16459,N_15896,N_15181);
nand U16460 (N_16460,N_14746,N_15363);
nor U16461 (N_16461,N_14906,N_14421);
or U16462 (N_16462,N_15739,N_14207);
nor U16463 (N_16463,N_14849,N_15520);
nand U16464 (N_16464,N_15895,N_14558);
nor U16465 (N_16465,N_14600,N_15908);
nand U16466 (N_16466,N_14561,N_15208);
and U16467 (N_16467,N_15170,N_14546);
nand U16468 (N_16468,N_14740,N_14499);
and U16469 (N_16469,N_15939,N_14120);
and U16470 (N_16470,N_14635,N_14618);
nor U16471 (N_16471,N_14616,N_14068);
or U16472 (N_16472,N_15937,N_14963);
nand U16473 (N_16473,N_15599,N_14629);
nor U16474 (N_16474,N_15180,N_15510);
nor U16475 (N_16475,N_14307,N_15641);
nor U16476 (N_16476,N_14788,N_15398);
xor U16477 (N_16477,N_14909,N_14125);
and U16478 (N_16478,N_15044,N_15509);
xnor U16479 (N_16479,N_14551,N_14162);
nand U16480 (N_16480,N_15616,N_14864);
nand U16481 (N_16481,N_14043,N_15972);
nor U16482 (N_16482,N_15736,N_15163);
xnor U16483 (N_16483,N_15665,N_14830);
and U16484 (N_16484,N_14805,N_14296);
and U16485 (N_16485,N_15907,N_15538);
or U16486 (N_16486,N_15925,N_14048);
or U16487 (N_16487,N_14340,N_14794);
and U16488 (N_16488,N_14476,N_14047);
or U16489 (N_16489,N_14811,N_15351);
or U16490 (N_16490,N_14783,N_14359);
nand U16491 (N_16491,N_15890,N_14129);
and U16492 (N_16492,N_15809,N_15316);
xor U16493 (N_16493,N_15525,N_15344);
nor U16494 (N_16494,N_15774,N_15512);
nand U16495 (N_16495,N_14096,N_15421);
nor U16496 (N_16496,N_14152,N_14912);
xnor U16497 (N_16497,N_14071,N_14233);
nand U16498 (N_16498,N_14406,N_15380);
nor U16499 (N_16499,N_14535,N_14024);
and U16500 (N_16500,N_14781,N_15132);
and U16501 (N_16501,N_14901,N_15422);
nor U16502 (N_16502,N_14195,N_15102);
nand U16503 (N_16503,N_14574,N_15244);
or U16504 (N_16504,N_14851,N_14088);
nand U16505 (N_16505,N_15487,N_14400);
or U16506 (N_16506,N_15799,N_14888);
nor U16507 (N_16507,N_15596,N_15213);
xor U16508 (N_16508,N_15107,N_14274);
and U16509 (N_16509,N_15651,N_15906);
nand U16510 (N_16510,N_14015,N_14455);
xnor U16511 (N_16511,N_14968,N_15947);
and U16512 (N_16512,N_15642,N_14178);
nor U16513 (N_16513,N_15949,N_14355);
and U16514 (N_16514,N_15700,N_15469);
nand U16515 (N_16515,N_15816,N_14980);
xor U16516 (N_16516,N_15914,N_14054);
nand U16517 (N_16517,N_15747,N_14329);
nand U16518 (N_16518,N_15699,N_14852);
and U16519 (N_16519,N_15805,N_14081);
xor U16520 (N_16520,N_15822,N_14926);
and U16521 (N_16521,N_14422,N_14334);
nor U16522 (N_16522,N_15390,N_15484);
nor U16523 (N_16523,N_14537,N_15221);
and U16524 (N_16524,N_14445,N_14277);
nand U16525 (N_16525,N_14997,N_14153);
or U16526 (N_16526,N_14763,N_14703);
and U16527 (N_16527,N_14664,N_15675);
xnor U16528 (N_16528,N_14782,N_15495);
and U16529 (N_16529,N_15303,N_14490);
and U16530 (N_16530,N_14659,N_14745);
or U16531 (N_16531,N_14973,N_15368);
and U16532 (N_16532,N_14147,N_15045);
or U16533 (N_16533,N_15598,N_15414);
nand U16534 (N_16534,N_14306,N_15263);
nand U16535 (N_16535,N_14528,N_14960);
nor U16536 (N_16536,N_15667,N_14737);
or U16537 (N_16537,N_14472,N_14510);
nand U16538 (N_16538,N_14322,N_14385);
and U16539 (N_16539,N_15703,N_15337);
and U16540 (N_16540,N_14253,N_15265);
nand U16541 (N_16541,N_14952,N_14381);
nand U16542 (N_16542,N_14030,N_14285);
or U16543 (N_16543,N_15784,N_14470);
nor U16544 (N_16544,N_15875,N_14769);
or U16545 (N_16545,N_15991,N_15188);
xnor U16546 (N_16546,N_15969,N_15142);
and U16547 (N_16547,N_15049,N_15040);
or U16548 (N_16548,N_14766,N_14484);
nand U16549 (N_16549,N_15539,N_15935);
xnor U16550 (N_16550,N_15253,N_14500);
nor U16551 (N_16551,N_14232,N_15674);
nor U16552 (N_16552,N_15698,N_15440);
nor U16553 (N_16553,N_15964,N_15282);
nor U16554 (N_16554,N_14364,N_15987);
xnor U16555 (N_16555,N_14491,N_15302);
or U16556 (N_16556,N_14032,N_14666);
and U16557 (N_16557,N_14000,N_15313);
or U16558 (N_16558,N_15094,N_14137);
or U16559 (N_16559,N_15647,N_14168);
and U16560 (N_16560,N_14736,N_15862);
and U16561 (N_16561,N_14739,N_14380);
and U16562 (N_16562,N_15227,N_15005);
and U16563 (N_16563,N_15968,N_15919);
and U16564 (N_16564,N_14240,N_15990);
nand U16565 (N_16565,N_15817,N_15463);
or U16566 (N_16566,N_14655,N_15210);
and U16567 (N_16567,N_15915,N_15806);
or U16568 (N_16568,N_15770,N_15152);
and U16569 (N_16569,N_14461,N_14206);
nor U16570 (N_16570,N_14079,N_14518);
and U16571 (N_16571,N_14956,N_15194);
nor U16572 (N_16572,N_14640,N_14050);
and U16573 (N_16573,N_14283,N_14361);
or U16574 (N_16574,N_15511,N_14700);
nor U16575 (N_16575,N_15825,N_15873);
or U16576 (N_16576,N_14753,N_15569);
nor U16577 (N_16577,N_15139,N_15158);
or U16578 (N_16578,N_14244,N_15453);
or U16579 (N_16579,N_15863,N_14483);
nor U16580 (N_16580,N_15090,N_15426);
nor U16581 (N_16581,N_15197,N_14905);
nor U16582 (N_16582,N_14440,N_14471);
or U16583 (N_16583,N_15772,N_15775);
nand U16584 (N_16584,N_15627,N_14577);
nor U16585 (N_16585,N_15024,N_15016);
nor U16586 (N_16586,N_15352,N_14569);
nand U16587 (N_16587,N_15884,N_14205);
or U16588 (N_16588,N_15611,N_14184);
and U16589 (N_16589,N_15424,N_15289);
nor U16590 (N_16590,N_14313,N_14839);
nand U16591 (N_16591,N_15269,N_15006);
nor U16592 (N_16592,N_14812,N_14291);
and U16593 (N_16593,N_14858,N_15066);
xor U16594 (N_16594,N_15500,N_14133);
nor U16595 (N_16595,N_15683,N_14356);
nand U16596 (N_16596,N_14899,N_14016);
and U16597 (N_16597,N_15315,N_15583);
or U16598 (N_16598,N_15297,N_14813);
or U16599 (N_16599,N_15252,N_14610);
or U16600 (N_16600,N_14726,N_15450);
nor U16601 (N_16601,N_14160,N_15685);
or U16602 (N_16602,N_14368,N_15026);
nand U16603 (N_16603,N_14486,N_14683);
and U16604 (N_16604,N_14148,N_15325);
nor U16605 (N_16605,N_15942,N_14010);
nor U16606 (N_16606,N_15638,N_15117);
nor U16607 (N_16607,N_15012,N_15249);
nor U16608 (N_16608,N_15948,N_15780);
nor U16609 (N_16609,N_14245,N_15716);
nor U16610 (N_16610,N_15189,N_14458);
nor U16611 (N_16611,N_14756,N_15334);
and U16612 (N_16612,N_14859,N_15338);
nor U16613 (N_16613,N_15727,N_15746);
or U16614 (N_16614,N_14869,N_15499);
nand U16615 (N_16615,N_14211,N_15447);
or U16616 (N_16616,N_15028,N_15018);
or U16617 (N_16617,N_15720,N_15916);
xor U16618 (N_16618,N_15140,N_14064);
xnor U16619 (N_16619,N_15432,N_14744);
xnor U16620 (N_16620,N_15429,N_15036);
nor U16621 (N_16621,N_15941,N_14947);
or U16622 (N_16622,N_15127,N_14902);
and U16623 (N_16623,N_14673,N_14132);
or U16624 (N_16624,N_15136,N_15802);
xnor U16625 (N_16625,N_14970,N_14702);
or U16626 (N_16626,N_15385,N_15400);
and U16627 (N_16627,N_15560,N_14770);
nor U16628 (N_16628,N_15035,N_15882);
nand U16629 (N_16629,N_15278,N_15489);
xnor U16630 (N_16630,N_14128,N_14154);
and U16631 (N_16631,N_15962,N_15940);
and U16632 (N_16632,N_15382,N_15250);
or U16633 (N_16633,N_14931,N_15138);
and U16634 (N_16634,N_15621,N_15177);
or U16635 (N_16635,N_14863,N_15821);
nand U16636 (N_16636,N_15791,N_15446);
nor U16637 (N_16637,N_14430,N_15692);
nand U16638 (N_16638,N_14878,N_15759);
or U16639 (N_16639,N_15166,N_14848);
xor U16640 (N_16640,N_15314,N_14423);
or U16641 (N_16641,N_14023,N_15865);
or U16642 (N_16642,N_14661,N_15839);
nor U16643 (N_16643,N_14547,N_15209);
nand U16644 (N_16644,N_15742,N_15425);
xnor U16645 (N_16645,N_14602,N_14866);
or U16646 (N_16646,N_15384,N_15963);
or U16647 (N_16647,N_15153,N_14199);
nor U16648 (N_16648,N_14021,N_14117);
nor U16649 (N_16649,N_14710,N_15643);
nor U16650 (N_16650,N_14001,N_14687);
and U16651 (N_16651,N_14994,N_14140);
nor U16652 (N_16652,N_15847,N_14601);
nand U16653 (N_16653,N_14810,N_14747);
nand U16654 (N_16654,N_14127,N_15119);
or U16655 (N_16655,N_14150,N_15020);
nand U16656 (N_16656,N_15733,N_14924);
xnor U16657 (N_16657,N_15660,N_15661);
or U16658 (N_16658,N_14286,N_15904);
nor U16659 (N_16659,N_15529,N_14799);
and U16660 (N_16660,N_15899,N_14668);
or U16661 (N_16661,N_14197,N_14641);
or U16662 (N_16662,N_14512,N_14959);
nor U16663 (N_16663,N_14442,N_14311);
or U16664 (N_16664,N_15794,N_15796);
nor U16665 (N_16665,N_14834,N_15679);
and U16666 (N_16666,N_15004,N_15258);
nand U16667 (N_16667,N_15609,N_15299);
nand U16668 (N_16668,N_15548,N_15149);
nand U16669 (N_16669,N_14250,N_14619);
and U16670 (N_16670,N_15008,N_14748);
or U16671 (N_16671,N_14750,N_14183);
nor U16672 (N_16672,N_15475,N_15042);
nand U16673 (N_16673,N_14976,N_14007);
nor U16674 (N_16674,N_15239,N_14333);
nor U16675 (N_16675,N_14690,N_15361);
xor U16676 (N_16676,N_15501,N_15223);
and U16677 (N_16677,N_14713,N_15321);
nor U16678 (N_16678,N_15695,N_14896);
nand U16679 (N_16679,N_14169,N_14139);
and U16680 (N_16680,N_15287,N_15427);
or U16681 (N_16681,N_15984,N_15449);
or U16682 (N_16682,N_15106,N_14914);
or U16683 (N_16683,N_15485,N_14111);
or U16684 (N_16684,N_15123,N_15910);
nor U16685 (N_16685,N_14940,N_14776);
nand U16686 (N_16686,N_14180,N_15043);
nand U16687 (N_16687,N_15790,N_14058);
nor U16688 (N_16688,N_15358,N_15696);
nor U16689 (N_16689,N_15064,N_14991);
or U16690 (N_16690,N_14995,N_15783);
nand U16691 (N_16691,N_14831,N_14591);
nor U16692 (N_16692,N_14397,N_15625);
xnor U16693 (N_16693,N_15257,N_15576);
and U16694 (N_16694,N_14375,N_15523);
xor U16695 (N_16695,N_15917,N_15273);
nor U16696 (N_16696,N_14444,N_14779);
nand U16697 (N_16697,N_14818,N_15934);
nand U16698 (N_16698,N_14972,N_14468);
and U16699 (N_16699,N_14570,N_15038);
nor U16700 (N_16700,N_14441,N_14815);
or U16701 (N_16701,N_14067,N_14049);
and U16702 (N_16702,N_15517,N_14479);
nand U16703 (N_16703,N_15932,N_14646);
or U16704 (N_16704,N_14118,N_14022);
or U16705 (N_16705,N_15290,N_15804);
or U16706 (N_16706,N_15228,N_14060);
nand U16707 (N_16707,N_14325,N_15900);
xnor U16708 (N_16708,N_15168,N_14543);
nand U16709 (N_16709,N_14607,N_14409);
or U16710 (N_16710,N_14263,N_14757);
nor U16711 (N_16711,N_15305,N_14989);
nand U16712 (N_16712,N_14246,N_15318);
and U16713 (N_16713,N_14056,N_14352);
and U16714 (N_16714,N_14219,N_14113);
nor U16715 (N_16715,N_15633,N_14281);
nand U16716 (N_16716,N_14063,N_14808);
or U16717 (N_16717,N_15100,N_15901);
or U16718 (N_16718,N_15922,N_14407);
nand U16719 (N_16719,N_14242,N_15231);
nor U16720 (N_16720,N_14013,N_15676);
nand U16721 (N_16721,N_15371,N_14443);
or U16722 (N_16722,N_14532,N_14045);
xor U16723 (N_16723,N_14267,N_14765);
or U16724 (N_16724,N_14345,N_14833);
and U16725 (N_16725,N_15826,N_15069);
and U16726 (N_16726,N_15866,N_15557);
nor U16727 (N_16727,N_15717,N_15787);
nor U16728 (N_16728,N_15859,N_14797);
or U16729 (N_16729,N_15076,N_14883);
or U16730 (N_16730,N_15454,N_15369);
and U16731 (N_16731,N_14087,N_15632);
nand U16732 (N_16732,N_14227,N_15120);
nor U16733 (N_16733,N_14636,N_15894);
and U16734 (N_16734,N_14792,N_15402);
nand U16735 (N_16735,N_15381,N_14280);
and U16736 (N_16736,N_15434,N_15886);
xnor U16737 (N_16737,N_15514,N_15124);
or U16738 (N_16738,N_14946,N_14854);
nand U16739 (N_16739,N_15254,N_14662);
nand U16740 (N_16740,N_14625,N_14382);
nand U16741 (N_16741,N_14101,N_15730);
or U16742 (N_16742,N_15977,N_14708);
and U16743 (N_16743,N_15578,N_15897);
and U16744 (N_16744,N_14141,N_15423);
nand U16745 (N_16745,N_15740,N_14019);
or U16746 (N_16746,N_14121,N_15684);
or U16747 (N_16747,N_15519,N_15518);
and U16748 (N_16748,N_14383,N_14828);
and U16749 (N_16749,N_15007,N_14480);
and U16750 (N_16750,N_15751,N_15571);
or U16751 (N_16751,N_15670,N_14069);
or U16752 (N_16752,N_14432,N_15460);
nand U16753 (N_16753,N_14279,N_14115);
nor U16754 (N_16754,N_15885,N_15707);
nand U16755 (N_16755,N_14733,N_15161);
and U16756 (N_16756,N_15323,N_15031);
or U16757 (N_16757,N_15553,N_15346);
nand U16758 (N_16758,N_14665,N_15754);
and U16759 (N_16759,N_14873,N_15236);
nand U16760 (N_16760,N_14872,N_15248);
and U16761 (N_16761,N_15931,N_15159);
and U16762 (N_16762,N_15841,N_14335);
or U16763 (N_16763,N_14332,N_14210);
and U16764 (N_16764,N_15680,N_14214);
or U16765 (N_16765,N_14731,N_15849);
or U16766 (N_16766,N_14606,N_15420);
or U16767 (N_16767,N_14076,N_14971);
nand U16768 (N_16768,N_15365,N_15888);
nor U16769 (N_16769,N_14228,N_14882);
or U16770 (N_16770,N_14755,N_14401);
and U16771 (N_16771,N_14289,N_14474);
or U16772 (N_16772,N_14316,N_14897);
or U16773 (N_16773,N_15160,N_15593);
or U16774 (N_16774,N_15678,N_14092);
or U16775 (N_16775,N_15322,N_15918);
or U16776 (N_16776,N_15105,N_14221);
nand U16777 (N_16777,N_14845,N_15268);
nand U16778 (N_16778,N_15312,N_14389);
and U16779 (N_16779,N_14363,N_14679);
nor U16780 (N_16780,N_14519,N_14405);
nand U16781 (N_16781,N_14312,N_14464);
or U16782 (N_16782,N_15172,N_15550);
and U16783 (N_16783,N_14482,N_14435);
nor U16784 (N_16784,N_14396,N_15929);
nand U16785 (N_16785,N_15309,N_15492);
nor U16786 (N_16786,N_14785,N_14749);
or U16787 (N_16787,N_14151,N_15793);
or U16788 (N_16788,N_14774,N_15810);
and U16789 (N_16789,N_14784,N_15836);
nand U16790 (N_16790,N_15668,N_15909);
xor U16791 (N_16791,N_15110,N_14456);
nor U16792 (N_16792,N_14082,N_14590);
nand U16793 (N_16793,N_14806,N_15846);
xor U16794 (N_16794,N_14507,N_14594);
xnor U16795 (N_16795,N_14974,N_15014);
or U16796 (N_16796,N_14235,N_14714);
or U16797 (N_16797,N_15304,N_14891);
nand U16798 (N_16798,N_14173,N_14085);
or U16799 (N_16799,N_14672,N_15488);
nand U16800 (N_16800,N_15436,N_15370);
or U16801 (N_16801,N_15298,N_15532);
nor U16802 (N_16802,N_14564,N_15577);
nand U16803 (N_16803,N_14634,N_15230);
or U16804 (N_16804,N_15662,N_14175);
and U16805 (N_16805,N_15620,N_14586);
nor U16806 (N_16806,N_14230,N_14028);
nand U16807 (N_16807,N_15803,N_15920);
and U16808 (N_16808,N_15669,N_14026);
and U16809 (N_16809,N_14597,N_14730);
or U16810 (N_16810,N_14884,N_14261);
and U16811 (N_16811,N_14260,N_15439);
nand U16812 (N_16812,N_15205,N_15798);
or U16813 (N_16813,N_15174,N_14103);
and U16814 (N_16814,N_15677,N_15214);
xor U16815 (N_16815,N_14156,N_15443);
nand U16816 (N_16816,N_14538,N_14106);
nand U16817 (N_16817,N_14231,N_14734);
nor U16818 (N_16818,N_14225,N_14615);
or U16819 (N_16819,N_14604,N_14916);
nor U16820 (N_16820,N_14020,N_14516);
or U16821 (N_16821,N_14465,N_14922);
nor U16822 (N_16822,N_14420,N_14303);
nor U16823 (N_16823,N_15141,N_14846);
or U16824 (N_16824,N_15348,N_15721);
nor U16825 (N_16825,N_15379,N_14695);
and U16826 (N_16826,N_14953,N_14724);
and U16827 (N_16827,N_14514,N_14582);
or U16828 (N_16828,N_15776,N_14164);
nand U16829 (N_16829,N_14181,N_15418);
and U16830 (N_16830,N_15961,N_14800);
and U16831 (N_16831,N_14377,N_15600);
or U16832 (N_16832,N_14977,N_15047);
nand U16833 (N_16833,N_15157,N_14494);
and U16834 (N_16834,N_15547,N_15623);
xnor U16835 (N_16835,N_15686,N_15838);
and U16836 (N_16836,N_15445,N_14138);
and U16837 (N_16837,N_15283,N_15491);
nor U16838 (N_16838,N_15339,N_15151);
and U16839 (N_16839,N_15360,N_15536);
or U16840 (N_16840,N_14354,N_14264);
xnor U16841 (N_16841,N_14346,N_15101);
and U16842 (N_16842,N_14768,N_15735);
nor U16843 (N_16843,N_14282,N_14370);
nand U16844 (N_16844,N_15533,N_14426);
nand U16845 (N_16845,N_15891,N_15526);
nor U16846 (N_16846,N_14319,N_14143);
nor U16847 (N_16847,N_14678,N_14676);
and U16848 (N_16848,N_15950,N_15395);
nand U16849 (N_16849,N_15029,N_14624);
nor U16850 (N_16850,N_14170,N_14287);
nor U16851 (N_16851,N_14320,N_15203);
and U16852 (N_16852,N_15478,N_14576);
or U16853 (N_16853,N_14224,N_14353);
nand U16854 (N_16854,N_14536,N_15274);
nand U16855 (N_16855,N_14773,N_14348);
nand U16856 (N_16856,N_15187,N_14950);
nand U16857 (N_16857,N_15353,N_14208);
xor U16858 (N_16858,N_14741,N_14270);
and U16859 (N_16859,N_14803,N_14910);
nor U16860 (N_16860,N_15310,N_14827);
and U16861 (N_16861,N_15288,N_14948);
or U16862 (N_16862,N_15327,N_14647);
nand U16863 (N_16863,N_14822,N_15480);
nor U16864 (N_16864,N_15581,N_14575);
and U16865 (N_16865,N_14009,N_15072);
and U16866 (N_16866,N_14326,N_15502);
nor U16867 (N_16867,N_15779,N_14256);
and U16868 (N_16868,N_15145,N_15068);
nand U16869 (N_16869,N_14366,N_15967);
nor U16870 (N_16870,N_15845,N_15970);
or U16871 (N_16871,N_15926,N_15945);
and U16872 (N_16872,N_15435,N_15657);
nor U16873 (N_16873,N_15921,N_14003);
nand U16874 (N_16874,N_15459,N_14617);
nand U16875 (N_16875,N_15084,N_14254);
nor U16876 (N_16876,N_14418,N_14550);
or U16877 (N_16877,N_15854,N_14653);
xor U16878 (N_16878,N_15640,N_15342);
nand U16879 (N_16879,N_14961,N_15689);
or U16880 (N_16880,N_14520,N_15568);
nand U16881 (N_16881,N_14194,N_14985);
or U16882 (N_16882,N_15413,N_15843);
nand U16883 (N_16883,N_15830,N_15508);
nor U16884 (N_16884,N_14881,N_15393);
nand U16885 (N_16885,N_15419,N_15762);
or U16886 (N_16886,N_15591,N_15618);
nor U16887 (N_16887,N_15220,N_15311);
or U16888 (N_16888,N_15749,N_15615);
nor U16889 (N_16889,N_15766,N_15367);
nand U16890 (N_16890,N_14919,N_15349);
nand U16891 (N_16891,N_15201,N_14328);
or U16892 (N_16892,N_15988,N_14452);
or U16893 (N_16893,N_14347,N_14628);
nand U16894 (N_16894,N_15131,N_15033);
nand U16895 (N_16895,N_15955,N_15409);
xnor U16896 (N_16896,N_14262,N_15978);
or U16897 (N_16897,N_15953,N_14310);
and U16898 (N_16898,N_15629,N_14593);
nand U16899 (N_16899,N_15458,N_14809);
nand U16900 (N_16900,N_15829,N_14540);
and U16901 (N_16901,N_15556,N_14650);
xor U16902 (N_16902,N_14031,N_14621);
nor U16903 (N_16903,N_15034,N_14074);
nor U16904 (N_16904,N_14840,N_14707);
and U16905 (N_16905,N_15722,N_14671);
xnor U16906 (N_16906,N_15467,N_15778);
nand U16907 (N_16907,N_14290,N_14622);
and U16908 (N_16908,N_15009,N_14743);
or U16909 (N_16909,N_14823,N_14969);
nand U16910 (N_16910,N_15000,N_14627);
or U16911 (N_16911,N_15087,N_15986);
or U16912 (N_16912,N_15750,N_15431);
and U16913 (N_16913,N_14416,N_15777);
nor U16914 (N_16914,N_15391,N_14993);
or U16915 (N_16915,N_15743,N_15867);
nor U16916 (N_16916,N_14498,N_15493);
and U16917 (N_16917,N_15555,N_15565);
and U16918 (N_16918,N_14165,N_15575);
and U16919 (N_16919,N_14337,N_14034);
nand U16920 (N_16920,N_14572,N_15284);
and U16921 (N_16921,N_15605,N_15295);
nor U16922 (N_16922,N_15893,N_15959);
xnor U16923 (N_16923,N_15225,N_15183);
nor U16924 (N_16924,N_14933,N_14996);
nand U16925 (N_16925,N_14860,N_14771);
or U16926 (N_16926,N_15457,N_15630);
or U16927 (N_16927,N_15200,N_15182);
and U16928 (N_16928,N_14712,N_15840);
nand U16929 (N_16929,N_14459,N_15095);
nand U16930 (N_16930,N_15405,N_15649);
or U16931 (N_16931,N_15800,N_15808);
and U16932 (N_16932,N_15116,N_15708);
nand U16933 (N_16933,N_15115,N_14824);
nor U16934 (N_16934,N_14539,N_15444);
nand U16935 (N_16935,N_15185,N_14318);
xnor U16936 (N_16936,N_15078,N_14517);
xor U16937 (N_16937,N_15441,N_14694);
and U16938 (N_16938,N_15376,N_14819);
nor U16939 (N_16939,N_15701,N_14506);
nand U16940 (N_16940,N_15588,N_14378);
nand U16941 (N_16941,N_15912,N_14149);
nor U16942 (N_16942,N_14252,N_15663);
and U16943 (N_16943,N_14660,N_14344);
and U16944 (N_16944,N_15760,N_14309);
or U16945 (N_16945,N_15744,N_15010);
and U16946 (N_16946,N_14110,N_15877);
xnor U16947 (N_16947,N_14218,N_14203);
or U16948 (N_16948,N_14485,N_15541);
nand U16949 (N_16949,N_15374,N_14871);
nor U16950 (N_16950,N_15694,N_14080);
or U16951 (N_16951,N_14534,N_14711);
nor U16952 (N_16952,N_14294,N_15490);
and U16953 (N_16953,N_14857,N_15960);
nand U16954 (N_16954,N_15898,N_15652);
and U16955 (N_16955,N_15468,N_15582);
nor U16956 (N_16956,N_15712,N_15835);
xor U16957 (N_16957,N_15291,N_14688);
xor U16958 (N_16958,N_14090,N_15831);
or U16959 (N_16959,N_15307,N_15061);
nor U16960 (N_16960,N_15324,N_14158);
nand U16961 (N_16961,N_15146,N_14358);
nor U16962 (N_16962,N_15089,N_14675);
or U16963 (N_16963,N_15807,N_14503);
and U16964 (N_16964,N_15328,N_15165);
xnor U16965 (N_16965,N_14638,N_15062);
nor U16966 (N_16966,N_14131,N_15129);
nor U16967 (N_16967,N_14826,N_15190);
nor U16968 (N_16968,N_15503,N_14033);
or U16969 (N_16969,N_14119,N_15494);
nor U16970 (N_16970,N_15067,N_15483);
nor U16971 (N_16971,N_14642,N_15497);
nand U16972 (N_16972,N_15092,N_14135);
and U16973 (N_16973,N_15118,N_15041);
nor U16974 (N_16974,N_14751,N_15202);
or U16975 (N_16975,N_15448,N_15654);
nor U16976 (N_16976,N_14467,N_14798);
or U16977 (N_16977,N_14780,N_14454);
nor U16978 (N_16978,N_15229,N_15465);
nand U16979 (N_16979,N_14802,N_15531);
nand U16980 (N_16980,N_15355,N_15881);
or U16981 (N_16981,N_14513,N_14317);
nand U16982 (N_16982,N_14086,N_14035);
nand U16983 (N_16983,N_15671,N_14632);
or U16984 (N_16984,N_14202,N_14109);
xnor U16985 (N_16985,N_14425,N_14257);
or U16986 (N_16986,N_14608,N_15561);
or U16987 (N_16987,N_15876,N_14742);
xnor U16988 (N_16988,N_14786,N_14890);
nor U16989 (N_16989,N_15911,N_14917);
nor U16990 (N_16990,N_15993,N_15073);
nor U16991 (N_16991,N_15317,N_15590);
xor U16992 (N_16992,N_14393,N_15655);
and U16993 (N_16993,N_15025,N_14585);
nand U16994 (N_16994,N_14704,N_15451);
xor U16995 (N_16995,N_15150,N_14336);
and U16996 (N_16996,N_15650,N_15343);
and U16997 (N_16997,N_14511,N_14072);
or U16998 (N_16998,N_14578,N_14330);
nand U16999 (N_16999,N_15537,N_15566);
xnor U17000 (N_17000,N_14344,N_14205);
xor U17001 (N_17001,N_15631,N_15405);
nand U17002 (N_17002,N_15443,N_14918);
or U17003 (N_17003,N_14308,N_15466);
and U17004 (N_17004,N_14553,N_15755);
and U17005 (N_17005,N_14597,N_15834);
or U17006 (N_17006,N_14962,N_14171);
or U17007 (N_17007,N_15716,N_15129);
nand U17008 (N_17008,N_14123,N_15894);
and U17009 (N_17009,N_14402,N_14954);
and U17010 (N_17010,N_15473,N_14667);
nor U17011 (N_17011,N_14813,N_15218);
nor U17012 (N_17012,N_14583,N_15744);
nor U17013 (N_17013,N_15860,N_15551);
or U17014 (N_17014,N_15836,N_14691);
and U17015 (N_17015,N_15164,N_14103);
nand U17016 (N_17016,N_15729,N_14953);
and U17017 (N_17017,N_15878,N_14889);
xor U17018 (N_17018,N_15208,N_14888);
or U17019 (N_17019,N_14233,N_14274);
nor U17020 (N_17020,N_15215,N_14013);
and U17021 (N_17021,N_15355,N_14523);
or U17022 (N_17022,N_15533,N_14013);
nand U17023 (N_17023,N_14785,N_15859);
nand U17024 (N_17024,N_15691,N_15328);
nor U17025 (N_17025,N_15249,N_15234);
nand U17026 (N_17026,N_15288,N_14387);
xor U17027 (N_17027,N_14196,N_15280);
nor U17028 (N_17028,N_14093,N_15970);
xor U17029 (N_17029,N_15436,N_15554);
nand U17030 (N_17030,N_15874,N_15479);
or U17031 (N_17031,N_14380,N_15804);
nand U17032 (N_17032,N_14319,N_14174);
xor U17033 (N_17033,N_15906,N_14798);
and U17034 (N_17034,N_15600,N_15599);
nand U17035 (N_17035,N_15349,N_15532);
and U17036 (N_17036,N_14764,N_14559);
nand U17037 (N_17037,N_14654,N_15745);
and U17038 (N_17038,N_14809,N_14775);
nor U17039 (N_17039,N_14339,N_15366);
xor U17040 (N_17040,N_15429,N_15025);
nor U17041 (N_17041,N_15126,N_15715);
or U17042 (N_17042,N_14045,N_15328);
nor U17043 (N_17043,N_14272,N_15234);
or U17044 (N_17044,N_15625,N_15560);
xnor U17045 (N_17045,N_14836,N_15228);
nor U17046 (N_17046,N_15631,N_14302);
and U17047 (N_17047,N_15477,N_15862);
nor U17048 (N_17048,N_15501,N_15204);
nor U17049 (N_17049,N_15843,N_15584);
and U17050 (N_17050,N_15867,N_15697);
nor U17051 (N_17051,N_14678,N_15689);
or U17052 (N_17052,N_15873,N_14820);
nand U17053 (N_17053,N_15138,N_15589);
xor U17054 (N_17054,N_14821,N_14204);
or U17055 (N_17055,N_15737,N_14866);
xor U17056 (N_17056,N_14660,N_15122);
or U17057 (N_17057,N_14004,N_14904);
nor U17058 (N_17058,N_15379,N_14003);
nand U17059 (N_17059,N_14074,N_15662);
nand U17060 (N_17060,N_15863,N_15637);
xnor U17061 (N_17061,N_14454,N_15326);
and U17062 (N_17062,N_14280,N_14186);
nand U17063 (N_17063,N_15294,N_15407);
and U17064 (N_17064,N_14484,N_15254);
and U17065 (N_17065,N_15829,N_15812);
xor U17066 (N_17066,N_14275,N_14101);
or U17067 (N_17067,N_14222,N_14512);
nor U17068 (N_17068,N_14948,N_14081);
nor U17069 (N_17069,N_14232,N_15728);
or U17070 (N_17070,N_14396,N_14356);
nor U17071 (N_17071,N_14081,N_15727);
xnor U17072 (N_17072,N_15324,N_14427);
and U17073 (N_17073,N_14063,N_14748);
and U17074 (N_17074,N_14338,N_14889);
nor U17075 (N_17075,N_14561,N_15936);
and U17076 (N_17076,N_15227,N_14686);
and U17077 (N_17077,N_14352,N_15004);
xor U17078 (N_17078,N_15853,N_15284);
and U17079 (N_17079,N_14562,N_15066);
or U17080 (N_17080,N_15076,N_15167);
or U17081 (N_17081,N_15814,N_15633);
or U17082 (N_17082,N_15770,N_15253);
nand U17083 (N_17083,N_15466,N_15489);
nor U17084 (N_17084,N_15562,N_15503);
nor U17085 (N_17085,N_14028,N_15010);
xor U17086 (N_17086,N_15134,N_15733);
and U17087 (N_17087,N_15678,N_15004);
nand U17088 (N_17088,N_15569,N_15346);
nand U17089 (N_17089,N_14648,N_15352);
or U17090 (N_17090,N_15365,N_15750);
nand U17091 (N_17091,N_15451,N_14163);
nand U17092 (N_17092,N_14149,N_15304);
nand U17093 (N_17093,N_14460,N_15503);
or U17094 (N_17094,N_15234,N_15598);
nand U17095 (N_17095,N_14091,N_14953);
or U17096 (N_17096,N_15812,N_14018);
xnor U17097 (N_17097,N_14845,N_15316);
nand U17098 (N_17098,N_15485,N_14689);
nand U17099 (N_17099,N_14611,N_14395);
nor U17100 (N_17100,N_14870,N_14395);
nand U17101 (N_17101,N_14500,N_14869);
or U17102 (N_17102,N_14802,N_15173);
and U17103 (N_17103,N_15360,N_14616);
nand U17104 (N_17104,N_14808,N_15033);
or U17105 (N_17105,N_15627,N_14163);
nor U17106 (N_17106,N_15851,N_14191);
nand U17107 (N_17107,N_14955,N_14607);
or U17108 (N_17108,N_15110,N_15229);
or U17109 (N_17109,N_15169,N_15210);
xor U17110 (N_17110,N_14714,N_15981);
or U17111 (N_17111,N_14513,N_15849);
nor U17112 (N_17112,N_15466,N_15668);
or U17113 (N_17113,N_14069,N_15335);
nand U17114 (N_17114,N_14167,N_15344);
and U17115 (N_17115,N_14168,N_14909);
or U17116 (N_17116,N_14806,N_15789);
and U17117 (N_17117,N_14583,N_14720);
or U17118 (N_17118,N_14582,N_15860);
nand U17119 (N_17119,N_15213,N_15174);
or U17120 (N_17120,N_14507,N_15544);
and U17121 (N_17121,N_15732,N_14696);
nor U17122 (N_17122,N_14542,N_14599);
nand U17123 (N_17123,N_15115,N_14870);
and U17124 (N_17124,N_15584,N_14068);
or U17125 (N_17125,N_15951,N_15952);
nand U17126 (N_17126,N_15384,N_15066);
and U17127 (N_17127,N_14688,N_14244);
and U17128 (N_17128,N_15685,N_14005);
nand U17129 (N_17129,N_14892,N_14594);
or U17130 (N_17130,N_15775,N_14695);
or U17131 (N_17131,N_14115,N_15450);
xnor U17132 (N_17132,N_14512,N_14188);
or U17133 (N_17133,N_15233,N_14230);
nand U17134 (N_17134,N_15923,N_15621);
nand U17135 (N_17135,N_14040,N_14631);
nand U17136 (N_17136,N_14154,N_14385);
nor U17137 (N_17137,N_15045,N_14571);
or U17138 (N_17138,N_15690,N_14018);
and U17139 (N_17139,N_14368,N_15552);
nand U17140 (N_17140,N_14094,N_14690);
nor U17141 (N_17141,N_14407,N_15154);
xor U17142 (N_17142,N_14834,N_15955);
or U17143 (N_17143,N_14404,N_14564);
nand U17144 (N_17144,N_15588,N_15567);
nor U17145 (N_17145,N_14056,N_14625);
or U17146 (N_17146,N_15142,N_15993);
nor U17147 (N_17147,N_15515,N_14622);
and U17148 (N_17148,N_15372,N_15302);
and U17149 (N_17149,N_14051,N_15991);
nand U17150 (N_17150,N_15077,N_14213);
nor U17151 (N_17151,N_15445,N_14416);
nor U17152 (N_17152,N_14168,N_15259);
nand U17153 (N_17153,N_14048,N_15001);
or U17154 (N_17154,N_15776,N_14339);
nor U17155 (N_17155,N_15083,N_14798);
nor U17156 (N_17156,N_15449,N_14733);
xor U17157 (N_17157,N_14070,N_14889);
nor U17158 (N_17158,N_15081,N_15929);
nor U17159 (N_17159,N_15086,N_14104);
and U17160 (N_17160,N_14981,N_14455);
nor U17161 (N_17161,N_14524,N_14502);
nor U17162 (N_17162,N_14068,N_14691);
nor U17163 (N_17163,N_15465,N_15887);
and U17164 (N_17164,N_14564,N_14010);
nor U17165 (N_17165,N_15429,N_15837);
nor U17166 (N_17166,N_14918,N_14020);
or U17167 (N_17167,N_15502,N_15688);
nand U17168 (N_17168,N_14762,N_15466);
xnor U17169 (N_17169,N_14231,N_15085);
and U17170 (N_17170,N_15200,N_14077);
or U17171 (N_17171,N_14848,N_15786);
and U17172 (N_17172,N_15873,N_15703);
nand U17173 (N_17173,N_15229,N_14193);
and U17174 (N_17174,N_15909,N_15565);
or U17175 (N_17175,N_14633,N_14807);
or U17176 (N_17176,N_14369,N_14971);
and U17177 (N_17177,N_15297,N_14691);
nor U17178 (N_17178,N_14363,N_15319);
and U17179 (N_17179,N_15605,N_14391);
nand U17180 (N_17180,N_14241,N_14513);
or U17181 (N_17181,N_14999,N_14916);
nor U17182 (N_17182,N_15649,N_15797);
or U17183 (N_17183,N_14441,N_15712);
nand U17184 (N_17184,N_15952,N_15499);
nand U17185 (N_17185,N_15482,N_14872);
or U17186 (N_17186,N_14080,N_15730);
nor U17187 (N_17187,N_14580,N_15550);
nand U17188 (N_17188,N_14500,N_14695);
nor U17189 (N_17189,N_14328,N_15099);
nand U17190 (N_17190,N_15839,N_15949);
nand U17191 (N_17191,N_14540,N_15129);
or U17192 (N_17192,N_15918,N_14946);
xor U17193 (N_17193,N_15901,N_14438);
and U17194 (N_17194,N_15635,N_14546);
and U17195 (N_17195,N_14023,N_14944);
nor U17196 (N_17196,N_14270,N_15936);
and U17197 (N_17197,N_15106,N_15223);
or U17198 (N_17198,N_15810,N_15226);
or U17199 (N_17199,N_15305,N_15773);
nand U17200 (N_17200,N_14949,N_14277);
nand U17201 (N_17201,N_15023,N_15507);
nor U17202 (N_17202,N_15157,N_15760);
nor U17203 (N_17203,N_15048,N_14268);
and U17204 (N_17204,N_14871,N_15442);
nand U17205 (N_17205,N_14810,N_15304);
nand U17206 (N_17206,N_14558,N_15975);
nand U17207 (N_17207,N_15130,N_15053);
and U17208 (N_17208,N_15389,N_14439);
or U17209 (N_17209,N_14945,N_15841);
nand U17210 (N_17210,N_14468,N_14188);
or U17211 (N_17211,N_14681,N_15274);
xor U17212 (N_17212,N_15794,N_14664);
xor U17213 (N_17213,N_14234,N_15951);
and U17214 (N_17214,N_14459,N_14028);
xor U17215 (N_17215,N_15030,N_14140);
xor U17216 (N_17216,N_14942,N_14796);
nor U17217 (N_17217,N_15743,N_14840);
xnor U17218 (N_17218,N_14981,N_15758);
or U17219 (N_17219,N_14167,N_15944);
and U17220 (N_17220,N_15689,N_15535);
xnor U17221 (N_17221,N_14989,N_14455);
nand U17222 (N_17222,N_14643,N_15253);
nand U17223 (N_17223,N_15922,N_14136);
nand U17224 (N_17224,N_14875,N_15314);
or U17225 (N_17225,N_15975,N_14294);
and U17226 (N_17226,N_14092,N_14215);
and U17227 (N_17227,N_15416,N_15490);
nor U17228 (N_17228,N_14602,N_14795);
or U17229 (N_17229,N_15561,N_14796);
or U17230 (N_17230,N_15534,N_15034);
or U17231 (N_17231,N_14120,N_15430);
and U17232 (N_17232,N_14262,N_15478);
nor U17233 (N_17233,N_15142,N_14775);
or U17234 (N_17234,N_14698,N_14842);
nor U17235 (N_17235,N_15935,N_14142);
or U17236 (N_17236,N_15179,N_14530);
and U17237 (N_17237,N_14862,N_14840);
and U17238 (N_17238,N_15328,N_14014);
or U17239 (N_17239,N_14078,N_15464);
or U17240 (N_17240,N_15649,N_14342);
nand U17241 (N_17241,N_15951,N_15462);
or U17242 (N_17242,N_15887,N_15242);
nand U17243 (N_17243,N_15419,N_14542);
and U17244 (N_17244,N_15142,N_14358);
or U17245 (N_17245,N_15482,N_15442);
or U17246 (N_17246,N_14758,N_15771);
nor U17247 (N_17247,N_14305,N_15201);
xnor U17248 (N_17248,N_14513,N_14125);
xnor U17249 (N_17249,N_15099,N_14078);
nand U17250 (N_17250,N_14841,N_15830);
and U17251 (N_17251,N_14011,N_14003);
nand U17252 (N_17252,N_15206,N_14828);
nand U17253 (N_17253,N_14909,N_15832);
and U17254 (N_17254,N_14891,N_14328);
nand U17255 (N_17255,N_14757,N_15904);
xnor U17256 (N_17256,N_14834,N_14103);
nor U17257 (N_17257,N_14778,N_15499);
nor U17258 (N_17258,N_14942,N_15752);
nand U17259 (N_17259,N_15323,N_14196);
and U17260 (N_17260,N_14573,N_15503);
and U17261 (N_17261,N_15580,N_14783);
and U17262 (N_17262,N_15144,N_15259);
nor U17263 (N_17263,N_15756,N_15239);
xor U17264 (N_17264,N_14017,N_14684);
and U17265 (N_17265,N_15806,N_15626);
or U17266 (N_17266,N_15619,N_15489);
or U17267 (N_17267,N_15991,N_14370);
xnor U17268 (N_17268,N_14223,N_15172);
and U17269 (N_17269,N_15717,N_15884);
or U17270 (N_17270,N_15493,N_14800);
nand U17271 (N_17271,N_15613,N_15671);
nand U17272 (N_17272,N_15860,N_14772);
nand U17273 (N_17273,N_14927,N_15090);
or U17274 (N_17274,N_14662,N_15266);
or U17275 (N_17275,N_15943,N_14600);
nand U17276 (N_17276,N_14228,N_15548);
and U17277 (N_17277,N_14640,N_15156);
nor U17278 (N_17278,N_14505,N_15113);
nand U17279 (N_17279,N_14022,N_15645);
xor U17280 (N_17280,N_14264,N_14095);
nand U17281 (N_17281,N_14934,N_14964);
or U17282 (N_17282,N_15897,N_14561);
nand U17283 (N_17283,N_15964,N_14163);
nor U17284 (N_17284,N_15459,N_15040);
and U17285 (N_17285,N_14931,N_14218);
or U17286 (N_17286,N_14513,N_15496);
nor U17287 (N_17287,N_15834,N_14908);
or U17288 (N_17288,N_15755,N_14938);
and U17289 (N_17289,N_14939,N_14691);
nand U17290 (N_17290,N_15473,N_14648);
or U17291 (N_17291,N_14058,N_15993);
nor U17292 (N_17292,N_15457,N_15265);
and U17293 (N_17293,N_15293,N_14694);
and U17294 (N_17294,N_15659,N_15886);
nor U17295 (N_17295,N_14446,N_15484);
nor U17296 (N_17296,N_15952,N_14152);
nand U17297 (N_17297,N_14922,N_14862);
xor U17298 (N_17298,N_14786,N_15541);
nor U17299 (N_17299,N_14305,N_15689);
or U17300 (N_17300,N_15154,N_14462);
or U17301 (N_17301,N_14013,N_14709);
nor U17302 (N_17302,N_14020,N_15438);
nor U17303 (N_17303,N_14506,N_15301);
or U17304 (N_17304,N_14887,N_14815);
nand U17305 (N_17305,N_15792,N_15385);
nand U17306 (N_17306,N_15716,N_14402);
nand U17307 (N_17307,N_14064,N_15862);
or U17308 (N_17308,N_14214,N_14011);
or U17309 (N_17309,N_14852,N_14930);
nand U17310 (N_17310,N_14705,N_15637);
nand U17311 (N_17311,N_14560,N_14071);
and U17312 (N_17312,N_14615,N_15013);
nand U17313 (N_17313,N_15801,N_14042);
nor U17314 (N_17314,N_14727,N_15396);
and U17315 (N_17315,N_14044,N_15738);
or U17316 (N_17316,N_14465,N_15401);
xor U17317 (N_17317,N_14430,N_14446);
nor U17318 (N_17318,N_15945,N_14350);
or U17319 (N_17319,N_14952,N_15770);
or U17320 (N_17320,N_15045,N_15707);
or U17321 (N_17321,N_15447,N_14794);
and U17322 (N_17322,N_15031,N_15474);
and U17323 (N_17323,N_15460,N_15439);
nand U17324 (N_17324,N_15228,N_15058);
and U17325 (N_17325,N_15722,N_15321);
nand U17326 (N_17326,N_15734,N_15243);
nor U17327 (N_17327,N_15888,N_14128);
xnor U17328 (N_17328,N_14082,N_15922);
xor U17329 (N_17329,N_14594,N_15880);
nand U17330 (N_17330,N_14716,N_14758);
nor U17331 (N_17331,N_15105,N_14595);
nand U17332 (N_17332,N_14490,N_14244);
nor U17333 (N_17333,N_15669,N_14221);
nor U17334 (N_17334,N_15435,N_15213);
nor U17335 (N_17335,N_14896,N_14909);
or U17336 (N_17336,N_14863,N_15569);
and U17337 (N_17337,N_15336,N_15175);
or U17338 (N_17338,N_15323,N_15079);
nor U17339 (N_17339,N_15462,N_14260);
or U17340 (N_17340,N_15038,N_15763);
nand U17341 (N_17341,N_14776,N_15954);
nand U17342 (N_17342,N_14399,N_14906);
nand U17343 (N_17343,N_14312,N_14576);
nand U17344 (N_17344,N_15263,N_15224);
and U17345 (N_17345,N_14160,N_14141);
nor U17346 (N_17346,N_14732,N_15031);
nor U17347 (N_17347,N_14737,N_14905);
or U17348 (N_17348,N_14204,N_15921);
nand U17349 (N_17349,N_14337,N_14114);
nand U17350 (N_17350,N_14096,N_15621);
nor U17351 (N_17351,N_14180,N_15696);
nand U17352 (N_17352,N_14758,N_14234);
or U17353 (N_17353,N_14800,N_15812);
and U17354 (N_17354,N_15648,N_14853);
or U17355 (N_17355,N_14579,N_15297);
nand U17356 (N_17356,N_14420,N_15209);
nor U17357 (N_17357,N_14726,N_14971);
and U17358 (N_17358,N_15717,N_15081);
or U17359 (N_17359,N_15388,N_15529);
or U17360 (N_17360,N_14537,N_14136);
nand U17361 (N_17361,N_14380,N_15530);
nand U17362 (N_17362,N_14484,N_15919);
or U17363 (N_17363,N_14350,N_15636);
nand U17364 (N_17364,N_15363,N_14340);
and U17365 (N_17365,N_15453,N_15468);
and U17366 (N_17366,N_14728,N_14703);
nor U17367 (N_17367,N_14802,N_14703);
or U17368 (N_17368,N_14347,N_15087);
nand U17369 (N_17369,N_14012,N_15653);
nor U17370 (N_17370,N_14212,N_14461);
nand U17371 (N_17371,N_14271,N_14257);
xor U17372 (N_17372,N_15679,N_15315);
nor U17373 (N_17373,N_15739,N_15919);
or U17374 (N_17374,N_15828,N_14586);
and U17375 (N_17375,N_14230,N_14075);
nand U17376 (N_17376,N_15605,N_15639);
nor U17377 (N_17377,N_15248,N_14584);
nand U17378 (N_17378,N_15308,N_14754);
xnor U17379 (N_17379,N_14808,N_14789);
nand U17380 (N_17380,N_14723,N_14963);
and U17381 (N_17381,N_15752,N_15204);
and U17382 (N_17382,N_15983,N_14718);
xor U17383 (N_17383,N_15432,N_15162);
or U17384 (N_17384,N_15858,N_15386);
or U17385 (N_17385,N_14984,N_15949);
and U17386 (N_17386,N_14734,N_15434);
nand U17387 (N_17387,N_15698,N_15046);
or U17388 (N_17388,N_14437,N_14166);
nor U17389 (N_17389,N_14901,N_15377);
or U17390 (N_17390,N_14650,N_14655);
nor U17391 (N_17391,N_14611,N_14948);
nand U17392 (N_17392,N_14770,N_15665);
xnor U17393 (N_17393,N_14651,N_15675);
nand U17394 (N_17394,N_14783,N_14070);
and U17395 (N_17395,N_15383,N_14593);
or U17396 (N_17396,N_15641,N_14000);
and U17397 (N_17397,N_15496,N_15006);
nand U17398 (N_17398,N_14687,N_14204);
nor U17399 (N_17399,N_14123,N_14049);
nor U17400 (N_17400,N_15290,N_14344);
or U17401 (N_17401,N_15494,N_14362);
nor U17402 (N_17402,N_14824,N_15375);
and U17403 (N_17403,N_14171,N_14295);
nand U17404 (N_17404,N_14887,N_15421);
nand U17405 (N_17405,N_15917,N_14483);
nor U17406 (N_17406,N_15103,N_14259);
nor U17407 (N_17407,N_14663,N_14995);
nand U17408 (N_17408,N_15972,N_14352);
nand U17409 (N_17409,N_15397,N_14615);
nand U17410 (N_17410,N_15006,N_15585);
nor U17411 (N_17411,N_15894,N_15203);
or U17412 (N_17412,N_15622,N_14168);
nor U17413 (N_17413,N_15970,N_14275);
or U17414 (N_17414,N_15952,N_14813);
xnor U17415 (N_17415,N_15066,N_15175);
or U17416 (N_17416,N_14015,N_14264);
and U17417 (N_17417,N_15950,N_15775);
and U17418 (N_17418,N_14754,N_14698);
or U17419 (N_17419,N_15045,N_14336);
nor U17420 (N_17420,N_15006,N_15364);
nor U17421 (N_17421,N_14537,N_15201);
nor U17422 (N_17422,N_14764,N_15207);
nor U17423 (N_17423,N_15194,N_15612);
nor U17424 (N_17424,N_14352,N_14050);
or U17425 (N_17425,N_14061,N_14413);
xnor U17426 (N_17426,N_14930,N_15532);
or U17427 (N_17427,N_15728,N_15981);
nand U17428 (N_17428,N_14736,N_15958);
nand U17429 (N_17429,N_14907,N_14860);
or U17430 (N_17430,N_14167,N_15134);
nor U17431 (N_17431,N_15321,N_15037);
and U17432 (N_17432,N_14340,N_15748);
nor U17433 (N_17433,N_15518,N_15461);
and U17434 (N_17434,N_14637,N_15924);
nand U17435 (N_17435,N_14721,N_15712);
or U17436 (N_17436,N_14285,N_15674);
nor U17437 (N_17437,N_14852,N_15853);
or U17438 (N_17438,N_14759,N_15530);
nand U17439 (N_17439,N_15304,N_14620);
or U17440 (N_17440,N_14201,N_15801);
or U17441 (N_17441,N_14674,N_15549);
xor U17442 (N_17442,N_14012,N_14537);
or U17443 (N_17443,N_14367,N_15407);
nand U17444 (N_17444,N_14224,N_14137);
nor U17445 (N_17445,N_15915,N_14986);
nand U17446 (N_17446,N_15582,N_14045);
xor U17447 (N_17447,N_15100,N_14151);
nand U17448 (N_17448,N_15249,N_15317);
nor U17449 (N_17449,N_15130,N_15491);
nor U17450 (N_17450,N_15160,N_14412);
or U17451 (N_17451,N_15990,N_14637);
or U17452 (N_17452,N_15168,N_14755);
and U17453 (N_17453,N_15156,N_14924);
nor U17454 (N_17454,N_15567,N_15663);
and U17455 (N_17455,N_15407,N_14215);
nor U17456 (N_17456,N_14402,N_15572);
and U17457 (N_17457,N_15884,N_14586);
nor U17458 (N_17458,N_14429,N_14408);
and U17459 (N_17459,N_14119,N_15535);
nand U17460 (N_17460,N_14341,N_15047);
nor U17461 (N_17461,N_14044,N_15088);
and U17462 (N_17462,N_14787,N_15978);
nor U17463 (N_17463,N_15508,N_15192);
or U17464 (N_17464,N_14289,N_14685);
nor U17465 (N_17465,N_15127,N_15025);
or U17466 (N_17466,N_15729,N_15202);
and U17467 (N_17467,N_15722,N_14181);
nor U17468 (N_17468,N_15753,N_14555);
xnor U17469 (N_17469,N_15300,N_15291);
or U17470 (N_17470,N_14354,N_15762);
or U17471 (N_17471,N_14499,N_14910);
nor U17472 (N_17472,N_14572,N_15580);
xnor U17473 (N_17473,N_15264,N_14975);
or U17474 (N_17474,N_15528,N_14052);
nand U17475 (N_17475,N_15876,N_15872);
and U17476 (N_17476,N_15292,N_14504);
or U17477 (N_17477,N_14578,N_15958);
or U17478 (N_17478,N_15131,N_14254);
and U17479 (N_17479,N_15605,N_15022);
nand U17480 (N_17480,N_15793,N_15395);
or U17481 (N_17481,N_15805,N_14046);
xnor U17482 (N_17482,N_14511,N_14985);
nand U17483 (N_17483,N_14992,N_15601);
or U17484 (N_17484,N_14406,N_15830);
nor U17485 (N_17485,N_14101,N_15980);
and U17486 (N_17486,N_14707,N_14504);
nor U17487 (N_17487,N_14300,N_14086);
nand U17488 (N_17488,N_14851,N_14089);
xor U17489 (N_17489,N_15036,N_14196);
nor U17490 (N_17490,N_14058,N_14888);
and U17491 (N_17491,N_14371,N_14095);
nand U17492 (N_17492,N_14403,N_14192);
nand U17493 (N_17493,N_14912,N_14833);
nor U17494 (N_17494,N_14625,N_15056);
or U17495 (N_17495,N_14852,N_15420);
and U17496 (N_17496,N_15224,N_15005);
and U17497 (N_17497,N_14128,N_14429);
nand U17498 (N_17498,N_14164,N_14862);
xnor U17499 (N_17499,N_14892,N_15738);
xor U17500 (N_17500,N_14501,N_15638);
nand U17501 (N_17501,N_15274,N_15154);
and U17502 (N_17502,N_15846,N_15482);
and U17503 (N_17503,N_15256,N_14606);
or U17504 (N_17504,N_15488,N_14833);
and U17505 (N_17505,N_14250,N_14882);
xnor U17506 (N_17506,N_14034,N_15484);
nor U17507 (N_17507,N_15982,N_15604);
or U17508 (N_17508,N_15214,N_15266);
and U17509 (N_17509,N_14234,N_14514);
xor U17510 (N_17510,N_14015,N_15778);
nor U17511 (N_17511,N_14135,N_14275);
nand U17512 (N_17512,N_15186,N_15280);
or U17513 (N_17513,N_15075,N_14249);
or U17514 (N_17514,N_15746,N_14735);
or U17515 (N_17515,N_14376,N_15325);
nand U17516 (N_17516,N_15161,N_14545);
nand U17517 (N_17517,N_15795,N_14433);
and U17518 (N_17518,N_15530,N_14112);
nand U17519 (N_17519,N_15529,N_15679);
or U17520 (N_17520,N_15618,N_14843);
and U17521 (N_17521,N_15617,N_15844);
nor U17522 (N_17522,N_14134,N_14408);
or U17523 (N_17523,N_14560,N_15630);
or U17524 (N_17524,N_14656,N_15114);
and U17525 (N_17525,N_14145,N_14596);
nor U17526 (N_17526,N_15623,N_14829);
nand U17527 (N_17527,N_14546,N_15259);
nor U17528 (N_17528,N_14300,N_14231);
nor U17529 (N_17529,N_15020,N_15977);
nand U17530 (N_17530,N_15330,N_14196);
nor U17531 (N_17531,N_14332,N_14110);
or U17532 (N_17532,N_15106,N_14080);
or U17533 (N_17533,N_15492,N_14017);
and U17534 (N_17534,N_15208,N_15925);
nor U17535 (N_17535,N_14156,N_15150);
nand U17536 (N_17536,N_15703,N_14291);
and U17537 (N_17537,N_14243,N_14853);
or U17538 (N_17538,N_15104,N_14731);
nor U17539 (N_17539,N_14155,N_14967);
and U17540 (N_17540,N_15428,N_15926);
nand U17541 (N_17541,N_14638,N_14917);
nand U17542 (N_17542,N_14901,N_14100);
or U17543 (N_17543,N_15882,N_14719);
nand U17544 (N_17544,N_15501,N_15443);
and U17545 (N_17545,N_15686,N_15436);
nor U17546 (N_17546,N_14627,N_14237);
xor U17547 (N_17547,N_15410,N_14303);
or U17548 (N_17548,N_15887,N_14804);
nand U17549 (N_17549,N_15851,N_15286);
nand U17550 (N_17550,N_15727,N_14756);
nand U17551 (N_17551,N_15892,N_14766);
and U17552 (N_17552,N_14321,N_15096);
and U17553 (N_17553,N_15771,N_14048);
nor U17554 (N_17554,N_15783,N_15071);
and U17555 (N_17555,N_15164,N_15655);
and U17556 (N_17556,N_14604,N_14328);
and U17557 (N_17557,N_15609,N_14418);
nor U17558 (N_17558,N_15700,N_15077);
nor U17559 (N_17559,N_15378,N_14932);
or U17560 (N_17560,N_15480,N_14330);
nand U17561 (N_17561,N_15876,N_14887);
nand U17562 (N_17562,N_14142,N_15946);
nand U17563 (N_17563,N_15452,N_14644);
or U17564 (N_17564,N_15478,N_14013);
nor U17565 (N_17565,N_14619,N_15256);
and U17566 (N_17566,N_15242,N_14788);
nand U17567 (N_17567,N_14449,N_15165);
nor U17568 (N_17568,N_15109,N_15517);
or U17569 (N_17569,N_14549,N_15963);
or U17570 (N_17570,N_14498,N_14984);
or U17571 (N_17571,N_15067,N_14901);
and U17572 (N_17572,N_14909,N_15101);
nand U17573 (N_17573,N_15180,N_15234);
and U17574 (N_17574,N_14211,N_14591);
and U17575 (N_17575,N_15609,N_14912);
nand U17576 (N_17576,N_14389,N_15541);
or U17577 (N_17577,N_15582,N_15920);
or U17578 (N_17578,N_15092,N_14245);
and U17579 (N_17579,N_14638,N_15870);
or U17580 (N_17580,N_15798,N_14117);
and U17581 (N_17581,N_14112,N_14771);
nor U17582 (N_17582,N_15527,N_14497);
or U17583 (N_17583,N_15033,N_15586);
xor U17584 (N_17584,N_14848,N_15150);
or U17585 (N_17585,N_14990,N_14482);
or U17586 (N_17586,N_15410,N_14821);
or U17587 (N_17587,N_15780,N_14338);
and U17588 (N_17588,N_15096,N_14552);
xnor U17589 (N_17589,N_14422,N_15684);
and U17590 (N_17590,N_15654,N_15943);
xor U17591 (N_17591,N_14582,N_15735);
and U17592 (N_17592,N_15192,N_15409);
nor U17593 (N_17593,N_14764,N_15741);
xnor U17594 (N_17594,N_15742,N_15665);
or U17595 (N_17595,N_15076,N_14919);
and U17596 (N_17596,N_14758,N_14663);
or U17597 (N_17597,N_15276,N_15572);
nand U17598 (N_17598,N_14045,N_15580);
nand U17599 (N_17599,N_14455,N_15458);
and U17600 (N_17600,N_15240,N_14107);
or U17601 (N_17601,N_15407,N_14657);
xnor U17602 (N_17602,N_14259,N_14769);
xor U17603 (N_17603,N_15936,N_15576);
and U17604 (N_17604,N_14991,N_15710);
and U17605 (N_17605,N_14103,N_15112);
and U17606 (N_17606,N_15983,N_15486);
or U17607 (N_17607,N_14127,N_14899);
nor U17608 (N_17608,N_15322,N_15245);
nand U17609 (N_17609,N_15931,N_15891);
and U17610 (N_17610,N_14445,N_14004);
nand U17611 (N_17611,N_15860,N_15149);
nand U17612 (N_17612,N_14102,N_14439);
or U17613 (N_17613,N_15183,N_14790);
nand U17614 (N_17614,N_15208,N_15109);
and U17615 (N_17615,N_15556,N_15679);
or U17616 (N_17616,N_15125,N_15406);
or U17617 (N_17617,N_14126,N_14643);
xnor U17618 (N_17618,N_14059,N_15691);
and U17619 (N_17619,N_15850,N_14559);
nor U17620 (N_17620,N_15196,N_15903);
and U17621 (N_17621,N_15116,N_15399);
xor U17622 (N_17622,N_14512,N_14056);
nor U17623 (N_17623,N_14120,N_14483);
nor U17624 (N_17624,N_15510,N_15748);
and U17625 (N_17625,N_15573,N_15888);
or U17626 (N_17626,N_15997,N_14176);
or U17627 (N_17627,N_15842,N_14833);
nor U17628 (N_17628,N_15702,N_15162);
nor U17629 (N_17629,N_15097,N_14053);
and U17630 (N_17630,N_14205,N_15145);
and U17631 (N_17631,N_14662,N_15811);
xor U17632 (N_17632,N_15550,N_15880);
xnor U17633 (N_17633,N_15336,N_15250);
nand U17634 (N_17634,N_15413,N_14952);
or U17635 (N_17635,N_15597,N_15776);
and U17636 (N_17636,N_15797,N_15862);
and U17637 (N_17637,N_15106,N_14668);
xor U17638 (N_17638,N_15131,N_15954);
or U17639 (N_17639,N_15650,N_15776);
nand U17640 (N_17640,N_15620,N_15746);
nor U17641 (N_17641,N_15863,N_15646);
nand U17642 (N_17642,N_15222,N_14932);
and U17643 (N_17643,N_15129,N_15288);
or U17644 (N_17644,N_14438,N_14231);
nand U17645 (N_17645,N_15762,N_15642);
nand U17646 (N_17646,N_14153,N_15332);
xnor U17647 (N_17647,N_14164,N_14435);
nand U17648 (N_17648,N_15984,N_15739);
xnor U17649 (N_17649,N_14256,N_15119);
nor U17650 (N_17650,N_14997,N_15707);
nor U17651 (N_17651,N_15149,N_14989);
nor U17652 (N_17652,N_15571,N_14305);
nor U17653 (N_17653,N_15487,N_15453);
nand U17654 (N_17654,N_14866,N_15397);
nand U17655 (N_17655,N_15778,N_15871);
xnor U17656 (N_17656,N_15578,N_14911);
or U17657 (N_17657,N_14806,N_15850);
and U17658 (N_17658,N_14306,N_14406);
or U17659 (N_17659,N_15711,N_14488);
nand U17660 (N_17660,N_14859,N_15050);
and U17661 (N_17661,N_14976,N_15839);
xnor U17662 (N_17662,N_14630,N_15380);
or U17663 (N_17663,N_14670,N_15550);
and U17664 (N_17664,N_14339,N_15848);
and U17665 (N_17665,N_15818,N_14857);
and U17666 (N_17666,N_14872,N_15071);
nand U17667 (N_17667,N_14456,N_14800);
xor U17668 (N_17668,N_15332,N_14640);
nand U17669 (N_17669,N_15159,N_15117);
and U17670 (N_17670,N_14578,N_14222);
nor U17671 (N_17671,N_15938,N_14116);
or U17672 (N_17672,N_15392,N_15060);
and U17673 (N_17673,N_15137,N_15352);
nand U17674 (N_17674,N_14631,N_14635);
xnor U17675 (N_17675,N_14590,N_15987);
and U17676 (N_17676,N_15542,N_15900);
or U17677 (N_17677,N_15107,N_15518);
and U17678 (N_17678,N_15830,N_15206);
xor U17679 (N_17679,N_15263,N_14567);
or U17680 (N_17680,N_15743,N_15903);
and U17681 (N_17681,N_15861,N_15835);
xnor U17682 (N_17682,N_15727,N_15375);
or U17683 (N_17683,N_15091,N_15886);
nor U17684 (N_17684,N_14174,N_15746);
xnor U17685 (N_17685,N_14027,N_14213);
and U17686 (N_17686,N_15061,N_14215);
nand U17687 (N_17687,N_15382,N_14055);
or U17688 (N_17688,N_14901,N_15701);
and U17689 (N_17689,N_15826,N_15540);
or U17690 (N_17690,N_14105,N_14858);
xor U17691 (N_17691,N_14253,N_14960);
nor U17692 (N_17692,N_15311,N_14968);
nand U17693 (N_17693,N_14320,N_14957);
and U17694 (N_17694,N_14909,N_15496);
nand U17695 (N_17695,N_14996,N_14676);
nand U17696 (N_17696,N_14044,N_15872);
xor U17697 (N_17697,N_14498,N_14225);
nor U17698 (N_17698,N_14586,N_14890);
or U17699 (N_17699,N_14881,N_15160);
or U17700 (N_17700,N_15640,N_15907);
xor U17701 (N_17701,N_15115,N_15787);
nand U17702 (N_17702,N_14486,N_15304);
xnor U17703 (N_17703,N_15390,N_14615);
nand U17704 (N_17704,N_15342,N_14575);
and U17705 (N_17705,N_14642,N_14624);
xor U17706 (N_17706,N_15714,N_14086);
nor U17707 (N_17707,N_14079,N_15782);
nand U17708 (N_17708,N_15672,N_14234);
and U17709 (N_17709,N_14748,N_14694);
or U17710 (N_17710,N_14712,N_15391);
nand U17711 (N_17711,N_14020,N_15844);
or U17712 (N_17712,N_14698,N_15089);
or U17713 (N_17713,N_14688,N_14015);
nor U17714 (N_17714,N_14403,N_14013);
nor U17715 (N_17715,N_14567,N_15800);
and U17716 (N_17716,N_14716,N_15977);
nand U17717 (N_17717,N_14412,N_14929);
and U17718 (N_17718,N_14881,N_14249);
nor U17719 (N_17719,N_14887,N_14730);
or U17720 (N_17720,N_15494,N_15380);
and U17721 (N_17721,N_15470,N_15797);
or U17722 (N_17722,N_14220,N_15218);
and U17723 (N_17723,N_14321,N_15761);
nand U17724 (N_17724,N_14972,N_15096);
or U17725 (N_17725,N_14160,N_15166);
or U17726 (N_17726,N_15644,N_14601);
and U17727 (N_17727,N_15663,N_14666);
and U17728 (N_17728,N_14283,N_15320);
nand U17729 (N_17729,N_14864,N_15689);
xnor U17730 (N_17730,N_15305,N_14627);
and U17731 (N_17731,N_15403,N_15307);
and U17732 (N_17732,N_15580,N_15718);
or U17733 (N_17733,N_15941,N_15713);
or U17734 (N_17734,N_15498,N_14445);
or U17735 (N_17735,N_15394,N_15739);
or U17736 (N_17736,N_15925,N_15108);
and U17737 (N_17737,N_14171,N_14252);
or U17738 (N_17738,N_15074,N_15348);
nand U17739 (N_17739,N_14163,N_14547);
nand U17740 (N_17740,N_15033,N_15548);
nand U17741 (N_17741,N_14251,N_15786);
and U17742 (N_17742,N_14821,N_15690);
or U17743 (N_17743,N_15545,N_14863);
nand U17744 (N_17744,N_14929,N_15367);
or U17745 (N_17745,N_15678,N_14153);
nand U17746 (N_17746,N_14602,N_14759);
nand U17747 (N_17747,N_15435,N_15241);
nor U17748 (N_17748,N_14064,N_14568);
and U17749 (N_17749,N_15305,N_14001);
nor U17750 (N_17750,N_14830,N_14289);
nand U17751 (N_17751,N_14572,N_14432);
nor U17752 (N_17752,N_14258,N_15207);
nand U17753 (N_17753,N_14502,N_14375);
and U17754 (N_17754,N_15794,N_14159);
or U17755 (N_17755,N_14936,N_15598);
nor U17756 (N_17756,N_14659,N_15901);
nor U17757 (N_17757,N_15290,N_15642);
or U17758 (N_17758,N_15983,N_15383);
nand U17759 (N_17759,N_15826,N_14455);
and U17760 (N_17760,N_14409,N_14413);
or U17761 (N_17761,N_15549,N_15333);
and U17762 (N_17762,N_15446,N_15536);
nand U17763 (N_17763,N_14428,N_15854);
or U17764 (N_17764,N_14477,N_15463);
or U17765 (N_17765,N_15609,N_15145);
nand U17766 (N_17766,N_14727,N_15634);
nand U17767 (N_17767,N_14816,N_14633);
and U17768 (N_17768,N_15528,N_14629);
nand U17769 (N_17769,N_14371,N_14575);
nand U17770 (N_17770,N_14245,N_15622);
nor U17771 (N_17771,N_14077,N_15827);
or U17772 (N_17772,N_14107,N_14076);
nor U17773 (N_17773,N_14908,N_14134);
nand U17774 (N_17774,N_15172,N_14616);
or U17775 (N_17775,N_14029,N_15828);
nand U17776 (N_17776,N_14954,N_14318);
nand U17777 (N_17777,N_14466,N_15043);
nor U17778 (N_17778,N_15680,N_14660);
nor U17779 (N_17779,N_14089,N_14064);
nor U17780 (N_17780,N_15124,N_15047);
nor U17781 (N_17781,N_15677,N_14965);
and U17782 (N_17782,N_14377,N_14066);
nand U17783 (N_17783,N_14236,N_14355);
nand U17784 (N_17784,N_14770,N_14104);
or U17785 (N_17785,N_14957,N_15813);
nand U17786 (N_17786,N_14188,N_15000);
and U17787 (N_17787,N_15732,N_14734);
nor U17788 (N_17788,N_15576,N_14226);
xnor U17789 (N_17789,N_15672,N_14499);
nand U17790 (N_17790,N_15427,N_14703);
nor U17791 (N_17791,N_14522,N_14292);
nor U17792 (N_17792,N_14383,N_14713);
nand U17793 (N_17793,N_14030,N_14249);
or U17794 (N_17794,N_15862,N_14345);
and U17795 (N_17795,N_14259,N_14295);
or U17796 (N_17796,N_14584,N_15541);
nand U17797 (N_17797,N_14079,N_14949);
and U17798 (N_17798,N_15054,N_14571);
nand U17799 (N_17799,N_14434,N_15853);
or U17800 (N_17800,N_15719,N_15183);
and U17801 (N_17801,N_15428,N_14809);
xnor U17802 (N_17802,N_14026,N_14854);
nand U17803 (N_17803,N_15347,N_14066);
or U17804 (N_17804,N_15487,N_14057);
or U17805 (N_17805,N_14935,N_14301);
and U17806 (N_17806,N_15278,N_14287);
or U17807 (N_17807,N_15282,N_15598);
nor U17808 (N_17808,N_14504,N_14199);
and U17809 (N_17809,N_14320,N_14424);
nor U17810 (N_17810,N_15175,N_14659);
and U17811 (N_17811,N_15876,N_14318);
nor U17812 (N_17812,N_15759,N_15732);
and U17813 (N_17813,N_15156,N_14674);
xnor U17814 (N_17814,N_15775,N_15041);
nor U17815 (N_17815,N_15973,N_15923);
and U17816 (N_17816,N_14198,N_15150);
or U17817 (N_17817,N_15065,N_14191);
or U17818 (N_17818,N_14091,N_15512);
or U17819 (N_17819,N_14870,N_14882);
xor U17820 (N_17820,N_15072,N_14372);
nor U17821 (N_17821,N_14332,N_15047);
or U17822 (N_17822,N_15441,N_14930);
or U17823 (N_17823,N_14950,N_15591);
or U17824 (N_17824,N_14678,N_15497);
xnor U17825 (N_17825,N_14174,N_15363);
nand U17826 (N_17826,N_15333,N_14432);
nand U17827 (N_17827,N_15236,N_15523);
nor U17828 (N_17828,N_15074,N_15617);
or U17829 (N_17829,N_15894,N_15212);
or U17830 (N_17830,N_15833,N_14568);
xor U17831 (N_17831,N_14197,N_15066);
xor U17832 (N_17832,N_15966,N_15061);
and U17833 (N_17833,N_15243,N_14725);
nor U17834 (N_17834,N_15424,N_14971);
or U17835 (N_17835,N_15039,N_15204);
and U17836 (N_17836,N_14862,N_15146);
xor U17837 (N_17837,N_14764,N_15736);
nand U17838 (N_17838,N_14457,N_14423);
or U17839 (N_17839,N_14230,N_14602);
nand U17840 (N_17840,N_14968,N_14021);
and U17841 (N_17841,N_15449,N_15376);
xor U17842 (N_17842,N_14646,N_15761);
xnor U17843 (N_17843,N_15010,N_14628);
and U17844 (N_17844,N_15198,N_14088);
or U17845 (N_17845,N_15603,N_15388);
or U17846 (N_17846,N_15936,N_14197);
nor U17847 (N_17847,N_15316,N_14487);
xor U17848 (N_17848,N_14701,N_15330);
xnor U17849 (N_17849,N_15832,N_15229);
nor U17850 (N_17850,N_14686,N_14232);
and U17851 (N_17851,N_14160,N_14644);
and U17852 (N_17852,N_15046,N_15458);
and U17853 (N_17853,N_15222,N_15426);
nand U17854 (N_17854,N_14194,N_15712);
nand U17855 (N_17855,N_15312,N_15067);
nor U17856 (N_17856,N_15661,N_14340);
or U17857 (N_17857,N_15466,N_14176);
and U17858 (N_17858,N_15861,N_14315);
nor U17859 (N_17859,N_14456,N_15122);
nand U17860 (N_17860,N_15546,N_15765);
nor U17861 (N_17861,N_15239,N_14273);
xor U17862 (N_17862,N_15013,N_14086);
nand U17863 (N_17863,N_15376,N_14571);
and U17864 (N_17864,N_14839,N_14512);
and U17865 (N_17865,N_15597,N_15497);
or U17866 (N_17866,N_14624,N_15439);
or U17867 (N_17867,N_15085,N_14987);
and U17868 (N_17868,N_14730,N_15405);
or U17869 (N_17869,N_15419,N_14245);
nand U17870 (N_17870,N_14589,N_15516);
and U17871 (N_17871,N_15747,N_14120);
xor U17872 (N_17872,N_14807,N_15455);
or U17873 (N_17873,N_14088,N_14646);
and U17874 (N_17874,N_14291,N_14112);
nor U17875 (N_17875,N_15546,N_15349);
nand U17876 (N_17876,N_14995,N_14423);
or U17877 (N_17877,N_14380,N_15558);
nand U17878 (N_17878,N_15417,N_14488);
and U17879 (N_17879,N_14682,N_15379);
or U17880 (N_17880,N_14636,N_15791);
and U17881 (N_17881,N_15713,N_15754);
or U17882 (N_17882,N_15517,N_14610);
nand U17883 (N_17883,N_14748,N_15834);
or U17884 (N_17884,N_15025,N_14296);
xnor U17885 (N_17885,N_14057,N_14154);
and U17886 (N_17886,N_15124,N_14967);
nor U17887 (N_17887,N_15968,N_14483);
nand U17888 (N_17888,N_14289,N_14496);
or U17889 (N_17889,N_15865,N_14237);
or U17890 (N_17890,N_15076,N_14832);
nor U17891 (N_17891,N_15342,N_14321);
and U17892 (N_17892,N_15513,N_14289);
and U17893 (N_17893,N_15144,N_14410);
nand U17894 (N_17894,N_15846,N_14597);
nor U17895 (N_17895,N_14114,N_15434);
xnor U17896 (N_17896,N_15115,N_14518);
xnor U17897 (N_17897,N_14301,N_14974);
nor U17898 (N_17898,N_15577,N_15384);
or U17899 (N_17899,N_14966,N_14956);
nand U17900 (N_17900,N_14103,N_15594);
or U17901 (N_17901,N_15789,N_14249);
nand U17902 (N_17902,N_14963,N_14607);
nor U17903 (N_17903,N_15643,N_14900);
nand U17904 (N_17904,N_15969,N_15348);
and U17905 (N_17905,N_15215,N_15963);
nand U17906 (N_17906,N_14333,N_15410);
nor U17907 (N_17907,N_15234,N_14014);
nand U17908 (N_17908,N_14736,N_14017);
nand U17909 (N_17909,N_14871,N_14961);
nand U17910 (N_17910,N_14319,N_15787);
nor U17911 (N_17911,N_15882,N_14619);
or U17912 (N_17912,N_15827,N_15062);
xor U17913 (N_17913,N_15020,N_14974);
and U17914 (N_17914,N_15230,N_15434);
nor U17915 (N_17915,N_14377,N_14693);
or U17916 (N_17916,N_15488,N_15809);
nand U17917 (N_17917,N_14712,N_14222);
and U17918 (N_17918,N_15636,N_14765);
xnor U17919 (N_17919,N_14638,N_14662);
and U17920 (N_17920,N_14683,N_15408);
or U17921 (N_17921,N_14790,N_14907);
nor U17922 (N_17922,N_15185,N_15388);
nor U17923 (N_17923,N_14045,N_15584);
nor U17924 (N_17924,N_15014,N_14128);
nand U17925 (N_17925,N_14177,N_14938);
xor U17926 (N_17926,N_14980,N_14436);
nand U17927 (N_17927,N_14741,N_14972);
nand U17928 (N_17928,N_15315,N_14218);
and U17929 (N_17929,N_15254,N_14122);
and U17930 (N_17930,N_14525,N_14177);
nand U17931 (N_17931,N_15239,N_15099);
and U17932 (N_17932,N_14021,N_14411);
nor U17933 (N_17933,N_15442,N_14193);
nand U17934 (N_17934,N_15925,N_14854);
nor U17935 (N_17935,N_14321,N_15218);
nand U17936 (N_17936,N_15504,N_15737);
nor U17937 (N_17937,N_14594,N_14497);
nand U17938 (N_17938,N_15630,N_14540);
or U17939 (N_17939,N_15228,N_15640);
or U17940 (N_17940,N_15984,N_15693);
nor U17941 (N_17941,N_15919,N_15060);
nand U17942 (N_17942,N_15772,N_14901);
nor U17943 (N_17943,N_15332,N_14764);
or U17944 (N_17944,N_14771,N_14339);
nor U17945 (N_17945,N_14933,N_14305);
and U17946 (N_17946,N_14919,N_15713);
nor U17947 (N_17947,N_14846,N_15743);
nand U17948 (N_17948,N_15115,N_14897);
nor U17949 (N_17949,N_15430,N_15820);
or U17950 (N_17950,N_15597,N_14930);
or U17951 (N_17951,N_15415,N_14835);
and U17952 (N_17952,N_14662,N_14014);
and U17953 (N_17953,N_15074,N_14038);
or U17954 (N_17954,N_15858,N_14872);
nand U17955 (N_17955,N_15963,N_15123);
or U17956 (N_17956,N_14203,N_14712);
nor U17957 (N_17957,N_15087,N_15802);
nand U17958 (N_17958,N_15365,N_14776);
or U17959 (N_17959,N_15585,N_15014);
nor U17960 (N_17960,N_14084,N_15770);
nor U17961 (N_17961,N_14805,N_14801);
and U17962 (N_17962,N_15587,N_14826);
nand U17963 (N_17963,N_15254,N_14887);
and U17964 (N_17964,N_14224,N_14207);
xnor U17965 (N_17965,N_14569,N_15504);
nand U17966 (N_17966,N_15280,N_15301);
nand U17967 (N_17967,N_14790,N_14118);
nor U17968 (N_17968,N_15121,N_15790);
xnor U17969 (N_17969,N_14725,N_15010);
and U17970 (N_17970,N_14697,N_15782);
nor U17971 (N_17971,N_14532,N_15497);
nand U17972 (N_17972,N_15329,N_14546);
nand U17973 (N_17973,N_14650,N_15176);
nand U17974 (N_17974,N_14134,N_15528);
xnor U17975 (N_17975,N_15649,N_15340);
and U17976 (N_17976,N_14318,N_14127);
xor U17977 (N_17977,N_14928,N_15222);
nand U17978 (N_17978,N_14782,N_14731);
and U17979 (N_17979,N_14188,N_14632);
xnor U17980 (N_17980,N_15259,N_15812);
nand U17981 (N_17981,N_15866,N_14875);
or U17982 (N_17982,N_15039,N_15518);
and U17983 (N_17983,N_15640,N_15169);
and U17984 (N_17984,N_14511,N_15527);
and U17985 (N_17985,N_15390,N_15480);
nor U17986 (N_17986,N_14595,N_14579);
nor U17987 (N_17987,N_15258,N_14701);
nor U17988 (N_17988,N_15152,N_15448);
and U17989 (N_17989,N_15033,N_15902);
xor U17990 (N_17990,N_15191,N_15700);
or U17991 (N_17991,N_15066,N_14243);
and U17992 (N_17992,N_14400,N_15383);
xnor U17993 (N_17993,N_14885,N_14778);
or U17994 (N_17994,N_14134,N_14874);
nor U17995 (N_17995,N_14390,N_14363);
or U17996 (N_17996,N_14917,N_14874);
nor U17997 (N_17997,N_15216,N_14775);
nor U17998 (N_17998,N_15453,N_14595);
or U17999 (N_17999,N_15666,N_15394);
and U18000 (N_18000,N_16621,N_17354);
and U18001 (N_18001,N_17946,N_17811);
or U18002 (N_18002,N_16969,N_17311);
nand U18003 (N_18003,N_16538,N_16527);
nor U18004 (N_18004,N_16406,N_17225);
or U18005 (N_18005,N_17813,N_16235);
or U18006 (N_18006,N_16313,N_16619);
or U18007 (N_18007,N_16022,N_16351);
nand U18008 (N_18008,N_17032,N_17065);
and U18009 (N_18009,N_16506,N_16526);
and U18010 (N_18010,N_16257,N_17949);
or U18011 (N_18011,N_16971,N_17133);
and U18012 (N_18012,N_17304,N_16587);
xor U18013 (N_18013,N_17875,N_16123);
xnor U18014 (N_18014,N_17210,N_16599);
nand U18015 (N_18015,N_16845,N_16477);
or U18016 (N_18016,N_17978,N_17351);
or U18017 (N_18017,N_16899,N_16055);
nand U18018 (N_18018,N_17816,N_16069);
nand U18019 (N_18019,N_16705,N_16590);
and U18020 (N_18020,N_16081,N_16516);
or U18021 (N_18021,N_16226,N_16160);
and U18022 (N_18022,N_16949,N_16015);
nand U18023 (N_18023,N_16448,N_17888);
nor U18024 (N_18024,N_16132,N_17766);
nor U18025 (N_18025,N_17387,N_17879);
nand U18026 (N_18026,N_16445,N_17873);
nand U18027 (N_18027,N_16211,N_17805);
xor U18028 (N_18028,N_17395,N_17736);
or U18029 (N_18029,N_16286,N_17837);
nor U18030 (N_18030,N_17798,N_17625);
and U18031 (N_18031,N_16084,N_16752);
and U18032 (N_18032,N_17907,N_17493);
nand U18033 (N_18033,N_16467,N_17179);
nand U18034 (N_18034,N_17100,N_16718);
nor U18035 (N_18035,N_17572,N_16732);
xnor U18036 (N_18036,N_16058,N_16551);
and U18037 (N_18037,N_17325,N_16546);
or U18038 (N_18038,N_16871,N_17479);
and U18039 (N_18039,N_16418,N_16793);
nor U18040 (N_18040,N_17601,N_17668);
nand U18041 (N_18041,N_16288,N_16558);
nor U18042 (N_18042,N_16903,N_16495);
xnor U18043 (N_18043,N_16159,N_16509);
nor U18044 (N_18044,N_16016,N_16561);
and U18045 (N_18045,N_17147,N_17373);
and U18046 (N_18046,N_16644,N_16067);
and U18047 (N_18047,N_17633,N_17347);
or U18048 (N_18048,N_16011,N_17629);
nor U18049 (N_18049,N_17326,N_16580);
nand U18050 (N_18050,N_16152,N_17795);
nor U18051 (N_18051,N_16106,N_16236);
nor U18052 (N_18052,N_17704,N_16353);
nor U18053 (N_18053,N_17700,N_16191);
nand U18054 (N_18054,N_16733,N_17081);
nand U18055 (N_18055,N_17198,N_16806);
and U18056 (N_18056,N_17546,N_16839);
nand U18057 (N_18057,N_16396,N_16966);
nand U18058 (N_18058,N_17144,N_16409);
and U18059 (N_18059,N_16428,N_17063);
and U18060 (N_18060,N_16659,N_17696);
nand U18061 (N_18061,N_17787,N_17836);
and U18062 (N_18062,N_16175,N_17243);
xor U18063 (N_18063,N_16959,N_16988);
nand U18064 (N_18064,N_16884,N_17323);
or U18065 (N_18065,N_16105,N_17567);
or U18066 (N_18066,N_16151,N_16505);
or U18067 (N_18067,N_17404,N_16374);
xnor U18068 (N_18068,N_17454,N_17550);
and U18069 (N_18069,N_16332,N_17080);
and U18070 (N_18070,N_17592,N_17206);
nand U18071 (N_18071,N_17060,N_16260);
and U18072 (N_18072,N_16860,N_17173);
nor U18073 (N_18073,N_16715,N_17061);
xor U18074 (N_18074,N_17374,N_16673);
nand U18075 (N_18075,N_17077,N_17064);
and U18076 (N_18076,N_16810,N_17468);
and U18077 (N_18077,N_16277,N_17259);
nand U18078 (N_18078,N_17526,N_17918);
and U18079 (N_18079,N_16688,N_16869);
or U18080 (N_18080,N_16660,N_16820);
nor U18081 (N_18081,N_16711,N_17617);
nand U18082 (N_18082,N_17528,N_17934);
xnor U18083 (N_18083,N_16970,N_17832);
or U18084 (N_18084,N_16861,N_17130);
xnor U18085 (N_18085,N_17220,N_17166);
nand U18086 (N_18086,N_17000,N_16821);
nand U18087 (N_18087,N_17285,N_16847);
nand U18088 (N_18088,N_16642,N_16072);
nor U18089 (N_18089,N_17038,N_16179);
and U18090 (N_18090,N_16926,N_17585);
and U18091 (N_18091,N_17380,N_17737);
nor U18092 (N_18092,N_17009,N_17486);
nand U18093 (N_18093,N_17040,N_17959);
nor U18094 (N_18094,N_17103,N_16675);
or U18095 (N_18095,N_16734,N_17997);
nand U18096 (N_18096,N_17899,N_16371);
and U18097 (N_18097,N_16301,N_17525);
xnor U18098 (N_18098,N_16663,N_16932);
or U18099 (N_18099,N_17134,N_16744);
nand U18100 (N_18100,N_17093,N_16633);
and U18101 (N_18101,N_17726,N_17405);
nand U18102 (N_18102,N_17257,N_16457);
or U18103 (N_18103,N_16864,N_17624);
nand U18104 (N_18104,N_16309,N_17803);
nor U18105 (N_18105,N_16000,N_17970);
or U18106 (N_18106,N_17860,N_17738);
and U18107 (N_18107,N_16610,N_16798);
nor U18108 (N_18108,N_16762,N_17490);
and U18109 (N_18109,N_17375,N_17286);
nand U18110 (N_18110,N_16857,N_17903);
nor U18111 (N_18111,N_17070,N_16001);
nor U18112 (N_18112,N_17036,N_16426);
nor U18113 (N_18113,N_17841,N_17217);
xnor U18114 (N_18114,N_16608,N_17194);
and U18115 (N_18115,N_17322,N_17654);
nand U18116 (N_18116,N_17916,N_16614);
nor U18117 (N_18117,N_16087,N_17400);
or U18118 (N_18118,N_17928,N_16240);
nand U18119 (N_18119,N_17132,N_16367);
and U18120 (N_18120,N_17932,N_17341);
nor U18121 (N_18121,N_16483,N_16611);
and U18122 (N_18122,N_17510,N_17850);
nor U18123 (N_18123,N_17437,N_16153);
or U18124 (N_18124,N_17974,N_16440);
nand U18125 (N_18125,N_16343,N_17492);
and U18126 (N_18126,N_16287,N_16623);
nor U18127 (N_18127,N_17261,N_16243);
nand U18128 (N_18128,N_17889,N_17951);
or U18129 (N_18129,N_16756,N_16267);
and U18130 (N_18130,N_17174,N_16746);
and U18131 (N_18131,N_17947,N_16263);
nor U18132 (N_18132,N_17535,N_16731);
nand U18133 (N_18133,N_16612,N_16843);
and U18134 (N_18134,N_16816,N_16555);
and U18135 (N_18135,N_16080,N_17457);
nand U18136 (N_18136,N_17785,N_16462);
nand U18137 (N_18137,N_16995,N_17289);
nand U18138 (N_18138,N_16485,N_17744);
and U18139 (N_18139,N_16796,N_17845);
and U18140 (N_18140,N_16737,N_17965);
or U18141 (N_18141,N_16233,N_16888);
or U18142 (N_18142,N_17681,N_16355);
nor U18143 (N_18143,N_16817,N_16269);
nor U18144 (N_18144,N_17044,N_17478);
or U18145 (N_18145,N_16473,N_16964);
and U18146 (N_18146,N_16197,N_17610);
nand U18147 (N_18147,N_16522,N_17104);
nand U18148 (N_18148,N_17623,N_16951);
nor U18149 (N_18149,N_16136,N_17491);
xnor U18150 (N_18150,N_16024,N_17794);
nand U18151 (N_18151,N_16183,N_17033);
nor U18152 (N_18152,N_17301,N_16169);
or U18153 (N_18153,N_17135,N_16361);
and U18154 (N_18154,N_16767,N_17877);
and U18155 (N_18155,N_17588,N_16992);
or U18156 (N_18156,N_16478,N_17871);
or U18157 (N_18157,N_16248,N_17500);
nand U18158 (N_18158,N_17205,N_16830);
or U18159 (N_18159,N_16382,N_17338);
and U18160 (N_18160,N_17458,N_17267);
and U18161 (N_18161,N_17188,N_16866);
or U18162 (N_18162,N_17848,N_17838);
nor U18163 (N_18163,N_16071,N_16177);
nand U18164 (N_18164,N_16395,N_17112);
and U18165 (N_18165,N_16874,N_17919);
and U18166 (N_18166,N_17977,N_17117);
and U18167 (N_18167,N_16126,N_16196);
or U18168 (N_18168,N_16962,N_16828);
or U18169 (N_18169,N_16963,N_17141);
or U18170 (N_18170,N_17950,N_16381);
nand U18171 (N_18171,N_16968,N_16563);
and U18172 (N_18172,N_17644,N_16771);
nand U18173 (N_18173,N_16760,N_17534);
or U18174 (N_18174,N_16424,N_17808);
or U18175 (N_18175,N_17663,N_17756);
nor U18176 (N_18176,N_17319,N_17584);
nand U18177 (N_18177,N_16511,N_16616);
or U18178 (N_18178,N_16695,N_16836);
nor U18179 (N_18179,N_17772,N_16475);
and U18180 (N_18180,N_16609,N_16782);
nand U18181 (N_18181,N_17670,N_16981);
nor U18182 (N_18182,N_17758,N_17449);
nor U18183 (N_18183,N_16928,N_16685);
xnor U18184 (N_18184,N_16799,N_16157);
and U18185 (N_18185,N_16986,N_16348);
or U18186 (N_18186,N_17433,N_17391);
and U18187 (N_18187,N_16973,N_17591);
or U18188 (N_18188,N_17569,N_16772);
nand U18189 (N_18189,N_17968,N_16765);
nand U18190 (N_18190,N_17581,N_16867);
or U18191 (N_18191,N_17900,N_16579);
nand U18192 (N_18192,N_16524,N_16111);
nor U18193 (N_18193,N_17401,N_17779);
nor U18194 (N_18194,N_17632,N_16013);
or U18195 (N_18195,N_17752,N_17393);
and U18196 (N_18196,N_16434,N_16242);
or U18197 (N_18197,N_16541,N_17709);
and U18198 (N_18198,N_17332,N_17872);
or U18199 (N_18199,N_16238,N_16911);
and U18200 (N_18200,N_16094,N_17605);
nor U18201 (N_18201,N_17788,N_17005);
nand U18202 (N_18202,N_17991,N_17138);
nor U18203 (N_18203,N_16164,N_16496);
nand U18204 (N_18204,N_16914,N_17830);
and U18205 (N_18205,N_16597,N_17441);
nand U18206 (N_18206,N_16728,N_16007);
nor U18207 (N_18207,N_16076,N_16005);
nand U18208 (N_18208,N_16594,N_16578);
or U18209 (N_18209,N_16125,N_16996);
nand U18210 (N_18210,N_16295,N_17396);
nand U18211 (N_18211,N_16826,N_16559);
or U18212 (N_18212,N_16491,N_16221);
nor U18213 (N_18213,N_16209,N_16002);
and U18214 (N_18214,N_16178,N_16622);
or U18215 (N_18215,N_17762,N_17314);
or U18216 (N_18216,N_17673,N_16430);
and U18217 (N_18217,N_17204,N_17980);
and U18218 (N_18218,N_16170,N_16118);
or U18219 (N_18219,N_16676,N_17887);
nor U18220 (N_18220,N_17321,N_16003);
xor U18221 (N_18221,N_16965,N_17429);
and U18222 (N_18222,N_17678,N_17570);
or U18223 (N_18223,N_16827,N_17796);
or U18224 (N_18224,N_17662,N_16437);
or U18225 (N_18225,N_16513,N_16850);
xor U18226 (N_18226,N_16831,N_16730);
or U18227 (N_18227,N_17814,N_17034);
and U18228 (N_18228,N_17935,N_17690);
nand U18229 (N_18229,N_16444,N_16185);
or U18230 (N_18230,N_17529,N_16455);
xor U18231 (N_18231,N_17990,N_17313);
nor U18232 (N_18232,N_17833,N_17041);
or U18233 (N_18233,N_17810,N_17518);
nor U18234 (N_18234,N_16312,N_17541);
and U18235 (N_18235,N_17418,N_17818);
or U18236 (N_18236,N_16070,N_16726);
nor U18237 (N_18237,N_16905,N_17360);
nor U18238 (N_18238,N_16740,N_16357);
nor U18239 (N_18239,N_17003,N_17672);
and U18240 (N_18240,N_17784,N_16412);
nor U18241 (N_18241,N_17770,N_16637);
or U18242 (N_18242,N_17119,N_17504);
and U18243 (N_18243,N_17114,N_16502);
nand U18244 (N_18244,N_16484,N_17998);
xor U18245 (N_18245,N_17058,N_16630);
nor U18246 (N_18246,N_17544,N_16285);
or U18247 (N_18247,N_16163,N_17209);
and U18248 (N_18248,N_17767,N_16219);
or U18249 (N_18249,N_16341,N_16605);
nor U18250 (N_18250,N_17923,N_17022);
nand U18251 (N_18251,N_16413,N_17215);
nor U18252 (N_18252,N_16275,N_17240);
nand U18253 (N_18253,N_16499,N_17501);
or U18254 (N_18254,N_16150,N_17461);
nand U18255 (N_18255,N_17964,N_17634);
xor U18256 (N_18256,N_16112,N_16829);
and U18257 (N_18257,N_16133,N_16528);
nand U18258 (N_18258,N_16998,N_16227);
or U18259 (N_18259,N_17929,N_17576);
and U18260 (N_18260,N_16489,N_16729);
and U18261 (N_18261,N_17381,N_16408);
nand U18262 (N_18262,N_17503,N_17187);
or U18263 (N_18263,N_16043,N_16165);
or U18264 (N_18264,N_16942,N_17489);
nor U18265 (N_18265,N_16432,N_16463);
nand U18266 (N_18266,N_17336,N_16683);
or U18267 (N_18267,N_17012,N_16977);
nor U18268 (N_18268,N_16975,N_17986);
nand U18269 (N_18269,N_16140,N_17427);
nor U18270 (N_18270,N_17732,N_16936);
or U18271 (N_18271,N_16727,N_16337);
or U18272 (N_18272,N_17720,N_16701);
nand U18273 (N_18273,N_17880,N_16379);
xor U18274 (N_18274,N_17078,N_16270);
or U18275 (N_18275,N_17940,N_16745);
nor U18276 (N_18276,N_16725,N_17771);
or U18277 (N_18277,N_16751,N_16791);
xnor U18278 (N_18278,N_16201,N_16634);
nand U18279 (N_18279,N_16804,N_16738);
nor U18280 (N_18280,N_17902,N_16482);
and U18281 (N_18281,N_17214,N_17106);
xnor U18282 (N_18282,N_16237,N_17254);
nand U18283 (N_18283,N_17498,N_17255);
and U18284 (N_18284,N_17665,N_16019);
or U18285 (N_18285,N_17708,N_17062);
xor U18286 (N_18286,N_17410,N_16814);
and U18287 (N_18287,N_17494,N_17999);
or U18288 (N_18288,N_17515,N_17046);
and U18289 (N_18289,N_17120,N_16508);
and U18290 (N_18290,N_16655,N_17713);
and U18291 (N_18291,N_16638,N_17506);
xor U18292 (N_18292,N_17430,N_17777);
and U18293 (N_18293,N_17712,N_17780);
xor U18294 (N_18294,N_16360,N_17278);
or U18295 (N_18295,N_16576,N_17088);
nand U18296 (N_18296,N_17698,N_16758);
nor U18297 (N_18297,N_17552,N_16088);
nand U18298 (N_18298,N_17786,N_17972);
nand U18299 (N_18299,N_16537,N_16927);
nor U18300 (N_18300,N_17893,N_17340);
and U18301 (N_18301,N_17912,N_17438);
nand U18302 (N_18302,N_16060,N_16661);
and U18303 (N_18303,N_17072,N_16639);
nand U18304 (N_18304,N_17024,N_16114);
or U18305 (N_18305,N_17943,N_16452);
or U18306 (N_18306,N_17042,N_17357);
and U18307 (N_18307,N_16754,N_16419);
nor U18308 (N_18308,N_16389,N_16808);
nor U18309 (N_18309,N_16465,N_16856);
nand U18310 (N_18310,N_16581,N_17109);
nor U18311 (N_18311,N_16693,N_16410);
or U18312 (N_18312,N_16093,N_17442);
xor U18313 (N_18313,N_16443,N_17399);
nand U18314 (N_18314,N_16887,N_17091);
or U18315 (N_18315,N_16224,N_16636);
nor U18316 (N_18316,N_16770,N_17731);
and U18317 (N_18317,N_17327,N_16356);
and U18318 (N_18318,N_17957,N_17763);
and U18319 (N_18319,N_17342,N_16672);
nor U18320 (N_18320,N_16886,N_17260);
or U18321 (N_18321,N_17006,N_16848);
or U18322 (N_18322,N_16214,N_16607);
or U18323 (N_18323,N_16876,N_16784);
nand U18324 (N_18324,N_16451,N_16459);
nor U18325 (N_18325,N_17536,N_16124);
nor U18326 (N_18326,N_17343,N_16722);
nor U18327 (N_18327,N_16469,N_17435);
nor U18328 (N_18328,N_16865,N_17746);
or U18329 (N_18329,N_17791,N_16934);
or U18330 (N_18330,N_17010,N_16033);
and U18331 (N_18331,N_16853,N_16121);
nand U18332 (N_18332,N_17684,N_17013);
xor U18333 (N_18333,N_17637,N_16323);
nor U18334 (N_18334,N_16895,N_16891);
xor U18335 (N_18335,N_16340,N_16023);
and U18336 (N_18336,N_17178,N_16773);
or U18337 (N_18337,N_17249,N_16769);
nor U18338 (N_18338,N_16498,N_17250);
and U18339 (N_18339,N_17370,N_16249);
nor U18340 (N_18340,N_17711,N_17789);
or U18341 (N_18341,N_16851,N_16294);
or U18342 (N_18342,N_17149,N_16566);
or U18343 (N_18343,N_17397,N_16283);
nand U18344 (N_18344,N_16645,N_17107);
nor U18345 (N_18345,N_17695,N_17116);
or U18346 (N_18346,N_16147,N_17192);
nand U18347 (N_18347,N_17182,N_17706);
nor U18348 (N_18348,N_17008,N_17776);
nand U18349 (N_18349,N_17371,N_17566);
or U18350 (N_18350,N_17642,N_16362);
or U18351 (N_18351,N_16909,N_17066);
and U18352 (N_18352,N_17409,N_17275);
and U18353 (N_18353,N_17783,N_16667);
xnor U18354 (N_18354,N_16441,N_17764);
or U18355 (N_18355,N_17307,N_16858);
nand U18356 (N_18356,N_17897,N_16416);
or U18357 (N_18357,N_16394,N_17878);
nand U18358 (N_18358,N_16801,N_16296);
xnor U18359 (N_18359,N_16026,N_16304);
and U18360 (N_18360,N_17961,N_16460);
and U18361 (N_18361,N_16916,N_17864);
nand U18362 (N_18362,N_16359,N_17734);
or U18363 (N_18363,N_17241,N_17742);
or U18364 (N_18364,N_16689,N_16584);
xnor U18365 (N_18365,N_17604,N_17612);
nand U18366 (N_18366,N_16714,N_17554);
nor U18367 (N_18367,N_16464,N_16901);
or U18368 (N_18368,N_16047,N_17408);
or U18369 (N_18369,N_17511,N_17161);
nand U18370 (N_18370,N_17539,N_16068);
xnor U18371 (N_18371,N_17656,N_17029);
nand U18372 (N_18372,N_16560,N_17121);
xnor U18373 (N_18373,N_16282,N_17309);
nand U18374 (N_18374,N_17881,N_16273);
nor U18375 (N_18375,N_16339,N_17933);
nand U18376 (N_18376,N_16788,N_16199);
nand U18377 (N_18377,N_16512,N_16571);
and U18378 (N_18378,N_16564,N_16873);
or U18379 (N_18379,N_16422,N_17057);
nor U18380 (N_18380,N_16736,N_17098);
nand U18381 (N_18381,N_17385,N_17936);
nand U18382 (N_18382,N_17212,N_17287);
nand U18383 (N_18383,N_17587,N_17884);
nand U18384 (N_18384,N_16698,N_16053);
nor U18385 (N_18385,N_17335,N_16863);
and U18386 (N_18386,N_16918,N_16841);
nand U18387 (N_18387,N_16704,N_17037);
and U18388 (N_18388,N_16335,N_17775);
nand U18389 (N_18389,N_17755,N_17156);
and U18390 (N_18390,N_16948,N_17630);
xor U18391 (N_18391,N_17095,N_16652);
nand U18392 (N_18392,N_17575,N_17839);
nand U18393 (N_18393,N_17297,N_16085);
nor U18394 (N_18394,N_17985,N_16384);
and U18395 (N_18395,N_17703,N_17334);
or U18396 (N_18396,N_17025,N_17087);
and U18397 (N_18397,N_16035,N_17857);
and U18398 (N_18398,N_16447,N_17361);
and U18399 (N_18399,N_16220,N_17646);
and U18400 (N_18400,N_17626,N_17476);
nand U18401 (N_18401,N_16494,N_16044);
nor U18402 (N_18402,N_17555,N_17942);
or U18403 (N_18403,N_16562,N_16907);
or U18404 (N_18404,N_16129,N_16542);
or U18405 (N_18405,N_16099,N_17142);
nor U18406 (N_18406,N_17989,N_16893);
xnor U18407 (N_18407,N_17653,N_16329);
and U18408 (N_18408,N_17558,N_17749);
nand U18409 (N_18409,N_17747,N_17292);
nor U18410 (N_18410,N_16439,N_16453);
and U18411 (N_18411,N_16472,N_17128);
nand U18412 (N_18412,N_17915,N_16917);
or U18413 (N_18413,N_16091,N_17548);
xnor U18414 (N_18414,N_16691,N_17150);
and U18415 (N_18415,N_16984,N_17234);
nor U18416 (N_18416,N_16476,N_17298);
and U18417 (N_18417,N_17790,N_16401);
or U18418 (N_18418,N_16514,N_17751);
nor U18419 (N_18419,N_17898,N_17748);
nand U18420 (N_18420,N_16092,N_16588);
nor U18421 (N_18421,N_16520,N_16748);
xor U18422 (N_18422,N_17475,N_17428);
or U18423 (N_18423,N_17996,N_17853);
nor U18424 (N_18424,N_16859,N_16223);
nand U18425 (N_18425,N_16031,N_17627);
or U18426 (N_18426,N_17549,N_17901);
and U18427 (N_18427,N_17448,N_16780);
nand U18428 (N_18428,N_16781,N_17055);
and U18429 (N_18429,N_16497,N_17652);
xor U18430 (N_18430,N_17407,N_17369);
or U18431 (N_18431,N_16515,N_16504);
nor U18432 (N_18432,N_17237,N_16600);
nor U18433 (N_18433,N_17821,N_17453);
or U18434 (N_18434,N_17804,N_16852);
and U18435 (N_18435,N_17208,N_16318);
and U18436 (N_18436,N_17320,N_16703);
xor U18437 (N_18437,N_16017,N_17984);
or U18438 (N_18438,N_17079,N_16450);
and U18439 (N_18439,N_16254,N_17682);
or U18440 (N_18440,N_17602,N_17266);
or U18441 (N_18441,N_16545,N_16938);
xor U18442 (N_18442,N_16849,N_16687);
nor U18443 (N_18443,N_17590,N_17593);
and U18444 (N_18444,N_16774,N_17392);
xor U18445 (N_18445,N_16657,N_17222);
or U18446 (N_18446,N_17707,N_16189);
or U18447 (N_18447,N_17609,N_16042);
or U18448 (N_18448,N_16665,N_17530);
or U18449 (N_18449,N_17722,N_17701);
nor U18450 (N_18450,N_17051,N_16468);
and U18451 (N_18451,N_17086,N_17865);
xnor U18452 (N_18452,N_16435,N_17306);
nand U18453 (N_18453,N_17186,N_16205);
nor U18454 (N_18454,N_17913,N_16763);
xor U18455 (N_18455,N_17456,N_17450);
and U18456 (N_18456,N_17971,N_16979);
nand U18457 (N_18457,N_16550,N_16113);
nand U18458 (N_18458,N_16941,N_16706);
and U18459 (N_18459,N_17979,N_17621);
or U18460 (N_18460,N_16761,N_17127);
or U18461 (N_18461,N_16173,N_17184);
or U18462 (N_18462,N_16835,N_17379);
or U18463 (N_18463,N_17075,N_16997);
nand U18464 (N_18464,N_17577,N_16933);
or U18465 (N_18465,N_17469,N_17477);
and U18466 (N_18466,N_16102,N_17291);
nor U18467 (N_18467,N_16908,N_16116);
nand U18468 (N_18468,N_17517,N_17927);
and U18469 (N_18469,N_16570,N_17724);
and U18470 (N_18470,N_17890,N_17305);
nand U18471 (N_18471,N_16481,N_16048);
nor U18472 (N_18472,N_16976,N_17263);
and U18473 (N_18473,N_17922,N_17595);
nor U18474 (N_18474,N_17403,N_16338);
xnor U18475 (N_18475,N_16141,N_17389);
nor U18476 (N_18476,N_16368,N_17084);
and U18477 (N_18477,N_17739,N_16292);
nor U18478 (N_18478,N_17411,N_16879);
or U18479 (N_18479,N_16253,N_17781);
nand U18480 (N_18480,N_17412,N_16380);
nand U18481 (N_18481,N_16955,N_16717);
nand U18482 (N_18482,N_16983,N_17757);
xnor U18483 (N_18483,N_17917,N_17016);
nor U18484 (N_18484,N_17312,N_16912);
or U18485 (N_18485,N_17606,N_16265);
and U18486 (N_18486,N_17754,N_16083);
and U18487 (N_18487,N_17229,N_16074);
nand U18488 (N_18488,N_17048,N_16109);
nand U18489 (N_18489,N_16342,N_17140);
or U18490 (N_18490,N_17045,N_16834);
nand U18491 (N_18491,N_16187,N_17231);
nand U18492 (N_18492,N_17693,N_17446);
or U18493 (N_18493,N_17185,N_17768);
or U18494 (N_18494,N_17382,N_16119);
nand U18495 (N_18495,N_17825,N_17867);
and U18496 (N_18496,N_17248,N_17851);
nand U18497 (N_18497,N_17647,N_17608);
or U18498 (N_18498,N_17512,N_17676);
and U18499 (N_18499,N_16298,N_17728);
nand U18500 (N_18500,N_17155,N_16194);
and U18501 (N_18501,N_16230,N_17607);
or U18502 (N_18502,N_16872,N_16345);
nor U18503 (N_18503,N_17035,N_16776);
or U18504 (N_18504,N_17146,N_17963);
nor U18505 (N_18505,N_17895,N_17424);
nand U18506 (N_18506,N_16534,N_16952);
xor U18507 (N_18507,N_16707,N_17002);
nand U18508 (N_18508,N_17282,N_17858);
and U18509 (N_18509,N_16743,N_16768);
nor U18510 (N_18510,N_16790,N_16039);
nor U18511 (N_18511,N_17938,N_16583);
nor U18512 (N_18512,N_17924,N_16943);
nor U18513 (N_18513,N_17015,N_17521);
or U18514 (N_18514,N_16818,N_17018);
and U18515 (N_18515,N_16149,N_17740);
and U18516 (N_18516,N_16739,N_17294);
and U18517 (N_18517,N_16090,N_16823);
and U18518 (N_18518,N_17562,N_16530);
and U18519 (N_18519,N_17440,N_16100);
nor U18520 (N_18520,N_16103,N_17960);
and U18521 (N_18521,N_17097,N_17735);
or U18522 (N_18522,N_16982,N_16819);
and U18523 (N_18523,N_16628,N_16548);
nand U18524 (N_18524,N_16720,N_17007);
xor U18525 (N_18525,N_17068,N_16716);
or U18526 (N_18526,N_17508,N_17073);
or U18527 (N_18527,N_17199,N_16531);
xnor U18528 (N_18528,N_16032,N_17264);
or U18529 (N_18529,N_16500,N_16222);
and U18530 (N_18530,N_17540,N_17815);
or U18531 (N_18531,N_17168,N_16180);
nor U18532 (N_18532,N_16631,N_17281);
and U18533 (N_18533,N_17223,N_17402);
or U18534 (N_18534,N_17611,N_16897);
and U18535 (N_18535,N_16812,N_16256);
or U18536 (N_18536,N_17547,N_16961);
or U18537 (N_18537,N_16393,N_17822);
nand U18538 (N_18538,N_17823,N_16346);
xnor U18539 (N_18539,N_16247,N_17487);
and U18540 (N_18540,N_17302,N_17982);
nor U18541 (N_18541,N_16904,N_16148);
nor U18542 (N_18542,N_17896,N_16364);
and U18543 (N_18543,N_16846,N_16373);
and U18544 (N_18544,N_16245,N_17242);
and U18545 (N_18545,N_16742,N_17372);
and U18546 (N_18546,N_17967,N_16753);
nor U18547 (N_18547,N_16276,N_17499);
or U18548 (N_18548,N_16041,N_17145);
nand U18549 (N_18549,N_17284,N_17721);
xor U18550 (N_18550,N_16635,N_16320);
xor U18551 (N_18551,N_17619,N_17460);
xor U18552 (N_18552,N_17099,N_16931);
or U18553 (N_18553,N_17419,N_16025);
or U18554 (N_18554,N_16198,N_16615);
or U18555 (N_18555,N_17955,N_16438);
nor U18556 (N_18556,N_16388,N_16168);
nand U18557 (N_18557,N_17367,N_16135);
or U18558 (N_18558,N_17660,N_17666);
nor U18559 (N_18559,N_17216,N_17105);
or U18560 (N_18560,N_16671,N_16284);
nand U18561 (N_18561,N_17052,N_17447);
xor U18562 (N_18562,N_16319,N_16699);
nand U18563 (N_18563,N_17944,N_17488);
nand U18564 (N_18564,N_16783,N_16885);
nand U18565 (N_18565,N_16544,N_17280);
nor U18566 (N_18566,N_16953,N_16349);
nor U18567 (N_18567,N_17224,N_17452);
nand U18568 (N_18568,N_16794,N_17245);
nand U18569 (N_18569,N_16540,N_17589);
or U18570 (N_18570,N_16747,N_16898);
nand U18571 (N_18571,N_16334,N_16656);
or U18572 (N_18572,N_16210,N_16649);
nand U18573 (N_18573,N_17170,N_17497);
nor U18574 (N_18574,N_16490,N_16519);
nor U18575 (N_18575,N_16991,N_16066);
nor U18576 (N_18576,N_17718,N_17353);
nand U18577 (N_18577,N_17571,N_17376);
or U18578 (N_18578,N_16376,N_16552);
nor U18579 (N_18579,N_16073,N_16557);
or U18580 (N_18580,N_17840,N_16442);
xnor U18581 (N_18581,N_17994,N_17520);
xor U18582 (N_18582,N_16837,N_17434);
nand U18583 (N_18583,N_16987,N_16646);
or U18584 (N_18584,N_16574,N_17246);
nor U18585 (N_18585,N_17115,N_16789);
and U18586 (N_18586,N_16547,N_17180);
nor U18587 (N_18587,N_16417,N_17926);
nand U18588 (N_18588,N_16322,N_17580);
and U18589 (N_18589,N_16618,N_17561);
xnor U18590 (N_18590,N_17472,N_16372);
or U18591 (N_18591,N_16317,N_17514);
or U18592 (N_18592,N_16403,N_17330);
nand U18593 (N_18593,N_16461,N_16306);
and U18594 (N_18594,N_16466,N_17655);
nor U18595 (N_18595,N_17337,N_16855);
nor U18596 (N_18596,N_16700,N_17597);
nor U18597 (N_18597,N_16021,N_17874);
or U18598 (N_18598,N_16034,N_17689);
xor U18599 (N_18599,N_16940,N_17843);
nand U18600 (N_18600,N_16040,N_17969);
or U18601 (N_18601,N_17842,N_16363);
nand U18602 (N_18602,N_16398,N_16431);
or U18603 (N_18603,N_16881,N_17277);
xnor U18604 (N_18604,N_16045,N_16692);
and U18605 (N_18605,N_17089,N_16308);
and U18606 (N_18606,N_16064,N_17909);
nor U18607 (N_18607,N_17782,N_16488);
nand U18608 (N_18608,N_17293,N_16158);
or U18609 (N_18609,N_17047,N_17719);
or U18610 (N_18610,N_16251,N_17139);
and U18611 (N_18611,N_16078,N_16390);
nor U18612 (N_18612,N_17226,N_17258);
nor U18613 (N_18613,N_16479,N_16300);
or U18614 (N_18614,N_16449,N_17870);
nor U18615 (N_18615,N_16980,N_16586);
or U18616 (N_18616,N_16507,N_17773);
xnor U18617 (N_18617,N_17126,N_16833);
and U18618 (N_18618,N_17195,N_16186);
or U18619 (N_18619,N_17421,N_17911);
nor U18620 (N_18620,N_17640,N_17253);
nor U18621 (N_18621,N_17202,N_16213);
and U18622 (N_18622,N_17657,N_16596);
and U18623 (N_18623,N_16307,N_16311);
or U18624 (N_18624,N_16331,N_17350);
or U18625 (N_18625,N_16902,N_17664);
and U18626 (N_18626,N_16883,N_17948);
nor U18627 (N_18627,N_17573,N_16915);
or U18628 (N_18628,N_17675,N_17272);
xor U18629 (N_18629,N_16316,N_17981);
nor U18630 (N_18630,N_17993,N_16352);
nor U18631 (N_18631,N_17920,N_16261);
and U18632 (N_18632,N_16037,N_17868);
nand U18633 (N_18633,N_17053,N_17532);
nor U18634 (N_18634,N_16347,N_16138);
nand U18635 (N_18635,N_17574,N_16832);
nor U18636 (N_18636,N_17232,N_17705);
or U18637 (N_18637,N_17551,N_16458);
or U18638 (N_18638,N_16387,N_16679);
and U18639 (N_18639,N_17152,N_17648);
and U18640 (N_18640,N_16086,N_16258);
nor U18641 (N_18641,N_17233,N_17473);
nand U18642 (N_18642,N_17352,N_17014);
or U18643 (N_18643,N_16289,N_17542);
and U18644 (N_18644,N_16378,N_16420);
nor U18645 (N_18645,N_16302,N_16208);
and U18646 (N_18646,N_17310,N_16012);
xnor U18647 (N_18647,N_17213,N_17904);
or U18648 (N_18648,N_17683,N_17537);
and U18649 (N_18649,N_17743,N_16923);
xor U18650 (N_18650,N_16020,N_17221);
and U18651 (N_18651,N_16108,N_17043);
or U18652 (N_18652,N_17296,N_17159);
xor U18653 (N_18653,N_16327,N_16556);
or U18654 (N_18654,N_17344,N_16890);
or U18655 (N_18655,N_16427,N_17316);
or U18656 (N_18656,N_16553,N_17244);
nand U18657 (N_18657,N_16142,N_17160);
and U18658 (N_18658,N_17636,N_16517);
nand U18659 (N_18659,N_16697,N_17855);
and U18660 (N_18660,N_16595,N_16844);
xor U18661 (N_18661,N_16778,N_16215);
nor U18662 (N_18662,N_17157,N_17987);
nor U18663 (N_18663,N_17691,N_17792);
or U18664 (N_18664,N_17163,N_16122);
nor U18665 (N_18665,N_16960,N_17937);
nand U18666 (N_18666,N_17308,N_16662);
nand U18667 (N_18667,N_17467,N_16648);
or U18668 (N_18668,N_16056,N_17026);
or U18669 (N_18669,N_16429,N_16321);
xnor U18670 (N_18670,N_17480,N_17524);
nand U18671 (N_18671,N_16787,N_17355);
nand U18672 (N_18672,N_16350,N_17462);
and U18673 (N_18673,N_16501,N_16144);
xor U18674 (N_18674,N_16797,N_16096);
nand U18675 (N_18675,N_17483,N_17129);
nand U18676 (N_18676,N_17074,N_16813);
nor U18677 (N_18677,N_16095,N_17727);
xnor U18678 (N_18678,N_16684,N_16930);
nand U18679 (N_18679,N_16573,N_17714);
nand U18680 (N_18680,N_16470,N_16004);
and U18681 (N_18681,N_16075,N_16028);
or U18682 (N_18682,N_16492,N_17300);
and U18683 (N_18683,N_16681,N_17797);
nor U18684 (N_18684,N_16009,N_17820);
xnor U18685 (N_18685,N_17124,N_17413);
nand U18686 (N_18686,N_17028,N_16192);
nor U18687 (N_18687,N_17717,N_17586);
nor U18688 (N_18688,N_17578,N_17774);
or U18689 (N_18689,N_17290,N_16593);
nand U18690 (N_18690,N_16624,N_16062);
nor U18691 (N_18691,N_16143,N_17973);
or U18692 (N_18692,N_17560,N_16626);
nand U18693 (N_18693,N_16101,N_17614);
nand U18694 (N_18694,N_16724,N_17414);
or U18695 (N_18695,N_17019,N_17017);
xnor U18696 (N_18696,N_16894,N_16061);
nand U18697 (N_18697,N_16171,N_16206);
nand U18698 (N_18698,N_16549,N_16575);
and U18699 (N_18699,N_17276,N_16604);
nor U18700 (N_18700,N_17082,N_16710);
xor U18701 (N_18701,N_16708,N_17600);
xor U18702 (N_18702,N_16008,N_17398);
nor U18703 (N_18703,N_16330,N_17930);
nor U18704 (N_18704,N_17137,N_16400);
nand U18705 (N_18705,N_17349,N_17228);
or U18706 (N_18706,N_16315,N_16944);
nand U18707 (N_18707,N_17406,N_16259);
nor U18708 (N_18708,N_17680,N_16324);
and U18709 (N_18709,N_16182,N_17416);
nor U18710 (N_18710,N_16585,N_17886);
or U18711 (N_18711,N_16369,N_17463);
nand U18712 (N_18712,N_16231,N_17324);
xnor U18713 (N_18713,N_17616,N_16454);
and U18714 (N_18714,N_17765,N_17594);
and U18715 (N_18715,N_16436,N_16958);
and U18716 (N_18716,N_16525,N_17885);
nor U18717 (N_18717,N_16425,N_17001);
or U18718 (N_18718,N_17113,N_17553);
and U18719 (N_18719,N_17021,N_17181);
nand U18720 (N_18720,N_17778,N_16592);
nand U18721 (N_18721,N_17239,N_17191);
nor U18722 (N_18722,N_16870,N_16155);
xor U18723 (N_18723,N_16050,N_16935);
nor U18724 (N_18724,N_16036,N_17125);
nand U18725 (N_18725,N_17956,N_16079);
and U18726 (N_18726,N_17908,N_16800);
or U18727 (N_18727,N_17445,N_17800);
xor U18728 (N_18728,N_16139,N_17203);
or U18729 (N_18729,N_16218,N_16328);
nand U18730 (N_18730,N_17688,N_17069);
xor U18731 (N_18731,N_17645,N_16232);
nand U18732 (N_18732,N_16089,N_16910);
nand U18733 (N_18733,N_17366,N_16172);
or U18734 (N_18734,N_17102,N_17531);
or U18735 (N_18735,N_16862,N_16027);
nor U18736 (N_18736,N_17474,N_16386);
and U18737 (N_18737,N_17083,N_16415);
nand U18738 (N_18738,N_17426,N_17958);
and U18739 (N_18739,N_17677,N_17417);
nand U18740 (N_18740,N_16601,N_17582);
and U18741 (N_18741,N_16303,N_16446);
nor U18742 (N_18742,N_16246,N_17268);
nor U18743 (N_18743,N_17422,N_16880);
nor U18744 (N_18744,N_17238,N_17769);
or U18745 (N_18745,N_16137,N_17092);
nand U18746 (N_18746,N_17639,N_16994);
nor U18747 (N_18747,N_17172,N_16193);
nor U18748 (N_18748,N_17436,N_16117);
nand U18749 (N_18749,N_16059,N_17420);
nand U18750 (N_18750,N_16252,N_16385);
nor U18751 (N_18751,N_16176,N_17527);
nand U18752 (N_18752,N_17812,N_17641);
nor U18753 (N_18753,N_16203,N_16082);
and U18754 (N_18754,N_17861,N_16568);
nor U18755 (N_18755,N_16145,N_16641);
nand U18756 (N_18756,N_17533,N_16937);
or U18757 (N_18757,N_17733,N_16764);
and U18758 (N_18758,N_17158,N_17699);
nand U18759 (N_18759,N_16326,N_17891);
nor U18760 (N_18760,N_17030,N_17265);
or U18761 (N_18761,N_17484,N_17669);
or U18762 (N_18762,N_16627,N_17925);
or U18763 (N_18763,N_16404,N_16030);
nand U18764 (N_18764,N_17651,N_17844);
or U18765 (N_18765,N_16651,N_17201);
or U18766 (N_18766,N_16664,N_17151);
nor U18767 (N_18767,N_17027,N_16805);
xnor U18768 (N_18768,N_16811,N_16723);
nand U18769 (N_18769,N_16433,N_17377);
nor U18770 (N_18770,N_17279,N_17090);
or U18771 (N_18771,N_16650,N_16990);
nor U18772 (N_18772,N_17039,N_16272);
nand U18773 (N_18773,N_16278,N_17067);
nand U18774 (N_18774,N_16291,N_17638);
nand U18775 (N_18775,N_17945,N_16255);
and U18776 (N_18776,N_17011,N_16107);
nor U18777 (N_18777,N_17171,N_16134);
or U18778 (N_18778,N_17988,N_17905);
or U18779 (N_18779,N_16010,N_16539);
and U18780 (N_18780,N_17136,N_17723);
and U18781 (N_18781,N_16785,N_17315);
or U18782 (N_18782,N_16184,N_16456);
nor U18783 (N_18783,N_17004,N_16653);
or U18784 (N_18784,N_16200,N_16674);
nor U18785 (N_18785,N_17799,N_16204);
nor U18786 (N_18786,N_16521,N_17716);
nand U18787 (N_18787,N_16632,N_16554);
nor U18788 (N_18788,N_16518,N_17962);
or U18789 (N_18789,N_17495,N_17056);
and U18790 (N_18790,N_17674,N_16896);
nor U18791 (N_18791,N_17299,N_17059);
nand U18792 (N_18792,N_17523,N_16006);
or U18793 (N_18793,N_17557,N_17333);
nand U18794 (N_18794,N_16195,N_16925);
or U18795 (N_18795,N_16290,N_16620);
and U18796 (N_18796,N_17271,N_17694);
nor U18797 (N_18797,N_16755,N_17346);
xor U18798 (N_18798,N_16999,N_17288);
nand U18799 (N_18799,N_16188,N_17583);
nand U18800 (N_18800,N_17543,N_16166);
nor U18801 (N_18801,N_17835,N_16310);
or U18802 (N_18802,N_17863,N_17545);
nor U18803 (N_18803,N_17122,N_17819);
xnor U18804 (N_18804,N_17741,N_16493);
xnor U18805 (N_18805,N_17023,N_17622);
nand U18806 (N_18806,N_17931,N_17834);
nand U18807 (N_18807,N_17459,N_17892);
or U18808 (N_18808,N_17358,N_17565);
and U18809 (N_18809,N_16097,N_17378);
and U18810 (N_18810,N_17921,N_16877);
or U18811 (N_18811,N_16978,N_16694);
or U18812 (N_18812,N_17806,N_16947);
xnor U18813 (N_18813,N_16777,N_17598);
and U18814 (N_18814,N_16162,N_17169);
or U18815 (N_18815,N_16589,N_17162);
nand U18816 (N_18816,N_16625,N_17869);
nand U18817 (N_18817,N_16146,N_17667);
nand U18818 (N_18818,N_17076,N_16510);
nand U18819 (N_18819,N_16271,N_17363);
nor U18820 (N_18820,N_16474,N_17328);
nor U18821 (N_18821,N_17522,N_16229);
nand U18822 (N_18822,N_16104,N_16824);
and U18823 (N_18823,N_17827,N_17470);
or U18824 (N_18824,N_16131,N_16299);
nand U18825 (N_18825,N_16402,N_16190);
and U18826 (N_18826,N_16922,N_16569);
nor U18827 (N_18827,N_16532,N_16954);
nor U18828 (N_18828,N_16262,N_16274);
and U18829 (N_18829,N_17866,N_16336);
or U18830 (N_18830,N_16529,N_17348);
or U18831 (N_18831,N_17507,N_17910);
or U18832 (N_18832,N_17846,N_17110);
nand U18833 (N_18833,N_16825,N_17852);
and U18834 (N_18834,N_16719,N_16049);
and U18835 (N_18835,N_16029,N_16750);
nand U18836 (N_18836,N_16305,N_16234);
and U18837 (N_18837,N_16018,N_16766);
xnor U18838 (N_18838,N_17679,N_16749);
and U18839 (N_18839,N_16207,N_17193);
nand U18840 (N_18840,N_16640,N_17218);
nand U18841 (N_18841,N_16989,N_16567);
and U18842 (N_18842,N_16536,N_17364);
and U18843 (N_18843,N_17817,N_17983);
xor U18844 (N_18844,N_16967,N_17031);
or U18845 (N_18845,N_17465,N_17802);
nor U18846 (N_18846,N_17686,N_16582);
or U18847 (N_18847,N_17505,N_16690);
nand U18848 (N_18848,N_17455,N_17854);
or U18849 (N_18849,N_17050,N_17197);
and U18850 (N_18850,N_17164,N_16065);
and U18851 (N_18851,N_17167,N_17196);
nor U18852 (N_18852,N_16840,N_16052);
nand U18853 (N_18853,N_17715,N_16972);
and U18854 (N_18854,N_16250,N_17054);
nand U18855 (N_18855,N_17189,N_16775);
or U18856 (N_18856,N_17671,N_16423);
nand U18857 (N_18857,N_16054,N_17386);
or U18858 (N_18858,N_17143,N_16809);
nor U18859 (N_18859,N_17262,N_17801);
and U18860 (N_18860,N_16906,N_16156);
nand U18861 (N_18861,N_16411,N_17020);
nor U18862 (N_18862,N_17466,N_17939);
nand U18863 (N_18863,N_16077,N_17745);
nor U18864 (N_18864,N_16241,N_16629);
xnor U18865 (N_18865,N_17596,N_16957);
nor U18866 (N_18866,N_16154,N_16956);
nand U18867 (N_18867,N_17165,N_17725);
nand U18868 (N_18868,N_16945,N_17356);
nand U18869 (N_18869,N_17183,N_16414);
and U18870 (N_18870,N_17049,N_16110);
nand U18871 (N_18871,N_17658,N_16786);
nor U18872 (N_18872,N_17859,N_17952);
nand U18873 (N_18873,N_16228,N_16759);
nor U18874 (N_18874,N_17235,N_16815);
xnor U18875 (N_18875,N_16993,N_17760);
nand U18876 (N_18876,N_16358,N_16882);
nand U18877 (N_18877,N_16543,N_16680);
xor U18878 (N_18878,N_16889,N_16892);
nor U18879 (N_18879,N_17599,N_17190);
and U18880 (N_18880,N_17331,N_16128);
and U18881 (N_18881,N_16591,N_16666);
and U18882 (N_18882,N_17485,N_17131);
nand U18883 (N_18883,N_17650,N_17175);
nor U18884 (N_18884,N_17635,N_17269);
nand U18885 (N_18885,N_16127,N_16421);
nand U18886 (N_18886,N_17123,N_17538);
nor U18887 (N_18887,N_17519,N_16854);
and U18888 (N_18888,N_16344,N_17995);
and U18889 (N_18889,N_16792,N_16735);
nor U18890 (N_18890,N_17953,N_16795);
nand U18891 (N_18891,N_16974,N_17362);
nor U18892 (N_18892,N_17882,N_17200);
or U18893 (N_18893,N_16057,N_17730);
and U18894 (N_18894,N_16279,N_17251);
xnor U18895 (N_18895,N_16682,N_17826);
nand U18896 (N_18896,N_17439,N_17976);
and U18897 (N_18897,N_16598,N_17941);
and U18898 (N_18898,N_17482,N_16617);
nor U18899 (N_18899,N_17383,N_16535);
nor U18900 (N_18900,N_17876,N_17431);
nand U18901 (N_18901,N_16405,N_17975);
xor U18902 (N_18902,N_17425,N_16807);
or U18903 (N_18903,N_17809,N_17659);
or U18904 (N_18904,N_16370,N_16713);
nor U18905 (N_18905,N_17862,N_16654);
nor U18906 (N_18906,N_16281,N_16407);
and U18907 (N_18907,N_16802,N_17365);
or U18908 (N_18908,N_16115,N_17685);
and U18909 (N_18909,N_16900,N_17563);
xor U18910 (N_18910,N_17273,N_16397);
nand U18911 (N_18911,N_16130,N_17481);
or U18912 (N_18912,N_16677,N_17753);
nand U18913 (N_18913,N_16686,N_16668);
xnor U18914 (N_18914,N_17496,N_16822);
nand U18915 (N_18915,N_17750,N_17564);
or U18916 (N_18916,N_17329,N_17085);
and U18917 (N_18917,N_17556,N_16244);
nand U18918 (N_18918,N_17443,N_16174);
nand U18919 (N_18919,N_17154,N_16603);
or U18920 (N_18920,N_16365,N_16878);
xnor U18921 (N_18921,N_16924,N_17618);
or U18922 (N_18922,N_17702,N_17247);
nor U18923 (N_18923,N_17729,N_17317);
nor U18924 (N_18924,N_16950,N_17502);
nor U18925 (N_18925,N_16985,N_17643);
and U18926 (N_18926,N_17368,N_17807);
and U18927 (N_18927,N_16702,N_17631);
or U18928 (N_18928,N_17432,N_16314);
and U18929 (N_18929,N_16712,N_17516);
or U18930 (N_18930,N_17829,N_17111);
nor U18931 (N_18931,N_17303,N_17649);
or U18932 (N_18932,N_17847,N_16487);
xor U18933 (N_18933,N_17108,N_17824);
or U18934 (N_18934,N_17153,N_16669);
nand U18935 (N_18935,N_16217,N_16120);
and U18936 (N_18936,N_17270,N_17283);
or U18937 (N_18937,N_17423,N_16920);
nand U18938 (N_18938,N_16014,N_16647);
and U18939 (N_18939,N_16803,N_17628);
and U18940 (N_18940,N_17295,N_16572);
nor U18941 (N_18941,N_17603,N_16503);
nor U18942 (N_18942,N_16392,N_16779);
nor U18943 (N_18943,N_16757,N_17148);
nand U18944 (N_18944,N_16709,N_16280);
nand U18945 (N_18945,N_16741,N_17345);
or U18946 (N_18946,N_16333,N_17096);
nand U18947 (N_18947,N_16678,N_16565);
or U18948 (N_18948,N_16838,N_17828);
and U18949 (N_18949,N_17849,N_16051);
nand U18950 (N_18950,N_17883,N_16293);
nor U18951 (N_18951,N_17118,N_17914);
or U18952 (N_18952,N_16225,N_17252);
and U18953 (N_18953,N_16264,N_16391);
nor U18954 (N_18954,N_16602,N_16325);
nor U18955 (N_18955,N_16921,N_16929);
nor U18956 (N_18956,N_16875,N_17256);
nor U18957 (N_18957,N_16366,N_17415);
or U18958 (N_18958,N_17692,N_16399);
nand U18959 (N_18959,N_16471,N_17954);
and U18960 (N_18960,N_17509,N_17568);
and U18961 (N_18961,N_17697,N_16354);
or U18962 (N_18962,N_16297,N_17831);
or U18963 (N_18963,N_17620,N_17219);
and U18964 (N_18964,N_17710,N_17394);
nor U18965 (N_18965,N_17388,N_17894);
or U18966 (N_18966,N_17071,N_16670);
nand U18967 (N_18967,N_17559,N_16383);
or U18968 (N_18968,N_16643,N_17318);
nand U18969 (N_18969,N_16721,N_16919);
or U18970 (N_18970,N_17094,N_16696);
or U18971 (N_18971,N_17236,N_16533);
and U18972 (N_18972,N_16098,N_17759);
nand U18973 (N_18973,N_17274,N_16946);
and U18974 (N_18974,N_17177,N_17992);
nand U18975 (N_18975,N_17359,N_17230);
or U18976 (N_18976,N_17761,N_16202);
or U18977 (N_18977,N_16377,N_17339);
and U18978 (N_18978,N_17513,N_16523);
or U18979 (N_18979,N_16212,N_17390);
and U18980 (N_18980,N_16167,N_17906);
or U18981 (N_18981,N_17966,N_16868);
xor U18982 (N_18982,N_17661,N_16038);
and U18983 (N_18983,N_16063,N_17613);
nand U18984 (N_18984,N_16939,N_17856);
nand U18985 (N_18985,N_17101,N_17176);
nor U18986 (N_18986,N_16486,N_16239);
xor U18987 (N_18987,N_17227,N_16658);
or U18988 (N_18988,N_17384,N_17687);
nor U18989 (N_18989,N_16216,N_16913);
or U18990 (N_18990,N_17793,N_17615);
nand U18991 (N_18991,N_16480,N_16613);
or U18992 (N_18992,N_17211,N_16375);
nand U18993 (N_18993,N_16266,N_16046);
nor U18994 (N_18994,N_16181,N_17579);
xnor U18995 (N_18995,N_16577,N_17444);
nand U18996 (N_18996,N_16161,N_17207);
nand U18997 (N_18997,N_16268,N_17451);
nand U18998 (N_18998,N_17464,N_17471);
xor U18999 (N_18999,N_16606,N_16842);
or U19000 (N_19000,N_17064,N_16453);
nor U19001 (N_19001,N_16560,N_16290);
nand U19002 (N_19002,N_17619,N_17528);
and U19003 (N_19003,N_16956,N_16011);
or U19004 (N_19004,N_16062,N_16818);
nor U19005 (N_19005,N_16117,N_16852);
nor U19006 (N_19006,N_17226,N_16358);
nor U19007 (N_19007,N_16030,N_17041);
nand U19008 (N_19008,N_17337,N_16445);
and U19009 (N_19009,N_17772,N_16572);
nand U19010 (N_19010,N_16833,N_16900);
and U19011 (N_19011,N_17350,N_17784);
or U19012 (N_19012,N_16973,N_17556);
or U19013 (N_19013,N_16142,N_17017);
nand U19014 (N_19014,N_17871,N_16692);
nand U19015 (N_19015,N_17117,N_17266);
and U19016 (N_19016,N_17905,N_16758);
and U19017 (N_19017,N_16268,N_16406);
nor U19018 (N_19018,N_17779,N_17445);
nand U19019 (N_19019,N_17080,N_17156);
or U19020 (N_19020,N_16271,N_17522);
nor U19021 (N_19021,N_17205,N_16000);
and U19022 (N_19022,N_17329,N_17641);
nand U19023 (N_19023,N_16842,N_17366);
xor U19024 (N_19024,N_16519,N_16298);
and U19025 (N_19025,N_16901,N_17611);
nor U19026 (N_19026,N_17340,N_16319);
or U19027 (N_19027,N_16523,N_16776);
nor U19028 (N_19028,N_16609,N_17947);
xor U19029 (N_19029,N_17814,N_16035);
nor U19030 (N_19030,N_16484,N_16861);
nand U19031 (N_19031,N_17760,N_16322);
nand U19032 (N_19032,N_16072,N_16346);
or U19033 (N_19033,N_17172,N_16050);
nand U19034 (N_19034,N_16316,N_17022);
nand U19035 (N_19035,N_17668,N_16377);
or U19036 (N_19036,N_16904,N_17491);
xnor U19037 (N_19037,N_16279,N_16268);
nand U19038 (N_19038,N_17790,N_17745);
nor U19039 (N_19039,N_16999,N_16436);
or U19040 (N_19040,N_16826,N_16896);
nand U19041 (N_19041,N_17661,N_16471);
xor U19042 (N_19042,N_16386,N_16807);
nand U19043 (N_19043,N_17460,N_17695);
nor U19044 (N_19044,N_16357,N_17125);
and U19045 (N_19045,N_17859,N_17862);
nand U19046 (N_19046,N_17640,N_16868);
nor U19047 (N_19047,N_17442,N_17580);
xor U19048 (N_19048,N_17764,N_16243);
or U19049 (N_19049,N_17940,N_17973);
nand U19050 (N_19050,N_17048,N_17154);
and U19051 (N_19051,N_17664,N_17928);
nand U19052 (N_19052,N_17256,N_17547);
or U19053 (N_19053,N_16114,N_16176);
nand U19054 (N_19054,N_16727,N_16323);
or U19055 (N_19055,N_16622,N_16437);
nor U19056 (N_19056,N_16484,N_16665);
xnor U19057 (N_19057,N_16908,N_16258);
nor U19058 (N_19058,N_16499,N_16514);
nand U19059 (N_19059,N_17362,N_16993);
and U19060 (N_19060,N_16665,N_16351);
nor U19061 (N_19061,N_17047,N_16962);
or U19062 (N_19062,N_16909,N_16304);
or U19063 (N_19063,N_17177,N_16279);
or U19064 (N_19064,N_17266,N_16892);
xnor U19065 (N_19065,N_17300,N_17926);
nand U19066 (N_19066,N_17828,N_17144);
nand U19067 (N_19067,N_17926,N_17427);
and U19068 (N_19068,N_16329,N_16571);
nor U19069 (N_19069,N_16402,N_16035);
or U19070 (N_19070,N_17624,N_17765);
or U19071 (N_19071,N_17161,N_17041);
or U19072 (N_19072,N_16333,N_17053);
or U19073 (N_19073,N_16747,N_17182);
and U19074 (N_19074,N_17912,N_16960);
nor U19075 (N_19075,N_16633,N_16847);
and U19076 (N_19076,N_17039,N_16641);
and U19077 (N_19077,N_17403,N_17543);
nor U19078 (N_19078,N_17386,N_16468);
or U19079 (N_19079,N_16534,N_17553);
or U19080 (N_19080,N_16560,N_17750);
or U19081 (N_19081,N_17576,N_17683);
nor U19082 (N_19082,N_16940,N_16983);
and U19083 (N_19083,N_16127,N_16360);
nand U19084 (N_19084,N_16876,N_17099);
nor U19085 (N_19085,N_17461,N_16154);
or U19086 (N_19086,N_17010,N_17922);
or U19087 (N_19087,N_17442,N_16972);
and U19088 (N_19088,N_17043,N_17664);
or U19089 (N_19089,N_16083,N_17122);
or U19090 (N_19090,N_17952,N_16423);
or U19091 (N_19091,N_16974,N_17674);
and U19092 (N_19092,N_16661,N_17433);
or U19093 (N_19093,N_16503,N_17625);
and U19094 (N_19094,N_17747,N_17960);
nand U19095 (N_19095,N_17567,N_16484);
and U19096 (N_19096,N_16658,N_17114);
xnor U19097 (N_19097,N_17937,N_17918);
and U19098 (N_19098,N_16065,N_17753);
and U19099 (N_19099,N_17958,N_17416);
nand U19100 (N_19100,N_16668,N_17109);
and U19101 (N_19101,N_17409,N_16755);
nand U19102 (N_19102,N_16621,N_16832);
and U19103 (N_19103,N_16877,N_17681);
and U19104 (N_19104,N_17473,N_16844);
nand U19105 (N_19105,N_17621,N_17975);
nor U19106 (N_19106,N_17407,N_16583);
nand U19107 (N_19107,N_16150,N_17669);
and U19108 (N_19108,N_17348,N_17809);
nor U19109 (N_19109,N_17274,N_16568);
or U19110 (N_19110,N_17833,N_17162);
nand U19111 (N_19111,N_16812,N_17372);
nor U19112 (N_19112,N_16202,N_16742);
nor U19113 (N_19113,N_17299,N_16995);
or U19114 (N_19114,N_16913,N_16835);
and U19115 (N_19115,N_17742,N_17553);
xnor U19116 (N_19116,N_17430,N_16168);
nand U19117 (N_19117,N_17056,N_16303);
and U19118 (N_19118,N_17253,N_17841);
nor U19119 (N_19119,N_16947,N_17189);
xnor U19120 (N_19120,N_17049,N_16227);
or U19121 (N_19121,N_17574,N_17434);
nand U19122 (N_19122,N_16443,N_16491);
and U19123 (N_19123,N_16056,N_17863);
nor U19124 (N_19124,N_16978,N_16840);
xor U19125 (N_19125,N_16148,N_16607);
or U19126 (N_19126,N_17992,N_16956);
nor U19127 (N_19127,N_17737,N_16092);
or U19128 (N_19128,N_17016,N_17714);
xnor U19129 (N_19129,N_16975,N_17213);
nand U19130 (N_19130,N_17416,N_17438);
nor U19131 (N_19131,N_17483,N_16080);
nand U19132 (N_19132,N_16873,N_16344);
and U19133 (N_19133,N_17974,N_16277);
and U19134 (N_19134,N_16358,N_16308);
and U19135 (N_19135,N_16671,N_16254);
and U19136 (N_19136,N_17033,N_16172);
nand U19137 (N_19137,N_16190,N_16451);
nand U19138 (N_19138,N_16026,N_17775);
xnor U19139 (N_19139,N_16395,N_17771);
or U19140 (N_19140,N_17168,N_16025);
nor U19141 (N_19141,N_17268,N_16170);
xnor U19142 (N_19142,N_16663,N_16889);
or U19143 (N_19143,N_17459,N_16609);
or U19144 (N_19144,N_17913,N_17214);
or U19145 (N_19145,N_17737,N_17590);
nor U19146 (N_19146,N_17019,N_17263);
xor U19147 (N_19147,N_16341,N_17406);
nand U19148 (N_19148,N_17609,N_16763);
or U19149 (N_19149,N_17691,N_17828);
or U19150 (N_19150,N_17823,N_16522);
nor U19151 (N_19151,N_16926,N_17777);
and U19152 (N_19152,N_17169,N_16535);
and U19153 (N_19153,N_16711,N_17796);
or U19154 (N_19154,N_17800,N_16103);
nor U19155 (N_19155,N_16564,N_16474);
nor U19156 (N_19156,N_16359,N_16366);
and U19157 (N_19157,N_17604,N_17310);
and U19158 (N_19158,N_16164,N_17579);
nor U19159 (N_19159,N_16841,N_17134);
or U19160 (N_19160,N_17545,N_17081);
and U19161 (N_19161,N_16528,N_16544);
or U19162 (N_19162,N_17098,N_16014);
nand U19163 (N_19163,N_16386,N_17105);
nor U19164 (N_19164,N_17476,N_16453);
and U19165 (N_19165,N_17681,N_17130);
and U19166 (N_19166,N_16665,N_17545);
nand U19167 (N_19167,N_17376,N_16466);
or U19168 (N_19168,N_16341,N_16442);
nor U19169 (N_19169,N_16640,N_16738);
xnor U19170 (N_19170,N_17183,N_17388);
nor U19171 (N_19171,N_16515,N_16096);
nor U19172 (N_19172,N_17209,N_16349);
nor U19173 (N_19173,N_17437,N_17458);
nor U19174 (N_19174,N_17716,N_16765);
and U19175 (N_19175,N_17262,N_16143);
or U19176 (N_19176,N_16732,N_16102);
nor U19177 (N_19177,N_17957,N_16471);
and U19178 (N_19178,N_17158,N_17176);
or U19179 (N_19179,N_16483,N_17394);
nor U19180 (N_19180,N_17298,N_17425);
nand U19181 (N_19181,N_16088,N_17657);
nand U19182 (N_19182,N_16589,N_16592);
nand U19183 (N_19183,N_17060,N_17744);
and U19184 (N_19184,N_17674,N_17538);
nand U19185 (N_19185,N_16680,N_16382);
or U19186 (N_19186,N_17209,N_17327);
xor U19187 (N_19187,N_16213,N_16179);
nand U19188 (N_19188,N_16726,N_16201);
xnor U19189 (N_19189,N_17636,N_17961);
xnor U19190 (N_19190,N_17574,N_16221);
nand U19191 (N_19191,N_16646,N_17310);
and U19192 (N_19192,N_17275,N_17402);
nor U19193 (N_19193,N_17707,N_16462);
nor U19194 (N_19194,N_16066,N_16788);
and U19195 (N_19195,N_16674,N_16592);
nor U19196 (N_19196,N_17291,N_16488);
or U19197 (N_19197,N_16813,N_17857);
or U19198 (N_19198,N_16679,N_17785);
or U19199 (N_19199,N_16074,N_17847);
nand U19200 (N_19200,N_17122,N_16042);
and U19201 (N_19201,N_17702,N_16271);
nand U19202 (N_19202,N_16251,N_16025);
or U19203 (N_19203,N_17778,N_17493);
nor U19204 (N_19204,N_17431,N_17631);
or U19205 (N_19205,N_17823,N_17818);
or U19206 (N_19206,N_16070,N_16627);
xor U19207 (N_19207,N_16963,N_17656);
nand U19208 (N_19208,N_17449,N_16985);
xnor U19209 (N_19209,N_17791,N_17985);
or U19210 (N_19210,N_17225,N_17814);
or U19211 (N_19211,N_17701,N_17793);
nand U19212 (N_19212,N_17432,N_17974);
nand U19213 (N_19213,N_16716,N_16292);
or U19214 (N_19214,N_17170,N_16092);
nor U19215 (N_19215,N_17015,N_16397);
or U19216 (N_19216,N_16309,N_16487);
and U19217 (N_19217,N_16351,N_17185);
or U19218 (N_19218,N_17316,N_17143);
or U19219 (N_19219,N_17226,N_16611);
xor U19220 (N_19220,N_16738,N_16055);
nand U19221 (N_19221,N_16559,N_17596);
nor U19222 (N_19222,N_17341,N_16528);
and U19223 (N_19223,N_17183,N_16176);
and U19224 (N_19224,N_16778,N_16473);
nand U19225 (N_19225,N_16268,N_16526);
or U19226 (N_19226,N_17481,N_17061);
nand U19227 (N_19227,N_17303,N_16829);
and U19228 (N_19228,N_16935,N_17899);
and U19229 (N_19229,N_16071,N_16575);
nor U19230 (N_19230,N_16431,N_16651);
nor U19231 (N_19231,N_16860,N_17363);
or U19232 (N_19232,N_17065,N_17264);
nor U19233 (N_19233,N_17965,N_17485);
and U19234 (N_19234,N_17410,N_16014);
or U19235 (N_19235,N_17438,N_16247);
and U19236 (N_19236,N_17855,N_16917);
xnor U19237 (N_19237,N_17579,N_16734);
and U19238 (N_19238,N_16796,N_17210);
nand U19239 (N_19239,N_16107,N_17776);
and U19240 (N_19240,N_17633,N_17259);
nor U19241 (N_19241,N_17173,N_17436);
xnor U19242 (N_19242,N_17962,N_17730);
and U19243 (N_19243,N_17228,N_17943);
or U19244 (N_19244,N_17603,N_17970);
or U19245 (N_19245,N_16633,N_17338);
and U19246 (N_19246,N_16628,N_17262);
xor U19247 (N_19247,N_17152,N_17748);
nand U19248 (N_19248,N_17988,N_16216);
nor U19249 (N_19249,N_16077,N_17650);
nand U19250 (N_19250,N_16012,N_16081);
nor U19251 (N_19251,N_16778,N_16198);
nand U19252 (N_19252,N_17597,N_16476);
nand U19253 (N_19253,N_16080,N_17715);
and U19254 (N_19254,N_17528,N_17784);
xor U19255 (N_19255,N_16215,N_16873);
or U19256 (N_19256,N_17060,N_16761);
or U19257 (N_19257,N_16800,N_17758);
and U19258 (N_19258,N_17851,N_17657);
nand U19259 (N_19259,N_16526,N_16857);
nand U19260 (N_19260,N_17262,N_17788);
or U19261 (N_19261,N_17378,N_17197);
nand U19262 (N_19262,N_16998,N_17477);
or U19263 (N_19263,N_16401,N_17762);
and U19264 (N_19264,N_16341,N_16045);
xor U19265 (N_19265,N_17963,N_17316);
or U19266 (N_19266,N_16344,N_17672);
and U19267 (N_19267,N_17042,N_17051);
nor U19268 (N_19268,N_17818,N_17295);
nand U19269 (N_19269,N_17056,N_16448);
or U19270 (N_19270,N_17598,N_17449);
nor U19271 (N_19271,N_17010,N_16541);
or U19272 (N_19272,N_17228,N_16443);
xnor U19273 (N_19273,N_16289,N_16400);
or U19274 (N_19274,N_16743,N_17251);
and U19275 (N_19275,N_17811,N_16729);
nor U19276 (N_19276,N_17432,N_16913);
nor U19277 (N_19277,N_17120,N_16880);
nor U19278 (N_19278,N_17477,N_17894);
xor U19279 (N_19279,N_17432,N_16984);
or U19280 (N_19280,N_17838,N_16496);
or U19281 (N_19281,N_17492,N_17256);
xor U19282 (N_19282,N_16288,N_16805);
nand U19283 (N_19283,N_17858,N_17245);
xor U19284 (N_19284,N_16926,N_17219);
nor U19285 (N_19285,N_16799,N_16391);
nand U19286 (N_19286,N_17655,N_16106);
or U19287 (N_19287,N_16155,N_16319);
xor U19288 (N_19288,N_16139,N_17673);
nand U19289 (N_19289,N_17768,N_16943);
nand U19290 (N_19290,N_16171,N_17290);
nor U19291 (N_19291,N_17765,N_17296);
or U19292 (N_19292,N_16079,N_16183);
and U19293 (N_19293,N_17257,N_17180);
and U19294 (N_19294,N_17530,N_17121);
nor U19295 (N_19295,N_16304,N_17499);
or U19296 (N_19296,N_16644,N_17178);
nor U19297 (N_19297,N_16317,N_17226);
nand U19298 (N_19298,N_17881,N_17492);
nand U19299 (N_19299,N_17320,N_16712);
nand U19300 (N_19300,N_17275,N_17427);
xor U19301 (N_19301,N_16082,N_17515);
nor U19302 (N_19302,N_17088,N_17775);
and U19303 (N_19303,N_16654,N_16052);
nand U19304 (N_19304,N_17058,N_16650);
nor U19305 (N_19305,N_16649,N_17142);
nor U19306 (N_19306,N_16315,N_16966);
nor U19307 (N_19307,N_17560,N_17525);
nor U19308 (N_19308,N_16273,N_16880);
or U19309 (N_19309,N_16434,N_16121);
and U19310 (N_19310,N_16217,N_17598);
nand U19311 (N_19311,N_16615,N_17469);
nor U19312 (N_19312,N_16634,N_17964);
nand U19313 (N_19313,N_17846,N_16652);
nand U19314 (N_19314,N_16668,N_17731);
xor U19315 (N_19315,N_17110,N_17260);
nor U19316 (N_19316,N_17526,N_17134);
and U19317 (N_19317,N_16416,N_16904);
and U19318 (N_19318,N_16304,N_17590);
nor U19319 (N_19319,N_17694,N_16997);
nand U19320 (N_19320,N_16607,N_17486);
and U19321 (N_19321,N_17245,N_16191);
or U19322 (N_19322,N_17892,N_17321);
and U19323 (N_19323,N_17405,N_16523);
nand U19324 (N_19324,N_16760,N_16464);
and U19325 (N_19325,N_17228,N_17668);
or U19326 (N_19326,N_17782,N_17463);
and U19327 (N_19327,N_16351,N_16477);
nor U19328 (N_19328,N_17797,N_17896);
nand U19329 (N_19329,N_16206,N_16346);
nor U19330 (N_19330,N_17246,N_17437);
and U19331 (N_19331,N_16367,N_16785);
nand U19332 (N_19332,N_17612,N_17275);
and U19333 (N_19333,N_17377,N_17304);
xor U19334 (N_19334,N_17765,N_17962);
nor U19335 (N_19335,N_16219,N_17932);
and U19336 (N_19336,N_16676,N_17111);
xor U19337 (N_19337,N_16280,N_16548);
or U19338 (N_19338,N_17392,N_16356);
or U19339 (N_19339,N_17901,N_17942);
or U19340 (N_19340,N_17314,N_16166);
and U19341 (N_19341,N_17598,N_17832);
nor U19342 (N_19342,N_16907,N_16583);
or U19343 (N_19343,N_16378,N_16789);
nor U19344 (N_19344,N_16264,N_16732);
or U19345 (N_19345,N_17144,N_16578);
nand U19346 (N_19346,N_17162,N_17704);
nor U19347 (N_19347,N_17899,N_17221);
or U19348 (N_19348,N_17985,N_17027);
and U19349 (N_19349,N_16387,N_17201);
or U19350 (N_19350,N_16249,N_17816);
nand U19351 (N_19351,N_17671,N_16883);
xnor U19352 (N_19352,N_17216,N_17793);
or U19353 (N_19353,N_17899,N_17868);
nand U19354 (N_19354,N_17997,N_16360);
or U19355 (N_19355,N_17273,N_16240);
nor U19356 (N_19356,N_17716,N_16668);
nor U19357 (N_19357,N_17753,N_16718);
and U19358 (N_19358,N_16616,N_17421);
nor U19359 (N_19359,N_16685,N_17705);
or U19360 (N_19360,N_16335,N_16035);
or U19361 (N_19361,N_17217,N_16825);
and U19362 (N_19362,N_16875,N_16754);
or U19363 (N_19363,N_16046,N_16585);
xnor U19364 (N_19364,N_16331,N_16941);
nor U19365 (N_19365,N_17155,N_17300);
and U19366 (N_19366,N_17628,N_16245);
or U19367 (N_19367,N_17965,N_17210);
nor U19368 (N_19368,N_17098,N_16974);
and U19369 (N_19369,N_16801,N_17334);
nand U19370 (N_19370,N_16388,N_16191);
nand U19371 (N_19371,N_17104,N_17819);
xor U19372 (N_19372,N_16450,N_17469);
nor U19373 (N_19373,N_16421,N_16828);
or U19374 (N_19374,N_17009,N_16888);
or U19375 (N_19375,N_16093,N_16195);
nor U19376 (N_19376,N_16937,N_17997);
nor U19377 (N_19377,N_16159,N_16054);
and U19378 (N_19378,N_16811,N_16481);
nor U19379 (N_19379,N_17575,N_17387);
nor U19380 (N_19380,N_17195,N_16498);
nor U19381 (N_19381,N_17831,N_17340);
nor U19382 (N_19382,N_17398,N_16085);
or U19383 (N_19383,N_17511,N_16586);
xor U19384 (N_19384,N_17589,N_17859);
and U19385 (N_19385,N_16023,N_17651);
or U19386 (N_19386,N_16109,N_17511);
nor U19387 (N_19387,N_17166,N_16431);
and U19388 (N_19388,N_17362,N_17271);
nand U19389 (N_19389,N_16131,N_16776);
or U19390 (N_19390,N_17795,N_16670);
or U19391 (N_19391,N_16546,N_16217);
nand U19392 (N_19392,N_17222,N_17546);
and U19393 (N_19393,N_17180,N_17758);
nor U19394 (N_19394,N_17229,N_16259);
or U19395 (N_19395,N_16751,N_16485);
or U19396 (N_19396,N_16723,N_17870);
xnor U19397 (N_19397,N_16705,N_17181);
or U19398 (N_19398,N_17621,N_16075);
nor U19399 (N_19399,N_17004,N_17892);
or U19400 (N_19400,N_16765,N_16569);
or U19401 (N_19401,N_16300,N_17298);
xnor U19402 (N_19402,N_17111,N_17503);
nand U19403 (N_19403,N_16705,N_16764);
nor U19404 (N_19404,N_17430,N_17348);
or U19405 (N_19405,N_16467,N_17773);
nor U19406 (N_19406,N_17224,N_17565);
or U19407 (N_19407,N_16611,N_17460);
and U19408 (N_19408,N_17053,N_17693);
and U19409 (N_19409,N_16098,N_16126);
or U19410 (N_19410,N_16952,N_16893);
and U19411 (N_19411,N_17343,N_16075);
nor U19412 (N_19412,N_16752,N_17914);
or U19413 (N_19413,N_16674,N_16389);
nand U19414 (N_19414,N_17291,N_16030);
xor U19415 (N_19415,N_17943,N_16734);
nand U19416 (N_19416,N_16808,N_17529);
or U19417 (N_19417,N_17052,N_17857);
or U19418 (N_19418,N_17530,N_17445);
or U19419 (N_19419,N_16428,N_16429);
nor U19420 (N_19420,N_17907,N_17834);
or U19421 (N_19421,N_17889,N_16293);
and U19422 (N_19422,N_16474,N_16929);
xor U19423 (N_19423,N_16592,N_17437);
nor U19424 (N_19424,N_16474,N_16132);
nand U19425 (N_19425,N_17704,N_17713);
nor U19426 (N_19426,N_17466,N_16199);
or U19427 (N_19427,N_17589,N_17330);
or U19428 (N_19428,N_17557,N_17320);
or U19429 (N_19429,N_17037,N_17378);
nor U19430 (N_19430,N_17378,N_17266);
nand U19431 (N_19431,N_16838,N_17949);
nand U19432 (N_19432,N_16446,N_17508);
or U19433 (N_19433,N_17376,N_17321);
or U19434 (N_19434,N_16641,N_17109);
and U19435 (N_19435,N_17335,N_16340);
or U19436 (N_19436,N_16713,N_16968);
or U19437 (N_19437,N_17996,N_17894);
nand U19438 (N_19438,N_16629,N_16646);
or U19439 (N_19439,N_17976,N_17741);
nand U19440 (N_19440,N_16781,N_16536);
nor U19441 (N_19441,N_17888,N_17533);
or U19442 (N_19442,N_16456,N_16216);
or U19443 (N_19443,N_17250,N_17809);
xor U19444 (N_19444,N_17790,N_16017);
nor U19445 (N_19445,N_16402,N_16985);
and U19446 (N_19446,N_17102,N_17676);
and U19447 (N_19447,N_16683,N_16012);
or U19448 (N_19448,N_17074,N_17466);
nor U19449 (N_19449,N_17108,N_16836);
or U19450 (N_19450,N_16744,N_17766);
and U19451 (N_19451,N_16112,N_16676);
nor U19452 (N_19452,N_16792,N_16395);
xor U19453 (N_19453,N_17725,N_16370);
nand U19454 (N_19454,N_17538,N_17247);
and U19455 (N_19455,N_17004,N_16678);
or U19456 (N_19456,N_17555,N_16880);
nand U19457 (N_19457,N_16961,N_16259);
nand U19458 (N_19458,N_16237,N_17998);
nand U19459 (N_19459,N_17832,N_17560);
nor U19460 (N_19460,N_16083,N_16677);
and U19461 (N_19461,N_17483,N_16755);
or U19462 (N_19462,N_16291,N_16722);
nor U19463 (N_19463,N_17396,N_16287);
and U19464 (N_19464,N_16113,N_16769);
nor U19465 (N_19465,N_17430,N_17763);
nor U19466 (N_19466,N_17911,N_16845);
nand U19467 (N_19467,N_17413,N_17871);
or U19468 (N_19468,N_16783,N_17780);
nand U19469 (N_19469,N_17135,N_17380);
and U19470 (N_19470,N_17252,N_16001);
nor U19471 (N_19471,N_17990,N_16865);
or U19472 (N_19472,N_16613,N_16916);
xor U19473 (N_19473,N_16135,N_16369);
and U19474 (N_19474,N_16448,N_16484);
nor U19475 (N_19475,N_17552,N_16394);
or U19476 (N_19476,N_17352,N_16740);
and U19477 (N_19477,N_16613,N_17679);
nand U19478 (N_19478,N_17902,N_16204);
and U19479 (N_19479,N_17406,N_17108);
nand U19480 (N_19480,N_17029,N_16915);
nor U19481 (N_19481,N_16252,N_16989);
nand U19482 (N_19482,N_17002,N_17519);
nand U19483 (N_19483,N_16649,N_16134);
nor U19484 (N_19484,N_16484,N_16148);
or U19485 (N_19485,N_16804,N_16153);
or U19486 (N_19486,N_16376,N_17131);
nor U19487 (N_19487,N_17710,N_17126);
and U19488 (N_19488,N_16954,N_16347);
or U19489 (N_19489,N_17281,N_17622);
nor U19490 (N_19490,N_16683,N_16827);
nor U19491 (N_19491,N_17366,N_17995);
nand U19492 (N_19492,N_17079,N_16083);
nand U19493 (N_19493,N_16980,N_17303);
nor U19494 (N_19494,N_16229,N_16492);
nor U19495 (N_19495,N_17791,N_17037);
or U19496 (N_19496,N_17755,N_17936);
nand U19497 (N_19497,N_17270,N_17254);
nand U19498 (N_19498,N_17041,N_17162);
or U19499 (N_19499,N_16670,N_17859);
nor U19500 (N_19500,N_16961,N_17574);
xor U19501 (N_19501,N_16116,N_16625);
xnor U19502 (N_19502,N_16916,N_17106);
nor U19503 (N_19503,N_17556,N_17117);
nor U19504 (N_19504,N_16503,N_16294);
nand U19505 (N_19505,N_16908,N_17732);
and U19506 (N_19506,N_16336,N_17456);
nand U19507 (N_19507,N_17879,N_16886);
nor U19508 (N_19508,N_17705,N_17517);
nor U19509 (N_19509,N_16444,N_17234);
nor U19510 (N_19510,N_16635,N_16579);
nand U19511 (N_19511,N_16758,N_16309);
and U19512 (N_19512,N_16197,N_17946);
nand U19513 (N_19513,N_17257,N_17259);
or U19514 (N_19514,N_17601,N_16803);
xor U19515 (N_19515,N_17942,N_16154);
and U19516 (N_19516,N_16296,N_16627);
or U19517 (N_19517,N_16202,N_17072);
nor U19518 (N_19518,N_16896,N_16524);
or U19519 (N_19519,N_17112,N_17963);
nor U19520 (N_19520,N_16036,N_16255);
nand U19521 (N_19521,N_17628,N_17032);
nand U19522 (N_19522,N_16021,N_17433);
xor U19523 (N_19523,N_17529,N_16305);
or U19524 (N_19524,N_16631,N_16479);
and U19525 (N_19525,N_17649,N_17664);
nor U19526 (N_19526,N_17567,N_16229);
xnor U19527 (N_19527,N_16152,N_16722);
nor U19528 (N_19528,N_16384,N_16160);
nand U19529 (N_19529,N_17077,N_16757);
or U19530 (N_19530,N_17975,N_17879);
nor U19531 (N_19531,N_16277,N_17249);
nand U19532 (N_19532,N_17682,N_17251);
or U19533 (N_19533,N_17926,N_17416);
xor U19534 (N_19534,N_17831,N_16032);
xor U19535 (N_19535,N_17665,N_16086);
nor U19536 (N_19536,N_17842,N_17027);
nand U19537 (N_19537,N_16856,N_16731);
and U19538 (N_19538,N_17052,N_16745);
or U19539 (N_19539,N_16453,N_16873);
or U19540 (N_19540,N_16182,N_16438);
nand U19541 (N_19541,N_17833,N_17090);
or U19542 (N_19542,N_17519,N_16913);
and U19543 (N_19543,N_17356,N_16278);
nor U19544 (N_19544,N_17949,N_16052);
xnor U19545 (N_19545,N_16223,N_17832);
nand U19546 (N_19546,N_17767,N_16671);
nor U19547 (N_19547,N_17205,N_16010);
or U19548 (N_19548,N_16579,N_16158);
nor U19549 (N_19549,N_17399,N_17526);
nand U19550 (N_19550,N_16064,N_16424);
nand U19551 (N_19551,N_16831,N_17669);
or U19552 (N_19552,N_17885,N_17427);
nor U19553 (N_19553,N_17663,N_17688);
nor U19554 (N_19554,N_17657,N_17991);
and U19555 (N_19555,N_16663,N_17075);
or U19556 (N_19556,N_16364,N_16750);
or U19557 (N_19557,N_16591,N_16102);
nor U19558 (N_19558,N_17088,N_17508);
nand U19559 (N_19559,N_17945,N_17437);
nand U19560 (N_19560,N_17258,N_17993);
and U19561 (N_19561,N_16369,N_16308);
nor U19562 (N_19562,N_16366,N_16901);
and U19563 (N_19563,N_17641,N_17130);
nand U19564 (N_19564,N_17174,N_17209);
nand U19565 (N_19565,N_17893,N_17355);
xnor U19566 (N_19566,N_16885,N_16994);
nor U19567 (N_19567,N_17335,N_16380);
nor U19568 (N_19568,N_16047,N_16976);
nand U19569 (N_19569,N_16514,N_16817);
and U19570 (N_19570,N_17077,N_17749);
or U19571 (N_19571,N_16498,N_17976);
nand U19572 (N_19572,N_16764,N_17832);
or U19573 (N_19573,N_16140,N_17751);
and U19574 (N_19574,N_17422,N_16069);
nand U19575 (N_19575,N_16891,N_17123);
nand U19576 (N_19576,N_17678,N_16165);
nor U19577 (N_19577,N_17276,N_16699);
or U19578 (N_19578,N_17106,N_17009);
xor U19579 (N_19579,N_16976,N_16680);
nor U19580 (N_19580,N_16207,N_17980);
or U19581 (N_19581,N_16634,N_17987);
nor U19582 (N_19582,N_16016,N_16116);
or U19583 (N_19583,N_16982,N_17229);
xor U19584 (N_19584,N_16614,N_17039);
or U19585 (N_19585,N_16146,N_16901);
xor U19586 (N_19586,N_16910,N_17925);
nor U19587 (N_19587,N_17604,N_17416);
xor U19588 (N_19588,N_16101,N_16860);
or U19589 (N_19589,N_16933,N_17654);
or U19590 (N_19590,N_16571,N_17576);
or U19591 (N_19591,N_17018,N_16252);
and U19592 (N_19592,N_17723,N_16671);
or U19593 (N_19593,N_17067,N_16340);
and U19594 (N_19594,N_17970,N_17042);
nor U19595 (N_19595,N_16634,N_17546);
nand U19596 (N_19596,N_16908,N_16161);
and U19597 (N_19597,N_17037,N_17224);
nand U19598 (N_19598,N_17130,N_17883);
nor U19599 (N_19599,N_16185,N_17369);
nand U19600 (N_19600,N_16020,N_17216);
and U19601 (N_19601,N_16491,N_17886);
nand U19602 (N_19602,N_17510,N_17680);
nand U19603 (N_19603,N_16660,N_16278);
or U19604 (N_19604,N_16061,N_17768);
nor U19605 (N_19605,N_17971,N_17554);
nor U19606 (N_19606,N_17850,N_17141);
nor U19607 (N_19607,N_17924,N_16069);
and U19608 (N_19608,N_16362,N_17034);
nand U19609 (N_19609,N_17241,N_16588);
xor U19610 (N_19610,N_17125,N_17323);
nor U19611 (N_19611,N_16100,N_17895);
nand U19612 (N_19612,N_16723,N_16003);
nand U19613 (N_19613,N_17295,N_16922);
and U19614 (N_19614,N_16354,N_16768);
and U19615 (N_19615,N_17105,N_17985);
xor U19616 (N_19616,N_16877,N_17688);
nor U19617 (N_19617,N_17875,N_16314);
or U19618 (N_19618,N_17397,N_16259);
and U19619 (N_19619,N_16827,N_16080);
and U19620 (N_19620,N_17005,N_17267);
or U19621 (N_19621,N_17293,N_17429);
or U19622 (N_19622,N_17802,N_16463);
or U19623 (N_19623,N_16907,N_16877);
nor U19624 (N_19624,N_16534,N_17727);
nand U19625 (N_19625,N_16296,N_16451);
and U19626 (N_19626,N_16711,N_17466);
xnor U19627 (N_19627,N_17576,N_17868);
or U19628 (N_19628,N_17688,N_17855);
nand U19629 (N_19629,N_17893,N_16339);
nand U19630 (N_19630,N_16072,N_17951);
or U19631 (N_19631,N_16657,N_17395);
or U19632 (N_19632,N_16086,N_16454);
and U19633 (N_19633,N_17760,N_17700);
nor U19634 (N_19634,N_17986,N_16099);
xor U19635 (N_19635,N_17843,N_16647);
or U19636 (N_19636,N_17296,N_16734);
nand U19637 (N_19637,N_16712,N_17282);
or U19638 (N_19638,N_17348,N_17908);
or U19639 (N_19639,N_17680,N_16750);
nor U19640 (N_19640,N_17399,N_17447);
nor U19641 (N_19641,N_16107,N_16665);
nor U19642 (N_19642,N_16068,N_16502);
and U19643 (N_19643,N_17536,N_16595);
nand U19644 (N_19644,N_16505,N_16099);
nor U19645 (N_19645,N_17075,N_17682);
or U19646 (N_19646,N_16523,N_17582);
and U19647 (N_19647,N_17054,N_17914);
nor U19648 (N_19648,N_16696,N_17536);
xnor U19649 (N_19649,N_16016,N_17026);
and U19650 (N_19650,N_17826,N_17074);
and U19651 (N_19651,N_17771,N_17610);
nor U19652 (N_19652,N_17123,N_17681);
or U19653 (N_19653,N_16531,N_16141);
nor U19654 (N_19654,N_16837,N_16416);
nor U19655 (N_19655,N_16085,N_16786);
nor U19656 (N_19656,N_17430,N_16433);
nand U19657 (N_19657,N_16622,N_16571);
and U19658 (N_19658,N_17180,N_16019);
nand U19659 (N_19659,N_16715,N_17817);
nand U19660 (N_19660,N_16870,N_17638);
and U19661 (N_19661,N_17771,N_16793);
or U19662 (N_19662,N_17056,N_17583);
or U19663 (N_19663,N_16384,N_17182);
and U19664 (N_19664,N_16018,N_16840);
nand U19665 (N_19665,N_16238,N_17134);
and U19666 (N_19666,N_16189,N_16512);
and U19667 (N_19667,N_17271,N_16950);
xor U19668 (N_19668,N_16766,N_17093);
nor U19669 (N_19669,N_16354,N_17083);
and U19670 (N_19670,N_16103,N_17352);
nor U19671 (N_19671,N_17499,N_16699);
nor U19672 (N_19672,N_17662,N_17083);
nand U19673 (N_19673,N_16193,N_17579);
or U19674 (N_19674,N_17316,N_17851);
nor U19675 (N_19675,N_17767,N_17607);
or U19676 (N_19676,N_17180,N_17539);
and U19677 (N_19677,N_16001,N_16461);
or U19678 (N_19678,N_16641,N_17562);
nand U19679 (N_19679,N_16228,N_17969);
xnor U19680 (N_19680,N_17629,N_16858);
nor U19681 (N_19681,N_16272,N_17026);
nand U19682 (N_19682,N_17011,N_16224);
or U19683 (N_19683,N_16434,N_17551);
xor U19684 (N_19684,N_17176,N_16493);
nor U19685 (N_19685,N_17085,N_17353);
nand U19686 (N_19686,N_17362,N_16479);
and U19687 (N_19687,N_16856,N_16982);
or U19688 (N_19688,N_16198,N_16882);
and U19689 (N_19689,N_16930,N_17830);
nand U19690 (N_19690,N_17585,N_16661);
nor U19691 (N_19691,N_16357,N_16480);
nor U19692 (N_19692,N_17811,N_16173);
nand U19693 (N_19693,N_16358,N_17293);
nor U19694 (N_19694,N_17783,N_17147);
nor U19695 (N_19695,N_17295,N_17107);
nand U19696 (N_19696,N_17637,N_17376);
nor U19697 (N_19697,N_17705,N_16579);
xor U19698 (N_19698,N_17742,N_17769);
nor U19699 (N_19699,N_17979,N_17852);
or U19700 (N_19700,N_16285,N_16820);
and U19701 (N_19701,N_17050,N_17217);
and U19702 (N_19702,N_16051,N_17246);
xor U19703 (N_19703,N_17785,N_16383);
nand U19704 (N_19704,N_17254,N_17696);
xnor U19705 (N_19705,N_17702,N_17323);
and U19706 (N_19706,N_17112,N_16873);
and U19707 (N_19707,N_16778,N_16324);
xnor U19708 (N_19708,N_16603,N_16432);
nand U19709 (N_19709,N_16065,N_16095);
nor U19710 (N_19710,N_17904,N_16460);
nor U19711 (N_19711,N_16861,N_16275);
nand U19712 (N_19712,N_17314,N_17916);
nor U19713 (N_19713,N_16923,N_16946);
nand U19714 (N_19714,N_17823,N_17874);
or U19715 (N_19715,N_16804,N_16475);
and U19716 (N_19716,N_16190,N_17326);
nand U19717 (N_19717,N_17569,N_16252);
or U19718 (N_19718,N_16108,N_17022);
or U19719 (N_19719,N_17272,N_16974);
and U19720 (N_19720,N_17149,N_17929);
or U19721 (N_19721,N_17910,N_17697);
or U19722 (N_19722,N_16728,N_16186);
nor U19723 (N_19723,N_16145,N_16451);
or U19724 (N_19724,N_16275,N_17823);
nand U19725 (N_19725,N_16134,N_17252);
or U19726 (N_19726,N_16460,N_16591);
xor U19727 (N_19727,N_16283,N_17293);
and U19728 (N_19728,N_16489,N_16251);
nor U19729 (N_19729,N_17902,N_16288);
nand U19730 (N_19730,N_17993,N_16065);
and U19731 (N_19731,N_16461,N_17820);
or U19732 (N_19732,N_17029,N_17014);
xnor U19733 (N_19733,N_17326,N_17187);
and U19734 (N_19734,N_16014,N_16644);
or U19735 (N_19735,N_16112,N_17297);
and U19736 (N_19736,N_17696,N_17275);
nand U19737 (N_19737,N_17670,N_16481);
nand U19738 (N_19738,N_17747,N_16119);
or U19739 (N_19739,N_16878,N_16276);
nor U19740 (N_19740,N_17541,N_16464);
and U19741 (N_19741,N_17552,N_16985);
nand U19742 (N_19742,N_16520,N_17820);
or U19743 (N_19743,N_16902,N_16725);
and U19744 (N_19744,N_17008,N_17342);
xor U19745 (N_19745,N_16833,N_16035);
nand U19746 (N_19746,N_17510,N_17525);
and U19747 (N_19747,N_17172,N_16876);
nor U19748 (N_19748,N_16723,N_17699);
nor U19749 (N_19749,N_17121,N_17879);
nand U19750 (N_19750,N_17606,N_16979);
nor U19751 (N_19751,N_16580,N_17568);
and U19752 (N_19752,N_16750,N_16210);
nand U19753 (N_19753,N_17396,N_17908);
nor U19754 (N_19754,N_16698,N_17956);
nand U19755 (N_19755,N_16010,N_16943);
nor U19756 (N_19756,N_16805,N_16158);
and U19757 (N_19757,N_17000,N_16810);
nand U19758 (N_19758,N_16268,N_16159);
nand U19759 (N_19759,N_16746,N_17563);
xor U19760 (N_19760,N_17798,N_16014);
xnor U19761 (N_19761,N_17218,N_17015);
or U19762 (N_19762,N_16138,N_17041);
or U19763 (N_19763,N_16518,N_16834);
xnor U19764 (N_19764,N_16574,N_16343);
and U19765 (N_19765,N_16679,N_16169);
nor U19766 (N_19766,N_16707,N_17080);
and U19767 (N_19767,N_17924,N_17756);
nand U19768 (N_19768,N_16596,N_17526);
or U19769 (N_19769,N_17367,N_17827);
or U19770 (N_19770,N_16432,N_17684);
nor U19771 (N_19771,N_17332,N_16430);
nand U19772 (N_19772,N_16695,N_17083);
and U19773 (N_19773,N_17244,N_16972);
and U19774 (N_19774,N_16096,N_16331);
nor U19775 (N_19775,N_16831,N_17443);
nor U19776 (N_19776,N_17150,N_16504);
or U19777 (N_19777,N_17669,N_17533);
nor U19778 (N_19778,N_17764,N_17527);
and U19779 (N_19779,N_17382,N_17664);
or U19780 (N_19780,N_16304,N_16203);
and U19781 (N_19781,N_17638,N_16655);
or U19782 (N_19782,N_16575,N_17982);
nor U19783 (N_19783,N_17975,N_17586);
or U19784 (N_19784,N_16041,N_17976);
or U19785 (N_19785,N_16464,N_16451);
xnor U19786 (N_19786,N_16929,N_16688);
and U19787 (N_19787,N_16959,N_16651);
xor U19788 (N_19788,N_16301,N_16390);
nor U19789 (N_19789,N_17672,N_16248);
nand U19790 (N_19790,N_16357,N_16196);
or U19791 (N_19791,N_16347,N_16303);
nor U19792 (N_19792,N_16703,N_16483);
nor U19793 (N_19793,N_16146,N_16563);
or U19794 (N_19794,N_16703,N_17666);
nor U19795 (N_19795,N_17268,N_17778);
or U19796 (N_19796,N_17117,N_16871);
nand U19797 (N_19797,N_17440,N_17419);
and U19798 (N_19798,N_17588,N_17032);
nand U19799 (N_19799,N_16102,N_17848);
and U19800 (N_19800,N_16046,N_16010);
and U19801 (N_19801,N_17518,N_17517);
and U19802 (N_19802,N_16390,N_16774);
nand U19803 (N_19803,N_16605,N_16240);
nand U19804 (N_19804,N_17527,N_17661);
or U19805 (N_19805,N_17397,N_16764);
xor U19806 (N_19806,N_17970,N_16500);
or U19807 (N_19807,N_17891,N_16760);
and U19808 (N_19808,N_17744,N_16296);
nand U19809 (N_19809,N_16122,N_17499);
or U19810 (N_19810,N_17451,N_16397);
or U19811 (N_19811,N_16778,N_16130);
nor U19812 (N_19812,N_16603,N_17318);
and U19813 (N_19813,N_16817,N_17514);
and U19814 (N_19814,N_17416,N_17264);
and U19815 (N_19815,N_17455,N_17573);
nand U19816 (N_19816,N_16786,N_16264);
xnor U19817 (N_19817,N_17373,N_16169);
and U19818 (N_19818,N_16773,N_17889);
and U19819 (N_19819,N_17827,N_16421);
and U19820 (N_19820,N_17790,N_17701);
xnor U19821 (N_19821,N_16997,N_16577);
or U19822 (N_19822,N_16280,N_17624);
nor U19823 (N_19823,N_16368,N_17199);
xor U19824 (N_19824,N_16595,N_16276);
nand U19825 (N_19825,N_16955,N_17805);
nor U19826 (N_19826,N_16570,N_17380);
or U19827 (N_19827,N_17772,N_17331);
or U19828 (N_19828,N_16739,N_17488);
nand U19829 (N_19829,N_16430,N_16348);
nor U19830 (N_19830,N_17203,N_17086);
and U19831 (N_19831,N_16746,N_16908);
or U19832 (N_19832,N_16633,N_16204);
nor U19833 (N_19833,N_16513,N_17877);
and U19834 (N_19834,N_16860,N_17719);
xor U19835 (N_19835,N_17908,N_16603);
and U19836 (N_19836,N_17796,N_16835);
nand U19837 (N_19837,N_17078,N_17959);
nor U19838 (N_19838,N_17322,N_17401);
nor U19839 (N_19839,N_16825,N_16065);
and U19840 (N_19840,N_16302,N_17378);
nand U19841 (N_19841,N_17855,N_17086);
nand U19842 (N_19842,N_17531,N_16257);
nor U19843 (N_19843,N_17962,N_16711);
or U19844 (N_19844,N_16217,N_16135);
and U19845 (N_19845,N_17111,N_17847);
nor U19846 (N_19846,N_17279,N_16275);
or U19847 (N_19847,N_16599,N_17973);
nand U19848 (N_19848,N_17866,N_16297);
nand U19849 (N_19849,N_17619,N_16881);
and U19850 (N_19850,N_17651,N_17758);
nand U19851 (N_19851,N_16045,N_17946);
and U19852 (N_19852,N_17054,N_17978);
and U19853 (N_19853,N_17528,N_16343);
xor U19854 (N_19854,N_17150,N_16166);
nand U19855 (N_19855,N_17849,N_16339);
xnor U19856 (N_19856,N_17393,N_17728);
nand U19857 (N_19857,N_16445,N_16412);
or U19858 (N_19858,N_16507,N_17003);
or U19859 (N_19859,N_16911,N_17670);
nor U19860 (N_19860,N_17080,N_17960);
nand U19861 (N_19861,N_17727,N_16661);
or U19862 (N_19862,N_16378,N_16748);
and U19863 (N_19863,N_16499,N_16004);
or U19864 (N_19864,N_16084,N_16357);
nor U19865 (N_19865,N_17432,N_17829);
nand U19866 (N_19866,N_17373,N_17238);
or U19867 (N_19867,N_16945,N_17910);
or U19868 (N_19868,N_17496,N_17769);
or U19869 (N_19869,N_16806,N_17962);
or U19870 (N_19870,N_17253,N_17916);
nor U19871 (N_19871,N_17998,N_17120);
nor U19872 (N_19872,N_16462,N_17312);
or U19873 (N_19873,N_16381,N_16289);
nor U19874 (N_19874,N_16384,N_16218);
nand U19875 (N_19875,N_16384,N_16671);
and U19876 (N_19876,N_16212,N_17537);
or U19877 (N_19877,N_16468,N_16148);
nand U19878 (N_19878,N_17840,N_17811);
nor U19879 (N_19879,N_16507,N_17389);
and U19880 (N_19880,N_17485,N_17835);
nor U19881 (N_19881,N_16237,N_16745);
nor U19882 (N_19882,N_17331,N_16876);
and U19883 (N_19883,N_17214,N_17644);
xor U19884 (N_19884,N_16246,N_16572);
nand U19885 (N_19885,N_16879,N_16390);
and U19886 (N_19886,N_17930,N_17277);
and U19887 (N_19887,N_16457,N_17919);
nor U19888 (N_19888,N_17188,N_16869);
and U19889 (N_19889,N_16069,N_16341);
xnor U19890 (N_19890,N_16833,N_17052);
nand U19891 (N_19891,N_17285,N_16694);
or U19892 (N_19892,N_16178,N_17531);
nor U19893 (N_19893,N_16016,N_16087);
or U19894 (N_19894,N_16465,N_16905);
xor U19895 (N_19895,N_17262,N_17410);
and U19896 (N_19896,N_16178,N_16697);
and U19897 (N_19897,N_17335,N_16533);
nor U19898 (N_19898,N_16354,N_17075);
nor U19899 (N_19899,N_16780,N_17628);
and U19900 (N_19900,N_17352,N_17088);
or U19901 (N_19901,N_17152,N_16405);
and U19902 (N_19902,N_16475,N_17035);
nand U19903 (N_19903,N_17224,N_16247);
nand U19904 (N_19904,N_16372,N_16532);
or U19905 (N_19905,N_16235,N_16074);
nor U19906 (N_19906,N_16094,N_16012);
nand U19907 (N_19907,N_16405,N_16410);
xor U19908 (N_19908,N_16380,N_17057);
nand U19909 (N_19909,N_16753,N_17102);
and U19910 (N_19910,N_17918,N_16533);
nand U19911 (N_19911,N_16243,N_16130);
and U19912 (N_19912,N_16166,N_16721);
or U19913 (N_19913,N_16859,N_16456);
or U19914 (N_19914,N_17378,N_16035);
nand U19915 (N_19915,N_17437,N_17261);
or U19916 (N_19916,N_17344,N_16107);
and U19917 (N_19917,N_17884,N_16024);
xnor U19918 (N_19918,N_16233,N_16678);
nor U19919 (N_19919,N_16581,N_17480);
and U19920 (N_19920,N_16545,N_17891);
nor U19921 (N_19921,N_17406,N_16765);
nor U19922 (N_19922,N_16616,N_16360);
nor U19923 (N_19923,N_17013,N_16452);
or U19924 (N_19924,N_16787,N_16275);
or U19925 (N_19925,N_17714,N_17254);
or U19926 (N_19926,N_16381,N_16397);
nand U19927 (N_19927,N_16453,N_16811);
nand U19928 (N_19928,N_16323,N_17658);
or U19929 (N_19929,N_16461,N_17603);
and U19930 (N_19930,N_17814,N_16990);
or U19931 (N_19931,N_17948,N_16818);
nand U19932 (N_19932,N_16222,N_16094);
nand U19933 (N_19933,N_16729,N_17344);
nand U19934 (N_19934,N_17128,N_16956);
nor U19935 (N_19935,N_17039,N_17100);
nand U19936 (N_19936,N_16624,N_17808);
nor U19937 (N_19937,N_16108,N_16029);
or U19938 (N_19938,N_17293,N_17289);
or U19939 (N_19939,N_16168,N_16357);
nor U19940 (N_19940,N_16599,N_17866);
nor U19941 (N_19941,N_17482,N_17848);
nor U19942 (N_19942,N_17458,N_17359);
nor U19943 (N_19943,N_17372,N_16130);
nand U19944 (N_19944,N_17033,N_17920);
and U19945 (N_19945,N_16935,N_16639);
nor U19946 (N_19946,N_17863,N_16562);
xnor U19947 (N_19947,N_16390,N_16547);
nor U19948 (N_19948,N_16478,N_17285);
nor U19949 (N_19949,N_16113,N_17926);
or U19950 (N_19950,N_16087,N_17341);
and U19951 (N_19951,N_16406,N_16015);
or U19952 (N_19952,N_17285,N_17020);
nor U19953 (N_19953,N_17463,N_17269);
nor U19954 (N_19954,N_16662,N_16252);
or U19955 (N_19955,N_16186,N_16960);
nor U19956 (N_19956,N_16999,N_17488);
nand U19957 (N_19957,N_17814,N_16412);
xnor U19958 (N_19958,N_16260,N_17165);
or U19959 (N_19959,N_16504,N_17025);
or U19960 (N_19960,N_17309,N_16051);
and U19961 (N_19961,N_17046,N_17143);
or U19962 (N_19962,N_17116,N_17336);
nor U19963 (N_19963,N_16214,N_17213);
nor U19964 (N_19964,N_16632,N_17496);
xor U19965 (N_19965,N_16055,N_17478);
nand U19966 (N_19966,N_16755,N_16261);
nand U19967 (N_19967,N_16909,N_17504);
nand U19968 (N_19968,N_16842,N_17474);
or U19969 (N_19969,N_16003,N_16081);
or U19970 (N_19970,N_17588,N_17897);
or U19971 (N_19971,N_16373,N_17156);
and U19972 (N_19972,N_17152,N_16449);
nand U19973 (N_19973,N_17345,N_16770);
nor U19974 (N_19974,N_16495,N_17707);
and U19975 (N_19975,N_17735,N_16741);
nor U19976 (N_19976,N_17302,N_16374);
and U19977 (N_19977,N_17489,N_16337);
or U19978 (N_19978,N_17261,N_16869);
nor U19979 (N_19979,N_16312,N_17223);
and U19980 (N_19980,N_16954,N_17155);
nor U19981 (N_19981,N_17261,N_16438);
or U19982 (N_19982,N_16907,N_16155);
nor U19983 (N_19983,N_17101,N_17386);
or U19984 (N_19984,N_16540,N_16340);
or U19985 (N_19985,N_16621,N_17230);
xnor U19986 (N_19986,N_16369,N_16138);
nor U19987 (N_19987,N_16466,N_17119);
xnor U19988 (N_19988,N_16100,N_17598);
and U19989 (N_19989,N_16446,N_17642);
and U19990 (N_19990,N_16435,N_16432);
or U19991 (N_19991,N_17091,N_16160);
nand U19992 (N_19992,N_16784,N_16797);
and U19993 (N_19993,N_17686,N_17239);
xor U19994 (N_19994,N_17125,N_16632);
and U19995 (N_19995,N_16680,N_17777);
and U19996 (N_19996,N_16603,N_17199);
xnor U19997 (N_19997,N_17759,N_17811);
or U19998 (N_19998,N_16724,N_16411);
and U19999 (N_19999,N_16689,N_17396);
nand UO_0 (O_0,N_18297,N_18873);
nor UO_1 (O_1,N_18513,N_19428);
and UO_2 (O_2,N_18868,N_18518);
xor UO_3 (O_3,N_19856,N_18546);
or UO_4 (O_4,N_19095,N_19016);
and UO_5 (O_5,N_18285,N_19094);
or UO_6 (O_6,N_18826,N_18955);
nor UO_7 (O_7,N_18969,N_18569);
or UO_8 (O_8,N_19224,N_19763);
nand UO_9 (O_9,N_19340,N_19171);
nor UO_10 (O_10,N_19100,N_18005);
nor UO_11 (O_11,N_19329,N_19883);
and UO_12 (O_12,N_19425,N_19679);
and UO_13 (O_13,N_18422,N_19824);
and UO_14 (O_14,N_18773,N_18371);
or UO_15 (O_15,N_19130,N_18515);
and UO_16 (O_16,N_19910,N_19962);
or UO_17 (O_17,N_18666,N_18038);
or UO_18 (O_18,N_18935,N_18416);
and UO_19 (O_19,N_18676,N_19302);
xor UO_20 (O_20,N_18428,N_18477);
or UO_21 (O_21,N_18305,N_19288);
and UO_22 (O_22,N_19718,N_19027);
and UO_23 (O_23,N_19449,N_19595);
and UO_24 (O_24,N_18255,N_19010);
or UO_25 (O_25,N_18014,N_18975);
or UO_26 (O_26,N_18204,N_18957);
nor UO_27 (O_27,N_19989,N_19479);
and UO_28 (O_28,N_18349,N_19032);
nor UO_29 (O_29,N_19054,N_19212);
and UO_30 (O_30,N_18720,N_18397);
nand UO_31 (O_31,N_18965,N_18224);
nand UO_32 (O_32,N_19018,N_19904);
nand UO_33 (O_33,N_19167,N_19659);
nand UO_34 (O_34,N_19141,N_19771);
or UO_35 (O_35,N_19639,N_19324);
nor UO_36 (O_36,N_18690,N_18077);
xor UO_37 (O_37,N_18537,N_18335);
nor UO_38 (O_38,N_19124,N_18409);
nand UO_39 (O_39,N_19971,N_18697);
xor UO_40 (O_40,N_18925,N_19313);
and UO_41 (O_41,N_18391,N_19704);
and UO_42 (O_42,N_18509,N_18115);
and UO_43 (O_43,N_18384,N_18942);
xnor UO_44 (O_44,N_18628,N_19940);
and UO_45 (O_45,N_19678,N_19181);
nor UO_46 (O_46,N_19118,N_18577);
and UO_47 (O_47,N_18311,N_18402);
nand UO_48 (O_48,N_19119,N_18583);
or UO_49 (O_49,N_18644,N_19218);
nand UO_50 (O_50,N_19614,N_18652);
nand UO_51 (O_51,N_19539,N_18344);
or UO_52 (O_52,N_19490,N_18619);
nor UO_53 (O_53,N_18294,N_18387);
nor UO_54 (O_54,N_19781,N_19069);
or UO_55 (O_55,N_18341,N_19657);
and UO_56 (O_56,N_19993,N_18146);
xor UO_57 (O_57,N_18497,N_18367);
xor UO_58 (O_58,N_19246,N_18640);
nand UO_59 (O_59,N_18603,N_18951);
and UO_60 (O_60,N_19881,N_18700);
xnor UO_61 (O_61,N_18261,N_18623);
nand UO_62 (O_62,N_19626,N_19404);
nor UO_63 (O_63,N_18492,N_18823);
or UO_64 (O_64,N_18597,N_19629);
nor UO_65 (O_65,N_18370,N_19273);
or UO_66 (O_66,N_19295,N_18635);
nand UO_67 (O_67,N_18911,N_19000);
and UO_68 (O_68,N_18306,N_18553);
nand UO_69 (O_69,N_19685,N_18858);
nor UO_70 (O_70,N_19876,N_19353);
xor UO_71 (O_71,N_19031,N_19129);
or UO_72 (O_72,N_19241,N_19536);
and UO_73 (O_73,N_18173,N_18634);
or UO_74 (O_74,N_18704,N_19601);
or UO_75 (O_75,N_18326,N_18202);
or UO_76 (O_76,N_19366,N_18145);
or UO_77 (O_77,N_18753,N_19598);
and UO_78 (O_78,N_18070,N_18258);
nand UO_79 (O_79,N_19202,N_19476);
xnor UO_80 (O_80,N_19646,N_19277);
xor UO_81 (O_81,N_18209,N_19420);
nor UO_82 (O_82,N_19395,N_19761);
nor UO_83 (O_83,N_19645,N_18505);
nand UO_84 (O_84,N_19328,N_18804);
nor UO_85 (O_85,N_19445,N_19300);
and UO_86 (O_86,N_19801,N_18771);
nor UO_87 (O_87,N_19927,N_19928);
or UO_88 (O_88,N_19624,N_18315);
and UO_89 (O_89,N_18250,N_19930);
nand UO_90 (O_90,N_18502,N_18009);
nor UO_91 (O_91,N_19775,N_19529);
nor UO_92 (O_92,N_19486,N_19899);
or UO_93 (O_93,N_18671,N_19397);
nand UO_94 (O_94,N_19954,N_18716);
nand UO_95 (O_95,N_19905,N_19867);
and UO_96 (O_96,N_19534,N_18260);
or UO_97 (O_97,N_19964,N_19647);
xnor UO_98 (O_98,N_19034,N_19789);
or UO_99 (O_99,N_19333,N_18743);
xor UO_100 (O_100,N_18780,N_18986);
and UO_101 (O_101,N_19441,N_18216);
nor UO_102 (O_102,N_19496,N_18135);
and UO_103 (O_103,N_18223,N_19456);
nand UO_104 (O_104,N_18796,N_18061);
xor UO_105 (O_105,N_18050,N_19448);
nand UO_106 (O_106,N_18578,N_18020);
nor UO_107 (O_107,N_18721,N_18579);
or UO_108 (O_108,N_18920,N_18237);
xor UO_109 (O_109,N_18316,N_18827);
or UO_110 (O_110,N_19342,N_18760);
nor UO_111 (O_111,N_19274,N_18821);
and UO_112 (O_112,N_18724,N_18389);
xnor UO_113 (O_113,N_19713,N_19463);
nand UO_114 (O_114,N_19757,N_19041);
xor UO_115 (O_115,N_18133,N_19799);
nor UO_116 (O_116,N_18352,N_18775);
xor UO_117 (O_117,N_19430,N_19870);
nand UO_118 (O_118,N_19611,N_19363);
nand UO_119 (O_119,N_18803,N_18554);
and UO_120 (O_120,N_19874,N_19706);
and UO_121 (O_121,N_18762,N_19682);
nor UO_122 (O_122,N_18672,N_18067);
nor UO_123 (O_123,N_19811,N_18997);
or UO_124 (O_124,N_19432,N_18338);
nand UO_125 (O_125,N_19809,N_19773);
nand UO_126 (O_126,N_19816,N_19897);
nand UO_127 (O_127,N_18466,N_18137);
or UO_128 (O_128,N_19727,N_18144);
and UO_129 (O_129,N_19135,N_19879);
or UO_130 (O_130,N_18556,N_18914);
nor UO_131 (O_131,N_19569,N_19453);
xor UO_132 (O_132,N_18833,N_18369);
and UO_133 (O_133,N_18612,N_19409);
nand UO_134 (O_134,N_19935,N_19025);
xnor UO_135 (O_135,N_19527,N_18267);
nand UO_136 (O_136,N_18750,N_18439);
nor UO_137 (O_137,N_19146,N_18591);
and UO_138 (O_138,N_19908,N_18987);
xnor UO_139 (O_139,N_19631,N_18938);
nand UO_140 (O_140,N_18590,N_19513);
nand UO_141 (O_141,N_18586,N_18910);
xnor UO_142 (O_142,N_18820,N_19945);
or UO_143 (O_143,N_18811,N_18256);
xor UO_144 (O_144,N_19564,N_18484);
or UO_145 (O_145,N_19652,N_18318);
nor UO_146 (O_146,N_19958,N_19588);
nand UO_147 (O_147,N_18163,N_19132);
and UO_148 (O_148,N_19272,N_18878);
or UO_149 (O_149,N_19662,N_18795);
xor UO_150 (O_150,N_19755,N_18737);
or UO_151 (O_151,N_19518,N_18111);
nand UO_152 (O_152,N_18192,N_19907);
and UO_153 (O_153,N_18799,N_19963);
or UO_154 (O_154,N_19632,N_18874);
nand UO_155 (O_155,N_19081,N_19105);
and UO_156 (O_156,N_18363,N_18419);
xor UO_157 (O_157,N_19924,N_19177);
and UO_158 (O_158,N_18934,N_19627);
nor UO_159 (O_159,N_18931,N_18268);
or UO_160 (O_160,N_18296,N_18455);
or UO_161 (O_161,N_18980,N_18304);
and UO_162 (O_162,N_18128,N_18211);
xor UO_163 (O_163,N_18281,N_19866);
or UO_164 (O_164,N_19970,N_18968);
xnor UO_165 (O_165,N_19412,N_18136);
or UO_166 (O_166,N_19966,N_19644);
and UO_167 (O_167,N_18605,N_18901);
nand UO_168 (O_168,N_19304,N_18595);
nor UO_169 (O_169,N_18759,N_18127);
or UO_170 (O_170,N_19603,N_19190);
and UO_171 (O_171,N_18802,N_19509);
nor UO_172 (O_172,N_18152,N_19911);
nand UO_173 (O_173,N_19361,N_18731);
or UO_174 (O_174,N_18524,N_19394);
nand UO_175 (O_175,N_19919,N_18645);
xnor UO_176 (O_176,N_19227,N_18543);
nor UO_177 (O_177,N_19279,N_19591);
nand UO_178 (O_178,N_18824,N_19649);
or UO_179 (O_179,N_18200,N_19477);
nand UO_180 (O_180,N_19560,N_19112);
and UO_181 (O_181,N_19594,N_18157);
nor UO_182 (O_182,N_18435,N_18566);
or UO_183 (O_183,N_18024,N_19195);
xnor UO_184 (O_184,N_18138,N_19759);
or UO_185 (O_185,N_18186,N_18401);
or UO_186 (O_186,N_19111,N_19243);
nor UO_187 (O_187,N_19810,N_18169);
nand UO_188 (O_188,N_19680,N_18059);
or UO_189 (O_189,N_18060,N_18159);
nor UO_190 (O_190,N_19592,N_18573);
or UO_191 (O_191,N_19860,N_19040);
nor UO_192 (O_192,N_18673,N_18602);
and UO_193 (O_193,N_18840,N_19125);
or UO_194 (O_194,N_18984,N_19994);
nor UO_195 (O_195,N_19478,N_19826);
or UO_196 (O_196,N_19378,N_18839);
or UO_197 (O_197,N_18116,N_19869);
or UO_198 (O_198,N_19665,N_18065);
nand UO_199 (O_199,N_18610,N_19724);
or UO_200 (O_200,N_19732,N_18503);
nor UO_201 (O_201,N_19655,N_18426);
nand UO_202 (O_202,N_19312,N_19165);
or UO_203 (O_203,N_19499,N_18450);
and UO_204 (O_204,N_18630,N_19305);
nor UO_205 (O_205,N_19265,N_18461);
or UO_206 (O_206,N_19256,N_18632);
nand UO_207 (O_207,N_18471,N_18184);
nor UO_208 (O_208,N_19973,N_19712);
xor UO_209 (O_209,N_18860,N_19358);
nand UO_210 (O_210,N_19320,N_19127);
and UO_211 (O_211,N_18015,N_18841);
or UO_212 (O_212,N_19393,N_18896);
nor UO_213 (O_213,N_19604,N_18510);
nor UO_214 (O_214,N_19788,N_19939);
and UO_215 (O_215,N_18348,N_18629);
nor UO_216 (O_216,N_19049,N_19162);
nand UO_217 (O_217,N_19156,N_19991);
nand UO_218 (O_218,N_18617,N_19317);
or UO_219 (O_219,N_19668,N_19097);
and UO_220 (O_220,N_18310,N_19087);
and UO_221 (O_221,N_19019,N_18507);
and UO_222 (O_222,N_19500,N_19469);
xor UO_223 (O_223,N_18565,N_18606);
xnor UO_224 (O_224,N_19210,N_18276);
or UO_225 (O_225,N_18961,N_18754);
and UO_226 (O_226,N_18334,N_19546);
or UO_227 (O_227,N_18340,N_18793);
nand UO_228 (O_228,N_18846,N_18051);
nor UO_229 (O_229,N_18381,N_19798);
xnor UO_230 (O_230,N_19092,N_18319);
xor UO_231 (O_231,N_19610,N_18129);
xor UO_232 (O_232,N_19200,N_18149);
xor UO_233 (O_233,N_19259,N_19523);
nor UO_234 (O_234,N_19310,N_19290);
xnor UO_235 (O_235,N_19249,N_18359);
nand UO_236 (O_236,N_18506,N_18342);
and UO_237 (O_237,N_18870,N_19510);
and UO_238 (O_238,N_18108,N_19877);
or UO_239 (O_239,N_18308,N_19036);
and UO_240 (O_240,N_19191,N_19960);
and UO_241 (O_241,N_18345,N_18973);
and UO_242 (O_242,N_18862,N_19648);
or UO_243 (O_243,N_19756,N_19549);
nand UO_244 (O_244,N_18514,N_18217);
nand UO_245 (O_245,N_18722,N_18269);
or UO_246 (O_246,N_18527,N_19451);
nor UO_247 (O_247,N_18866,N_18443);
and UO_248 (O_248,N_18445,N_19944);
or UO_249 (O_249,N_19151,N_19214);
nand UO_250 (O_250,N_18396,N_18855);
nand UO_251 (O_251,N_18424,N_19319);
and UO_252 (O_252,N_18243,N_19121);
or UO_253 (O_253,N_19269,N_18323);
or UO_254 (O_254,N_19858,N_18932);
or UO_255 (O_255,N_19006,N_18286);
or UO_256 (O_256,N_18373,N_19720);
and UO_257 (O_257,N_18637,N_18887);
nor UO_258 (O_258,N_18499,N_18203);
and UO_259 (O_259,N_19433,N_18195);
nand UO_260 (O_260,N_18789,N_19489);
xnor UO_261 (O_261,N_18520,N_19029);
nor UO_262 (O_262,N_18420,N_19880);
or UO_263 (O_263,N_18616,N_18374);
and UO_264 (O_264,N_18403,N_19382);
nor UO_265 (O_265,N_19419,N_19884);
and UO_266 (O_266,N_19213,N_19379);
nor UO_267 (O_267,N_18360,N_18791);
or UO_268 (O_268,N_18245,N_18723);
and UO_269 (O_269,N_19238,N_18850);
nand UO_270 (O_270,N_19209,N_19050);
xor UO_271 (O_271,N_18552,N_19746);
nand UO_272 (O_272,N_19707,N_18498);
nor UO_273 (O_273,N_18131,N_18252);
nor UO_274 (O_274,N_19384,N_19110);
nand UO_275 (O_275,N_18819,N_19551);
nand UO_276 (O_276,N_18213,N_18784);
and UO_277 (O_277,N_19106,N_18247);
or UO_278 (O_278,N_18983,N_18098);
nor UO_279 (O_279,N_18738,N_19630);
or UO_280 (O_280,N_19373,N_19699);
and UO_281 (O_281,N_19573,N_18201);
or UO_282 (O_282,N_19817,N_18193);
xor UO_283 (O_283,N_18982,N_18154);
nor UO_284 (O_284,N_19839,N_18620);
and UO_285 (O_285,N_19946,N_18962);
or UO_286 (O_286,N_18758,N_19341);
nor UO_287 (O_287,N_19843,N_19008);
or UO_288 (O_288,N_18086,N_19847);
nand UO_289 (O_289,N_19444,N_18809);
nor UO_290 (O_290,N_19023,N_19354);
xor UO_291 (O_291,N_18103,N_18196);
or UO_292 (O_292,N_19088,N_18989);
nand UO_293 (O_293,N_18400,N_18429);
xor UO_294 (O_294,N_19108,N_18740);
nor UO_295 (O_295,N_18221,N_19056);
nand UO_296 (O_296,N_19605,N_19004);
and UO_297 (O_297,N_19690,N_19506);
or UO_298 (O_298,N_19637,N_19519);
and UO_299 (O_299,N_19959,N_19073);
nor UO_300 (O_300,N_19347,N_18110);
and UO_301 (O_301,N_19472,N_19696);
or UO_302 (O_302,N_18643,N_18661);
nor UO_303 (O_303,N_19807,N_18890);
or UO_304 (O_304,N_19795,N_19383);
and UO_305 (O_305,N_18080,N_19525);
nor UO_306 (O_306,N_19550,N_18454);
nand UO_307 (O_307,N_19410,N_18275);
nand UO_308 (O_308,N_19693,N_18083);
xor UO_309 (O_309,N_18684,N_19275);
or UO_310 (O_310,N_19454,N_19201);
or UO_311 (O_311,N_19217,N_18208);
xnor UO_312 (O_312,N_18769,N_19233);
nand UO_313 (O_313,N_19475,N_19571);
or UO_314 (O_314,N_18857,N_18230);
and UO_315 (O_315,N_19987,N_18004);
or UO_316 (O_316,N_19147,N_18447);
or UO_317 (O_317,N_18696,N_18667);
nor UO_318 (O_318,N_18440,N_19465);
nand UO_319 (O_319,N_18922,N_18134);
nor UO_320 (O_320,N_18885,N_18631);
or UO_321 (O_321,N_19661,N_19067);
nand UO_322 (O_322,N_19464,N_18027);
or UO_323 (O_323,N_18165,N_18037);
or UO_324 (O_324,N_18735,N_18607);
nand UO_325 (O_325,N_18829,N_19834);
nand UO_326 (O_326,N_19803,N_18448);
nand UO_327 (O_327,N_18831,N_19418);
nor UO_328 (O_328,N_19915,N_18898);
nor UO_329 (O_329,N_18411,N_18232);
and UO_330 (O_330,N_19044,N_19140);
nor UO_331 (O_331,N_19846,N_18879);
nor UO_332 (O_332,N_19381,N_18881);
nand UO_333 (O_333,N_18706,N_19576);
nand UO_334 (O_334,N_18057,N_19906);
and UO_335 (O_335,N_19658,N_19537);
nand UO_336 (O_336,N_19057,N_19683);
nor UO_337 (O_337,N_19485,N_19923);
or UO_338 (O_338,N_18864,N_18528);
nand UO_339 (O_339,N_18756,N_19709);
nor UO_340 (O_340,N_19671,N_19326);
and UO_341 (O_341,N_18996,N_19965);
and UO_342 (O_342,N_18550,N_19359);
or UO_343 (O_343,N_18413,N_19426);
nand UO_344 (O_344,N_18681,N_18877);
and UO_345 (O_345,N_18930,N_19046);
xnor UO_346 (O_346,N_19255,N_19813);
or UO_347 (O_347,N_19242,N_18474);
nor UO_348 (O_348,N_18670,N_18945);
xnor UO_349 (O_349,N_18273,N_18808);
nor UO_350 (O_350,N_18480,N_18473);
or UO_351 (O_351,N_18102,N_18785);
and UO_352 (O_352,N_18226,N_18582);
nand UO_353 (O_353,N_19903,N_19887);
and UO_354 (O_354,N_19873,N_18035);
nand UO_355 (O_355,N_19091,N_18488);
nand UO_356 (O_356,N_18044,N_18303);
nor UO_357 (O_357,N_18763,N_18284);
and UO_358 (O_358,N_19508,N_19390);
nand UO_359 (O_359,N_19833,N_19596);
xnor UO_360 (O_360,N_18282,N_19541);
nor UO_361 (O_361,N_19047,N_18251);
nor UO_362 (O_362,N_18346,N_18888);
or UO_363 (O_363,N_18006,N_18295);
and UO_364 (O_364,N_19331,N_19262);
xnor UO_365 (O_365,N_19995,N_19528);
and UO_366 (O_366,N_19122,N_19391);
or UO_367 (O_367,N_18790,N_19380);
nor UO_368 (O_368,N_19494,N_19408);
or UO_369 (O_369,N_18114,N_19231);
nand UO_370 (O_370,N_18314,N_18548);
nand UO_371 (O_371,N_18976,N_18814);
nor UO_372 (O_372,N_18683,N_18625);
nand UO_373 (O_373,N_19514,N_19521);
nor UO_374 (O_374,N_19731,N_19778);
nor UO_375 (O_375,N_19311,N_19078);
and UO_376 (O_376,N_18495,N_18180);
nand UO_377 (O_377,N_18433,N_19697);
and UO_378 (O_378,N_19398,N_18701);
nor UO_379 (O_379,N_18917,N_18010);
or UO_380 (O_380,N_18604,N_19028);
and UO_381 (O_381,N_18394,N_19252);
or UO_382 (O_382,N_19585,N_19612);
or UO_383 (O_383,N_18101,N_18399);
nor UO_384 (O_384,N_19711,N_18390);
nand UO_385 (O_385,N_18622,N_19216);
or UO_386 (O_386,N_19917,N_19862);
nand UO_387 (O_387,N_19396,N_18998);
nor UO_388 (O_388,N_18337,N_19769);
nor UO_389 (O_389,N_18655,N_19783);
or UO_390 (O_390,N_19996,N_19285);
xor UO_391 (O_391,N_19660,N_18772);
xor UO_392 (O_392,N_18869,N_19721);
nand UO_393 (O_393,N_18353,N_18199);
nor UO_394 (O_394,N_18654,N_19461);
or UO_395 (O_395,N_18692,N_18709);
nor UO_396 (O_396,N_18076,N_18395);
and UO_397 (O_397,N_19352,N_19104);
nor UO_398 (O_398,N_19026,N_18122);
or UO_399 (O_399,N_19972,N_18456);
and UO_400 (O_400,N_18921,N_19134);
or UO_401 (O_401,N_18956,N_18918);
xnor UO_402 (O_402,N_19411,N_18013);
nor UO_403 (O_403,N_19780,N_19770);
xor UO_404 (O_404,N_19371,N_18106);
and UO_405 (O_405,N_19875,N_19812);
or UO_406 (O_406,N_19938,N_18800);
or UO_407 (O_407,N_19708,N_19749);
nand UO_408 (O_408,N_19436,N_18609);
nor UO_409 (O_409,N_18845,N_19758);
nor UO_410 (O_410,N_18504,N_18327);
nand UO_411 (O_411,N_19345,N_19728);
xnor UO_412 (O_412,N_19702,N_19791);
xnor UO_413 (O_413,N_18233,N_19814);
nor UO_414 (O_414,N_19298,N_19442);
xor UO_415 (O_415,N_19416,N_18062);
xnor UO_416 (O_416,N_19116,N_19664);
and UO_417 (O_417,N_18810,N_19609);
nor UO_418 (O_418,N_19822,N_18551);
nor UO_419 (O_419,N_18562,N_19734);
xnor UO_420 (O_420,N_19051,N_18806);
or UO_421 (O_421,N_19686,N_18393);
nor UO_422 (O_422,N_18355,N_18534);
nand UO_423 (O_423,N_18570,N_18302);
or UO_424 (O_424,N_19531,N_19052);
and UO_425 (O_425,N_18262,N_19999);
and UO_426 (O_426,N_19787,N_18608);
nor UO_427 (O_427,N_19695,N_19955);
xor UO_428 (O_428,N_19303,N_19590);
or UO_429 (O_429,N_19608,N_18339);
or UO_430 (O_430,N_19062,N_18049);
and UO_431 (O_431,N_18786,N_18407);
nand UO_432 (O_432,N_19815,N_18172);
nor UO_433 (O_433,N_18185,N_18174);
and UO_434 (O_434,N_18465,N_19840);
xnor UO_435 (O_435,N_19703,N_19481);
and UO_436 (O_436,N_19248,N_19175);
and UO_437 (O_437,N_19957,N_19512);
nor UO_438 (O_438,N_18119,N_19301);
xor UO_439 (O_439,N_19714,N_19722);
or UO_440 (O_440,N_19673,N_19115);
nor UO_441 (O_441,N_18058,N_18457);
xnor UO_442 (O_442,N_18941,N_18047);
or UO_443 (O_443,N_19071,N_19178);
xor UO_444 (O_444,N_19684,N_19968);
and UO_445 (O_445,N_18688,N_19725);
nor UO_446 (O_446,N_18529,N_18019);
and UO_447 (O_447,N_19001,N_18832);
or UO_448 (O_448,N_18659,N_18828);
xnor UO_449 (O_449,N_19223,N_19325);
nor UO_450 (O_450,N_19942,N_19745);
nand UO_451 (O_451,N_19321,N_18746);
nand UO_452 (O_452,N_19517,N_18849);
or UO_453 (O_453,N_18179,N_18739);
and UO_454 (O_454,N_19375,N_19544);
nand UO_455 (O_455,N_19237,N_18292);
and UO_456 (O_456,N_18818,N_18293);
and UO_457 (O_457,N_19187,N_18535);
or UO_458 (O_458,N_18011,N_19895);
xnor UO_459 (O_459,N_19888,N_18089);
or UO_460 (O_460,N_19893,N_19131);
or UO_461 (O_461,N_18486,N_18139);
and UO_462 (O_462,N_19841,N_19562);
and UO_463 (O_463,N_19438,N_19587);
and UO_464 (O_464,N_18468,N_18494);
nor UO_465 (O_465,N_19886,N_19367);
and UO_466 (O_466,N_19823,N_18594);
and UO_467 (O_467,N_18151,N_18087);
or UO_468 (O_468,N_18970,N_19323);
and UO_469 (O_469,N_18410,N_18904);
and UO_470 (O_470,N_18899,N_19113);
or UO_471 (O_471,N_18693,N_18031);
nor UO_472 (O_472,N_18194,N_19796);
or UO_473 (O_473,N_18966,N_19838);
nand UO_474 (O_474,N_18248,N_19491);
and UO_475 (O_475,N_18099,N_18383);
or UO_476 (O_476,N_18298,N_18244);
xnor UO_477 (O_477,N_19507,N_19577);
and UO_478 (O_478,N_18979,N_19918);
nor UO_479 (O_479,N_19377,N_18459);
and UO_480 (O_480,N_18324,N_19542);
or UO_481 (O_481,N_18691,N_18588);
xor UO_482 (O_482,N_18000,N_19705);
nor UO_483 (O_483,N_19297,N_19974);
nand UO_484 (O_484,N_18483,N_18615);
or UO_485 (O_485,N_18096,N_19284);
or UO_486 (O_486,N_18647,N_18576);
nand UO_487 (O_487,N_19143,N_19183);
nand UO_488 (O_488,N_19535,N_19984);
or UO_489 (O_489,N_19386,N_19327);
nor UO_490 (O_490,N_19261,N_19997);
nand UO_491 (O_491,N_19022,N_18544);
nand UO_492 (O_492,N_19013,N_19744);
nand UO_493 (O_493,N_19651,N_19058);
nor UO_494 (O_494,N_19868,N_19422);
nor UO_495 (O_495,N_18142,N_19250);
nand UO_496 (O_496,N_19760,N_18388);
xor UO_497 (O_497,N_18757,N_18205);
and UO_498 (O_498,N_18689,N_18542);
or UO_499 (O_499,N_19565,N_19266);
nand UO_500 (O_500,N_19785,N_19158);
nand UO_501 (O_501,N_19155,N_18007);
and UO_502 (O_502,N_18909,N_19045);
nor UO_503 (O_503,N_18240,N_19492);
or UO_504 (O_504,N_19633,N_18018);
nand UO_505 (O_505,N_19522,N_18665);
nor UO_506 (O_506,N_18491,N_19459);
and UO_507 (O_507,N_18056,N_19174);
nand UO_508 (O_508,N_19098,N_18913);
nor UO_509 (O_509,N_18451,N_18708);
nand UO_510 (O_510,N_19179,N_18919);
xnor UO_511 (O_511,N_18707,N_19401);
nor UO_512 (O_512,N_18225,N_18717);
and UO_513 (O_513,N_19189,N_18581);
or UO_514 (O_514,N_18012,N_18329);
and UO_515 (O_515,N_18741,N_19914);
nor UO_516 (O_516,N_19689,N_19059);
nand UO_517 (O_517,N_18380,N_18093);
nor UO_518 (O_518,N_19936,N_18636);
nor UO_519 (O_519,N_19043,N_18002);
or UO_520 (O_520,N_19322,N_19003);
nand UO_521 (O_521,N_19204,N_19082);
or UO_522 (O_522,N_19932,N_19225);
nor UO_523 (O_523,N_18838,N_18745);
nor UO_524 (O_524,N_19079,N_18985);
and UO_525 (O_525,N_18834,N_18254);
nand UO_526 (O_526,N_19339,N_19497);
and UO_527 (O_527,N_18228,N_19399);
or UO_528 (O_528,N_18736,N_19589);
or UO_529 (O_529,N_18508,N_19532);
or UO_530 (O_530,N_18781,N_18054);
and UO_531 (O_531,N_18782,N_18668);
and UO_532 (O_532,N_19515,N_19159);
and UO_533 (O_533,N_19315,N_19878);
nor UO_534 (O_534,N_19730,N_18751);
or UO_535 (O_535,N_18458,N_18125);
nor UO_536 (O_536,N_19584,N_18977);
or UO_537 (O_537,N_19961,N_18729);
nor UO_538 (O_538,N_19621,N_18287);
xnor UO_539 (O_539,N_18081,N_18924);
or UO_540 (O_540,N_18414,N_18299);
nor UO_541 (O_541,N_18034,N_19455);
nand UO_542 (O_542,N_18032,N_19900);
nand UO_543 (O_543,N_18699,N_18734);
or UO_544 (O_544,N_19164,N_18437);
nor UO_545 (O_545,N_18022,N_18090);
or UO_546 (O_546,N_19617,N_19356);
nand UO_547 (O_547,N_19048,N_19754);
nand UO_548 (O_548,N_19417,N_19619);
xnor UO_549 (O_549,N_19694,N_19207);
xnor UO_550 (O_550,N_19622,N_19579);
and UO_551 (O_551,N_18698,N_19374);
nor UO_552 (O_552,N_19615,N_18449);
nand UO_553 (O_553,N_18442,N_19672);
xnor UO_554 (O_554,N_18452,N_19344);
and UO_555 (O_555,N_18218,N_18572);
nand UO_556 (O_556,N_19568,N_18220);
nor UO_557 (O_557,N_18798,N_18104);
and UO_558 (O_558,N_19199,N_18992);
and UO_559 (O_559,N_18994,N_18767);
and UO_560 (O_560,N_19540,N_19929);
xnor UO_561 (O_561,N_19260,N_18538);
nor UO_562 (O_562,N_18580,N_18415);
and UO_563 (O_563,N_18072,N_18549);
or UO_564 (O_564,N_19185,N_19413);
nor UO_565 (O_565,N_19263,N_19144);
nor UO_566 (O_566,N_19267,N_18843);
nand UO_567 (O_567,N_19251,N_19737);
nand UO_568 (O_568,N_19952,N_18066);
nand UO_569 (O_569,N_19009,N_18714);
and UO_570 (O_570,N_19574,N_19524);
nor UO_571 (O_571,N_18300,N_19075);
and UO_572 (O_572,N_19083,N_18990);
and UO_573 (O_573,N_18943,N_18682);
and UO_574 (O_574,N_18001,N_19934);
and UO_575 (O_575,N_19751,N_18479);
or UO_576 (O_576,N_18150,N_19656);
and UO_577 (O_577,N_18765,N_18117);
nand UO_578 (O_578,N_19520,N_19948);
and UO_579 (O_579,N_18624,N_19716);
nand UO_580 (O_580,N_19467,N_18875);
and UO_581 (O_581,N_18343,N_19196);
xnor UO_582 (O_582,N_18336,N_19318);
xor UO_583 (O_583,N_19240,N_18761);
nand UO_584 (O_584,N_19828,N_18658);
or UO_585 (O_585,N_19956,N_19885);
and UO_586 (O_586,N_18906,N_19450);
nand UO_587 (O_587,N_18253,N_18657);
or UO_588 (O_588,N_18613,N_19825);
and UO_589 (O_589,N_18462,N_19228);
or UO_590 (O_590,N_18993,N_19793);
nand UO_591 (O_591,N_18082,N_18307);
or UO_592 (O_592,N_18559,N_18533);
nand UO_593 (O_593,N_18981,N_19244);
or UO_594 (O_594,N_18675,N_18884);
or UO_595 (O_595,N_18126,N_18585);
xnor UO_596 (O_596,N_18571,N_18705);
or UO_597 (O_597,N_18197,N_18236);
nand UO_598 (O_598,N_18130,N_18436);
nor UO_599 (O_599,N_19931,N_18161);
nor UO_600 (O_600,N_19851,N_19452);
nor UO_601 (O_601,N_19152,N_18816);
or UO_602 (O_602,N_18872,N_19370);
nand UO_603 (O_603,N_18530,N_18678);
xor UO_604 (O_604,N_18778,N_19674);
nor UO_605 (O_605,N_18235,N_18141);
nand UO_606 (O_606,N_18805,N_19863);
nand UO_607 (O_607,N_18752,N_19767);
nor UO_608 (O_608,N_19504,N_19017);
or UO_609 (O_609,N_19063,N_18742);
nor UO_610 (O_610,N_18406,N_19501);
nor UO_611 (O_611,N_19636,N_19021);
and UO_612 (O_612,N_19427,N_19211);
and UO_613 (O_613,N_18728,N_19692);
nand UO_614 (O_614,N_18522,N_19953);
or UO_615 (O_615,N_19066,N_18905);
nand UO_616 (O_616,N_19268,N_19443);
or UO_617 (O_617,N_19593,N_19792);
or UO_618 (O_618,N_19640,N_18851);
nor UO_619 (O_619,N_18241,N_19480);
nand UO_620 (O_620,N_19282,N_18423);
and UO_621 (O_621,N_19077,N_18646);
nor UO_622 (O_622,N_19053,N_18444);
nand UO_623 (O_623,N_19458,N_19483);
and UO_624 (O_624,N_19222,N_19012);
nor UO_625 (O_625,N_19844,N_19715);
or UO_626 (O_626,N_18871,N_19064);
nand UO_627 (O_627,N_18430,N_19800);
nor UO_628 (O_628,N_19768,N_19670);
nor UO_629 (O_629,N_18487,N_18939);
xnor UO_630 (O_630,N_19276,N_19139);
or UO_631 (O_631,N_18813,N_19487);
xnor UO_632 (O_632,N_18954,N_18485);
or UO_633 (O_633,N_18835,N_18425);
nand UO_634 (O_634,N_18158,N_19992);
nor UO_635 (O_635,N_18427,N_19206);
nor UO_636 (O_636,N_19126,N_18601);
and UO_637 (O_637,N_19643,N_18215);
and UO_638 (O_638,N_19871,N_18189);
and UO_639 (O_639,N_19074,N_19447);
or UO_640 (O_640,N_19314,N_19530);
nand UO_641 (O_641,N_18183,N_19889);
nand UO_642 (O_642,N_19752,N_18687);
or UO_643 (O_643,N_18663,N_19581);
or UO_644 (O_644,N_18160,N_18974);
and UO_645 (O_645,N_18953,N_18988);
or UO_646 (O_646,N_19109,N_19986);
and UO_647 (O_647,N_18817,N_18749);
nor UO_648 (O_648,N_19086,N_18472);
or UO_649 (O_649,N_18949,N_19372);
nand UO_650 (O_650,N_18801,N_18071);
xor UO_651 (O_651,N_19117,N_18025);
nand UO_652 (O_652,N_18042,N_19677);
nor UO_653 (O_653,N_18475,N_19173);
or UO_654 (O_654,N_19597,N_18382);
nand UO_655 (O_655,N_18063,N_19623);
or UO_656 (O_656,N_18109,N_18916);
and UO_657 (O_657,N_19253,N_18596);
nand UO_658 (O_658,N_19613,N_19698);
xor UO_659 (O_659,N_19516,N_19892);
nand UO_660 (O_660,N_18113,N_18766);
xnor UO_661 (O_661,N_19570,N_19667);
or UO_662 (O_662,N_19364,N_19533);
or UO_663 (O_663,N_19271,N_19602);
xor UO_664 (O_664,N_19090,N_19435);
and UO_665 (O_665,N_18587,N_18948);
and UO_666 (O_666,N_18288,N_19457);
and UO_667 (O_667,N_19747,N_19488);
nand UO_668 (O_668,N_19719,N_19978);
and UO_669 (O_669,N_18021,N_19790);
or UO_670 (O_670,N_18886,N_19848);
nor UO_671 (O_671,N_18123,N_19857);
or UO_672 (O_672,N_18626,N_18270);
nand UO_673 (O_673,N_19292,N_19197);
or UO_674 (O_674,N_19750,N_19741);
or UO_675 (O_675,N_18212,N_18589);
and UO_676 (O_676,N_19264,N_18531);
nor UO_677 (O_677,N_19376,N_19599);
xor UO_678 (O_678,N_19424,N_19797);
and UO_679 (O_679,N_19580,N_19280);
nor UO_680 (O_680,N_19898,N_18660);
or UO_681 (O_681,N_19980,N_18118);
or UO_682 (O_682,N_19998,N_18611);
nand UO_683 (O_683,N_18952,N_19766);
or UO_684 (O_684,N_18033,N_19229);
and UO_685 (O_685,N_18787,N_18088);
or UO_686 (O_686,N_19198,N_19166);
nand UO_687 (O_687,N_18176,N_18599);
nor UO_688 (O_688,N_19101,N_18972);
nand UO_689 (O_689,N_18744,N_18836);
and UO_690 (O_690,N_19700,N_19055);
nor UO_691 (O_691,N_19020,N_19042);
nor UO_692 (O_692,N_18695,N_19406);
xnor UO_693 (O_693,N_19805,N_19423);
nor UO_694 (O_694,N_19710,N_19804);
and UO_695 (O_695,N_19913,N_18536);
nand UO_696 (O_696,N_18876,N_18277);
nand UO_697 (O_697,N_19538,N_18274);
nand UO_698 (O_698,N_18365,N_18181);
xor UO_699 (O_699,N_18564,N_19332);
xnor UO_700 (O_700,N_18815,N_19784);
and UO_701 (O_701,N_19169,N_18912);
and UO_702 (O_702,N_19157,N_18376);
and UO_703 (O_703,N_18198,N_19335);
or UO_704 (O_704,N_19563,N_18648);
and UO_705 (O_705,N_19782,N_18112);
and UO_706 (O_706,N_19355,N_19753);
and UO_707 (O_707,N_19462,N_19072);
nand UO_708 (O_708,N_19552,N_19736);
or UO_709 (O_709,N_18853,N_19471);
or UO_710 (O_710,N_19405,N_18431);
and UO_711 (O_711,N_18356,N_19360);
nand UO_712 (O_712,N_18140,N_19439);
xor UO_713 (O_713,N_18155,N_19896);
and UO_714 (O_714,N_18516,N_19299);
nand UO_715 (O_715,N_19819,N_18903);
nand UO_716 (O_716,N_18467,N_19307);
or UO_717 (O_717,N_19642,N_19717);
or UO_718 (O_718,N_18897,N_19133);
nand UO_719 (O_719,N_18156,N_19543);
nor UO_720 (O_720,N_19061,N_18460);
and UO_721 (O_721,N_19912,N_18385);
xnor UO_722 (O_722,N_18361,N_18521);
and UO_723 (O_723,N_18847,N_18331);
or UO_724 (O_724,N_18937,N_18350);
or UO_725 (O_725,N_19969,N_18470);
nand UO_726 (O_726,N_18404,N_18016);
nand UO_727 (O_727,N_19291,N_19890);
nand UO_728 (O_728,N_18206,N_19337);
nand UO_729 (O_729,N_18639,N_18656);
nand UO_730 (O_730,N_18971,N_19007);
nand UO_731 (O_731,N_19415,N_18322);
nor UO_732 (O_732,N_19470,N_18175);
nor UO_733 (O_733,N_18779,N_19578);
nor UO_734 (O_734,N_18895,N_19553);
and UO_735 (O_735,N_18822,N_18291);
xor UO_736 (O_736,N_18045,N_18614);
and UO_737 (O_737,N_18889,N_18064);
or UO_738 (O_738,N_18055,N_18592);
nor UO_739 (O_739,N_19723,N_18259);
or UO_740 (O_740,N_19035,N_18926);
nor UO_741 (O_741,N_19294,N_19607);
nor UO_742 (O_742,N_19837,N_19821);
xor UO_743 (O_743,N_18105,N_19502);
or UO_744 (O_744,N_18191,N_18263);
and UO_745 (O_745,N_18928,N_18664);
and UO_746 (O_746,N_18271,N_18377);
and UO_747 (O_747,N_19330,N_18069);
or UO_748 (O_748,N_18865,N_19920);
or UO_749 (O_749,N_19849,N_18190);
xor UO_750 (O_750,N_19278,N_19947);
and UO_751 (O_751,N_18283,N_18727);
and UO_752 (O_752,N_18547,N_19180);
nor UO_753 (O_753,N_18309,N_19033);
or UO_754 (O_754,N_19093,N_18068);
nand UO_755 (O_755,N_19922,N_19296);
or UO_756 (O_756,N_18074,N_19894);
and UO_757 (O_757,N_19545,N_19440);
nor UO_758 (O_758,N_19628,N_19350);
nand UO_759 (O_759,N_19193,N_19933);
nand UO_760 (O_760,N_19289,N_19160);
and UO_761 (O_761,N_19635,N_19065);
nand UO_762 (O_762,N_19188,N_18837);
nor UO_763 (O_763,N_18830,N_19852);
or UO_764 (O_764,N_18358,N_18525);
nor UO_765 (O_765,N_18496,N_19136);
xor UO_766 (O_766,N_19572,N_19286);
or UO_767 (O_767,N_18178,N_18950);
nand UO_768 (O_768,N_18464,N_19832);
or UO_769 (O_769,N_18641,N_18523);
nor UO_770 (O_770,N_18725,N_19368);
nand UO_771 (O_771,N_19343,N_18398);
and UO_772 (O_772,N_19567,N_18084);
nand UO_773 (O_773,N_18434,N_18713);
nand UO_774 (O_774,N_18929,N_18621);
and UO_775 (O_775,N_19385,N_18280);
or UO_776 (O_776,N_18540,N_18674);
and UO_777 (O_777,N_18168,N_19774);
and UO_778 (O_778,N_18854,N_18600);
or UO_779 (O_779,N_19434,N_18017);
nor UO_780 (O_780,N_19145,N_19123);
nor UO_781 (O_781,N_18642,N_18132);
or UO_782 (O_782,N_19281,N_18040);
and UO_783 (O_783,N_18222,N_18366);
nand UO_784 (O_784,N_18999,N_18257);
and UO_785 (O_785,N_19070,N_18043);
and UO_786 (O_786,N_19120,N_19128);
xor UO_787 (O_787,N_18153,N_18794);
or UO_788 (O_788,N_19831,N_18046);
or UO_789 (O_789,N_18618,N_19586);
nand UO_790 (O_790,N_19669,N_19060);
and UO_791 (O_791,N_19466,N_19691);
and UO_792 (O_792,N_18649,N_19748);
or UO_793 (O_793,N_18712,N_19926);
or UO_794 (O_794,N_18100,N_19921);
or UO_795 (O_795,N_19937,N_19149);
nand UO_796 (O_796,N_18933,N_19221);
nor UO_797 (O_797,N_18627,N_19979);
xnor UO_798 (O_798,N_18900,N_19015);
or UO_799 (O_799,N_18489,N_18927);
and UO_800 (O_800,N_18711,N_18797);
or UO_801 (O_801,N_18995,N_18863);
or UO_802 (O_802,N_18519,N_18418);
xnor UO_803 (O_803,N_18882,N_18482);
nand UO_804 (O_804,N_18768,N_19859);
nor UO_805 (O_805,N_19349,N_18008);
nor UO_806 (O_806,N_18167,N_19102);
nor UO_807 (O_807,N_18095,N_18555);
and UO_808 (O_808,N_19089,N_19176);
nand UO_809 (O_809,N_19293,N_19743);
or UO_810 (O_810,N_18598,N_19786);
or UO_811 (O_811,N_19554,N_18686);
or UO_812 (O_812,N_18679,N_18078);
or UO_813 (O_813,N_19583,N_19084);
or UO_814 (O_814,N_19739,N_18171);
and UO_815 (O_815,N_18891,N_18453);
or UO_816 (O_816,N_19215,N_18073);
nor UO_817 (O_817,N_18249,N_19402);
and UO_818 (O_818,N_18481,N_19547);
and UO_819 (O_819,N_19618,N_18964);
and UO_820 (O_820,N_18557,N_19258);
or UO_821 (O_821,N_18718,N_18770);
and UO_822 (O_822,N_18680,N_18379);
nand UO_823 (O_823,N_19038,N_18861);
or UO_824 (O_824,N_19735,N_18651);
or UO_825 (O_825,N_19153,N_19431);
nor UO_826 (O_826,N_19039,N_18368);
nand UO_827 (O_827,N_19983,N_19882);
or UO_828 (O_828,N_19283,N_19794);
nand UO_829 (O_829,N_18301,N_19687);
nand UO_830 (O_830,N_18333,N_19982);
xor UO_831 (O_831,N_18892,N_19338);
and UO_832 (O_832,N_18563,N_18246);
nor UO_833 (O_833,N_19024,N_18517);
or UO_834 (O_834,N_19654,N_19369);
and UO_835 (O_835,N_19861,N_19236);
nand UO_836 (O_836,N_18880,N_18575);
and UO_837 (O_837,N_18364,N_19854);
and UO_838 (O_838,N_19484,N_18493);
and UO_839 (O_839,N_18085,N_18867);
nor UO_840 (O_840,N_19901,N_19002);
or UO_841 (O_841,N_18317,N_18242);
or UO_842 (O_842,N_18372,N_18094);
or UO_843 (O_843,N_18726,N_19808);
xnor UO_844 (O_844,N_18777,N_19638);
nand UO_845 (O_845,N_19726,N_19005);
or UO_846 (O_846,N_19561,N_19827);
nor UO_847 (O_847,N_19287,N_19154);
nor UO_848 (O_848,N_19068,N_19421);
and UO_849 (O_849,N_19351,N_19080);
nand UO_850 (O_850,N_19864,N_19096);
and UO_851 (O_851,N_18730,N_19976);
nor UO_852 (O_852,N_18842,N_19988);
nor UO_853 (O_853,N_19148,N_18029);
nand UO_854 (O_854,N_19835,N_19845);
or UO_855 (O_855,N_18357,N_19990);
or UO_856 (O_856,N_19234,N_19437);
nand UO_857 (O_857,N_18325,N_18574);
and UO_858 (O_858,N_18036,N_19473);
xnor UO_859 (O_859,N_19762,N_18320);
nand UO_860 (O_860,N_19270,N_19334);
nand UO_861 (O_861,N_18694,N_19468);
or UO_862 (O_862,N_18561,N_18238);
or UO_863 (O_863,N_18733,N_19575);
nand UO_864 (O_864,N_19950,N_19772);
nand UO_865 (O_865,N_19245,N_18041);
or UO_866 (O_866,N_19076,N_18967);
xor UO_867 (O_867,N_18568,N_19765);
and UO_868 (O_868,N_19600,N_18023);
nor UO_869 (O_869,N_18421,N_18239);
xor UO_870 (O_870,N_18584,N_18662);
nand UO_871 (O_871,N_18170,N_18147);
xnor UO_872 (O_872,N_18702,N_18354);
nand UO_873 (O_873,N_19729,N_18638);
nand UO_874 (O_874,N_19526,N_19230);
and UO_875 (O_875,N_18289,N_19558);
or UO_876 (O_876,N_19981,N_19184);
or UO_877 (O_877,N_18265,N_18219);
and UO_878 (O_878,N_18030,N_19967);
nor UO_879 (O_879,N_19951,N_18053);
nand UO_880 (O_880,N_19037,N_18207);
nor UO_881 (O_881,N_18432,N_18476);
and UO_882 (O_882,N_19620,N_18075);
and UO_883 (O_883,N_18164,N_19505);
and UO_884 (O_884,N_19474,N_19336);
nand UO_885 (O_885,N_18026,N_18883);
nor UO_886 (O_886,N_18776,N_19232);
nand UO_887 (O_887,N_19733,N_18120);
nand UO_888 (O_888,N_19764,N_19829);
and UO_889 (O_889,N_19168,N_19346);
nand UO_890 (O_890,N_18844,N_18229);
nand UO_891 (O_891,N_18958,N_18266);
and UO_892 (O_892,N_19498,N_18210);
and UO_893 (O_893,N_18732,N_18048);
nand UO_894 (O_894,N_19357,N_18214);
nor UO_895 (O_895,N_19802,N_18378);
and UO_896 (O_896,N_19557,N_18558);
nor UO_897 (O_897,N_19555,N_19014);
or UO_898 (O_898,N_19742,N_19205);
or UO_899 (O_899,N_19666,N_19219);
or UO_900 (O_900,N_19985,N_18124);
nor UO_901 (O_901,N_19776,N_19650);
nand UO_902 (O_902,N_19203,N_19163);
nand UO_903 (O_903,N_18107,N_19182);
nor UO_904 (O_904,N_19138,N_18923);
nand UO_905 (O_905,N_18653,N_18490);
or UO_906 (O_906,N_19559,N_18960);
or UO_907 (O_907,N_18501,N_19011);
and UO_908 (O_908,N_18441,N_18856);
and UO_909 (O_909,N_19403,N_19830);
nand UO_910 (O_910,N_18321,N_19150);
nor UO_911 (O_911,N_19107,N_19114);
and UO_912 (O_912,N_19850,N_19806);
nor UO_913 (O_913,N_18408,N_18792);
or UO_914 (O_914,N_18312,N_19688);
and UO_915 (O_915,N_18097,N_19316);
and UO_916 (O_916,N_18092,N_19503);
and UO_917 (O_917,N_18351,N_19220);
nand UO_918 (O_918,N_18807,N_18386);
or UO_919 (O_919,N_19400,N_18783);
or UO_920 (O_920,N_19975,N_18187);
nor UO_921 (O_921,N_18539,N_19446);
nor UO_922 (O_922,N_18143,N_19192);
nand UO_923 (O_923,N_19247,N_18463);
nand UO_924 (O_924,N_19306,N_18541);
nor UO_925 (O_925,N_19701,N_19429);
nor UO_926 (O_926,N_18328,N_18079);
or UO_927 (O_927,N_19493,N_18362);
nand UO_928 (O_928,N_19740,N_18272);
xor UO_929 (O_929,N_18650,N_19226);
and UO_930 (O_930,N_18417,N_19556);
nor UO_931 (O_931,N_18446,N_18121);
or UO_932 (O_932,N_19606,N_19309);
nor UO_933 (O_933,N_18748,N_19820);
or UO_934 (O_934,N_18039,N_19254);
or UO_935 (O_935,N_18747,N_18290);
and UO_936 (O_936,N_19653,N_19235);
and UO_937 (O_937,N_18231,N_18375);
nand UO_938 (O_938,N_19548,N_18148);
xor UO_939 (O_939,N_18279,N_18512);
and UO_940 (O_940,N_19663,N_18332);
and UO_941 (O_941,N_19388,N_18392);
nor UO_942 (O_942,N_19977,N_18278);
nand UO_943 (O_943,N_18685,N_18669);
xnor UO_944 (O_944,N_18940,N_19777);
and UO_945 (O_945,N_19891,N_18703);
nand UO_946 (O_946,N_19943,N_18188);
xor UO_947 (O_947,N_18264,N_18234);
and UO_948 (O_948,N_18091,N_19482);
or UO_949 (O_949,N_18944,N_19495);
xor UO_950 (O_950,N_19865,N_19681);
nand UO_951 (O_951,N_19902,N_18177);
or UO_952 (O_952,N_18526,N_19392);
nor UO_953 (O_953,N_19511,N_18182);
nand UO_954 (O_954,N_18469,N_19582);
or UO_955 (O_955,N_19186,N_18978);
and UO_956 (O_956,N_19909,N_19407);
xor UO_957 (O_957,N_18166,N_18764);
nor UO_958 (O_958,N_18959,N_19387);
and UO_959 (O_959,N_18947,N_19170);
xor UO_960 (O_960,N_18894,N_19239);
nand UO_961 (O_961,N_19142,N_18313);
nor UO_962 (O_962,N_18511,N_18852);
nor UO_963 (O_963,N_19566,N_18859);
and UO_964 (O_964,N_18162,N_19208);
nor UO_965 (O_965,N_19460,N_18848);
nor UO_966 (O_966,N_19818,N_18227);
nand UO_967 (O_967,N_18907,N_18500);
nand UO_968 (O_968,N_18003,N_19872);
and UO_969 (O_969,N_19836,N_19365);
or UO_970 (O_970,N_18052,N_19348);
nand UO_971 (O_971,N_19842,N_19414);
and UO_972 (O_972,N_19675,N_19916);
and UO_973 (O_973,N_19641,N_18633);
nand UO_974 (O_974,N_19030,N_19362);
and UO_975 (O_975,N_18825,N_19161);
xor UO_976 (O_976,N_18478,N_19941);
nor UO_977 (O_977,N_18936,N_18946);
or UO_978 (O_978,N_19676,N_19172);
and UO_979 (O_979,N_19257,N_19925);
or UO_980 (O_980,N_18412,N_19855);
nor UO_981 (O_981,N_18438,N_19738);
and UO_982 (O_982,N_18710,N_18893);
nand UO_983 (O_983,N_18812,N_19194);
nor UO_984 (O_984,N_18593,N_18715);
and UO_985 (O_985,N_18545,N_18908);
and UO_986 (O_986,N_18028,N_18532);
xnor UO_987 (O_987,N_19634,N_19103);
or UO_988 (O_988,N_18991,N_18347);
nand UO_989 (O_989,N_18963,N_18677);
or UO_990 (O_990,N_19389,N_18560);
nor UO_991 (O_991,N_18902,N_19779);
or UO_992 (O_992,N_19137,N_18755);
or UO_993 (O_993,N_19625,N_19616);
or UO_994 (O_994,N_18567,N_18915);
nor UO_995 (O_995,N_19099,N_18719);
or UO_996 (O_996,N_19949,N_18330);
nand UO_997 (O_997,N_19308,N_18405);
nor UO_998 (O_998,N_18774,N_19853);
or UO_999 (O_999,N_19085,N_18788);
or UO_1000 (O_1000,N_19802,N_18685);
nand UO_1001 (O_1001,N_19822,N_18729);
nand UO_1002 (O_1002,N_19832,N_19257);
and UO_1003 (O_1003,N_19224,N_19782);
nor UO_1004 (O_1004,N_19248,N_19649);
nand UO_1005 (O_1005,N_19551,N_19004);
nand UO_1006 (O_1006,N_19956,N_18498);
and UO_1007 (O_1007,N_19544,N_19969);
and UO_1008 (O_1008,N_18107,N_19272);
xor UO_1009 (O_1009,N_19980,N_19549);
nand UO_1010 (O_1010,N_19267,N_19243);
and UO_1011 (O_1011,N_18539,N_19124);
nor UO_1012 (O_1012,N_18149,N_18450);
xor UO_1013 (O_1013,N_19117,N_19403);
xnor UO_1014 (O_1014,N_19401,N_18787);
nor UO_1015 (O_1015,N_19212,N_19563);
xor UO_1016 (O_1016,N_19906,N_18746);
nand UO_1017 (O_1017,N_18101,N_19863);
nand UO_1018 (O_1018,N_19675,N_19030);
and UO_1019 (O_1019,N_18778,N_19931);
nor UO_1020 (O_1020,N_18296,N_19159);
nand UO_1021 (O_1021,N_18542,N_18445);
nor UO_1022 (O_1022,N_18512,N_18320);
or UO_1023 (O_1023,N_19618,N_19976);
nor UO_1024 (O_1024,N_19333,N_18711);
nand UO_1025 (O_1025,N_18435,N_19975);
nor UO_1026 (O_1026,N_18260,N_19799);
nor UO_1027 (O_1027,N_18031,N_18808);
nand UO_1028 (O_1028,N_18400,N_19308);
nor UO_1029 (O_1029,N_18518,N_19508);
and UO_1030 (O_1030,N_18352,N_19100);
or UO_1031 (O_1031,N_18588,N_19177);
nand UO_1032 (O_1032,N_18116,N_18590);
nor UO_1033 (O_1033,N_19983,N_18553);
nor UO_1034 (O_1034,N_18623,N_19076);
xor UO_1035 (O_1035,N_19729,N_19647);
nor UO_1036 (O_1036,N_19704,N_18531);
nor UO_1037 (O_1037,N_18982,N_19534);
nor UO_1038 (O_1038,N_18108,N_19435);
nor UO_1039 (O_1039,N_18961,N_19388);
or UO_1040 (O_1040,N_19525,N_19888);
or UO_1041 (O_1041,N_18623,N_18605);
xor UO_1042 (O_1042,N_19122,N_19317);
or UO_1043 (O_1043,N_18037,N_19201);
and UO_1044 (O_1044,N_19125,N_19139);
nor UO_1045 (O_1045,N_18315,N_19518);
nand UO_1046 (O_1046,N_18325,N_18535);
nand UO_1047 (O_1047,N_19398,N_19131);
and UO_1048 (O_1048,N_18573,N_19919);
xnor UO_1049 (O_1049,N_18218,N_18396);
nand UO_1050 (O_1050,N_18471,N_18327);
nor UO_1051 (O_1051,N_18048,N_18874);
xnor UO_1052 (O_1052,N_19571,N_18366);
nand UO_1053 (O_1053,N_18839,N_18587);
and UO_1054 (O_1054,N_18323,N_18428);
nand UO_1055 (O_1055,N_18273,N_19746);
nor UO_1056 (O_1056,N_18798,N_18803);
or UO_1057 (O_1057,N_18486,N_19817);
xor UO_1058 (O_1058,N_19678,N_19302);
nand UO_1059 (O_1059,N_19275,N_19454);
nor UO_1060 (O_1060,N_19681,N_18698);
nand UO_1061 (O_1061,N_19878,N_19701);
or UO_1062 (O_1062,N_19796,N_19291);
xor UO_1063 (O_1063,N_18556,N_19252);
nor UO_1064 (O_1064,N_18638,N_18949);
nand UO_1065 (O_1065,N_18557,N_18858);
nand UO_1066 (O_1066,N_18973,N_18589);
xor UO_1067 (O_1067,N_18860,N_19350);
nor UO_1068 (O_1068,N_19077,N_19629);
nor UO_1069 (O_1069,N_19409,N_18130);
nor UO_1070 (O_1070,N_19896,N_18764);
and UO_1071 (O_1071,N_18740,N_18309);
or UO_1072 (O_1072,N_19227,N_18142);
nand UO_1073 (O_1073,N_18368,N_19584);
nand UO_1074 (O_1074,N_18259,N_18190);
nor UO_1075 (O_1075,N_19150,N_19142);
xor UO_1076 (O_1076,N_19362,N_18156);
nand UO_1077 (O_1077,N_18489,N_19411);
nand UO_1078 (O_1078,N_19577,N_19527);
nand UO_1079 (O_1079,N_19540,N_19040);
and UO_1080 (O_1080,N_18514,N_19741);
and UO_1081 (O_1081,N_18140,N_19034);
nor UO_1082 (O_1082,N_19646,N_19372);
nor UO_1083 (O_1083,N_18036,N_18984);
nor UO_1084 (O_1084,N_18289,N_19598);
or UO_1085 (O_1085,N_18935,N_19636);
and UO_1086 (O_1086,N_19945,N_19994);
nand UO_1087 (O_1087,N_18810,N_19121);
or UO_1088 (O_1088,N_19954,N_18115);
or UO_1089 (O_1089,N_19824,N_19913);
and UO_1090 (O_1090,N_19316,N_19500);
nor UO_1091 (O_1091,N_18276,N_19624);
nand UO_1092 (O_1092,N_19508,N_19064);
nor UO_1093 (O_1093,N_19453,N_18070);
or UO_1094 (O_1094,N_18547,N_18227);
nor UO_1095 (O_1095,N_18903,N_19431);
or UO_1096 (O_1096,N_19405,N_19901);
nor UO_1097 (O_1097,N_19964,N_19291);
nor UO_1098 (O_1098,N_19615,N_19432);
nor UO_1099 (O_1099,N_18263,N_18380);
or UO_1100 (O_1100,N_18991,N_19460);
nor UO_1101 (O_1101,N_18298,N_19699);
or UO_1102 (O_1102,N_18512,N_18945);
nand UO_1103 (O_1103,N_19039,N_19464);
or UO_1104 (O_1104,N_18186,N_18909);
or UO_1105 (O_1105,N_19096,N_19263);
and UO_1106 (O_1106,N_18840,N_19347);
nand UO_1107 (O_1107,N_19165,N_19164);
or UO_1108 (O_1108,N_19239,N_18249);
and UO_1109 (O_1109,N_19052,N_19241);
and UO_1110 (O_1110,N_18004,N_19889);
nor UO_1111 (O_1111,N_19485,N_18698);
nor UO_1112 (O_1112,N_18288,N_19951);
and UO_1113 (O_1113,N_19649,N_19358);
nor UO_1114 (O_1114,N_18778,N_19419);
or UO_1115 (O_1115,N_19754,N_18538);
or UO_1116 (O_1116,N_19581,N_18186);
xor UO_1117 (O_1117,N_18050,N_18222);
nor UO_1118 (O_1118,N_19751,N_18877);
nor UO_1119 (O_1119,N_19921,N_19497);
and UO_1120 (O_1120,N_18930,N_18191);
or UO_1121 (O_1121,N_19254,N_18632);
and UO_1122 (O_1122,N_18358,N_19366);
or UO_1123 (O_1123,N_18988,N_19879);
or UO_1124 (O_1124,N_19900,N_19521);
or UO_1125 (O_1125,N_18094,N_18656);
xor UO_1126 (O_1126,N_18430,N_18017);
or UO_1127 (O_1127,N_19161,N_19194);
nor UO_1128 (O_1128,N_19942,N_18641);
nand UO_1129 (O_1129,N_19090,N_18418);
xor UO_1130 (O_1130,N_19704,N_19694);
nand UO_1131 (O_1131,N_18835,N_18936);
nor UO_1132 (O_1132,N_19571,N_18767);
or UO_1133 (O_1133,N_18200,N_18994);
and UO_1134 (O_1134,N_19444,N_19935);
nor UO_1135 (O_1135,N_18798,N_19826);
nor UO_1136 (O_1136,N_19894,N_18413);
nor UO_1137 (O_1137,N_18616,N_18014);
nor UO_1138 (O_1138,N_18091,N_19160);
and UO_1139 (O_1139,N_19894,N_18914);
or UO_1140 (O_1140,N_18575,N_18289);
and UO_1141 (O_1141,N_18416,N_19711);
nand UO_1142 (O_1142,N_19844,N_18537);
and UO_1143 (O_1143,N_19099,N_19061);
and UO_1144 (O_1144,N_18975,N_18485);
nor UO_1145 (O_1145,N_18710,N_19826);
nor UO_1146 (O_1146,N_19245,N_19823);
nand UO_1147 (O_1147,N_18354,N_19696);
or UO_1148 (O_1148,N_19019,N_18795);
nand UO_1149 (O_1149,N_18544,N_18413);
nor UO_1150 (O_1150,N_19041,N_19480);
nand UO_1151 (O_1151,N_18271,N_18403);
nand UO_1152 (O_1152,N_19318,N_19394);
xor UO_1153 (O_1153,N_19594,N_18017);
nor UO_1154 (O_1154,N_18982,N_18258);
nor UO_1155 (O_1155,N_19160,N_18383);
or UO_1156 (O_1156,N_18458,N_19282);
nand UO_1157 (O_1157,N_18071,N_18609);
and UO_1158 (O_1158,N_19280,N_18533);
nor UO_1159 (O_1159,N_18548,N_18200);
or UO_1160 (O_1160,N_19030,N_19165);
and UO_1161 (O_1161,N_18006,N_19865);
nand UO_1162 (O_1162,N_19553,N_19265);
and UO_1163 (O_1163,N_18729,N_19287);
or UO_1164 (O_1164,N_19665,N_19777);
and UO_1165 (O_1165,N_18733,N_19293);
nand UO_1166 (O_1166,N_19830,N_19867);
nand UO_1167 (O_1167,N_19301,N_18155);
or UO_1168 (O_1168,N_19572,N_19115);
or UO_1169 (O_1169,N_19513,N_18205);
nor UO_1170 (O_1170,N_18614,N_19851);
nand UO_1171 (O_1171,N_19638,N_19947);
nor UO_1172 (O_1172,N_19738,N_19342);
nand UO_1173 (O_1173,N_19596,N_19614);
xor UO_1174 (O_1174,N_19183,N_19741);
or UO_1175 (O_1175,N_19184,N_18633);
nand UO_1176 (O_1176,N_18674,N_19033);
and UO_1177 (O_1177,N_19490,N_18919);
nand UO_1178 (O_1178,N_18498,N_19539);
nand UO_1179 (O_1179,N_18376,N_19981);
nor UO_1180 (O_1180,N_19773,N_18349);
or UO_1181 (O_1181,N_19446,N_19031);
or UO_1182 (O_1182,N_18377,N_19476);
or UO_1183 (O_1183,N_19574,N_19916);
or UO_1184 (O_1184,N_19383,N_19703);
or UO_1185 (O_1185,N_18794,N_18467);
or UO_1186 (O_1186,N_18684,N_19495);
nor UO_1187 (O_1187,N_19462,N_18224);
and UO_1188 (O_1188,N_19124,N_18444);
nor UO_1189 (O_1189,N_18028,N_18240);
and UO_1190 (O_1190,N_18019,N_18630);
or UO_1191 (O_1191,N_18779,N_18512);
nand UO_1192 (O_1192,N_18770,N_18160);
xor UO_1193 (O_1193,N_19447,N_19465);
and UO_1194 (O_1194,N_18206,N_19623);
nor UO_1195 (O_1195,N_18746,N_18819);
xor UO_1196 (O_1196,N_19689,N_19088);
xor UO_1197 (O_1197,N_18149,N_18741);
or UO_1198 (O_1198,N_18738,N_18193);
and UO_1199 (O_1199,N_18189,N_18692);
and UO_1200 (O_1200,N_18306,N_19699);
or UO_1201 (O_1201,N_19168,N_18135);
xnor UO_1202 (O_1202,N_18735,N_19185);
and UO_1203 (O_1203,N_18700,N_19735);
or UO_1204 (O_1204,N_19287,N_18454);
and UO_1205 (O_1205,N_18860,N_19156);
xor UO_1206 (O_1206,N_19233,N_19746);
and UO_1207 (O_1207,N_19909,N_18627);
nand UO_1208 (O_1208,N_19058,N_18997);
nor UO_1209 (O_1209,N_18795,N_19788);
nor UO_1210 (O_1210,N_18426,N_19335);
nor UO_1211 (O_1211,N_18536,N_18175);
nand UO_1212 (O_1212,N_18640,N_18562);
nand UO_1213 (O_1213,N_18348,N_18099);
xor UO_1214 (O_1214,N_19281,N_18735);
nand UO_1215 (O_1215,N_19635,N_19206);
and UO_1216 (O_1216,N_18831,N_18644);
or UO_1217 (O_1217,N_18698,N_18578);
nand UO_1218 (O_1218,N_19467,N_19832);
or UO_1219 (O_1219,N_18396,N_19136);
nor UO_1220 (O_1220,N_18795,N_18728);
nor UO_1221 (O_1221,N_19720,N_19882);
nor UO_1222 (O_1222,N_19930,N_19077);
nand UO_1223 (O_1223,N_19749,N_18056);
and UO_1224 (O_1224,N_18106,N_18858);
or UO_1225 (O_1225,N_19814,N_18134);
or UO_1226 (O_1226,N_19210,N_18188);
or UO_1227 (O_1227,N_19911,N_18799);
or UO_1228 (O_1228,N_18513,N_18668);
nand UO_1229 (O_1229,N_18206,N_18988);
nand UO_1230 (O_1230,N_18386,N_19440);
or UO_1231 (O_1231,N_19617,N_19173);
and UO_1232 (O_1232,N_18973,N_19334);
nor UO_1233 (O_1233,N_18822,N_18850);
nand UO_1234 (O_1234,N_19134,N_18941);
or UO_1235 (O_1235,N_19910,N_18085);
or UO_1236 (O_1236,N_19592,N_19803);
and UO_1237 (O_1237,N_19237,N_18735);
xnor UO_1238 (O_1238,N_18984,N_19406);
nor UO_1239 (O_1239,N_18161,N_18537);
nor UO_1240 (O_1240,N_18520,N_18151);
and UO_1241 (O_1241,N_18520,N_18110);
and UO_1242 (O_1242,N_18056,N_18493);
or UO_1243 (O_1243,N_19145,N_18004);
or UO_1244 (O_1244,N_18690,N_19244);
nand UO_1245 (O_1245,N_19983,N_18342);
or UO_1246 (O_1246,N_19532,N_19395);
or UO_1247 (O_1247,N_19340,N_18021);
nor UO_1248 (O_1248,N_18556,N_19124);
nand UO_1249 (O_1249,N_18275,N_18366);
nand UO_1250 (O_1250,N_19737,N_18552);
nor UO_1251 (O_1251,N_19955,N_18749);
nand UO_1252 (O_1252,N_19786,N_18160);
xor UO_1253 (O_1253,N_19859,N_19593);
or UO_1254 (O_1254,N_19740,N_18675);
xnor UO_1255 (O_1255,N_18942,N_19347);
nand UO_1256 (O_1256,N_18871,N_19923);
or UO_1257 (O_1257,N_19008,N_18587);
xor UO_1258 (O_1258,N_19040,N_18505);
and UO_1259 (O_1259,N_19840,N_19066);
or UO_1260 (O_1260,N_18156,N_19743);
and UO_1261 (O_1261,N_18014,N_18502);
or UO_1262 (O_1262,N_18798,N_18776);
nand UO_1263 (O_1263,N_19787,N_18600);
nor UO_1264 (O_1264,N_19319,N_19127);
xnor UO_1265 (O_1265,N_19914,N_19376);
and UO_1266 (O_1266,N_18008,N_18259);
or UO_1267 (O_1267,N_19110,N_18758);
and UO_1268 (O_1268,N_18740,N_18395);
or UO_1269 (O_1269,N_19593,N_18608);
nand UO_1270 (O_1270,N_19901,N_18530);
or UO_1271 (O_1271,N_18736,N_19148);
nand UO_1272 (O_1272,N_19116,N_18099);
or UO_1273 (O_1273,N_18976,N_19210);
nor UO_1274 (O_1274,N_19823,N_18504);
nor UO_1275 (O_1275,N_18588,N_18842);
nor UO_1276 (O_1276,N_19517,N_19732);
nand UO_1277 (O_1277,N_18776,N_19242);
xnor UO_1278 (O_1278,N_18410,N_19729);
nand UO_1279 (O_1279,N_19425,N_18904);
and UO_1280 (O_1280,N_18482,N_19348);
nand UO_1281 (O_1281,N_18301,N_18421);
or UO_1282 (O_1282,N_19484,N_18380);
nor UO_1283 (O_1283,N_19326,N_19563);
nor UO_1284 (O_1284,N_18978,N_18105);
nor UO_1285 (O_1285,N_19273,N_18093);
and UO_1286 (O_1286,N_19840,N_18448);
xor UO_1287 (O_1287,N_18147,N_19504);
or UO_1288 (O_1288,N_18283,N_18951);
and UO_1289 (O_1289,N_19412,N_18154);
nor UO_1290 (O_1290,N_19068,N_19452);
or UO_1291 (O_1291,N_18454,N_19294);
and UO_1292 (O_1292,N_18964,N_18056);
and UO_1293 (O_1293,N_19589,N_19690);
xor UO_1294 (O_1294,N_19716,N_19732);
nand UO_1295 (O_1295,N_19107,N_19895);
and UO_1296 (O_1296,N_19878,N_18222);
nor UO_1297 (O_1297,N_19722,N_19030);
nand UO_1298 (O_1298,N_18630,N_19220);
nand UO_1299 (O_1299,N_18686,N_18495);
or UO_1300 (O_1300,N_18301,N_18487);
and UO_1301 (O_1301,N_19757,N_19321);
nor UO_1302 (O_1302,N_18171,N_18897);
xnor UO_1303 (O_1303,N_18588,N_19798);
and UO_1304 (O_1304,N_18876,N_19824);
and UO_1305 (O_1305,N_19977,N_19406);
nor UO_1306 (O_1306,N_18154,N_19102);
or UO_1307 (O_1307,N_19807,N_19381);
and UO_1308 (O_1308,N_18370,N_18542);
or UO_1309 (O_1309,N_18438,N_19053);
and UO_1310 (O_1310,N_18931,N_18390);
or UO_1311 (O_1311,N_18827,N_18684);
xor UO_1312 (O_1312,N_18182,N_18564);
nand UO_1313 (O_1313,N_19210,N_19585);
nor UO_1314 (O_1314,N_18637,N_18448);
xnor UO_1315 (O_1315,N_18483,N_18604);
nand UO_1316 (O_1316,N_19478,N_19956);
nor UO_1317 (O_1317,N_18172,N_19018);
and UO_1318 (O_1318,N_19185,N_18366);
nand UO_1319 (O_1319,N_19177,N_19237);
and UO_1320 (O_1320,N_18846,N_18272);
or UO_1321 (O_1321,N_18310,N_18428);
and UO_1322 (O_1322,N_18930,N_19646);
or UO_1323 (O_1323,N_18321,N_18539);
and UO_1324 (O_1324,N_18428,N_18479);
and UO_1325 (O_1325,N_19885,N_19831);
nor UO_1326 (O_1326,N_18644,N_19851);
nand UO_1327 (O_1327,N_19767,N_18524);
xnor UO_1328 (O_1328,N_19427,N_19463);
or UO_1329 (O_1329,N_19539,N_19685);
nand UO_1330 (O_1330,N_19393,N_18332);
or UO_1331 (O_1331,N_18395,N_19270);
or UO_1332 (O_1332,N_18369,N_19919);
and UO_1333 (O_1333,N_19468,N_18611);
nor UO_1334 (O_1334,N_18800,N_19374);
and UO_1335 (O_1335,N_19621,N_19815);
xor UO_1336 (O_1336,N_18942,N_18876);
nor UO_1337 (O_1337,N_19295,N_19417);
and UO_1338 (O_1338,N_19689,N_18970);
nand UO_1339 (O_1339,N_18975,N_19988);
xnor UO_1340 (O_1340,N_19950,N_19920);
nor UO_1341 (O_1341,N_18167,N_18471);
nand UO_1342 (O_1342,N_19021,N_18530);
or UO_1343 (O_1343,N_19210,N_19611);
nor UO_1344 (O_1344,N_19203,N_18908);
nor UO_1345 (O_1345,N_18187,N_19074);
and UO_1346 (O_1346,N_18643,N_18008);
or UO_1347 (O_1347,N_18927,N_19569);
and UO_1348 (O_1348,N_18922,N_19036);
nor UO_1349 (O_1349,N_18771,N_19138);
and UO_1350 (O_1350,N_19521,N_18345);
or UO_1351 (O_1351,N_18047,N_18697);
nand UO_1352 (O_1352,N_18898,N_19384);
xnor UO_1353 (O_1353,N_18533,N_19628);
nand UO_1354 (O_1354,N_19537,N_18573);
xnor UO_1355 (O_1355,N_18849,N_19873);
nor UO_1356 (O_1356,N_19311,N_18099);
or UO_1357 (O_1357,N_19369,N_19931);
nand UO_1358 (O_1358,N_19662,N_18241);
xor UO_1359 (O_1359,N_19024,N_19397);
and UO_1360 (O_1360,N_19591,N_19117);
nand UO_1361 (O_1361,N_19311,N_19510);
nand UO_1362 (O_1362,N_19713,N_19543);
xnor UO_1363 (O_1363,N_18256,N_18973);
xor UO_1364 (O_1364,N_19413,N_19203);
nand UO_1365 (O_1365,N_18114,N_19404);
and UO_1366 (O_1366,N_19152,N_19269);
nand UO_1367 (O_1367,N_18612,N_18975);
and UO_1368 (O_1368,N_19257,N_18925);
nor UO_1369 (O_1369,N_18397,N_19675);
nand UO_1370 (O_1370,N_19694,N_18734);
nor UO_1371 (O_1371,N_19683,N_19950);
or UO_1372 (O_1372,N_18726,N_18401);
xor UO_1373 (O_1373,N_19905,N_18231);
nand UO_1374 (O_1374,N_19856,N_18228);
and UO_1375 (O_1375,N_18669,N_19186);
and UO_1376 (O_1376,N_19520,N_18447);
nand UO_1377 (O_1377,N_19469,N_18165);
xnor UO_1378 (O_1378,N_18426,N_18044);
nor UO_1379 (O_1379,N_19583,N_19118);
nor UO_1380 (O_1380,N_19735,N_19763);
xnor UO_1381 (O_1381,N_19550,N_19343);
or UO_1382 (O_1382,N_18756,N_18550);
nand UO_1383 (O_1383,N_19405,N_18830);
nor UO_1384 (O_1384,N_19857,N_18035);
or UO_1385 (O_1385,N_18726,N_18902);
or UO_1386 (O_1386,N_18841,N_18007);
xor UO_1387 (O_1387,N_18661,N_19573);
and UO_1388 (O_1388,N_19949,N_19654);
nor UO_1389 (O_1389,N_19653,N_19940);
or UO_1390 (O_1390,N_18983,N_19122);
nand UO_1391 (O_1391,N_18029,N_19884);
and UO_1392 (O_1392,N_18530,N_18884);
nand UO_1393 (O_1393,N_18861,N_19545);
nand UO_1394 (O_1394,N_18479,N_18869);
nand UO_1395 (O_1395,N_18684,N_19650);
nand UO_1396 (O_1396,N_18006,N_19108);
xnor UO_1397 (O_1397,N_18040,N_19168);
and UO_1398 (O_1398,N_19943,N_19655);
nor UO_1399 (O_1399,N_18969,N_18691);
nor UO_1400 (O_1400,N_18336,N_19722);
and UO_1401 (O_1401,N_18937,N_18774);
nor UO_1402 (O_1402,N_18997,N_18772);
and UO_1403 (O_1403,N_19729,N_19918);
and UO_1404 (O_1404,N_19525,N_18708);
nor UO_1405 (O_1405,N_19344,N_18648);
and UO_1406 (O_1406,N_19284,N_19859);
xnor UO_1407 (O_1407,N_19055,N_19013);
xnor UO_1408 (O_1408,N_19202,N_19597);
and UO_1409 (O_1409,N_18191,N_19186);
or UO_1410 (O_1410,N_19810,N_18352);
or UO_1411 (O_1411,N_18245,N_19460);
xnor UO_1412 (O_1412,N_18242,N_18454);
nand UO_1413 (O_1413,N_18555,N_19399);
and UO_1414 (O_1414,N_19887,N_19657);
or UO_1415 (O_1415,N_18902,N_19890);
or UO_1416 (O_1416,N_19221,N_18699);
nor UO_1417 (O_1417,N_18818,N_19449);
xnor UO_1418 (O_1418,N_18055,N_18887);
and UO_1419 (O_1419,N_18544,N_18570);
nor UO_1420 (O_1420,N_19247,N_18191);
and UO_1421 (O_1421,N_18342,N_19788);
and UO_1422 (O_1422,N_18419,N_19706);
or UO_1423 (O_1423,N_18992,N_19037);
nor UO_1424 (O_1424,N_19034,N_18880);
and UO_1425 (O_1425,N_19960,N_19602);
or UO_1426 (O_1426,N_19160,N_18839);
xnor UO_1427 (O_1427,N_18561,N_19347);
nor UO_1428 (O_1428,N_19904,N_18257);
or UO_1429 (O_1429,N_18995,N_18165);
and UO_1430 (O_1430,N_19259,N_19406);
or UO_1431 (O_1431,N_19638,N_19958);
and UO_1432 (O_1432,N_19103,N_19684);
and UO_1433 (O_1433,N_18434,N_19820);
or UO_1434 (O_1434,N_19786,N_19433);
xnor UO_1435 (O_1435,N_19600,N_18277);
nand UO_1436 (O_1436,N_18150,N_18173);
and UO_1437 (O_1437,N_18657,N_19855);
nor UO_1438 (O_1438,N_19687,N_18315);
and UO_1439 (O_1439,N_19632,N_18986);
and UO_1440 (O_1440,N_19276,N_19603);
or UO_1441 (O_1441,N_19925,N_19761);
nor UO_1442 (O_1442,N_18080,N_18200);
and UO_1443 (O_1443,N_18591,N_19149);
nor UO_1444 (O_1444,N_19969,N_18828);
and UO_1445 (O_1445,N_19885,N_18962);
and UO_1446 (O_1446,N_18672,N_18718);
and UO_1447 (O_1447,N_18148,N_18857);
nor UO_1448 (O_1448,N_18171,N_18517);
nand UO_1449 (O_1449,N_19176,N_19518);
and UO_1450 (O_1450,N_19161,N_19148);
nor UO_1451 (O_1451,N_19577,N_18614);
and UO_1452 (O_1452,N_18680,N_19662);
nor UO_1453 (O_1453,N_19472,N_18067);
and UO_1454 (O_1454,N_19749,N_19469);
and UO_1455 (O_1455,N_18598,N_19270);
nand UO_1456 (O_1456,N_18632,N_19673);
and UO_1457 (O_1457,N_19467,N_19282);
and UO_1458 (O_1458,N_19985,N_18439);
nand UO_1459 (O_1459,N_19877,N_18950);
nand UO_1460 (O_1460,N_18269,N_18989);
or UO_1461 (O_1461,N_18682,N_18105);
or UO_1462 (O_1462,N_18254,N_19417);
and UO_1463 (O_1463,N_18867,N_18539);
nor UO_1464 (O_1464,N_19625,N_19477);
or UO_1465 (O_1465,N_19521,N_19748);
and UO_1466 (O_1466,N_18840,N_19565);
xor UO_1467 (O_1467,N_18416,N_19061);
nor UO_1468 (O_1468,N_19438,N_18354);
nand UO_1469 (O_1469,N_19162,N_19651);
or UO_1470 (O_1470,N_18126,N_18547);
nand UO_1471 (O_1471,N_18511,N_18948);
nand UO_1472 (O_1472,N_19674,N_18504);
or UO_1473 (O_1473,N_19188,N_19838);
nand UO_1474 (O_1474,N_19410,N_19971);
nor UO_1475 (O_1475,N_19273,N_18008);
nand UO_1476 (O_1476,N_19267,N_19972);
nand UO_1477 (O_1477,N_18184,N_18296);
or UO_1478 (O_1478,N_18787,N_19150);
or UO_1479 (O_1479,N_18169,N_19575);
or UO_1480 (O_1480,N_19953,N_19690);
xor UO_1481 (O_1481,N_19499,N_18170);
nor UO_1482 (O_1482,N_18452,N_19614);
nor UO_1483 (O_1483,N_18793,N_19932);
nor UO_1484 (O_1484,N_18053,N_18600);
or UO_1485 (O_1485,N_19478,N_19041);
or UO_1486 (O_1486,N_19385,N_18286);
nand UO_1487 (O_1487,N_18326,N_18124);
or UO_1488 (O_1488,N_18833,N_18048);
and UO_1489 (O_1489,N_19343,N_18025);
xor UO_1490 (O_1490,N_19925,N_19201);
nor UO_1491 (O_1491,N_19866,N_19415);
nor UO_1492 (O_1492,N_19163,N_19906);
nor UO_1493 (O_1493,N_18882,N_19180);
and UO_1494 (O_1494,N_19112,N_18853);
and UO_1495 (O_1495,N_19855,N_19556);
nand UO_1496 (O_1496,N_18207,N_19977);
nor UO_1497 (O_1497,N_18834,N_18904);
and UO_1498 (O_1498,N_18567,N_18304);
nand UO_1499 (O_1499,N_19466,N_18997);
and UO_1500 (O_1500,N_18195,N_19638);
nand UO_1501 (O_1501,N_18030,N_19632);
nand UO_1502 (O_1502,N_19313,N_19285);
nor UO_1503 (O_1503,N_19368,N_19720);
nand UO_1504 (O_1504,N_18577,N_18270);
nand UO_1505 (O_1505,N_18643,N_19790);
nand UO_1506 (O_1506,N_18158,N_19839);
or UO_1507 (O_1507,N_18185,N_18402);
nor UO_1508 (O_1508,N_18463,N_19644);
xnor UO_1509 (O_1509,N_19769,N_18145);
nand UO_1510 (O_1510,N_18945,N_18022);
xor UO_1511 (O_1511,N_18099,N_18247);
nand UO_1512 (O_1512,N_19616,N_18990);
nor UO_1513 (O_1513,N_18374,N_19962);
nor UO_1514 (O_1514,N_19483,N_19289);
and UO_1515 (O_1515,N_18374,N_18007);
nor UO_1516 (O_1516,N_18676,N_18344);
nor UO_1517 (O_1517,N_18708,N_19258);
or UO_1518 (O_1518,N_18024,N_19391);
or UO_1519 (O_1519,N_18047,N_18234);
or UO_1520 (O_1520,N_18523,N_18418);
or UO_1521 (O_1521,N_18114,N_18671);
or UO_1522 (O_1522,N_19022,N_19528);
nand UO_1523 (O_1523,N_18480,N_18476);
or UO_1524 (O_1524,N_19195,N_18115);
nand UO_1525 (O_1525,N_19214,N_18940);
nand UO_1526 (O_1526,N_19523,N_19974);
nand UO_1527 (O_1527,N_18697,N_18305);
nand UO_1528 (O_1528,N_19293,N_18318);
nand UO_1529 (O_1529,N_19762,N_18779);
or UO_1530 (O_1530,N_18370,N_19945);
nand UO_1531 (O_1531,N_19048,N_18526);
or UO_1532 (O_1532,N_19763,N_18072);
nand UO_1533 (O_1533,N_18040,N_19940);
xor UO_1534 (O_1534,N_19631,N_19160);
and UO_1535 (O_1535,N_19814,N_19635);
nand UO_1536 (O_1536,N_18663,N_18638);
nor UO_1537 (O_1537,N_19490,N_19735);
nor UO_1538 (O_1538,N_18576,N_19973);
or UO_1539 (O_1539,N_19333,N_18724);
nor UO_1540 (O_1540,N_18835,N_19644);
and UO_1541 (O_1541,N_19516,N_18843);
or UO_1542 (O_1542,N_19534,N_19243);
nand UO_1543 (O_1543,N_18166,N_18483);
nand UO_1544 (O_1544,N_19638,N_19885);
and UO_1545 (O_1545,N_18666,N_19488);
nor UO_1546 (O_1546,N_19757,N_19091);
and UO_1547 (O_1547,N_19974,N_19562);
nor UO_1548 (O_1548,N_18643,N_18817);
nand UO_1549 (O_1549,N_19968,N_18219);
or UO_1550 (O_1550,N_18815,N_18621);
or UO_1551 (O_1551,N_18578,N_18795);
xnor UO_1552 (O_1552,N_18554,N_18351);
nor UO_1553 (O_1553,N_18726,N_19940);
nor UO_1554 (O_1554,N_18082,N_18309);
nor UO_1555 (O_1555,N_19458,N_19486);
and UO_1556 (O_1556,N_18967,N_18070);
and UO_1557 (O_1557,N_18951,N_18251);
and UO_1558 (O_1558,N_19058,N_18202);
xor UO_1559 (O_1559,N_19826,N_19707);
and UO_1560 (O_1560,N_18165,N_19912);
and UO_1561 (O_1561,N_19934,N_19111);
nand UO_1562 (O_1562,N_19463,N_18629);
and UO_1563 (O_1563,N_18932,N_19439);
nand UO_1564 (O_1564,N_18401,N_18987);
nor UO_1565 (O_1565,N_19908,N_19016);
and UO_1566 (O_1566,N_19914,N_19281);
and UO_1567 (O_1567,N_19951,N_19694);
and UO_1568 (O_1568,N_18421,N_18790);
and UO_1569 (O_1569,N_19079,N_19063);
and UO_1570 (O_1570,N_19691,N_18676);
nand UO_1571 (O_1571,N_19893,N_18512);
or UO_1572 (O_1572,N_19188,N_18539);
nand UO_1573 (O_1573,N_19517,N_19010);
xor UO_1574 (O_1574,N_19114,N_18346);
nand UO_1575 (O_1575,N_18329,N_19951);
xor UO_1576 (O_1576,N_18808,N_19480);
nand UO_1577 (O_1577,N_18999,N_19022);
and UO_1578 (O_1578,N_19344,N_18595);
nand UO_1579 (O_1579,N_18511,N_19072);
nor UO_1580 (O_1580,N_18091,N_18052);
or UO_1581 (O_1581,N_19707,N_18174);
nor UO_1582 (O_1582,N_18238,N_19513);
nor UO_1583 (O_1583,N_19744,N_18436);
nor UO_1584 (O_1584,N_18448,N_18492);
nand UO_1585 (O_1585,N_19133,N_18226);
xor UO_1586 (O_1586,N_18153,N_19030);
and UO_1587 (O_1587,N_18502,N_18993);
or UO_1588 (O_1588,N_18555,N_19702);
or UO_1589 (O_1589,N_18430,N_18636);
nor UO_1590 (O_1590,N_19084,N_19743);
nand UO_1591 (O_1591,N_19058,N_18504);
xor UO_1592 (O_1592,N_19326,N_19123);
nand UO_1593 (O_1593,N_18280,N_19196);
nand UO_1594 (O_1594,N_18184,N_18297);
nand UO_1595 (O_1595,N_19179,N_19562);
and UO_1596 (O_1596,N_18423,N_19335);
and UO_1597 (O_1597,N_19130,N_19210);
nand UO_1598 (O_1598,N_18266,N_19815);
and UO_1599 (O_1599,N_18290,N_19146);
or UO_1600 (O_1600,N_18571,N_19503);
or UO_1601 (O_1601,N_19128,N_18206);
and UO_1602 (O_1602,N_18406,N_18742);
or UO_1603 (O_1603,N_19870,N_18811);
nor UO_1604 (O_1604,N_18236,N_18569);
or UO_1605 (O_1605,N_19184,N_19749);
nor UO_1606 (O_1606,N_19316,N_19445);
and UO_1607 (O_1607,N_18727,N_19818);
nand UO_1608 (O_1608,N_19415,N_19400);
nor UO_1609 (O_1609,N_19140,N_19480);
or UO_1610 (O_1610,N_19438,N_19106);
xnor UO_1611 (O_1611,N_18671,N_19018);
nand UO_1612 (O_1612,N_19080,N_19474);
or UO_1613 (O_1613,N_19288,N_19993);
or UO_1614 (O_1614,N_19232,N_19705);
nand UO_1615 (O_1615,N_18310,N_19273);
and UO_1616 (O_1616,N_18728,N_18027);
or UO_1617 (O_1617,N_19565,N_19457);
and UO_1618 (O_1618,N_19639,N_19638);
and UO_1619 (O_1619,N_19020,N_18359);
nand UO_1620 (O_1620,N_19308,N_18160);
xnor UO_1621 (O_1621,N_19128,N_18903);
and UO_1622 (O_1622,N_18430,N_18322);
or UO_1623 (O_1623,N_19815,N_19017);
nand UO_1624 (O_1624,N_18286,N_19525);
or UO_1625 (O_1625,N_18435,N_19538);
and UO_1626 (O_1626,N_19952,N_19832);
nand UO_1627 (O_1627,N_18741,N_19656);
nand UO_1628 (O_1628,N_19350,N_18391);
and UO_1629 (O_1629,N_18820,N_18762);
and UO_1630 (O_1630,N_19906,N_18796);
and UO_1631 (O_1631,N_19866,N_18373);
nand UO_1632 (O_1632,N_19011,N_18149);
and UO_1633 (O_1633,N_18582,N_18322);
and UO_1634 (O_1634,N_19898,N_19383);
or UO_1635 (O_1635,N_19937,N_18406);
nand UO_1636 (O_1636,N_19867,N_19841);
and UO_1637 (O_1637,N_19912,N_18901);
nand UO_1638 (O_1638,N_19077,N_18667);
nand UO_1639 (O_1639,N_19431,N_18948);
or UO_1640 (O_1640,N_19645,N_19670);
or UO_1641 (O_1641,N_19334,N_19289);
nand UO_1642 (O_1642,N_19722,N_19396);
and UO_1643 (O_1643,N_19918,N_19493);
or UO_1644 (O_1644,N_19884,N_18446);
or UO_1645 (O_1645,N_18956,N_19015);
xor UO_1646 (O_1646,N_18050,N_18585);
or UO_1647 (O_1647,N_19565,N_18740);
nand UO_1648 (O_1648,N_18358,N_18536);
or UO_1649 (O_1649,N_18746,N_19141);
nand UO_1650 (O_1650,N_18458,N_19957);
and UO_1651 (O_1651,N_18209,N_18623);
nand UO_1652 (O_1652,N_19503,N_18832);
or UO_1653 (O_1653,N_18796,N_18342);
nor UO_1654 (O_1654,N_19878,N_18192);
or UO_1655 (O_1655,N_18475,N_18478);
and UO_1656 (O_1656,N_19930,N_19319);
and UO_1657 (O_1657,N_19132,N_18463);
nand UO_1658 (O_1658,N_18097,N_18903);
and UO_1659 (O_1659,N_18984,N_19055);
xor UO_1660 (O_1660,N_18653,N_18588);
xnor UO_1661 (O_1661,N_19017,N_19243);
nand UO_1662 (O_1662,N_18110,N_18338);
nand UO_1663 (O_1663,N_19253,N_18974);
and UO_1664 (O_1664,N_18437,N_19068);
nand UO_1665 (O_1665,N_19437,N_19886);
nor UO_1666 (O_1666,N_19320,N_19100);
nand UO_1667 (O_1667,N_18040,N_18447);
nor UO_1668 (O_1668,N_18904,N_18591);
nand UO_1669 (O_1669,N_18050,N_19738);
and UO_1670 (O_1670,N_19376,N_18811);
nor UO_1671 (O_1671,N_18336,N_19161);
nand UO_1672 (O_1672,N_18459,N_19529);
or UO_1673 (O_1673,N_19588,N_19668);
nand UO_1674 (O_1674,N_18936,N_18874);
nor UO_1675 (O_1675,N_18163,N_18729);
and UO_1676 (O_1676,N_19072,N_18689);
xnor UO_1677 (O_1677,N_19106,N_19600);
xor UO_1678 (O_1678,N_19020,N_18829);
or UO_1679 (O_1679,N_18152,N_18361);
nor UO_1680 (O_1680,N_19787,N_19437);
or UO_1681 (O_1681,N_19995,N_19490);
or UO_1682 (O_1682,N_19574,N_18884);
or UO_1683 (O_1683,N_18804,N_18236);
or UO_1684 (O_1684,N_18088,N_18020);
and UO_1685 (O_1685,N_19253,N_19451);
nand UO_1686 (O_1686,N_19385,N_19151);
xor UO_1687 (O_1687,N_19873,N_19110);
and UO_1688 (O_1688,N_19875,N_18207);
xor UO_1689 (O_1689,N_19842,N_18301);
or UO_1690 (O_1690,N_18029,N_19877);
xor UO_1691 (O_1691,N_19921,N_18706);
or UO_1692 (O_1692,N_19751,N_19221);
nor UO_1693 (O_1693,N_18088,N_19228);
and UO_1694 (O_1694,N_19362,N_18968);
nand UO_1695 (O_1695,N_19476,N_18761);
nor UO_1696 (O_1696,N_19634,N_19912);
nor UO_1697 (O_1697,N_19271,N_18139);
nor UO_1698 (O_1698,N_19244,N_18004);
and UO_1699 (O_1699,N_18345,N_19704);
nand UO_1700 (O_1700,N_19961,N_19190);
nand UO_1701 (O_1701,N_19265,N_19024);
nor UO_1702 (O_1702,N_18785,N_19572);
or UO_1703 (O_1703,N_18671,N_18387);
or UO_1704 (O_1704,N_19229,N_19322);
and UO_1705 (O_1705,N_19489,N_18911);
nand UO_1706 (O_1706,N_18775,N_19854);
xnor UO_1707 (O_1707,N_18961,N_19718);
nor UO_1708 (O_1708,N_18595,N_19473);
xor UO_1709 (O_1709,N_18443,N_19076);
nand UO_1710 (O_1710,N_18985,N_19246);
or UO_1711 (O_1711,N_19931,N_18667);
xor UO_1712 (O_1712,N_19116,N_18609);
nand UO_1713 (O_1713,N_18500,N_18539);
and UO_1714 (O_1714,N_19592,N_19923);
or UO_1715 (O_1715,N_19058,N_18333);
or UO_1716 (O_1716,N_19550,N_18000);
or UO_1717 (O_1717,N_19035,N_19379);
or UO_1718 (O_1718,N_18437,N_19293);
nor UO_1719 (O_1719,N_19432,N_18012);
nor UO_1720 (O_1720,N_19832,N_18380);
xnor UO_1721 (O_1721,N_19830,N_19077);
nand UO_1722 (O_1722,N_19318,N_19480);
and UO_1723 (O_1723,N_18456,N_19135);
and UO_1724 (O_1724,N_18438,N_18227);
or UO_1725 (O_1725,N_18909,N_19609);
nor UO_1726 (O_1726,N_19989,N_18905);
nor UO_1727 (O_1727,N_18955,N_18882);
nor UO_1728 (O_1728,N_19289,N_18265);
xor UO_1729 (O_1729,N_19406,N_19852);
xnor UO_1730 (O_1730,N_19892,N_18078);
xor UO_1731 (O_1731,N_19911,N_19044);
nand UO_1732 (O_1732,N_19353,N_18127);
nor UO_1733 (O_1733,N_18784,N_18612);
and UO_1734 (O_1734,N_19529,N_18984);
and UO_1735 (O_1735,N_19940,N_19904);
or UO_1736 (O_1736,N_19491,N_19323);
and UO_1737 (O_1737,N_19444,N_18299);
nor UO_1738 (O_1738,N_18653,N_19801);
and UO_1739 (O_1739,N_19882,N_19146);
nand UO_1740 (O_1740,N_19088,N_19521);
nand UO_1741 (O_1741,N_18329,N_18951);
or UO_1742 (O_1742,N_18791,N_18001);
xnor UO_1743 (O_1743,N_19298,N_18369);
or UO_1744 (O_1744,N_19852,N_18419);
and UO_1745 (O_1745,N_18828,N_18736);
nor UO_1746 (O_1746,N_19472,N_18236);
nor UO_1747 (O_1747,N_18400,N_18927);
nand UO_1748 (O_1748,N_18923,N_18740);
xnor UO_1749 (O_1749,N_19135,N_18208);
or UO_1750 (O_1750,N_18940,N_19553);
or UO_1751 (O_1751,N_19160,N_19944);
or UO_1752 (O_1752,N_18661,N_19854);
nand UO_1753 (O_1753,N_19465,N_18311);
nand UO_1754 (O_1754,N_18001,N_18666);
or UO_1755 (O_1755,N_19551,N_18160);
or UO_1756 (O_1756,N_18737,N_19347);
or UO_1757 (O_1757,N_19388,N_19431);
nand UO_1758 (O_1758,N_19392,N_18928);
xnor UO_1759 (O_1759,N_19686,N_19242);
or UO_1760 (O_1760,N_19999,N_18197);
and UO_1761 (O_1761,N_18261,N_18187);
or UO_1762 (O_1762,N_19980,N_18918);
or UO_1763 (O_1763,N_19241,N_19742);
nor UO_1764 (O_1764,N_19305,N_19594);
and UO_1765 (O_1765,N_19867,N_18353);
xor UO_1766 (O_1766,N_18748,N_19273);
or UO_1767 (O_1767,N_18898,N_18023);
or UO_1768 (O_1768,N_18515,N_19547);
nor UO_1769 (O_1769,N_19392,N_19873);
nand UO_1770 (O_1770,N_18161,N_19978);
and UO_1771 (O_1771,N_18503,N_18688);
and UO_1772 (O_1772,N_19584,N_19559);
or UO_1773 (O_1773,N_18012,N_19975);
nor UO_1774 (O_1774,N_19770,N_18788);
nand UO_1775 (O_1775,N_18967,N_18425);
or UO_1776 (O_1776,N_18942,N_19253);
and UO_1777 (O_1777,N_19655,N_19105);
nand UO_1778 (O_1778,N_18898,N_18391);
nor UO_1779 (O_1779,N_18709,N_19189);
nor UO_1780 (O_1780,N_19156,N_18187);
nor UO_1781 (O_1781,N_18476,N_19195);
and UO_1782 (O_1782,N_18879,N_18507);
xnor UO_1783 (O_1783,N_18280,N_18218);
or UO_1784 (O_1784,N_19262,N_19648);
nand UO_1785 (O_1785,N_19322,N_19691);
and UO_1786 (O_1786,N_18978,N_18554);
or UO_1787 (O_1787,N_19006,N_18796);
and UO_1788 (O_1788,N_19625,N_18633);
nand UO_1789 (O_1789,N_19005,N_19440);
xor UO_1790 (O_1790,N_19823,N_19504);
nor UO_1791 (O_1791,N_18849,N_18348);
and UO_1792 (O_1792,N_19162,N_19289);
nand UO_1793 (O_1793,N_18679,N_19582);
nor UO_1794 (O_1794,N_19681,N_19955);
nand UO_1795 (O_1795,N_18810,N_19638);
and UO_1796 (O_1796,N_18435,N_18696);
nand UO_1797 (O_1797,N_19888,N_19623);
or UO_1798 (O_1798,N_19235,N_19303);
and UO_1799 (O_1799,N_19015,N_18483);
nand UO_1800 (O_1800,N_18866,N_18661);
xor UO_1801 (O_1801,N_19931,N_19246);
xor UO_1802 (O_1802,N_19741,N_18033);
nand UO_1803 (O_1803,N_19995,N_18363);
nor UO_1804 (O_1804,N_19206,N_18017);
nand UO_1805 (O_1805,N_19516,N_18186);
nand UO_1806 (O_1806,N_18016,N_19981);
nor UO_1807 (O_1807,N_18071,N_18863);
nor UO_1808 (O_1808,N_19053,N_19718);
nor UO_1809 (O_1809,N_18300,N_18717);
nand UO_1810 (O_1810,N_19887,N_18595);
and UO_1811 (O_1811,N_18163,N_19044);
xnor UO_1812 (O_1812,N_19823,N_19954);
and UO_1813 (O_1813,N_19916,N_19663);
nand UO_1814 (O_1814,N_19884,N_18764);
xor UO_1815 (O_1815,N_19067,N_18723);
and UO_1816 (O_1816,N_19709,N_18499);
nor UO_1817 (O_1817,N_18871,N_18636);
nand UO_1818 (O_1818,N_19188,N_19654);
nand UO_1819 (O_1819,N_18806,N_18249);
xnor UO_1820 (O_1820,N_19249,N_19686);
and UO_1821 (O_1821,N_18655,N_18168);
or UO_1822 (O_1822,N_18566,N_18693);
nor UO_1823 (O_1823,N_19569,N_19028);
or UO_1824 (O_1824,N_19471,N_19463);
and UO_1825 (O_1825,N_18958,N_19076);
or UO_1826 (O_1826,N_18152,N_18388);
nand UO_1827 (O_1827,N_19704,N_19035);
or UO_1828 (O_1828,N_19603,N_18506);
or UO_1829 (O_1829,N_18635,N_19407);
nor UO_1830 (O_1830,N_19334,N_18109);
and UO_1831 (O_1831,N_18458,N_18967);
nand UO_1832 (O_1832,N_19957,N_18616);
nor UO_1833 (O_1833,N_18544,N_18319);
or UO_1834 (O_1834,N_19998,N_19801);
nor UO_1835 (O_1835,N_18514,N_19674);
nor UO_1836 (O_1836,N_18129,N_19981);
and UO_1837 (O_1837,N_18293,N_18609);
nor UO_1838 (O_1838,N_19821,N_18848);
nand UO_1839 (O_1839,N_18157,N_19377);
nand UO_1840 (O_1840,N_19186,N_19932);
nor UO_1841 (O_1841,N_19895,N_19123);
nand UO_1842 (O_1842,N_18758,N_19945);
nor UO_1843 (O_1843,N_19572,N_19025);
or UO_1844 (O_1844,N_19032,N_18094);
nand UO_1845 (O_1845,N_19389,N_18374);
and UO_1846 (O_1846,N_19933,N_19246);
nor UO_1847 (O_1847,N_19424,N_19102);
and UO_1848 (O_1848,N_19476,N_19558);
or UO_1849 (O_1849,N_18747,N_19271);
and UO_1850 (O_1850,N_19432,N_19237);
nor UO_1851 (O_1851,N_18086,N_19646);
nor UO_1852 (O_1852,N_18415,N_19944);
or UO_1853 (O_1853,N_19609,N_18218);
and UO_1854 (O_1854,N_18585,N_19319);
nand UO_1855 (O_1855,N_19952,N_19005);
nor UO_1856 (O_1856,N_19077,N_19325);
or UO_1857 (O_1857,N_18143,N_18658);
or UO_1858 (O_1858,N_18073,N_19975);
and UO_1859 (O_1859,N_19722,N_19865);
nor UO_1860 (O_1860,N_18927,N_18662);
and UO_1861 (O_1861,N_18023,N_18056);
and UO_1862 (O_1862,N_19884,N_18668);
or UO_1863 (O_1863,N_19816,N_18447);
xnor UO_1864 (O_1864,N_19919,N_18563);
and UO_1865 (O_1865,N_19790,N_18401);
xor UO_1866 (O_1866,N_19328,N_18366);
nor UO_1867 (O_1867,N_19429,N_18183);
or UO_1868 (O_1868,N_19173,N_18367);
nand UO_1869 (O_1869,N_19975,N_18747);
nor UO_1870 (O_1870,N_18151,N_19123);
or UO_1871 (O_1871,N_19224,N_18638);
nor UO_1872 (O_1872,N_18393,N_19216);
xnor UO_1873 (O_1873,N_19152,N_19615);
nor UO_1874 (O_1874,N_19213,N_18619);
nor UO_1875 (O_1875,N_19231,N_18052);
nor UO_1876 (O_1876,N_19324,N_18860);
and UO_1877 (O_1877,N_19595,N_18228);
xor UO_1878 (O_1878,N_18215,N_19793);
nand UO_1879 (O_1879,N_18240,N_19058);
and UO_1880 (O_1880,N_19163,N_18913);
or UO_1881 (O_1881,N_18772,N_19310);
nor UO_1882 (O_1882,N_18681,N_19632);
nor UO_1883 (O_1883,N_19519,N_19931);
xnor UO_1884 (O_1884,N_19331,N_19947);
and UO_1885 (O_1885,N_19994,N_18111);
and UO_1886 (O_1886,N_18118,N_19313);
or UO_1887 (O_1887,N_18055,N_18610);
nor UO_1888 (O_1888,N_19470,N_19655);
and UO_1889 (O_1889,N_18334,N_19652);
nand UO_1890 (O_1890,N_19781,N_19026);
and UO_1891 (O_1891,N_18317,N_18882);
and UO_1892 (O_1892,N_19010,N_19780);
nand UO_1893 (O_1893,N_18669,N_18316);
nor UO_1894 (O_1894,N_19399,N_18932);
xor UO_1895 (O_1895,N_18669,N_18599);
nand UO_1896 (O_1896,N_19473,N_19908);
nor UO_1897 (O_1897,N_19867,N_19478);
and UO_1898 (O_1898,N_19904,N_19683);
nand UO_1899 (O_1899,N_19614,N_18614);
or UO_1900 (O_1900,N_18829,N_19820);
xor UO_1901 (O_1901,N_19735,N_18197);
nor UO_1902 (O_1902,N_19090,N_19793);
nor UO_1903 (O_1903,N_18760,N_18832);
or UO_1904 (O_1904,N_19712,N_19394);
nor UO_1905 (O_1905,N_18930,N_18254);
and UO_1906 (O_1906,N_18001,N_19967);
nand UO_1907 (O_1907,N_19401,N_18188);
or UO_1908 (O_1908,N_19556,N_19613);
nand UO_1909 (O_1909,N_18181,N_18633);
nand UO_1910 (O_1910,N_19673,N_19846);
or UO_1911 (O_1911,N_18698,N_19931);
and UO_1912 (O_1912,N_18769,N_18983);
nand UO_1913 (O_1913,N_18220,N_19106);
or UO_1914 (O_1914,N_18980,N_18004);
or UO_1915 (O_1915,N_19645,N_19332);
nor UO_1916 (O_1916,N_19939,N_19832);
nor UO_1917 (O_1917,N_18747,N_19692);
xnor UO_1918 (O_1918,N_19435,N_19535);
nor UO_1919 (O_1919,N_19561,N_19915);
nor UO_1920 (O_1920,N_19493,N_19026);
nor UO_1921 (O_1921,N_18407,N_19752);
nand UO_1922 (O_1922,N_19856,N_19039);
and UO_1923 (O_1923,N_19216,N_18064);
nand UO_1924 (O_1924,N_18328,N_18669);
or UO_1925 (O_1925,N_18873,N_19462);
or UO_1926 (O_1926,N_18689,N_18966);
and UO_1927 (O_1927,N_18282,N_19236);
or UO_1928 (O_1928,N_19634,N_18077);
nor UO_1929 (O_1929,N_19857,N_18723);
or UO_1930 (O_1930,N_19521,N_18760);
nand UO_1931 (O_1931,N_19577,N_18724);
xnor UO_1932 (O_1932,N_18737,N_18857);
xnor UO_1933 (O_1933,N_19279,N_19141);
nor UO_1934 (O_1934,N_18567,N_19183);
nor UO_1935 (O_1935,N_19111,N_19196);
nand UO_1936 (O_1936,N_19934,N_18506);
and UO_1937 (O_1937,N_19942,N_18488);
xnor UO_1938 (O_1938,N_19174,N_18702);
nor UO_1939 (O_1939,N_19080,N_18919);
nor UO_1940 (O_1940,N_19800,N_18364);
nand UO_1941 (O_1941,N_19916,N_18548);
or UO_1942 (O_1942,N_19261,N_19583);
nor UO_1943 (O_1943,N_19032,N_18047);
nand UO_1944 (O_1944,N_19139,N_19421);
or UO_1945 (O_1945,N_19723,N_19654);
nor UO_1946 (O_1946,N_18936,N_18841);
and UO_1947 (O_1947,N_18125,N_19759);
xor UO_1948 (O_1948,N_19133,N_18928);
nand UO_1949 (O_1949,N_19800,N_19727);
nor UO_1950 (O_1950,N_19160,N_19781);
nand UO_1951 (O_1951,N_18186,N_19820);
or UO_1952 (O_1952,N_18470,N_19460);
nor UO_1953 (O_1953,N_19962,N_19489);
nor UO_1954 (O_1954,N_18683,N_18441);
or UO_1955 (O_1955,N_18286,N_18436);
nand UO_1956 (O_1956,N_18412,N_19525);
or UO_1957 (O_1957,N_19031,N_19798);
and UO_1958 (O_1958,N_18667,N_18963);
nand UO_1959 (O_1959,N_19720,N_18561);
and UO_1960 (O_1960,N_19972,N_19297);
nor UO_1961 (O_1961,N_18219,N_18216);
nor UO_1962 (O_1962,N_19309,N_19914);
nor UO_1963 (O_1963,N_19621,N_18628);
and UO_1964 (O_1964,N_18738,N_19986);
or UO_1965 (O_1965,N_19659,N_18169);
and UO_1966 (O_1966,N_18788,N_18150);
xor UO_1967 (O_1967,N_18226,N_19337);
xnor UO_1968 (O_1968,N_19573,N_19210);
or UO_1969 (O_1969,N_18192,N_19035);
xor UO_1970 (O_1970,N_19811,N_18044);
or UO_1971 (O_1971,N_18190,N_19565);
or UO_1972 (O_1972,N_18708,N_19647);
nor UO_1973 (O_1973,N_19496,N_18937);
and UO_1974 (O_1974,N_19739,N_18459);
nand UO_1975 (O_1975,N_19738,N_18861);
and UO_1976 (O_1976,N_19399,N_19660);
nor UO_1977 (O_1977,N_18941,N_19133);
xor UO_1978 (O_1978,N_18624,N_18302);
nor UO_1979 (O_1979,N_18681,N_18851);
nand UO_1980 (O_1980,N_19290,N_19569);
and UO_1981 (O_1981,N_19164,N_18239);
nand UO_1982 (O_1982,N_18726,N_18621);
and UO_1983 (O_1983,N_18562,N_19254);
and UO_1984 (O_1984,N_18282,N_19190);
xnor UO_1985 (O_1985,N_18168,N_19951);
nand UO_1986 (O_1986,N_18080,N_18189);
nor UO_1987 (O_1987,N_19102,N_18259);
nand UO_1988 (O_1988,N_19250,N_19419);
and UO_1989 (O_1989,N_19879,N_18464);
and UO_1990 (O_1990,N_19854,N_19455);
or UO_1991 (O_1991,N_19032,N_19620);
nor UO_1992 (O_1992,N_18537,N_19365);
nor UO_1993 (O_1993,N_18490,N_18222);
or UO_1994 (O_1994,N_18478,N_19733);
nor UO_1995 (O_1995,N_19368,N_18832);
nand UO_1996 (O_1996,N_19521,N_18016);
nor UO_1997 (O_1997,N_19176,N_18517);
xnor UO_1998 (O_1998,N_19818,N_19342);
nand UO_1999 (O_1999,N_19745,N_19254);
nand UO_2000 (O_2000,N_19933,N_18748);
and UO_2001 (O_2001,N_18022,N_19544);
nand UO_2002 (O_2002,N_19139,N_19640);
nor UO_2003 (O_2003,N_18351,N_18658);
nor UO_2004 (O_2004,N_19159,N_19581);
xor UO_2005 (O_2005,N_18216,N_19502);
and UO_2006 (O_2006,N_19484,N_18160);
or UO_2007 (O_2007,N_19934,N_19396);
or UO_2008 (O_2008,N_19691,N_18329);
nand UO_2009 (O_2009,N_19852,N_19184);
nand UO_2010 (O_2010,N_19258,N_19125);
and UO_2011 (O_2011,N_19189,N_19811);
and UO_2012 (O_2012,N_19454,N_18848);
or UO_2013 (O_2013,N_18665,N_18555);
nor UO_2014 (O_2014,N_19984,N_18453);
nand UO_2015 (O_2015,N_19119,N_19581);
or UO_2016 (O_2016,N_19727,N_18150);
xnor UO_2017 (O_2017,N_19894,N_18645);
nor UO_2018 (O_2018,N_19467,N_18993);
nor UO_2019 (O_2019,N_19309,N_18703);
nor UO_2020 (O_2020,N_18016,N_18031);
or UO_2021 (O_2021,N_19693,N_19106);
or UO_2022 (O_2022,N_18938,N_18276);
and UO_2023 (O_2023,N_18685,N_19742);
nand UO_2024 (O_2024,N_19480,N_19063);
nor UO_2025 (O_2025,N_19658,N_18291);
or UO_2026 (O_2026,N_18722,N_18159);
xnor UO_2027 (O_2027,N_19740,N_18769);
or UO_2028 (O_2028,N_19364,N_19228);
nand UO_2029 (O_2029,N_18126,N_19019);
nand UO_2030 (O_2030,N_19614,N_18171);
and UO_2031 (O_2031,N_18936,N_18259);
nand UO_2032 (O_2032,N_18643,N_18870);
xnor UO_2033 (O_2033,N_19227,N_19824);
xor UO_2034 (O_2034,N_18607,N_18574);
or UO_2035 (O_2035,N_19875,N_19100);
or UO_2036 (O_2036,N_18497,N_18471);
and UO_2037 (O_2037,N_18693,N_18662);
and UO_2038 (O_2038,N_18558,N_19062);
nand UO_2039 (O_2039,N_19162,N_18566);
nor UO_2040 (O_2040,N_19690,N_19067);
or UO_2041 (O_2041,N_19087,N_18304);
or UO_2042 (O_2042,N_18289,N_19146);
or UO_2043 (O_2043,N_18001,N_19724);
and UO_2044 (O_2044,N_18687,N_18646);
nor UO_2045 (O_2045,N_18822,N_19017);
nand UO_2046 (O_2046,N_18721,N_18318);
nand UO_2047 (O_2047,N_18103,N_19014);
or UO_2048 (O_2048,N_18359,N_18585);
nor UO_2049 (O_2049,N_18911,N_18714);
and UO_2050 (O_2050,N_19609,N_18382);
or UO_2051 (O_2051,N_18585,N_19389);
or UO_2052 (O_2052,N_18253,N_18903);
and UO_2053 (O_2053,N_19164,N_19340);
nand UO_2054 (O_2054,N_18710,N_18745);
xor UO_2055 (O_2055,N_19000,N_19597);
or UO_2056 (O_2056,N_18826,N_19599);
xor UO_2057 (O_2057,N_18196,N_19410);
nand UO_2058 (O_2058,N_19913,N_18184);
nor UO_2059 (O_2059,N_18198,N_18337);
nor UO_2060 (O_2060,N_19163,N_18694);
nor UO_2061 (O_2061,N_18727,N_19930);
nand UO_2062 (O_2062,N_18639,N_19858);
or UO_2063 (O_2063,N_18824,N_19515);
or UO_2064 (O_2064,N_19436,N_19217);
or UO_2065 (O_2065,N_18142,N_19438);
nor UO_2066 (O_2066,N_18448,N_18961);
or UO_2067 (O_2067,N_18817,N_18044);
nand UO_2068 (O_2068,N_18058,N_18080);
nand UO_2069 (O_2069,N_19122,N_18320);
xnor UO_2070 (O_2070,N_18981,N_18185);
nand UO_2071 (O_2071,N_19840,N_19047);
nand UO_2072 (O_2072,N_19362,N_18265);
nand UO_2073 (O_2073,N_19154,N_19617);
nor UO_2074 (O_2074,N_19350,N_19536);
nand UO_2075 (O_2075,N_18052,N_19110);
xor UO_2076 (O_2076,N_18019,N_18407);
and UO_2077 (O_2077,N_18962,N_18161);
nand UO_2078 (O_2078,N_18964,N_18744);
or UO_2079 (O_2079,N_19240,N_18858);
nand UO_2080 (O_2080,N_18306,N_19015);
nand UO_2081 (O_2081,N_19106,N_19404);
nand UO_2082 (O_2082,N_18973,N_18943);
xnor UO_2083 (O_2083,N_19702,N_18627);
and UO_2084 (O_2084,N_18366,N_19171);
nand UO_2085 (O_2085,N_19171,N_18179);
and UO_2086 (O_2086,N_18824,N_19402);
nand UO_2087 (O_2087,N_18608,N_18452);
and UO_2088 (O_2088,N_19606,N_18969);
and UO_2089 (O_2089,N_18750,N_19209);
nor UO_2090 (O_2090,N_19992,N_18030);
nor UO_2091 (O_2091,N_19022,N_18638);
and UO_2092 (O_2092,N_19367,N_18868);
nor UO_2093 (O_2093,N_18605,N_18447);
xor UO_2094 (O_2094,N_19848,N_18185);
or UO_2095 (O_2095,N_19175,N_18582);
or UO_2096 (O_2096,N_19862,N_18128);
nor UO_2097 (O_2097,N_18661,N_19927);
and UO_2098 (O_2098,N_18215,N_19056);
and UO_2099 (O_2099,N_19851,N_19854);
nor UO_2100 (O_2100,N_18705,N_18334);
or UO_2101 (O_2101,N_18956,N_18066);
or UO_2102 (O_2102,N_19893,N_19327);
nand UO_2103 (O_2103,N_18001,N_19083);
or UO_2104 (O_2104,N_18903,N_18913);
or UO_2105 (O_2105,N_18508,N_18726);
xnor UO_2106 (O_2106,N_18448,N_18002);
or UO_2107 (O_2107,N_19525,N_19989);
nor UO_2108 (O_2108,N_19183,N_19310);
or UO_2109 (O_2109,N_18589,N_18481);
and UO_2110 (O_2110,N_18261,N_18616);
xnor UO_2111 (O_2111,N_19822,N_18704);
or UO_2112 (O_2112,N_19903,N_18596);
and UO_2113 (O_2113,N_18201,N_19016);
or UO_2114 (O_2114,N_19868,N_19616);
nand UO_2115 (O_2115,N_18730,N_19700);
or UO_2116 (O_2116,N_18210,N_19016);
and UO_2117 (O_2117,N_19599,N_18915);
nand UO_2118 (O_2118,N_19926,N_19596);
nand UO_2119 (O_2119,N_19578,N_18660);
and UO_2120 (O_2120,N_18021,N_18352);
xor UO_2121 (O_2121,N_18489,N_19608);
nor UO_2122 (O_2122,N_19847,N_19254);
nand UO_2123 (O_2123,N_18704,N_18586);
or UO_2124 (O_2124,N_19837,N_19384);
or UO_2125 (O_2125,N_18550,N_18559);
and UO_2126 (O_2126,N_19404,N_18846);
nor UO_2127 (O_2127,N_18288,N_19505);
xnor UO_2128 (O_2128,N_19769,N_19946);
and UO_2129 (O_2129,N_18425,N_19080);
or UO_2130 (O_2130,N_18827,N_18152);
or UO_2131 (O_2131,N_18425,N_18485);
nand UO_2132 (O_2132,N_18756,N_18368);
nor UO_2133 (O_2133,N_18512,N_19960);
nand UO_2134 (O_2134,N_18545,N_18351);
or UO_2135 (O_2135,N_18025,N_19113);
nor UO_2136 (O_2136,N_19696,N_18524);
xnor UO_2137 (O_2137,N_18511,N_18686);
nor UO_2138 (O_2138,N_18219,N_18537);
or UO_2139 (O_2139,N_19296,N_18294);
or UO_2140 (O_2140,N_19025,N_18086);
or UO_2141 (O_2141,N_19242,N_19271);
or UO_2142 (O_2142,N_19125,N_18629);
nand UO_2143 (O_2143,N_19551,N_18939);
or UO_2144 (O_2144,N_19383,N_19153);
and UO_2145 (O_2145,N_18158,N_18013);
nor UO_2146 (O_2146,N_19767,N_18682);
nor UO_2147 (O_2147,N_18431,N_18960);
and UO_2148 (O_2148,N_19720,N_18016);
or UO_2149 (O_2149,N_18431,N_18188);
nand UO_2150 (O_2150,N_18205,N_18156);
and UO_2151 (O_2151,N_19492,N_19371);
or UO_2152 (O_2152,N_18639,N_18092);
and UO_2153 (O_2153,N_18510,N_19718);
nand UO_2154 (O_2154,N_18035,N_19218);
or UO_2155 (O_2155,N_18353,N_19837);
nand UO_2156 (O_2156,N_19137,N_19370);
or UO_2157 (O_2157,N_19884,N_18478);
xor UO_2158 (O_2158,N_18017,N_19877);
nand UO_2159 (O_2159,N_19325,N_19722);
xor UO_2160 (O_2160,N_19689,N_18236);
and UO_2161 (O_2161,N_19156,N_18957);
and UO_2162 (O_2162,N_19128,N_18107);
nor UO_2163 (O_2163,N_19380,N_19142);
or UO_2164 (O_2164,N_18504,N_18829);
nand UO_2165 (O_2165,N_18843,N_18304);
or UO_2166 (O_2166,N_18175,N_18130);
and UO_2167 (O_2167,N_19415,N_18444);
nor UO_2168 (O_2168,N_19679,N_19516);
xor UO_2169 (O_2169,N_19571,N_18740);
nand UO_2170 (O_2170,N_18740,N_19256);
nand UO_2171 (O_2171,N_19210,N_18747);
nand UO_2172 (O_2172,N_19953,N_18853);
and UO_2173 (O_2173,N_19959,N_19229);
nand UO_2174 (O_2174,N_18353,N_19280);
nand UO_2175 (O_2175,N_19540,N_19607);
nand UO_2176 (O_2176,N_19834,N_19804);
or UO_2177 (O_2177,N_19888,N_18257);
nand UO_2178 (O_2178,N_19568,N_18760);
and UO_2179 (O_2179,N_19023,N_19579);
or UO_2180 (O_2180,N_19155,N_18780);
nand UO_2181 (O_2181,N_18702,N_18174);
nor UO_2182 (O_2182,N_19938,N_18751);
and UO_2183 (O_2183,N_19614,N_18802);
nor UO_2184 (O_2184,N_18298,N_18941);
and UO_2185 (O_2185,N_18634,N_19986);
and UO_2186 (O_2186,N_18529,N_18642);
or UO_2187 (O_2187,N_19102,N_18559);
xor UO_2188 (O_2188,N_18301,N_18467);
or UO_2189 (O_2189,N_18211,N_19897);
nor UO_2190 (O_2190,N_19458,N_18334);
nand UO_2191 (O_2191,N_19569,N_19562);
nor UO_2192 (O_2192,N_18018,N_19483);
nand UO_2193 (O_2193,N_19661,N_19057);
and UO_2194 (O_2194,N_19618,N_19424);
nor UO_2195 (O_2195,N_18708,N_18426);
or UO_2196 (O_2196,N_18663,N_19525);
nand UO_2197 (O_2197,N_19083,N_19452);
and UO_2198 (O_2198,N_18560,N_19761);
and UO_2199 (O_2199,N_19597,N_19572);
or UO_2200 (O_2200,N_18493,N_19859);
nand UO_2201 (O_2201,N_18805,N_18807);
or UO_2202 (O_2202,N_19624,N_19076);
and UO_2203 (O_2203,N_18881,N_18891);
or UO_2204 (O_2204,N_19318,N_19824);
or UO_2205 (O_2205,N_18959,N_18578);
xor UO_2206 (O_2206,N_19635,N_18273);
or UO_2207 (O_2207,N_18905,N_18213);
xnor UO_2208 (O_2208,N_19227,N_18551);
or UO_2209 (O_2209,N_18540,N_19218);
nand UO_2210 (O_2210,N_19149,N_18838);
xnor UO_2211 (O_2211,N_18003,N_18790);
or UO_2212 (O_2212,N_18925,N_19879);
nor UO_2213 (O_2213,N_18841,N_18329);
and UO_2214 (O_2214,N_19103,N_18571);
or UO_2215 (O_2215,N_19468,N_18672);
xnor UO_2216 (O_2216,N_19027,N_18287);
nand UO_2217 (O_2217,N_18353,N_19174);
nor UO_2218 (O_2218,N_18696,N_19333);
nor UO_2219 (O_2219,N_18755,N_18168);
and UO_2220 (O_2220,N_18342,N_18250);
and UO_2221 (O_2221,N_19690,N_19592);
or UO_2222 (O_2222,N_18390,N_18120);
or UO_2223 (O_2223,N_19625,N_18322);
and UO_2224 (O_2224,N_19749,N_19388);
nand UO_2225 (O_2225,N_19917,N_18424);
and UO_2226 (O_2226,N_18302,N_18304);
and UO_2227 (O_2227,N_19767,N_18591);
and UO_2228 (O_2228,N_19511,N_18563);
and UO_2229 (O_2229,N_19142,N_19620);
or UO_2230 (O_2230,N_19812,N_18429);
nand UO_2231 (O_2231,N_19243,N_18430);
nand UO_2232 (O_2232,N_19033,N_18826);
or UO_2233 (O_2233,N_18484,N_19267);
nand UO_2234 (O_2234,N_18018,N_19134);
and UO_2235 (O_2235,N_18987,N_18730);
or UO_2236 (O_2236,N_19604,N_18645);
nor UO_2237 (O_2237,N_19613,N_19890);
and UO_2238 (O_2238,N_18610,N_19280);
or UO_2239 (O_2239,N_18938,N_19902);
nand UO_2240 (O_2240,N_19319,N_19922);
or UO_2241 (O_2241,N_19650,N_18493);
or UO_2242 (O_2242,N_19150,N_18562);
and UO_2243 (O_2243,N_18675,N_18888);
or UO_2244 (O_2244,N_18512,N_19679);
and UO_2245 (O_2245,N_19646,N_19342);
and UO_2246 (O_2246,N_19364,N_19657);
and UO_2247 (O_2247,N_18642,N_18717);
and UO_2248 (O_2248,N_18455,N_18526);
or UO_2249 (O_2249,N_18399,N_19426);
and UO_2250 (O_2250,N_18318,N_18795);
nor UO_2251 (O_2251,N_19613,N_19702);
and UO_2252 (O_2252,N_18613,N_18642);
or UO_2253 (O_2253,N_19132,N_19098);
nand UO_2254 (O_2254,N_19675,N_18856);
nor UO_2255 (O_2255,N_19316,N_18049);
or UO_2256 (O_2256,N_18826,N_18866);
nand UO_2257 (O_2257,N_18501,N_19870);
nand UO_2258 (O_2258,N_19081,N_18697);
or UO_2259 (O_2259,N_19536,N_19091);
nor UO_2260 (O_2260,N_19002,N_18294);
or UO_2261 (O_2261,N_18430,N_18556);
nand UO_2262 (O_2262,N_18112,N_18205);
nor UO_2263 (O_2263,N_19996,N_19515);
or UO_2264 (O_2264,N_19443,N_18550);
nor UO_2265 (O_2265,N_19841,N_18076);
or UO_2266 (O_2266,N_19455,N_18072);
nand UO_2267 (O_2267,N_19948,N_19195);
or UO_2268 (O_2268,N_19334,N_19933);
and UO_2269 (O_2269,N_18724,N_19236);
nor UO_2270 (O_2270,N_19392,N_18150);
and UO_2271 (O_2271,N_19020,N_18255);
and UO_2272 (O_2272,N_19500,N_19752);
xnor UO_2273 (O_2273,N_18393,N_18695);
and UO_2274 (O_2274,N_19784,N_19714);
and UO_2275 (O_2275,N_19014,N_19603);
or UO_2276 (O_2276,N_19111,N_19203);
nand UO_2277 (O_2277,N_18283,N_19690);
nor UO_2278 (O_2278,N_19765,N_19418);
nor UO_2279 (O_2279,N_18920,N_18144);
or UO_2280 (O_2280,N_19123,N_19149);
or UO_2281 (O_2281,N_18507,N_19732);
nand UO_2282 (O_2282,N_19841,N_18200);
nand UO_2283 (O_2283,N_19163,N_18699);
nor UO_2284 (O_2284,N_18515,N_18429);
nand UO_2285 (O_2285,N_19395,N_18206);
nand UO_2286 (O_2286,N_19131,N_19861);
and UO_2287 (O_2287,N_19635,N_18660);
and UO_2288 (O_2288,N_18607,N_18857);
or UO_2289 (O_2289,N_19743,N_19571);
or UO_2290 (O_2290,N_18238,N_18118);
xnor UO_2291 (O_2291,N_19327,N_19061);
nor UO_2292 (O_2292,N_19762,N_18959);
nand UO_2293 (O_2293,N_19991,N_18103);
and UO_2294 (O_2294,N_19269,N_18027);
nor UO_2295 (O_2295,N_19291,N_19927);
or UO_2296 (O_2296,N_19387,N_19430);
xnor UO_2297 (O_2297,N_18339,N_19157);
and UO_2298 (O_2298,N_19877,N_18980);
nand UO_2299 (O_2299,N_19653,N_18081);
nand UO_2300 (O_2300,N_18927,N_18711);
xnor UO_2301 (O_2301,N_18319,N_19219);
nand UO_2302 (O_2302,N_18974,N_19072);
and UO_2303 (O_2303,N_19264,N_19567);
nand UO_2304 (O_2304,N_19338,N_18751);
and UO_2305 (O_2305,N_18283,N_18207);
nor UO_2306 (O_2306,N_18344,N_19187);
nor UO_2307 (O_2307,N_19252,N_18359);
nand UO_2308 (O_2308,N_19937,N_18918);
and UO_2309 (O_2309,N_18502,N_18018);
nand UO_2310 (O_2310,N_18523,N_19739);
nor UO_2311 (O_2311,N_18499,N_19556);
xnor UO_2312 (O_2312,N_19879,N_18146);
and UO_2313 (O_2313,N_18499,N_19503);
xor UO_2314 (O_2314,N_19835,N_18004);
and UO_2315 (O_2315,N_19164,N_19769);
nor UO_2316 (O_2316,N_18086,N_19607);
or UO_2317 (O_2317,N_19179,N_19559);
or UO_2318 (O_2318,N_18098,N_19565);
nor UO_2319 (O_2319,N_18451,N_18590);
or UO_2320 (O_2320,N_18309,N_19242);
and UO_2321 (O_2321,N_19166,N_19137);
and UO_2322 (O_2322,N_18899,N_19042);
or UO_2323 (O_2323,N_19037,N_19345);
and UO_2324 (O_2324,N_18360,N_19514);
nor UO_2325 (O_2325,N_19559,N_19634);
and UO_2326 (O_2326,N_19346,N_19185);
nand UO_2327 (O_2327,N_19505,N_18664);
or UO_2328 (O_2328,N_18820,N_18427);
nand UO_2329 (O_2329,N_19527,N_19780);
nor UO_2330 (O_2330,N_19917,N_18969);
nand UO_2331 (O_2331,N_18767,N_19504);
or UO_2332 (O_2332,N_18059,N_19799);
nor UO_2333 (O_2333,N_18049,N_19733);
xor UO_2334 (O_2334,N_18926,N_19875);
or UO_2335 (O_2335,N_19848,N_18059);
or UO_2336 (O_2336,N_18333,N_19787);
and UO_2337 (O_2337,N_19322,N_19119);
nor UO_2338 (O_2338,N_18795,N_19181);
or UO_2339 (O_2339,N_18129,N_19593);
nand UO_2340 (O_2340,N_19848,N_18921);
nor UO_2341 (O_2341,N_18851,N_18882);
or UO_2342 (O_2342,N_19979,N_18038);
and UO_2343 (O_2343,N_19420,N_18420);
or UO_2344 (O_2344,N_18330,N_18109);
or UO_2345 (O_2345,N_19632,N_19470);
nor UO_2346 (O_2346,N_18064,N_18860);
or UO_2347 (O_2347,N_19748,N_18315);
nor UO_2348 (O_2348,N_18457,N_18087);
nor UO_2349 (O_2349,N_18133,N_19878);
and UO_2350 (O_2350,N_18238,N_19136);
nor UO_2351 (O_2351,N_18815,N_18040);
or UO_2352 (O_2352,N_19251,N_19442);
nor UO_2353 (O_2353,N_18207,N_18175);
nor UO_2354 (O_2354,N_19688,N_19120);
and UO_2355 (O_2355,N_18656,N_19701);
nor UO_2356 (O_2356,N_19216,N_18270);
or UO_2357 (O_2357,N_18394,N_18803);
nand UO_2358 (O_2358,N_18117,N_18988);
nand UO_2359 (O_2359,N_18135,N_18173);
nor UO_2360 (O_2360,N_18683,N_19415);
xnor UO_2361 (O_2361,N_19956,N_18850);
nor UO_2362 (O_2362,N_18308,N_18682);
nor UO_2363 (O_2363,N_18297,N_19349);
nor UO_2364 (O_2364,N_18373,N_18720);
nand UO_2365 (O_2365,N_18047,N_19543);
or UO_2366 (O_2366,N_19487,N_18506);
or UO_2367 (O_2367,N_19944,N_18103);
nor UO_2368 (O_2368,N_18133,N_19282);
nor UO_2369 (O_2369,N_19581,N_19745);
and UO_2370 (O_2370,N_18066,N_19463);
and UO_2371 (O_2371,N_18777,N_18892);
and UO_2372 (O_2372,N_18213,N_18209);
or UO_2373 (O_2373,N_19600,N_19429);
and UO_2374 (O_2374,N_18703,N_19814);
or UO_2375 (O_2375,N_18495,N_19536);
nor UO_2376 (O_2376,N_19126,N_18987);
or UO_2377 (O_2377,N_19863,N_18095);
or UO_2378 (O_2378,N_18463,N_18435);
xnor UO_2379 (O_2379,N_18938,N_19155);
and UO_2380 (O_2380,N_18425,N_18802);
and UO_2381 (O_2381,N_18826,N_19525);
nor UO_2382 (O_2382,N_18728,N_19146);
and UO_2383 (O_2383,N_18766,N_19728);
nand UO_2384 (O_2384,N_18560,N_18461);
and UO_2385 (O_2385,N_19061,N_18307);
and UO_2386 (O_2386,N_19339,N_19148);
or UO_2387 (O_2387,N_19031,N_19281);
nor UO_2388 (O_2388,N_18941,N_18570);
and UO_2389 (O_2389,N_18013,N_19590);
and UO_2390 (O_2390,N_18210,N_19695);
nand UO_2391 (O_2391,N_18754,N_19674);
nor UO_2392 (O_2392,N_19587,N_19148);
or UO_2393 (O_2393,N_18292,N_19340);
nand UO_2394 (O_2394,N_18302,N_18901);
nor UO_2395 (O_2395,N_18696,N_19970);
and UO_2396 (O_2396,N_19518,N_19257);
and UO_2397 (O_2397,N_19958,N_19973);
and UO_2398 (O_2398,N_19131,N_18678);
or UO_2399 (O_2399,N_18453,N_19324);
or UO_2400 (O_2400,N_19334,N_19765);
nand UO_2401 (O_2401,N_19855,N_19611);
or UO_2402 (O_2402,N_18262,N_18916);
and UO_2403 (O_2403,N_18111,N_18193);
or UO_2404 (O_2404,N_19171,N_18655);
xnor UO_2405 (O_2405,N_18255,N_19941);
nor UO_2406 (O_2406,N_18298,N_19025);
nor UO_2407 (O_2407,N_18673,N_19519);
nand UO_2408 (O_2408,N_18843,N_19245);
nand UO_2409 (O_2409,N_18192,N_18649);
xnor UO_2410 (O_2410,N_19576,N_18991);
and UO_2411 (O_2411,N_19297,N_18266);
nand UO_2412 (O_2412,N_19325,N_19526);
nand UO_2413 (O_2413,N_19330,N_19008);
or UO_2414 (O_2414,N_18444,N_19714);
and UO_2415 (O_2415,N_18675,N_18687);
nor UO_2416 (O_2416,N_19013,N_19265);
and UO_2417 (O_2417,N_18875,N_19600);
nor UO_2418 (O_2418,N_19781,N_19278);
xor UO_2419 (O_2419,N_19359,N_18310);
nand UO_2420 (O_2420,N_18773,N_19880);
and UO_2421 (O_2421,N_19747,N_19975);
and UO_2422 (O_2422,N_18393,N_18142);
xor UO_2423 (O_2423,N_18748,N_18678);
nor UO_2424 (O_2424,N_19463,N_19147);
and UO_2425 (O_2425,N_19240,N_19940);
or UO_2426 (O_2426,N_18536,N_19585);
nor UO_2427 (O_2427,N_18645,N_18281);
nand UO_2428 (O_2428,N_18234,N_19834);
or UO_2429 (O_2429,N_18966,N_18956);
or UO_2430 (O_2430,N_19685,N_18302);
or UO_2431 (O_2431,N_18998,N_18369);
nor UO_2432 (O_2432,N_19865,N_18584);
nand UO_2433 (O_2433,N_19651,N_18937);
or UO_2434 (O_2434,N_18793,N_18990);
or UO_2435 (O_2435,N_19351,N_18451);
nor UO_2436 (O_2436,N_19644,N_18243);
nor UO_2437 (O_2437,N_18960,N_19388);
nand UO_2438 (O_2438,N_18961,N_18836);
nor UO_2439 (O_2439,N_19113,N_19139);
and UO_2440 (O_2440,N_18457,N_18749);
and UO_2441 (O_2441,N_18095,N_19925);
nor UO_2442 (O_2442,N_19335,N_18878);
and UO_2443 (O_2443,N_19266,N_19520);
nor UO_2444 (O_2444,N_18559,N_18398);
nor UO_2445 (O_2445,N_18541,N_18913);
and UO_2446 (O_2446,N_18086,N_18541);
or UO_2447 (O_2447,N_19178,N_18144);
and UO_2448 (O_2448,N_18791,N_18359);
or UO_2449 (O_2449,N_18410,N_18358);
nor UO_2450 (O_2450,N_19293,N_18872);
nand UO_2451 (O_2451,N_19181,N_19176);
nor UO_2452 (O_2452,N_18796,N_18851);
nand UO_2453 (O_2453,N_19639,N_18242);
nor UO_2454 (O_2454,N_19811,N_18012);
and UO_2455 (O_2455,N_18012,N_19992);
and UO_2456 (O_2456,N_18759,N_19980);
or UO_2457 (O_2457,N_18455,N_18077);
nand UO_2458 (O_2458,N_18861,N_19278);
nand UO_2459 (O_2459,N_18235,N_19098);
and UO_2460 (O_2460,N_19286,N_19107);
nand UO_2461 (O_2461,N_18958,N_18414);
nor UO_2462 (O_2462,N_19444,N_18985);
nand UO_2463 (O_2463,N_18614,N_18022);
or UO_2464 (O_2464,N_19650,N_19722);
or UO_2465 (O_2465,N_18480,N_18828);
xnor UO_2466 (O_2466,N_19165,N_18011);
or UO_2467 (O_2467,N_18123,N_18064);
nor UO_2468 (O_2468,N_18916,N_19947);
and UO_2469 (O_2469,N_19202,N_18487);
or UO_2470 (O_2470,N_18856,N_18660);
nor UO_2471 (O_2471,N_19729,N_19136);
nand UO_2472 (O_2472,N_19652,N_18998);
and UO_2473 (O_2473,N_18090,N_18673);
and UO_2474 (O_2474,N_18075,N_19056);
and UO_2475 (O_2475,N_19943,N_19066);
or UO_2476 (O_2476,N_18230,N_18052);
and UO_2477 (O_2477,N_19650,N_18855);
nor UO_2478 (O_2478,N_18554,N_18126);
or UO_2479 (O_2479,N_18277,N_18243);
nor UO_2480 (O_2480,N_19027,N_18846);
and UO_2481 (O_2481,N_19109,N_19627);
nor UO_2482 (O_2482,N_19553,N_19659);
and UO_2483 (O_2483,N_18734,N_19288);
or UO_2484 (O_2484,N_18688,N_19303);
and UO_2485 (O_2485,N_18614,N_19052);
and UO_2486 (O_2486,N_18140,N_18811);
nor UO_2487 (O_2487,N_19065,N_18259);
or UO_2488 (O_2488,N_19944,N_19034);
xor UO_2489 (O_2489,N_19178,N_19855);
nand UO_2490 (O_2490,N_18586,N_18271);
and UO_2491 (O_2491,N_19964,N_18640);
or UO_2492 (O_2492,N_18104,N_18509);
nand UO_2493 (O_2493,N_18218,N_18123);
or UO_2494 (O_2494,N_18377,N_19561);
nor UO_2495 (O_2495,N_19249,N_19618);
nand UO_2496 (O_2496,N_19463,N_18428);
and UO_2497 (O_2497,N_18107,N_19706);
nor UO_2498 (O_2498,N_19948,N_18125);
and UO_2499 (O_2499,N_18918,N_19563);
endmodule