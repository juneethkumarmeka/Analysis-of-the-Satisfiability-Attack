module basic_3000_30000_3500_6_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
and U0 (N_0,In_378,In_2377);
and U1 (N_1,In_193,In_2558);
or U2 (N_2,In_670,In_837);
nor U3 (N_3,In_793,In_1745);
or U4 (N_4,In_778,In_1563);
and U5 (N_5,In_106,In_1165);
nor U6 (N_6,In_1914,In_1013);
or U7 (N_7,In_506,In_2840);
nand U8 (N_8,In_1225,In_886);
xor U9 (N_9,In_2704,In_1111);
and U10 (N_10,In_2506,In_121);
nand U11 (N_11,In_1016,In_2887);
nand U12 (N_12,In_100,In_57);
or U13 (N_13,In_2318,In_437);
nor U14 (N_14,In_810,In_842);
or U15 (N_15,In_2729,In_2111);
nand U16 (N_16,In_2742,In_1180);
or U17 (N_17,In_690,In_1654);
nand U18 (N_18,In_538,In_13);
or U19 (N_19,In_333,In_1542);
or U20 (N_20,In_1200,In_1717);
nor U21 (N_21,In_1272,In_631);
nor U22 (N_22,In_327,In_2096);
nor U23 (N_23,In_1499,In_1515);
nand U24 (N_24,In_801,In_2267);
nand U25 (N_25,In_2329,In_2241);
or U26 (N_26,In_1065,In_963);
or U27 (N_27,In_2387,In_2850);
nand U28 (N_28,In_2958,In_1678);
nor U29 (N_29,In_1084,In_1374);
or U30 (N_30,In_526,In_1436);
nor U31 (N_31,In_427,In_453);
or U32 (N_32,In_621,In_1904);
and U33 (N_33,In_2295,In_1158);
nor U34 (N_34,In_668,In_2595);
and U35 (N_35,In_1629,In_940);
and U36 (N_36,In_2332,In_1591);
nand U37 (N_37,In_562,In_2327);
nor U38 (N_38,In_2409,In_527);
and U39 (N_39,In_2259,In_2581);
nor U40 (N_40,In_779,In_658);
or U41 (N_41,In_1283,In_183);
or U42 (N_42,In_235,In_2619);
or U43 (N_43,In_698,In_2445);
xnor U44 (N_44,In_2817,In_2833);
nor U45 (N_45,In_2779,In_2977);
or U46 (N_46,In_2083,In_2510);
nand U47 (N_47,In_1316,In_1141);
xor U48 (N_48,In_1514,In_1523);
xor U49 (N_49,In_1752,In_2163);
nand U50 (N_50,In_1834,In_175);
nand U51 (N_51,In_962,In_1659);
and U52 (N_52,In_1387,In_1566);
nor U53 (N_53,In_1781,In_2518);
nand U54 (N_54,In_1192,In_191);
or U55 (N_55,In_696,In_1427);
or U56 (N_56,In_870,In_2678);
xnor U57 (N_57,In_1991,In_802);
or U58 (N_58,In_2413,In_90);
xor U59 (N_59,In_326,In_1707);
xor U60 (N_60,In_1056,In_1277);
nand U61 (N_61,In_1619,In_62);
or U62 (N_62,In_917,In_1811);
nor U63 (N_63,In_70,In_2194);
and U64 (N_64,In_1950,In_117);
or U65 (N_65,In_888,In_284);
or U66 (N_66,In_401,In_663);
nor U67 (N_67,In_914,In_1400);
xor U68 (N_68,In_313,In_923);
nor U69 (N_69,In_2179,In_1160);
xnor U70 (N_70,In_1430,In_2247);
nor U71 (N_71,In_721,In_2443);
nand U72 (N_72,In_2156,In_375);
nand U73 (N_73,In_1869,In_2546);
nand U74 (N_74,In_1250,In_1244);
or U75 (N_75,In_69,In_39);
nand U76 (N_76,In_2109,In_274);
or U77 (N_77,In_32,In_283);
nor U78 (N_78,In_1445,In_282);
nor U79 (N_79,In_820,In_1600);
nor U80 (N_80,In_2098,In_1024);
nand U81 (N_81,In_1575,In_2561);
nand U82 (N_82,In_1741,In_1094);
nor U83 (N_83,In_881,In_2356);
nand U84 (N_84,In_2079,In_1519);
or U85 (N_85,In_2401,In_2000);
or U86 (N_86,In_776,In_474);
and U87 (N_87,In_404,In_2522);
nor U88 (N_88,In_347,In_549);
nor U89 (N_89,In_1044,In_760);
and U90 (N_90,In_1130,In_2812);
or U91 (N_91,In_1458,In_2822);
nor U92 (N_92,In_1486,In_171);
nand U93 (N_93,In_2408,In_2759);
nand U94 (N_94,In_2040,In_1011);
or U95 (N_95,In_1794,In_1832);
nor U96 (N_96,In_2298,In_364);
nand U97 (N_97,In_352,In_1596);
nor U98 (N_98,In_869,In_1046);
or U99 (N_99,In_1916,In_74);
or U100 (N_100,In_1399,In_2544);
nor U101 (N_101,In_699,In_531);
nor U102 (N_102,In_2069,In_2149);
nand U103 (N_103,In_1997,In_2775);
nor U104 (N_104,In_1749,In_151);
nor U105 (N_105,In_2613,In_392);
or U106 (N_106,In_596,In_119);
xor U107 (N_107,In_942,In_1410);
or U108 (N_108,In_684,In_1122);
or U109 (N_109,In_2235,In_2285);
nor U110 (N_110,In_357,In_1977);
nand U111 (N_111,In_1908,In_2893);
nand U112 (N_112,In_1354,In_2154);
nand U113 (N_113,In_635,In_706);
or U114 (N_114,In_1716,In_2867);
xnor U115 (N_115,In_2453,In_1304);
and U116 (N_116,In_2207,In_983);
or U117 (N_117,In_2392,In_2080);
nor U118 (N_118,In_542,In_1669);
nor U119 (N_119,In_348,In_744);
or U120 (N_120,In_467,In_1995);
nor U121 (N_121,In_2450,In_918);
and U122 (N_122,In_92,In_665);
xnor U123 (N_123,In_1763,In_834);
nand U124 (N_124,In_2916,In_1552);
and U125 (N_125,In_1118,In_1818);
nand U126 (N_126,In_1714,In_1090);
or U127 (N_127,In_2287,In_1784);
nand U128 (N_128,In_2343,In_297);
and U129 (N_129,In_2168,In_500);
nand U130 (N_130,In_1392,In_2672);
or U131 (N_131,In_2664,In_1762);
or U132 (N_132,In_1696,In_2917);
nand U133 (N_133,In_594,In_2342);
xor U134 (N_134,In_1797,In_145);
and U135 (N_135,In_2752,In_494);
and U136 (N_136,In_1722,In_2441);
or U137 (N_137,In_1379,In_2844);
xnor U138 (N_138,In_464,In_1537);
or U139 (N_139,In_2010,In_734);
xnor U140 (N_140,In_2283,In_125);
nand U141 (N_141,In_2877,In_109);
nand U142 (N_142,In_1107,In_215);
nand U143 (N_143,In_2810,In_1527);
xnor U144 (N_144,In_152,In_536);
and U145 (N_145,In_1189,In_391);
nand U146 (N_146,In_1670,In_1814);
nand U147 (N_147,In_2592,In_1455);
nor U148 (N_148,In_196,In_1822);
xnor U149 (N_149,In_28,In_525);
nor U150 (N_150,In_2036,In_1069);
nand U151 (N_151,In_1,In_1885);
nor U152 (N_152,In_20,In_1498);
nor U153 (N_153,In_372,In_2918);
nand U154 (N_154,In_476,In_1932);
or U155 (N_155,In_1650,In_764);
and U156 (N_156,In_169,In_156);
nor U157 (N_157,In_2766,In_2007);
nor U158 (N_158,In_1196,In_2731);
nor U159 (N_159,In_2262,In_2717);
nor U160 (N_160,In_896,In_2559);
xor U161 (N_161,In_1859,In_73);
or U162 (N_162,In_2881,In_2525);
nand U163 (N_163,In_2030,In_2202);
xnor U164 (N_164,In_1391,In_2999);
and U165 (N_165,In_2464,In_311);
nor U166 (N_166,In_578,In_2824);
and U167 (N_167,In_2683,In_2136);
and U168 (N_168,In_2728,In_2276);
nor U169 (N_169,In_2665,In_2716);
nor U170 (N_170,In_2784,In_131);
or U171 (N_171,In_2903,In_898);
or U172 (N_172,In_529,In_2930);
nand U173 (N_173,In_632,In_651);
nand U174 (N_174,In_2987,In_419);
or U175 (N_175,In_1831,In_2151);
or U176 (N_176,In_1906,In_724);
and U177 (N_177,In_1689,In_2735);
and U178 (N_178,In_996,In_1723);
xor U179 (N_179,In_2352,In_2077);
nand U180 (N_180,In_345,In_2300);
and U181 (N_181,In_1078,In_239);
xor U182 (N_182,In_2739,In_1656);
and U183 (N_183,In_1414,In_831);
and U184 (N_184,In_1367,In_103);
or U185 (N_185,In_1861,In_1481);
nand U186 (N_186,In_960,In_210);
and U187 (N_187,In_16,In_1351);
or U188 (N_188,In_505,In_1027);
xor U189 (N_189,In_2004,In_1381);
nor U190 (N_190,In_1688,In_2796);
xnor U191 (N_191,In_1406,In_2442);
nand U192 (N_192,In_2153,In_563);
xnor U193 (N_193,In_315,In_2745);
and U194 (N_194,In_2684,In_2063);
and U195 (N_195,In_1708,In_79);
nand U196 (N_196,In_934,In_901);
nand U197 (N_197,In_2690,In_250);
xnor U198 (N_198,In_1518,In_1594);
nor U199 (N_199,In_507,In_2639);
and U200 (N_200,In_2033,In_2384);
nand U201 (N_201,In_1418,In_807);
or U202 (N_202,In_67,In_438);
nor U203 (N_203,In_1910,In_2424);
xnor U204 (N_204,In_452,In_1203);
nor U205 (N_205,In_2048,In_784);
nor U206 (N_206,In_747,In_2847);
nor U207 (N_207,In_1170,In_2865);
or U208 (N_208,In_2886,In_2514);
or U209 (N_209,In_451,In_2491);
nand U210 (N_210,In_133,In_2702);
and U211 (N_211,In_1630,In_875);
nor U212 (N_212,In_2406,In_2128);
or U213 (N_213,In_1676,In_848);
nor U214 (N_214,In_2334,In_1247);
and U215 (N_215,In_1735,In_2148);
nand U216 (N_216,In_2931,In_1778);
nor U217 (N_217,In_2860,In_600);
nor U218 (N_218,In_1234,In_2452);
or U219 (N_219,In_1962,In_715);
and U220 (N_220,In_1655,In_2949);
nor U221 (N_221,In_31,In_324);
xor U222 (N_222,In_1242,In_136);
or U223 (N_223,In_612,In_1388);
nor U224 (N_224,In_2538,In_754);
and U225 (N_225,In_1288,In_2302);
nor U226 (N_226,In_1759,In_2046);
and U227 (N_227,In_1363,In_1557);
nor U228 (N_228,In_2434,In_1903);
nand U229 (N_229,In_927,In_1724);
and U230 (N_230,In_1750,In_2573);
and U231 (N_231,In_1467,In_2531);
nand U232 (N_232,In_2969,In_157);
or U233 (N_233,In_2505,In_1251);
nor U234 (N_234,In_54,In_1441);
and U235 (N_235,In_2551,In_2269);
or U236 (N_236,In_2853,In_1053);
xor U237 (N_237,In_617,In_1560);
nand U238 (N_238,In_504,In_1732);
or U239 (N_239,In_1266,In_2189);
nand U240 (N_240,In_1343,In_2806);
nor U241 (N_241,In_442,In_94);
nand U242 (N_242,In_1621,In_654);
nand U243 (N_243,In_84,In_2997);
nand U244 (N_244,In_2839,In_2448);
or U245 (N_245,In_2092,In_2962);
nand U246 (N_246,In_388,In_445);
or U247 (N_247,In_473,In_214);
nor U248 (N_248,In_1555,In_1975);
xor U249 (N_249,In_2520,In_178);
nor U250 (N_250,In_1758,In_1808);
nand U251 (N_251,In_1968,In_532);
nand U252 (N_252,In_66,In_303);
and U253 (N_253,In_255,In_742);
xor U254 (N_254,In_240,In_769);
nand U255 (N_255,In_1915,In_2773);
nand U256 (N_256,In_607,In_711);
nor U257 (N_257,In_271,In_325);
nor U258 (N_258,In_371,In_1772);
nor U259 (N_259,In_1726,In_1711);
or U260 (N_260,In_1093,In_2072);
nor U261 (N_261,In_141,In_2980);
nand U262 (N_262,In_547,In_633);
nand U263 (N_263,In_1699,In_2908);
or U264 (N_264,In_1156,In_2625);
and U265 (N_265,In_1145,In_2420);
nand U266 (N_266,In_17,In_314);
nand U267 (N_267,In_259,In_338);
and U268 (N_268,In_1369,In_503);
nand U269 (N_269,In_995,In_1095);
nor U270 (N_270,In_1018,In_1401);
or U271 (N_271,In_429,In_195);
nand U272 (N_272,In_534,In_2305);
or U273 (N_273,In_1012,In_1980);
xor U274 (N_274,In_2515,In_281);
nor U275 (N_275,In_789,In_2826);
and U276 (N_276,In_2959,In_154);
nor U277 (N_277,In_1548,In_1287);
and U278 (N_278,In_548,In_1827);
xnor U279 (N_279,In_1175,In_605);
nand U280 (N_280,In_2624,In_2301);
and U281 (N_281,In_1059,In_30);
or U282 (N_282,In_301,In_1826);
nand U283 (N_283,In_2017,In_2682);
or U284 (N_284,In_1474,In_546);
or U285 (N_285,In_277,In_2929);
nor U286 (N_286,In_691,In_973);
or U287 (N_287,In_2360,In_209);
nand U288 (N_288,In_1309,In_863);
xnor U289 (N_289,In_2854,In_107);
and U290 (N_290,In_188,In_2873);
nor U291 (N_291,In_2073,In_2379);
nand U292 (N_292,In_1588,In_762);
nand U293 (N_293,In_2834,In_1934);
nand U294 (N_294,In_1993,In_305);
nand U295 (N_295,In_2855,In_2020);
or U296 (N_296,In_2937,In_2229);
nor U297 (N_297,In_367,In_2757);
and U298 (N_298,In_1589,In_2673);
and U299 (N_299,In_160,In_459);
nand U300 (N_300,In_1503,In_774);
xnor U301 (N_301,In_2225,In_406);
nand U302 (N_302,In_2463,In_513);
or U303 (N_303,In_1380,In_1804);
nand U304 (N_304,In_2339,In_2133);
nand U305 (N_305,In_2688,In_1449);
and U306 (N_306,In_626,In_2169);
and U307 (N_307,In_1315,In_435);
nand U308 (N_308,In_614,In_220);
or U309 (N_309,In_83,In_921);
nor U310 (N_310,In_2082,In_1155);
or U311 (N_311,In_269,In_1782);
and U312 (N_312,In_2906,In_2642);
nand U313 (N_313,In_1883,In_713);
nand U314 (N_314,In_1029,In_1477);
nand U315 (N_315,In_2347,In_1256);
nand U316 (N_316,In_134,In_49);
nor U317 (N_317,In_29,In_867);
nor U318 (N_318,In_1489,In_2950);
and U319 (N_319,In_2274,In_186);
or U320 (N_320,In_2388,In_1751);
nor U321 (N_321,In_821,In_2957);
or U322 (N_322,In_1798,In_2280);
nor U323 (N_323,In_1715,In_2963);
nor U324 (N_324,In_1360,In_181);
and U325 (N_325,In_892,In_2412);
and U326 (N_326,In_1417,In_756);
or U327 (N_327,In_2393,In_2830);
nor U328 (N_328,In_2076,In_709);
nor U329 (N_329,In_1033,In_2602);
nor U330 (N_330,In_1108,In_335);
nand U331 (N_331,In_1528,In_611);
or U332 (N_332,In_829,In_714);
or U333 (N_333,In_1395,In_2206);
and U334 (N_334,In_471,In_2024);
and U335 (N_335,In_1598,In_2674);
nand U336 (N_336,In_229,In_1216);
or U337 (N_337,In_2053,In_480);
and U338 (N_338,In_738,In_1949);
nand U339 (N_339,In_965,In_1599);
and U340 (N_340,In_948,In_428);
nor U341 (N_341,In_1157,In_48);
nand U342 (N_342,In_2284,In_618);
nor U343 (N_343,In_2667,In_1963);
and U344 (N_344,In_561,In_1021);
nor U345 (N_345,In_2547,In_2576);
or U346 (N_346,In_272,In_140);
xnor U347 (N_347,In_2669,In_1839);
or U348 (N_348,In_415,In_556);
nand U349 (N_349,In_2121,In_1545);
or U350 (N_350,In_86,In_757);
nand U351 (N_351,In_1790,In_2219);
nor U352 (N_352,In_405,In_2772);
or U353 (N_353,In_18,In_1181);
xnor U354 (N_354,In_2363,In_1341);
nand U355 (N_355,In_2939,In_828);
nand U356 (N_356,In_1681,In_2701);
or U357 (N_357,In_2019,In_827);
nand U358 (N_358,In_2549,In_653);
or U359 (N_359,In_2116,In_1705);
nand U360 (N_360,In_2042,In_2099);
nand U361 (N_361,In_1526,In_153);
xor U362 (N_362,In_2774,In_887);
or U363 (N_363,In_499,In_2878);
or U364 (N_364,In_523,In_76);
nand U365 (N_365,In_1397,In_2323);
or U366 (N_366,In_1960,In_727);
or U367 (N_367,In_2045,In_2135);
or U368 (N_368,In_2216,In_1362);
or U369 (N_369,In_839,In_2988);
and U370 (N_370,In_298,In_2956);
and U371 (N_371,In_2923,In_1734);
nand U372 (N_372,In_2970,In_2186);
and U373 (N_373,In_2719,In_1052);
nand U374 (N_374,In_1258,In_1923);
and U375 (N_375,In_1768,In_859);
nor U376 (N_376,In_957,In_2802);
xor U377 (N_377,In_2440,In_1439);
or U378 (N_378,In_1821,In_1359);
or U379 (N_379,In_920,In_1253);
nand U380 (N_380,In_1941,In_1330);
or U381 (N_381,In_75,In_337);
or U382 (N_382,In_2814,In_1985);
or U383 (N_383,In_2037,In_1692);
nor U384 (N_384,In_2791,In_985);
and U385 (N_385,In_2800,In_2105);
and U386 (N_386,In_819,In_64);
or U387 (N_387,In_1593,In_2627);
nand U388 (N_388,In_2859,In_567);
nand U389 (N_389,In_2748,In_2730);
nand U390 (N_390,In_1124,In_959);
and U391 (N_391,In_1269,In_999);
nor U392 (N_392,In_2540,In_798);
and U393 (N_393,In_2655,In_123);
or U394 (N_394,In_1132,In_279);
and U395 (N_395,In_377,In_443);
or U396 (N_396,In_1082,In_1000);
or U397 (N_397,In_1119,In_2516);
nand U398 (N_398,In_683,In_2606);
or U399 (N_399,In_1796,In_836);
or U400 (N_400,In_2102,In_584);
and U401 (N_401,In_1473,In_2785);
and U402 (N_402,In_987,In_2885);
nand U403 (N_403,In_2499,In_1907);
nand U404 (N_404,In_340,In_430);
nand U405 (N_405,In_516,In_1882);
nand U406 (N_406,In_1553,In_382);
nor U407 (N_407,In_2575,In_180);
or U408 (N_408,In_2433,In_2473);
nand U409 (N_409,In_890,In_1459);
nand U410 (N_410,In_813,In_1658);
nand U411 (N_411,In_1178,In_2761);
or U412 (N_412,In_1435,In_2178);
and U413 (N_413,In_550,In_219);
nand U414 (N_414,In_1389,In_2150);
nand U415 (N_415,In_22,In_1565);
nand U416 (N_416,In_2691,In_1986);
and U417 (N_417,In_1008,In_1100);
or U418 (N_418,In_60,In_483);
or U419 (N_419,In_1215,In_2103);
xor U420 (N_420,In_1856,In_42);
and U421 (N_421,In_1973,In_816);
nand U422 (N_422,In_2776,In_455);
nor U423 (N_423,In_558,In_1767);
and U424 (N_424,In_1294,In_1125);
or U425 (N_425,In_1134,In_2203);
xnor U426 (N_426,In_2770,In_1524);
nand U427 (N_427,In_399,In_497);
nand U428 (N_428,In_937,In_2373);
and U429 (N_429,In_2411,In_393);
or U430 (N_430,In_2058,In_2948);
nor U431 (N_431,In_2699,In_1701);
nor U432 (N_432,In_2967,In_1002);
or U433 (N_433,In_521,In_2979);
nor U434 (N_434,In_216,In_1644);
or U435 (N_435,In_1313,In_1642);
nor U436 (N_436,In_588,In_1660);
and U437 (N_437,In_1836,In_2749);
nand U438 (N_438,In_2933,In_1135);
and U439 (N_439,In_1695,In_2951);
and U440 (N_440,In_1206,In_1466);
or U441 (N_441,In_840,In_285);
and U442 (N_442,In_2804,In_1079);
or U443 (N_443,In_189,In_788);
nand U444 (N_444,In_369,In_2404);
xor U445 (N_445,In_2849,In_379);
nor U446 (N_446,In_1501,In_876);
nand U447 (N_447,In_2539,In_1857);
nor U448 (N_448,In_2474,In_1533);
nand U449 (N_449,In_2620,In_23);
or U450 (N_450,In_2112,In_412);
xnor U451 (N_451,In_2454,In_939);
or U452 (N_452,In_1721,In_1824);
xnor U453 (N_453,In_1844,In_2501);
nor U454 (N_454,In_2056,In_582);
and U455 (N_455,In_2255,In_458);
and U456 (N_456,In_852,In_394);
and U457 (N_457,In_2243,In_2793);
or U458 (N_458,In_2656,In_318);
or U459 (N_459,In_1951,In_2155);
xnor U460 (N_460,In_2369,In_687);
or U461 (N_461,In_1979,In_708);
nor U462 (N_462,In_1933,In_954);
or U463 (N_463,In_1372,In_291);
or U464 (N_464,In_2944,In_2626);
or U465 (N_465,In_1366,In_2011);
nand U466 (N_466,In_1030,In_2245);
nand U467 (N_467,In_2580,In_2126);
nor U468 (N_468,In_2823,In_1273);
nand U469 (N_469,In_481,In_830);
nand U470 (N_470,In_2199,In_252);
and U471 (N_471,In_2909,In_1195);
and U472 (N_472,In_1789,In_675);
nand U473 (N_473,In_113,In_2726);
nand U474 (N_474,In_595,In_2789);
nor U475 (N_475,In_1274,In_1218);
nor U476 (N_476,In_931,In_1227);
nand U477 (N_477,In_2237,In_2687);
nor U478 (N_478,In_1162,In_718);
or U479 (N_479,In_1081,In_2264);
nand U480 (N_480,In_1590,In_2158);
nor U481 (N_481,In_469,In_2059);
and U482 (N_482,In_2394,In_599);
nand U483 (N_483,In_763,In_2480);
or U484 (N_484,In_1248,In_2012);
nor U485 (N_485,In_2500,In_253);
xnor U486 (N_486,In_710,In_1085);
nand U487 (N_487,In_2054,In_2649);
nor U488 (N_488,In_2493,In_743);
and U489 (N_489,In_2523,In_782);
or U490 (N_490,In_1217,In_349);
and U491 (N_491,In_306,In_137);
nand U492 (N_492,In_1208,In_2085);
and U493 (N_493,In_1864,In_1390);
xor U494 (N_494,In_1431,In_1054);
xnor U495 (N_495,In_278,In_729);
nand U496 (N_496,In_434,In_2043);
nand U497 (N_497,In_346,In_1226);
nor U498 (N_498,In_135,In_1129);
xor U499 (N_499,In_63,In_2344);
nor U500 (N_500,In_1006,In_1199);
nand U501 (N_501,In_1035,In_1314);
and U502 (N_502,In_93,In_1413);
nand U503 (N_503,In_2115,In_2876);
and U504 (N_504,In_2733,In_2553);
or U505 (N_505,In_2494,In_2663);
nor U506 (N_506,In_2820,In_2217);
or U507 (N_507,In_1163,In_1522);
xnor U508 (N_508,In_1948,In_128);
and U509 (N_509,In_1601,In_2910);
nand U510 (N_510,In_2273,In_204);
and U511 (N_511,In_1558,In_496);
nor U512 (N_512,In_147,In_1026);
or U513 (N_513,In_700,In_685);
nand U514 (N_514,In_1485,In_2478);
nand U515 (N_515,In_843,In_751);
and U516 (N_516,In_1817,In_408);
and U517 (N_517,In_1576,In_1633);
or U518 (N_518,In_2212,In_1879);
nand U519 (N_519,In_108,In_2934);
and U520 (N_520,In_3,In_1585);
nor U521 (N_521,In_1887,In_1113);
nor U522 (N_522,In_1376,In_244);
xnor U523 (N_523,In_2293,In_2591);
or U524 (N_524,In_2160,In_2661);
nand U525 (N_525,In_1302,In_2249);
and U526 (N_526,In_395,In_1546);
or U527 (N_527,In_753,In_1945);
and U528 (N_528,In_2797,In_2799);
xnor U529 (N_529,In_439,In_2755);
nor U530 (N_530,In_1318,In_1894);
xnor U531 (N_531,In_1770,In_1222);
nand U532 (N_532,In_2488,In_1866);
or U533 (N_533,In_1268,In_1592);
and U534 (N_534,In_120,In_225);
and U535 (N_535,In_2090,In_885);
xor U536 (N_536,In_1262,In_2303);
xnor U537 (N_537,In_688,In_1312);
and U538 (N_538,In_2660,In_2882);
nand U539 (N_539,In_1264,In_190);
xnor U540 (N_540,In_400,In_2061);
xor U541 (N_541,In_915,In_2922);
nor U542 (N_542,In_2942,In_833);
nand U543 (N_543,In_2952,In_2657);
nor U544 (N_544,In_581,In_1952);
nor U545 (N_545,In_111,In_845);
or U546 (N_546,In_2071,In_1978);
and U547 (N_547,In_2608,In_912);
nor U548 (N_548,In_2197,In_1086);
nor U549 (N_549,In_1547,In_2961);
and U550 (N_550,In_1561,In_2215);
nor U551 (N_551,In_319,In_2803);
nor U552 (N_552,In_803,In_1231);
and U553 (N_553,In_2915,In_844);
nor U554 (N_554,In_1204,In_280);
nor U555 (N_555,In_417,In_1730);
and U556 (N_556,In_1014,In_309);
nand U557 (N_557,In_1091,In_1944);
nor U558 (N_558,In_288,In_2087);
and U559 (N_559,In_2982,In_1674);
or U560 (N_560,In_1183,In_2486);
or U561 (N_561,In_2432,In_2981);
or U562 (N_562,In_1425,In_619);
or U563 (N_563,In_970,In_299);
xnor U564 (N_564,In_849,In_138);
or U565 (N_565,In_468,In_2485);
nand U566 (N_566,In_2870,In_2795);
nand U567 (N_567,In_817,In_1614);
or U568 (N_568,In_2914,In_666);
nand U569 (N_569,In_2596,In_1207);
nor U570 (N_570,In_968,In_1099);
nand U571 (N_571,In_2794,In_1853);
or U572 (N_572,In_1047,In_1648);
nand U573 (N_573,In_2894,In_2556);
or U574 (N_574,In_1295,In_2960);
and U575 (N_575,In_2975,In_644);
and U576 (N_576,In_1815,In_1820);
nor U577 (N_577,In_1877,In_1513);
and U578 (N_578,In_2224,In_1638);
nand U579 (N_579,In_1300,In_2921);
nand U580 (N_580,In_45,In_2006);
and U581 (N_581,In_1625,In_1847);
nor U582 (N_582,In_454,In_241);
nor U583 (N_583,In_650,In_1437);
and U584 (N_584,In_1888,In_1370);
and U585 (N_585,In_2132,In_341);
nand U586 (N_586,In_2631,In_2279);
nor U587 (N_587,In_2171,In_1843);
or U588 (N_588,In_112,In_1463);
nand U589 (N_589,In_1775,In_1912);
nor U590 (N_590,In_2599,In_441);
nor U591 (N_591,In_966,In_2543);
nor U592 (N_592,In_41,In_440);
nor U593 (N_593,In_2386,In_2187);
or U594 (N_594,In_1460,In_1550);
nor U595 (N_595,In_1899,In_2813);
nand U596 (N_596,In_2422,In_498);
nand U597 (N_597,In_2750,In_1456);
xnor U598 (N_598,In_902,In_2325);
or U599 (N_599,In_2764,In_2477);
or U600 (N_600,In_1061,In_946);
xor U601 (N_601,In_1036,In_2723);
nor U602 (N_602,In_1121,In_1209);
and U603 (N_603,In_580,In_1641);
and U604 (N_604,In_1067,In_1610);
or U605 (N_605,In_2519,In_329);
or U606 (N_606,In_2052,In_1371);
or U607 (N_607,In_2891,In_170);
xnor U608 (N_608,In_2114,In_358);
nand U609 (N_609,In_65,In_997);
nand U610 (N_610,In_1502,In_2913);
and U611 (N_611,In_938,In_1737);
and U612 (N_612,In_1464,In_493);
or U613 (N_613,In_1422,In_1517);
nor U614 (N_614,In_1606,In_1780);
and U615 (N_615,In_2190,In_2296);
or U616 (N_616,In_2188,In_770);
nand U617 (N_617,In_124,In_530);
xnor U618 (N_618,In_1846,In_637);
nor U619 (N_619,In_1308,In_448);
nand U620 (N_620,In_511,In_862);
nor U621 (N_621,In_2227,In_491);
and U622 (N_622,In_2711,In_1976);
nor U623 (N_623,In_1896,In_2471);
and U624 (N_624,In_1905,In_1495);
nand U625 (N_625,In_2467,In_489);
and U626 (N_626,In_2399,In_2868);
nand U627 (N_627,In_1404,In_1743);
nor U628 (N_628,In_1005,In_2176);
or U629 (N_629,In_1506,In_613);
nor U630 (N_630,In_555,In_2120);
nor U631 (N_631,In_1988,In_2695);
nand U632 (N_632,In_2781,In_33);
or U633 (N_633,In_2223,In_1511);
nor U634 (N_634,In_569,In_2195);
and U635 (N_635,In_1813,In_822);
xnor U636 (N_636,In_2292,In_689);
nand U637 (N_637,In_775,In_1494);
or U638 (N_638,In_1173,In_449);
nor U639 (N_639,In_1870,In_1339);
nor U640 (N_640,In_2686,In_2680);
nand U641 (N_641,In_114,In_1525);
xnor U642 (N_642,In_2277,In_27);
nor U643 (N_643,In_1551,In_986);
and U644 (N_644,In_2465,In_1322);
or U645 (N_645,In_1480,In_2286);
nand U646 (N_646,In_1761,In_46);
xor U647 (N_647,In_262,In_576);
nand U648 (N_648,In_1265,In_2306);
xnor U649 (N_649,In_1336,In_200);
nor U650 (N_650,In_143,In_1411);
and U651 (N_651,In_492,In_641);
nand U652 (N_652,In_1352,In_1837);
or U653 (N_653,In_38,In_1845);
nor U654 (N_654,In_1972,In_1408);
or U655 (N_655,In_1092,In_2792);
nand U656 (N_656,In_1911,In_672);
or U657 (N_657,In_575,In_514);
nor U658 (N_658,In_615,In_475);
nand U659 (N_659,In_1937,In_230);
nor U660 (N_660,In_1740,In_1805);
nand U661 (N_661,In_1578,In_166);
or U662 (N_662,In_2593,In_2233);
or U663 (N_663,In_2895,In_2736);
or U664 (N_664,In_2358,In_1971);
and U665 (N_665,In_2616,In_2668);
nor U666 (N_666,In_2288,In_1967);
or U667 (N_667,In_1996,In_2439);
nand U668 (N_668,In_126,In_851);
or U669 (N_669,In_1512,In_1051);
nor U670 (N_670,In_2307,In_2449);
or U671 (N_671,In_1854,In_947);
and U672 (N_672,In_2641,In_1275);
or U673 (N_673,In_130,In_2618);
and U674 (N_674,In_608,In_2679);
and U675 (N_675,In_1850,In_351);
or U676 (N_676,In_2466,In_316);
nor U677 (N_677,In_1194,In_387);
and U678 (N_678,In_2100,In_759);
nand U679 (N_679,In_1177,In_2238);
or U680 (N_680,In_1332,In_1120);
nand U681 (N_681,In_261,In_2320);
or U682 (N_682,In_1434,In_1801);
nor U683 (N_683,In_2741,In_223);
nor U684 (N_684,In_755,In_245);
xnor U685 (N_685,In_1544,In_105);
nor U686 (N_686,In_717,In_630);
xor U687 (N_687,In_1677,In_1731);
nor U688 (N_688,In_2181,In_2370);
or U689 (N_689,In_2692,In_872);
and U690 (N_690,In_929,In_1637);
or U691 (N_691,In_208,In_2715);
and U692 (N_692,In_2763,In_2455);
and U693 (N_693,In_374,In_2429);
xor U694 (N_694,In_2527,In_750);
or U695 (N_695,In_2650,In_976);
nand U696 (N_696,In_930,In_815);
nand U697 (N_697,In_1549,In_2562);
nand U698 (N_698,In_14,In_647);
nand U699 (N_699,In_2589,In_265);
nor U700 (N_700,In_461,In_353);
xor U701 (N_701,In_2014,In_2583);
nor U702 (N_702,In_1580,In_2481);
nor U703 (N_703,In_2414,In_602);
nand U704 (N_704,In_12,In_681);
nor U705 (N_705,In_2138,In_2435);
and U706 (N_706,In_1573,In_1657);
or U707 (N_707,In_81,In_1581);
nand U708 (N_708,In_1440,In_1974);
nor U709 (N_709,In_179,In_977);
and U710 (N_710,In_1444,In_1438);
and U711 (N_711,In_2248,In_407);
or U712 (N_712,In_2253,In_224);
nand U713 (N_713,In_118,In_155);
or U714 (N_714,In_1616,In_2359);
nand U715 (N_715,In_1632,In_2577);
and U716 (N_716,In_2568,In_1803);
and U717 (N_717,In_466,In_2629);
xor U718 (N_718,In_2978,In_1365);
and U719 (N_719,In_1034,In_2382);
xnor U720 (N_720,In_1510,In_1159);
xor U721 (N_721,In_2275,In_692);
nand U722 (N_722,In_2060,In_933);
xor U723 (N_723,In_794,In_44);
and U724 (N_724,In_2220,In_2545);
nand U725 (N_725,In_2456,In_71);
or U726 (N_726,In_1902,In_2355);
nor U727 (N_727,In_1709,In_2638);
nand U728 (N_728,In_791,In_339);
nand U729 (N_729,In_1210,In_1484);
or U730 (N_730,In_1881,In_2582);
nand U731 (N_731,In_15,In_2610);
and U732 (N_732,In_1793,In_1127);
or U733 (N_733,In_2191,In_1375);
nor U734 (N_734,In_2110,In_2991);
or U735 (N_735,In_310,In_2331);
nand U736 (N_736,In_1166,In_1338);
and U737 (N_737,In_1964,In_1983);
or U738 (N_738,In_2911,In_1211);
or U739 (N_739,In_846,In_1415);
or U740 (N_740,In_1571,In_2364);
and U741 (N_741,In_402,In_403);
or U742 (N_742,In_1516,In_432);
nand U743 (N_743,In_510,In_956);
and U744 (N_744,In_1534,In_1829);
nand U745 (N_745,In_463,In_139);
or U746 (N_746,In_1640,In_2920);
xor U747 (N_747,In_249,In_99);
or U748 (N_748,In_2685,In_515);
nor U749 (N_749,In_1663,In_2118);
nand U750 (N_750,In_2140,In_2572);
nand U751 (N_751,In_972,In_2039);
nand U752 (N_752,In_1326,In_697);
nor U753 (N_753,In_1151,In_2722);
and U754 (N_754,In_2049,In_1687);
nor U755 (N_755,In_1539,In_98);
nand U756 (N_756,In_385,In_2945);
or U757 (N_757,In_1101,In_2315);
nor U758 (N_758,In_276,In_719);
or U759 (N_759,In_2862,In_1328);
nor U760 (N_760,In_2503,In_1197);
nand U761 (N_761,In_1096,In_543);
nand U762 (N_762,In_1788,In_792);
and U763 (N_763,In_951,In_1873);
or U764 (N_764,In_2210,In_2706);
or U765 (N_765,In_2727,In_1405);
nand U766 (N_766,In_176,In_1167);
and U767 (N_767,In_2968,In_10);
and U768 (N_768,In_577,In_838);
and U769 (N_769,In_2879,In_1691);
xor U770 (N_770,In_2851,In_2174);
or U771 (N_771,In_2438,In_162);
xor U772 (N_772,In_772,In_495);
nand U773 (N_773,In_2354,In_2966);
xor U774 (N_774,In_2511,In_2430);
or U775 (N_775,In_2483,In_2263);
nand U776 (N_776,In_1174,In_1080);
nor U777 (N_777,In_2177,In_1671);
and U778 (N_778,In_1144,In_2598);
nor U779 (N_779,In_2935,In_77);
or U780 (N_780,In_1507,In_2407);
or U781 (N_781,In_686,In_1791);
xor U782 (N_782,In_2446,In_1355);
nand U783 (N_783,In_2996,In_597);
xnor U784 (N_784,In_557,In_2437);
or U785 (N_785,In_2240,In_1626);
nand U786 (N_786,In_1835,In_856);
nand U787 (N_787,In_1628,In_1862);
nor U788 (N_788,In_2837,In_568);
nand U789 (N_789,In_2533,In_381);
and U790 (N_790,In_1618,In_2383);
nand U791 (N_791,In_1462,In_1554);
xnor U792 (N_792,In_266,In_880);
nor U793 (N_793,In_958,In_2848);
nand U794 (N_794,In_922,In_1848);
or U795 (N_795,In_1307,In_1182);
xnor U796 (N_796,In_552,In_1252);
or U797 (N_797,In_907,In_1257);
nor U798 (N_798,In_1984,In_1320);
or U799 (N_799,In_953,In_991);
nor U800 (N_800,In_1538,In_2390);
nand U801 (N_801,In_2925,In_1483);
or U802 (N_802,In_936,In_11);
nor U803 (N_803,In_640,In_1298);
nor U804 (N_804,In_1738,In_2758);
xor U805 (N_805,In_1682,In_1833);
nor U806 (N_806,In_1423,In_2815);
nand U807 (N_807,In_2846,In_1520);
or U808 (N_808,In_518,In_2097);
or U809 (N_809,In_998,In_508);
and U810 (N_810,In_1668,In_2351);
xor U811 (N_811,In_1868,In_2496);
or U812 (N_812,In_211,In_2713);
or U813 (N_813,In_2863,In_1356);
and U814 (N_814,In_36,In_2350);
nor U815 (N_815,In_2783,In_573);
nand U816 (N_816,In_1959,In_2927);
and U817 (N_817,In_2236,In_2209);
and U818 (N_818,In_1942,In_1123);
nor U819 (N_819,In_418,In_1876);
and U820 (N_820,In_332,In_2754);
and U821 (N_821,In_487,In_2932);
and U822 (N_822,In_1799,In_509);
nor U823 (N_823,In_1311,In_1492);
nand U824 (N_824,In_2395,In_2330);
or U825 (N_825,In_465,In_722);
nor U826 (N_826,In_1443,In_773);
xor U827 (N_827,In_2571,In_2208);
and U828 (N_828,In_82,In_2309);
or U829 (N_829,In_571,In_1102);
and U830 (N_830,In_545,In_1243);
and U831 (N_831,In_2765,In_409);
nor U832 (N_832,In_2947,In_1193);
nand U833 (N_833,In_1386,In_1872);
xor U834 (N_834,In_2172,In_857);
nor U835 (N_835,In_264,In_1116);
nand U836 (N_836,In_25,In_362);
nand U837 (N_837,In_1891,In_1747);
xor U838 (N_838,In_2953,In_1001);
and U839 (N_839,In_422,In_1994);
or U840 (N_840,In_292,In_520);
nor U841 (N_841,In_2468,In_2936);
nor U842 (N_842,In_251,In_1536);
and U843 (N_843,In_1347,In_1450);
and U844 (N_844,In_1087,In_2336);
and U845 (N_845,In_1003,In_363);
nor U846 (N_846,In_671,In_716);
and U847 (N_847,In_2025,In_818);
or U848 (N_848,In_2319,In_2998);
nand U849 (N_849,In_2622,In_1429);
nand U850 (N_850,In_2231,In_1451);
and U851 (N_851,In_24,In_95);
nand U852 (N_852,In_2992,In_1310);
nor U853 (N_853,In_2828,In_2643);
and U854 (N_854,In_296,In_1152);
or U855 (N_855,In_1068,In_1825);
or U856 (N_856,In_1622,In_2818);
xor U857 (N_857,In_806,In_2565);
nand U858 (N_858,In_2143,In_1057);
nand U859 (N_859,In_1947,In_1567);
nor U860 (N_860,In_1333,In_2459);
nand U861 (N_861,In_2747,In_1077);
nor U862 (N_862,In_1331,In_1324);
nor U863 (N_863,In_1461,In_1299);
and U864 (N_864,In_1595,In_847);
xor U865 (N_865,In_1246,In_809);
nand U866 (N_866,In_217,In_2416);
or U867 (N_867,In_1679,In_1966);
nand U868 (N_868,In_97,In_1285);
nand U869 (N_869,In_601,In_1773);
or U870 (N_870,In_796,In_2578);
nor U871 (N_871,In_8,In_1179);
nor U872 (N_872,In_1039,In_2009);
or U873 (N_873,In_1666,In_2035);
nand U874 (N_874,In_1920,In_2611);
or U875 (N_875,In_1229,In_2064);
nand U876 (N_876,In_2504,In_553);
nand U877 (N_877,In_2057,In_1482);
or U878 (N_878,In_752,In_1897);
or U879 (N_879,In_1713,In_2031);
nand U880 (N_880,In_2564,In_1871);
nor U881 (N_881,In_2905,In_850);
nand U882 (N_882,In_795,In_2645);
and U883 (N_883,In_1249,In_739);
nand U884 (N_884,In_1577,In_616);
and U885 (N_885,In_1969,In_589);
nand U886 (N_886,In_43,In_304);
xnor U887 (N_887,In_785,In_1076);
or U888 (N_888,In_425,In_470);
and U889 (N_889,In_1508,In_1004);
or U890 (N_890,In_674,In_2297);
and U891 (N_891,In_964,In_177);
nand U892 (N_892,In_450,In_825);
nand U893 (N_893,In_2900,In_1472);
nand U894 (N_894,In_2694,In_122);
or U895 (N_895,In_2201,In_1587);
xnor U896 (N_896,In_916,In_1653);
and U897 (N_897,In_1424,In_2896);
and U898 (N_898,In_2537,In_368);
and U899 (N_899,In_416,In_2075);
nor U900 (N_900,In_1323,In_384);
or U901 (N_901,In_1452,In_2084);
nor U902 (N_902,In_649,In_2801);
nor U903 (N_903,In_424,In_2807);
and U904 (N_904,In_1953,In_2086);
nand U905 (N_905,In_758,In_2228);
nand U906 (N_906,In_2470,In_2357);
and U907 (N_907,In_2603,In_620);
nor U908 (N_908,In_9,In_158);
nor U909 (N_909,In_1704,In_1137);
nand U910 (N_910,In_566,In_142);
or U911 (N_911,In_2234,In_2164);
xor U912 (N_912,In_1361,In_1342);
or U913 (N_913,In_1958,In_173);
xor U914 (N_914,In_2512,In_2548);
nand U915 (N_915,In_2832,In_1394);
nand U916 (N_916,In_2391,In_2226);
nor U917 (N_917,In_1358,In_1198);
nor U918 (N_918,In_4,In_702);
xnor U919 (N_919,In_1828,In_1783);
xor U920 (N_920,In_2495,In_218);
xor U921 (N_921,In_592,In_2689);
and U922 (N_922,In_2451,In_2502);
nand U923 (N_923,In_2574,In_78);
nor U924 (N_924,In_1884,In_559);
and U925 (N_925,In_89,In_102);
or U926 (N_926,In_1267,In_456);
xnor U927 (N_927,In_1729,In_2698);
nor U928 (N_928,In_799,In_1421);
nor U929 (N_929,In_1058,In_2811);
nand U930 (N_930,In_1048,In_380);
nand U931 (N_931,In_1184,In_2983);
nand U932 (N_932,In_1842,In_1631);
or U933 (N_933,In_2008,In_101);
xnor U934 (N_934,In_1368,In_1150);
or U935 (N_935,In_804,In_748);
nor U936 (N_936,In_1521,In_2532);
nand U937 (N_937,In_2001,In_2898);
nor U938 (N_938,In_680,In_206);
and U939 (N_939,In_2213,In_1702);
nor U940 (N_940,In_1171,In_1213);
nor U941 (N_941,In_2938,In_275);
nor U942 (N_942,In_1851,In_2068);
nor U943 (N_943,In_373,In_1568);
nor U944 (N_944,In_660,In_1926);
or U945 (N_945,In_1756,In_2421);
nor U946 (N_946,In_436,In_2185);
and U947 (N_947,In_2659,In_1931);
nand U948 (N_948,In_0,In_2094);
nor U949 (N_949,In_308,In_625);
or U950 (N_950,In_2607,In_1109);
and U951 (N_951,In_2184,In_2193);
nor U952 (N_952,In_2380,In_1860);
and U953 (N_953,In_227,In_2993);
and U954 (N_954,In_236,In_485);
and U955 (N_955,In_2732,In_1627);
nor U956 (N_956,In_2652,In_1924);
xnor U957 (N_957,In_1040,In_1987);
or U958 (N_958,In_421,In_1720);
or U959 (N_959,In_1412,In_1050);
and U960 (N_960,In_2093,In_2609);
nand U961 (N_961,In_2926,In_1042);
nor U962 (N_962,In_2314,In_2904);
nand U963 (N_963,In_232,In_2521);
nor U964 (N_964,In_2990,In_2144);
or U965 (N_965,In_1769,In_720);
and U966 (N_966,In_1909,In_85);
and U967 (N_967,In_254,In_572);
nand U968 (N_968,In_2594,In_1296);
xnor U969 (N_969,In_992,In_2845);
and U970 (N_970,In_2646,In_2985);
nand U971 (N_971,In_221,In_1325);
nand U972 (N_972,In_1865,In_2230);
and U973 (N_973,In_1838,In_88);
and U974 (N_974,In_1223,In_2605);
nand U975 (N_975,In_1074,In_1940);
nor U976 (N_976,In_2419,In_167);
and U977 (N_977,In_2427,In_583);
nor U978 (N_978,In_1718,In_1739);
xnor U979 (N_979,In_1214,In_591);
and U980 (N_980,In_814,In_359);
xnor U981 (N_981,In_34,In_1383);
nand U982 (N_982,In_1488,In_1736);
or U983 (N_983,In_2353,In_2244);
nor U984 (N_984,In_2771,In_2955);
nand U985 (N_985,In_978,In_302);
nand U986 (N_986,In_1652,In_414);
nand U987 (N_987,In_2693,In_2836);
or U988 (N_988,In_2167,In_662);
nand U989 (N_989,In_1569,In_1572);
nor U990 (N_990,In_740,In_1680);
nand U991 (N_991,In_484,In_1271);
and U992 (N_992,In_585,In_1071);
xnor U993 (N_993,In_1901,In_1496);
and U994 (N_994,In_1635,In_1291);
xor U995 (N_995,In_2047,In_1453);
or U996 (N_996,In_2378,In_730);
or U997 (N_997,In_226,In_205);
nand U998 (N_998,In_2710,In_1072);
and U999 (N_999,In_1041,In_1292);
and U1000 (N_1000,In_643,In_2567);
nand U1001 (N_1001,In_2261,In_1031);
nand U1002 (N_1002,In_2487,In_741);
or U1003 (N_1003,In_2402,In_622);
and U1004 (N_1004,In_1776,In_2152);
nand U1005 (N_1005,In_246,In_656);
nand U1006 (N_1006,In_2299,In_1645);
and U1007 (N_1007,In_2023,In_1140);
nor U1008 (N_1008,In_1841,In_1487);
nor U1009 (N_1009,In_1191,In_1792);
xnor U1010 (N_1010,In_2196,In_969);
xnor U1011 (N_1011,In_1938,In_2821);
nand U1012 (N_1012,In_1470,In_2091);
nor U1013 (N_1013,In_1240,In_800);
nand U1014 (N_1014,In_835,In_2884);
and U1015 (N_1015,In_1661,In_2778);
and U1016 (N_1016,In_2708,In_540);
nor U1017 (N_1017,In_1465,In_1066);
nand U1018 (N_1018,In_551,In_2038);
nor U1019 (N_1019,In_1607,In_1777);
nor U1020 (N_1020,In_2316,In_636);
nand U1021 (N_1021,In_2246,In_642);
nor U1022 (N_1022,In_1114,In_2055);
or U1023 (N_1023,In_2397,In_1917);
or U1024 (N_1024,In_1505,In_2703);
or U1025 (N_1025,In_2971,In_1613);
or U1026 (N_1026,In_579,In_1276);
nand U1027 (N_1027,In_1700,In_343);
nand U1028 (N_1028,In_2417,In_234);
and U1029 (N_1029,In_726,In_1143);
and U1030 (N_1030,In_974,In_2113);
xnor U1031 (N_1031,In_2200,In_627);
and U1032 (N_1032,In_2871,In_2560);
nand U1033 (N_1033,In_2769,In_1787);
nor U1034 (N_1034,In_606,In_80);
nor U1035 (N_1035,In_2808,In_1690);
and U1036 (N_1036,In_1918,In_2290);
or U1037 (N_1037,In_1929,In_47);
nor U1038 (N_1038,In_2070,In_477);
xnor U1039 (N_1039,In_2428,In_397);
nor U1040 (N_1040,In_1685,In_2912);
xor U1041 (N_1041,In_1733,In_2805);
or U1042 (N_1042,In_199,In_420);
nor U1043 (N_1043,In_2050,In_1855);
nor U1044 (N_1044,In_1686,In_1454);
nor U1045 (N_1045,In_2866,In_623);
nor U1046 (N_1046,In_879,In_1377);
and U1047 (N_1047,In_2976,In_1245);
or U1048 (N_1048,In_767,In_2677);
xnor U1049 (N_1049,In_2964,In_2122);
and U1050 (N_1050,In_1615,In_238);
or U1051 (N_1051,In_1290,In_1946);
nor U1052 (N_1052,In_2989,In_2550);
or U1053 (N_1053,In_1237,In_482);
or U1054 (N_1054,In_766,In_182);
nor U1055 (N_1055,In_365,In_376);
nor U1056 (N_1056,In_2654,In_2016);
or U1057 (N_1057,In_639,In_883);
nand U1058 (N_1058,In_2340,In_2841);
or U1059 (N_1059,In_1457,In_1138);
or U1060 (N_1060,In_486,In_2368);
or U1061 (N_1061,In_1297,In_2946);
nand U1062 (N_1062,In_1874,In_2372);
xnor U1063 (N_1063,In_565,In_1476);
or U1064 (N_1064,In_2943,In_2027);
and U1065 (N_1065,In_1939,In_2530);
and U1066 (N_1066,In_904,In_1755);
and U1067 (N_1067,In_2490,In_2460);
or U1068 (N_1068,In_1497,In_2426);
nand U1069 (N_1069,In_609,In_1442);
xnor U1070 (N_1070,In_2218,In_1169);
or U1071 (N_1071,In_945,In_990);
nand U1072 (N_1072,In_2541,In_1063);
nor U1073 (N_1073,In_2536,In_2492);
nand U1074 (N_1074,In_1602,In_2141);
nor U1075 (N_1075,In_1329,In_1420);
and U1076 (N_1076,In_893,In_519);
and U1077 (N_1077,In_673,In_873);
and U1078 (N_1078,In_1992,In_1712);
or U1079 (N_1079,In_2204,In_2697);
nand U1080 (N_1080,In_1281,In_1279);
and U1081 (N_1081,In_1744,In_2324);
or U1082 (N_1082,In_1694,In_1321);
and U1083 (N_1083,In_87,In_2108);
nor U1084 (N_1084,In_257,In_198);
or U1085 (N_1085,In_2705,In_1261);
and U1086 (N_1086,In_192,In_159);
nor U1087 (N_1087,In_805,In_1922);
nor U1088 (N_1088,In_2221,In_91);
nand U1089 (N_1089,In_2901,In_926);
or U1090 (N_1090,In_2475,In_287);
nand U1091 (N_1091,In_2002,In_2809);
nand U1092 (N_1092,In_655,In_1146);
nor U1093 (N_1093,In_457,In_1961);
nand U1094 (N_1094,In_2875,In_2337);
and U1095 (N_1095,In_2326,In_812);
or U1096 (N_1096,In_1212,In_2137);
nand U1097 (N_1097,In_808,In_524);
or U1098 (N_1098,In_144,In_2222);
or U1099 (N_1099,In_2563,In_1490);
and U1100 (N_1100,In_1925,In_1532);
or U1101 (N_1101,In_1771,In_1955);
and U1102 (N_1102,In_1139,In_2670);
or U1103 (N_1103,In_2145,In_746);
or U1104 (N_1104,In_1706,In_1280);
nor U1105 (N_1105,In_197,In_2767);
nor U1106 (N_1106,In_1989,In_115);
nor U1107 (N_1107,In_1785,In_360);
or U1108 (N_1108,In_648,In_522);
or U1109 (N_1109,In_1345,In_1982);
nor U1110 (N_1110,In_1045,In_433);
nand U1111 (N_1111,In_860,In_2051);
nand U1112 (N_1112,In_212,In_2088);
or U1113 (N_1113,In_1617,In_2425);
xnor U1114 (N_1114,In_1176,In_853);
and U1115 (N_1115,In_2954,In_2322);
nor U1116 (N_1116,In_1816,In_2304);
nor U1117 (N_1117,In_826,In_2786);
and U1118 (N_1118,In_132,In_2067);
nor U1119 (N_1119,In_2555,In_2874);
nand U1120 (N_1120,In_479,In_149);
xnor U1121 (N_1121,In_2600,In_1293);
and U1122 (N_1122,In_2597,In_858);
xor U1123 (N_1123,In_2415,In_909);
or U1124 (N_1124,In_2919,In_1104);
and U1125 (N_1125,In_2032,In_2266);
nand U1126 (N_1126,In_2570,In_1062);
or U1127 (N_1127,In_676,In_2029);
nor U1128 (N_1128,In_2165,In_949);
or U1129 (N_1129,In_2676,In_704);
and U1130 (N_1130,In_2183,In_344);
or U1131 (N_1131,In_603,In_2381);
nor U1132 (N_1132,In_293,In_1840);
nor U1133 (N_1133,In_1800,In_979);
nor U1134 (N_1134,In_2310,In_1089);
nor U1135 (N_1135,In_765,In_2173);
and U1136 (N_1136,In_5,In_2476);
or U1137 (N_1137,In_1270,In_1020);
or U1138 (N_1138,In_2484,In_1126);
and U1139 (N_1139,In_1998,In_1867);
nand U1140 (N_1140,In_289,In_1471);
or U1141 (N_1141,In_1895,In_2129);
and U1142 (N_1142,In_2718,In_771);
nor U1143 (N_1143,In_1584,In_321);
and U1144 (N_1144,In_2857,In_1893);
nor U1145 (N_1145,In_258,In_1064);
nor U1146 (N_1146,In_2489,In_2825);
nor U1147 (N_1147,In_661,In_528);
nand U1148 (N_1148,In_2892,In_1684);
nor U1149 (N_1149,In_705,In_2756);
or U1150 (N_1150,In_2457,In_1469);
and U1151 (N_1151,In_1106,In_1136);
nor U1152 (N_1152,In_1010,In_2130);
and U1153 (N_1153,In_370,In_1889);
or U1154 (N_1154,In_1305,In_2211);
nor U1155 (N_1155,In_1235,In_2198);
nor U1156 (N_1156,In_286,In_2861);
nor U1157 (N_1157,In_2651,In_1233);
nand U1158 (N_1158,In_2447,In_2497);
or U1159 (N_1159,In_52,In_1403);
and U1160 (N_1160,In_2258,In_1728);
nor U1161 (N_1161,In_1254,In_2856);
xor U1162 (N_1162,In_1201,In_2251);
or U1163 (N_1163,In_164,In_1396);
or U1164 (N_1164,In_1603,In_1753);
nand U1165 (N_1165,In_2146,In_865);
nor U1166 (N_1166,In_2579,In_624);
nor U1167 (N_1167,In_1807,In_1543);
and U1168 (N_1168,In_1863,In_984);
and U1169 (N_1169,In_2768,In_203);
and U1170 (N_1170,In_478,In_488);
and U1171 (N_1171,In_1186,In_1172);
nand U1172 (N_1172,In_679,In_2507);
nand U1173 (N_1173,In_2312,In_2065);
and U1174 (N_1174,In_2018,In_1921);
xor U1175 (N_1175,In_37,In_1378);
and U1176 (N_1176,In_1900,In_2743);
nor U1177 (N_1177,In_2345,In_2139);
or U1178 (N_1178,In_2636,In_1913);
and U1179 (N_1179,In_1110,In_2418);
nand U1180 (N_1180,In_2250,In_2941);
nand U1181 (N_1181,In_2294,In_2333);
and U1182 (N_1182,In_2282,In_2902);
or U1183 (N_1183,In_1766,In_731);
nand U1184 (N_1184,In_694,In_2623);
and U1185 (N_1185,In_2986,In_1990);
xor U1186 (N_1186,In_1683,In_2897);
nor U1187 (N_1187,In_2534,In_72);
xnor U1188 (N_1188,In_2104,In_2740);
and U1189 (N_1189,In_737,In_645);
nand U1190 (N_1190,In_2308,In_2095);
nor U1191 (N_1191,In_861,In_2760);
nor U1192 (N_1192,In_1133,In_1075);
nand U1193 (N_1193,In_1647,In_268);
and U1194 (N_1194,In_1446,In_1954);
or U1195 (N_1195,In_2444,In_336);
or U1196 (N_1196,In_919,In_2242);
nand U1197 (N_1197,In_1936,In_1530);
or U1198 (N_1198,In_541,In_2232);
and U1199 (N_1199,In_1556,In_1886);
nor U1200 (N_1200,In_1019,In_1965);
nor U1201 (N_1201,In_129,In_1540);
or U1202 (N_1202,In_1719,In_2124);
xor U1203 (N_1203,In_2317,In_19);
or U1204 (N_1204,In_207,In_2700);
nor U1205 (N_1205,In_1479,In_2182);
nand U1206 (N_1206,In_2777,In_194);
and U1207 (N_1207,In_628,In_307);
nor U1208 (N_1208,In_1220,In_2291);
or U1209 (N_1209,In_1115,In_878);
nand U1210 (N_1210,In_1239,In_1823);
nor U1211 (N_1211,In_2089,In_1570);
nand U1212 (N_1212,In_2712,In_1230);
nor U1213 (N_1213,In_604,In_2831);
xnor U1214 (N_1214,In_174,In_2634);
xor U1215 (N_1215,In_989,In_797);
nor U1216 (N_1216,In_2436,In_590);
nand U1217 (N_1217,In_1402,In_444);
and U1218 (N_1218,In_1703,In_554);
nand U1219 (N_1219,In_723,In_1981);
nor U1220 (N_1220,In_728,In_2738);
nor U1221 (N_1221,In_1128,In_1649);
xor U1222 (N_1222,In_1795,In_1284);
nand U1223 (N_1223,In_2410,In_163);
nand U1224 (N_1224,In_2341,In_2321);
or U1225 (N_1225,In_1149,In_2431);
nand U1226 (N_1226,In_1335,In_903);
or U1227 (N_1227,In_2586,In_1970);
nor U1228 (N_1228,In_501,In_2101);
xnor U1229 (N_1229,In_2366,In_1812);
and U1230 (N_1230,In_866,In_2338);
xor U1231 (N_1231,In_1943,In_1646);
and U1232 (N_1232,In_242,In_935);
nor U1233 (N_1233,In_2162,In_1350);
nor U1234 (N_1234,In_871,In_537);
nor U1235 (N_1235,In_2081,In_2744);
and U1236 (N_1236,In_2974,In_472);
nand U1237 (N_1237,In_354,In_895);
nand U1238 (N_1238,In_517,In_2376);
xor U1239 (N_1239,In_110,In_2022);
xor U1240 (N_1240,In_841,In_2254);
nor U1241 (N_1241,In_2724,In_1009);
nand U1242 (N_1242,In_2640,In_2753);
nand U1243 (N_1243,In_2005,In_2180);
nand U1244 (N_1244,In_1260,In_669);
nor U1245 (N_1245,In_1662,In_2313);
nor U1246 (N_1246,In_900,In_2899);
nor U1247 (N_1247,In_925,In_2872);
and U1248 (N_1248,In_2965,In_1725);
nand U1249 (N_1249,In_2782,In_889);
nand U1250 (N_1250,In_1809,In_693);
and U1251 (N_1251,In_2790,In_1060);
nand U1252 (N_1252,In_58,In_1597);
nand U1253 (N_1253,In_749,In_342);
nand U1254 (N_1254,In_2268,In_2517);
and U1255 (N_1255,In_910,In_1742);
nor U1256 (N_1256,In_2479,In_1509);
nor U1257 (N_1257,In_161,In_1748);
or U1258 (N_1258,In_943,In_1478);
and U1259 (N_1259,In_1148,In_2371);
or U1260 (N_1260,In_1491,In_1168);
or U1261 (N_1261,In_2367,In_2192);
nand U1262 (N_1262,In_811,In_1892);
xor U1263 (N_1263,In_677,In_781);
nand U1264 (N_1264,In_2106,In_1806);
and U1265 (N_1265,In_1337,In_882);
and U1266 (N_1266,In_1032,In_2972);
or U1267 (N_1267,In_899,In_462);
or U1268 (N_1268,In_184,In_1919);
nand U1269 (N_1269,In_2396,In_1608);
and U1270 (N_1270,In_413,In_2159);
and U1271 (N_1271,In_981,In_1898);
nor U1272 (N_1272,In_2013,In_2041);
or U1273 (N_1273,In_2034,In_423);
nor U1274 (N_1274,In_1672,In_761);
nand U1275 (N_1275,In_1675,In_1432);
and U1276 (N_1276,In_993,In_735);
nor U1277 (N_1277,In_894,In_270);
nand U1278 (N_1278,In_1409,In_1353);
or U1279 (N_1279,In_1043,In_2271);
nor U1280 (N_1280,In_786,In_267);
and U1281 (N_1281,In_2362,In_334);
nand U1282 (N_1282,In_593,In_2349);
nor U1283 (N_1283,In_1754,In_411);
xor U1284 (N_1284,In_447,In_1131);
nor U1285 (N_1285,In_1710,In_1154);
or U1286 (N_1286,In_1319,In_913);
and U1287 (N_1287,In_1774,In_955);
or U1288 (N_1288,In_2940,In_2635);
xor U1289 (N_1289,In_646,In_908);
xor U1290 (N_1290,In_564,In_410);
nand U1291 (N_1291,In_1117,In_634);
nor U1292 (N_1292,In_2142,In_2257);
and U1293 (N_1293,In_2816,In_1562);
or U1294 (N_1294,In_1802,In_2984);
nand U1295 (N_1295,In_570,In_202);
nand U1296 (N_1296,In_300,In_1639);
or U1297 (N_1297,In_1289,In_1957);
and U1298 (N_1298,In_168,In_1022);
xnor U1299 (N_1299,In_1636,In_1357);
nor U1300 (N_1300,In_2405,In_824);
nand U1301 (N_1301,In_1611,In_790);
nor U1302 (N_1302,In_1612,In_1185);
or U1303 (N_1303,In_2385,In_1531);
nand U1304 (N_1304,In_201,In_460);
xor U1305 (N_1305,In_2780,In_59);
and U1306 (N_1306,In_2587,In_2161);
or U1307 (N_1307,In_868,In_2907);
nor U1308 (N_1308,In_2681,In_1205);
nor U1309 (N_1309,In_2632,In_330);
nor U1310 (N_1310,In_1609,In_1605);
nor U1311 (N_1311,In_1373,In_356);
or U1312 (N_1312,In_2015,In_2062);
or U1313 (N_1313,In_1665,In_2335);
nor U1314 (N_1314,In_884,In_1579);
nand U1315 (N_1315,In_2524,In_2542);
nor U1316 (N_1316,In_897,In_924);
and U1317 (N_1317,In_331,In_2633);
nor U1318 (N_1318,In_317,In_682);
and U1319 (N_1319,In_61,In_2864);
nand U1320 (N_1320,In_1112,In_2612);
nand U1321 (N_1321,In_322,In_736);
nand U1322 (N_1322,In_2469,In_712);
nor U1323 (N_1323,In_2852,In_2278);
or U1324 (N_1324,In_2026,In_1049);
nand U1325 (N_1325,In_1007,In_248);
or U1326 (N_1326,In_1634,In_1364);
nor U1327 (N_1327,In_2131,In_2696);
or U1328 (N_1328,In_172,In_980);
nand U1329 (N_1329,In_2528,In_539);
xor U1330 (N_1330,In_323,In_260);
and U1331 (N_1331,In_932,In_2513);
or U1332 (N_1332,In_2028,In_2);
and U1333 (N_1333,In_1188,In_1232);
or U1334 (N_1334,In_273,In_2858);
nand U1335 (N_1335,In_2074,In_1344);
xnor U1336 (N_1336,In_1583,In_2924);
or U1337 (N_1337,In_988,In_1228);
and U1338 (N_1338,In_975,In_2125);
nor U1339 (N_1339,In_1221,In_1219);
nand U1340 (N_1340,In_832,In_2658);
or U1341 (N_1341,In_1999,In_1673);
or U1342 (N_1342,In_328,In_366);
and U1343 (N_1343,In_490,In_967);
or U1344 (N_1344,In_2272,In_35);
nand U1345 (N_1345,In_294,In_1564);
and U1346 (N_1346,In_53,In_2647);
nand U1347 (N_1347,In_1306,In_1083);
and U1348 (N_1348,In_2403,In_1384);
nor U1349 (N_1349,In_783,In_1190);
nand U1350 (N_1350,In_854,In_2707);
and U1351 (N_1351,In_2928,In_2166);
or U1352 (N_1352,In_2066,In_2615);
nor U1353 (N_1353,In_1493,In_535);
or U1354 (N_1354,In_745,In_2256);
nand U1355 (N_1355,In_2973,In_2346);
or U1356 (N_1356,In_96,In_768);
or U1357 (N_1357,In_2584,In_512);
and U1358 (N_1358,In_1088,In_2205);
xnor U1359 (N_1359,In_2044,In_1760);
nor U1360 (N_1360,In_233,In_1037);
or U1361 (N_1361,In_2721,In_678);
or U1362 (N_1362,In_1153,In_1224);
nand U1363 (N_1363,In_2472,In_7);
nor U1364 (N_1364,In_2585,In_1764);
or U1365 (N_1365,In_263,In_1393);
nor U1366 (N_1366,In_2883,In_2554);
xor U1367 (N_1367,In_2869,In_533);
nor U1368 (N_1368,In_1426,In_51);
nor U1369 (N_1369,In_148,In_1398);
or U1370 (N_1370,In_2117,In_2734);
nand U1371 (N_1371,In_2361,In_2289);
and U1372 (N_1372,In_2509,In_2021);
and U1373 (N_1373,In_243,In_1529);
nand U1374 (N_1374,In_1698,In_2498);
or U1375 (N_1375,In_355,In_386);
or U1376 (N_1376,In_40,In_1098);
nand U1377 (N_1377,In_146,In_2175);
and U1378 (N_1378,In_2365,In_1346);
and U1379 (N_1379,In_2601,In_1928);
nor U1380 (N_1380,In_104,In_1852);
and U1381 (N_1381,In_787,In_2829);
nor U1382 (N_1382,In_598,In_2630);
or U1383 (N_1383,In_2994,In_2819);
and U1384 (N_1384,In_1241,In_1025);
nand U1385 (N_1385,In_502,In_2788);
nor U1386 (N_1386,In_2389,In_1875);
or U1387 (N_1387,In_50,In_2529);
nor U1388 (N_1388,In_1849,In_703);
nor U1389 (N_1389,In_1746,In_1428);
and U1390 (N_1390,In_941,In_574);
or U1391 (N_1391,In_2400,In_2671);
and U1392 (N_1392,In_2078,In_1382);
and U1393 (N_1393,In_237,In_1878);
or U1394 (N_1394,In_874,In_1097);
and U1395 (N_1395,In_1202,In_68);
and U1396 (N_1396,In_2588,In_777);
nor U1397 (N_1397,In_1620,In_1810);
and U1398 (N_1398,In_187,In_1105);
nand U1399 (N_1399,In_222,In_544);
xor U1400 (N_1400,In_2843,In_2888);
or U1401 (N_1401,In_1765,In_2746);
or U1402 (N_1402,In_2675,In_2644);
nand U1403 (N_1403,In_1447,In_2890);
nor U1404 (N_1404,In_587,In_2147);
nor U1405 (N_1405,In_652,In_1103);
nand U1406 (N_1406,In_2995,In_707);
nor U1407 (N_1407,In_1890,In_2835);
nor U1408 (N_1408,In_398,In_2889);
or U1409 (N_1409,In_2827,In_2653);
nor U1410 (N_1410,In_2123,In_1327);
or U1411 (N_1411,In_928,In_2107);
nand U1412 (N_1412,In_1073,In_21);
nand U1413 (N_1413,In_2526,In_228);
nand U1414 (N_1414,In_446,In_2725);
nor U1415 (N_1415,In_906,In_2374);
or U1416 (N_1416,In_891,In_2239);
nor U1417 (N_1417,In_1340,In_1407);
xnor U1418 (N_1418,In_629,In_2119);
xor U1419 (N_1419,In_971,In_638);
and U1420 (N_1420,In_2127,In_877);
and U1421 (N_1421,In_1956,In_1623);
or U1422 (N_1422,In_864,In_1349);
or U1423 (N_1423,In_2423,In_1286);
xor U1424 (N_1424,In_2604,In_994);
nor U1425 (N_1425,In_1930,In_2662);
or U1426 (N_1426,In_1385,In_2458);
and U1427 (N_1427,In_1779,In_1586);
nor U1428 (N_1428,In_952,In_1448);
nor U1429 (N_1429,In_2328,In_26);
and U1430 (N_1430,In_1282,In_2787);
and U1431 (N_1431,In_361,In_1236);
and U1432 (N_1432,In_2762,In_1259);
or U1433 (N_1433,In_944,In_390);
nor U1434 (N_1434,In_982,In_1038);
nor U1435 (N_1435,In_127,In_905);
nand U1436 (N_1436,In_823,In_2880);
and U1437 (N_1437,In_695,In_290);
nor U1438 (N_1438,In_1819,In_1468);
or U1439 (N_1439,In_1693,In_1017);
nor U1440 (N_1440,In_1255,In_2348);
nand U1441 (N_1441,In_2557,In_733);
and U1442 (N_1442,In_701,In_1187);
and U1443 (N_1443,In_2637,In_2134);
nand U1444 (N_1444,In_1348,In_56);
or U1445 (N_1445,In_1263,In_855);
and U1446 (N_1446,In_586,In_295);
and U1447 (N_1447,In_732,In_431);
nand U1448 (N_1448,In_657,In_396);
or U1449 (N_1449,In_560,In_1535);
nand U1450 (N_1450,In_1582,In_2842);
and U1451 (N_1451,In_1559,In_2838);
and U1452 (N_1452,In_961,In_2720);
or U1453 (N_1453,In_1697,In_55);
or U1454 (N_1454,In_426,In_2614);
nand U1455 (N_1455,In_2621,In_383);
nor U1456 (N_1456,In_780,In_2270);
and U1457 (N_1457,In_1935,In_2566);
or U1458 (N_1458,In_659,In_350);
or U1459 (N_1459,In_2535,In_1667);
nor U1460 (N_1460,In_312,In_610);
nor U1461 (N_1461,In_2552,In_2737);
or U1462 (N_1462,In_667,In_2508);
nor U1463 (N_1463,In_1624,In_2617);
nor U1464 (N_1464,In_1643,In_2398);
xor U1465 (N_1465,In_2375,In_1278);
and U1466 (N_1466,In_1015,In_1830);
nand U1467 (N_1467,In_6,In_2666);
xor U1468 (N_1468,In_2311,In_2648);
or U1469 (N_1469,In_2157,In_2569);
and U1470 (N_1470,In_2709,In_1504);
nor U1471 (N_1471,In_725,In_165);
or U1472 (N_1472,In_2798,In_2214);
and U1473 (N_1473,In_2265,In_911);
xor U1474 (N_1474,In_2714,In_185);
nor U1475 (N_1475,In_1317,In_213);
and U1476 (N_1476,In_1147,In_1023);
and U1477 (N_1477,In_1651,In_1574);
and U1478 (N_1478,In_247,In_950);
nand U1479 (N_1479,In_2482,In_1604);
nand U1480 (N_1480,In_1927,In_1858);
xor U1481 (N_1481,In_2252,In_1880);
nand U1482 (N_1482,In_1164,In_1055);
nand U1483 (N_1483,In_1070,In_1028);
xnor U1484 (N_1484,In_1664,In_2170);
xnor U1485 (N_1485,In_1161,In_231);
nand U1486 (N_1486,In_2590,In_1475);
or U1487 (N_1487,In_150,In_1142);
and U1488 (N_1488,In_116,In_2461);
nor U1489 (N_1489,In_1786,In_2462);
nor U1490 (N_1490,In_664,In_1419);
or U1491 (N_1491,In_2281,In_2628);
nor U1492 (N_1492,In_1433,In_1301);
and U1493 (N_1493,In_320,In_1541);
and U1494 (N_1494,In_1757,In_2003);
nor U1495 (N_1495,In_1238,In_1303);
nor U1496 (N_1496,In_1334,In_1500);
and U1497 (N_1497,In_2751,In_389);
xnor U1498 (N_1498,In_1416,In_1727);
and U1499 (N_1499,In_256,In_2260);
or U1500 (N_1500,In_1190,In_2622);
xnor U1501 (N_1501,In_398,In_155);
and U1502 (N_1502,In_2432,In_2966);
nand U1503 (N_1503,In_2999,In_2731);
or U1504 (N_1504,In_2108,In_1291);
nor U1505 (N_1505,In_1963,In_1058);
and U1506 (N_1506,In_2407,In_1386);
nand U1507 (N_1507,In_419,In_2828);
and U1508 (N_1508,In_2869,In_2266);
or U1509 (N_1509,In_2296,In_370);
nand U1510 (N_1510,In_1562,In_642);
xor U1511 (N_1511,In_114,In_2526);
and U1512 (N_1512,In_976,In_969);
or U1513 (N_1513,In_495,In_2398);
or U1514 (N_1514,In_2319,In_2176);
nand U1515 (N_1515,In_2644,In_1801);
nor U1516 (N_1516,In_2957,In_2080);
nor U1517 (N_1517,In_1864,In_1734);
nand U1518 (N_1518,In_1758,In_674);
nor U1519 (N_1519,In_295,In_1);
and U1520 (N_1520,In_2581,In_1389);
nand U1521 (N_1521,In_325,In_2849);
and U1522 (N_1522,In_787,In_1232);
nand U1523 (N_1523,In_2435,In_1954);
nand U1524 (N_1524,In_872,In_901);
nand U1525 (N_1525,In_2880,In_2912);
nand U1526 (N_1526,In_1914,In_123);
or U1527 (N_1527,In_1990,In_1471);
nand U1528 (N_1528,In_1098,In_1453);
or U1529 (N_1529,In_518,In_347);
or U1530 (N_1530,In_765,In_2243);
and U1531 (N_1531,In_1973,In_2758);
nand U1532 (N_1532,In_2848,In_1489);
or U1533 (N_1533,In_351,In_2605);
or U1534 (N_1534,In_2870,In_1499);
xor U1535 (N_1535,In_126,In_247);
nor U1536 (N_1536,In_228,In_1024);
nand U1537 (N_1537,In_11,In_2681);
nand U1538 (N_1538,In_129,In_1346);
xnor U1539 (N_1539,In_2655,In_2183);
and U1540 (N_1540,In_473,In_2810);
nor U1541 (N_1541,In_758,In_48);
and U1542 (N_1542,In_2997,In_2500);
nor U1543 (N_1543,In_1079,In_1666);
nor U1544 (N_1544,In_872,In_2536);
nor U1545 (N_1545,In_725,In_1548);
and U1546 (N_1546,In_436,In_2380);
and U1547 (N_1547,In_79,In_1410);
and U1548 (N_1548,In_1907,In_1106);
nand U1549 (N_1549,In_2628,In_1914);
and U1550 (N_1550,In_1590,In_548);
or U1551 (N_1551,In_2528,In_398);
nand U1552 (N_1552,In_1818,In_939);
nand U1553 (N_1553,In_710,In_915);
and U1554 (N_1554,In_1230,In_2236);
or U1555 (N_1555,In_2526,In_2760);
nor U1556 (N_1556,In_156,In_1605);
and U1557 (N_1557,In_2959,In_1818);
or U1558 (N_1558,In_548,In_554);
or U1559 (N_1559,In_355,In_1641);
xor U1560 (N_1560,In_2483,In_2121);
or U1561 (N_1561,In_214,In_1306);
nor U1562 (N_1562,In_1341,In_2298);
nor U1563 (N_1563,In_3,In_2571);
xnor U1564 (N_1564,In_494,In_2482);
nand U1565 (N_1565,In_2135,In_487);
nor U1566 (N_1566,In_75,In_2094);
nand U1567 (N_1567,In_2420,In_63);
nand U1568 (N_1568,In_1,In_2258);
or U1569 (N_1569,In_2708,In_1649);
nor U1570 (N_1570,In_176,In_773);
xor U1571 (N_1571,In_2393,In_1693);
and U1572 (N_1572,In_1190,In_2350);
nand U1573 (N_1573,In_1251,In_42);
nand U1574 (N_1574,In_2293,In_1557);
and U1575 (N_1575,In_2404,In_625);
or U1576 (N_1576,In_652,In_2017);
nor U1577 (N_1577,In_347,In_1243);
nand U1578 (N_1578,In_1693,In_884);
or U1579 (N_1579,In_2057,In_1850);
and U1580 (N_1580,In_2834,In_984);
nand U1581 (N_1581,In_899,In_2034);
nor U1582 (N_1582,In_747,In_407);
nand U1583 (N_1583,In_1728,In_730);
nand U1584 (N_1584,In_2814,In_256);
nand U1585 (N_1585,In_2825,In_2094);
nor U1586 (N_1586,In_2647,In_1922);
nand U1587 (N_1587,In_2830,In_2240);
xor U1588 (N_1588,In_294,In_2013);
xor U1589 (N_1589,In_2392,In_1248);
xor U1590 (N_1590,In_734,In_480);
or U1591 (N_1591,In_1944,In_1048);
or U1592 (N_1592,In_1606,In_1201);
nor U1593 (N_1593,In_1366,In_529);
nand U1594 (N_1594,In_1506,In_409);
or U1595 (N_1595,In_2417,In_1056);
nor U1596 (N_1596,In_1690,In_1403);
and U1597 (N_1597,In_713,In_614);
nand U1598 (N_1598,In_2905,In_68);
or U1599 (N_1599,In_2888,In_271);
and U1600 (N_1600,In_2233,In_513);
nor U1601 (N_1601,In_1951,In_1955);
nor U1602 (N_1602,In_617,In_316);
or U1603 (N_1603,In_1548,In_2105);
or U1604 (N_1604,In_2394,In_171);
nor U1605 (N_1605,In_2575,In_1464);
or U1606 (N_1606,In_2901,In_1133);
xnor U1607 (N_1607,In_1318,In_1794);
xnor U1608 (N_1608,In_2524,In_1995);
and U1609 (N_1609,In_9,In_2892);
or U1610 (N_1610,In_2288,In_1893);
nor U1611 (N_1611,In_2085,In_2598);
nor U1612 (N_1612,In_2871,In_2342);
and U1613 (N_1613,In_207,In_1872);
nor U1614 (N_1614,In_2275,In_484);
nand U1615 (N_1615,In_1662,In_144);
or U1616 (N_1616,In_2917,In_2680);
and U1617 (N_1617,In_440,In_667);
nor U1618 (N_1618,In_1681,In_72);
nand U1619 (N_1619,In_726,In_1260);
nand U1620 (N_1620,In_2045,In_970);
nor U1621 (N_1621,In_2688,In_62);
nor U1622 (N_1622,In_730,In_2402);
nor U1623 (N_1623,In_304,In_891);
nor U1624 (N_1624,In_2551,In_22);
nor U1625 (N_1625,In_2703,In_2194);
and U1626 (N_1626,In_1270,In_2671);
nor U1627 (N_1627,In_833,In_1967);
xnor U1628 (N_1628,In_409,In_2835);
nor U1629 (N_1629,In_2852,In_679);
nand U1630 (N_1630,In_1256,In_2267);
or U1631 (N_1631,In_1863,In_2299);
or U1632 (N_1632,In_1907,In_1381);
nand U1633 (N_1633,In_787,In_1408);
nand U1634 (N_1634,In_2524,In_2923);
nand U1635 (N_1635,In_191,In_2131);
or U1636 (N_1636,In_2466,In_587);
or U1637 (N_1637,In_718,In_2757);
and U1638 (N_1638,In_1574,In_600);
nor U1639 (N_1639,In_1064,In_2466);
and U1640 (N_1640,In_32,In_2817);
or U1641 (N_1641,In_1278,In_1905);
and U1642 (N_1642,In_533,In_1637);
and U1643 (N_1643,In_2801,In_495);
or U1644 (N_1644,In_2720,In_2483);
nand U1645 (N_1645,In_1392,In_2239);
and U1646 (N_1646,In_474,In_434);
xor U1647 (N_1647,In_2279,In_1416);
xor U1648 (N_1648,In_2395,In_525);
or U1649 (N_1649,In_2800,In_2034);
nor U1650 (N_1650,In_1156,In_2989);
nand U1651 (N_1651,In_1074,In_1198);
nand U1652 (N_1652,In_1486,In_2761);
nor U1653 (N_1653,In_2778,In_2782);
and U1654 (N_1654,In_1522,In_1503);
and U1655 (N_1655,In_2387,In_1523);
nand U1656 (N_1656,In_2449,In_35);
and U1657 (N_1657,In_2984,In_1513);
nand U1658 (N_1658,In_2000,In_2463);
nand U1659 (N_1659,In_560,In_2070);
nand U1660 (N_1660,In_1122,In_2778);
and U1661 (N_1661,In_1139,In_553);
or U1662 (N_1662,In_783,In_1568);
and U1663 (N_1663,In_1473,In_141);
and U1664 (N_1664,In_843,In_2073);
nor U1665 (N_1665,In_257,In_2395);
nor U1666 (N_1666,In_2285,In_241);
and U1667 (N_1667,In_2248,In_2902);
or U1668 (N_1668,In_819,In_865);
nand U1669 (N_1669,In_2448,In_300);
or U1670 (N_1670,In_274,In_1460);
nor U1671 (N_1671,In_2073,In_2623);
nand U1672 (N_1672,In_2463,In_1239);
and U1673 (N_1673,In_1492,In_203);
nand U1674 (N_1674,In_1173,In_1318);
and U1675 (N_1675,In_2538,In_2972);
or U1676 (N_1676,In_1301,In_2714);
nand U1677 (N_1677,In_766,In_2310);
nand U1678 (N_1678,In_1158,In_922);
xor U1679 (N_1679,In_1056,In_22);
nand U1680 (N_1680,In_2004,In_1983);
or U1681 (N_1681,In_714,In_2463);
or U1682 (N_1682,In_2260,In_2873);
nor U1683 (N_1683,In_2238,In_633);
nor U1684 (N_1684,In_2023,In_2360);
or U1685 (N_1685,In_2845,In_159);
nor U1686 (N_1686,In_2560,In_2637);
and U1687 (N_1687,In_1017,In_1286);
xnor U1688 (N_1688,In_497,In_2121);
or U1689 (N_1689,In_1314,In_2788);
and U1690 (N_1690,In_2464,In_1302);
and U1691 (N_1691,In_2310,In_1519);
or U1692 (N_1692,In_2954,In_1374);
nor U1693 (N_1693,In_752,In_2228);
xnor U1694 (N_1694,In_530,In_2576);
xor U1695 (N_1695,In_2196,In_678);
nor U1696 (N_1696,In_40,In_2672);
nand U1697 (N_1697,In_1937,In_1202);
xnor U1698 (N_1698,In_1875,In_1281);
nand U1699 (N_1699,In_2347,In_1102);
and U1700 (N_1700,In_2563,In_2379);
and U1701 (N_1701,In_2075,In_2711);
and U1702 (N_1702,In_1830,In_1643);
nand U1703 (N_1703,In_1504,In_870);
nand U1704 (N_1704,In_2272,In_150);
and U1705 (N_1705,In_157,In_2305);
nor U1706 (N_1706,In_2248,In_835);
nand U1707 (N_1707,In_2094,In_1902);
or U1708 (N_1708,In_2972,In_1391);
nand U1709 (N_1709,In_2356,In_2970);
nor U1710 (N_1710,In_2001,In_1078);
or U1711 (N_1711,In_868,In_2990);
and U1712 (N_1712,In_564,In_126);
nor U1713 (N_1713,In_1796,In_2186);
nand U1714 (N_1714,In_131,In_2788);
nor U1715 (N_1715,In_1428,In_1859);
or U1716 (N_1716,In_1059,In_2284);
nand U1717 (N_1717,In_2158,In_1632);
xor U1718 (N_1718,In_1019,In_869);
or U1719 (N_1719,In_1608,In_2491);
nor U1720 (N_1720,In_893,In_2752);
and U1721 (N_1721,In_1951,In_2691);
and U1722 (N_1722,In_1767,In_585);
nor U1723 (N_1723,In_2989,In_1460);
or U1724 (N_1724,In_1012,In_2124);
nand U1725 (N_1725,In_2874,In_578);
or U1726 (N_1726,In_749,In_331);
nand U1727 (N_1727,In_2592,In_2479);
or U1728 (N_1728,In_1171,In_1974);
or U1729 (N_1729,In_1375,In_2858);
nand U1730 (N_1730,In_891,In_2623);
and U1731 (N_1731,In_2783,In_2885);
nand U1732 (N_1732,In_2948,In_489);
xor U1733 (N_1733,In_1750,In_1575);
nor U1734 (N_1734,In_2304,In_2242);
nand U1735 (N_1735,In_2002,In_11);
nand U1736 (N_1736,In_1855,In_1701);
nor U1737 (N_1737,In_2937,In_2031);
or U1738 (N_1738,In_2483,In_2729);
nand U1739 (N_1739,In_580,In_984);
nand U1740 (N_1740,In_1490,In_2422);
nor U1741 (N_1741,In_1919,In_2413);
or U1742 (N_1742,In_2449,In_1764);
or U1743 (N_1743,In_97,In_953);
or U1744 (N_1744,In_44,In_2681);
xor U1745 (N_1745,In_2114,In_849);
and U1746 (N_1746,In_1268,In_1027);
nand U1747 (N_1747,In_2893,In_605);
nand U1748 (N_1748,In_1040,In_782);
nor U1749 (N_1749,In_2313,In_2520);
xnor U1750 (N_1750,In_1180,In_438);
nor U1751 (N_1751,In_921,In_1317);
nor U1752 (N_1752,In_1342,In_487);
or U1753 (N_1753,In_1767,In_959);
nor U1754 (N_1754,In_1987,In_1705);
nand U1755 (N_1755,In_2520,In_108);
and U1756 (N_1756,In_2996,In_813);
and U1757 (N_1757,In_135,In_728);
nor U1758 (N_1758,In_1073,In_2138);
or U1759 (N_1759,In_334,In_2186);
or U1760 (N_1760,In_1843,In_2078);
or U1761 (N_1761,In_307,In_2114);
nor U1762 (N_1762,In_1962,In_2514);
and U1763 (N_1763,In_2489,In_602);
or U1764 (N_1764,In_2501,In_2324);
nand U1765 (N_1765,In_348,In_2295);
and U1766 (N_1766,In_1796,In_275);
and U1767 (N_1767,In_2063,In_2245);
nor U1768 (N_1768,In_1519,In_2281);
and U1769 (N_1769,In_944,In_616);
and U1770 (N_1770,In_504,In_2343);
xnor U1771 (N_1771,In_653,In_2214);
nand U1772 (N_1772,In_2869,In_1697);
or U1773 (N_1773,In_1171,In_851);
or U1774 (N_1774,In_265,In_2449);
or U1775 (N_1775,In_461,In_2998);
nand U1776 (N_1776,In_1768,In_2906);
nand U1777 (N_1777,In_1195,In_275);
or U1778 (N_1778,In_319,In_878);
nand U1779 (N_1779,In_2046,In_132);
nand U1780 (N_1780,In_635,In_2541);
or U1781 (N_1781,In_1422,In_1479);
xor U1782 (N_1782,In_2398,In_13);
and U1783 (N_1783,In_2839,In_2774);
or U1784 (N_1784,In_1508,In_2301);
or U1785 (N_1785,In_2950,In_1488);
nand U1786 (N_1786,In_289,In_192);
and U1787 (N_1787,In_62,In_1421);
nand U1788 (N_1788,In_973,In_2244);
or U1789 (N_1789,In_329,In_461);
nor U1790 (N_1790,In_682,In_1624);
and U1791 (N_1791,In_672,In_2832);
nand U1792 (N_1792,In_1097,In_203);
xor U1793 (N_1793,In_1939,In_1972);
or U1794 (N_1794,In_1162,In_2538);
nor U1795 (N_1795,In_2364,In_290);
or U1796 (N_1796,In_2974,In_1620);
nand U1797 (N_1797,In_2073,In_1656);
and U1798 (N_1798,In_1402,In_1652);
and U1799 (N_1799,In_1965,In_1570);
or U1800 (N_1800,In_2365,In_1267);
nand U1801 (N_1801,In_2505,In_2202);
nor U1802 (N_1802,In_1450,In_585);
or U1803 (N_1803,In_1131,In_2621);
nand U1804 (N_1804,In_155,In_1487);
and U1805 (N_1805,In_1222,In_1529);
nor U1806 (N_1806,In_1844,In_1309);
nor U1807 (N_1807,In_2454,In_2136);
nor U1808 (N_1808,In_2329,In_917);
nand U1809 (N_1809,In_242,In_2708);
nand U1810 (N_1810,In_2685,In_818);
xor U1811 (N_1811,In_2856,In_2117);
nand U1812 (N_1812,In_2142,In_2968);
or U1813 (N_1813,In_244,In_1373);
and U1814 (N_1814,In_2312,In_2614);
nand U1815 (N_1815,In_1589,In_1568);
nor U1816 (N_1816,In_89,In_2274);
or U1817 (N_1817,In_2857,In_1851);
and U1818 (N_1818,In_161,In_285);
and U1819 (N_1819,In_1334,In_327);
and U1820 (N_1820,In_1717,In_2070);
xnor U1821 (N_1821,In_2312,In_695);
nor U1822 (N_1822,In_1056,In_1589);
or U1823 (N_1823,In_2024,In_2742);
nand U1824 (N_1824,In_2534,In_1413);
or U1825 (N_1825,In_396,In_1893);
or U1826 (N_1826,In_1009,In_1631);
nor U1827 (N_1827,In_817,In_32);
nand U1828 (N_1828,In_973,In_2489);
nand U1829 (N_1829,In_1779,In_1855);
nor U1830 (N_1830,In_516,In_597);
nand U1831 (N_1831,In_421,In_132);
or U1832 (N_1832,In_322,In_2212);
and U1833 (N_1833,In_704,In_2704);
nor U1834 (N_1834,In_1490,In_609);
or U1835 (N_1835,In_1269,In_1564);
or U1836 (N_1836,In_896,In_2296);
and U1837 (N_1837,In_1629,In_306);
xnor U1838 (N_1838,In_2801,In_2719);
or U1839 (N_1839,In_725,In_1634);
or U1840 (N_1840,In_979,In_2677);
nor U1841 (N_1841,In_616,In_1409);
nand U1842 (N_1842,In_2620,In_1478);
or U1843 (N_1843,In_1773,In_1673);
or U1844 (N_1844,In_198,In_920);
and U1845 (N_1845,In_1476,In_2262);
or U1846 (N_1846,In_930,In_2613);
nor U1847 (N_1847,In_2771,In_2894);
nand U1848 (N_1848,In_2063,In_2614);
nor U1849 (N_1849,In_2873,In_2943);
or U1850 (N_1850,In_1567,In_2667);
and U1851 (N_1851,In_1467,In_834);
and U1852 (N_1852,In_2957,In_2969);
or U1853 (N_1853,In_228,In_4);
or U1854 (N_1854,In_109,In_2349);
nand U1855 (N_1855,In_2835,In_373);
or U1856 (N_1856,In_367,In_2096);
and U1857 (N_1857,In_1232,In_253);
and U1858 (N_1858,In_1955,In_1172);
nor U1859 (N_1859,In_1592,In_73);
and U1860 (N_1860,In_2421,In_257);
and U1861 (N_1861,In_1549,In_756);
nor U1862 (N_1862,In_438,In_2560);
nand U1863 (N_1863,In_1832,In_24);
nand U1864 (N_1864,In_2586,In_159);
nor U1865 (N_1865,In_908,In_91);
nand U1866 (N_1866,In_1275,In_2115);
and U1867 (N_1867,In_627,In_2282);
nand U1868 (N_1868,In_2249,In_2166);
and U1869 (N_1869,In_2303,In_2378);
nor U1870 (N_1870,In_1071,In_1670);
and U1871 (N_1871,In_2694,In_2534);
or U1872 (N_1872,In_839,In_620);
or U1873 (N_1873,In_509,In_887);
or U1874 (N_1874,In_113,In_2398);
and U1875 (N_1875,In_1295,In_364);
xor U1876 (N_1876,In_1895,In_1030);
nand U1877 (N_1877,In_395,In_1433);
nand U1878 (N_1878,In_634,In_1055);
nor U1879 (N_1879,In_1623,In_477);
xor U1880 (N_1880,In_1672,In_1852);
and U1881 (N_1881,In_898,In_1486);
nand U1882 (N_1882,In_1308,In_308);
nor U1883 (N_1883,In_862,In_393);
xnor U1884 (N_1884,In_1543,In_2316);
and U1885 (N_1885,In_2792,In_296);
or U1886 (N_1886,In_865,In_2974);
nor U1887 (N_1887,In_1442,In_1699);
nand U1888 (N_1888,In_2997,In_669);
xor U1889 (N_1889,In_652,In_2639);
and U1890 (N_1890,In_1999,In_727);
nor U1891 (N_1891,In_49,In_1750);
xor U1892 (N_1892,In_2528,In_160);
nand U1893 (N_1893,In_620,In_586);
and U1894 (N_1894,In_1269,In_2304);
xor U1895 (N_1895,In_395,In_2605);
nor U1896 (N_1896,In_1426,In_2649);
or U1897 (N_1897,In_2915,In_71);
nor U1898 (N_1898,In_2366,In_2518);
or U1899 (N_1899,In_1327,In_227);
nand U1900 (N_1900,In_1912,In_33);
nor U1901 (N_1901,In_411,In_1575);
nor U1902 (N_1902,In_1144,In_2611);
nor U1903 (N_1903,In_940,In_2675);
nor U1904 (N_1904,In_2840,In_1669);
nand U1905 (N_1905,In_1807,In_2183);
nand U1906 (N_1906,In_121,In_600);
or U1907 (N_1907,In_653,In_2726);
and U1908 (N_1908,In_1384,In_2874);
nand U1909 (N_1909,In_90,In_2645);
nor U1910 (N_1910,In_2490,In_2654);
and U1911 (N_1911,In_1573,In_856);
nor U1912 (N_1912,In_387,In_2128);
and U1913 (N_1913,In_1417,In_2196);
nor U1914 (N_1914,In_2975,In_1423);
and U1915 (N_1915,In_1837,In_1913);
nor U1916 (N_1916,In_1707,In_1923);
or U1917 (N_1917,In_2187,In_1462);
or U1918 (N_1918,In_2932,In_2750);
or U1919 (N_1919,In_346,In_549);
nand U1920 (N_1920,In_1585,In_2985);
and U1921 (N_1921,In_1063,In_964);
and U1922 (N_1922,In_2465,In_1391);
nor U1923 (N_1923,In_2345,In_1514);
nand U1924 (N_1924,In_806,In_1702);
nor U1925 (N_1925,In_173,In_2737);
nor U1926 (N_1926,In_533,In_2110);
nand U1927 (N_1927,In_2173,In_2509);
and U1928 (N_1928,In_1326,In_853);
xor U1929 (N_1929,In_2952,In_2121);
nand U1930 (N_1930,In_2822,In_2830);
nand U1931 (N_1931,In_2809,In_1875);
and U1932 (N_1932,In_1335,In_1883);
xnor U1933 (N_1933,In_1192,In_425);
nand U1934 (N_1934,In_2277,In_2649);
nand U1935 (N_1935,In_1175,In_2890);
nor U1936 (N_1936,In_215,In_387);
xor U1937 (N_1937,In_1844,In_2748);
nor U1938 (N_1938,In_767,In_168);
or U1939 (N_1939,In_1383,In_913);
nor U1940 (N_1940,In_1889,In_2529);
nor U1941 (N_1941,In_2436,In_364);
nor U1942 (N_1942,In_2522,In_852);
nor U1943 (N_1943,In_2301,In_665);
nand U1944 (N_1944,In_1049,In_340);
nor U1945 (N_1945,In_1719,In_939);
nor U1946 (N_1946,In_1444,In_2194);
nand U1947 (N_1947,In_1275,In_1748);
and U1948 (N_1948,In_172,In_632);
nor U1949 (N_1949,In_1479,In_2172);
or U1950 (N_1950,In_1808,In_1177);
and U1951 (N_1951,In_601,In_994);
and U1952 (N_1952,In_2109,In_2857);
and U1953 (N_1953,In_1688,In_694);
or U1954 (N_1954,In_88,In_1915);
nor U1955 (N_1955,In_2879,In_2597);
nor U1956 (N_1956,In_1420,In_1848);
nand U1957 (N_1957,In_2574,In_1040);
xor U1958 (N_1958,In_2747,In_491);
nand U1959 (N_1959,In_1283,In_2785);
nand U1960 (N_1960,In_1732,In_619);
nand U1961 (N_1961,In_2067,In_2063);
nand U1962 (N_1962,In_429,In_2619);
nor U1963 (N_1963,In_2103,In_2622);
nor U1964 (N_1964,In_1641,In_1518);
or U1965 (N_1965,In_1152,In_1885);
nand U1966 (N_1966,In_1156,In_73);
or U1967 (N_1967,In_2434,In_222);
xnor U1968 (N_1968,In_1251,In_2281);
nand U1969 (N_1969,In_1856,In_1879);
nand U1970 (N_1970,In_2651,In_2232);
nand U1971 (N_1971,In_466,In_864);
or U1972 (N_1972,In_621,In_2888);
nand U1973 (N_1973,In_794,In_2540);
or U1974 (N_1974,In_977,In_2009);
and U1975 (N_1975,In_2526,In_2755);
nand U1976 (N_1976,In_2312,In_395);
and U1977 (N_1977,In_2086,In_31);
xnor U1978 (N_1978,In_956,In_559);
nor U1979 (N_1979,In_2547,In_102);
xor U1980 (N_1980,In_1841,In_2525);
nand U1981 (N_1981,In_2079,In_1194);
nor U1982 (N_1982,In_1494,In_2772);
xnor U1983 (N_1983,In_1271,In_2015);
and U1984 (N_1984,In_122,In_1728);
and U1985 (N_1985,In_2658,In_284);
nor U1986 (N_1986,In_248,In_1632);
or U1987 (N_1987,In_2982,In_2697);
nand U1988 (N_1988,In_685,In_1289);
nor U1989 (N_1989,In_109,In_592);
nand U1990 (N_1990,In_1645,In_345);
and U1991 (N_1991,In_718,In_786);
or U1992 (N_1992,In_2531,In_1601);
nor U1993 (N_1993,In_752,In_2634);
or U1994 (N_1994,In_2792,In_734);
or U1995 (N_1995,In_840,In_1024);
nand U1996 (N_1996,In_2114,In_1396);
or U1997 (N_1997,In_2967,In_2608);
nand U1998 (N_1998,In_2369,In_2749);
and U1999 (N_1999,In_1881,In_1132);
nor U2000 (N_2000,In_2641,In_2584);
nand U2001 (N_2001,In_334,In_1794);
and U2002 (N_2002,In_1465,In_2439);
nand U2003 (N_2003,In_102,In_2453);
xnor U2004 (N_2004,In_571,In_607);
and U2005 (N_2005,In_916,In_1439);
or U2006 (N_2006,In_776,In_1454);
nor U2007 (N_2007,In_2294,In_1438);
nor U2008 (N_2008,In_2977,In_2642);
or U2009 (N_2009,In_2260,In_2369);
nor U2010 (N_2010,In_2304,In_2490);
nor U2011 (N_2011,In_2774,In_1825);
nor U2012 (N_2012,In_1670,In_169);
nor U2013 (N_2013,In_2532,In_802);
or U2014 (N_2014,In_222,In_2719);
and U2015 (N_2015,In_876,In_2924);
or U2016 (N_2016,In_2151,In_2610);
nor U2017 (N_2017,In_728,In_2676);
and U2018 (N_2018,In_2904,In_119);
nand U2019 (N_2019,In_2535,In_563);
or U2020 (N_2020,In_897,In_2727);
and U2021 (N_2021,In_2271,In_2212);
and U2022 (N_2022,In_1430,In_139);
nand U2023 (N_2023,In_866,In_638);
nor U2024 (N_2024,In_80,In_951);
nand U2025 (N_2025,In_210,In_1709);
and U2026 (N_2026,In_2744,In_1026);
or U2027 (N_2027,In_204,In_2095);
or U2028 (N_2028,In_2686,In_25);
xnor U2029 (N_2029,In_671,In_1383);
xor U2030 (N_2030,In_1095,In_2545);
nor U2031 (N_2031,In_305,In_833);
and U2032 (N_2032,In_1161,In_568);
nor U2033 (N_2033,In_497,In_482);
nand U2034 (N_2034,In_941,In_583);
nor U2035 (N_2035,In_825,In_1730);
or U2036 (N_2036,In_2910,In_2950);
nand U2037 (N_2037,In_163,In_2833);
nor U2038 (N_2038,In_666,In_2419);
nor U2039 (N_2039,In_2934,In_307);
and U2040 (N_2040,In_2434,In_2400);
nor U2041 (N_2041,In_864,In_843);
or U2042 (N_2042,In_736,In_557);
and U2043 (N_2043,In_1627,In_1939);
nor U2044 (N_2044,In_472,In_1433);
nor U2045 (N_2045,In_1679,In_1620);
or U2046 (N_2046,In_2042,In_1594);
and U2047 (N_2047,In_226,In_898);
and U2048 (N_2048,In_2434,In_643);
or U2049 (N_2049,In_2398,In_672);
or U2050 (N_2050,In_158,In_911);
and U2051 (N_2051,In_1761,In_374);
nor U2052 (N_2052,In_2588,In_2861);
xnor U2053 (N_2053,In_1883,In_1005);
nand U2054 (N_2054,In_1690,In_481);
or U2055 (N_2055,In_2689,In_1181);
nor U2056 (N_2056,In_1398,In_814);
or U2057 (N_2057,In_2305,In_1356);
and U2058 (N_2058,In_1103,In_1631);
or U2059 (N_2059,In_1393,In_833);
or U2060 (N_2060,In_554,In_656);
or U2061 (N_2061,In_159,In_2532);
nor U2062 (N_2062,In_2605,In_83);
nor U2063 (N_2063,In_676,In_2965);
and U2064 (N_2064,In_1461,In_2421);
and U2065 (N_2065,In_1149,In_106);
nor U2066 (N_2066,In_530,In_2445);
or U2067 (N_2067,In_1208,In_1297);
and U2068 (N_2068,In_834,In_1182);
nand U2069 (N_2069,In_2992,In_1815);
nand U2070 (N_2070,In_2588,In_2806);
and U2071 (N_2071,In_2448,In_2571);
or U2072 (N_2072,In_2548,In_2414);
nand U2073 (N_2073,In_2597,In_2834);
nor U2074 (N_2074,In_1380,In_2262);
and U2075 (N_2075,In_661,In_2048);
xor U2076 (N_2076,In_2808,In_2287);
or U2077 (N_2077,In_2148,In_1235);
or U2078 (N_2078,In_618,In_1216);
nor U2079 (N_2079,In_2429,In_818);
nor U2080 (N_2080,In_1477,In_2744);
nor U2081 (N_2081,In_1422,In_2538);
nand U2082 (N_2082,In_1349,In_2578);
xnor U2083 (N_2083,In_216,In_2520);
xnor U2084 (N_2084,In_512,In_1039);
nand U2085 (N_2085,In_1490,In_185);
or U2086 (N_2086,In_2613,In_1620);
nand U2087 (N_2087,In_1390,In_1459);
and U2088 (N_2088,In_1653,In_2524);
nor U2089 (N_2089,In_1981,In_1558);
and U2090 (N_2090,In_2607,In_1142);
and U2091 (N_2091,In_2797,In_1557);
or U2092 (N_2092,In_781,In_2302);
nor U2093 (N_2093,In_2690,In_988);
nand U2094 (N_2094,In_1373,In_1276);
or U2095 (N_2095,In_1012,In_1652);
nand U2096 (N_2096,In_1157,In_188);
nand U2097 (N_2097,In_2862,In_609);
nor U2098 (N_2098,In_2123,In_1704);
nor U2099 (N_2099,In_1986,In_372);
nand U2100 (N_2100,In_329,In_1258);
xnor U2101 (N_2101,In_773,In_1535);
and U2102 (N_2102,In_345,In_2415);
nand U2103 (N_2103,In_1117,In_881);
and U2104 (N_2104,In_455,In_804);
nor U2105 (N_2105,In_1266,In_1398);
xor U2106 (N_2106,In_564,In_2643);
xnor U2107 (N_2107,In_1114,In_772);
and U2108 (N_2108,In_2218,In_1842);
nand U2109 (N_2109,In_1125,In_449);
nor U2110 (N_2110,In_2714,In_47);
or U2111 (N_2111,In_1872,In_708);
nand U2112 (N_2112,In_826,In_2587);
nor U2113 (N_2113,In_1313,In_2875);
and U2114 (N_2114,In_131,In_2556);
nand U2115 (N_2115,In_855,In_1619);
or U2116 (N_2116,In_144,In_2461);
nor U2117 (N_2117,In_630,In_1150);
nor U2118 (N_2118,In_2493,In_1528);
nand U2119 (N_2119,In_1365,In_186);
nand U2120 (N_2120,In_1875,In_1965);
or U2121 (N_2121,In_1979,In_2562);
xor U2122 (N_2122,In_1074,In_805);
nand U2123 (N_2123,In_2157,In_2510);
nand U2124 (N_2124,In_1903,In_88);
and U2125 (N_2125,In_2121,In_1869);
or U2126 (N_2126,In_2879,In_2996);
and U2127 (N_2127,In_2520,In_357);
or U2128 (N_2128,In_2502,In_946);
and U2129 (N_2129,In_2561,In_751);
or U2130 (N_2130,In_413,In_1649);
nand U2131 (N_2131,In_2854,In_1597);
nor U2132 (N_2132,In_704,In_1925);
or U2133 (N_2133,In_2002,In_339);
nor U2134 (N_2134,In_107,In_2780);
and U2135 (N_2135,In_635,In_2654);
xnor U2136 (N_2136,In_185,In_400);
nand U2137 (N_2137,In_48,In_2337);
or U2138 (N_2138,In_2704,In_1308);
or U2139 (N_2139,In_1334,In_1010);
and U2140 (N_2140,In_1812,In_2758);
nand U2141 (N_2141,In_1887,In_2527);
xnor U2142 (N_2142,In_2680,In_2618);
nor U2143 (N_2143,In_2846,In_1205);
or U2144 (N_2144,In_2961,In_1208);
or U2145 (N_2145,In_2656,In_305);
or U2146 (N_2146,In_358,In_91);
nor U2147 (N_2147,In_2975,In_1851);
xnor U2148 (N_2148,In_2682,In_550);
and U2149 (N_2149,In_2056,In_2563);
xnor U2150 (N_2150,In_1206,In_2286);
xnor U2151 (N_2151,In_262,In_1842);
xor U2152 (N_2152,In_2226,In_2914);
or U2153 (N_2153,In_1139,In_1367);
and U2154 (N_2154,In_1591,In_691);
and U2155 (N_2155,In_873,In_1388);
nand U2156 (N_2156,In_1834,In_1365);
xnor U2157 (N_2157,In_615,In_2916);
and U2158 (N_2158,In_1385,In_312);
nor U2159 (N_2159,In_787,In_1439);
nand U2160 (N_2160,In_977,In_686);
or U2161 (N_2161,In_1029,In_1348);
nand U2162 (N_2162,In_2010,In_2566);
and U2163 (N_2163,In_230,In_2038);
nor U2164 (N_2164,In_1931,In_1372);
or U2165 (N_2165,In_648,In_351);
nor U2166 (N_2166,In_1286,In_2216);
or U2167 (N_2167,In_1190,In_396);
and U2168 (N_2168,In_2129,In_1229);
xor U2169 (N_2169,In_1467,In_1389);
xnor U2170 (N_2170,In_888,In_991);
and U2171 (N_2171,In_2335,In_2555);
or U2172 (N_2172,In_836,In_450);
nor U2173 (N_2173,In_463,In_592);
xor U2174 (N_2174,In_672,In_2042);
xnor U2175 (N_2175,In_1742,In_382);
and U2176 (N_2176,In_1578,In_772);
nand U2177 (N_2177,In_346,In_1377);
nand U2178 (N_2178,In_2253,In_2154);
nand U2179 (N_2179,In_2490,In_2231);
nand U2180 (N_2180,In_2887,In_2215);
nand U2181 (N_2181,In_2854,In_2406);
and U2182 (N_2182,In_1330,In_381);
or U2183 (N_2183,In_1372,In_1588);
nand U2184 (N_2184,In_1872,In_2707);
nand U2185 (N_2185,In_1480,In_1375);
nand U2186 (N_2186,In_318,In_247);
nor U2187 (N_2187,In_93,In_1197);
nand U2188 (N_2188,In_1986,In_1959);
and U2189 (N_2189,In_1110,In_2966);
or U2190 (N_2190,In_1376,In_778);
xor U2191 (N_2191,In_1538,In_660);
nor U2192 (N_2192,In_2127,In_225);
and U2193 (N_2193,In_869,In_1050);
xor U2194 (N_2194,In_2152,In_1475);
nor U2195 (N_2195,In_449,In_782);
and U2196 (N_2196,In_1093,In_731);
nor U2197 (N_2197,In_1919,In_2700);
nand U2198 (N_2198,In_1772,In_954);
or U2199 (N_2199,In_1596,In_287);
or U2200 (N_2200,In_446,In_2158);
and U2201 (N_2201,In_829,In_1672);
and U2202 (N_2202,In_1741,In_2823);
xor U2203 (N_2203,In_438,In_2129);
nor U2204 (N_2204,In_583,In_2802);
or U2205 (N_2205,In_76,In_2268);
nand U2206 (N_2206,In_1612,In_945);
nor U2207 (N_2207,In_889,In_2313);
and U2208 (N_2208,In_2978,In_596);
nand U2209 (N_2209,In_2758,In_57);
nor U2210 (N_2210,In_996,In_1248);
xor U2211 (N_2211,In_636,In_2357);
nand U2212 (N_2212,In_604,In_2100);
nand U2213 (N_2213,In_447,In_2155);
nand U2214 (N_2214,In_1443,In_206);
nand U2215 (N_2215,In_2238,In_415);
or U2216 (N_2216,In_36,In_2750);
and U2217 (N_2217,In_2014,In_339);
and U2218 (N_2218,In_2362,In_649);
nor U2219 (N_2219,In_1332,In_1560);
xor U2220 (N_2220,In_1204,In_1533);
xnor U2221 (N_2221,In_779,In_1874);
nor U2222 (N_2222,In_838,In_2618);
xnor U2223 (N_2223,In_95,In_1140);
nor U2224 (N_2224,In_1146,In_284);
and U2225 (N_2225,In_1653,In_697);
and U2226 (N_2226,In_2367,In_300);
and U2227 (N_2227,In_2104,In_1800);
and U2228 (N_2228,In_2984,In_1721);
nand U2229 (N_2229,In_1942,In_1150);
or U2230 (N_2230,In_1885,In_1999);
and U2231 (N_2231,In_2400,In_2983);
and U2232 (N_2232,In_2186,In_2346);
or U2233 (N_2233,In_1285,In_544);
and U2234 (N_2234,In_2047,In_419);
and U2235 (N_2235,In_1770,In_2181);
and U2236 (N_2236,In_58,In_2965);
and U2237 (N_2237,In_1236,In_1988);
and U2238 (N_2238,In_1921,In_2712);
or U2239 (N_2239,In_2887,In_1814);
nor U2240 (N_2240,In_599,In_1885);
nor U2241 (N_2241,In_891,In_2038);
nand U2242 (N_2242,In_296,In_2295);
or U2243 (N_2243,In_881,In_2228);
nor U2244 (N_2244,In_900,In_304);
nor U2245 (N_2245,In_686,In_1393);
nor U2246 (N_2246,In_1023,In_2352);
and U2247 (N_2247,In_990,In_2337);
xor U2248 (N_2248,In_2905,In_2431);
or U2249 (N_2249,In_2453,In_2545);
and U2250 (N_2250,In_1241,In_847);
or U2251 (N_2251,In_1223,In_2674);
and U2252 (N_2252,In_2814,In_63);
nor U2253 (N_2253,In_2628,In_2262);
nor U2254 (N_2254,In_1795,In_2676);
and U2255 (N_2255,In_1863,In_787);
xnor U2256 (N_2256,In_798,In_338);
nand U2257 (N_2257,In_599,In_1302);
nor U2258 (N_2258,In_500,In_1331);
and U2259 (N_2259,In_548,In_830);
and U2260 (N_2260,In_2113,In_1188);
nor U2261 (N_2261,In_432,In_317);
and U2262 (N_2262,In_367,In_2076);
nand U2263 (N_2263,In_1333,In_2992);
xnor U2264 (N_2264,In_2384,In_808);
or U2265 (N_2265,In_824,In_2220);
nand U2266 (N_2266,In_2153,In_2437);
and U2267 (N_2267,In_1158,In_1864);
nand U2268 (N_2268,In_1428,In_874);
and U2269 (N_2269,In_682,In_1246);
or U2270 (N_2270,In_2681,In_1177);
xnor U2271 (N_2271,In_833,In_2092);
and U2272 (N_2272,In_625,In_290);
xor U2273 (N_2273,In_2876,In_2479);
and U2274 (N_2274,In_360,In_1129);
nor U2275 (N_2275,In_84,In_2697);
nor U2276 (N_2276,In_929,In_2054);
or U2277 (N_2277,In_72,In_1111);
nand U2278 (N_2278,In_363,In_2535);
and U2279 (N_2279,In_2519,In_1907);
or U2280 (N_2280,In_2809,In_1565);
and U2281 (N_2281,In_1275,In_2261);
or U2282 (N_2282,In_480,In_1666);
nor U2283 (N_2283,In_146,In_2987);
nor U2284 (N_2284,In_2401,In_2292);
nand U2285 (N_2285,In_1586,In_1985);
or U2286 (N_2286,In_1969,In_2433);
nor U2287 (N_2287,In_1911,In_982);
nor U2288 (N_2288,In_1489,In_40);
and U2289 (N_2289,In_754,In_1560);
or U2290 (N_2290,In_1819,In_1477);
xor U2291 (N_2291,In_678,In_732);
and U2292 (N_2292,In_1915,In_232);
nand U2293 (N_2293,In_1725,In_1164);
nor U2294 (N_2294,In_30,In_1859);
nor U2295 (N_2295,In_1600,In_2322);
and U2296 (N_2296,In_611,In_2671);
nand U2297 (N_2297,In_1503,In_2624);
nor U2298 (N_2298,In_73,In_2332);
nor U2299 (N_2299,In_2969,In_2091);
nand U2300 (N_2300,In_2165,In_740);
or U2301 (N_2301,In_331,In_1518);
or U2302 (N_2302,In_2639,In_289);
and U2303 (N_2303,In_909,In_1631);
and U2304 (N_2304,In_588,In_1726);
nand U2305 (N_2305,In_127,In_1051);
and U2306 (N_2306,In_325,In_158);
nand U2307 (N_2307,In_2266,In_2382);
or U2308 (N_2308,In_67,In_1497);
or U2309 (N_2309,In_2275,In_2303);
nand U2310 (N_2310,In_851,In_1558);
and U2311 (N_2311,In_1220,In_2952);
nand U2312 (N_2312,In_1725,In_2113);
nor U2313 (N_2313,In_2872,In_2658);
nor U2314 (N_2314,In_123,In_931);
nor U2315 (N_2315,In_417,In_1311);
or U2316 (N_2316,In_1471,In_311);
nor U2317 (N_2317,In_1909,In_1275);
or U2318 (N_2318,In_2839,In_2815);
xnor U2319 (N_2319,In_263,In_486);
or U2320 (N_2320,In_1821,In_2377);
xnor U2321 (N_2321,In_1785,In_1698);
nand U2322 (N_2322,In_1998,In_1759);
or U2323 (N_2323,In_1521,In_282);
or U2324 (N_2324,In_2743,In_1203);
xnor U2325 (N_2325,In_593,In_207);
and U2326 (N_2326,In_1293,In_627);
or U2327 (N_2327,In_2002,In_2404);
nand U2328 (N_2328,In_721,In_1473);
or U2329 (N_2329,In_2769,In_2100);
xnor U2330 (N_2330,In_2301,In_787);
nand U2331 (N_2331,In_2565,In_2745);
nand U2332 (N_2332,In_844,In_2874);
nand U2333 (N_2333,In_693,In_881);
nor U2334 (N_2334,In_1065,In_487);
nor U2335 (N_2335,In_2027,In_711);
nor U2336 (N_2336,In_1712,In_629);
nand U2337 (N_2337,In_481,In_2181);
or U2338 (N_2338,In_1996,In_1695);
nand U2339 (N_2339,In_1036,In_2569);
nand U2340 (N_2340,In_1274,In_2667);
or U2341 (N_2341,In_2454,In_69);
and U2342 (N_2342,In_292,In_1073);
nor U2343 (N_2343,In_2158,In_1014);
xor U2344 (N_2344,In_2217,In_1762);
xor U2345 (N_2345,In_1808,In_2319);
or U2346 (N_2346,In_819,In_1105);
nor U2347 (N_2347,In_208,In_854);
and U2348 (N_2348,In_2663,In_810);
and U2349 (N_2349,In_1852,In_2697);
and U2350 (N_2350,In_2353,In_2605);
nand U2351 (N_2351,In_329,In_568);
nor U2352 (N_2352,In_33,In_2490);
nand U2353 (N_2353,In_2457,In_1388);
and U2354 (N_2354,In_469,In_1240);
nor U2355 (N_2355,In_1586,In_420);
and U2356 (N_2356,In_1528,In_1222);
nor U2357 (N_2357,In_1857,In_1627);
nand U2358 (N_2358,In_1214,In_95);
nor U2359 (N_2359,In_935,In_2497);
or U2360 (N_2360,In_472,In_1023);
and U2361 (N_2361,In_387,In_878);
and U2362 (N_2362,In_331,In_935);
or U2363 (N_2363,In_309,In_82);
nor U2364 (N_2364,In_2327,In_2886);
nand U2365 (N_2365,In_1786,In_766);
nor U2366 (N_2366,In_51,In_673);
xor U2367 (N_2367,In_357,In_66);
nand U2368 (N_2368,In_73,In_1784);
xor U2369 (N_2369,In_2671,In_1786);
or U2370 (N_2370,In_774,In_2517);
nor U2371 (N_2371,In_2116,In_912);
nor U2372 (N_2372,In_277,In_2719);
nand U2373 (N_2373,In_1172,In_2900);
and U2374 (N_2374,In_2448,In_2693);
xnor U2375 (N_2375,In_1751,In_647);
and U2376 (N_2376,In_1942,In_365);
and U2377 (N_2377,In_1256,In_591);
and U2378 (N_2378,In_1723,In_1725);
nand U2379 (N_2379,In_1866,In_405);
xnor U2380 (N_2380,In_2334,In_2097);
xnor U2381 (N_2381,In_2114,In_1221);
or U2382 (N_2382,In_1349,In_1770);
nor U2383 (N_2383,In_2444,In_2714);
or U2384 (N_2384,In_2081,In_2981);
or U2385 (N_2385,In_246,In_50);
nand U2386 (N_2386,In_1489,In_703);
nor U2387 (N_2387,In_2863,In_2015);
nor U2388 (N_2388,In_1307,In_1028);
nor U2389 (N_2389,In_2842,In_2419);
nor U2390 (N_2390,In_1450,In_199);
nor U2391 (N_2391,In_1226,In_1690);
nor U2392 (N_2392,In_2462,In_645);
nor U2393 (N_2393,In_2494,In_1146);
nor U2394 (N_2394,In_495,In_1191);
nand U2395 (N_2395,In_2281,In_393);
nor U2396 (N_2396,In_1170,In_1429);
xnor U2397 (N_2397,In_914,In_1197);
xor U2398 (N_2398,In_2219,In_46);
nand U2399 (N_2399,In_2787,In_446);
or U2400 (N_2400,In_269,In_1139);
or U2401 (N_2401,In_221,In_74);
xnor U2402 (N_2402,In_1801,In_2796);
nand U2403 (N_2403,In_366,In_2270);
and U2404 (N_2404,In_121,In_1948);
nand U2405 (N_2405,In_138,In_611);
and U2406 (N_2406,In_2228,In_671);
or U2407 (N_2407,In_1196,In_745);
or U2408 (N_2408,In_2613,In_2875);
nor U2409 (N_2409,In_1040,In_2079);
and U2410 (N_2410,In_2652,In_930);
and U2411 (N_2411,In_174,In_2024);
nor U2412 (N_2412,In_2643,In_821);
nor U2413 (N_2413,In_2863,In_1320);
or U2414 (N_2414,In_306,In_2645);
nor U2415 (N_2415,In_1109,In_1219);
nor U2416 (N_2416,In_2512,In_2285);
or U2417 (N_2417,In_299,In_1924);
nand U2418 (N_2418,In_1075,In_1266);
nand U2419 (N_2419,In_1750,In_1846);
and U2420 (N_2420,In_1138,In_2594);
or U2421 (N_2421,In_2037,In_2399);
nor U2422 (N_2422,In_1195,In_1062);
nor U2423 (N_2423,In_1560,In_1830);
and U2424 (N_2424,In_1579,In_2572);
nor U2425 (N_2425,In_980,In_1773);
nand U2426 (N_2426,In_2668,In_1773);
nand U2427 (N_2427,In_781,In_641);
nor U2428 (N_2428,In_1821,In_60);
or U2429 (N_2429,In_818,In_1344);
nor U2430 (N_2430,In_234,In_1825);
or U2431 (N_2431,In_2984,In_27);
nor U2432 (N_2432,In_1396,In_2340);
and U2433 (N_2433,In_1127,In_2942);
nand U2434 (N_2434,In_568,In_2629);
and U2435 (N_2435,In_82,In_2321);
xor U2436 (N_2436,In_1917,In_1176);
nand U2437 (N_2437,In_453,In_202);
or U2438 (N_2438,In_2846,In_660);
and U2439 (N_2439,In_2490,In_2315);
xor U2440 (N_2440,In_2614,In_929);
or U2441 (N_2441,In_786,In_2224);
nor U2442 (N_2442,In_47,In_613);
and U2443 (N_2443,In_952,In_1195);
xor U2444 (N_2444,In_198,In_2765);
and U2445 (N_2445,In_378,In_2479);
and U2446 (N_2446,In_2482,In_631);
nor U2447 (N_2447,In_2109,In_2909);
nand U2448 (N_2448,In_367,In_2392);
nand U2449 (N_2449,In_1557,In_751);
or U2450 (N_2450,In_2479,In_2000);
nand U2451 (N_2451,In_2981,In_2008);
nor U2452 (N_2452,In_2919,In_1701);
or U2453 (N_2453,In_2173,In_392);
nand U2454 (N_2454,In_2596,In_595);
and U2455 (N_2455,In_2119,In_1799);
or U2456 (N_2456,In_1426,In_2607);
nand U2457 (N_2457,In_1267,In_1967);
and U2458 (N_2458,In_567,In_814);
nand U2459 (N_2459,In_445,In_441);
nand U2460 (N_2460,In_803,In_1754);
nand U2461 (N_2461,In_98,In_1980);
or U2462 (N_2462,In_608,In_1335);
nor U2463 (N_2463,In_2396,In_1077);
and U2464 (N_2464,In_2339,In_1584);
nor U2465 (N_2465,In_641,In_2843);
nand U2466 (N_2466,In_467,In_1925);
or U2467 (N_2467,In_859,In_1612);
nor U2468 (N_2468,In_2752,In_1128);
nor U2469 (N_2469,In_767,In_2278);
and U2470 (N_2470,In_1827,In_2301);
xnor U2471 (N_2471,In_2540,In_2877);
or U2472 (N_2472,In_900,In_2996);
nor U2473 (N_2473,In_2186,In_2287);
or U2474 (N_2474,In_1261,In_2424);
nor U2475 (N_2475,In_966,In_1490);
nand U2476 (N_2476,In_607,In_2533);
nor U2477 (N_2477,In_1434,In_1914);
nor U2478 (N_2478,In_91,In_988);
xor U2479 (N_2479,In_2251,In_2352);
nand U2480 (N_2480,In_158,In_836);
or U2481 (N_2481,In_1299,In_1430);
xor U2482 (N_2482,In_602,In_2014);
nor U2483 (N_2483,In_1405,In_2140);
and U2484 (N_2484,In_950,In_187);
nand U2485 (N_2485,In_1074,In_1786);
and U2486 (N_2486,In_2442,In_131);
and U2487 (N_2487,In_2105,In_716);
nand U2488 (N_2488,In_1737,In_1907);
nor U2489 (N_2489,In_1755,In_1500);
nand U2490 (N_2490,In_485,In_1241);
and U2491 (N_2491,In_958,In_2033);
and U2492 (N_2492,In_1247,In_345);
xnor U2493 (N_2493,In_2211,In_2448);
nand U2494 (N_2494,In_2228,In_1402);
or U2495 (N_2495,In_2602,In_2539);
nor U2496 (N_2496,In_2271,In_1282);
or U2497 (N_2497,In_2555,In_1439);
nand U2498 (N_2498,In_1502,In_1403);
or U2499 (N_2499,In_2455,In_626);
nand U2500 (N_2500,In_462,In_264);
or U2501 (N_2501,In_2951,In_1432);
xnor U2502 (N_2502,In_2159,In_2324);
and U2503 (N_2503,In_707,In_2961);
or U2504 (N_2504,In_2374,In_1725);
nor U2505 (N_2505,In_286,In_341);
nand U2506 (N_2506,In_286,In_1536);
and U2507 (N_2507,In_982,In_2640);
or U2508 (N_2508,In_103,In_2321);
or U2509 (N_2509,In_2787,In_318);
and U2510 (N_2510,In_67,In_602);
or U2511 (N_2511,In_1419,In_2687);
and U2512 (N_2512,In_642,In_1355);
xor U2513 (N_2513,In_2586,In_531);
and U2514 (N_2514,In_1072,In_1075);
and U2515 (N_2515,In_1730,In_2938);
xnor U2516 (N_2516,In_1003,In_1313);
xnor U2517 (N_2517,In_197,In_532);
or U2518 (N_2518,In_1983,In_1996);
nor U2519 (N_2519,In_2251,In_1137);
or U2520 (N_2520,In_2691,In_30);
and U2521 (N_2521,In_2973,In_484);
xnor U2522 (N_2522,In_2468,In_942);
or U2523 (N_2523,In_2906,In_1972);
or U2524 (N_2524,In_1401,In_2240);
nor U2525 (N_2525,In_1667,In_83);
or U2526 (N_2526,In_2916,In_1804);
nor U2527 (N_2527,In_1636,In_948);
and U2528 (N_2528,In_2614,In_2790);
nor U2529 (N_2529,In_2062,In_871);
xnor U2530 (N_2530,In_1483,In_643);
nand U2531 (N_2531,In_2715,In_1443);
nand U2532 (N_2532,In_242,In_6);
nand U2533 (N_2533,In_1621,In_1000);
and U2534 (N_2534,In_933,In_1417);
nand U2535 (N_2535,In_1535,In_2151);
and U2536 (N_2536,In_1903,In_1485);
and U2537 (N_2537,In_1012,In_2672);
or U2538 (N_2538,In_760,In_861);
nand U2539 (N_2539,In_2554,In_2605);
nand U2540 (N_2540,In_1343,In_500);
nand U2541 (N_2541,In_1672,In_1417);
nor U2542 (N_2542,In_1153,In_2282);
nand U2543 (N_2543,In_2054,In_2162);
nand U2544 (N_2544,In_2731,In_1978);
or U2545 (N_2545,In_251,In_1281);
or U2546 (N_2546,In_438,In_528);
xnor U2547 (N_2547,In_1242,In_2262);
and U2548 (N_2548,In_373,In_2498);
xnor U2549 (N_2549,In_855,In_1566);
and U2550 (N_2550,In_987,In_1402);
and U2551 (N_2551,In_2484,In_2835);
nand U2552 (N_2552,In_393,In_135);
xor U2553 (N_2553,In_2338,In_1007);
and U2554 (N_2554,In_2701,In_1743);
and U2555 (N_2555,In_420,In_287);
nor U2556 (N_2556,In_2545,In_2749);
nand U2557 (N_2557,In_2918,In_1042);
or U2558 (N_2558,In_342,In_1977);
nand U2559 (N_2559,In_33,In_2199);
and U2560 (N_2560,In_518,In_2861);
nor U2561 (N_2561,In_1468,In_1628);
nor U2562 (N_2562,In_910,In_2988);
nor U2563 (N_2563,In_2710,In_2818);
nand U2564 (N_2564,In_138,In_226);
xnor U2565 (N_2565,In_1578,In_2220);
nand U2566 (N_2566,In_241,In_415);
or U2567 (N_2567,In_1009,In_502);
or U2568 (N_2568,In_1112,In_1067);
nor U2569 (N_2569,In_1919,In_95);
or U2570 (N_2570,In_2740,In_2668);
nor U2571 (N_2571,In_2010,In_2464);
or U2572 (N_2572,In_67,In_2399);
nand U2573 (N_2573,In_1147,In_1653);
nand U2574 (N_2574,In_903,In_636);
nor U2575 (N_2575,In_883,In_1241);
nand U2576 (N_2576,In_2105,In_2604);
nor U2577 (N_2577,In_2377,In_1061);
xnor U2578 (N_2578,In_1393,In_727);
nand U2579 (N_2579,In_2007,In_1040);
or U2580 (N_2580,In_2241,In_76);
and U2581 (N_2581,In_1899,In_1697);
or U2582 (N_2582,In_2356,In_1370);
and U2583 (N_2583,In_2985,In_2068);
nand U2584 (N_2584,In_1428,In_1705);
xor U2585 (N_2585,In_2191,In_1997);
or U2586 (N_2586,In_2046,In_1235);
or U2587 (N_2587,In_2714,In_305);
nor U2588 (N_2588,In_1592,In_1590);
nor U2589 (N_2589,In_2690,In_1400);
nor U2590 (N_2590,In_664,In_1215);
nand U2591 (N_2591,In_210,In_253);
and U2592 (N_2592,In_2612,In_254);
nand U2593 (N_2593,In_844,In_242);
or U2594 (N_2594,In_1083,In_931);
or U2595 (N_2595,In_1655,In_1341);
or U2596 (N_2596,In_1866,In_2057);
xnor U2597 (N_2597,In_2308,In_279);
and U2598 (N_2598,In_379,In_2539);
nor U2599 (N_2599,In_1916,In_855);
nand U2600 (N_2600,In_1650,In_2657);
nand U2601 (N_2601,In_644,In_401);
nand U2602 (N_2602,In_1337,In_2456);
nand U2603 (N_2603,In_486,In_2093);
nor U2604 (N_2604,In_1349,In_2895);
nor U2605 (N_2605,In_2384,In_2323);
nor U2606 (N_2606,In_1814,In_2429);
or U2607 (N_2607,In_191,In_56);
or U2608 (N_2608,In_1016,In_1919);
nand U2609 (N_2609,In_1748,In_90);
or U2610 (N_2610,In_2534,In_1476);
nor U2611 (N_2611,In_1365,In_2822);
nand U2612 (N_2612,In_1771,In_1637);
and U2613 (N_2613,In_1403,In_1699);
xnor U2614 (N_2614,In_189,In_2400);
nand U2615 (N_2615,In_263,In_589);
or U2616 (N_2616,In_702,In_345);
nor U2617 (N_2617,In_2499,In_2119);
nand U2618 (N_2618,In_785,In_671);
and U2619 (N_2619,In_2004,In_2826);
nand U2620 (N_2620,In_1935,In_1817);
nor U2621 (N_2621,In_973,In_2735);
nor U2622 (N_2622,In_2517,In_1729);
or U2623 (N_2623,In_2314,In_1300);
nor U2624 (N_2624,In_1983,In_1477);
nand U2625 (N_2625,In_1516,In_422);
xnor U2626 (N_2626,In_2173,In_2847);
nand U2627 (N_2627,In_1130,In_2728);
nand U2628 (N_2628,In_1316,In_2166);
and U2629 (N_2629,In_1055,In_2698);
and U2630 (N_2630,In_388,In_374);
or U2631 (N_2631,In_479,In_2393);
nor U2632 (N_2632,In_1565,In_128);
and U2633 (N_2633,In_2977,In_1243);
xnor U2634 (N_2634,In_587,In_500);
nor U2635 (N_2635,In_2545,In_1608);
nand U2636 (N_2636,In_2756,In_674);
and U2637 (N_2637,In_653,In_480);
nor U2638 (N_2638,In_487,In_1239);
nand U2639 (N_2639,In_496,In_933);
nand U2640 (N_2640,In_2852,In_1419);
xnor U2641 (N_2641,In_530,In_1579);
and U2642 (N_2642,In_2032,In_1684);
or U2643 (N_2643,In_21,In_1643);
nand U2644 (N_2644,In_1378,In_1570);
and U2645 (N_2645,In_316,In_2540);
nand U2646 (N_2646,In_1339,In_1572);
nand U2647 (N_2647,In_1194,In_1189);
or U2648 (N_2648,In_499,In_2078);
xnor U2649 (N_2649,In_333,In_2385);
and U2650 (N_2650,In_767,In_351);
and U2651 (N_2651,In_853,In_1765);
and U2652 (N_2652,In_2611,In_2807);
nor U2653 (N_2653,In_2249,In_1556);
and U2654 (N_2654,In_1361,In_992);
or U2655 (N_2655,In_1418,In_2103);
and U2656 (N_2656,In_2486,In_1809);
or U2657 (N_2657,In_2331,In_2437);
or U2658 (N_2658,In_2998,In_1730);
nand U2659 (N_2659,In_1519,In_2522);
nor U2660 (N_2660,In_1980,In_694);
and U2661 (N_2661,In_2423,In_1981);
nor U2662 (N_2662,In_629,In_2751);
or U2663 (N_2663,In_1151,In_1342);
nand U2664 (N_2664,In_1158,In_1800);
nor U2665 (N_2665,In_1554,In_1147);
or U2666 (N_2666,In_84,In_964);
nor U2667 (N_2667,In_1466,In_1828);
and U2668 (N_2668,In_2174,In_1893);
nand U2669 (N_2669,In_2281,In_2022);
xor U2670 (N_2670,In_2779,In_1295);
nor U2671 (N_2671,In_347,In_2636);
and U2672 (N_2672,In_2755,In_2464);
and U2673 (N_2673,In_1876,In_2684);
or U2674 (N_2674,In_2714,In_2366);
or U2675 (N_2675,In_1875,In_417);
xnor U2676 (N_2676,In_2103,In_2476);
nand U2677 (N_2677,In_2397,In_2250);
nor U2678 (N_2678,In_243,In_2330);
nor U2679 (N_2679,In_2920,In_343);
nor U2680 (N_2680,In_1173,In_1177);
xnor U2681 (N_2681,In_580,In_1053);
or U2682 (N_2682,In_338,In_1098);
and U2683 (N_2683,In_291,In_719);
nand U2684 (N_2684,In_1541,In_544);
or U2685 (N_2685,In_918,In_2357);
or U2686 (N_2686,In_1183,In_2140);
nor U2687 (N_2687,In_2736,In_296);
and U2688 (N_2688,In_337,In_530);
xor U2689 (N_2689,In_2315,In_891);
nor U2690 (N_2690,In_1017,In_1469);
and U2691 (N_2691,In_197,In_688);
and U2692 (N_2692,In_2543,In_848);
and U2693 (N_2693,In_307,In_1950);
or U2694 (N_2694,In_1528,In_1626);
nand U2695 (N_2695,In_488,In_734);
nor U2696 (N_2696,In_2792,In_211);
xnor U2697 (N_2697,In_325,In_1223);
or U2698 (N_2698,In_228,In_2280);
and U2699 (N_2699,In_260,In_489);
nor U2700 (N_2700,In_1793,In_538);
and U2701 (N_2701,In_2578,In_1180);
and U2702 (N_2702,In_2131,In_662);
nand U2703 (N_2703,In_2617,In_2141);
nand U2704 (N_2704,In_632,In_427);
and U2705 (N_2705,In_695,In_191);
xor U2706 (N_2706,In_2052,In_177);
and U2707 (N_2707,In_1959,In_855);
nor U2708 (N_2708,In_640,In_2500);
nor U2709 (N_2709,In_1137,In_1127);
xor U2710 (N_2710,In_2614,In_2683);
and U2711 (N_2711,In_1689,In_1024);
nor U2712 (N_2712,In_1658,In_547);
nand U2713 (N_2713,In_742,In_736);
or U2714 (N_2714,In_914,In_2081);
nor U2715 (N_2715,In_929,In_503);
nand U2716 (N_2716,In_2573,In_2735);
nand U2717 (N_2717,In_1845,In_159);
and U2718 (N_2718,In_1633,In_2899);
nor U2719 (N_2719,In_2032,In_2076);
or U2720 (N_2720,In_997,In_1710);
nand U2721 (N_2721,In_2891,In_1157);
and U2722 (N_2722,In_178,In_775);
or U2723 (N_2723,In_2925,In_857);
nor U2724 (N_2724,In_1161,In_2875);
nand U2725 (N_2725,In_2435,In_2304);
xnor U2726 (N_2726,In_97,In_1834);
nor U2727 (N_2727,In_1212,In_1299);
and U2728 (N_2728,In_914,In_252);
and U2729 (N_2729,In_2019,In_476);
xnor U2730 (N_2730,In_136,In_2330);
or U2731 (N_2731,In_620,In_2457);
or U2732 (N_2732,In_2782,In_1671);
or U2733 (N_2733,In_1617,In_483);
xnor U2734 (N_2734,In_910,In_1804);
nor U2735 (N_2735,In_1061,In_1650);
or U2736 (N_2736,In_1359,In_1618);
nand U2737 (N_2737,In_2673,In_2432);
nand U2738 (N_2738,In_29,In_723);
and U2739 (N_2739,In_134,In_1950);
nor U2740 (N_2740,In_653,In_1721);
and U2741 (N_2741,In_257,In_1178);
nor U2742 (N_2742,In_1325,In_904);
and U2743 (N_2743,In_2070,In_682);
nor U2744 (N_2744,In_726,In_1855);
and U2745 (N_2745,In_1521,In_2519);
nand U2746 (N_2746,In_2145,In_1039);
nand U2747 (N_2747,In_537,In_32);
xor U2748 (N_2748,In_186,In_2286);
nand U2749 (N_2749,In_1626,In_366);
and U2750 (N_2750,In_1146,In_2007);
nor U2751 (N_2751,In_2716,In_2879);
or U2752 (N_2752,In_1672,In_832);
nor U2753 (N_2753,In_2366,In_1273);
nand U2754 (N_2754,In_2300,In_104);
and U2755 (N_2755,In_1620,In_2584);
nand U2756 (N_2756,In_2121,In_2663);
and U2757 (N_2757,In_451,In_52);
or U2758 (N_2758,In_1271,In_1021);
or U2759 (N_2759,In_1997,In_611);
or U2760 (N_2760,In_87,In_2229);
xnor U2761 (N_2761,In_2068,In_911);
nand U2762 (N_2762,In_2738,In_2297);
nor U2763 (N_2763,In_1448,In_2985);
or U2764 (N_2764,In_532,In_2345);
nand U2765 (N_2765,In_1156,In_2550);
nand U2766 (N_2766,In_1479,In_281);
and U2767 (N_2767,In_2474,In_2573);
or U2768 (N_2768,In_703,In_1179);
or U2769 (N_2769,In_1442,In_348);
and U2770 (N_2770,In_556,In_760);
nand U2771 (N_2771,In_69,In_2310);
nor U2772 (N_2772,In_633,In_2680);
nand U2773 (N_2773,In_1366,In_1824);
nor U2774 (N_2774,In_1307,In_647);
xnor U2775 (N_2775,In_2936,In_2191);
or U2776 (N_2776,In_2207,In_1746);
nor U2777 (N_2777,In_2505,In_1221);
and U2778 (N_2778,In_2585,In_2051);
and U2779 (N_2779,In_2056,In_405);
nor U2780 (N_2780,In_709,In_2531);
nand U2781 (N_2781,In_1511,In_551);
xnor U2782 (N_2782,In_2254,In_2523);
nor U2783 (N_2783,In_2204,In_2171);
nand U2784 (N_2784,In_1650,In_1413);
or U2785 (N_2785,In_1726,In_1819);
and U2786 (N_2786,In_2621,In_2801);
and U2787 (N_2787,In_1236,In_2455);
nor U2788 (N_2788,In_1703,In_1986);
nand U2789 (N_2789,In_2974,In_1306);
nor U2790 (N_2790,In_2131,In_824);
and U2791 (N_2791,In_1448,In_2902);
nor U2792 (N_2792,In_2108,In_1246);
nand U2793 (N_2793,In_2367,In_1126);
xor U2794 (N_2794,In_2492,In_367);
nor U2795 (N_2795,In_2930,In_2923);
xnor U2796 (N_2796,In_2259,In_2145);
or U2797 (N_2797,In_2629,In_513);
and U2798 (N_2798,In_1622,In_2190);
nand U2799 (N_2799,In_2526,In_2850);
nor U2800 (N_2800,In_1825,In_407);
and U2801 (N_2801,In_1829,In_495);
and U2802 (N_2802,In_661,In_684);
or U2803 (N_2803,In_1401,In_734);
nand U2804 (N_2804,In_1829,In_822);
and U2805 (N_2805,In_1821,In_827);
nor U2806 (N_2806,In_1285,In_2362);
and U2807 (N_2807,In_1869,In_567);
xnor U2808 (N_2808,In_1253,In_1176);
or U2809 (N_2809,In_2394,In_601);
or U2810 (N_2810,In_1937,In_622);
nand U2811 (N_2811,In_774,In_2716);
xor U2812 (N_2812,In_2494,In_1269);
xnor U2813 (N_2813,In_1516,In_1439);
xor U2814 (N_2814,In_1368,In_1018);
nand U2815 (N_2815,In_253,In_950);
nand U2816 (N_2816,In_2970,In_1896);
nand U2817 (N_2817,In_292,In_1879);
or U2818 (N_2818,In_2888,In_206);
and U2819 (N_2819,In_383,In_1277);
nor U2820 (N_2820,In_652,In_1467);
nor U2821 (N_2821,In_2976,In_587);
or U2822 (N_2822,In_2449,In_2853);
and U2823 (N_2823,In_636,In_1278);
or U2824 (N_2824,In_1296,In_532);
nand U2825 (N_2825,In_1376,In_1316);
xnor U2826 (N_2826,In_2365,In_2676);
nand U2827 (N_2827,In_1471,In_2956);
nand U2828 (N_2828,In_125,In_1588);
nor U2829 (N_2829,In_1776,In_2435);
nor U2830 (N_2830,In_959,In_187);
and U2831 (N_2831,In_1937,In_1355);
and U2832 (N_2832,In_314,In_2180);
and U2833 (N_2833,In_780,In_1220);
and U2834 (N_2834,In_575,In_1566);
or U2835 (N_2835,In_1360,In_27);
nand U2836 (N_2836,In_1023,In_1991);
or U2837 (N_2837,In_519,In_2306);
nand U2838 (N_2838,In_2597,In_2224);
nor U2839 (N_2839,In_2164,In_1039);
nand U2840 (N_2840,In_2399,In_2943);
or U2841 (N_2841,In_1832,In_419);
nand U2842 (N_2842,In_1378,In_2880);
xor U2843 (N_2843,In_897,In_1721);
or U2844 (N_2844,In_1260,In_2949);
xnor U2845 (N_2845,In_398,In_2291);
xnor U2846 (N_2846,In_437,In_151);
nand U2847 (N_2847,In_2853,In_2880);
and U2848 (N_2848,In_2512,In_688);
nand U2849 (N_2849,In_2788,In_1278);
or U2850 (N_2850,In_30,In_2477);
and U2851 (N_2851,In_249,In_2591);
and U2852 (N_2852,In_1485,In_1405);
or U2853 (N_2853,In_975,In_670);
xor U2854 (N_2854,In_2,In_945);
and U2855 (N_2855,In_748,In_966);
or U2856 (N_2856,In_954,In_544);
nor U2857 (N_2857,In_1807,In_1091);
nor U2858 (N_2858,In_1756,In_1494);
nor U2859 (N_2859,In_2933,In_1265);
and U2860 (N_2860,In_419,In_1709);
or U2861 (N_2861,In_2032,In_2146);
or U2862 (N_2862,In_1978,In_2905);
nor U2863 (N_2863,In_82,In_2279);
nor U2864 (N_2864,In_1569,In_439);
xor U2865 (N_2865,In_2067,In_2415);
nor U2866 (N_2866,In_339,In_1410);
xnor U2867 (N_2867,In_1113,In_1281);
nor U2868 (N_2868,In_1073,In_2537);
xnor U2869 (N_2869,In_1098,In_842);
and U2870 (N_2870,In_2218,In_1174);
or U2871 (N_2871,In_930,In_733);
or U2872 (N_2872,In_2874,In_2069);
xor U2873 (N_2873,In_781,In_2450);
or U2874 (N_2874,In_726,In_2636);
and U2875 (N_2875,In_1516,In_1482);
or U2876 (N_2876,In_1522,In_1062);
or U2877 (N_2877,In_865,In_2583);
xor U2878 (N_2878,In_563,In_1194);
nor U2879 (N_2879,In_73,In_311);
and U2880 (N_2880,In_1621,In_1956);
nand U2881 (N_2881,In_2388,In_51);
or U2882 (N_2882,In_2414,In_378);
nor U2883 (N_2883,In_129,In_1202);
xnor U2884 (N_2884,In_1000,In_2454);
nor U2885 (N_2885,In_781,In_996);
and U2886 (N_2886,In_2066,In_1829);
and U2887 (N_2887,In_2961,In_627);
or U2888 (N_2888,In_2446,In_268);
xor U2889 (N_2889,In_1674,In_1354);
and U2890 (N_2890,In_537,In_1550);
xnor U2891 (N_2891,In_274,In_2290);
nand U2892 (N_2892,In_385,In_865);
nor U2893 (N_2893,In_261,In_213);
nor U2894 (N_2894,In_57,In_2985);
xor U2895 (N_2895,In_2224,In_395);
nand U2896 (N_2896,In_920,In_2849);
and U2897 (N_2897,In_1985,In_11);
nand U2898 (N_2898,In_2056,In_1255);
or U2899 (N_2899,In_597,In_1184);
nand U2900 (N_2900,In_1339,In_1217);
nor U2901 (N_2901,In_1652,In_1390);
nand U2902 (N_2902,In_274,In_2928);
nor U2903 (N_2903,In_2839,In_1463);
and U2904 (N_2904,In_1763,In_1051);
nor U2905 (N_2905,In_1245,In_366);
nand U2906 (N_2906,In_2722,In_161);
or U2907 (N_2907,In_2091,In_258);
nand U2908 (N_2908,In_741,In_1358);
nand U2909 (N_2909,In_2235,In_1126);
nand U2910 (N_2910,In_2312,In_1145);
and U2911 (N_2911,In_202,In_2769);
nor U2912 (N_2912,In_2810,In_2704);
or U2913 (N_2913,In_2536,In_1840);
nor U2914 (N_2914,In_1552,In_1192);
nand U2915 (N_2915,In_116,In_497);
nor U2916 (N_2916,In_2799,In_33);
nand U2917 (N_2917,In_1359,In_512);
xnor U2918 (N_2918,In_1532,In_2656);
nor U2919 (N_2919,In_1990,In_2548);
nor U2920 (N_2920,In_1173,In_2313);
nand U2921 (N_2921,In_2876,In_550);
and U2922 (N_2922,In_2665,In_264);
or U2923 (N_2923,In_2658,In_546);
or U2924 (N_2924,In_350,In_226);
and U2925 (N_2925,In_233,In_1684);
or U2926 (N_2926,In_1122,In_140);
and U2927 (N_2927,In_2979,In_363);
and U2928 (N_2928,In_317,In_673);
nand U2929 (N_2929,In_2456,In_48);
nand U2930 (N_2930,In_1046,In_1944);
nand U2931 (N_2931,In_399,In_2253);
xor U2932 (N_2932,In_2698,In_1034);
xor U2933 (N_2933,In_1423,In_1611);
or U2934 (N_2934,In_330,In_2593);
nor U2935 (N_2935,In_2017,In_202);
nand U2936 (N_2936,In_1460,In_39);
nand U2937 (N_2937,In_1825,In_2628);
or U2938 (N_2938,In_1959,In_940);
nand U2939 (N_2939,In_1258,In_733);
and U2940 (N_2940,In_1133,In_127);
xor U2941 (N_2941,In_60,In_1392);
and U2942 (N_2942,In_336,In_192);
and U2943 (N_2943,In_275,In_1082);
or U2944 (N_2944,In_1537,In_2708);
xor U2945 (N_2945,In_455,In_2749);
xnor U2946 (N_2946,In_1944,In_1146);
and U2947 (N_2947,In_2893,In_2117);
xor U2948 (N_2948,In_2098,In_2515);
or U2949 (N_2949,In_2913,In_2947);
nor U2950 (N_2950,In_2069,In_2825);
and U2951 (N_2951,In_119,In_600);
nand U2952 (N_2952,In_886,In_2648);
nor U2953 (N_2953,In_1840,In_2484);
xnor U2954 (N_2954,In_575,In_2093);
nand U2955 (N_2955,In_130,In_1028);
or U2956 (N_2956,In_2549,In_900);
xnor U2957 (N_2957,In_1130,In_252);
nand U2958 (N_2958,In_1951,In_2881);
nand U2959 (N_2959,In_2208,In_2939);
and U2960 (N_2960,In_336,In_2771);
nor U2961 (N_2961,In_1356,In_2248);
or U2962 (N_2962,In_2869,In_1382);
nor U2963 (N_2963,In_1199,In_55);
nand U2964 (N_2964,In_911,In_433);
or U2965 (N_2965,In_2780,In_749);
nor U2966 (N_2966,In_1615,In_1344);
nand U2967 (N_2967,In_2834,In_2607);
and U2968 (N_2968,In_903,In_995);
nor U2969 (N_2969,In_2458,In_967);
nor U2970 (N_2970,In_1754,In_2595);
and U2971 (N_2971,In_418,In_2199);
or U2972 (N_2972,In_1017,In_2452);
nand U2973 (N_2973,In_1169,In_19);
and U2974 (N_2974,In_2359,In_1556);
or U2975 (N_2975,In_790,In_1004);
or U2976 (N_2976,In_1605,In_2319);
or U2977 (N_2977,In_464,In_1283);
and U2978 (N_2978,In_1426,In_215);
and U2979 (N_2979,In_1447,In_1032);
nor U2980 (N_2980,In_2400,In_1125);
nor U2981 (N_2981,In_626,In_2548);
nor U2982 (N_2982,In_1059,In_622);
or U2983 (N_2983,In_2901,In_2638);
and U2984 (N_2984,In_1608,In_836);
nand U2985 (N_2985,In_495,In_729);
xnor U2986 (N_2986,In_1092,In_1754);
nor U2987 (N_2987,In_1489,In_36);
or U2988 (N_2988,In_1502,In_2737);
nand U2989 (N_2989,In_1829,In_2179);
nor U2990 (N_2990,In_1158,In_822);
and U2991 (N_2991,In_85,In_2996);
nand U2992 (N_2992,In_2471,In_367);
xnor U2993 (N_2993,In_2585,In_2384);
or U2994 (N_2994,In_1525,In_2307);
and U2995 (N_2995,In_2871,In_2505);
and U2996 (N_2996,In_747,In_2558);
and U2997 (N_2997,In_2119,In_359);
and U2998 (N_2998,In_2963,In_2971);
xnor U2999 (N_2999,In_2964,In_2776);
nand U3000 (N_3000,In_2440,In_142);
or U3001 (N_3001,In_1966,In_1001);
and U3002 (N_3002,In_1187,In_52);
and U3003 (N_3003,In_1724,In_2079);
nand U3004 (N_3004,In_885,In_1819);
xnor U3005 (N_3005,In_1390,In_1862);
xor U3006 (N_3006,In_2309,In_261);
nor U3007 (N_3007,In_1618,In_1474);
and U3008 (N_3008,In_1679,In_2035);
nand U3009 (N_3009,In_2862,In_1713);
and U3010 (N_3010,In_2156,In_266);
xnor U3011 (N_3011,In_2333,In_2671);
nand U3012 (N_3012,In_1107,In_1225);
nor U3013 (N_3013,In_1392,In_449);
nand U3014 (N_3014,In_2301,In_1146);
xor U3015 (N_3015,In_954,In_365);
or U3016 (N_3016,In_2487,In_2139);
and U3017 (N_3017,In_1676,In_2666);
and U3018 (N_3018,In_2130,In_851);
or U3019 (N_3019,In_567,In_2327);
nand U3020 (N_3020,In_865,In_472);
or U3021 (N_3021,In_1496,In_367);
nand U3022 (N_3022,In_816,In_2018);
and U3023 (N_3023,In_621,In_862);
and U3024 (N_3024,In_2114,In_1034);
nor U3025 (N_3025,In_2915,In_1221);
and U3026 (N_3026,In_2346,In_421);
nor U3027 (N_3027,In_2101,In_1311);
nand U3028 (N_3028,In_622,In_1556);
or U3029 (N_3029,In_1257,In_874);
nor U3030 (N_3030,In_535,In_1369);
or U3031 (N_3031,In_1771,In_765);
and U3032 (N_3032,In_1373,In_2909);
xor U3033 (N_3033,In_726,In_389);
and U3034 (N_3034,In_1625,In_184);
xnor U3035 (N_3035,In_609,In_53);
or U3036 (N_3036,In_2778,In_895);
and U3037 (N_3037,In_1530,In_1112);
or U3038 (N_3038,In_1505,In_2305);
xnor U3039 (N_3039,In_1993,In_128);
nand U3040 (N_3040,In_2589,In_206);
or U3041 (N_3041,In_2193,In_1799);
xor U3042 (N_3042,In_2212,In_2443);
xor U3043 (N_3043,In_353,In_2461);
and U3044 (N_3044,In_142,In_2824);
or U3045 (N_3045,In_2021,In_2396);
nor U3046 (N_3046,In_201,In_925);
xnor U3047 (N_3047,In_53,In_1776);
nor U3048 (N_3048,In_814,In_1651);
or U3049 (N_3049,In_1733,In_2210);
or U3050 (N_3050,In_2685,In_356);
nor U3051 (N_3051,In_2069,In_1475);
or U3052 (N_3052,In_2446,In_1157);
nand U3053 (N_3053,In_2829,In_959);
nor U3054 (N_3054,In_2749,In_2733);
and U3055 (N_3055,In_745,In_1773);
nor U3056 (N_3056,In_2297,In_2165);
xor U3057 (N_3057,In_1038,In_2888);
and U3058 (N_3058,In_1786,In_2117);
nor U3059 (N_3059,In_2816,In_845);
and U3060 (N_3060,In_198,In_1654);
xnor U3061 (N_3061,In_2425,In_2595);
nand U3062 (N_3062,In_1412,In_1341);
nand U3063 (N_3063,In_1698,In_236);
xor U3064 (N_3064,In_2423,In_1182);
nor U3065 (N_3065,In_1775,In_1946);
nand U3066 (N_3066,In_671,In_1924);
nor U3067 (N_3067,In_2187,In_1467);
nor U3068 (N_3068,In_1012,In_2045);
nor U3069 (N_3069,In_1730,In_2452);
and U3070 (N_3070,In_1535,In_2558);
nor U3071 (N_3071,In_2088,In_1090);
nor U3072 (N_3072,In_319,In_1995);
nor U3073 (N_3073,In_1597,In_2894);
or U3074 (N_3074,In_1931,In_2578);
nor U3075 (N_3075,In_2375,In_1998);
and U3076 (N_3076,In_2433,In_652);
nand U3077 (N_3077,In_2238,In_1428);
and U3078 (N_3078,In_161,In_1650);
nor U3079 (N_3079,In_1846,In_2811);
and U3080 (N_3080,In_359,In_2353);
nor U3081 (N_3081,In_1928,In_1243);
nand U3082 (N_3082,In_721,In_2137);
nor U3083 (N_3083,In_44,In_1787);
nor U3084 (N_3084,In_422,In_1520);
or U3085 (N_3085,In_1432,In_1365);
and U3086 (N_3086,In_1906,In_2606);
and U3087 (N_3087,In_2804,In_2556);
nor U3088 (N_3088,In_446,In_1264);
or U3089 (N_3089,In_2784,In_2713);
nor U3090 (N_3090,In_1462,In_381);
nand U3091 (N_3091,In_1059,In_2976);
or U3092 (N_3092,In_28,In_1083);
or U3093 (N_3093,In_1812,In_2517);
nor U3094 (N_3094,In_2775,In_1093);
nand U3095 (N_3095,In_2921,In_2117);
nor U3096 (N_3096,In_2047,In_1312);
or U3097 (N_3097,In_1866,In_2653);
and U3098 (N_3098,In_2115,In_2458);
and U3099 (N_3099,In_2775,In_555);
nor U3100 (N_3100,In_1819,In_2800);
xnor U3101 (N_3101,In_1554,In_188);
nor U3102 (N_3102,In_1717,In_469);
and U3103 (N_3103,In_1793,In_1783);
nor U3104 (N_3104,In_1774,In_415);
nor U3105 (N_3105,In_264,In_134);
nor U3106 (N_3106,In_872,In_1287);
nand U3107 (N_3107,In_1791,In_798);
or U3108 (N_3108,In_1677,In_1704);
nor U3109 (N_3109,In_592,In_786);
xor U3110 (N_3110,In_1414,In_2400);
xor U3111 (N_3111,In_237,In_2110);
xnor U3112 (N_3112,In_2267,In_116);
or U3113 (N_3113,In_2622,In_2060);
or U3114 (N_3114,In_1447,In_992);
and U3115 (N_3115,In_1103,In_2837);
and U3116 (N_3116,In_20,In_1284);
or U3117 (N_3117,In_2483,In_1551);
xor U3118 (N_3118,In_417,In_2635);
and U3119 (N_3119,In_2048,In_1186);
nand U3120 (N_3120,In_725,In_2609);
nor U3121 (N_3121,In_2461,In_2670);
nor U3122 (N_3122,In_1451,In_1683);
nand U3123 (N_3123,In_2312,In_1973);
or U3124 (N_3124,In_1618,In_1154);
xnor U3125 (N_3125,In_954,In_2964);
or U3126 (N_3126,In_1707,In_313);
or U3127 (N_3127,In_2575,In_2108);
and U3128 (N_3128,In_1878,In_2619);
nor U3129 (N_3129,In_916,In_1393);
and U3130 (N_3130,In_2293,In_2952);
nor U3131 (N_3131,In_1753,In_1547);
nor U3132 (N_3132,In_285,In_2578);
and U3133 (N_3133,In_825,In_2627);
nand U3134 (N_3134,In_2396,In_1607);
and U3135 (N_3135,In_1496,In_2112);
or U3136 (N_3136,In_2190,In_1754);
nor U3137 (N_3137,In_2172,In_146);
nor U3138 (N_3138,In_2588,In_1336);
or U3139 (N_3139,In_1632,In_308);
nand U3140 (N_3140,In_200,In_2159);
or U3141 (N_3141,In_719,In_153);
and U3142 (N_3142,In_2366,In_229);
or U3143 (N_3143,In_200,In_2116);
nand U3144 (N_3144,In_2272,In_2318);
or U3145 (N_3145,In_440,In_1238);
nor U3146 (N_3146,In_2623,In_897);
nor U3147 (N_3147,In_745,In_91);
or U3148 (N_3148,In_243,In_1387);
or U3149 (N_3149,In_2966,In_1286);
and U3150 (N_3150,In_2284,In_884);
nor U3151 (N_3151,In_1434,In_316);
nand U3152 (N_3152,In_1850,In_2341);
nor U3153 (N_3153,In_2581,In_2206);
nor U3154 (N_3154,In_1199,In_830);
nor U3155 (N_3155,In_395,In_1823);
nor U3156 (N_3156,In_2139,In_2900);
nor U3157 (N_3157,In_1457,In_1716);
or U3158 (N_3158,In_2334,In_2080);
or U3159 (N_3159,In_1677,In_2693);
and U3160 (N_3160,In_2612,In_419);
nor U3161 (N_3161,In_2598,In_2979);
or U3162 (N_3162,In_82,In_582);
and U3163 (N_3163,In_2895,In_1397);
or U3164 (N_3164,In_2598,In_2421);
or U3165 (N_3165,In_1406,In_676);
nor U3166 (N_3166,In_100,In_1388);
nor U3167 (N_3167,In_2729,In_132);
nor U3168 (N_3168,In_97,In_1751);
and U3169 (N_3169,In_1961,In_1622);
and U3170 (N_3170,In_1534,In_2231);
xor U3171 (N_3171,In_2986,In_1328);
nor U3172 (N_3172,In_603,In_423);
nor U3173 (N_3173,In_2173,In_1603);
nand U3174 (N_3174,In_1972,In_2293);
and U3175 (N_3175,In_975,In_2588);
or U3176 (N_3176,In_1801,In_2697);
nand U3177 (N_3177,In_1879,In_303);
nand U3178 (N_3178,In_1366,In_1901);
or U3179 (N_3179,In_2900,In_822);
nand U3180 (N_3180,In_656,In_2163);
nor U3181 (N_3181,In_821,In_2102);
or U3182 (N_3182,In_1334,In_2842);
nor U3183 (N_3183,In_2800,In_2147);
and U3184 (N_3184,In_204,In_524);
nand U3185 (N_3185,In_2800,In_1089);
nor U3186 (N_3186,In_1769,In_1253);
nor U3187 (N_3187,In_647,In_893);
nor U3188 (N_3188,In_799,In_900);
xor U3189 (N_3189,In_2316,In_2817);
xor U3190 (N_3190,In_263,In_2065);
or U3191 (N_3191,In_2676,In_1951);
and U3192 (N_3192,In_2207,In_2226);
nor U3193 (N_3193,In_1451,In_308);
nand U3194 (N_3194,In_2951,In_2517);
and U3195 (N_3195,In_2250,In_1186);
or U3196 (N_3196,In_2067,In_804);
nor U3197 (N_3197,In_2391,In_1141);
nor U3198 (N_3198,In_873,In_1171);
and U3199 (N_3199,In_2486,In_901);
and U3200 (N_3200,In_1361,In_2327);
and U3201 (N_3201,In_1274,In_2661);
nand U3202 (N_3202,In_2863,In_1755);
nand U3203 (N_3203,In_255,In_1529);
or U3204 (N_3204,In_1795,In_990);
and U3205 (N_3205,In_2374,In_2291);
nand U3206 (N_3206,In_1752,In_1349);
nand U3207 (N_3207,In_2540,In_2076);
nand U3208 (N_3208,In_575,In_488);
nand U3209 (N_3209,In_584,In_888);
and U3210 (N_3210,In_902,In_1642);
or U3211 (N_3211,In_2101,In_711);
or U3212 (N_3212,In_2051,In_529);
or U3213 (N_3213,In_2782,In_218);
or U3214 (N_3214,In_365,In_2350);
and U3215 (N_3215,In_2042,In_873);
nor U3216 (N_3216,In_262,In_270);
or U3217 (N_3217,In_450,In_1044);
nand U3218 (N_3218,In_877,In_504);
and U3219 (N_3219,In_1201,In_975);
and U3220 (N_3220,In_467,In_911);
or U3221 (N_3221,In_2341,In_1848);
nand U3222 (N_3222,In_1979,In_1404);
and U3223 (N_3223,In_193,In_1605);
or U3224 (N_3224,In_664,In_887);
nand U3225 (N_3225,In_927,In_2615);
or U3226 (N_3226,In_1779,In_2963);
xor U3227 (N_3227,In_1061,In_2171);
and U3228 (N_3228,In_2601,In_623);
and U3229 (N_3229,In_494,In_1491);
xor U3230 (N_3230,In_925,In_701);
nand U3231 (N_3231,In_1819,In_555);
or U3232 (N_3232,In_2249,In_2112);
nand U3233 (N_3233,In_2241,In_823);
xor U3234 (N_3234,In_240,In_1867);
nor U3235 (N_3235,In_1987,In_969);
and U3236 (N_3236,In_337,In_737);
xnor U3237 (N_3237,In_2053,In_2678);
nor U3238 (N_3238,In_1858,In_2096);
and U3239 (N_3239,In_732,In_1805);
nor U3240 (N_3240,In_366,In_1154);
xnor U3241 (N_3241,In_2387,In_1186);
nand U3242 (N_3242,In_1154,In_460);
or U3243 (N_3243,In_2888,In_1931);
or U3244 (N_3244,In_2746,In_2842);
nor U3245 (N_3245,In_1686,In_602);
nand U3246 (N_3246,In_2114,In_949);
and U3247 (N_3247,In_2769,In_2998);
nor U3248 (N_3248,In_2927,In_1948);
or U3249 (N_3249,In_805,In_317);
nor U3250 (N_3250,In_1943,In_2132);
nand U3251 (N_3251,In_2406,In_2663);
nor U3252 (N_3252,In_1745,In_852);
nand U3253 (N_3253,In_1969,In_2612);
nor U3254 (N_3254,In_318,In_72);
or U3255 (N_3255,In_486,In_31);
nor U3256 (N_3256,In_543,In_533);
or U3257 (N_3257,In_2888,In_2912);
nand U3258 (N_3258,In_1817,In_2620);
and U3259 (N_3259,In_2508,In_639);
and U3260 (N_3260,In_834,In_513);
nor U3261 (N_3261,In_2979,In_2332);
nand U3262 (N_3262,In_1474,In_2154);
nor U3263 (N_3263,In_405,In_2402);
and U3264 (N_3264,In_524,In_14);
nor U3265 (N_3265,In_2156,In_1305);
xor U3266 (N_3266,In_2697,In_2684);
xnor U3267 (N_3267,In_2425,In_413);
and U3268 (N_3268,In_32,In_1357);
nor U3269 (N_3269,In_1941,In_2346);
nand U3270 (N_3270,In_910,In_1152);
or U3271 (N_3271,In_1947,In_815);
xor U3272 (N_3272,In_201,In_646);
and U3273 (N_3273,In_795,In_1120);
nand U3274 (N_3274,In_2604,In_2627);
nor U3275 (N_3275,In_1754,In_514);
and U3276 (N_3276,In_2592,In_102);
nor U3277 (N_3277,In_547,In_1329);
or U3278 (N_3278,In_2628,In_903);
and U3279 (N_3279,In_2619,In_832);
nor U3280 (N_3280,In_941,In_1756);
nor U3281 (N_3281,In_1747,In_2657);
nor U3282 (N_3282,In_2400,In_1724);
or U3283 (N_3283,In_1980,In_2843);
nand U3284 (N_3284,In_629,In_53);
and U3285 (N_3285,In_660,In_202);
and U3286 (N_3286,In_2619,In_1428);
nor U3287 (N_3287,In_1403,In_2462);
and U3288 (N_3288,In_1841,In_1337);
or U3289 (N_3289,In_2356,In_2779);
nor U3290 (N_3290,In_1000,In_848);
or U3291 (N_3291,In_1089,In_1694);
or U3292 (N_3292,In_1080,In_2336);
or U3293 (N_3293,In_1921,In_328);
or U3294 (N_3294,In_1743,In_2426);
and U3295 (N_3295,In_1050,In_2633);
or U3296 (N_3296,In_1335,In_1999);
or U3297 (N_3297,In_1659,In_2382);
and U3298 (N_3298,In_1205,In_923);
nor U3299 (N_3299,In_2572,In_178);
and U3300 (N_3300,In_1328,In_1454);
nand U3301 (N_3301,In_1714,In_2307);
or U3302 (N_3302,In_693,In_1568);
or U3303 (N_3303,In_831,In_2129);
or U3304 (N_3304,In_1456,In_1811);
or U3305 (N_3305,In_2710,In_371);
nand U3306 (N_3306,In_484,In_1068);
nand U3307 (N_3307,In_1580,In_739);
nand U3308 (N_3308,In_1135,In_2242);
nand U3309 (N_3309,In_1736,In_2357);
or U3310 (N_3310,In_2823,In_327);
and U3311 (N_3311,In_1834,In_741);
and U3312 (N_3312,In_1947,In_2006);
and U3313 (N_3313,In_1026,In_255);
nand U3314 (N_3314,In_230,In_2205);
nand U3315 (N_3315,In_1881,In_1342);
nor U3316 (N_3316,In_1547,In_87);
or U3317 (N_3317,In_2018,In_1001);
and U3318 (N_3318,In_2859,In_1478);
xnor U3319 (N_3319,In_1837,In_0);
nor U3320 (N_3320,In_1883,In_70);
and U3321 (N_3321,In_324,In_2060);
and U3322 (N_3322,In_1763,In_2094);
nand U3323 (N_3323,In_31,In_1215);
and U3324 (N_3324,In_2202,In_1867);
or U3325 (N_3325,In_1214,In_1812);
nand U3326 (N_3326,In_1926,In_2765);
nor U3327 (N_3327,In_343,In_1372);
and U3328 (N_3328,In_2561,In_2446);
or U3329 (N_3329,In_2125,In_2772);
nor U3330 (N_3330,In_525,In_2599);
and U3331 (N_3331,In_2426,In_2518);
nand U3332 (N_3332,In_1264,In_1689);
nand U3333 (N_3333,In_2892,In_1038);
nand U3334 (N_3334,In_2598,In_1553);
or U3335 (N_3335,In_1508,In_79);
or U3336 (N_3336,In_1575,In_2412);
nor U3337 (N_3337,In_866,In_70);
or U3338 (N_3338,In_2535,In_1082);
nand U3339 (N_3339,In_885,In_1902);
nand U3340 (N_3340,In_2534,In_2609);
or U3341 (N_3341,In_1429,In_1541);
nor U3342 (N_3342,In_544,In_1616);
xnor U3343 (N_3343,In_2433,In_1390);
and U3344 (N_3344,In_1459,In_1500);
and U3345 (N_3345,In_205,In_2465);
and U3346 (N_3346,In_1618,In_686);
or U3347 (N_3347,In_1953,In_735);
nor U3348 (N_3348,In_2447,In_2017);
nand U3349 (N_3349,In_2382,In_18);
nand U3350 (N_3350,In_2107,In_2775);
or U3351 (N_3351,In_977,In_1547);
nand U3352 (N_3352,In_2176,In_1479);
nor U3353 (N_3353,In_1571,In_2675);
nand U3354 (N_3354,In_858,In_2635);
nand U3355 (N_3355,In_1060,In_331);
nor U3356 (N_3356,In_2445,In_695);
nor U3357 (N_3357,In_2967,In_362);
and U3358 (N_3358,In_2932,In_809);
or U3359 (N_3359,In_1041,In_2860);
nand U3360 (N_3360,In_2385,In_136);
nor U3361 (N_3361,In_1523,In_2324);
or U3362 (N_3362,In_233,In_2797);
nor U3363 (N_3363,In_1666,In_642);
and U3364 (N_3364,In_922,In_997);
xnor U3365 (N_3365,In_151,In_677);
nand U3366 (N_3366,In_825,In_843);
or U3367 (N_3367,In_36,In_1046);
nand U3368 (N_3368,In_770,In_1338);
or U3369 (N_3369,In_1135,In_2208);
nand U3370 (N_3370,In_139,In_38);
nor U3371 (N_3371,In_902,In_2911);
nand U3372 (N_3372,In_868,In_2824);
nand U3373 (N_3373,In_2502,In_911);
and U3374 (N_3374,In_1840,In_1054);
or U3375 (N_3375,In_2066,In_1882);
nor U3376 (N_3376,In_228,In_121);
nor U3377 (N_3377,In_2897,In_317);
and U3378 (N_3378,In_2157,In_1923);
and U3379 (N_3379,In_2449,In_549);
and U3380 (N_3380,In_1861,In_2523);
nand U3381 (N_3381,In_997,In_431);
nand U3382 (N_3382,In_90,In_935);
or U3383 (N_3383,In_474,In_1367);
and U3384 (N_3384,In_1238,In_2409);
nor U3385 (N_3385,In_2910,In_553);
nor U3386 (N_3386,In_448,In_365);
nand U3387 (N_3387,In_230,In_2187);
nor U3388 (N_3388,In_2414,In_1092);
nor U3389 (N_3389,In_2484,In_2313);
or U3390 (N_3390,In_1061,In_2598);
and U3391 (N_3391,In_1368,In_1752);
nand U3392 (N_3392,In_667,In_2325);
xor U3393 (N_3393,In_513,In_1867);
xnor U3394 (N_3394,In_2457,In_2736);
or U3395 (N_3395,In_2641,In_1091);
nor U3396 (N_3396,In_1680,In_586);
nand U3397 (N_3397,In_510,In_1092);
and U3398 (N_3398,In_341,In_1217);
or U3399 (N_3399,In_2158,In_2949);
nand U3400 (N_3400,In_541,In_1350);
or U3401 (N_3401,In_2924,In_1003);
and U3402 (N_3402,In_1423,In_2736);
nor U3403 (N_3403,In_1300,In_1003);
and U3404 (N_3404,In_1016,In_117);
or U3405 (N_3405,In_269,In_1259);
or U3406 (N_3406,In_2824,In_2573);
nand U3407 (N_3407,In_1396,In_1156);
and U3408 (N_3408,In_2755,In_1270);
and U3409 (N_3409,In_826,In_2539);
nand U3410 (N_3410,In_1103,In_1657);
and U3411 (N_3411,In_478,In_1788);
nor U3412 (N_3412,In_1074,In_910);
nor U3413 (N_3413,In_2778,In_2833);
nand U3414 (N_3414,In_280,In_324);
or U3415 (N_3415,In_637,In_1876);
nand U3416 (N_3416,In_394,In_256);
and U3417 (N_3417,In_2027,In_1011);
nand U3418 (N_3418,In_2997,In_1578);
nor U3419 (N_3419,In_2350,In_2253);
or U3420 (N_3420,In_2791,In_1225);
nand U3421 (N_3421,In_2820,In_640);
nand U3422 (N_3422,In_2331,In_2763);
nand U3423 (N_3423,In_1018,In_365);
or U3424 (N_3424,In_715,In_2929);
or U3425 (N_3425,In_2294,In_63);
nand U3426 (N_3426,In_2607,In_1713);
xor U3427 (N_3427,In_2738,In_201);
or U3428 (N_3428,In_773,In_924);
nand U3429 (N_3429,In_387,In_2022);
nand U3430 (N_3430,In_2995,In_685);
xnor U3431 (N_3431,In_4,In_817);
or U3432 (N_3432,In_1198,In_440);
nand U3433 (N_3433,In_2646,In_1388);
and U3434 (N_3434,In_295,In_1993);
and U3435 (N_3435,In_2712,In_2077);
nor U3436 (N_3436,In_1085,In_109);
nor U3437 (N_3437,In_2521,In_2230);
and U3438 (N_3438,In_776,In_211);
nand U3439 (N_3439,In_13,In_1602);
nand U3440 (N_3440,In_285,In_2300);
and U3441 (N_3441,In_2751,In_792);
nor U3442 (N_3442,In_2866,In_2904);
xor U3443 (N_3443,In_185,In_2420);
and U3444 (N_3444,In_2971,In_2043);
nor U3445 (N_3445,In_2406,In_1863);
nand U3446 (N_3446,In_71,In_1876);
or U3447 (N_3447,In_2109,In_1941);
nor U3448 (N_3448,In_20,In_1560);
or U3449 (N_3449,In_1343,In_568);
and U3450 (N_3450,In_2894,In_2046);
or U3451 (N_3451,In_547,In_236);
nand U3452 (N_3452,In_2078,In_914);
and U3453 (N_3453,In_76,In_869);
xor U3454 (N_3454,In_2993,In_2466);
nor U3455 (N_3455,In_1123,In_1731);
nor U3456 (N_3456,In_2093,In_1255);
or U3457 (N_3457,In_2118,In_355);
nand U3458 (N_3458,In_1095,In_2643);
nor U3459 (N_3459,In_2673,In_792);
nand U3460 (N_3460,In_2799,In_2131);
or U3461 (N_3461,In_2731,In_2494);
nor U3462 (N_3462,In_2011,In_1799);
nor U3463 (N_3463,In_1096,In_1397);
nand U3464 (N_3464,In_513,In_1222);
xor U3465 (N_3465,In_232,In_2696);
or U3466 (N_3466,In_345,In_0);
nand U3467 (N_3467,In_374,In_609);
and U3468 (N_3468,In_1077,In_2465);
nor U3469 (N_3469,In_1836,In_2351);
xor U3470 (N_3470,In_1689,In_2944);
or U3471 (N_3471,In_2323,In_934);
and U3472 (N_3472,In_1910,In_1323);
nand U3473 (N_3473,In_214,In_695);
nand U3474 (N_3474,In_2670,In_1395);
nor U3475 (N_3475,In_913,In_1733);
and U3476 (N_3476,In_1851,In_1203);
nor U3477 (N_3477,In_1007,In_1067);
nor U3478 (N_3478,In_2159,In_2034);
nor U3479 (N_3479,In_2231,In_736);
or U3480 (N_3480,In_2459,In_2046);
and U3481 (N_3481,In_27,In_272);
nor U3482 (N_3482,In_754,In_2370);
nor U3483 (N_3483,In_1653,In_2949);
or U3484 (N_3484,In_2048,In_327);
nor U3485 (N_3485,In_2946,In_2914);
or U3486 (N_3486,In_147,In_2768);
and U3487 (N_3487,In_1292,In_1697);
xnor U3488 (N_3488,In_1353,In_1917);
nand U3489 (N_3489,In_1458,In_2132);
or U3490 (N_3490,In_1558,In_1546);
nand U3491 (N_3491,In_2643,In_1493);
nor U3492 (N_3492,In_786,In_973);
nor U3493 (N_3493,In_647,In_2755);
xnor U3494 (N_3494,In_1937,In_685);
or U3495 (N_3495,In_452,In_1562);
nor U3496 (N_3496,In_2355,In_2011);
or U3497 (N_3497,In_485,In_2682);
and U3498 (N_3498,In_384,In_941);
and U3499 (N_3499,In_376,In_1949);
or U3500 (N_3500,In_311,In_2127);
and U3501 (N_3501,In_1603,In_878);
nand U3502 (N_3502,In_1421,In_1145);
or U3503 (N_3503,In_87,In_572);
nor U3504 (N_3504,In_608,In_2783);
and U3505 (N_3505,In_1178,In_2283);
nand U3506 (N_3506,In_1684,In_1430);
or U3507 (N_3507,In_18,In_1889);
nor U3508 (N_3508,In_85,In_1570);
or U3509 (N_3509,In_230,In_1375);
or U3510 (N_3510,In_2171,In_1877);
nand U3511 (N_3511,In_2281,In_994);
and U3512 (N_3512,In_1874,In_2118);
and U3513 (N_3513,In_960,In_1929);
xnor U3514 (N_3514,In_2132,In_325);
nand U3515 (N_3515,In_1714,In_1506);
or U3516 (N_3516,In_1734,In_2196);
nor U3517 (N_3517,In_1353,In_2935);
nand U3518 (N_3518,In_1582,In_434);
or U3519 (N_3519,In_2331,In_1291);
nand U3520 (N_3520,In_2770,In_1239);
or U3521 (N_3521,In_1581,In_1517);
nand U3522 (N_3522,In_591,In_1263);
nand U3523 (N_3523,In_589,In_1421);
and U3524 (N_3524,In_874,In_420);
nor U3525 (N_3525,In_2857,In_2874);
nor U3526 (N_3526,In_351,In_326);
and U3527 (N_3527,In_2693,In_487);
nand U3528 (N_3528,In_275,In_2779);
and U3529 (N_3529,In_2858,In_2088);
or U3530 (N_3530,In_2063,In_1066);
nand U3531 (N_3531,In_1156,In_41);
nand U3532 (N_3532,In_2389,In_581);
or U3533 (N_3533,In_2016,In_210);
nor U3534 (N_3534,In_247,In_268);
nand U3535 (N_3535,In_1811,In_861);
and U3536 (N_3536,In_396,In_292);
and U3537 (N_3537,In_2260,In_1340);
nand U3538 (N_3538,In_937,In_2089);
nor U3539 (N_3539,In_2678,In_1715);
nand U3540 (N_3540,In_2621,In_1943);
and U3541 (N_3541,In_731,In_310);
nand U3542 (N_3542,In_2403,In_2445);
xor U3543 (N_3543,In_1811,In_1142);
nor U3544 (N_3544,In_2092,In_1712);
and U3545 (N_3545,In_310,In_1799);
nand U3546 (N_3546,In_2899,In_2428);
and U3547 (N_3547,In_1682,In_1993);
nor U3548 (N_3548,In_424,In_2306);
nand U3549 (N_3549,In_844,In_1882);
xnor U3550 (N_3550,In_78,In_504);
and U3551 (N_3551,In_2317,In_1810);
nor U3552 (N_3552,In_1305,In_2954);
nor U3553 (N_3553,In_1008,In_997);
and U3554 (N_3554,In_1170,In_2863);
nand U3555 (N_3555,In_2214,In_1057);
and U3556 (N_3556,In_1730,In_2294);
nor U3557 (N_3557,In_690,In_1226);
and U3558 (N_3558,In_972,In_2671);
nor U3559 (N_3559,In_1455,In_1340);
or U3560 (N_3560,In_591,In_267);
xnor U3561 (N_3561,In_607,In_2026);
and U3562 (N_3562,In_1697,In_1879);
nand U3563 (N_3563,In_2423,In_1470);
nor U3564 (N_3564,In_1668,In_1950);
nor U3565 (N_3565,In_587,In_2775);
nand U3566 (N_3566,In_2760,In_633);
nor U3567 (N_3567,In_787,In_837);
or U3568 (N_3568,In_2943,In_38);
or U3569 (N_3569,In_1534,In_822);
nand U3570 (N_3570,In_56,In_2855);
and U3571 (N_3571,In_2598,In_1263);
and U3572 (N_3572,In_1057,In_848);
nand U3573 (N_3573,In_1921,In_86);
nor U3574 (N_3574,In_1604,In_2752);
nor U3575 (N_3575,In_1651,In_1595);
or U3576 (N_3576,In_2617,In_1171);
nor U3577 (N_3577,In_453,In_2996);
and U3578 (N_3578,In_269,In_2017);
nand U3579 (N_3579,In_1684,In_579);
or U3580 (N_3580,In_1011,In_2955);
nor U3581 (N_3581,In_679,In_448);
nor U3582 (N_3582,In_2848,In_642);
and U3583 (N_3583,In_781,In_2172);
xor U3584 (N_3584,In_811,In_672);
and U3585 (N_3585,In_1857,In_2558);
nor U3586 (N_3586,In_1716,In_2837);
or U3587 (N_3587,In_924,In_2036);
nor U3588 (N_3588,In_2900,In_135);
xor U3589 (N_3589,In_746,In_412);
and U3590 (N_3590,In_2298,In_2741);
or U3591 (N_3591,In_1028,In_214);
or U3592 (N_3592,In_2066,In_343);
or U3593 (N_3593,In_2479,In_1375);
nor U3594 (N_3594,In_2517,In_1365);
nor U3595 (N_3595,In_1730,In_1489);
xnor U3596 (N_3596,In_75,In_379);
and U3597 (N_3597,In_956,In_2085);
and U3598 (N_3598,In_2742,In_696);
or U3599 (N_3599,In_2770,In_1811);
nand U3600 (N_3600,In_704,In_2854);
nor U3601 (N_3601,In_1431,In_1144);
and U3602 (N_3602,In_1121,In_962);
nand U3603 (N_3603,In_486,In_1774);
nand U3604 (N_3604,In_1611,In_1277);
nor U3605 (N_3605,In_2742,In_201);
nand U3606 (N_3606,In_1729,In_742);
nand U3607 (N_3607,In_1207,In_1008);
nor U3608 (N_3608,In_1679,In_1683);
xor U3609 (N_3609,In_1426,In_1381);
nand U3610 (N_3610,In_2565,In_1230);
or U3611 (N_3611,In_652,In_2838);
nor U3612 (N_3612,In_598,In_1673);
nand U3613 (N_3613,In_1016,In_1179);
and U3614 (N_3614,In_2348,In_868);
nand U3615 (N_3615,In_1123,In_318);
and U3616 (N_3616,In_1219,In_2838);
xor U3617 (N_3617,In_1425,In_155);
or U3618 (N_3618,In_376,In_1283);
nor U3619 (N_3619,In_289,In_794);
nand U3620 (N_3620,In_1791,In_2790);
nor U3621 (N_3621,In_2231,In_1306);
and U3622 (N_3622,In_497,In_711);
nand U3623 (N_3623,In_814,In_1521);
and U3624 (N_3624,In_2345,In_2069);
nand U3625 (N_3625,In_1448,In_458);
nand U3626 (N_3626,In_831,In_608);
nor U3627 (N_3627,In_489,In_1882);
and U3628 (N_3628,In_1762,In_137);
or U3629 (N_3629,In_2380,In_2842);
and U3630 (N_3630,In_1766,In_2987);
or U3631 (N_3631,In_2372,In_29);
nand U3632 (N_3632,In_1190,In_2458);
or U3633 (N_3633,In_2696,In_690);
nor U3634 (N_3634,In_2908,In_1363);
nand U3635 (N_3635,In_2918,In_1161);
and U3636 (N_3636,In_244,In_1705);
or U3637 (N_3637,In_1975,In_2733);
nand U3638 (N_3638,In_2508,In_632);
xor U3639 (N_3639,In_1078,In_480);
or U3640 (N_3640,In_1673,In_2332);
and U3641 (N_3641,In_315,In_265);
and U3642 (N_3642,In_1874,In_291);
nor U3643 (N_3643,In_1597,In_231);
nor U3644 (N_3644,In_626,In_413);
nor U3645 (N_3645,In_2774,In_468);
nor U3646 (N_3646,In_1205,In_707);
or U3647 (N_3647,In_2098,In_2114);
or U3648 (N_3648,In_1400,In_531);
or U3649 (N_3649,In_1500,In_1054);
nand U3650 (N_3650,In_2487,In_614);
and U3651 (N_3651,In_343,In_341);
nand U3652 (N_3652,In_420,In_1764);
nand U3653 (N_3653,In_1038,In_2383);
and U3654 (N_3654,In_1289,In_1475);
xor U3655 (N_3655,In_1197,In_955);
and U3656 (N_3656,In_2603,In_682);
and U3657 (N_3657,In_1146,In_2304);
and U3658 (N_3658,In_2832,In_433);
or U3659 (N_3659,In_2920,In_997);
or U3660 (N_3660,In_1487,In_488);
nor U3661 (N_3661,In_1986,In_2163);
nand U3662 (N_3662,In_963,In_1967);
nand U3663 (N_3663,In_307,In_895);
nor U3664 (N_3664,In_2121,In_1638);
nor U3665 (N_3665,In_340,In_2410);
nand U3666 (N_3666,In_2361,In_1926);
and U3667 (N_3667,In_802,In_2820);
nor U3668 (N_3668,In_1139,In_2248);
and U3669 (N_3669,In_2054,In_59);
nand U3670 (N_3670,In_966,In_2577);
nand U3671 (N_3671,In_2988,In_847);
or U3672 (N_3672,In_844,In_631);
or U3673 (N_3673,In_1111,In_1835);
nor U3674 (N_3674,In_2025,In_2689);
and U3675 (N_3675,In_1011,In_24);
nand U3676 (N_3676,In_1219,In_2344);
or U3677 (N_3677,In_431,In_2599);
nor U3678 (N_3678,In_155,In_2573);
or U3679 (N_3679,In_1545,In_375);
or U3680 (N_3680,In_2211,In_1517);
and U3681 (N_3681,In_836,In_2891);
or U3682 (N_3682,In_2524,In_1599);
nor U3683 (N_3683,In_485,In_1695);
xor U3684 (N_3684,In_705,In_2172);
or U3685 (N_3685,In_839,In_535);
or U3686 (N_3686,In_2082,In_600);
xor U3687 (N_3687,In_1177,In_918);
nor U3688 (N_3688,In_2766,In_1572);
nand U3689 (N_3689,In_208,In_2663);
nor U3690 (N_3690,In_2763,In_2120);
or U3691 (N_3691,In_2003,In_1041);
nor U3692 (N_3692,In_2099,In_1347);
xnor U3693 (N_3693,In_1698,In_767);
and U3694 (N_3694,In_263,In_1258);
and U3695 (N_3695,In_1789,In_449);
and U3696 (N_3696,In_338,In_356);
nor U3697 (N_3697,In_1621,In_2930);
xnor U3698 (N_3698,In_1582,In_1586);
and U3699 (N_3699,In_438,In_934);
and U3700 (N_3700,In_689,In_725);
nand U3701 (N_3701,In_1060,In_2257);
and U3702 (N_3702,In_2610,In_350);
or U3703 (N_3703,In_1303,In_428);
nand U3704 (N_3704,In_2938,In_2607);
and U3705 (N_3705,In_1619,In_2495);
or U3706 (N_3706,In_2047,In_439);
nor U3707 (N_3707,In_2491,In_562);
nand U3708 (N_3708,In_347,In_1573);
and U3709 (N_3709,In_691,In_700);
nand U3710 (N_3710,In_523,In_1247);
and U3711 (N_3711,In_940,In_2728);
and U3712 (N_3712,In_1030,In_551);
and U3713 (N_3713,In_1107,In_2810);
nor U3714 (N_3714,In_2636,In_1934);
nor U3715 (N_3715,In_187,In_852);
nor U3716 (N_3716,In_491,In_2985);
or U3717 (N_3717,In_1438,In_2836);
and U3718 (N_3718,In_2743,In_2419);
or U3719 (N_3719,In_2285,In_1454);
and U3720 (N_3720,In_774,In_466);
and U3721 (N_3721,In_783,In_2736);
or U3722 (N_3722,In_1161,In_2359);
and U3723 (N_3723,In_1375,In_2565);
or U3724 (N_3724,In_1692,In_609);
nand U3725 (N_3725,In_246,In_1725);
xnor U3726 (N_3726,In_539,In_415);
nor U3727 (N_3727,In_2455,In_1886);
or U3728 (N_3728,In_286,In_2047);
or U3729 (N_3729,In_2617,In_1289);
and U3730 (N_3730,In_2175,In_2070);
nand U3731 (N_3731,In_2628,In_2941);
or U3732 (N_3732,In_1334,In_2109);
nand U3733 (N_3733,In_1998,In_621);
or U3734 (N_3734,In_2387,In_1217);
or U3735 (N_3735,In_2777,In_141);
nor U3736 (N_3736,In_1501,In_337);
and U3737 (N_3737,In_1634,In_1126);
nor U3738 (N_3738,In_2691,In_1252);
and U3739 (N_3739,In_2456,In_57);
or U3740 (N_3740,In_724,In_2714);
or U3741 (N_3741,In_19,In_2139);
and U3742 (N_3742,In_1113,In_2188);
or U3743 (N_3743,In_337,In_700);
or U3744 (N_3744,In_1719,In_1021);
or U3745 (N_3745,In_2926,In_1207);
nand U3746 (N_3746,In_963,In_2599);
nand U3747 (N_3747,In_1550,In_2474);
nor U3748 (N_3748,In_2475,In_1937);
and U3749 (N_3749,In_2321,In_2548);
nand U3750 (N_3750,In_1356,In_1730);
or U3751 (N_3751,In_2361,In_2833);
nand U3752 (N_3752,In_1703,In_174);
nor U3753 (N_3753,In_2335,In_2735);
xor U3754 (N_3754,In_1014,In_41);
nand U3755 (N_3755,In_147,In_2955);
and U3756 (N_3756,In_1158,In_47);
nor U3757 (N_3757,In_786,In_1549);
and U3758 (N_3758,In_1557,In_1866);
nor U3759 (N_3759,In_461,In_2099);
or U3760 (N_3760,In_169,In_1531);
nand U3761 (N_3761,In_584,In_1496);
nand U3762 (N_3762,In_210,In_2495);
nand U3763 (N_3763,In_2758,In_226);
or U3764 (N_3764,In_2731,In_293);
nor U3765 (N_3765,In_1192,In_2946);
nor U3766 (N_3766,In_2416,In_64);
and U3767 (N_3767,In_2191,In_322);
nand U3768 (N_3768,In_2158,In_960);
nor U3769 (N_3769,In_792,In_2135);
nand U3770 (N_3770,In_164,In_410);
or U3771 (N_3771,In_785,In_51);
nand U3772 (N_3772,In_1303,In_2063);
and U3773 (N_3773,In_1099,In_1938);
nand U3774 (N_3774,In_691,In_2236);
and U3775 (N_3775,In_1113,In_2839);
nand U3776 (N_3776,In_2789,In_160);
nand U3777 (N_3777,In_1168,In_1045);
nand U3778 (N_3778,In_233,In_324);
or U3779 (N_3779,In_2458,In_2480);
or U3780 (N_3780,In_70,In_1131);
nand U3781 (N_3781,In_2482,In_917);
and U3782 (N_3782,In_238,In_1706);
and U3783 (N_3783,In_1233,In_2095);
and U3784 (N_3784,In_606,In_2502);
xnor U3785 (N_3785,In_2756,In_2237);
and U3786 (N_3786,In_1384,In_2227);
and U3787 (N_3787,In_1101,In_375);
nand U3788 (N_3788,In_887,In_2962);
or U3789 (N_3789,In_1831,In_660);
or U3790 (N_3790,In_1995,In_1974);
xnor U3791 (N_3791,In_1187,In_1771);
or U3792 (N_3792,In_2530,In_1166);
or U3793 (N_3793,In_2559,In_2647);
and U3794 (N_3794,In_673,In_1150);
nor U3795 (N_3795,In_2746,In_2195);
xnor U3796 (N_3796,In_2906,In_1167);
nand U3797 (N_3797,In_1781,In_1027);
xnor U3798 (N_3798,In_903,In_2752);
nand U3799 (N_3799,In_481,In_2708);
nand U3800 (N_3800,In_56,In_1922);
xor U3801 (N_3801,In_1411,In_1468);
nand U3802 (N_3802,In_1057,In_2375);
and U3803 (N_3803,In_168,In_2103);
or U3804 (N_3804,In_837,In_706);
and U3805 (N_3805,In_2153,In_1891);
nand U3806 (N_3806,In_2399,In_1690);
nand U3807 (N_3807,In_1919,In_2275);
and U3808 (N_3808,In_1150,In_1670);
or U3809 (N_3809,In_1792,In_389);
nand U3810 (N_3810,In_492,In_2520);
nand U3811 (N_3811,In_2224,In_1886);
or U3812 (N_3812,In_923,In_107);
nor U3813 (N_3813,In_812,In_814);
or U3814 (N_3814,In_1091,In_2100);
or U3815 (N_3815,In_303,In_593);
or U3816 (N_3816,In_1449,In_2018);
nand U3817 (N_3817,In_430,In_1960);
nor U3818 (N_3818,In_169,In_2087);
nand U3819 (N_3819,In_2,In_19);
nand U3820 (N_3820,In_2173,In_1147);
nand U3821 (N_3821,In_1174,In_989);
and U3822 (N_3822,In_1697,In_2655);
and U3823 (N_3823,In_870,In_1263);
nand U3824 (N_3824,In_1537,In_24);
and U3825 (N_3825,In_696,In_57);
xnor U3826 (N_3826,In_1833,In_1295);
nor U3827 (N_3827,In_746,In_1500);
nand U3828 (N_3828,In_1474,In_1604);
nor U3829 (N_3829,In_123,In_540);
xor U3830 (N_3830,In_382,In_1034);
or U3831 (N_3831,In_909,In_2272);
xnor U3832 (N_3832,In_447,In_515);
and U3833 (N_3833,In_1164,In_2051);
or U3834 (N_3834,In_148,In_2784);
xnor U3835 (N_3835,In_1814,In_67);
and U3836 (N_3836,In_1682,In_52);
and U3837 (N_3837,In_1012,In_629);
and U3838 (N_3838,In_872,In_1047);
or U3839 (N_3839,In_1345,In_2184);
xor U3840 (N_3840,In_2683,In_2294);
nand U3841 (N_3841,In_762,In_53);
or U3842 (N_3842,In_1196,In_1331);
nor U3843 (N_3843,In_2209,In_737);
or U3844 (N_3844,In_2158,In_208);
and U3845 (N_3845,In_1835,In_2209);
nor U3846 (N_3846,In_1220,In_201);
or U3847 (N_3847,In_2160,In_2063);
nor U3848 (N_3848,In_1240,In_1605);
xor U3849 (N_3849,In_581,In_685);
xor U3850 (N_3850,In_2208,In_2696);
and U3851 (N_3851,In_1502,In_903);
and U3852 (N_3852,In_1143,In_990);
nand U3853 (N_3853,In_730,In_33);
nand U3854 (N_3854,In_2347,In_414);
nand U3855 (N_3855,In_761,In_1451);
nor U3856 (N_3856,In_2036,In_105);
and U3857 (N_3857,In_809,In_1190);
nor U3858 (N_3858,In_2607,In_2478);
and U3859 (N_3859,In_2331,In_2114);
or U3860 (N_3860,In_385,In_2029);
nand U3861 (N_3861,In_614,In_914);
and U3862 (N_3862,In_330,In_1539);
nor U3863 (N_3863,In_38,In_803);
and U3864 (N_3864,In_517,In_2337);
nor U3865 (N_3865,In_2454,In_1779);
and U3866 (N_3866,In_1353,In_1434);
nor U3867 (N_3867,In_250,In_2350);
or U3868 (N_3868,In_1202,In_2266);
and U3869 (N_3869,In_995,In_2235);
or U3870 (N_3870,In_818,In_1813);
nor U3871 (N_3871,In_26,In_2882);
nand U3872 (N_3872,In_843,In_453);
nand U3873 (N_3873,In_2851,In_2435);
and U3874 (N_3874,In_1886,In_2243);
nand U3875 (N_3875,In_796,In_1518);
and U3876 (N_3876,In_2702,In_2451);
nand U3877 (N_3877,In_2397,In_1090);
or U3878 (N_3878,In_2918,In_790);
nor U3879 (N_3879,In_1892,In_1537);
and U3880 (N_3880,In_195,In_1741);
nand U3881 (N_3881,In_1432,In_1506);
nand U3882 (N_3882,In_323,In_554);
or U3883 (N_3883,In_41,In_1658);
and U3884 (N_3884,In_1063,In_2030);
nor U3885 (N_3885,In_50,In_709);
nand U3886 (N_3886,In_2009,In_197);
and U3887 (N_3887,In_597,In_1565);
or U3888 (N_3888,In_2131,In_900);
xnor U3889 (N_3889,In_33,In_2719);
nand U3890 (N_3890,In_1899,In_2184);
and U3891 (N_3891,In_1160,In_201);
and U3892 (N_3892,In_2887,In_1546);
xnor U3893 (N_3893,In_132,In_2122);
nor U3894 (N_3894,In_1847,In_969);
nor U3895 (N_3895,In_1951,In_2966);
or U3896 (N_3896,In_1191,In_1781);
and U3897 (N_3897,In_251,In_701);
nand U3898 (N_3898,In_483,In_2843);
and U3899 (N_3899,In_2861,In_2746);
and U3900 (N_3900,In_1377,In_34);
nor U3901 (N_3901,In_1398,In_1920);
and U3902 (N_3902,In_23,In_1226);
xnor U3903 (N_3903,In_2776,In_970);
xnor U3904 (N_3904,In_2743,In_218);
xnor U3905 (N_3905,In_2108,In_1336);
and U3906 (N_3906,In_46,In_2454);
xor U3907 (N_3907,In_848,In_1691);
xor U3908 (N_3908,In_2559,In_43);
and U3909 (N_3909,In_745,In_1923);
and U3910 (N_3910,In_564,In_2585);
nor U3911 (N_3911,In_746,In_1063);
nor U3912 (N_3912,In_779,In_2884);
nand U3913 (N_3913,In_287,In_2092);
nor U3914 (N_3914,In_2542,In_1864);
and U3915 (N_3915,In_395,In_1911);
xor U3916 (N_3916,In_1529,In_2165);
nor U3917 (N_3917,In_1175,In_2495);
xor U3918 (N_3918,In_587,In_2421);
and U3919 (N_3919,In_2245,In_927);
or U3920 (N_3920,In_2089,In_1741);
nor U3921 (N_3921,In_2377,In_2856);
nor U3922 (N_3922,In_187,In_2352);
or U3923 (N_3923,In_1527,In_1960);
and U3924 (N_3924,In_2197,In_483);
nand U3925 (N_3925,In_652,In_1495);
or U3926 (N_3926,In_2655,In_2386);
nand U3927 (N_3927,In_2008,In_2677);
and U3928 (N_3928,In_232,In_432);
xnor U3929 (N_3929,In_1743,In_1709);
and U3930 (N_3930,In_1835,In_1709);
or U3931 (N_3931,In_2527,In_861);
xnor U3932 (N_3932,In_1834,In_326);
or U3933 (N_3933,In_462,In_470);
nor U3934 (N_3934,In_1243,In_1190);
nor U3935 (N_3935,In_826,In_2718);
and U3936 (N_3936,In_2865,In_670);
and U3937 (N_3937,In_523,In_1808);
nor U3938 (N_3938,In_2925,In_1743);
nor U3939 (N_3939,In_1252,In_537);
xor U3940 (N_3940,In_2972,In_2307);
and U3941 (N_3941,In_1531,In_2475);
nor U3942 (N_3942,In_1073,In_86);
and U3943 (N_3943,In_2926,In_1045);
nand U3944 (N_3944,In_2184,In_73);
nand U3945 (N_3945,In_1879,In_2466);
or U3946 (N_3946,In_2052,In_2429);
nand U3947 (N_3947,In_705,In_191);
nand U3948 (N_3948,In_435,In_462);
nor U3949 (N_3949,In_2658,In_2117);
xnor U3950 (N_3950,In_2195,In_1929);
nand U3951 (N_3951,In_401,In_2225);
xnor U3952 (N_3952,In_127,In_2440);
nor U3953 (N_3953,In_2340,In_1054);
and U3954 (N_3954,In_994,In_2796);
or U3955 (N_3955,In_2802,In_2652);
nor U3956 (N_3956,In_1497,In_343);
or U3957 (N_3957,In_1052,In_1459);
nand U3958 (N_3958,In_1508,In_2887);
nor U3959 (N_3959,In_2105,In_937);
or U3960 (N_3960,In_383,In_852);
and U3961 (N_3961,In_1773,In_32);
nor U3962 (N_3962,In_2032,In_1537);
nand U3963 (N_3963,In_1206,In_225);
nand U3964 (N_3964,In_1838,In_2463);
nand U3965 (N_3965,In_1891,In_704);
nor U3966 (N_3966,In_1647,In_36);
or U3967 (N_3967,In_254,In_266);
nor U3968 (N_3968,In_1258,In_2170);
and U3969 (N_3969,In_2926,In_1964);
or U3970 (N_3970,In_336,In_645);
or U3971 (N_3971,In_1361,In_892);
nor U3972 (N_3972,In_1533,In_394);
or U3973 (N_3973,In_1001,In_1370);
or U3974 (N_3974,In_1060,In_378);
or U3975 (N_3975,In_1180,In_1704);
nand U3976 (N_3976,In_2326,In_746);
nand U3977 (N_3977,In_760,In_1127);
or U3978 (N_3978,In_1642,In_2724);
or U3979 (N_3979,In_1139,In_477);
nand U3980 (N_3980,In_1832,In_931);
nor U3981 (N_3981,In_2419,In_1139);
xnor U3982 (N_3982,In_222,In_1570);
or U3983 (N_3983,In_754,In_462);
xor U3984 (N_3984,In_2109,In_449);
nand U3985 (N_3985,In_481,In_2648);
and U3986 (N_3986,In_2746,In_1793);
xnor U3987 (N_3987,In_909,In_1882);
nand U3988 (N_3988,In_2670,In_2480);
and U3989 (N_3989,In_2042,In_2046);
nor U3990 (N_3990,In_1435,In_103);
nor U3991 (N_3991,In_1963,In_917);
and U3992 (N_3992,In_748,In_2329);
or U3993 (N_3993,In_1813,In_364);
nand U3994 (N_3994,In_853,In_1371);
or U3995 (N_3995,In_2544,In_2337);
or U3996 (N_3996,In_1131,In_478);
nor U3997 (N_3997,In_371,In_405);
and U3998 (N_3998,In_983,In_2494);
and U3999 (N_3999,In_339,In_2659);
nand U4000 (N_4000,In_1203,In_1782);
and U4001 (N_4001,In_1209,In_2084);
xnor U4002 (N_4002,In_229,In_919);
or U4003 (N_4003,In_2576,In_1124);
or U4004 (N_4004,In_2352,In_2213);
nand U4005 (N_4005,In_1739,In_904);
or U4006 (N_4006,In_1470,In_921);
nand U4007 (N_4007,In_977,In_289);
and U4008 (N_4008,In_235,In_2776);
nand U4009 (N_4009,In_1364,In_2353);
nand U4010 (N_4010,In_1611,In_628);
or U4011 (N_4011,In_1679,In_1868);
nor U4012 (N_4012,In_969,In_2966);
nor U4013 (N_4013,In_2193,In_2253);
nor U4014 (N_4014,In_2208,In_1429);
xnor U4015 (N_4015,In_217,In_145);
or U4016 (N_4016,In_718,In_2460);
and U4017 (N_4017,In_1988,In_1727);
and U4018 (N_4018,In_2322,In_2140);
and U4019 (N_4019,In_1931,In_2902);
nor U4020 (N_4020,In_897,In_2746);
or U4021 (N_4021,In_1382,In_979);
nand U4022 (N_4022,In_2727,In_2572);
nand U4023 (N_4023,In_2765,In_130);
nand U4024 (N_4024,In_2447,In_2663);
nor U4025 (N_4025,In_1316,In_1580);
or U4026 (N_4026,In_1296,In_2404);
or U4027 (N_4027,In_548,In_1725);
nand U4028 (N_4028,In_2336,In_1551);
nor U4029 (N_4029,In_376,In_2776);
nor U4030 (N_4030,In_1398,In_378);
or U4031 (N_4031,In_611,In_1632);
or U4032 (N_4032,In_2848,In_1600);
and U4033 (N_4033,In_2938,In_646);
or U4034 (N_4034,In_761,In_125);
and U4035 (N_4035,In_987,In_608);
and U4036 (N_4036,In_73,In_2042);
and U4037 (N_4037,In_2882,In_25);
and U4038 (N_4038,In_2617,In_2467);
and U4039 (N_4039,In_2328,In_1980);
or U4040 (N_4040,In_1580,In_2553);
nand U4041 (N_4041,In_1262,In_1041);
nor U4042 (N_4042,In_1943,In_2776);
and U4043 (N_4043,In_2876,In_842);
or U4044 (N_4044,In_1630,In_2024);
and U4045 (N_4045,In_1937,In_321);
nor U4046 (N_4046,In_745,In_2543);
or U4047 (N_4047,In_1374,In_1252);
nor U4048 (N_4048,In_776,In_2081);
xor U4049 (N_4049,In_2907,In_1707);
nand U4050 (N_4050,In_462,In_1161);
nor U4051 (N_4051,In_173,In_1371);
nor U4052 (N_4052,In_1872,In_415);
nor U4053 (N_4053,In_1953,In_1754);
or U4054 (N_4054,In_2220,In_523);
nand U4055 (N_4055,In_1724,In_2850);
and U4056 (N_4056,In_2642,In_1880);
nand U4057 (N_4057,In_1950,In_516);
or U4058 (N_4058,In_2773,In_1707);
and U4059 (N_4059,In_111,In_1232);
nand U4060 (N_4060,In_2798,In_2774);
nor U4061 (N_4061,In_2696,In_2297);
nand U4062 (N_4062,In_2138,In_2512);
nand U4063 (N_4063,In_521,In_2314);
or U4064 (N_4064,In_1570,In_2830);
or U4065 (N_4065,In_2060,In_771);
and U4066 (N_4066,In_153,In_317);
nand U4067 (N_4067,In_1658,In_1351);
xor U4068 (N_4068,In_2454,In_2796);
or U4069 (N_4069,In_2994,In_1768);
nor U4070 (N_4070,In_2668,In_2820);
nor U4071 (N_4071,In_2186,In_2366);
and U4072 (N_4072,In_1960,In_2825);
nor U4073 (N_4073,In_2652,In_1807);
or U4074 (N_4074,In_1454,In_1881);
nor U4075 (N_4075,In_2314,In_1456);
or U4076 (N_4076,In_2462,In_617);
and U4077 (N_4077,In_2192,In_803);
or U4078 (N_4078,In_969,In_638);
or U4079 (N_4079,In_587,In_132);
or U4080 (N_4080,In_1212,In_1373);
or U4081 (N_4081,In_2991,In_64);
nor U4082 (N_4082,In_1968,In_2943);
or U4083 (N_4083,In_1330,In_1187);
nand U4084 (N_4084,In_187,In_1284);
or U4085 (N_4085,In_2750,In_499);
and U4086 (N_4086,In_0,In_2612);
nor U4087 (N_4087,In_113,In_2941);
and U4088 (N_4088,In_306,In_373);
or U4089 (N_4089,In_2146,In_2554);
or U4090 (N_4090,In_2599,In_1098);
nand U4091 (N_4091,In_2578,In_1737);
nor U4092 (N_4092,In_2836,In_929);
or U4093 (N_4093,In_1679,In_2432);
nand U4094 (N_4094,In_2480,In_2060);
nand U4095 (N_4095,In_1587,In_81);
nor U4096 (N_4096,In_1605,In_268);
and U4097 (N_4097,In_1942,In_266);
and U4098 (N_4098,In_816,In_1114);
and U4099 (N_4099,In_111,In_2533);
xnor U4100 (N_4100,In_1922,In_817);
nor U4101 (N_4101,In_1002,In_1416);
nand U4102 (N_4102,In_669,In_1625);
nor U4103 (N_4103,In_317,In_845);
and U4104 (N_4104,In_811,In_904);
nor U4105 (N_4105,In_2980,In_1282);
nand U4106 (N_4106,In_2803,In_200);
or U4107 (N_4107,In_2887,In_1987);
nor U4108 (N_4108,In_518,In_2443);
or U4109 (N_4109,In_1495,In_1824);
nand U4110 (N_4110,In_878,In_1475);
and U4111 (N_4111,In_1148,In_416);
nor U4112 (N_4112,In_2488,In_11);
or U4113 (N_4113,In_737,In_1680);
or U4114 (N_4114,In_256,In_578);
or U4115 (N_4115,In_2840,In_367);
xnor U4116 (N_4116,In_1762,In_2269);
nand U4117 (N_4117,In_2290,In_1705);
nor U4118 (N_4118,In_1692,In_2724);
and U4119 (N_4119,In_1908,In_1986);
or U4120 (N_4120,In_1111,In_1864);
nand U4121 (N_4121,In_2904,In_1144);
nor U4122 (N_4122,In_784,In_2805);
nor U4123 (N_4123,In_1565,In_1153);
xnor U4124 (N_4124,In_500,In_305);
nand U4125 (N_4125,In_1254,In_1974);
xor U4126 (N_4126,In_1106,In_653);
xor U4127 (N_4127,In_2295,In_2);
nand U4128 (N_4128,In_369,In_192);
nor U4129 (N_4129,In_2213,In_482);
and U4130 (N_4130,In_1641,In_1680);
and U4131 (N_4131,In_2123,In_504);
nand U4132 (N_4132,In_129,In_1585);
nor U4133 (N_4133,In_2954,In_1355);
nand U4134 (N_4134,In_1781,In_2592);
or U4135 (N_4135,In_1722,In_1549);
or U4136 (N_4136,In_1569,In_1080);
nand U4137 (N_4137,In_144,In_1227);
nor U4138 (N_4138,In_2910,In_1326);
nor U4139 (N_4139,In_2200,In_2508);
nor U4140 (N_4140,In_1887,In_1671);
nor U4141 (N_4141,In_627,In_1751);
nor U4142 (N_4142,In_2340,In_728);
nand U4143 (N_4143,In_2502,In_1569);
nand U4144 (N_4144,In_927,In_2020);
nand U4145 (N_4145,In_1289,In_2487);
and U4146 (N_4146,In_2210,In_243);
or U4147 (N_4147,In_2580,In_2505);
nand U4148 (N_4148,In_1796,In_2051);
or U4149 (N_4149,In_1817,In_312);
nor U4150 (N_4150,In_2488,In_2680);
and U4151 (N_4151,In_459,In_2639);
or U4152 (N_4152,In_2935,In_2136);
nor U4153 (N_4153,In_601,In_1209);
nor U4154 (N_4154,In_2583,In_2350);
and U4155 (N_4155,In_1577,In_2437);
nand U4156 (N_4156,In_787,In_2045);
and U4157 (N_4157,In_2360,In_521);
and U4158 (N_4158,In_2008,In_2067);
or U4159 (N_4159,In_1826,In_2942);
nand U4160 (N_4160,In_2727,In_1445);
nor U4161 (N_4161,In_1030,In_1169);
nand U4162 (N_4162,In_1726,In_1600);
and U4163 (N_4163,In_770,In_1152);
nor U4164 (N_4164,In_399,In_1629);
or U4165 (N_4165,In_1155,In_2211);
and U4166 (N_4166,In_2329,In_793);
nor U4167 (N_4167,In_838,In_2599);
and U4168 (N_4168,In_303,In_970);
or U4169 (N_4169,In_632,In_55);
or U4170 (N_4170,In_1955,In_2456);
nand U4171 (N_4171,In_237,In_1100);
or U4172 (N_4172,In_1131,In_1523);
nor U4173 (N_4173,In_2966,In_2072);
nor U4174 (N_4174,In_765,In_2623);
nand U4175 (N_4175,In_363,In_455);
nand U4176 (N_4176,In_1909,In_2389);
and U4177 (N_4177,In_96,In_1136);
nor U4178 (N_4178,In_2467,In_1288);
and U4179 (N_4179,In_106,In_1161);
and U4180 (N_4180,In_1692,In_666);
or U4181 (N_4181,In_1686,In_1568);
and U4182 (N_4182,In_1385,In_947);
and U4183 (N_4183,In_1838,In_2968);
nand U4184 (N_4184,In_1809,In_2831);
or U4185 (N_4185,In_471,In_2375);
or U4186 (N_4186,In_823,In_1444);
and U4187 (N_4187,In_2089,In_1311);
xnor U4188 (N_4188,In_720,In_2141);
nand U4189 (N_4189,In_592,In_1462);
or U4190 (N_4190,In_68,In_1655);
nand U4191 (N_4191,In_2466,In_2808);
and U4192 (N_4192,In_1686,In_2858);
or U4193 (N_4193,In_1454,In_2998);
or U4194 (N_4194,In_1838,In_2362);
nor U4195 (N_4195,In_171,In_1580);
nand U4196 (N_4196,In_2104,In_1339);
or U4197 (N_4197,In_259,In_2519);
nand U4198 (N_4198,In_2693,In_894);
and U4199 (N_4199,In_2491,In_1694);
xnor U4200 (N_4200,In_1756,In_973);
nand U4201 (N_4201,In_1289,In_1360);
and U4202 (N_4202,In_2141,In_2001);
or U4203 (N_4203,In_2311,In_2012);
xnor U4204 (N_4204,In_589,In_2584);
or U4205 (N_4205,In_418,In_1661);
xor U4206 (N_4206,In_558,In_2703);
nand U4207 (N_4207,In_581,In_1231);
or U4208 (N_4208,In_57,In_1765);
or U4209 (N_4209,In_800,In_1058);
nor U4210 (N_4210,In_2242,In_2984);
or U4211 (N_4211,In_2361,In_1561);
or U4212 (N_4212,In_332,In_674);
or U4213 (N_4213,In_299,In_2825);
nor U4214 (N_4214,In_1034,In_1628);
nor U4215 (N_4215,In_2809,In_74);
nand U4216 (N_4216,In_2048,In_949);
or U4217 (N_4217,In_1594,In_1905);
nand U4218 (N_4218,In_395,In_2741);
and U4219 (N_4219,In_587,In_2187);
nor U4220 (N_4220,In_1757,In_2062);
nor U4221 (N_4221,In_744,In_2812);
nand U4222 (N_4222,In_1474,In_1086);
nand U4223 (N_4223,In_900,In_2643);
nor U4224 (N_4224,In_2022,In_400);
nor U4225 (N_4225,In_74,In_2368);
xnor U4226 (N_4226,In_399,In_1403);
or U4227 (N_4227,In_2608,In_2713);
or U4228 (N_4228,In_2093,In_973);
or U4229 (N_4229,In_2757,In_453);
or U4230 (N_4230,In_1567,In_1588);
and U4231 (N_4231,In_6,In_1527);
nand U4232 (N_4232,In_1406,In_672);
and U4233 (N_4233,In_2599,In_1617);
xnor U4234 (N_4234,In_2830,In_1544);
and U4235 (N_4235,In_2712,In_40);
or U4236 (N_4236,In_2155,In_1614);
xor U4237 (N_4237,In_1446,In_1834);
and U4238 (N_4238,In_1294,In_2583);
xnor U4239 (N_4239,In_1980,In_2421);
nand U4240 (N_4240,In_2959,In_1952);
nand U4241 (N_4241,In_877,In_1467);
nor U4242 (N_4242,In_88,In_986);
nor U4243 (N_4243,In_2349,In_1861);
or U4244 (N_4244,In_1351,In_2808);
nor U4245 (N_4245,In_1848,In_995);
and U4246 (N_4246,In_1395,In_1315);
nor U4247 (N_4247,In_2587,In_1485);
and U4248 (N_4248,In_1151,In_732);
or U4249 (N_4249,In_828,In_621);
and U4250 (N_4250,In_2316,In_1405);
xnor U4251 (N_4251,In_1685,In_1418);
or U4252 (N_4252,In_2371,In_2075);
nand U4253 (N_4253,In_1863,In_1649);
xnor U4254 (N_4254,In_2307,In_898);
nand U4255 (N_4255,In_1578,In_105);
xnor U4256 (N_4256,In_1989,In_1785);
and U4257 (N_4257,In_2864,In_1901);
nand U4258 (N_4258,In_465,In_1661);
or U4259 (N_4259,In_19,In_477);
nor U4260 (N_4260,In_2361,In_678);
nand U4261 (N_4261,In_245,In_2438);
and U4262 (N_4262,In_2720,In_460);
xor U4263 (N_4263,In_1972,In_468);
and U4264 (N_4264,In_702,In_160);
nand U4265 (N_4265,In_2560,In_2699);
and U4266 (N_4266,In_1007,In_115);
or U4267 (N_4267,In_2128,In_706);
or U4268 (N_4268,In_2070,In_1659);
nand U4269 (N_4269,In_2733,In_2024);
and U4270 (N_4270,In_435,In_1314);
nand U4271 (N_4271,In_1954,In_1435);
or U4272 (N_4272,In_692,In_1474);
or U4273 (N_4273,In_295,In_711);
xnor U4274 (N_4274,In_1221,In_389);
nand U4275 (N_4275,In_1121,In_2730);
or U4276 (N_4276,In_2111,In_1365);
nor U4277 (N_4277,In_188,In_247);
nor U4278 (N_4278,In_1078,In_2114);
nand U4279 (N_4279,In_2401,In_17);
nor U4280 (N_4280,In_1312,In_942);
or U4281 (N_4281,In_891,In_2577);
xor U4282 (N_4282,In_2849,In_1930);
and U4283 (N_4283,In_2610,In_2681);
nor U4284 (N_4284,In_2731,In_915);
nand U4285 (N_4285,In_163,In_1904);
nand U4286 (N_4286,In_2664,In_82);
and U4287 (N_4287,In_2897,In_2240);
nand U4288 (N_4288,In_2986,In_656);
nor U4289 (N_4289,In_2674,In_2425);
nand U4290 (N_4290,In_2764,In_648);
nand U4291 (N_4291,In_1034,In_502);
nor U4292 (N_4292,In_1356,In_2771);
xnor U4293 (N_4293,In_1197,In_1625);
nand U4294 (N_4294,In_1121,In_2638);
or U4295 (N_4295,In_993,In_742);
nor U4296 (N_4296,In_1426,In_2999);
and U4297 (N_4297,In_1140,In_359);
and U4298 (N_4298,In_936,In_428);
nand U4299 (N_4299,In_2039,In_2248);
and U4300 (N_4300,In_2066,In_183);
or U4301 (N_4301,In_848,In_685);
or U4302 (N_4302,In_459,In_1727);
nor U4303 (N_4303,In_2431,In_2352);
xor U4304 (N_4304,In_1109,In_349);
or U4305 (N_4305,In_2749,In_2792);
or U4306 (N_4306,In_350,In_1998);
xor U4307 (N_4307,In_650,In_1737);
nor U4308 (N_4308,In_564,In_2236);
or U4309 (N_4309,In_2352,In_1073);
and U4310 (N_4310,In_2696,In_263);
nand U4311 (N_4311,In_2872,In_1938);
xor U4312 (N_4312,In_1962,In_1319);
nand U4313 (N_4313,In_2190,In_951);
nand U4314 (N_4314,In_666,In_2853);
nand U4315 (N_4315,In_2190,In_2590);
nor U4316 (N_4316,In_903,In_1828);
nand U4317 (N_4317,In_1578,In_324);
xnor U4318 (N_4318,In_1421,In_1589);
nor U4319 (N_4319,In_1498,In_46);
nor U4320 (N_4320,In_2911,In_88);
or U4321 (N_4321,In_1510,In_726);
nand U4322 (N_4322,In_1027,In_2663);
nand U4323 (N_4323,In_2978,In_1225);
and U4324 (N_4324,In_547,In_2266);
xor U4325 (N_4325,In_947,In_681);
nand U4326 (N_4326,In_484,In_1442);
or U4327 (N_4327,In_2889,In_419);
and U4328 (N_4328,In_730,In_1394);
and U4329 (N_4329,In_158,In_1444);
or U4330 (N_4330,In_799,In_1652);
nor U4331 (N_4331,In_2377,In_1397);
and U4332 (N_4332,In_2433,In_419);
and U4333 (N_4333,In_644,In_525);
and U4334 (N_4334,In_2119,In_1334);
nand U4335 (N_4335,In_2300,In_829);
and U4336 (N_4336,In_1291,In_2244);
and U4337 (N_4337,In_241,In_885);
or U4338 (N_4338,In_2161,In_2702);
nand U4339 (N_4339,In_2147,In_1970);
or U4340 (N_4340,In_2636,In_2898);
or U4341 (N_4341,In_1767,In_1716);
and U4342 (N_4342,In_1367,In_2970);
and U4343 (N_4343,In_199,In_425);
or U4344 (N_4344,In_842,In_716);
nand U4345 (N_4345,In_1534,In_2533);
or U4346 (N_4346,In_2227,In_1411);
and U4347 (N_4347,In_2957,In_490);
or U4348 (N_4348,In_826,In_1560);
and U4349 (N_4349,In_228,In_223);
and U4350 (N_4350,In_1436,In_1135);
nor U4351 (N_4351,In_1410,In_746);
and U4352 (N_4352,In_1627,In_2785);
nand U4353 (N_4353,In_2761,In_2666);
nand U4354 (N_4354,In_2863,In_2521);
or U4355 (N_4355,In_2484,In_330);
nor U4356 (N_4356,In_238,In_2038);
and U4357 (N_4357,In_409,In_2628);
or U4358 (N_4358,In_645,In_839);
and U4359 (N_4359,In_287,In_2628);
nor U4360 (N_4360,In_241,In_1273);
nand U4361 (N_4361,In_552,In_499);
or U4362 (N_4362,In_111,In_2267);
nand U4363 (N_4363,In_1459,In_1441);
and U4364 (N_4364,In_308,In_2854);
or U4365 (N_4365,In_62,In_283);
nor U4366 (N_4366,In_2370,In_1620);
and U4367 (N_4367,In_1159,In_2982);
nor U4368 (N_4368,In_2998,In_1491);
nor U4369 (N_4369,In_132,In_1404);
or U4370 (N_4370,In_676,In_0);
nor U4371 (N_4371,In_2318,In_1626);
xnor U4372 (N_4372,In_2778,In_2718);
and U4373 (N_4373,In_2251,In_1027);
or U4374 (N_4374,In_2860,In_2883);
and U4375 (N_4375,In_334,In_1437);
and U4376 (N_4376,In_793,In_2549);
xor U4377 (N_4377,In_747,In_171);
nand U4378 (N_4378,In_697,In_1831);
and U4379 (N_4379,In_1400,In_1477);
or U4380 (N_4380,In_1992,In_1834);
or U4381 (N_4381,In_2151,In_2384);
nor U4382 (N_4382,In_676,In_997);
and U4383 (N_4383,In_286,In_2386);
or U4384 (N_4384,In_1978,In_2164);
nor U4385 (N_4385,In_2844,In_687);
and U4386 (N_4386,In_1718,In_702);
nor U4387 (N_4387,In_231,In_2989);
or U4388 (N_4388,In_2219,In_259);
and U4389 (N_4389,In_2898,In_2498);
nand U4390 (N_4390,In_2800,In_1140);
nor U4391 (N_4391,In_2815,In_352);
nand U4392 (N_4392,In_2132,In_2050);
nand U4393 (N_4393,In_2600,In_300);
nand U4394 (N_4394,In_1488,In_746);
or U4395 (N_4395,In_2970,In_789);
or U4396 (N_4396,In_293,In_1550);
and U4397 (N_4397,In_1840,In_2305);
nor U4398 (N_4398,In_2059,In_2647);
nor U4399 (N_4399,In_1152,In_1802);
or U4400 (N_4400,In_691,In_139);
nand U4401 (N_4401,In_1652,In_1568);
nor U4402 (N_4402,In_931,In_986);
and U4403 (N_4403,In_2746,In_1675);
nor U4404 (N_4404,In_2550,In_2528);
nor U4405 (N_4405,In_726,In_2474);
xor U4406 (N_4406,In_102,In_2594);
nand U4407 (N_4407,In_2621,In_1865);
or U4408 (N_4408,In_2940,In_2169);
and U4409 (N_4409,In_2449,In_2080);
and U4410 (N_4410,In_2485,In_2423);
nand U4411 (N_4411,In_146,In_2084);
or U4412 (N_4412,In_1563,In_934);
or U4413 (N_4413,In_290,In_2852);
and U4414 (N_4414,In_341,In_2748);
nor U4415 (N_4415,In_1565,In_2160);
nand U4416 (N_4416,In_1749,In_1490);
nand U4417 (N_4417,In_2374,In_2437);
xor U4418 (N_4418,In_680,In_2417);
nor U4419 (N_4419,In_804,In_2121);
or U4420 (N_4420,In_2002,In_1483);
and U4421 (N_4421,In_1044,In_144);
nand U4422 (N_4422,In_340,In_2873);
xnor U4423 (N_4423,In_1964,In_633);
nor U4424 (N_4424,In_2792,In_396);
nand U4425 (N_4425,In_265,In_975);
or U4426 (N_4426,In_2723,In_572);
nor U4427 (N_4427,In_767,In_2655);
nand U4428 (N_4428,In_942,In_621);
or U4429 (N_4429,In_725,In_544);
nor U4430 (N_4430,In_1823,In_88);
or U4431 (N_4431,In_1184,In_1471);
or U4432 (N_4432,In_736,In_1877);
nand U4433 (N_4433,In_2930,In_837);
nor U4434 (N_4434,In_1091,In_1394);
nor U4435 (N_4435,In_1614,In_1988);
and U4436 (N_4436,In_1411,In_1519);
or U4437 (N_4437,In_2103,In_2930);
xnor U4438 (N_4438,In_895,In_1126);
and U4439 (N_4439,In_784,In_2720);
or U4440 (N_4440,In_1669,In_7);
or U4441 (N_4441,In_1117,In_2022);
nor U4442 (N_4442,In_2812,In_969);
nand U4443 (N_4443,In_1939,In_1415);
nand U4444 (N_4444,In_424,In_2551);
or U4445 (N_4445,In_410,In_917);
nor U4446 (N_4446,In_2725,In_1700);
nand U4447 (N_4447,In_2627,In_2880);
nor U4448 (N_4448,In_2964,In_51);
or U4449 (N_4449,In_2542,In_849);
or U4450 (N_4450,In_119,In_1732);
xnor U4451 (N_4451,In_1447,In_1922);
nand U4452 (N_4452,In_1124,In_275);
nand U4453 (N_4453,In_1314,In_434);
or U4454 (N_4454,In_1345,In_1742);
or U4455 (N_4455,In_1704,In_1438);
and U4456 (N_4456,In_2938,In_2066);
nand U4457 (N_4457,In_1842,In_430);
nor U4458 (N_4458,In_2403,In_35);
or U4459 (N_4459,In_1289,In_507);
xnor U4460 (N_4460,In_227,In_1321);
nor U4461 (N_4461,In_1302,In_2021);
xor U4462 (N_4462,In_229,In_1002);
and U4463 (N_4463,In_539,In_2328);
and U4464 (N_4464,In_2373,In_487);
or U4465 (N_4465,In_2248,In_2119);
or U4466 (N_4466,In_489,In_1812);
nand U4467 (N_4467,In_2993,In_454);
or U4468 (N_4468,In_2502,In_1713);
or U4469 (N_4469,In_2313,In_1657);
nor U4470 (N_4470,In_2537,In_1324);
and U4471 (N_4471,In_1857,In_875);
and U4472 (N_4472,In_2717,In_2633);
or U4473 (N_4473,In_203,In_1716);
and U4474 (N_4474,In_2681,In_977);
nand U4475 (N_4475,In_2446,In_78);
or U4476 (N_4476,In_2794,In_2812);
and U4477 (N_4477,In_1511,In_179);
nand U4478 (N_4478,In_2787,In_434);
or U4479 (N_4479,In_17,In_2042);
and U4480 (N_4480,In_1658,In_707);
or U4481 (N_4481,In_2129,In_2048);
nand U4482 (N_4482,In_882,In_1886);
nand U4483 (N_4483,In_780,In_1962);
and U4484 (N_4484,In_2976,In_1019);
nand U4485 (N_4485,In_1681,In_518);
nor U4486 (N_4486,In_140,In_771);
or U4487 (N_4487,In_2699,In_1063);
and U4488 (N_4488,In_709,In_2636);
nor U4489 (N_4489,In_159,In_2788);
nor U4490 (N_4490,In_317,In_1636);
nand U4491 (N_4491,In_571,In_2323);
nand U4492 (N_4492,In_1785,In_132);
nand U4493 (N_4493,In_878,In_1706);
xor U4494 (N_4494,In_1102,In_1071);
xor U4495 (N_4495,In_1391,In_2621);
nand U4496 (N_4496,In_2572,In_184);
and U4497 (N_4497,In_1470,In_2378);
nor U4498 (N_4498,In_1283,In_2323);
nor U4499 (N_4499,In_143,In_606);
xnor U4500 (N_4500,In_245,In_2105);
nor U4501 (N_4501,In_64,In_1556);
or U4502 (N_4502,In_2541,In_2515);
xnor U4503 (N_4503,In_558,In_537);
nor U4504 (N_4504,In_2049,In_761);
or U4505 (N_4505,In_811,In_2379);
nor U4506 (N_4506,In_206,In_2312);
and U4507 (N_4507,In_2943,In_469);
or U4508 (N_4508,In_2343,In_1707);
nor U4509 (N_4509,In_2812,In_2717);
and U4510 (N_4510,In_1675,In_1579);
and U4511 (N_4511,In_1498,In_375);
or U4512 (N_4512,In_255,In_2514);
nand U4513 (N_4513,In_1149,In_1443);
and U4514 (N_4514,In_485,In_2085);
or U4515 (N_4515,In_1440,In_1429);
and U4516 (N_4516,In_2844,In_1094);
and U4517 (N_4517,In_1998,In_1110);
nor U4518 (N_4518,In_613,In_1635);
nand U4519 (N_4519,In_1398,In_2036);
nor U4520 (N_4520,In_2017,In_844);
nor U4521 (N_4521,In_1581,In_2619);
and U4522 (N_4522,In_2486,In_118);
xor U4523 (N_4523,In_1698,In_2087);
and U4524 (N_4524,In_706,In_1830);
nor U4525 (N_4525,In_2018,In_1522);
and U4526 (N_4526,In_1232,In_1206);
and U4527 (N_4527,In_1182,In_829);
and U4528 (N_4528,In_2759,In_1515);
and U4529 (N_4529,In_2642,In_2390);
and U4530 (N_4530,In_1277,In_595);
and U4531 (N_4531,In_2538,In_2643);
nor U4532 (N_4532,In_1158,In_504);
xor U4533 (N_4533,In_2917,In_1924);
and U4534 (N_4534,In_223,In_423);
nand U4535 (N_4535,In_1915,In_176);
nand U4536 (N_4536,In_705,In_1028);
or U4537 (N_4537,In_208,In_2872);
and U4538 (N_4538,In_614,In_2688);
or U4539 (N_4539,In_1365,In_566);
or U4540 (N_4540,In_2296,In_2939);
or U4541 (N_4541,In_1327,In_485);
or U4542 (N_4542,In_1423,In_936);
and U4543 (N_4543,In_466,In_2205);
and U4544 (N_4544,In_352,In_451);
xnor U4545 (N_4545,In_1341,In_826);
nor U4546 (N_4546,In_813,In_734);
nand U4547 (N_4547,In_2349,In_2070);
or U4548 (N_4548,In_2800,In_1321);
or U4549 (N_4549,In_104,In_2649);
and U4550 (N_4550,In_1878,In_1286);
or U4551 (N_4551,In_1139,In_819);
and U4552 (N_4552,In_2211,In_2277);
nand U4553 (N_4553,In_723,In_1457);
nand U4554 (N_4554,In_257,In_1620);
or U4555 (N_4555,In_433,In_2490);
or U4556 (N_4556,In_2876,In_52);
nor U4557 (N_4557,In_880,In_2124);
nor U4558 (N_4558,In_2663,In_2773);
and U4559 (N_4559,In_1403,In_1902);
or U4560 (N_4560,In_1384,In_693);
nand U4561 (N_4561,In_909,In_450);
and U4562 (N_4562,In_2588,In_1441);
xor U4563 (N_4563,In_259,In_1795);
nor U4564 (N_4564,In_2865,In_2165);
nand U4565 (N_4565,In_355,In_491);
or U4566 (N_4566,In_1162,In_161);
nand U4567 (N_4567,In_2642,In_690);
or U4568 (N_4568,In_2677,In_2611);
nand U4569 (N_4569,In_359,In_2426);
nor U4570 (N_4570,In_1955,In_740);
xnor U4571 (N_4571,In_2240,In_2737);
nand U4572 (N_4572,In_598,In_2903);
nor U4573 (N_4573,In_2019,In_948);
or U4574 (N_4574,In_1593,In_1769);
and U4575 (N_4575,In_2672,In_2357);
or U4576 (N_4576,In_913,In_807);
or U4577 (N_4577,In_2124,In_2476);
or U4578 (N_4578,In_266,In_835);
nor U4579 (N_4579,In_960,In_947);
or U4580 (N_4580,In_2190,In_1670);
and U4581 (N_4581,In_1352,In_2606);
nor U4582 (N_4582,In_1539,In_759);
xnor U4583 (N_4583,In_1030,In_972);
nand U4584 (N_4584,In_622,In_102);
nand U4585 (N_4585,In_1095,In_1022);
and U4586 (N_4586,In_2847,In_2161);
or U4587 (N_4587,In_2190,In_2589);
or U4588 (N_4588,In_2100,In_2852);
nor U4589 (N_4589,In_3,In_1386);
or U4590 (N_4590,In_1837,In_1076);
xor U4591 (N_4591,In_515,In_819);
nand U4592 (N_4592,In_2545,In_2717);
and U4593 (N_4593,In_698,In_1092);
nand U4594 (N_4594,In_616,In_1270);
or U4595 (N_4595,In_2256,In_2146);
nand U4596 (N_4596,In_1426,In_518);
or U4597 (N_4597,In_703,In_769);
nor U4598 (N_4598,In_26,In_100);
or U4599 (N_4599,In_780,In_1504);
or U4600 (N_4600,In_215,In_2686);
and U4601 (N_4601,In_1066,In_2422);
and U4602 (N_4602,In_888,In_1073);
and U4603 (N_4603,In_2617,In_2170);
nand U4604 (N_4604,In_2261,In_2908);
nor U4605 (N_4605,In_2748,In_1317);
nand U4606 (N_4606,In_1742,In_2887);
nand U4607 (N_4607,In_888,In_2862);
nor U4608 (N_4608,In_2050,In_549);
nand U4609 (N_4609,In_2739,In_1681);
nand U4610 (N_4610,In_2041,In_2557);
or U4611 (N_4611,In_0,In_17);
nor U4612 (N_4612,In_1937,In_94);
nor U4613 (N_4613,In_2536,In_1802);
nor U4614 (N_4614,In_678,In_851);
and U4615 (N_4615,In_805,In_1529);
nand U4616 (N_4616,In_2621,In_1280);
nand U4617 (N_4617,In_1303,In_2699);
xnor U4618 (N_4618,In_207,In_2943);
and U4619 (N_4619,In_2738,In_1399);
xnor U4620 (N_4620,In_890,In_2625);
and U4621 (N_4621,In_943,In_537);
xor U4622 (N_4622,In_2314,In_1694);
nor U4623 (N_4623,In_2080,In_2695);
nor U4624 (N_4624,In_117,In_2733);
nor U4625 (N_4625,In_2577,In_1598);
or U4626 (N_4626,In_1270,In_1983);
nor U4627 (N_4627,In_534,In_2291);
and U4628 (N_4628,In_17,In_2853);
and U4629 (N_4629,In_1564,In_276);
or U4630 (N_4630,In_275,In_2197);
or U4631 (N_4631,In_633,In_1421);
xor U4632 (N_4632,In_2709,In_2588);
and U4633 (N_4633,In_926,In_43);
or U4634 (N_4634,In_2242,In_707);
nor U4635 (N_4635,In_532,In_2082);
nor U4636 (N_4636,In_2677,In_2380);
nand U4637 (N_4637,In_2978,In_1606);
nor U4638 (N_4638,In_83,In_239);
nand U4639 (N_4639,In_1594,In_589);
nand U4640 (N_4640,In_1383,In_137);
or U4641 (N_4641,In_2525,In_659);
or U4642 (N_4642,In_2080,In_1321);
xnor U4643 (N_4643,In_583,In_2586);
nand U4644 (N_4644,In_2840,In_1848);
and U4645 (N_4645,In_605,In_1476);
and U4646 (N_4646,In_1991,In_170);
or U4647 (N_4647,In_1878,In_2403);
nor U4648 (N_4648,In_726,In_1340);
nand U4649 (N_4649,In_431,In_2839);
and U4650 (N_4650,In_2546,In_1022);
nor U4651 (N_4651,In_1623,In_553);
and U4652 (N_4652,In_591,In_1420);
and U4653 (N_4653,In_2145,In_959);
nor U4654 (N_4654,In_441,In_272);
nor U4655 (N_4655,In_2957,In_2990);
and U4656 (N_4656,In_800,In_2890);
and U4657 (N_4657,In_1332,In_1990);
nor U4658 (N_4658,In_1589,In_1521);
and U4659 (N_4659,In_875,In_159);
and U4660 (N_4660,In_2747,In_2563);
and U4661 (N_4661,In_1108,In_686);
and U4662 (N_4662,In_543,In_1256);
nand U4663 (N_4663,In_2621,In_2866);
or U4664 (N_4664,In_2552,In_2704);
or U4665 (N_4665,In_138,In_695);
or U4666 (N_4666,In_1904,In_1056);
and U4667 (N_4667,In_16,In_161);
and U4668 (N_4668,In_2007,In_179);
or U4669 (N_4669,In_1732,In_1960);
xor U4670 (N_4670,In_2904,In_1855);
nand U4671 (N_4671,In_1042,In_102);
nand U4672 (N_4672,In_2657,In_1150);
xor U4673 (N_4673,In_2452,In_1174);
nor U4674 (N_4674,In_2391,In_684);
nand U4675 (N_4675,In_552,In_2918);
and U4676 (N_4676,In_1373,In_2320);
nand U4677 (N_4677,In_1820,In_2325);
and U4678 (N_4678,In_247,In_481);
and U4679 (N_4679,In_1562,In_2285);
nor U4680 (N_4680,In_1907,In_95);
or U4681 (N_4681,In_2827,In_1768);
or U4682 (N_4682,In_846,In_1981);
nor U4683 (N_4683,In_2278,In_2875);
and U4684 (N_4684,In_311,In_2966);
xnor U4685 (N_4685,In_1684,In_1948);
nand U4686 (N_4686,In_2680,In_1424);
xor U4687 (N_4687,In_805,In_2296);
nor U4688 (N_4688,In_1463,In_1255);
nor U4689 (N_4689,In_1967,In_251);
or U4690 (N_4690,In_2131,In_2281);
or U4691 (N_4691,In_2367,In_2263);
nand U4692 (N_4692,In_774,In_2481);
nand U4693 (N_4693,In_2577,In_968);
and U4694 (N_4694,In_548,In_2648);
or U4695 (N_4695,In_1071,In_2435);
nand U4696 (N_4696,In_1275,In_866);
nand U4697 (N_4697,In_2966,In_2918);
nand U4698 (N_4698,In_1387,In_1580);
nor U4699 (N_4699,In_1092,In_2186);
nor U4700 (N_4700,In_1224,In_1792);
and U4701 (N_4701,In_650,In_1054);
and U4702 (N_4702,In_2162,In_2090);
nor U4703 (N_4703,In_1309,In_2404);
nor U4704 (N_4704,In_2952,In_2523);
xor U4705 (N_4705,In_202,In_2577);
and U4706 (N_4706,In_225,In_423);
and U4707 (N_4707,In_2780,In_502);
nor U4708 (N_4708,In_78,In_214);
and U4709 (N_4709,In_1903,In_203);
or U4710 (N_4710,In_86,In_2648);
xnor U4711 (N_4711,In_2408,In_114);
nor U4712 (N_4712,In_539,In_2445);
nor U4713 (N_4713,In_2558,In_739);
nor U4714 (N_4714,In_2161,In_1993);
nand U4715 (N_4715,In_2223,In_1327);
nor U4716 (N_4716,In_214,In_1933);
and U4717 (N_4717,In_1346,In_42);
nor U4718 (N_4718,In_290,In_758);
or U4719 (N_4719,In_733,In_1448);
nand U4720 (N_4720,In_1295,In_2334);
nand U4721 (N_4721,In_1857,In_1915);
nor U4722 (N_4722,In_105,In_2803);
nor U4723 (N_4723,In_1471,In_2222);
nor U4724 (N_4724,In_2879,In_167);
or U4725 (N_4725,In_576,In_1627);
nand U4726 (N_4726,In_1628,In_2520);
or U4727 (N_4727,In_898,In_2512);
nor U4728 (N_4728,In_1042,In_2423);
and U4729 (N_4729,In_2269,In_2125);
or U4730 (N_4730,In_988,In_1357);
nor U4731 (N_4731,In_2145,In_311);
nor U4732 (N_4732,In_2239,In_2077);
or U4733 (N_4733,In_126,In_320);
or U4734 (N_4734,In_524,In_558);
or U4735 (N_4735,In_2485,In_218);
nor U4736 (N_4736,In_2775,In_2332);
xor U4737 (N_4737,In_811,In_576);
nand U4738 (N_4738,In_930,In_2560);
xor U4739 (N_4739,In_952,In_1629);
nor U4740 (N_4740,In_408,In_1729);
and U4741 (N_4741,In_495,In_269);
nand U4742 (N_4742,In_2614,In_1162);
or U4743 (N_4743,In_179,In_2550);
and U4744 (N_4744,In_1583,In_2316);
and U4745 (N_4745,In_232,In_346);
and U4746 (N_4746,In_2711,In_467);
nor U4747 (N_4747,In_464,In_3);
nand U4748 (N_4748,In_869,In_2433);
and U4749 (N_4749,In_1012,In_2842);
xor U4750 (N_4750,In_2704,In_435);
nand U4751 (N_4751,In_1261,In_2175);
nor U4752 (N_4752,In_1848,In_574);
or U4753 (N_4753,In_2514,In_2614);
nor U4754 (N_4754,In_1344,In_2485);
nand U4755 (N_4755,In_152,In_741);
and U4756 (N_4756,In_2459,In_2421);
nand U4757 (N_4757,In_2415,In_1177);
xor U4758 (N_4758,In_2208,In_560);
and U4759 (N_4759,In_2021,In_165);
or U4760 (N_4760,In_1702,In_369);
xnor U4761 (N_4761,In_2249,In_2165);
nor U4762 (N_4762,In_1188,In_1286);
and U4763 (N_4763,In_609,In_611);
xor U4764 (N_4764,In_75,In_553);
and U4765 (N_4765,In_2613,In_487);
and U4766 (N_4766,In_2689,In_17);
nor U4767 (N_4767,In_2677,In_1516);
nand U4768 (N_4768,In_1970,In_791);
and U4769 (N_4769,In_1361,In_778);
or U4770 (N_4770,In_2043,In_1630);
nand U4771 (N_4771,In_892,In_2654);
nand U4772 (N_4772,In_514,In_1397);
or U4773 (N_4773,In_197,In_675);
nor U4774 (N_4774,In_1963,In_2724);
and U4775 (N_4775,In_66,In_1076);
nor U4776 (N_4776,In_1877,In_2895);
nor U4777 (N_4777,In_18,In_605);
and U4778 (N_4778,In_1307,In_2759);
nand U4779 (N_4779,In_433,In_1412);
xor U4780 (N_4780,In_677,In_962);
nor U4781 (N_4781,In_2159,In_1575);
and U4782 (N_4782,In_1463,In_1596);
nor U4783 (N_4783,In_191,In_1022);
xnor U4784 (N_4784,In_2723,In_2372);
or U4785 (N_4785,In_1687,In_638);
xnor U4786 (N_4786,In_1869,In_2789);
xnor U4787 (N_4787,In_1602,In_2396);
nor U4788 (N_4788,In_1125,In_1663);
nor U4789 (N_4789,In_2366,In_1286);
or U4790 (N_4790,In_1786,In_1954);
nand U4791 (N_4791,In_2396,In_2962);
and U4792 (N_4792,In_1662,In_1514);
nand U4793 (N_4793,In_1574,In_1792);
and U4794 (N_4794,In_1040,In_2208);
or U4795 (N_4795,In_2971,In_2610);
nor U4796 (N_4796,In_2135,In_364);
nor U4797 (N_4797,In_1800,In_1277);
and U4798 (N_4798,In_366,In_1513);
and U4799 (N_4799,In_2082,In_864);
nand U4800 (N_4800,In_1137,In_1767);
and U4801 (N_4801,In_1441,In_1785);
nand U4802 (N_4802,In_1587,In_2015);
or U4803 (N_4803,In_1919,In_826);
nor U4804 (N_4804,In_2907,In_2252);
nand U4805 (N_4805,In_330,In_811);
xor U4806 (N_4806,In_193,In_2988);
nand U4807 (N_4807,In_1038,In_54);
nor U4808 (N_4808,In_2778,In_2418);
and U4809 (N_4809,In_2004,In_602);
or U4810 (N_4810,In_945,In_2208);
nand U4811 (N_4811,In_902,In_1516);
nand U4812 (N_4812,In_1010,In_824);
and U4813 (N_4813,In_1146,In_1939);
nand U4814 (N_4814,In_1538,In_522);
nand U4815 (N_4815,In_507,In_159);
or U4816 (N_4816,In_1074,In_613);
and U4817 (N_4817,In_316,In_2915);
and U4818 (N_4818,In_2540,In_1676);
nand U4819 (N_4819,In_2663,In_658);
xnor U4820 (N_4820,In_487,In_2229);
and U4821 (N_4821,In_622,In_581);
or U4822 (N_4822,In_2560,In_2838);
nor U4823 (N_4823,In_1232,In_2279);
and U4824 (N_4824,In_1075,In_2690);
nor U4825 (N_4825,In_1300,In_928);
and U4826 (N_4826,In_2171,In_1046);
and U4827 (N_4827,In_50,In_1565);
nor U4828 (N_4828,In_2160,In_1097);
and U4829 (N_4829,In_1233,In_2472);
and U4830 (N_4830,In_933,In_2083);
nand U4831 (N_4831,In_365,In_321);
xor U4832 (N_4832,In_2224,In_1445);
nand U4833 (N_4833,In_2878,In_2711);
nor U4834 (N_4834,In_2626,In_681);
nand U4835 (N_4835,In_2321,In_402);
xor U4836 (N_4836,In_2017,In_1361);
or U4837 (N_4837,In_2842,In_2461);
nor U4838 (N_4838,In_2345,In_846);
xor U4839 (N_4839,In_1911,In_1053);
or U4840 (N_4840,In_344,In_1840);
and U4841 (N_4841,In_1703,In_1928);
or U4842 (N_4842,In_503,In_248);
nor U4843 (N_4843,In_2423,In_268);
or U4844 (N_4844,In_1132,In_1866);
nor U4845 (N_4845,In_2475,In_2820);
nor U4846 (N_4846,In_2068,In_678);
or U4847 (N_4847,In_750,In_331);
and U4848 (N_4848,In_2549,In_1507);
and U4849 (N_4849,In_1219,In_1298);
or U4850 (N_4850,In_2832,In_2668);
and U4851 (N_4851,In_215,In_1183);
nor U4852 (N_4852,In_1585,In_1440);
or U4853 (N_4853,In_2539,In_270);
and U4854 (N_4854,In_1448,In_2079);
nand U4855 (N_4855,In_2105,In_278);
and U4856 (N_4856,In_831,In_1439);
or U4857 (N_4857,In_484,In_2773);
or U4858 (N_4858,In_1991,In_2258);
nand U4859 (N_4859,In_1121,In_2643);
nand U4860 (N_4860,In_1947,In_602);
nor U4861 (N_4861,In_1959,In_271);
or U4862 (N_4862,In_1291,In_1222);
or U4863 (N_4863,In_1097,In_1498);
nor U4864 (N_4864,In_1459,In_2479);
or U4865 (N_4865,In_904,In_101);
or U4866 (N_4866,In_2146,In_2796);
and U4867 (N_4867,In_2161,In_1035);
and U4868 (N_4868,In_1760,In_2724);
and U4869 (N_4869,In_412,In_1915);
and U4870 (N_4870,In_2758,In_2115);
nand U4871 (N_4871,In_2013,In_1720);
nand U4872 (N_4872,In_2765,In_506);
xor U4873 (N_4873,In_2281,In_1917);
nand U4874 (N_4874,In_1364,In_2122);
and U4875 (N_4875,In_2143,In_256);
or U4876 (N_4876,In_1849,In_1824);
and U4877 (N_4877,In_540,In_544);
or U4878 (N_4878,In_2014,In_268);
xor U4879 (N_4879,In_1791,In_733);
nor U4880 (N_4880,In_890,In_1583);
nor U4881 (N_4881,In_1857,In_1156);
nor U4882 (N_4882,In_122,In_642);
nor U4883 (N_4883,In_2600,In_1771);
and U4884 (N_4884,In_1826,In_2151);
and U4885 (N_4885,In_2432,In_25);
xnor U4886 (N_4886,In_2845,In_2262);
nor U4887 (N_4887,In_168,In_2699);
and U4888 (N_4888,In_2007,In_687);
nand U4889 (N_4889,In_747,In_2338);
or U4890 (N_4890,In_2014,In_2355);
nand U4891 (N_4891,In_2491,In_2346);
nor U4892 (N_4892,In_1280,In_2668);
nor U4893 (N_4893,In_1198,In_1877);
nor U4894 (N_4894,In_2667,In_2815);
nor U4895 (N_4895,In_1740,In_408);
and U4896 (N_4896,In_452,In_2139);
and U4897 (N_4897,In_359,In_2198);
or U4898 (N_4898,In_813,In_2607);
or U4899 (N_4899,In_1602,In_1553);
and U4900 (N_4900,In_1703,In_2438);
nand U4901 (N_4901,In_1338,In_2389);
or U4902 (N_4902,In_1268,In_2160);
nor U4903 (N_4903,In_1813,In_1585);
nand U4904 (N_4904,In_2564,In_1018);
and U4905 (N_4905,In_908,In_2711);
nor U4906 (N_4906,In_1002,In_355);
nor U4907 (N_4907,In_935,In_2527);
and U4908 (N_4908,In_338,In_394);
and U4909 (N_4909,In_2096,In_1580);
or U4910 (N_4910,In_422,In_2139);
and U4911 (N_4911,In_2935,In_645);
nand U4912 (N_4912,In_1219,In_1538);
and U4913 (N_4913,In_459,In_2134);
or U4914 (N_4914,In_2561,In_2652);
or U4915 (N_4915,In_2849,In_1033);
and U4916 (N_4916,In_2669,In_907);
xnor U4917 (N_4917,In_1191,In_409);
or U4918 (N_4918,In_2131,In_2947);
and U4919 (N_4919,In_2140,In_714);
xnor U4920 (N_4920,In_792,In_1628);
and U4921 (N_4921,In_1192,In_1775);
nor U4922 (N_4922,In_1967,In_127);
nand U4923 (N_4923,In_1064,In_2122);
nor U4924 (N_4924,In_2923,In_553);
and U4925 (N_4925,In_1172,In_2766);
or U4926 (N_4926,In_1429,In_931);
and U4927 (N_4927,In_508,In_1324);
nand U4928 (N_4928,In_2705,In_214);
nor U4929 (N_4929,In_883,In_2041);
and U4930 (N_4930,In_2681,In_2759);
or U4931 (N_4931,In_320,In_1313);
nand U4932 (N_4932,In_2465,In_72);
and U4933 (N_4933,In_1127,In_1109);
xor U4934 (N_4934,In_795,In_858);
nand U4935 (N_4935,In_75,In_2060);
and U4936 (N_4936,In_996,In_2836);
or U4937 (N_4937,In_1770,In_1610);
nor U4938 (N_4938,In_2740,In_1776);
xor U4939 (N_4939,In_1306,In_2530);
and U4940 (N_4940,In_206,In_377);
and U4941 (N_4941,In_201,In_815);
nor U4942 (N_4942,In_1533,In_1036);
xor U4943 (N_4943,In_1908,In_898);
xor U4944 (N_4944,In_1480,In_202);
xor U4945 (N_4945,In_1956,In_199);
nand U4946 (N_4946,In_2983,In_2171);
and U4947 (N_4947,In_1594,In_2743);
and U4948 (N_4948,In_845,In_882);
nor U4949 (N_4949,In_2678,In_863);
and U4950 (N_4950,In_2615,In_126);
or U4951 (N_4951,In_581,In_382);
nand U4952 (N_4952,In_298,In_2713);
nor U4953 (N_4953,In_1522,In_2960);
and U4954 (N_4954,In_62,In_2331);
xnor U4955 (N_4955,In_758,In_1295);
nand U4956 (N_4956,In_1385,In_867);
or U4957 (N_4957,In_426,In_714);
or U4958 (N_4958,In_267,In_150);
nor U4959 (N_4959,In_238,In_2835);
nand U4960 (N_4960,In_1201,In_1540);
nor U4961 (N_4961,In_1038,In_1327);
nand U4962 (N_4962,In_301,In_1397);
and U4963 (N_4963,In_2682,In_1385);
and U4964 (N_4964,In_1772,In_1759);
xor U4965 (N_4965,In_1474,In_2886);
and U4966 (N_4966,In_1213,In_538);
nor U4967 (N_4967,In_820,In_2970);
or U4968 (N_4968,In_2906,In_1999);
and U4969 (N_4969,In_2813,In_54);
nand U4970 (N_4970,In_2052,In_2672);
nor U4971 (N_4971,In_2492,In_120);
and U4972 (N_4972,In_174,In_257);
nand U4973 (N_4973,In_1738,In_1951);
nor U4974 (N_4974,In_1317,In_464);
and U4975 (N_4975,In_1148,In_1708);
xor U4976 (N_4976,In_1066,In_2611);
nand U4977 (N_4977,In_132,In_2038);
or U4978 (N_4978,In_2480,In_431);
nand U4979 (N_4979,In_92,In_866);
nor U4980 (N_4980,In_2191,In_902);
and U4981 (N_4981,In_546,In_1393);
and U4982 (N_4982,In_2632,In_1784);
and U4983 (N_4983,In_2094,In_2664);
nand U4984 (N_4984,In_1234,In_1815);
and U4985 (N_4985,In_721,In_2116);
and U4986 (N_4986,In_2056,In_644);
or U4987 (N_4987,In_1181,In_728);
nor U4988 (N_4988,In_2956,In_1724);
nor U4989 (N_4989,In_1787,In_2959);
xor U4990 (N_4990,In_1686,In_2006);
and U4991 (N_4991,In_1263,In_251);
xnor U4992 (N_4992,In_2161,In_1864);
and U4993 (N_4993,In_1871,In_412);
nand U4994 (N_4994,In_2994,In_1763);
nand U4995 (N_4995,In_2046,In_2602);
or U4996 (N_4996,In_755,In_2578);
or U4997 (N_4997,In_2941,In_2318);
nand U4998 (N_4998,In_1334,In_56);
nor U4999 (N_4999,In_452,In_2278);
nor U5000 (N_5000,N_4932,N_1368);
nand U5001 (N_5001,N_3899,N_930);
nor U5002 (N_5002,N_3359,N_3988);
nor U5003 (N_5003,N_3986,N_1390);
nand U5004 (N_5004,N_4058,N_4758);
and U5005 (N_5005,N_1352,N_394);
nor U5006 (N_5006,N_4878,N_4757);
nand U5007 (N_5007,N_4000,N_1687);
nand U5008 (N_5008,N_246,N_2139);
nand U5009 (N_5009,N_3865,N_2463);
xnor U5010 (N_5010,N_4671,N_2330);
nand U5011 (N_5011,N_1730,N_2771);
nor U5012 (N_5012,N_1196,N_4836);
xnor U5013 (N_5013,N_1870,N_3692);
nand U5014 (N_5014,N_964,N_2650);
nand U5015 (N_5015,N_4755,N_4214);
and U5016 (N_5016,N_79,N_265);
nor U5017 (N_5017,N_1770,N_1978);
xnor U5018 (N_5018,N_2690,N_445);
and U5019 (N_5019,N_1972,N_3488);
or U5020 (N_5020,N_4578,N_4929);
nor U5021 (N_5021,N_4653,N_645);
nor U5022 (N_5022,N_3546,N_832);
and U5023 (N_5023,N_738,N_3177);
nand U5024 (N_5024,N_739,N_1737);
xnor U5025 (N_5025,N_617,N_4864);
nand U5026 (N_5026,N_3111,N_4262);
nor U5027 (N_5027,N_1965,N_1066);
or U5028 (N_5028,N_4496,N_227);
nand U5029 (N_5029,N_2806,N_4588);
nor U5030 (N_5030,N_3621,N_2216);
xnor U5031 (N_5031,N_2737,N_2765);
or U5032 (N_5032,N_1320,N_81);
or U5033 (N_5033,N_2816,N_4279);
nand U5034 (N_5034,N_4123,N_3374);
nand U5035 (N_5035,N_1,N_328);
and U5036 (N_5036,N_101,N_3946);
xnor U5037 (N_5037,N_268,N_1051);
or U5038 (N_5038,N_1553,N_4253);
nor U5039 (N_5039,N_4295,N_1597);
and U5040 (N_5040,N_973,N_1173);
or U5041 (N_5041,N_1588,N_2408);
nor U5042 (N_5042,N_2697,N_4226);
nand U5043 (N_5043,N_3218,N_2836);
or U5044 (N_5044,N_2554,N_562);
or U5045 (N_5045,N_2295,N_2963);
or U5046 (N_5046,N_1925,N_821);
nor U5047 (N_5047,N_3388,N_1873);
nor U5048 (N_5048,N_1487,N_4767);
or U5049 (N_5049,N_3225,N_2629);
nor U5050 (N_5050,N_4851,N_377);
nand U5051 (N_5051,N_1935,N_4773);
and U5052 (N_5052,N_3530,N_1828);
nand U5053 (N_5053,N_1706,N_747);
and U5054 (N_5054,N_4739,N_3879);
nor U5055 (N_5055,N_321,N_446);
or U5056 (N_5056,N_4259,N_1260);
nor U5057 (N_5057,N_3471,N_197);
nor U5058 (N_5058,N_2222,N_4078);
nor U5059 (N_5059,N_1938,N_3615);
or U5060 (N_5060,N_3492,N_274);
and U5061 (N_5061,N_4893,N_184);
nor U5062 (N_5062,N_3289,N_3393);
nor U5063 (N_5063,N_4621,N_2179);
and U5064 (N_5064,N_857,N_983);
xor U5065 (N_5065,N_4114,N_1946);
nor U5066 (N_5066,N_2522,N_4868);
nand U5067 (N_5067,N_3964,N_2521);
nand U5068 (N_5068,N_1958,N_2882);
xnor U5069 (N_5069,N_2280,N_833);
and U5070 (N_5070,N_4187,N_4507);
and U5071 (N_5071,N_4592,N_914);
or U5072 (N_5072,N_4941,N_4813);
nand U5073 (N_5073,N_3222,N_41);
nand U5074 (N_5074,N_3079,N_1874);
xnor U5075 (N_5075,N_4514,N_228);
xor U5076 (N_5076,N_1461,N_968);
nand U5077 (N_5077,N_178,N_3073);
xor U5078 (N_5078,N_3,N_143);
and U5079 (N_5079,N_135,N_2721);
nand U5080 (N_5080,N_3658,N_421);
or U5081 (N_5081,N_1495,N_782);
nor U5082 (N_5082,N_1323,N_1435);
nor U5083 (N_5083,N_4989,N_2596);
nand U5084 (N_5084,N_3528,N_4701);
and U5085 (N_5085,N_3877,N_2504);
nand U5086 (N_5086,N_1454,N_493);
and U5087 (N_5087,N_3258,N_4736);
nor U5088 (N_5088,N_1559,N_3751);
nand U5089 (N_5089,N_4024,N_1085);
or U5090 (N_5090,N_3957,N_1816);
nand U5091 (N_5091,N_2687,N_4471);
and U5092 (N_5092,N_504,N_4321);
xnor U5093 (N_5093,N_1557,N_3547);
and U5094 (N_5094,N_820,N_1902);
xor U5095 (N_5095,N_4324,N_2660);
and U5096 (N_5096,N_2838,N_234);
nor U5097 (N_5097,N_1305,N_3826);
nand U5098 (N_5098,N_2525,N_3399);
or U5099 (N_5099,N_4013,N_3197);
nand U5100 (N_5100,N_2586,N_2112);
xor U5101 (N_5101,N_1418,N_2275);
nand U5102 (N_5102,N_1008,N_42);
nand U5103 (N_5103,N_4064,N_126);
or U5104 (N_5104,N_3053,N_1239);
xnor U5105 (N_5105,N_3854,N_4768);
nor U5106 (N_5106,N_839,N_2964);
nand U5107 (N_5107,N_1378,N_2953);
nor U5108 (N_5108,N_4745,N_2253);
and U5109 (N_5109,N_3541,N_3990);
and U5110 (N_5110,N_2855,N_3713);
or U5111 (N_5111,N_4860,N_1826);
or U5112 (N_5112,N_429,N_2908);
or U5113 (N_5113,N_4798,N_3945);
nor U5114 (N_5114,N_3228,N_2927);
xor U5115 (N_5115,N_3357,N_1625);
nand U5116 (N_5116,N_1739,N_1395);
xnor U5117 (N_5117,N_931,N_4030);
nor U5118 (N_5118,N_1824,N_4116);
nor U5119 (N_5119,N_3319,N_3277);
or U5120 (N_5120,N_4317,N_1459);
nor U5121 (N_5121,N_4695,N_1410);
and U5122 (N_5122,N_3119,N_2287);
and U5123 (N_5123,N_4314,N_4051);
or U5124 (N_5124,N_2160,N_2221);
xor U5125 (N_5125,N_975,N_4610);
nor U5126 (N_5126,N_1855,N_3639);
xnor U5127 (N_5127,N_4502,N_1000);
xnor U5128 (N_5128,N_1974,N_1227);
nor U5129 (N_5129,N_4707,N_4367);
nor U5130 (N_5130,N_3507,N_3013);
nand U5131 (N_5131,N_4923,N_1984);
or U5132 (N_5132,N_3041,N_354);
nor U5133 (N_5133,N_192,N_2546);
nand U5134 (N_5134,N_1614,N_253);
nand U5135 (N_5135,N_3366,N_2950);
nand U5136 (N_5136,N_2294,N_342);
nand U5137 (N_5137,N_2945,N_3993);
xnor U5138 (N_5138,N_2892,N_825);
or U5139 (N_5139,N_654,N_4270);
xor U5140 (N_5140,N_3424,N_4774);
nor U5141 (N_5141,N_2700,N_3750);
and U5142 (N_5142,N_1396,N_608);
nand U5143 (N_5143,N_4733,N_1391);
and U5144 (N_5144,N_530,N_3351);
nor U5145 (N_5145,N_27,N_392);
and U5146 (N_5146,N_2471,N_4043);
nand U5147 (N_5147,N_3102,N_2155);
xnor U5148 (N_5148,N_2211,N_1302);
nor U5149 (N_5149,N_1119,N_4600);
nand U5150 (N_5150,N_2503,N_3311);
or U5151 (N_5151,N_353,N_3634);
xnor U5152 (N_5152,N_1895,N_1463);
and U5153 (N_5153,N_2915,N_2020);
nand U5154 (N_5154,N_3076,N_1186);
nand U5155 (N_5155,N_4389,N_4935);
nor U5156 (N_5156,N_1638,N_4955);
or U5157 (N_5157,N_3014,N_695);
nor U5158 (N_5158,N_660,N_2844);
nand U5159 (N_5159,N_2207,N_4155);
nand U5160 (N_5160,N_4406,N_701);
nor U5161 (N_5161,N_4092,N_3917);
and U5162 (N_5162,N_4917,N_2972);
nand U5163 (N_5163,N_2192,N_1424);
xnor U5164 (N_5164,N_1922,N_3989);
nand U5165 (N_5165,N_1993,N_3731);
and U5166 (N_5166,N_3836,N_687);
and U5167 (N_5167,N_2724,N_4292);
nor U5168 (N_5168,N_1684,N_3601);
nand U5169 (N_5169,N_2616,N_4056);
and U5170 (N_5170,N_3510,N_3770);
nand U5171 (N_5171,N_2173,N_4005);
nor U5172 (N_5172,N_2223,N_218);
or U5173 (N_5173,N_865,N_1631);
or U5174 (N_5174,N_2602,N_1982);
nand U5175 (N_5175,N_4760,N_4053);
or U5176 (N_5176,N_1213,N_1483);
and U5177 (N_5177,N_4237,N_207);
or U5178 (N_5178,N_3938,N_1132);
xnor U5179 (N_5179,N_4085,N_3007);
nor U5180 (N_5180,N_2854,N_1866);
nor U5181 (N_5181,N_3443,N_162);
nand U5182 (N_5182,N_1711,N_2931);
and U5183 (N_5183,N_3320,N_2262);
nand U5184 (N_5184,N_2313,N_515);
nor U5185 (N_5185,N_1152,N_665);
or U5186 (N_5186,N_3650,N_1637);
or U5187 (N_5187,N_4103,N_3091);
nand U5188 (N_5188,N_760,N_1226);
nor U5189 (N_5189,N_4985,N_3331);
nand U5190 (N_5190,N_3147,N_2130);
and U5191 (N_5191,N_4029,N_3752);
and U5192 (N_5192,N_2068,N_72);
or U5193 (N_5193,N_2532,N_4119);
nor U5194 (N_5194,N_2792,N_160);
or U5195 (N_5195,N_4120,N_3392);
nor U5196 (N_5196,N_804,N_2191);
nand U5197 (N_5197,N_1298,N_575);
xor U5198 (N_5198,N_3195,N_3201);
nor U5199 (N_5199,N_479,N_1832);
or U5200 (N_5200,N_355,N_1791);
xnor U5201 (N_5201,N_4657,N_2888);
nor U5202 (N_5202,N_1210,N_1114);
xor U5203 (N_5203,N_4529,N_3644);
nor U5204 (N_5204,N_508,N_2877);
or U5205 (N_5205,N_1010,N_1412);
nand U5206 (N_5206,N_3573,N_3354);
nand U5207 (N_5207,N_849,N_1878);
and U5208 (N_5208,N_3684,N_3685);
nor U5209 (N_5209,N_4151,N_4345);
or U5210 (N_5210,N_3848,N_1886);
nand U5211 (N_5211,N_4892,N_4459);
nor U5212 (N_5212,N_4271,N_198);
and U5213 (N_5213,N_1350,N_777);
nand U5214 (N_5214,N_2449,N_781);
nor U5215 (N_5215,N_2392,N_991);
or U5216 (N_5216,N_4559,N_33);
and U5217 (N_5217,N_3061,N_1515);
nand U5218 (N_5218,N_1273,N_1995);
nor U5219 (N_5219,N_3813,N_1250);
or U5220 (N_5220,N_3950,N_2583);
xor U5221 (N_5221,N_4210,N_3120);
or U5222 (N_5222,N_2605,N_3696);
nor U5223 (N_5223,N_3974,N_3485);
and U5224 (N_5224,N_1147,N_2121);
nor U5225 (N_5225,N_1903,N_800);
nor U5226 (N_5226,N_3868,N_4705);
or U5227 (N_5227,N_2233,N_2367);
or U5228 (N_5228,N_3861,N_190);
or U5229 (N_5229,N_2328,N_3429);
nor U5230 (N_5230,N_4313,N_634);
nand U5231 (N_5231,N_2590,N_1278);
or U5232 (N_5232,N_3063,N_1564);
xnor U5233 (N_5233,N_113,N_620);
or U5234 (N_5234,N_3211,N_402);
or U5235 (N_5235,N_1952,N_3844);
nor U5236 (N_5236,N_1530,N_2540);
nor U5237 (N_5237,N_2579,N_55);
or U5238 (N_5238,N_4518,N_668);
nand U5239 (N_5239,N_2309,N_1635);
xnor U5240 (N_5240,N_1098,N_1802);
nand U5241 (N_5241,N_3155,N_1703);
xor U5242 (N_5242,N_2929,N_859);
or U5243 (N_5243,N_4238,N_2807);
nor U5244 (N_5244,N_1823,N_2990);
xnor U5245 (N_5245,N_2418,N_2597);
or U5246 (N_5246,N_4659,N_1441);
and U5247 (N_5247,N_548,N_1808);
or U5248 (N_5248,N_3935,N_329);
and U5249 (N_5249,N_2035,N_2960);
nand U5250 (N_5250,N_790,N_4797);
and U5251 (N_5251,N_1837,N_58);
or U5252 (N_5252,N_4280,N_2077);
nor U5253 (N_5253,N_4138,N_1231);
and U5254 (N_5254,N_4796,N_963);
nand U5255 (N_5255,N_2264,N_2243);
nor U5256 (N_5256,N_4627,N_2249);
and U5257 (N_5257,N_3720,N_288);
nand U5258 (N_5258,N_3379,N_212);
or U5259 (N_5259,N_2943,N_2870);
nor U5260 (N_5260,N_4023,N_3240);
nand U5261 (N_5261,N_908,N_3569);
nand U5262 (N_5262,N_270,N_1279);
nor U5263 (N_5263,N_626,N_1343);
nor U5264 (N_5264,N_524,N_3298);
or U5265 (N_5265,N_3845,N_2909);
nor U5266 (N_5266,N_2865,N_3828);
and U5267 (N_5267,N_1203,N_662);
nand U5268 (N_5268,N_2234,N_3166);
or U5269 (N_5269,N_3288,N_2875);
and U5270 (N_5270,N_4579,N_4719);
or U5271 (N_5271,N_2588,N_1095);
and U5272 (N_5272,N_1087,N_2305);
nand U5273 (N_5273,N_555,N_1924);
or U5274 (N_5274,N_4127,N_59);
nor U5275 (N_5275,N_3971,N_2251);
and U5276 (N_5276,N_2417,N_538);
nor U5277 (N_5277,N_3801,N_320);
and U5278 (N_5278,N_692,N_3800);
nand U5279 (N_5279,N_133,N_436);
or U5280 (N_5280,N_4354,N_4890);
and U5281 (N_5281,N_764,N_1516);
nor U5282 (N_5282,N_3436,N_1247);
and U5283 (N_5283,N_4034,N_3884);
or U5284 (N_5284,N_2144,N_1310);
nand U5285 (N_5285,N_1243,N_3985);
xor U5286 (N_5286,N_2566,N_1282);
and U5287 (N_5287,N_4953,N_393);
nand U5288 (N_5288,N_3815,N_2686);
nor U5289 (N_5289,N_2947,N_2889);
nand U5290 (N_5290,N_4224,N_439);
nor U5291 (N_5291,N_407,N_3416);
or U5292 (N_5292,N_1472,N_2147);
nor U5293 (N_5293,N_4776,N_3760);
or U5294 (N_5294,N_4623,N_4785);
nor U5295 (N_5295,N_3793,N_840);
xor U5296 (N_5296,N_2618,N_3239);
nor U5297 (N_5297,N_2767,N_3797);
xnor U5298 (N_5298,N_3653,N_1399);
and U5299 (N_5299,N_4910,N_3723);
nand U5300 (N_5300,N_2850,N_2493);
nor U5301 (N_5301,N_1723,N_1827);
nor U5302 (N_5302,N_1224,N_3663);
nor U5303 (N_5303,N_813,N_1176);
or U5304 (N_5304,N_4423,N_4699);
or U5305 (N_5305,N_4972,N_1766);
and U5306 (N_5306,N_2815,N_3018);
and U5307 (N_5307,N_1128,N_1208);
or U5308 (N_5308,N_2201,N_2928);
nand U5309 (N_5309,N_4337,N_4427);
and U5310 (N_5310,N_3338,N_664);
or U5311 (N_5311,N_3009,N_263);
and U5312 (N_5312,N_3033,N_3323);
xor U5313 (N_5313,N_3247,N_275);
or U5314 (N_5314,N_1541,N_2872);
and U5315 (N_5315,N_744,N_301);
nor U5316 (N_5316,N_1756,N_2980);
or U5317 (N_5317,N_433,N_4647);
nor U5318 (N_5318,N_4149,N_3386);
nand U5319 (N_5319,N_1835,N_2006);
nand U5320 (N_5320,N_1782,N_1550);
or U5321 (N_5321,N_1311,N_1618);
nor U5322 (N_5322,N_4981,N_3857);
or U5323 (N_5323,N_3817,N_1328);
xor U5324 (N_5324,N_4183,N_2527);
or U5325 (N_5325,N_3486,N_4914);
nand U5326 (N_5326,N_1380,N_1107);
or U5327 (N_5327,N_3806,N_3415);
nand U5328 (N_5328,N_171,N_4918);
nor U5329 (N_5329,N_629,N_3339);
nor U5330 (N_5330,N_3114,N_3852);
xor U5331 (N_5331,N_2483,N_724);
and U5332 (N_5332,N_336,N_2492);
or U5333 (N_5333,N_958,N_693);
or U5334 (N_5334,N_3505,N_2741);
nor U5335 (N_5335,N_2707,N_1376);
nor U5336 (N_5336,N_2636,N_1634);
nand U5337 (N_5337,N_2433,N_2303);
or U5338 (N_5338,N_3786,N_4749);
nor U5339 (N_5339,N_4865,N_2536);
nand U5340 (N_5340,N_3688,N_1434);
nor U5341 (N_5341,N_3671,N_3918);
or U5342 (N_5342,N_4930,N_2117);
and U5343 (N_5343,N_3635,N_3104);
xnor U5344 (N_5344,N_3315,N_2695);
nand U5345 (N_5345,N_2106,N_4572);
nor U5346 (N_5346,N_4885,N_3941);
nand U5347 (N_5347,N_837,N_1414);
or U5348 (N_5348,N_2907,N_1889);
nand U5349 (N_5349,N_2839,N_1382);
nor U5350 (N_5350,N_2027,N_82);
nor U5351 (N_5351,N_823,N_1928);
or U5352 (N_5352,N_1740,N_2712);
nand U5353 (N_5353,N_3862,N_3292);
nand U5354 (N_5354,N_4505,N_4526);
xor U5355 (N_5355,N_102,N_2852);
nor U5356 (N_5356,N_391,N_231);
nand U5357 (N_5357,N_2312,N_4152);
and U5358 (N_5358,N_1612,N_2282);
and U5359 (N_5359,N_3140,N_4576);
xnor U5360 (N_5360,N_1222,N_1182);
nand U5361 (N_5361,N_4681,N_2893);
nand U5362 (N_5362,N_1754,N_343);
or U5363 (N_5363,N_352,N_4702);
and U5364 (N_5364,N_667,N_4492);
and U5365 (N_5365,N_3340,N_381);
and U5366 (N_5366,N_1348,N_792);
or U5367 (N_5367,N_2977,N_405);
or U5368 (N_5368,N_3494,N_831);
nand U5369 (N_5369,N_3876,N_3252);
nand U5370 (N_5370,N_3972,N_1174);
nor U5371 (N_5371,N_732,N_2814);
and U5372 (N_5372,N_3039,N_211);
nand U5373 (N_5373,N_1170,N_960);
nand U5374 (N_5374,N_116,N_2246);
and U5375 (N_5375,N_1052,N_3164);
nor U5376 (N_5376,N_826,N_2250);
or U5377 (N_5377,N_1709,N_296);
nand U5378 (N_5378,N_3452,N_1292);
and U5379 (N_5379,N_89,N_1523);
xnor U5380 (N_5380,N_4522,N_4975);
or U5381 (N_5381,N_1804,N_242);
or U5382 (N_5382,N_3882,N_3210);
and U5383 (N_5383,N_87,N_4834);
or U5384 (N_5384,N_2646,N_2582);
and U5385 (N_5385,N_1954,N_638);
and U5386 (N_5386,N_1096,N_1616);
and U5387 (N_5387,N_3788,N_1266);
nand U5388 (N_5388,N_1807,N_206);
or U5389 (N_5389,N_3501,N_2466);
nand U5390 (N_5390,N_678,N_1043);
nand U5391 (N_5391,N_3058,N_2320);
and U5392 (N_5392,N_2033,N_4231);
and U5393 (N_5393,N_2694,N_4566);
xnor U5394 (N_5394,N_1568,N_2018);
nand U5395 (N_5395,N_2188,N_2097);
or U5396 (N_5396,N_3450,N_943);
nor U5397 (N_5397,N_1644,N_4268);
xor U5398 (N_5398,N_4063,N_2886);
xnor U5399 (N_5399,N_3117,N_4338);
xnor U5400 (N_5400,N_2353,N_2072);
nand U5401 (N_5401,N_3512,N_1326);
and U5402 (N_5402,N_588,N_3444);
nand U5403 (N_5403,N_2967,N_2555);
and U5404 (N_5404,N_1769,N_4590);
or U5405 (N_5405,N_1191,N_372);
nor U5406 (N_5406,N_276,N_2567);
nor U5407 (N_5407,N_1421,N_1621);
xor U5408 (N_5408,N_3762,N_2199);
and U5409 (N_5409,N_4694,N_690);
nand U5410 (N_5410,N_3477,N_2802);
and U5411 (N_5411,N_786,N_2951);
nand U5412 (N_5412,N_2428,N_1899);
nand U5413 (N_5413,N_426,N_2834);
nand U5414 (N_5414,N_3398,N_2780);
nand U5415 (N_5415,N_2113,N_4071);
or U5416 (N_5416,N_2400,N_302);
and U5417 (N_5417,N_3095,N_4761);
nor U5418 (N_5418,N_3270,N_3765);
or U5419 (N_5419,N_1175,N_4408);
or U5420 (N_5420,N_717,N_3235);
and U5421 (N_5421,N_1760,N_2701);
nand U5422 (N_5422,N_4753,N_2911);
nor U5423 (N_5423,N_416,N_1012);
and U5424 (N_5424,N_3141,N_512);
nand U5425 (N_5425,N_1476,N_2708);
and U5426 (N_5426,N_2515,N_560);
xor U5427 (N_5427,N_1753,N_4105);
nor U5428 (N_5428,N_1697,N_1624);
nor U5429 (N_5429,N_4528,N_3369);
or U5430 (N_5430,N_4744,N_3256);
xnor U5431 (N_5431,N_628,N_1027);
nand U5432 (N_5432,N_4091,N_1058);
nor U5433 (N_5433,N_4751,N_877);
and U5434 (N_5434,N_715,N_4436);
nand U5435 (N_5435,N_152,N_3321);
xnor U5436 (N_5436,N_595,N_2285);
or U5437 (N_5437,N_173,N_4450);
nor U5438 (N_5438,N_3417,N_4136);
xor U5439 (N_5439,N_3717,N_2993);
nand U5440 (N_5440,N_2704,N_4319);
and U5441 (N_5441,N_2772,N_1367);
xor U5442 (N_5442,N_3608,N_66);
or U5443 (N_5443,N_3345,N_1933);
and U5444 (N_5444,N_224,N_2946);
nor U5445 (N_5445,N_1876,N_1055);
nand U5446 (N_5446,N_3397,N_3174);
nor U5447 (N_5447,N_539,N_4115);
and U5448 (N_5448,N_2603,N_3458);
xor U5449 (N_5449,N_985,N_2307);
nor U5450 (N_5450,N_4188,N_3944);
nor U5451 (N_5451,N_812,N_4900);
nor U5452 (N_5452,N_3272,N_43);
nor U5453 (N_5453,N_2561,N_4942);
or U5454 (N_5454,N_4011,N_2109);
and U5455 (N_5455,N_704,N_125);
and U5456 (N_5456,N_16,N_1751);
and U5457 (N_5457,N_996,N_1927);
and U5458 (N_5458,N_4684,N_3565);
nand U5459 (N_5459,N_3632,N_3960);
or U5460 (N_5460,N_3693,N_1726);
nor U5461 (N_5461,N_4551,N_145);
or U5462 (N_5462,N_2659,N_2187);
or U5463 (N_5463,N_2528,N_3795);
and U5464 (N_5464,N_3987,N_2920);
or U5465 (N_5465,N_2323,N_1124);
nand U5466 (N_5466,N_4440,N_2738);
nor U5467 (N_5467,N_4686,N_3404);
xnor U5468 (N_5468,N_4858,N_4494);
nor U5469 (N_5469,N_3207,N_1145);
and U5470 (N_5470,N_3858,N_2666);
nor U5471 (N_5471,N_1825,N_469);
and U5472 (N_5472,N_4346,N_3582);
and U5473 (N_5473,N_3309,N_4672);
or U5474 (N_5474,N_4593,N_1345);
or U5475 (N_5475,N_3866,N_1657);
nand U5476 (N_5476,N_647,N_1332);
and U5477 (N_5477,N_4061,N_3187);
nor U5478 (N_5478,N_653,N_4067);
and U5479 (N_5479,N_4108,N_4047);
or U5480 (N_5480,N_803,N_4388);
nand U5481 (N_5481,N_2257,N_2052);
and U5482 (N_5482,N_2661,N_1403);
and U5483 (N_5483,N_2564,N_3782);
or U5484 (N_5484,N_1443,N_4144);
and U5485 (N_5485,N_1736,N_492);
or U5486 (N_5486,N_2611,N_546);
nor U5487 (N_5487,N_1301,N_4947);
or U5488 (N_5488,N_4888,N_1950);
and U5489 (N_5489,N_3025,N_1543);
xnor U5490 (N_5490,N_3203,N_2581);
and U5491 (N_5491,N_2864,N_1235);
and U5492 (N_5492,N_4752,N_1576);
nor U5493 (N_5493,N_1806,N_709);
xor U5494 (N_5494,N_1022,N_204);
nand U5495 (N_5495,N_107,N_4607);
or U5496 (N_5496,N_1202,N_3375);
or U5497 (N_5497,N_2210,N_3912);
or U5498 (N_5498,N_4978,N_1408);
nand U5499 (N_5499,N_4299,N_890);
nand U5500 (N_5500,N_2029,N_2364);
or U5501 (N_5501,N_1551,N_4220);
nor U5502 (N_5502,N_86,N_3695);
nor U5503 (N_5503,N_2797,N_3134);
nor U5504 (N_5504,N_3840,N_935);
nand U5505 (N_5505,N_2628,N_2128);
xnor U5506 (N_5506,N_362,N_1659);
nor U5507 (N_5507,N_3342,N_1296);
nand U5508 (N_5508,N_4812,N_1427);
xnor U5509 (N_5509,N_1455,N_604);
nand U5510 (N_5510,N_700,N_309);
and U5511 (N_5511,N_2718,N_2637);
nor U5512 (N_5512,N_4163,N_3967);
nand U5513 (N_5513,N_2550,N_3426);
and U5514 (N_5514,N_2366,N_1801);
nand U5515 (N_5515,N_3839,N_4218);
or U5516 (N_5516,N_1667,N_3778);
nand U5517 (N_5517,N_809,N_1536);
nor U5518 (N_5518,N_1148,N_2079);
or U5519 (N_5519,N_4339,N_4870);
nand U5520 (N_5520,N_2385,N_1445);
nand U5521 (N_5521,N_2456,N_1812);
xor U5522 (N_5522,N_4251,N_3431);
or U5523 (N_5523,N_2338,N_2560);
or U5524 (N_5524,N_4984,N_83);
and U5525 (N_5525,N_2162,N_3057);
nand U5526 (N_5526,N_3665,N_3301);
and U5527 (N_5527,N_4819,N_4779);
nand U5528 (N_5528,N_3128,N_2026);
nand U5529 (N_5529,N_789,N_2010);
nor U5530 (N_5530,N_4612,N_239);
nor U5531 (N_5531,N_600,N_643);
nor U5532 (N_5532,N_2553,N_2389);
xor U5533 (N_5533,N_3641,N_2009);
or U5534 (N_5534,N_646,N_4206);
nor U5535 (N_5535,N_29,N_3003);
nand U5536 (N_5536,N_3097,N_264);
or U5537 (N_5537,N_2325,N_370);
nand U5538 (N_5538,N_3682,N_1696);
xnor U5539 (N_5539,N_1771,N_4204);
nor U5540 (N_5540,N_680,N_30);
and U5541 (N_5541,N_1962,N_255);
xnor U5542 (N_5542,N_1589,N_307);
nand U5543 (N_5543,N_4791,N_2332);
nand U5544 (N_5544,N_4198,N_2511);
nand U5545 (N_5545,N_449,N_3503);
nor U5546 (N_5546,N_4057,N_4400);
and U5547 (N_5547,N_1907,N_1172);
xor U5548 (N_5548,N_1727,N_2677);
or U5549 (N_5549,N_3405,N_2895);
nand U5550 (N_5550,N_933,N_1194);
and U5551 (N_5551,N_3005,N_495);
nand U5552 (N_5552,N_3580,N_1780);
and U5553 (N_5553,N_75,N_4560);
and U5554 (N_5554,N_104,N_3052);
xnor U5555 (N_5555,N_4173,N_2301);
xor U5556 (N_5556,N_1779,N_3980);
or U5557 (N_5557,N_2081,N_4591);
nand U5558 (N_5558,N_1669,N_3089);
and U5559 (N_5559,N_4994,N_3457);
or U5560 (N_5560,N_273,N_765);
xnor U5561 (N_5561,N_2415,N_2500);
or U5562 (N_5562,N_2803,N_108);
or U5563 (N_5563,N_2692,N_4619);
and U5564 (N_5564,N_291,N_2310);
nor U5565 (N_5565,N_1694,N_2432);
and U5566 (N_5566,N_486,N_1115);
and U5567 (N_5567,N_1997,N_2619);
nand U5568 (N_5568,N_4154,N_4537);
or U5569 (N_5569,N_1569,N_4874);
or U5570 (N_5570,N_4582,N_2942);
nand U5571 (N_5571,N_3299,N_559);
nand U5572 (N_5572,N_3463,N_4117);
or U5573 (N_5573,N_2516,N_3425);
and U5574 (N_5574,N_1357,N_774);
and U5575 (N_5575,N_209,N_4781);
and U5576 (N_5576,N_24,N_1469);
nand U5577 (N_5577,N_3587,N_435);
nand U5578 (N_5578,N_4307,N_237);
or U5579 (N_5579,N_4233,N_4033);
nand U5580 (N_5580,N_369,N_3885);
nand U5581 (N_5581,N_936,N_2324);
nand U5582 (N_5582,N_2386,N_1864);
or U5583 (N_5583,N_3433,N_1003);
or U5584 (N_5584,N_3544,N_1337);
nor U5585 (N_5585,N_4962,N_182);
nand U5586 (N_5586,N_1195,N_1539);
or U5587 (N_5587,N_2453,N_1014);
xnor U5588 (N_5588,N_3567,N_528);
and U5589 (N_5589,N_1805,N_3662);
nand U5590 (N_5590,N_4355,N_2085);
and U5591 (N_5591,N_4987,N_2326);
xnor U5592 (N_5592,N_2204,N_2119);
xor U5593 (N_5593,N_1558,N_2762);
and U5594 (N_5594,N_4194,N_4926);
nor U5595 (N_5595,N_1875,N_3624);
nor U5596 (N_5596,N_3557,N_199);
nor U5597 (N_5597,N_3083,N_4140);
nor U5598 (N_5598,N_466,N_3763);
or U5599 (N_5599,N_1628,N_4843);
nor U5600 (N_5600,N_4157,N_3543);
nand U5601 (N_5601,N_4968,N_889);
nor U5602 (N_5602,N_4372,N_3344);
and U5603 (N_5603,N_2159,N_3764);
and U5604 (N_5604,N_2867,N_3548);
nor U5605 (N_5605,N_3754,N_1708);
nor U5606 (N_5606,N_4539,N_3919);
or U5607 (N_5607,N_2431,N_549);
or U5608 (N_5608,N_4754,N_3698);
nand U5609 (N_5609,N_4958,N_1139);
nor U5610 (N_5610,N_3791,N_3798);
nand U5611 (N_5611,N_2623,N_581);
xnor U5612 (N_5612,N_3875,N_4920);
xnor U5613 (N_5613,N_3153,N_1759);
and U5614 (N_5614,N_4825,N_785);
nand U5615 (N_5615,N_897,N_3887);
xnor U5616 (N_5616,N_817,N_4244);
nand U5617 (N_5617,N_3343,N_875);
or U5618 (N_5618,N_1293,N_1620);
xnor U5619 (N_5619,N_4993,N_1090);
nor U5620 (N_5620,N_189,N_3745);
nor U5621 (N_5621,N_3531,N_90);
nand U5622 (N_5622,N_1656,N_3743);
nor U5623 (N_5623,N_4899,N_3768);
and U5624 (N_5624,N_4996,N_2534);
xor U5625 (N_5625,N_248,N_1129);
or U5626 (N_5626,N_4069,N_4081);
nand U5627 (N_5627,N_2357,N_4131);
nor U5628 (N_5628,N_751,N_1917);
and U5629 (N_5629,N_2343,N_1241);
or U5630 (N_5630,N_4500,N_997);
and U5631 (N_5631,N_1265,N_2570);
and U5632 (N_5632,N_3572,N_2949);
nor U5633 (N_5633,N_670,N_4668);
nand U5634 (N_5634,N_1862,N_1707);
nand U5635 (N_5635,N_2464,N_1748);
or U5636 (N_5636,N_2781,N_4125);
and U5637 (N_5637,N_2145,N_1503);
and U5638 (N_5638,N_1583,N_2149);
or U5639 (N_5639,N_2535,N_4650);
and U5640 (N_5640,N_745,N_3186);
xor U5641 (N_5641,N_2594,N_2088);
nand U5642 (N_5642,N_584,N_1071);
nor U5643 (N_5643,N_1402,N_4806);
nor U5644 (N_5644,N_696,N_2423);
or U5645 (N_5645,N_2165,N_3420);
or U5646 (N_5646,N_2054,N_1686);
and U5647 (N_5647,N_1480,N_366);
nor U5648 (N_5648,N_119,N_312);
and U5649 (N_5649,N_1973,N_1381);
and U5650 (N_5650,N_2391,N_4616);
and U5651 (N_5651,N_4208,N_131);
and U5652 (N_5652,N_1444,N_4635);
nor U5653 (N_5653,N_522,N_2208);
nand U5654 (N_5654,N_3080,N_2584);
nand U5655 (N_5655,N_3250,N_2656);
nand U5656 (N_5656,N_4782,N_4207);
and U5657 (N_5657,N_3677,N_250);
nand U5658 (N_5658,N_2252,N_4312);
or U5659 (N_5659,N_2048,N_2465);
nor U5660 (N_5660,N_1762,N_597);
or U5661 (N_5661,N_3954,N_953);
xnor U5662 (N_5662,N_2489,N_4666);
nand U5663 (N_5663,N_4944,N_2904);
xor U5664 (N_5664,N_689,N_3522);
nor U5665 (N_5665,N_2627,N_4146);
nand U5666 (N_5666,N_1765,N_713);
nor U5667 (N_5667,N_2485,N_2209);
and U5668 (N_5668,N_3337,N_1284);
nand U5669 (N_5669,N_4988,N_990);
nor U5670 (N_5670,N_3465,N_961);
and U5671 (N_5671,N_4288,N_3468);
nand U5672 (N_5672,N_2734,N_2176);
nand U5673 (N_5673,N_3895,N_2399);
and U5674 (N_5674,N_1829,N_503);
or U5675 (N_5675,N_437,N_4168);
or U5676 (N_5676,N_23,N_3378);
or U5677 (N_5677,N_1580,N_2484);
or U5678 (N_5678,N_3892,N_2377);
or U5679 (N_5679,N_3300,N_3112);
nand U5680 (N_5680,N_2057,N_2729);
nand U5681 (N_5681,N_2926,N_4689);
nand U5682 (N_5682,N_1057,N_1041);
nand U5683 (N_5683,N_1668,N_972);
nand U5684 (N_5684,N_2722,N_2641);
and U5685 (N_5685,N_4004,N_470);
and U5686 (N_5686,N_4905,N_1920);
xnor U5687 (N_5687,N_3026,N_2643);
nor U5688 (N_5688,N_2425,N_1312);
nand U5689 (N_5689,N_3729,N_4297);
and U5690 (N_5690,N_1389,N_3708);
nand U5691 (N_5691,N_3084,N_2095);
nor U5692 (N_5692,N_1246,N_3412);
or U5693 (N_5693,N_4990,N_3317);
and U5694 (N_5694,N_1223,N_3737);
nor U5695 (N_5695,N_4784,N_583);
and U5696 (N_5696,N_3976,N_4083);
or U5697 (N_5697,N_4192,N_2426);
nor U5698 (N_5698,N_1957,N_1141);
and U5699 (N_5699,N_2011,N_4629);
nand U5700 (N_5700,N_4951,N_1948);
or U5701 (N_5701,N_1103,N_159);
nor U5702 (N_5702,N_4141,N_360);
xor U5703 (N_5703,N_2083,N_2137);
or U5704 (N_5704,N_3915,N_2640);
nor U5705 (N_5705,N_3208,N_4250);
and U5706 (N_5706,N_324,N_3287);
xor U5707 (N_5707,N_2678,N_2441);
nand U5708 (N_5708,N_3711,N_419);
or U5709 (N_5709,N_3995,N_1275);
nand U5710 (N_5710,N_1209,N_4946);
nor U5711 (N_5711,N_2265,N_3821);
and U5712 (N_5712,N_513,N_2120);
nand U5713 (N_5713,N_2256,N_1489);
nor U5714 (N_5714,N_2622,N_3516);
nand U5715 (N_5715,N_1548,N_1199);
xor U5716 (N_5716,N_1729,N_3519);
nand U5717 (N_5717,N_3925,N_4002);
and U5718 (N_5718,N_2374,N_1187);
nand U5719 (N_5719,N_2731,N_4249);
and U5720 (N_5720,N_280,N_2938);
or U5721 (N_5721,N_2573,N_165);
and U5722 (N_5722,N_4881,N_938);
or U5723 (N_5723,N_4611,N_2045);
nand U5724 (N_5724,N_2370,N_901);
nor U5725 (N_5725,N_3360,N_623);
and U5726 (N_5726,N_11,N_862);
and U5727 (N_5727,N_3655,N_4001);
nand U5728 (N_5728,N_2458,N_3755);
nand U5729 (N_5729,N_2847,N_843);
nor U5730 (N_5730,N_4457,N_884);
xor U5731 (N_5731,N_4829,N_3962);
nor U5732 (N_5732,N_4816,N_561);
nor U5733 (N_5733,N_2181,N_1673);
nand U5734 (N_5734,N_404,N_1288);
and U5735 (N_5735,N_3487,N_2140);
nor U5736 (N_5736,N_1662,N_4762);
nand U5737 (N_5737,N_532,N_1217);
nand U5738 (N_5738,N_1977,N_3143);
nor U5739 (N_5739,N_3271,N_4508);
xor U5740 (N_5740,N_2270,N_758);
nand U5741 (N_5741,N_2163,N_97);
nor U5742 (N_5742,N_906,N_364);
nand U5743 (N_5743,N_3932,N_3159);
and U5744 (N_5744,N_1144,N_3447);
nand U5745 (N_5745,N_2342,N_2099);
and U5746 (N_5746,N_1884,N_3859);
nand U5747 (N_5747,N_4476,N_31);
nor U5748 (N_5748,N_1392,N_3952);
and U5749 (N_5749,N_3064,N_589);
or U5750 (N_5750,N_2114,N_3700);
nor U5751 (N_5751,N_4006,N_4234);
nand U5752 (N_5752,N_2064,N_4282);
and U5753 (N_5753,N_4129,N_2956);
nand U5754 (N_5754,N_1493,N_3062);
or U5755 (N_5755,N_4568,N_4052);
xnor U5756 (N_5756,N_3322,N_2340);
and U5757 (N_5757,N_1354,N_2625);
nor U5758 (N_5758,N_3618,N_3335);
and U5759 (N_5759,N_325,N_2202);
or U5760 (N_5760,N_2254,N_3157);
xor U5761 (N_5761,N_577,N_1256);
nor U5762 (N_5762,N_2070,N_920);
or U5763 (N_5763,N_1852,N_4254);
or U5764 (N_5764,N_3332,N_3410);
or U5765 (N_5765,N_3726,N_1510);
or U5766 (N_5766,N_3841,N_810);
nand U5767 (N_5767,N_596,N_1893);
nand U5768 (N_5768,N_2190,N_2129);
nor U5769 (N_5769,N_4166,N_1712);
nor U5770 (N_5770,N_4236,N_34);
xor U5771 (N_5771,N_2647,N_1774);
nor U5772 (N_5772,N_855,N_3540);
and U5773 (N_5773,N_1793,N_386);
and U5774 (N_5774,N_3678,N_3734);
and U5775 (N_5775,N_1994,N_2796);
xor U5776 (N_5776,N_537,N_60);
nand U5777 (N_5777,N_3842,N_208);
and U5778 (N_5778,N_4770,N_1364);
or U5779 (N_5779,N_1790,N_4937);
nand U5780 (N_5780,N_1371,N_140);
nor U5781 (N_5781,N_2615,N_2791);
nand U5782 (N_5782,N_1358,N_3637);
and U5783 (N_5783,N_3390,N_50);
nand U5784 (N_5784,N_822,N_1623);
nor U5785 (N_5785,N_2958,N_1642);
and U5786 (N_5786,N_2347,N_2930);
nor U5787 (N_5787,N_4371,N_2060);
xor U5788 (N_5788,N_379,N_3180);
xor U5789 (N_5789,N_3672,N_952);
or U5790 (N_5790,N_2713,N_2043);
nand U5791 (N_5791,N_4609,N_2524);
nand U5792 (N_5792,N_1238,N_4349);
xor U5793 (N_5793,N_25,N_1522);
and U5794 (N_5794,N_180,N_2049);
and U5795 (N_5795,N_3365,N_1912);
nor U5796 (N_5796,N_878,N_2266);
xnor U5797 (N_5797,N_2268,N_518);
and U5798 (N_5798,N_4227,N_3829);
nor U5799 (N_5799,N_3480,N_134);
and U5800 (N_5800,N_2420,N_1494);
or U5801 (N_5801,N_1230,N_2635);
or U5802 (N_5802,N_438,N_215);
nor U5803 (N_5803,N_4599,N_3121);
xor U5804 (N_5804,N_3261,N_1215);
and U5805 (N_5805,N_2664,N_4383);
nand U5806 (N_5806,N_525,N_3206);
or U5807 (N_5807,N_1404,N_2012);
and U5808 (N_5808,N_3432,N_3096);
nor U5809 (N_5809,N_3689,N_2720);
or U5810 (N_5810,N_3355,N_4109);
nor U5811 (N_5811,N_284,N_1023);
nand U5812 (N_5812,N_956,N_3105);
nor U5813 (N_5813,N_4342,N_2632);
nand U5814 (N_5814,N_2080,N_475);
and U5815 (N_5815,N_4919,N_3537);
or U5816 (N_5816,N_1401,N_247);
and U5817 (N_5817,N_4902,N_1613);
or U5818 (N_5818,N_4425,N_3285);
or U5819 (N_5819,N_1622,N_153);
nor U5820 (N_5820,N_3616,N_2830);
nand U5821 (N_5821,N_4232,N_2082);
xnor U5822 (N_5822,N_2379,N_1626);
or U5823 (N_5823,N_4997,N_293);
nor U5824 (N_5824,N_2983,N_3732);
nor U5825 (N_5825,N_4716,N_2196);
nand U5826 (N_5826,N_3449,N_4561);
xor U5827 (N_5827,N_3747,N_4169);
or U5828 (N_5828,N_4601,N_149);
nor U5829 (N_5829,N_409,N_2100);
or U5830 (N_5830,N_491,N_2004);
and U5831 (N_5831,N_1918,N_4414);
nor U5832 (N_5832,N_155,N_3596);
nor U5833 (N_5833,N_4266,N_4645);
nor U5834 (N_5834,N_2809,N_4894);
nor U5835 (N_5835,N_3136,N_2373);
nor U5836 (N_5836,N_4306,N_2799);
or U5837 (N_5837,N_361,N_1897);
nand U5838 (N_5838,N_2259,N_2461);
nand U5839 (N_5839,N_4170,N_1287);
or U5840 (N_5840,N_1157,N_6);
nor U5841 (N_5841,N_161,N_2078);
nand U5842 (N_5842,N_1333,N_3939);
nand U5843 (N_5843,N_4658,N_4417);
nor U5844 (N_5844,N_547,N_2490);
and U5845 (N_5845,N_2823,N_4300);
nor U5846 (N_5846,N_2754,N_4841);
or U5847 (N_5847,N_3937,N_2236);
or U5848 (N_5848,N_3328,N_1219);
nor U5849 (N_5849,N_4692,N_2092);
nand U5850 (N_5850,N_4554,N_3586);
or U5851 (N_5851,N_946,N_1356);
nor U5852 (N_5852,N_705,N_1650);
and U5853 (N_5853,N_1122,N_599);
nor U5854 (N_5854,N_401,N_856);
nor U5855 (N_5855,N_2916,N_1386);
or U5856 (N_5856,N_3617,N_3931);
and U5857 (N_5857,N_736,N_4803);
and U5858 (N_5858,N_2868,N_3467);
and U5859 (N_5859,N_3257,N_318);
nand U5860 (N_5860,N_4780,N_4866);
nor U5861 (N_5861,N_3576,N_2407);
nor U5862 (N_5862,N_4277,N_2529);
or U5863 (N_5863,N_740,N_463);
or U5864 (N_5864,N_4597,N_1883);
nor U5865 (N_5865,N_904,N_2742);
or U5866 (N_5866,N_3329,N_241);
nand U5867 (N_5867,N_3538,N_819);
and U5868 (N_5868,N_1819,N_3706);
nor U5869 (N_5869,N_2316,N_2194);
xnor U5870 (N_5870,N_640,N_1340);
nor U5871 (N_5871,N_3229,N_669);
nor U5872 (N_5872,N_3922,N_2022);
nand U5873 (N_5873,N_1573,N_151);
nor U5874 (N_5874,N_2273,N_4833);
nand U5875 (N_5875,N_3724,N_2198);
xnor U5876 (N_5876,N_1277,N_1987);
xor U5877 (N_5877,N_1716,N_4323);
nor U5878 (N_5878,N_962,N_766);
and U5879 (N_5879,N_4973,N_1777);
nand U5880 (N_5880,N_633,N_3552);
and U5881 (N_5881,N_26,N_1167);
and U5882 (N_5882,N_2028,N_3198);
or U5883 (N_5883,N_2702,N_3231);
and U5884 (N_5884,N_3048,N_842);
and U5885 (N_5885,N_4680,N_4014);
or U5886 (N_5886,N_4382,N_4969);
nand U5887 (N_5887,N_1869,N_3138);
or U5888 (N_5888,N_4511,N_3738);
xnor U5889 (N_5889,N_4172,N_4709);
xnor U5890 (N_5890,N_681,N_326);
xnor U5891 (N_5891,N_3490,N_4135);
nand U5892 (N_5892,N_3040,N_3645);
or U5893 (N_5893,N_4712,N_456);
nor U5894 (N_5894,N_1009,N_3757);
and U5895 (N_5895,N_1934,N_4482);
or U5896 (N_5896,N_2884,N_4394);
nor U5897 (N_5897,N_3736,N_490);
nor U5898 (N_5898,N_3389,N_4901);
nor U5899 (N_5899,N_727,N_3914);
nand U5900 (N_5900,N_331,N_3897);
or U5901 (N_5901,N_3316,N_3881);
nor U5902 (N_5902,N_887,N_2107);
xor U5903 (N_5903,N_2617,N_4276);
nor U5904 (N_5904,N_3181,N_4533);
nand U5905 (N_5905,N_907,N_2843);
or U5906 (N_5906,N_2517,N_4087);
or U5907 (N_5907,N_1185,N_948);
nand U5908 (N_5908,N_3959,N_2786);
nor U5909 (N_5909,N_4506,N_4704);
nor U5910 (N_5910,N_4221,N_1989);
and U5911 (N_5911,N_4661,N_2059);
nand U5912 (N_5912,N_2102,N_3496);
and U5913 (N_5913,N_4648,N_2189);
nand U5914 (N_5914,N_4341,N_3071);
nor U5915 (N_5915,N_127,N_4358);
and U5916 (N_5916,N_2205,N_163);
or U5917 (N_5917,N_1184,N_4097);
and U5918 (N_5918,N_2115,N_3010);
nor U5919 (N_5919,N_4316,N_2750);
or U5920 (N_5920,N_459,N_1750);
and U5921 (N_5921,N_4452,N_3205);
xor U5922 (N_5922,N_1856,N_3464);
xor U5923 (N_5923,N_4583,N_3419);
nand U5924 (N_5924,N_510,N_734);
nor U5925 (N_5925,N_2753,N_2154);
or U5926 (N_5926,N_3030,N_2901);
or U5927 (N_5927,N_2624,N_4497);
and U5928 (N_5928,N_441,N_3438);
nor U5929 (N_5929,N_2443,N_4831);
nand U5930 (N_5930,N_3916,N_971);
nand U5931 (N_5931,N_1908,N_1422);
nor U5932 (N_5932,N_1574,N_1646);
or U5933 (N_5933,N_3871,N_3352);
or U5934 (N_5934,N_2812,N_2329);
and U5935 (N_5935,N_1415,N_1232);
nand U5936 (N_5936,N_2291,N_2861);
or U5937 (N_5937,N_4260,N_1930);
nand U5938 (N_5938,N_3116,N_905);
nand U5939 (N_5939,N_1068,N_1504);
or U5940 (N_5940,N_1044,N_4971);
nor U5941 (N_5941,N_4632,N_2419);
xor U5942 (N_5942,N_2539,N_2369);
nand U5943 (N_5943,N_4008,N_4096);
and U5944 (N_5944,N_2569,N_1931);
nand U5945 (N_5945,N_2481,N_3019);
or U5946 (N_5946,N_1169,N_3204);
nor U5947 (N_5947,N_4364,N_891);
and U5948 (N_5948,N_3042,N_1116);
or U5949 (N_5949,N_791,N_3772);
and U5950 (N_5950,N_1586,N_4553);
nand U5951 (N_5951,N_36,N_2831);
and U5952 (N_5952,N_229,N_1944);
and U5953 (N_5953,N_4577,N_795);
or U5954 (N_5954,N_4189,N_721);
nand U5955 (N_5955,N_611,N_4764);
nor U5956 (N_5956,N_1242,N_691);
nand U5957 (N_5957,N_4272,N_1362);
nor U5958 (N_5958,N_1015,N_389);
and U5959 (N_5959,N_4088,N_4448);
nand U5960 (N_5960,N_3305,N_53);
nor U5961 (N_5961,N_2132,N_912);
nand U5962 (N_5962,N_1506,N_776);
or U5963 (N_5963,N_4887,N_4983);
nor U5964 (N_5964,N_3564,N_4099);
or U5965 (N_5965,N_141,N_886);
nor U5966 (N_5966,N_3059,N_652);
nor U5967 (N_5967,N_3851,N_3346);
and U5968 (N_5968,N_415,N_1082);
and U5969 (N_5969,N_221,N_978);
nand U5970 (N_5970,N_4401,N_3721);
or U5971 (N_5971,N_2639,N_726);
nor U5972 (N_5972,N_4242,N_1649);
or U5973 (N_5973,N_2696,N_497);
or U5974 (N_5974,N_1200,N_2037);
nand U5975 (N_5975,N_2067,N_2869);
or U5976 (N_5976,N_3293,N_573);
or U5977 (N_5977,N_698,N_2055);
xnor U5978 (N_5978,N_3896,N_3853);
and U5979 (N_5979,N_4945,N_1212);
and U5980 (N_5980,N_3521,N_3661);
and U5981 (N_5981,N_1783,N_1142);
nor U5982 (N_5982,N_3785,N_1229);
and U5983 (N_5983,N_1505,N_332);
or U5984 (N_5984,N_723,N_2510);
and U5985 (N_5985,N_4956,N_450);
nand U5986 (N_5986,N_3371,N_613);
or U5987 (N_5987,N_3683,N_4606);
xor U5988 (N_5988,N_3864,N_1681);
nor U5989 (N_5989,N_1315,N_4848);
nand U5990 (N_5990,N_2981,N_4229);
and U5991 (N_5991,N_2723,N_3087);
nor U5992 (N_5992,N_3101,N_2853);
nand U5993 (N_5993,N_3669,N_679);
xnor U5994 (N_5994,N_4015,N_2138);
nand U5995 (N_5995,N_420,N_3623);
or U5996 (N_5996,N_4060,N_310);
nor U5997 (N_5997,N_3822,N_482);
and U5998 (N_5998,N_1619,N_222);
or U5999 (N_5999,N_913,N_1795);
or U6000 (N_6000,N_2378,N_4512);
and U6001 (N_6001,N_4032,N_1741);
xnor U6002 (N_6002,N_3810,N_1865);
nand U6003 (N_6003,N_3607,N_2726);
or U6004 (N_6004,N_4347,N_1538);
or U6005 (N_6005,N_4721,N_1787);
or U6006 (N_6006,N_3780,N_3442);
nand U6007 (N_6007,N_1595,N_1960);
nand U6008 (N_6008,N_3730,N_4193);
nand U6009 (N_6009,N_2574,N_297);
and U6010 (N_6010,N_1013,N_796);
xor U6011 (N_6011,N_2710,N_1037);
nor U6012 (N_6012,N_3188,N_3192);
nand U6013 (N_6013,N_390,N_3045);
nor U6014 (N_6014,N_880,N_3921);
nand U6015 (N_6015,N_755,N_4243);
xor U6016 (N_6016,N_4441,N_3441);
xnor U6017 (N_6017,N_4284,N_3015);
and U6018 (N_6018,N_2171,N_3869);
or U6019 (N_6019,N_3122,N_2496);
nor U6020 (N_6020,N_3094,N_2747);
nand U6021 (N_6021,N_1911,N_1743);
or U6022 (N_6022,N_4817,N_2298);
nand U6023 (N_6023,N_1674,N_2784);
nor U6024 (N_6024,N_203,N_1839);
and U6025 (N_6025,N_61,N_2362);
xnor U6026 (N_6026,N_4510,N_4444);
xor U6027 (N_6027,N_3891,N_2308);
nor U6028 (N_6028,N_885,N_1527);
nand U6029 (N_6029,N_818,N_3578);
or U6030 (N_6030,N_601,N_1841);
or U6031 (N_6031,N_1641,N_1871);
and U6032 (N_6032,N_1904,N_1125);
nand U6033 (N_6033,N_3255,N_2665);
or U6034 (N_6034,N_3408,N_2039);
and U6035 (N_6035,N_3773,N_2317);
nor U6036 (N_6036,N_2744,N_1094);
nand U6037 (N_6037,N_873,N_570);
and U6038 (N_6038,N_945,N_1975);
nand U6039 (N_6039,N_4420,N_2883);
or U6040 (N_6040,N_4563,N_949);
xnor U6041 (N_6041,N_4714,N_2881);
or U6042 (N_6042,N_3036,N_658);
nor U6043 (N_6043,N_1112,N_4748);
or U6044 (N_6044,N_3004,N_650);
and U6045 (N_6045,N_1325,N_1035);
and U6046 (N_6046,N_3199,N_2360);
or U6047 (N_6047,N_3476,N_2968);
and U6048 (N_6048,N_3158,N_509);
nand U6049 (N_6049,N_1458,N_282);
nand U6050 (N_6050,N_1130,N_3575);
nor U6051 (N_6051,N_4737,N_2444);
or U6052 (N_6052,N_1498,N_816);
nor U6053 (N_6053,N_2591,N_1915);
and U6054 (N_6054,N_96,N_465);
nor U6055 (N_6055,N_4844,N_3709);
nor U6056 (N_6056,N_448,N_3535);
or U6057 (N_6057,N_4543,N_4548);
and U6058 (N_6058,N_3603,N_4333);
and U6059 (N_6059,N_2538,N_77);
or U6060 (N_6060,N_2848,N_4211);
nand U6061 (N_6061,N_410,N_3466);
or U6062 (N_6062,N_278,N_4574);
nand U6063 (N_6063,N_2486,N_625);
and U6064 (N_6064,N_2768,N_2827);
or U6065 (N_6065,N_586,N_2689);
nand U6066 (N_6066,N_4974,N_78);
nand U6067 (N_6067,N_3982,N_4380);
or U6068 (N_6068,N_2435,N_3579);
nand U6069 (N_6069,N_2242,N_3597);
xor U6070 (N_6070,N_164,N_4741);
xnor U6071 (N_6071,N_176,N_4134);
or U6072 (N_6072,N_3832,N_2932);
xor U6073 (N_6073,N_1537,N_3570);
nor U6074 (N_6074,N_2998,N_3926);
and U6075 (N_6075,N_2987,N_916);
nor U6076 (N_6076,N_2182,N_500);
nor U6077 (N_6077,N_2434,N_2894);
and U6078 (N_6078,N_674,N_4637);
nor U6079 (N_6079,N_4734,N_2682);
and U6080 (N_6080,N_4385,N_3536);
or U6081 (N_6081,N_1341,N_1749);
nand U6082 (N_6082,N_1581,N_4195);
nand U6083 (N_6083,N_637,N_2151);
nand U6084 (N_6084,N_3230,N_1137);
or U6085 (N_6085,N_202,N_683);
xnor U6086 (N_6086,N_3913,N_544);
nand U6087 (N_6087,N_1064,N_4732);
nand U6088 (N_6088,N_802,N_1181);
or U6089 (N_6089,N_1482,N_4089);
or U6090 (N_6090,N_729,N_2996);
or U6091 (N_6091,N_319,N_4344);
nor U6092 (N_6092,N_3308,N_4907);
nand U6093 (N_6093,N_1143,N_4378);
nand U6094 (N_6094,N_3551,N_3969);
and U6095 (N_6095,N_3511,N_1460);
nand U6096 (N_6096,N_4361,N_3182);
nand U6097 (N_6097,N_4565,N_4222);
and U6098 (N_6098,N_2454,N_1996);
or U6099 (N_6099,N_4515,N_1881);
nor U6100 (N_6100,N_841,N_3819);
or U6101 (N_6101,N_3283,N_699);
nor U6102 (N_6102,N_4743,N_1258);
and U6103 (N_6103,N_951,N_4162);
nand U6104 (N_6104,N_112,N_2587);
xnor U6105 (N_6105,N_3560,N_2513);
and U6106 (N_6106,N_1761,N_2514);
and U6107 (N_6107,N_2969,N_869);
nand U6108 (N_6108,N_1747,N_576);
or U6109 (N_6109,N_2153,N_4334);
and U6110 (N_6110,N_3699,N_2898);
nand U6111 (N_6111,N_2933,N_2790);
xor U6112 (N_6112,N_1407,N_408);
or U6113 (N_6113,N_2448,N_2498);
or U6114 (N_6114,N_1734,N_1084);
xnor U6115 (N_6115,N_2703,N_1156);
nand U6116 (N_6116,N_283,N_1690);
and U6117 (N_6117,N_4294,N_3834);
nor U6118 (N_6118,N_2631,N_3901);
xnor U6119 (N_6119,N_917,N_28);
nor U6120 (N_6120,N_1655,N_4891);
nor U6121 (N_6121,N_3908,N_3595);
and U6122 (N_6122,N_4800,N_2568);
nor U6123 (N_6123,N_4031,N_4100);
nor U6124 (N_6124,N_1263,N_4718);
or U6125 (N_6125,N_4203,N_266);
nor U6126 (N_6126,N_1796,N_395);
nor U6127 (N_6127,N_4302,N_1813);
or U6128 (N_6128,N_1968,N_1453);
and U6129 (N_6129,N_260,N_3370);
nor U6130 (N_6130,N_4738,N_1803);
nor U6131 (N_6131,N_2971,N_4558);
and U6132 (N_6132,N_1370,N_3304);
nand U6133 (N_6133,N_4594,N_3681);
nand U6134 (N_6134,N_1385,N_4048);
or U6135 (N_6135,N_4729,N_2284);
nor U6136 (N_6136,N_3127,N_1449);
or U6137 (N_6137,N_2499,N_2756);
xor U6138 (N_6138,N_3383,N_4628);
xor U6139 (N_6139,N_1006,N_286);
nand U6140 (N_6140,N_1702,N_624);
nand U6141 (N_6141,N_2669,N_2698);
and U6142 (N_6142,N_12,N_1081);
nand U6143 (N_6143,N_2982,N_2674);
and U6144 (N_6144,N_2751,N_4557);
nor U6145 (N_6145,N_3701,N_1910);
nand U6146 (N_6146,N_367,N_99);
or U6147 (N_6147,N_114,N_4309);
or U6148 (N_6148,N_4291,N_4393);
xnor U6149 (N_6149,N_2395,N_3628);
nand U6150 (N_6150,N_188,N_4180);
nand U6151 (N_6151,N_1146,N_2921);
nor U6152 (N_6152,N_2788,N_4595);
nor U6153 (N_6153,N_440,N_836);
nor U6154 (N_6154,N_3867,N_3259);
nor U6155 (N_6155,N_1861,N_4713);
or U6156 (N_6156,N_3789,N_4722);
xor U6157 (N_6157,N_9,N_1833);
nand U6158 (N_6158,N_3414,N_2811);
nor U6159 (N_6159,N_40,N_1981);
xnor U6160 (N_6160,N_2116,N_3735);
and U6161 (N_6161,N_3710,N_471);
nand U6162 (N_6162,N_1397,N_3651);
xor U6163 (N_6163,N_3368,N_2685);
nor U6164 (N_6164,N_2231,N_4039);
or U6165 (N_6165,N_3125,N_3380);
or U6166 (N_6166,N_3553,N_1545);
or U6167 (N_6167,N_4631,N_1789);
or U6168 (N_6168,N_4126,N_425);
or U6169 (N_6169,N_2267,N_2424);
or U6170 (N_6170,N_1860,N_4055);
or U6171 (N_6171,N_3361,N_3622);
nand U6172 (N_6172,N_1817,N_2512);
and U6173 (N_6173,N_4756,N_3975);
nor U6174 (N_6174,N_4027,N_3715);
or U6175 (N_6175,N_1126,N_3604);
nand U6176 (N_6176,N_462,N_3555);
or U6177 (N_6177,N_4073,N_195);
and U6178 (N_6178,N_4261,N_3626);
nand U6179 (N_6179,N_3483,N_1764);
xor U6180 (N_6180,N_3883,N_3313);
nand U6181 (N_6181,N_2272,N_85);
xor U6182 (N_6182,N_1318,N_1688);
xor U6183 (N_6183,N_4391,N_4145);
or U6184 (N_6184,N_1276,N_957);
and U6185 (N_6185,N_1294,N_1150);
and U6186 (N_6186,N_256,N_2170);
nor U6187 (N_6187,N_3787,N_4473);
xnor U6188 (N_6188,N_752,N_2215);
nand U6189 (N_6189,N_564,N_1359);
and U6190 (N_6190,N_730,N_3372);
nor U6191 (N_6191,N_3401,N_2547);
nand U6192 (N_6192,N_4792,N_898);
and U6193 (N_6193,N_557,N_1369);
nor U6194 (N_6194,N_4965,N_671);
nor U6195 (N_6195,N_4463,N_2896);
nand U6196 (N_6196,N_4462,N_3148);
and U6197 (N_6197,N_998,N_814);
nor U6198 (N_6198,N_3933,N_3081);
nand U6199 (N_6199,N_2371,N_3167);
and U6200 (N_6200,N_2217,N_4960);
and U6201 (N_6201,N_2497,N_2654);
nor U6202 (N_6202,N_1138,N_4952);
or U6203 (N_6203,N_854,N_2821);
nand U6204 (N_6204,N_3992,N_3888);
or U6205 (N_6205,N_451,N_2003);
nand U6206 (N_6206,N_39,N_2150);
nand U6207 (N_6207,N_969,N_3281);
nor U6208 (N_6208,N_2405,N_3924);
and U6209 (N_6209,N_2469,N_269);
nand U6210 (N_6210,N_1111,N_428);
and U6211 (N_6211,N_892,N_3758);
nor U6212 (N_6212,N_1500,N_876);
xnor U6213 (N_6213,N_3090,N_3783);
and U6214 (N_6214,N_2372,N_4934);
and U6215 (N_6215,N_4010,N_3002);
xor U6216 (N_6216,N_3756,N_2606);
and U6217 (N_6217,N_3647,N_136);
and U6218 (N_6218,N_1346,N_2589);
nor U6219 (N_6219,N_1582,N_2447);
nor U6220 (N_6220,N_1300,N_4228);
nor U6221 (N_6221,N_2571,N_714);
and U6222 (N_6222,N_3611,N_4585);
and U6223 (N_6223,N_552,N_649);
and U6224 (N_6224,N_2858,N_1155);
or U6225 (N_6225,N_56,N_2409);
or U6226 (N_6226,N_65,N_1890);
xnor U6227 (N_6227,N_4571,N_3910);
xor U6228 (N_6228,N_3561,N_3106);
nor U6229 (N_6229,N_2548,N_4062);
or U6230 (N_6230,N_2411,N_1937);
xor U6231 (N_6231,N_3652,N_2053);
xnor U6232 (N_6232,N_3583,N_921);
nor U6233 (N_6233,N_2691,N_719);
and U6234 (N_6234,N_2558,N_2075);
or U6235 (N_6235,N_1715,N_1514);
and U6236 (N_6236,N_3563,N_2655);
or U6237 (N_6237,N_3781,N_1528);
nand U6238 (N_6238,N_4998,N_4904);
nor U6239 (N_6239,N_2094,N_3725);
and U6240 (N_6240,N_2299,N_925);
and U6241 (N_6241,N_4622,N_3707);
xor U6242 (N_6242,N_4943,N_2773);
or U6243 (N_6243,N_3246,N_2862);
nand U6244 (N_6244,N_3670,N_2565);
and U6245 (N_6245,N_4596,N_3395);
or U6246 (N_6246,N_927,N_863);
and U6247 (N_6247,N_4475,N_4465);
nand U6248 (N_6248,N_458,N_2652);
or U6249 (N_6249,N_4068,N_1233);
nor U6250 (N_6250,N_2344,N_4828);
and U6251 (N_6251,N_1940,N_3175);
or U6252 (N_6252,N_4788,N_2335);
nand U6253 (N_6253,N_2897,N_3264);
nor U6254 (N_6254,N_22,N_1892);
nor U6255 (N_6255,N_685,N_4484);
xnor U6256 (N_6256,N_1815,N_981);
nor U6257 (N_6257,N_69,N_4021);
xnor U6258 (N_6258,N_294,N_4186);
and U6259 (N_6259,N_553,N_4869);
or U6260 (N_6260,N_249,N_4999);
or U6261 (N_6261,N_4493,N_2101);
and U6262 (N_6262,N_339,N_1289);
and U6263 (N_6263,N_1383,N_4499);
or U6264 (N_6264,N_1467,N_4285);
nor U6265 (N_6265,N_4810,N_4898);
xnor U6266 (N_6266,N_2965,N_753);
xor U6267 (N_6267,N_1951,N_1313);
nor U6268 (N_6268,N_4527,N_1101);
xnor U6269 (N_6269,N_2031,N_166);
and U6270 (N_6270,N_4370,N_3599);
and U6271 (N_6271,N_2776,N_1336);
or U6272 (N_6272,N_3016,N_2476);
or U6273 (N_6273,N_1021,N_656);
and U6274 (N_6274,N_1092,N_150);
nor U6275 (N_6275,N_868,N_4915);
or U6276 (N_6276,N_2475,N_993);
or U6277 (N_6277,N_3554,N_1671);
nor U6278 (N_6278,N_4075,N_2519);
and U6279 (N_6279,N_3792,N_4142);
nor U6280 (N_6280,N_3075,N_121);
xnor U6281 (N_6281,N_834,N_1083);
nand U6282 (N_6282,N_3767,N_4386);
nand U6283 (N_6283,N_523,N_3489);
xnor U6284 (N_6284,N_2978,N_3200);
nor U6285 (N_6285,N_73,N_893);
nor U6286 (N_6286,N_252,N_1109);
nor U6287 (N_6287,N_4415,N_2684);
or U6288 (N_6288,N_4703,N_1133);
nand U6289 (N_6289,N_1286,N_1274);
nor U6290 (N_6290,N_3627,N_572);
xor U6291 (N_6291,N_1329,N_232);
nand U6292 (N_6292,N_2728,N_4437);
and U6293 (N_6293,N_258,N_992);
and U6294 (N_6294,N_519,N_403);
xor U6295 (N_6295,N_3956,N_3226);
nor U6296 (N_6296,N_4348,N_2089);
or U6297 (N_6297,N_2959,N_3584);
or U6298 (N_6298,N_1755,N_4422);
and U6299 (N_6299,N_3527,N_1600);
xor U6300 (N_6300,N_3348,N_4811);
nand U6301 (N_6301,N_4269,N_2074);
nor U6302 (N_6302,N_2013,N_3499);
nor U6303 (N_6303,N_3929,N_2380);
xnor U6304 (N_6304,N_3407,N_4209);
and U6305 (N_6305,N_1430,N_3178);
nand U6306 (N_6306,N_1452,N_4634);
xnor U6307 (N_6307,N_3660,N_1375);
nand U6308 (N_6308,N_2017,N_4889);
nor U6309 (N_6309,N_3194,N_398);
nand U6310 (N_6310,N_4158,N_1240);
and U6311 (N_6311,N_4018,N_1428);
or U6312 (N_6312,N_2166,N_1450);
and U6313 (N_6313,N_2633,N_3620);
and U6314 (N_6314,N_2413,N_606);
nand U6315 (N_6315,N_1093,N_2363);
and U6316 (N_6316,N_2906,N_4461);
nand U6317 (N_6317,N_3664,N_330);
xor U6318 (N_6318,N_4706,N_1165);
xnor U6319 (N_6319,N_80,N_1388);
nor U6320 (N_6320,N_797,N_4534);
xnor U6321 (N_6321,N_3609,N_514);
and U6322 (N_6322,N_829,N_1110);
nor U6323 (N_6323,N_3269,N_488);
nand U6324 (N_6324,N_2760,N_3238);
or U6325 (N_6325,N_4801,N_1030);
nor U6326 (N_6326,N_1005,N_3484);
and U6327 (N_6327,N_1113,N_3190);
nand U6328 (N_6328,N_1393,N_1178);
nor U6329 (N_6329,N_2135,N_220);
nor U6330 (N_6330,N_4840,N_3078);
nand U6331 (N_6331,N_1024,N_2376);
and U6332 (N_6332,N_424,N_4765);
nor U6333 (N_6333,N_91,N_3631);
nand U6334 (N_6334,N_4664,N_92);
and U6335 (N_6335,N_3227,N_2038);
and U6336 (N_6336,N_1080,N_3676);
nor U6337 (N_6337,N_4488,N_3799);
xor U6338 (N_6338,N_569,N_4164);
nor U6339 (N_6339,N_3874,N_4311);
nand U6340 (N_6340,N_3549,N_1643);
and U6341 (N_6341,N_1261,N_4327);
and U6342 (N_6342,N_4303,N_3223);
and U6343 (N_6343,N_317,N_748);
or U6344 (N_6344,N_3454,N_2177);
nand U6345 (N_6345,N_2758,N_4957);
nor U6346 (N_6346,N_4392,N_327);
xor U6347 (N_6347,N_351,N_2127);
nor U6348 (N_6348,N_1998,N_3263);
or U6349 (N_6349,N_3977,N_1660);
and U6350 (N_6350,N_2062,N_2131);
and U6351 (N_6351,N_2626,N_236);
nor U6352 (N_6352,N_271,N_630);
nor U6353 (N_6353,N_3532,N_3542);
xnor U6354 (N_6354,N_4696,N_7);
nor U6355 (N_6355,N_4603,N_3905);
nor U6356 (N_6356,N_3034,N_4098);
or U6357 (N_6357,N_1939,N_2999);
nor U6358 (N_6358,N_1799,N_4466);
and U6359 (N_6359,N_725,N_1608);
and U6360 (N_6360,N_778,N_380);
and U6361 (N_6361,N_2910,N_3437);
nand U6362 (N_6362,N_4620,N_4643);
nor U6363 (N_6363,N_3568,N_3212);
nor U6364 (N_6364,N_4205,N_292);
and U6365 (N_6365,N_3029,N_385);
and U6366 (N_6366,N_673,N_3347);
or U6367 (N_6367,N_872,N_2761);
and U6368 (N_6368,N_2549,N_3593);
or U6369 (N_6369,N_467,N_4970);
or U6370 (N_6370,N_2526,N_2832);
nand U6371 (N_6371,N_2663,N_3103);
and U6372 (N_6372,N_3099,N_4153);
and U6373 (N_6373,N_2752,N_694);
or U6374 (N_6374,N_3878,N_2903);
nor U6375 (N_6375,N_4613,N_2224);
and U6376 (N_6376,N_3759,N_4682);
and U6377 (N_6377,N_3838,N_1757);
and U6378 (N_6378,N_2086,N_2966);
or U6379 (N_6379,N_2000,N_2402);
nand U6380 (N_6380,N_3649,N_780);
nor U6381 (N_6381,N_3126,N_1032);
nand U6382 (N_6382,N_3124,N_3265);
and U6383 (N_6383,N_2156,N_4961);
nand U6384 (N_6384,N_4352,N_4472);
nand U6385 (N_6385,N_4185,N_1327);
nand U6386 (N_6386,N_929,N_4750);
and U6387 (N_6387,N_2345,N_2244);
or U6388 (N_6388,N_244,N_1887);
and U6389 (N_6389,N_2676,N_431);
or U6390 (N_6390,N_4517,N_627);
or U6391 (N_6391,N_731,N_1529);
or U6392 (N_6392,N_1955,N_2662);
nor U6393 (N_6393,N_1502,N_3142);
nor U6394 (N_6394,N_1629,N_2725);
nand U6395 (N_6395,N_4490,N_2683);
and U6396 (N_6396,N_3132,N_2557);
and U6397 (N_6397,N_967,N_2829);
or U6398 (N_6398,N_2203,N_1598);
nand U6399 (N_6399,N_430,N_2263);
or U6400 (N_6400,N_1205,N_4790);
and U6401 (N_6401,N_3880,N_4433);
or U6402 (N_6402,N_1710,N_3716);
and U6403 (N_6403,N_1571,N_4350);
nor U6404 (N_6404,N_1949,N_494);
nand U6405 (N_6405,N_728,N_340);
xor U6406 (N_6406,N_4305,N_4219);
nand U6407 (N_6407,N_3242,N_3176);
nor U6408 (N_6408,N_460,N_636);
or U6409 (N_6409,N_989,N_1088);
or U6410 (N_6410,N_2261,N_4871);
and U6411 (N_6411,N_4019,N_4700);
xor U6412 (N_6412,N_2306,N_3566);
xnor U6413 (N_6413,N_2543,N_641);
and U6414 (N_6414,N_4740,N_2779);
nand U6415 (N_6415,N_117,N_2349);
or U6416 (N_6416,N_1682,N_1183);
and U6417 (N_6417,N_2005,N_2061);
nor U6418 (N_6418,N_4980,N_357);
xnor U6419 (N_6419,N_535,N_4184);
nand U6420 (N_6420,N_1214,N_3072);
and U6421 (N_6421,N_1479,N_3113);
or U6422 (N_6422,N_3382,N_3439);
or U6423 (N_6423,N_52,N_784);
or U6424 (N_6424,N_1546,N_1177);
nor U6425 (N_6425,N_1077,N_49);
xnor U6426 (N_6426,N_1675,N_4486);
nor U6427 (N_6427,N_3109,N_3953);
or U6428 (N_6428,N_4298,N_1894);
and U6429 (N_6429,N_976,N_169);
and U6430 (N_6430,N_2899,N_2562);
and U6431 (N_6431,N_18,N_2348);
nand U6432 (N_6432,N_1017,N_2509);
and U6433 (N_6433,N_1689,N_4003);
xnor U6434 (N_6434,N_251,N_3550);
or U6435 (N_6435,N_894,N_2185);
nor U6436 (N_6436,N_1773,N_2576);
nor U6437 (N_6437,N_4263,N_1752);
or U6438 (N_6438,N_2206,N_4042);
or U6439 (N_6439,N_4084,N_4624);
or U6440 (N_6440,N_1867,N_1025);
nor U6441 (N_6441,N_2477,N_2505);
xnor U6442 (N_6442,N_3802,N_1406);
and U6443 (N_6443,N_1149,N_770);
nand U6444 (N_6444,N_3843,N_287);
nand U6445 (N_6445,N_4045,N_1471);
nor U6446 (N_6446,N_454,N_4283);
nand U6447 (N_6447,N_3850,N_194);
and U6448 (N_6448,N_400,N_1647);
nor U6449 (N_6449,N_879,N_798);
nor U6450 (N_6450,N_1033,N_3396);
nor U6451 (N_6451,N_3185,N_374);
or U6452 (N_6452,N_4377,N_1372);
nand U6453 (N_6453,N_4255,N_4453);
nor U6454 (N_6454,N_1160,N_4016);
or U6455 (N_6455,N_1425,N_262);
nand U6456 (N_6456,N_4256,N_3961);
nand U6457 (N_6457,N_1936,N_954);
nand U6458 (N_6458,N_2460,N_4660);
and U6459 (N_6459,N_3903,N_2015);
or U6460 (N_6460,N_4586,N_793);
nand U6461 (N_6461,N_167,N_688);
and U6462 (N_6462,N_1980,N_2785);
and U6463 (N_6463,N_4196,N_3286);
nor U6464 (N_6464,N_2736,N_4649);
or U6465 (N_6465,N_2430,N_3054);
and U6466 (N_6466,N_1151,N_977);
xnor U6467 (N_6467,N_707,N_2296);
and U6468 (N_6468,N_2572,N_1338);
or U6469 (N_6469,N_1499,N_799);
and U6470 (N_6470,N_1718,N_3149);
and U6471 (N_6471,N_2356,N_1969);
nor U6472 (N_6472,N_1501,N_1491);
and U6473 (N_6473,N_3712,N_1228);
or U6474 (N_6474,N_2879,N_45);
and U6475 (N_6475,N_2820,N_3943);
nor U6476 (N_6476,N_2955,N_2186);
nand U6477 (N_6477,N_2008,N_2321);
and U6478 (N_6478,N_1438,N_1896);
and U6479 (N_6479,N_3777,N_4697);
or U6480 (N_6480,N_3703,N_238);
and U6481 (N_6481,N_2794,N_3890);
nand U6482 (N_6482,N_1474,N_3294);
or U6483 (N_6483,N_2918,N_3241);
nand U6484 (N_6484,N_4959,N_3590);
nand U6485 (N_6485,N_1919,N_2457);
or U6486 (N_6486,N_306,N_2609);
nor U6487 (N_6487,N_3193,N_1704);
or U6488 (N_6488,N_4267,N_3697);
nand U6489 (N_6489,N_3894,N_4161);
nand U6490 (N_6490,N_4381,N_4458);
nand U6491 (N_6491,N_3107,N_1314);
and U6492 (N_6492,N_186,N_4884);
nand U6493 (N_6493,N_3893,N_2178);
nand U6494 (N_6494,N_3704,N_3460);
and U6495 (N_6495,N_3744,N_3667);
nor U6496 (N_6496,N_4655,N_1042);
nor U6497 (N_6497,N_4673,N_2644);
nor U6498 (N_6498,N_2289,N_1384);
and U6499 (N_6499,N_455,N_937);
nand U6500 (N_6500,N_120,N_2143);
nor U6501 (N_6501,N_4133,N_4587);
nand U6502 (N_6502,N_3559,N_947);
nor U6503 (N_6503,N_257,N_2551);
and U6504 (N_6504,N_1159,N_850);
nor U6505 (N_6505,N_3234,N_1738);
and U6506 (N_6506,N_3302,N_1591);
and U6507 (N_6507,N_2658,N_768);
nor U6508 (N_6508,N_1029,N_3411);
or U6509 (N_6509,N_111,N_1065);
xnor U6510 (N_6510,N_2032,N_4470);
nor U6511 (N_6511,N_412,N_4691);
or U6512 (N_6512,N_2401,N_861);
or U6513 (N_6513,N_3165,N_4979);
and U6514 (N_6514,N_2351,N_2084);
xnor U6515 (N_6515,N_3636,N_2141);
or U6516 (N_6516,N_2164,N_3278);
xor U6517 (N_6517,N_4911,N_4468);
or U6518 (N_6518,N_3051,N_2240);
or U6519 (N_6519,N_3139,N_1377);
and U6520 (N_6520,N_4882,N_2817);
or U6521 (N_6521,N_4273,N_3524);
and U6522 (N_6522,N_2091,N_4906);
nor U6523 (N_6523,N_2822,N_1617);
and U6524 (N_6524,N_2671,N_2941);
nor U6525 (N_6525,N_2030,N_219);
xor U6526 (N_6526,N_4174,N_4759);
or U6527 (N_6527,N_4598,N_4102);
and U6528 (N_6528,N_359,N_3470);
nand U6529 (N_6529,N_3779,N_4171);
nor U6530 (N_6530,N_3936,N_105);
nand U6531 (N_6531,N_4439,N_2346);
nand U6532 (N_6532,N_2542,N_3600);
nand U6533 (N_6533,N_4688,N_3811);
and U6534 (N_6534,N_2023,N_3680);
nor U6535 (N_6535,N_225,N_1594);
or U6536 (N_6536,N_2382,N_3927);
nand U6537 (N_6537,N_2749,N_1526);
and U6538 (N_6538,N_1732,N_3606);
and U6539 (N_6539,N_677,N_2711);
or U6540 (N_6540,N_3475,N_4552);
and U6541 (N_6541,N_240,N_783);
and U6542 (N_6542,N_4608,N_1683);
nor U6543 (N_6543,N_3478,N_1168);
and U6544 (N_6544,N_2613,N_3364);
nand U6545 (N_6545,N_1413,N_1117);
nor U6546 (N_6546,N_542,N_3930);
nand U6547 (N_6547,N_1843,N_1844);
nor U6548 (N_6548,N_1914,N_2642);
xnor U6549 (N_6549,N_4405,N_3809);
nor U6550 (N_6550,N_3958,N_594);
and U6551 (N_6551,N_2740,N_2331);
nand U6552 (N_6552,N_2598,N_2069);
nand U6553 (N_6553,N_2948,N_4541);
nor U6554 (N_6554,N_2871,N_1719);
nand U6555 (N_6555,N_2917,N_1123);
or U6556 (N_6556,N_371,N_3657);
nand U6557 (N_6557,N_1592,N_4175);
nand U6558 (N_6558,N_1648,N_4165);
and U6559 (N_6559,N_4373,N_1863);
and U6560 (N_6560,N_2984,N_858);
xor U6561 (N_6561,N_4723,N_3280);
and U6562 (N_6562,N_170,N_3970);
or U6563 (N_6563,N_2040,N_4190);
nor U6564 (N_6564,N_4795,N_1038);
and U6565 (N_6565,N_3668,N_4446);
nor U6566 (N_6566,N_3462,N_4147);
nor U6567 (N_6567,N_4320,N_4399);
and U6568 (N_6568,N_3086,N_1136);
xnor U6569 (N_6569,N_1563,N_3775);
or U6570 (N_6570,N_4413,N_2863);
nand U6571 (N_6571,N_1497,N_1520);
nand U6572 (N_6572,N_2680,N_2278);
and U6573 (N_6573,N_1237,N_659);
or U6574 (N_6574,N_3529,N_4435);
and U6575 (N_6575,N_1877,N_4398);
and U6576 (N_6576,N_2472,N_1409);
nand U6577 (N_6577,N_129,N_1106);
nand U6578 (N_6578,N_1763,N_4429);
or U6579 (N_6579,N_2912,N_3066);
nor U6580 (N_6580,N_1339,N_2668);
nor U6581 (N_6581,N_4491,N_3069);
nor U6582 (N_6582,N_3520,N_4963);
or U6583 (N_6583,N_1063,N_4504);
nand U6584 (N_6584,N_3509,N_4808);
nor U6585 (N_6585,N_4215,N_4823);
or U6586 (N_6586,N_3739,N_1045);
and U6587 (N_6587,N_3753,N_1054);
nand U6588 (N_6588,N_1836,N_2819);
and U6589 (N_6589,N_88,N_4849);
xnor U6590 (N_6590,N_4802,N_2495);
nand U6591 (N_6591,N_201,N_2866);
nand U6592 (N_6592,N_4711,N_3666);
nand U6593 (N_6593,N_3184,N_3421);
or U6594 (N_6594,N_4451,N_3093);
or U6595 (N_6595,N_1701,N_46);
nor U6596 (N_6596,N_4191,N_1532);
or U6597 (N_6597,N_2612,N_895);
or U6598 (N_6598,N_1809,N_1699);
nand U6599 (N_6599,N_4720,N_4665);
or U6600 (N_6600,N_122,N_115);
nor U6601 (N_6601,N_2954,N_1693);
and U6602 (N_6602,N_3358,N_1906);
or U6603 (N_6603,N_148,N_3873);
or U6604 (N_6604,N_2142,N_2979);
or U6605 (N_6605,N_642,N_2578);
and U6606 (N_6606,N_1432,N_1517);
xnor U6607 (N_6607,N_1373,N_3137);
nor U6608 (N_6608,N_815,N_1846);
nand U6609 (N_6609,N_540,N_2427);
xnor U6610 (N_6610,N_3999,N_47);
nand U6611 (N_6611,N_2359,N_2225);
and U6612 (N_6612,N_2180,N_847);
or U6613 (N_6613,N_1069,N_1078);
nor U6614 (N_6614,N_3151,N_1164);
and U6615 (N_6615,N_3373,N_3526);
nand U6616 (N_6616,N_461,N_4257);
nand U6617 (N_6617,N_1347,N_3172);
nand U6618 (N_6618,N_4617,N_2600);
and U6619 (N_6619,N_3863,N_4651);
nand U6620 (N_6620,N_3434,N_520);
and U6621 (N_6621,N_2478,N_1776);
and U6622 (N_6622,N_3856,N_3245);
xor U6623 (N_6623,N_1512,N_2649);
or U6624 (N_6624,N_346,N_1540);
or U6625 (N_6625,N_2645,N_1360);
and U6626 (N_6626,N_2446,N_3998);
xnor U6627 (N_6627,N_1280,N_214);
nand U6628 (N_6628,N_4421,N_74);
and U6629 (N_6629,N_2667,N_267);
nand U6630 (N_6630,N_860,N_2808);
or U6631 (N_6631,N_3216,N_68);
nand U6632 (N_6632,N_1518,N_333);
nand U6633 (N_6633,N_1511,N_2914);
and U6634 (N_6634,N_4826,N_3686);
nand U6635 (N_6635,N_3077,N_1961);
xor U6636 (N_6636,N_4419,N_3562);
or U6637 (N_6637,N_3928,N_44);
and U6638 (N_6638,N_2220,N_2383);
nor U6639 (N_6639,N_1464,N_4530);
nand U6640 (N_6640,N_1953,N_4156);
or U6641 (N_6641,N_563,N_345);
and U6642 (N_6642,N_1330,N_1692);
and U6643 (N_6643,N_2793,N_1253);
nor U6644 (N_6644,N_771,N_3498);
or U6645 (N_6645,N_1488,N_3455);
nor U6646 (N_6646,N_1932,N_14);
nand U6647 (N_6647,N_1334,N_2620);
nand U6648 (N_6648,N_4852,N_2601);
or U6649 (N_6649,N_2103,N_3808);
nor U6650 (N_6650,N_598,N_138);
nand U6651 (N_6651,N_3472,N_4536);
nand U6652 (N_6652,N_3189,N_4216);
nor U6653 (N_6653,N_4020,N_4159);
or U6654 (N_6654,N_807,N_846);
nand U6655 (N_6655,N_2277,N_1433);
xnor U6656 (N_6656,N_603,N_2404);
and U6657 (N_6657,N_4286,N_1304);
nand U6658 (N_6658,N_4880,N_4059);
and U6659 (N_6659,N_4026,N_3469);
and U6660 (N_6660,N_4814,N_3131);
nor U6661 (N_6661,N_181,N_1587);
nand U6662 (N_6662,N_1606,N_4245);
and U6663 (N_6663,N_1577,N_1916);
and U6664 (N_6664,N_4418,N_2397);
xor U6665 (N_6665,N_2390,N_2473);
or U6666 (N_6666,N_4331,N_3156);
or U6667 (N_6667,N_4217,N_3446);
nand U6668 (N_6668,N_3984,N_4351);
and U6669 (N_6669,N_1521,N_2936);
nor U6670 (N_6670,N_2384,N_1048);
xnor U6671 (N_6671,N_4769,N_2255);
nor U6672 (N_6672,N_2260,N_304);
xor U6673 (N_6673,N_845,N_2286);
nor U6674 (N_6674,N_2919,N_3435);
nand U6675 (N_6675,N_2533,N_1365);
nor U6676 (N_6676,N_1611,N_3070);
nor U6677 (N_6677,N_835,N_2986);
or U6678 (N_6678,N_2988,N_2782);
and U6679 (N_6679,N_3495,N_2857);
nor U6680 (N_6680,N_4789,N_871);
xnor U6681 (N_6681,N_2388,N_3191);
xor U6682 (N_6682,N_761,N_4886);
nand U6683 (N_6683,N_2279,N_4839);
nor U6684 (N_6684,N_3849,N_3949);
and U6685 (N_6685,N_4332,N_10);
nor U6686 (N_6686,N_1026,N_1785);
nand U6687 (N_6687,N_3297,N_3387);
nand U6688 (N_6688,N_2315,N_2846);
nor U6689 (N_6689,N_2774,N_1236);
nand U6690 (N_6690,N_3948,N_4044);
and U6691 (N_6691,N_1331,N_3920);
nand U6692 (N_6692,N_1218,N_3805);
and U6693 (N_6693,N_63,N_2992);
nand U6694 (N_6694,N_3497,N_733);
nor U6695 (N_6695,N_2825,N_1728);
nand U6696 (N_6696,N_1636,N_2403);
and U6697 (N_6697,N_2770,N_1834);
and U6698 (N_6698,N_3325,N_4717);
nand U6699 (N_6699,N_1811,N_2108);
and U6700 (N_6700,N_4575,N_1281);
nand U6701 (N_6701,N_432,N_1394);
nor U6702 (N_6702,N_4804,N_3214);
nor U6703 (N_6703,N_3219,N_582);
or U6704 (N_6704,N_3047,N_4786);
nor U6705 (N_6705,N_1271,N_994);
nand U6706 (N_6706,N_21,N_754);
and U6707 (N_6707,N_477,N_3687);
and U6708 (N_6708,N_4991,N_4679);
xnor U6709 (N_6709,N_2422,N_4130);
nand U6710 (N_6710,N_399,N_2705);
nand U6711 (N_6711,N_2066,N_4281);
and U6712 (N_6712,N_1792,N_987);
and U6713 (N_6713,N_3243,N_1419);
or U6714 (N_6714,N_828,N_794);
and U6715 (N_6715,N_1560,N_1967);
or U6716 (N_6716,N_4139,N_230);
nand U6717 (N_6717,N_1420,N_3160);
or U6718 (N_6718,N_2334,N_4783);
nor U6719 (N_6719,N_2501,N_2651);
nor U6720 (N_6720,N_1267,N_2995);
nand U6721 (N_6721,N_388,N_118);
nor U6722 (N_6722,N_591,N_4438);
and U6723 (N_6723,N_4853,N_501);
nand U6724 (N_6724,N_423,N_4807);
and U6725 (N_6725,N_2452,N_4763);
nor U6726 (N_6726,N_4065,N_1695);
nor U6727 (N_6727,N_4454,N_1651);
nor U6728 (N_6728,N_1197,N_4009);
nor U6729 (N_6729,N_4412,N_3968);
and U6730 (N_6730,N_1735,N_1850);
xnor U6731 (N_6731,N_375,N_4432);
and U6732 (N_6732,N_4054,N_1154);
xnor U6733 (N_6733,N_1926,N_4654);
nand U6734 (N_6734,N_3237,N_1909);
nor U6735 (N_6735,N_3769,N_2440);
or U6736 (N_6736,N_2090,N_3367);
xnor U6737 (N_6737,N_474,N_4710);
or U6738 (N_6738,N_3872,N_483);
nand U6739 (N_6739,N_4199,N_2050);
xnor U6740 (N_6740,N_644,N_4455);
or U6741 (N_6741,N_1705,N_1245);
or U6742 (N_6742,N_3027,N_710);
and U6743 (N_6743,N_290,N_2318);
nor U6744 (N_6744,N_4040,N_3221);
or U6745 (N_6745,N_1366,N_4580);
and U6746 (N_6746,N_568,N_4310);
or U6747 (N_6747,N_1848,N_1351);
nand U6748 (N_6748,N_3171,N_1158);
or U6749 (N_6749,N_896,N_3803);
or U6750 (N_6750,N_511,N_2925);
and U6751 (N_6751,N_1162,N_4876);
nor U6752 (N_6752,N_2387,N_2675);
nand U6753 (N_6753,N_363,N_4374);
xnor U6754 (N_6754,N_1252,N_4093);
nand U6755 (N_6755,N_543,N_2226);
nand U6756 (N_6756,N_4546,N_1361);
or U6757 (N_6757,N_585,N_866);
or U6758 (N_6758,N_2653,N_746);
xnor U6759 (N_6759,N_4086,N_2288);
nor U6760 (N_6760,N_1508,N_2608);
nor U6761 (N_6761,N_655,N_95);
and U6762 (N_6762,N_261,N_2970);
and U6763 (N_6763,N_3728,N_1891);
nor U6764 (N_6764,N_1677,N_1120);
and U6765 (N_6765,N_2118,N_4082);
nor U6766 (N_6766,N_1562,N_1986);
nand U6767 (N_6767,N_1678,N_882);
or U6768 (N_6768,N_4842,N_2518);
and U6769 (N_6769,N_464,N_4090);
xor U6770 (N_6770,N_2124,N_130);
nand U6771 (N_6771,N_1788,N_4111);
and U6772 (N_6772,N_4070,N_3963);
nand U6773 (N_6773,N_3909,N_4730);
and U6774 (N_6774,N_3814,N_2837);
nand U6775 (N_6775,N_1535,N_3021);
or U6776 (N_6776,N_3284,N_1830);
nor U6777 (N_6777,N_2110,N_1309);
or U6778 (N_6778,N_191,N_1448);
nor U6779 (N_6779,N_4838,N_2748);
nor U6780 (N_6780,N_2672,N_2859);
nand U6781 (N_6781,N_980,N_2341);
nand U6782 (N_6782,N_4200,N_3748);
nor U6783 (N_6783,N_1405,N_1121);
or U6784 (N_6784,N_3377,N_2235);
and U6785 (N_6785,N_1002,N_4477);
and U6786 (N_6786,N_3812,N_3006);
and U6787 (N_6787,N_3017,N_2891);
nand U6788 (N_6788,N_566,N_2046);
xnor U6789 (N_6789,N_2237,N_1439);
xor U6790 (N_6790,N_1820,N_910);
nand U6791 (N_6791,N_1473,N_1322);
nor U6792 (N_6792,N_4555,N_2874);
or U6793 (N_6793,N_3152,N_4916);
and U6794 (N_6794,N_1249,N_4827);
and U6795 (N_6795,N_545,N_1670);
or U6796 (N_6796,N_4646,N_1744);
and U6797 (N_6797,N_2900,N_158);
or U6798 (N_6798,N_1851,N_4687);
nand U6799 (N_6799,N_4246,N_1552);
xnor U6800 (N_6800,N_350,N_580);
or U6801 (N_6801,N_718,N_4675);
or U6802 (N_6802,N_4410,N_2311);
or U6803 (N_6803,N_128,N_2421);
nor U6804 (N_6804,N_2887,N_4521);
and U6805 (N_6805,N_2732,N_3162);
or U6806 (N_6806,N_3037,N_558);
nor U6807 (N_6807,N_716,N_609);
and U6808 (N_6808,N_2470,N_1640);
nand U6809 (N_6809,N_2439,N_54);
and U6810 (N_6810,N_2810,N_3705);
nor U6811 (N_6811,N_4896,N_735);
or U6812 (N_6812,N_4778,N_870);
and U6813 (N_6813,N_1991,N_2239);
or U6814 (N_6814,N_444,N_1039);
nand U6815 (N_6815,N_3202,N_4982);
or U6816 (N_6816,N_4449,N_3060);
and U6817 (N_6817,N_779,N_4535);
nand U6818 (N_6818,N_950,N_3306);
nor U6819 (N_6819,N_4402,N_1316);
or U6820 (N_6820,N_3907,N_1604);
and U6821 (N_6821,N_3654,N_3400);
nor U6822 (N_6822,N_1872,N_1062);
and U6823 (N_6823,N_1470,N_4264);
nand U6824 (N_6824,N_3742,N_3491);
nand U6825 (N_6825,N_2585,N_4201);
nor U6826 (N_6826,N_4479,N_2104);
or U6827 (N_6827,N_2073,N_1810);
xnor U6828 (N_6828,N_3092,N_3074);
and U6829 (N_6829,N_1970,N_1193);
and U6830 (N_6830,N_4301,N_4567);
nand U6831 (N_6831,N_4938,N_4662);
nor U6832 (N_6832,N_2991,N_1956);
nand U6833 (N_6833,N_934,N_314);
nand U6834 (N_6834,N_3588,N_1821);
and U6835 (N_6835,N_2835,N_4498);
or U6836 (N_6836,N_1086,N_1091);
nand U6837 (N_6837,N_3168,N_3385);
nand U6838 (N_6838,N_4467,N_1416);
nand U6839 (N_6839,N_1579,N_1632);
and U6840 (N_6840,N_3150,N_1451);
and U6841 (N_6841,N_4239,N_4304);
xnor U6842 (N_6842,N_2416,N_4483);
nand U6843 (N_6843,N_2398,N_2058);
nor U6844 (N_6844,N_767,N_4845);
and U6845 (N_6845,N_2293,N_801);
nand U6846 (N_6846,N_2368,N_3067);
or U6847 (N_6847,N_3825,N_3790);
nand U6848 (N_6848,N_1429,N_3381);
nand U6849 (N_6849,N_900,N_4724);
nor U6850 (N_6850,N_4095,N_2905);
nand U6851 (N_6851,N_2973,N_2719);
nor U6852 (N_6852,N_2148,N_534);
nand U6853 (N_6853,N_3135,N_722);
and U6854 (N_6854,N_3427,N_2175);
and U6855 (N_6855,N_4376,N_4625);
or U6856 (N_6856,N_1251,N_4248);
nor U6857 (N_6857,N_851,N_959);
nor U6858 (N_6858,N_413,N_3675);
or U6859 (N_6859,N_427,N_3282);
nor U6860 (N_6860,N_4747,N_2730);
nor U6861 (N_6861,N_2994,N_2746);
and U6862 (N_6862,N_3406,N_2436);
nand U6863 (N_6863,N_1853,N_661);
nand U6864 (N_6864,N_4992,N_316);
nor U6865 (N_6865,N_2098,N_1596);
xnor U6866 (N_6866,N_3923,N_3088);
nand U6867 (N_6867,N_2630,N_811);
nor U6868 (N_6868,N_2002,N_1047);
xor U6869 (N_6869,N_4883,N_2716);
and U6870 (N_6870,N_35,N_3213);
nand U6871 (N_6871,N_4480,N_4112);
nor U6872 (N_6872,N_3244,N_1665);
or U6873 (N_6873,N_2269,N_243);
nand U6874 (N_6874,N_2087,N_4343);
nor U6875 (N_6875,N_3951,N_2795);
nor U6876 (N_6876,N_883,N_3161);
nand U6877 (N_6877,N_1607,N_743);
nor U6878 (N_6878,N_3310,N_2479);
nor U6879 (N_6879,N_2763,N_2197);
nand U6880 (N_6880,N_612,N_1036);
nor U6881 (N_6881,N_1179,N_3115);
or U6882 (N_6882,N_1658,N_1555);
nor U6883 (N_6883,N_3118,N_3741);
or U6884 (N_6884,N_4028,N_3614);
and U6885 (N_6885,N_2849,N_940);
nor U6886 (N_6886,N_3296,N_1207);
or U6887 (N_6887,N_2961,N_2302);
xnor U6888 (N_6888,N_775,N_2714);
nor U6889 (N_6889,N_2025,N_1885);
and U6890 (N_6890,N_2047,N_676);
nor U6891 (N_6891,N_4481,N_2860);
nand U6892 (N_6892,N_1349,N_4725);
nand U6893 (N_6893,N_1079,N_4964);
xor U6894 (N_6894,N_2125,N_919);
nand U6895 (N_6895,N_2902,N_132);
and U6896 (N_6896,N_2974,N_3330);
and U6897 (N_6897,N_3674,N_1898);
nor U6898 (N_6898,N_4771,N_1999);
xnor U6899 (N_6899,N_1868,N_484);
nor U6900 (N_6900,N_720,N_397);
xor U6901 (N_6901,N_3179,N_741);
nor U6902 (N_6902,N_602,N_3459);
or U6903 (N_6903,N_4474,N_2657);
nor U6904 (N_6904,N_4927,N_805);
and U6905 (N_6905,N_1073,N_4513);
and U6906 (N_6906,N_3312,N_848);
and U6907 (N_6907,N_4822,N_4683);
and U6908 (N_6908,N_593,N_1306);
nor U6909 (N_6909,N_217,N_3267);
nor U6910 (N_6910,N_756,N_2365);
or U6911 (N_6911,N_1963,N_3592);
nand U6912 (N_6912,N_4357,N_2845);
nor U6913 (N_6913,N_110,N_1490);
or U6914 (N_6914,N_4742,N_4867);
nand U6915 (N_6915,N_1020,N_2056);
nand U6916 (N_6916,N_1321,N_2034);
nand U6917 (N_6917,N_2232,N_1988);
and U6918 (N_6918,N_4549,N_2412);
nand U6919 (N_6919,N_4516,N_1234);
and U6920 (N_6920,N_365,N_13);
or U6921 (N_6921,N_3170,N_3031);
nor U6922 (N_6922,N_358,N_663);
and U6923 (N_6923,N_4072,N_4794);
nor U6924 (N_6924,N_103,N_434);
and U6925 (N_6925,N_1220,N_3774);
xor U6926 (N_6926,N_4936,N_1056);
or U6927 (N_6927,N_4727,N_3589);
and U6928 (N_6928,N_4365,N_3714);
or U6929 (N_6929,N_615,N_2544);
xnor U6930 (N_6930,N_2828,N_3163);
nor U6931 (N_6931,N_3220,N_3991);
nor U6932 (N_6932,N_3831,N_2136);
and U6933 (N_6933,N_4225,N_1513);
and U6934 (N_6934,N_235,N_3860);
or U6935 (N_6935,N_196,N_200);
nor U6936 (N_6936,N_4818,N_2396);
or U6937 (N_6937,N_4080,N_2976);
nor U6938 (N_6938,N_827,N_4107);
nand U6939 (N_6939,N_3276,N_928);
nand U6940 (N_6940,N_480,N_772);
or U6941 (N_6941,N_1299,N_2193);
or U6942 (N_6942,N_1108,N_348);
nand U6943 (N_6943,N_3403,N_4113);
nand U6944 (N_6944,N_1921,N_2679);
or U6945 (N_6945,N_1605,N_1486);
nand U6946 (N_6946,N_1567,N_2507);
and U6947 (N_6947,N_4456,N_447);
or U6948 (N_6948,N_32,N_2826);
or U6949 (N_6949,N_2271,N_1046);
or U6950 (N_6950,N_3558,N_1800);
and U6951 (N_6951,N_2935,N_2219);
nand U6952 (N_6952,N_2123,N_1784);
nor U6953 (N_6953,N_1880,N_2508);
nand U6954 (N_6954,N_1778,N_216);
nor U6955 (N_6955,N_550,N_3065);
nand U6956 (N_6956,N_1714,N_3001);
nor U6957 (N_6957,N_70,N_1485);
nand U6958 (N_6958,N_3870,N_4950);
nand U6959 (N_6959,N_1040,N_3056);
and U6960 (N_6960,N_453,N_387);
nand U6961 (N_6961,N_1436,N_3500);
nor U6962 (N_6962,N_2322,N_373);
xor U6963 (N_6963,N_487,N_3100);
or U6964 (N_6964,N_1411,N_773);
or U6965 (N_6965,N_1786,N_4614);
nand U6966 (N_6966,N_277,N_533);
and U6967 (N_6967,N_172,N_414);
and U6968 (N_6968,N_442,N_2474);
and U6969 (N_6969,N_4076,N_3215);
and U6970 (N_6970,N_1457,N_3295);
or U6971 (N_6971,N_2939,N_942);
nor U6972 (N_6972,N_4379,N_1797);
and U6973 (N_6973,N_4532,N_4041);
and U6974 (N_6974,N_3173,N_3886);
nor U6975 (N_6975,N_2228,N_2491);
and U6976 (N_6976,N_1639,N_4564);
nor U6977 (N_6977,N_4241,N_1447);
nand U6978 (N_6978,N_830,N_788);
or U6979 (N_6979,N_2957,N_3479);
or U6980 (N_6980,N_1966,N_1163);
or U6981 (N_6981,N_305,N_651);
nor U6982 (N_6982,N_1720,N_2467);
and U6983 (N_6983,N_1725,N_703);
xor U6984 (N_6984,N_3581,N_4805);
or U6985 (N_6985,N_1544,N_124);
nand U6986 (N_6986,N_2545,N_3638);
or U6987 (N_6987,N_4542,N_51);
and U6988 (N_6988,N_2733,N_1344);
nor U6989 (N_6989,N_3046,N_3268);
or U6990 (N_6990,N_4584,N_2759);
xor U6991 (N_6991,N_1259,N_2019);
and U6992 (N_6992,N_3055,N_2693);
nand U6993 (N_6993,N_3979,N_1099);
nand U6994 (N_6994,N_2885,N_1363);
nor U6995 (N_6995,N_2200,N_1105);
or U6996 (N_6996,N_3248,N_4933);
xor U6997 (N_6997,N_2241,N_3290);
xnor U6998 (N_6998,N_3612,N_2406);
nor U6999 (N_6999,N_1342,N_3353);
nor U7000 (N_7000,N_213,N_48);
nor U7001 (N_7001,N_313,N_4847);
and U7002 (N_7002,N_139,N_3633);
nand U7003 (N_7003,N_4690,N_1601);
nor U7004 (N_7004,N_1031,N_3643);
and U7005 (N_7005,N_1019,N_4939);
nor U7006 (N_7006,N_1713,N_4799);
nor U7007 (N_7007,N_3691,N_1135);
nand U7008 (N_7008,N_506,N_1426);
nor U7009 (N_7009,N_2715,N_4384);
xnor U7010 (N_7010,N_0,N_2989);
nor U7011 (N_7011,N_915,N_1590);
nor U7012 (N_7012,N_1633,N_2036);
or U7013 (N_7013,N_3110,N_4677);
nand U7014 (N_7014,N_3349,N_536);
or U7015 (N_7015,N_1446,N_4928);
xor U7016 (N_7016,N_521,N_4820);
or U7017 (N_7017,N_2292,N_3902);
and U7018 (N_7018,N_2111,N_1746);
nand U7019 (N_7019,N_2063,N_1676);
nand U7020 (N_7020,N_4322,N_3023);
or U7021 (N_7021,N_1225,N_622);
nand U7022 (N_7022,N_965,N_4431);
nor U7023 (N_7023,N_1269,N_3327);
and U7024 (N_7024,N_852,N_67);
nor U7025 (N_7025,N_3749,N_4489);
nand U7026 (N_7026,N_4642,N_168);
xnor U7027 (N_7027,N_485,N_2126);
nor U7028 (N_7028,N_911,N_4235);
or U7029 (N_7029,N_4977,N_1685);
nand U7030 (N_7030,N_3818,N_422);
and U7031 (N_7031,N_3493,N_2798);
nor U7032 (N_7032,N_1324,N_347);
or U7033 (N_7033,N_4366,N_1615);
and U7034 (N_7034,N_3613,N_639);
xnor U7035 (N_7035,N_2227,N_1556);
nand U7036 (N_7036,N_4447,N_4731);
and U7037 (N_7037,N_4230,N_2314);
or U7038 (N_7038,N_1901,N_1189);
xor U7039 (N_7039,N_4873,N_3625);
nor U7040 (N_7040,N_4931,N_4430);
xor U7041 (N_7041,N_2134,N_3504);
or U7042 (N_7042,N_1979,N_3804);
and U7043 (N_7043,N_2212,N_1983);
and U7044 (N_7044,N_3981,N_1496);
nand U7045 (N_7045,N_986,N_4179);
and U7046 (N_7046,N_1645,N_4605);
xor U7047 (N_7047,N_1475,N_3740);
and U7048 (N_7048,N_4177,N_4360);
and U7049 (N_7049,N_4223,N_4837);
nor U7050 (N_7050,N_295,N_3574);
and U7051 (N_7051,N_4296,N_4202);
or U7052 (N_7052,N_4387,N_4640);
or U7053 (N_7053,N_4626,N_2673);
nor U7054 (N_7054,N_1854,N_1721);
nand U7055 (N_7055,N_4877,N_4547);
and U7056 (N_7056,N_356,N_3690);
or U7057 (N_7057,N_1561,N_3224);
nor U7058 (N_7058,N_1772,N_2997);
nand U7059 (N_7059,N_3350,N_505);
or U7060 (N_7060,N_4967,N_2488);
or U7061 (N_7061,N_259,N_4325);
or U7062 (N_7062,N_279,N_4538);
nand U7063 (N_7063,N_3940,N_3996);
xnor U7064 (N_7064,N_2238,N_2014);
or U7065 (N_7065,N_4025,N_3508);
and U7066 (N_7066,N_3776,N_210);
and U7067 (N_7067,N_4604,N_3456);
or U7068 (N_7068,N_697,N_1255);
nand U7069 (N_7069,N_1923,N_4569);
xor U7070 (N_7070,N_2769,N_1672);
and U7071 (N_7071,N_4909,N_4148);
or U7072 (N_7072,N_1857,N_396);
nand U7073 (N_7073,N_2482,N_708);
nand U7074 (N_7074,N_2076,N_3571);
and U7075 (N_7075,N_1627,N_2709);
nand U7076 (N_7076,N_3274,N_3394);
nor U7077 (N_7077,N_742,N_19);
nor U7078 (N_7078,N_3032,N_4735);
or U7079 (N_7079,N_4663,N_867);
nor U7080 (N_7080,N_1295,N_2610);
or U7081 (N_7081,N_3898,N_452);
nor U7082 (N_7082,N_1947,N_3376);
nor U7083 (N_7083,N_2437,N_1465);
or U7084 (N_7084,N_4922,N_1533);
nand U7085 (N_7085,N_1992,N_3428);
and U7086 (N_7086,N_2438,N_4293);
nor U7087 (N_7087,N_932,N_3473);
and U7088 (N_7088,N_1524,N_2);
nor U7089 (N_7089,N_1102,N_3533);
nand U7090 (N_7090,N_4178,N_84);
nor U7091 (N_7091,N_4676,N_1034);
nor U7092 (N_7092,N_899,N_300);
nand U7093 (N_7093,N_4850,N_315);
nand U7094 (N_7094,N_3648,N_1717);
or U7095 (N_7095,N_1398,N_4728);
xnor U7096 (N_7096,N_2161,N_4636);
nor U7097 (N_7097,N_2537,N_3517);
and U7098 (N_7098,N_3942,N_3020);
nor U7099 (N_7099,N_2105,N_874);
nor U7100 (N_7100,N_2021,N_4698);
nand U7101 (N_7101,N_2913,N_498);
and U7102 (N_7102,N_1319,N_3545);
nand U7103 (N_7103,N_2184,N_2880);
and U7104 (N_7104,N_2520,N_2146);
xnor U7105 (N_7105,N_3445,N_335);
and U7106 (N_7106,N_57,N_1679);
or U7107 (N_7107,N_2468,N_2429);
or U7108 (N_7108,N_4861,N_289);
nor U7109 (N_7109,N_4775,N_824);
and U7110 (N_7110,N_3440,N_1547);
nor U7111 (N_7111,N_1849,N_3679);
nor U7112 (N_7112,N_507,N_1067);
and U7113 (N_7113,N_3978,N_4037);
nand U7114 (N_7114,N_175,N_2851);
nor U7115 (N_7115,N_4369,N_1270);
nor U7116 (N_7116,N_337,N_590);
and U7117 (N_7117,N_4639,N_565);
nand U7118 (N_7118,N_4495,N_3642);
nand U7119 (N_7119,N_2375,N_368);
and U7120 (N_7120,N_1171,N_1423);
and U7121 (N_7121,N_3515,N_2878);
and U7122 (N_7122,N_2638,N_3610);
xnor U7123 (N_7123,N_4940,N_144);
nand U7124 (N_7124,N_4390,N_574);
or U7125 (N_7125,N_1201,N_3028);
or U7126 (N_7126,N_2333,N_924);
nand U7127 (N_7127,N_3807,N_2739);
or U7128 (N_7128,N_383,N_3275);
nand U7129 (N_7129,N_1204,N_1768);
or U7130 (N_7130,N_3038,N_2944);
or U7131 (N_7131,N_2230,N_1290);
or U7132 (N_7132,N_918,N_174);
or U7133 (N_7133,N_8,N_4396);
and U7134 (N_7134,N_1374,N_3955);
nor U7135 (N_7135,N_4856,N_3012);
nand U7136 (N_7136,N_1477,N_1941);
and U7137 (N_7137,N_4442,N_3602);
nor U7138 (N_7138,N_1731,N_4315);
xnor U7139 (N_7139,N_1845,N_71);
xor U7140 (N_7140,N_2856,N_4274);
or U7141 (N_7141,N_98,N_4362);
or U7142 (N_7142,N_4862,N_76);
xnor U7143 (N_7143,N_982,N_2414);
or U7144 (N_7144,N_4038,N_4487);
nand U7145 (N_7145,N_3217,N_109);
nand U7146 (N_7146,N_382,N_2530);
nand U7147 (N_7147,N_2168,N_1153);
nand U7148 (N_7148,N_2648,N_3146);
xnor U7149 (N_7149,N_2381,N_1781);
and U7150 (N_7150,N_457,N_1059);
nor U7151 (N_7151,N_3594,N_763);
or U7152 (N_7152,N_334,N_3254);
and U7153 (N_7153,N_3656,N_3911);
or U7154 (N_7154,N_527,N_1858);
and U7155 (N_7155,N_3391,N_4330);
nand U7156 (N_7156,N_1492,N_2841);
and U7157 (N_7157,N_1531,N_2699);
nor U7158 (N_7158,N_1985,N_1722);
or U7159 (N_7159,N_3333,N_2410);
nor U7160 (N_7160,N_2922,N_4411);
nand U7161 (N_7161,N_4726,N_3629);
or U7162 (N_7162,N_4948,N_4469);
or U7163 (N_7163,N_2634,N_1216);
nor U7164 (N_7164,N_4693,N_3129);
nor U7165 (N_7165,N_3303,N_4252);
nor U7166 (N_7166,N_2044,N_2218);
and U7167 (N_7167,N_4212,N_233);
nor U7168 (N_7168,N_4403,N_2024);
or U7169 (N_7169,N_2563,N_3362);
and U7170 (N_7170,N_2304,N_4615);
nor U7171 (N_7171,N_1076,N_4835);
nor U7172 (N_7172,N_1254,N_3422);
nor U7173 (N_7173,N_712,N_4633);
nor U7174 (N_7174,N_4335,N_1285);
nand U7175 (N_7175,N_3766,N_2559);
and U7176 (N_7176,N_1016,N_2757);
nand U7177 (N_7177,N_1206,N_4540);
or U7178 (N_7178,N_2336,N_1262);
nor U7179 (N_7179,N_2556,N_4630);
nand U7180 (N_7180,N_1100,N_2213);
and U7181 (N_7181,N_3384,N_2487);
or U7182 (N_7182,N_2789,N_1007);
nor U7183 (N_7183,N_4531,N_4077);
and U7184 (N_7184,N_4581,N_2172);
nand U7185 (N_7185,N_3236,N_1680);
nor U7186 (N_7186,N_516,N_3525);
nor U7187 (N_7187,N_4017,N_4049);
and U7188 (N_7188,N_3145,N_838);
nor U7189 (N_7189,N_2706,N_15);
nand U7190 (N_7190,N_2041,N_4562);
and U7191 (N_7191,N_349,N_4674);
and U7192 (N_7192,N_806,N_2276);
nand U7193 (N_7193,N_2442,N_2258);
nand U7194 (N_7194,N_3169,N_4121);
or U7195 (N_7195,N_4150,N_3085);
xor U7196 (N_7196,N_4275,N_3513);
nand U7197 (N_7197,N_995,N_4602);
and U7198 (N_7198,N_4924,N_2245);
nand U7199 (N_7199,N_3965,N_3827);
nor U7200 (N_7200,N_864,N_554);
nand U7201 (N_7201,N_3889,N_1700);
and U7202 (N_7202,N_476,N_1468);
nor U7203 (N_7203,N_2777,N_2727);
and U7204 (N_7204,N_2451,N_1053);
nor U7205 (N_7205,N_926,N_4685);
or U7206 (N_7206,N_3108,N_1127);
nand U7207 (N_7207,N_3539,N_1353);
nor U7208 (N_7208,N_1879,N_3082);
and U7209 (N_7209,N_3830,N_944);
or U7210 (N_7210,N_4066,N_3318);
and U7211 (N_7211,N_1534,N_489);
or U7212 (N_7212,N_185,N_4240);
and U7213 (N_7213,N_3356,N_62);
nor U7214 (N_7214,N_4160,N_254);
nand U7215 (N_7215,N_3453,N_502);
or U7216 (N_7216,N_4908,N_4854);
and U7217 (N_7217,N_2494,N_666);
or U7218 (N_7218,N_1456,N_4954);
nand U7219 (N_7219,N_1565,N_3934);
and U7220 (N_7220,N_378,N_417);
xor U7221 (N_7221,N_2775,N_3585);
and U7222 (N_7222,N_4859,N_619);
xor U7223 (N_7223,N_4897,N_4167);
and U7224 (N_7224,N_1180,N_4872);
and U7225 (N_7225,N_272,N_4359);
and U7226 (N_7226,N_106,N_344);
nand U7227 (N_7227,N_2093,N_2681);
nand U7228 (N_7228,N_955,N_4519);
or U7229 (N_7229,N_1272,N_1257);
nand U7230 (N_7230,N_1089,N_2001);
or U7231 (N_7231,N_1307,N_3430);
and U7232 (N_7232,N_3796,N_706);
nand U7233 (N_7233,N_888,N_2065);
or U7234 (N_7234,N_3659,N_3502);
nand U7235 (N_7235,N_1572,N_1814);
xnor U7236 (N_7236,N_1061,N_1913);
nand U7237 (N_7237,N_3846,N_1593);
xor U7238 (N_7238,N_1745,N_183);
and U7239 (N_7239,N_4336,N_4570);
or U7240 (N_7240,N_64,N_4787);
xor U7241 (N_7241,N_4128,N_285);
nand U7242 (N_7242,N_1943,N_3718);
and U7243 (N_7243,N_3000,N_1664);
xor U7244 (N_7244,N_1481,N_4509);
or U7245 (N_7245,N_2247,N_2248);
nand U7246 (N_7246,N_468,N_3900);
xor U7247 (N_7247,N_4416,N_4106);
nor U7248 (N_7248,N_481,N_3640);
nor U7249 (N_7249,N_376,N_1355);
nand U7250 (N_7250,N_3262,N_3514);
nand U7251 (N_7251,N_1507,N_1166);
nand U7252 (N_7252,N_2755,N_2158);
and U7253 (N_7253,N_4669,N_2778);
and U7254 (N_7254,N_4124,N_3341);
or U7255 (N_7255,N_100,N_551);
or U7256 (N_7256,N_3523,N_3820);
and U7257 (N_7257,N_4409,N_2300);
nor U7258 (N_7258,N_17,N_2621);
and U7259 (N_7259,N_2743,N_4857);
or U7260 (N_7260,N_1630,N_2350);
nor U7261 (N_7261,N_1118,N_3049);
nand U7262 (N_7262,N_2599,N_2480);
nor U7263 (N_7263,N_4667,N_3154);
nor U7264 (N_7264,N_3363,N_177);
or U7265 (N_7265,N_2975,N_2783);
nor U7266 (N_7266,N_1542,N_3266);
nand U7267 (N_7267,N_384,N_2985);
nand U7268 (N_7268,N_4912,N_4863);
nand U7269 (N_7269,N_3336,N_2962);
nor U7270 (N_7270,N_187,N_3423);
or U7271 (N_7271,N_1417,N_3043);
nand U7272 (N_7272,N_684,N_614);
nand U7273 (N_7273,N_3556,N_2506);
nand U7274 (N_7274,N_2133,N_1074);
nand U7275 (N_7275,N_4879,N_4110);
or U7276 (N_7276,N_94,N_2281);
nand U7277 (N_7277,N_4046,N_2575);
nor U7278 (N_7278,N_2577,N_2167);
nand U7279 (N_7279,N_2042,N_4846);
or U7280 (N_7280,N_3249,N_4550);
and U7281 (N_7281,N_4182,N_123);
and U7282 (N_7282,N_769,N_1442);
or U7283 (N_7283,N_1964,N_3906);
and U7284 (N_7284,N_193,N_1097);
nand U7285 (N_7285,N_635,N_3232);
and U7286 (N_7286,N_2152,N_881);
or U7287 (N_7287,N_4503,N_4181);
nand U7288 (N_7288,N_1942,N_2604);
or U7289 (N_7289,N_4375,N_3855);
and U7290 (N_7290,N_711,N_4478);
xnor U7291 (N_7291,N_979,N_3233);
nor U7292 (N_7292,N_1400,N_675);
nor U7293 (N_7293,N_4326,N_3904);
nand U7294 (N_7294,N_1818,N_1335);
xor U7295 (N_7295,N_1484,N_587);
and U7296 (N_7296,N_3794,N_4278);
or U7297 (N_7297,N_4670,N_2327);
or U7298 (N_7298,N_3761,N_2717);
or U7299 (N_7299,N_3733,N_4363);
or U7300 (N_7300,N_4976,N_2833);
and U7301 (N_7301,N_3702,N_541);
nor U7302 (N_7302,N_2735,N_4007);
and U7303 (N_7303,N_4424,N_1859);
nor U7304 (N_7304,N_311,N_531);
nand U7305 (N_7305,N_567,N_607);
or U7306 (N_7306,N_1661,N_2096);
nor U7307 (N_7307,N_3011,N_3413);
nand U7308 (N_7308,N_4766,N_1248);
xor U7309 (N_7309,N_3518,N_147);
nand U7310 (N_7310,N_1317,N_4678);
nand U7311 (N_7311,N_4903,N_2801);
xnor U7312 (N_7312,N_4809,N_2824);
nor U7313 (N_7313,N_1698,N_303);
xnor U7314 (N_7314,N_3481,N_1888);
and U7315 (N_7315,N_2593,N_632);
nand U7316 (N_7316,N_3771,N_93);
or U7317 (N_7317,N_2354,N_3024);
or U7318 (N_7318,N_223,N_556);
nor U7319 (N_7319,N_3260,N_1724);
nand U7320 (N_7320,N_137,N_4445);
xnor U7321 (N_7321,N_4426,N_686);
or U7322 (N_7322,N_4913,N_970);
nor U7323 (N_7323,N_3044,N_4340);
nor U7324 (N_7324,N_4197,N_3098);
and U7325 (N_7325,N_1134,N_4644);
nand U7326 (N_7326,N_2923,N_517);
and U7327 (N_7327,N_2274,N_1387);
nand U7328 (N_7328,N_3719,N_2462);
nand U7329 (N_7329,N_1244,N_1478);
nand U7330 (N_7330,N_4079,N_1028);
nand U7331 (N_7331,N_4556,N_38);
nand U7332 (N_7332,N_1959,N_909);
nor U7333 (N_7333,N_4485,N_2229);
nand U7334 (N_7334,N_1584,N_1283);
and U7335 (N_7335,N_322,N_2290);
or U7336 (N_7336,N_3619,N_4708);
or U7337 (N_7337,N_1575,N_1509);
nand U7338 (N_7338,N_762,N_2450);
nand U7339 (N_7339,N_1190,N_4395);
nor U7340 (N_7340,N_157,N_1519);
nand U7341 (N_7341,N_2122,N_4265);
nand U7342 (N_7342,N_853,N_3722);
nand U7343 (N_7343,N_903,N_3273);
xor U7344 (N_7344,N_1666,N_749);
xnor U7345 (N_7345,N_1847,N_2169);
or U7346 (N_7346,N_3746,N_341);
and U7347 (N_7347,N_2393,N_966);
or U7348 (N_7348,N_4443,N_648);
or U7349 (N_7349,N_2445,N_1654);
xnor U7350 (N_7350,N_1211,N_3833);
or U7351 (N_7351,N_2541,N_2787);
nand U7352 (N_7352,N_2174,N_299);
nor U7353 (N_7353,N_2195,N_4777);
xor U7354 (N_7354,N_922,N_4995);
and U7355 (N_7355,N_1976,N_4589);
nor U7356 (N_7356,N_3183,N_281);
nand U7357 (N_7357,N_2805,N_808);
nand U7358 (N_7358,N_146,N_1842);
or U7359 (N_7359,N_3694,N_621);
or U7360 (N_7360,N_1758,N_2361);
nor U7361 (N_7361,N_1609,N_4715);
nand U7362 (N_7362,N_1691,N_4921);
xnor U7363 (N_7363,N_1431,N_4137);
nor U7364 (N_7364,N_2818,N_3847);
nor U7365 (N_7365,N_1905,N_1001);
and U7366 (N_7366,N_4821,N_672);
and U7367 (N_7367,N_4397,N_1652);
and U7368 (N_7368,N_4101,N_2876);
nor U7369 (N_7369,N_616,N_418);
nor U7370 (N_7370,N_3196,N_2339);
nand U7371 (N_7371,N_3402,N_4641);
nand U7372 (N_7372,N_1566,N_1462);
nor U7373 (N_7373,N_1929,N_4094);
and U7374 (N_7374,N_1742,N_496);
nand U7375 (N_7375,N_3824,N_2352);
or U7376 (N_7376,N_4772,N_154);
nor U7377 (N_7377,N_3506,N_4258);
nor U7378 (N_7378,N_1264,N_759);
nand U7379 (N_7379,N_2595,N_1602);
nand U7380 (N_7380,N_3973,N_702);
xnor U7381 (N_7381,N_1900,N_2157);
xnor U7382 (N_7382,N_1140,N_3418);
nand U7383 (N_7383,N_2934,N_3068);
and U7384 (N_7384,N_3022,N_3673);
nand U7385 (N_7385,N_1018,N_3035);
or U7386 (N_7386,N_4036,N_1663);
nand U7387 (N_7387,N_4050,N_1525);
or U7388 (N_7388,N_1653,N_3008);
nand U7389 (N_7389,N_2614,N_3630);
or U7390 (N_7390,N_4118,N_1840);
or U7391 (N_7391,N_4290,N_2873);
nor U7392 (N_7392,N_4925,N_844);
nor U7393 (N_7393,N_2016,N_3144);
or U7394 (N_7394,N_3451,N_2670);
and U7395 (N_7395,N_3251,N_3307);
nand U7396 (N_7396,N_1060,N_3130);
or U7397 (N_7397,N_411,N_4328);
nand U7398 (N_7398,N_298,N_1570);
or U7399 (N_7399,N_529,N_4523);
or U7400 (N_7400,N_4074,N_4986);
and U7401 (N_7401,N_2358,N_3253);
and U7402 (N_7402,N_3997,N_226);
nand U7403 (N_7403,N_1831,N_3823);
xor U7404 (N_7404,N_1990,N_1971);
nand U7405 (N_7405,N_4460,N_3646);
xnor U7406 (N_7406,N_323,N_657);
or U7407 (N_7407,N_2804,N_2840);
nand U7408 (N_7408,N_2283,N_179);
nor U7409 (N_7409,N_4830,N_1578);
or U7410 (N_7410,N_988,N_2607);
xor U7411 (N_7411,N_4356,N_941);
nor U7412 (N_7412,N_3727,N_3461);
or U7413 (N_7413,N_2319,N_1308);
xor U7414 (N_7414,N_1610,N_1011);
xnor U7415 (N_7415,N_592,N_1554);
and U7416 (N_7416,N_3837,N_4308);
nand U7417 (N_7417,N_443,N_1221);
or U7418 (N_7418,N_4404,N_245);
or U7419 (N_7419,N_4875,N_902);
nor U7420 (N_7420,N_4287,N_4132);
or U7421 (N_7421,N_3133,N_1822);
nor U7422 (N_7422,N_1767,N_1072);
and U7423 (N_7423,N_757,N_142);
xnor U7424 (N_7424,N_499,N_4104);
nand U7425 (N_7425,N_2051,N_4247);
xor U7426 (N_7426,N_156,N_2764);
nand U7427 (N_7427,N_2890,N_1882);
xnor U7428 (N_7428,N_571,N_1733);
xor U7429 (N_7429,N_1161,N_605);
and U7430 (N_7430,N_3983,N_3947);
nand U7431 (N_7431,N_1775,N_4022);
and U7432 (N_7432,N_4501,N_3598);
xor U7433 (N_7433,N_2355,N_472);
nand U7434 (N_7434,N_478,N_4122);
nor U7435 (N_7435,N_4966,N_4545);
nor U7436 (N_7436,N_4318,N_1603);
nor U7437 (N_7437,N_3966,N_1297);
or U7438 (N_7438,N_1466,N_4815);
and U7439 (N_7439,N_2688,N_3209);
or U7440 (N_7440,N_1549,N_4652);
nand U7441 (N_7441,N_3334,N_3591);
nor U7442 (N_7442,N_2952,N_923);
nand U7443 (N_7443,N_3474,N_2297);
and U7444 (N_7444,N_4895,N_4143);
xnor U7445 (N_7445,N_473,N_999);
nor U7446 (N_7446,N_4638,N_4);
or U7447 (N_7447,N_4544,N_2745);
or U7448 (N_7448,N_4832,N_4353);
and U7449 (N_7449,N_2924,N_579);
nor U7450 (N_7450,N_4329,N_3784);
and U7451 (N_7451,N_3050,N_5);
nor U7452 (N_7452,N_2214,N_2813);
nand U7453 (N_7453,N_3816,N_2940);
nand U7454 (N_7454,N_2071,N_4573);
and U7455 (N_7455,N_3314,N_4746);
nand U7456 (N_7456,N_338,N_1268);
or U7457 (N_7457,N_526,N_2459);
nand U7458 (N_7458,N_4793,N_4618);
xor U7459 (N_7459,N_3448,N_1440);
nor U7460 (N_7460,N_3326,N_2531);
nor U7461 (N_7461,N_4368,N_1798);
or U7462 (N_7462,N_2455,N_1291);
or U7463 (N_7463,N_3324,N_3409);
or U7464 (N_7464,N_1198,N_2552);
and U7465 (N_7465,N_4176,N_631);
nand U7466 (N_7466,N_3994,N_2394);
or U7467 (N_7467,N_308,N_1192);
or U7468 (N_7468,N_1437,N_1379);
and U7469 (N_7469,N_4524,N_4012);
or U7470 (N_7470,N_2523,N_1188);
and U7471 (N_7471,N_406,N_3123);
or U7472 (N_7472,N_1075,N_1794);
nor U7473 (N_7473,N_787,N_974);
nor U7474 (N_7474,N_3605,N_1004);
nor U7475 (N_7475,N_4656,N_2580);
nor U7476 (N_7476,N_2800,N_3291);
and U7477 (N_7477,N_1945,N_1104);
xnor U7478 (N_7478,N_1585,N_4824);
and U7479 (N_7479,N_4035,N_618);
nand U7480 (N_7480,N_1838,N_578);
nor U7481 (N_7481,N_4520,N_20);
xnor U7482 (N_7482,N_4407,N_939);
and U7483 (N_7483,N_4855,N_1049);
or U7484 (N_7484,N_1131,N_2592);
xor U7485 (N_7485,N_737,N_4289);
nor U7486 (N_7486,N_1050,N_4949);
or U7487 (N_7487,N_3482,N_3577);
or U7488 (N_7488,N_2842,N_610);
nand U7489 (N_7489,N_2337,N_3279);
or U7490 (N_7490,N_750,N_3835);
and U7491 (N_7491,N_1599,N_4434);
nand U7492 (N_7492,N_2766,N_4428);
or U7493 (N_7493,N_2502,N_2937);
and U7494 (N_7494,N_2007,N_682);
xnor U7495 (N_7495,N_4464,N_2183);
nand U7496 (N_7496,N_37,N_1303);
nor U7497 (N_7497,N_984,N_205);
nor U7498 (N_7498,N_1070,N_4213);
or U7499 (N_7499,N_4525,N_3534);
and U7500 (N_7500,N_3910,N_3160);
or U7501 (N_7501,N_2504,N_4587);
nor U7502 (N_7502,N_2595,N_347);
nor U7503 (N_7503,N_827,N_674);
and U7504 (N_7504,N_2453,N_2805);
nand U7505 (N_7505,N_2224,N_2849);
or U7506 (N_7506,N_2459,N_2007);
nand U7507 (N_7507,N_2761,N_4227);
nand U7508 (N_7508,N_1908,N_1576);
and U7509 (N_7509,N_932,N_4820);
nand U7510 (N_7510,N_562,N_3164);
nor U7511 (N_7511,N_1009,N_4367);
or U7512 (N_7512,N_1773,N_4444);
and U7513 (N_7513,N_829,N_3945);
nor U7514 (N_7514,N_1313,N_1470);
and U7515 (N_7515,N_2666,N_3200);
or U7516 (N_7516,N_4382,N_4885);
and U7517 (N_7517,N_106,N_503);
or U7518 (N_7518,N_3404,N_899);
and U7519 (N_7519,N_459,N_2402);
and U7520 (N_7520,N_1009,N_430);
nand U7521 (N_7521,N_849,N_3345);
nand U7522 (N_7522,N_1982,N_706);
nor U7523 (N_7523,N_952,N_3847);
xnor U7524 (N_7524,N_4691,N_1524);
nand U7525 (N_7525,N_4188,N_1270);
or U7526 (N_7526,N_295,N_278);
and U7527 (N_7527,N_68,N_1582);
or U7528 (N_7528,N_3257,N_2413);
nand U7529 (N_7529,N_1637,N_2849);
or U7530 (N_7530,N_312,N_1690);
nor U7531 (N_7531,N_2582,N_4965);
nor U7532 (N_7532,N_3069,N_2026);
nand U7533 (N_7533,N_408,N_3665);
xnor U7534 (N_7534,N_593,N_820);
or U7535 (N_7535,N_2176,N_2941);
or U7536 (N_7536,N_1973,N_4857);
or U7537 (N_7537,N_1546,N_1448);
xor U7538 (N_7538,N_2088,N_3910);
nor U7539 (N_7539,N_2765,N_3861);
nand U7540 (N_7540,N_2649,N_4609);
and U7541 (N_7541,N_1761,N_3751);
nor U7542 (N_7542,N_634,N_201);
xor U7543 (N_7543,N_2562,N_2085);
xor U7544 (N_7544,N_4872,N_883);
or U7545 (N_7545,N_3776,N_3019);
or U7546 (N_7546,N_497,N_1240);
nor U7547 (N_7547,N_3579,N_3380);
nor U7548 (N_7548,N_3928,N_1720);
and U7549 (N_7549,N_922,N_2674);
or U7550 (N_7550,N_2943,N_3523);
or U7551 (N_7551,N_3791,N_1449);
or U7552 (N_7552,N_2886,N_1947);
or U7553 (N_7553,N_4787,N_102);
or U7554 (N_7554,N_4891,N_496);
nor U7555 (N_7555,N_1325,N_49);
nor U7556 (N_7556,N_98,N_2454);
nand U7557 (N_7557,N_2883,N_2762);
nor U7558 (N_7558,N_2397,N_4063);
and U7559 (N_7559,N_1196,N_4259);
nor U7560 (N_7560,N_4012,N_1454);
xor U7561 (N_7561,N_485,N_510);
and U7562 (N_7562,N_233,N_4222);
or U7563 (N_7563,N_1398,N_3230);
nand U7564 (N_7564,N_3297,N_2787);
and U7565 (N_7565,N_3496,N_2758);
and U7566 (N_7566,N_225,N_2791);
xor U7567 (N_7567,N_291,N_592);
xnor U7568 (N_7568,N_1542,N_310);
nand U7569 (N_7569,N_3911,N_3172);
or U7570 (N_7570,N_1101,N_4742);
and U7571 (N_7571,N_4,N_972);
or U7572 (N_7572,N_657,N_3528);
nand U7573 (N_7573,N_117,N_3649);
nor U7574 (N_7574,N_1946,N_152);
nor U7575 (N_7575,N_4598,N_803);
or U7576 (N_7576,N_2218,N_2441);
and U7577 (N_7577,N_4032,N_1488);
and U7578 (N_7578,N_1686,N_669);
or U7579 (N_7579,N_2423,N_1360);
nand U7580 (N_7580,N_329,N_3657);
xor U7581 (N_7581,N_2904,N_3830);
or U7582 (N_7582,N_1489,N_4233);
nor U7583 (N_7583,N_664,N_3287);
nand U7584 (N_7584,N_3909,N_518);
and U7585 (N_7585,N_2559,N_4387);
xor U7586 (N_7586,N_771,N_4061);
and U7587 (N_7587,N_3015,N_3556);
or U7588 (N_7588,N_3218,N_4233);
or U7589 (N_7589,N_3061,N_1725);
nor U7590 (N_7590,N_1780,N_931);
and U7591 (N_7591,N_1036,N_622);
or U7592 (N_7592,N_2769,N_1495);
nor U7593 (N_7593,N_706,N_3972);
xor U7594 (N_7594,N_1307,N_4159);
xor U7595 (N_7595,N_3649,N_2894);
nand U7596 (N_7596,N_2333,N_2943);
nand U7597 (N_7597,N_2005,N_1503);
nor U7598 (N_7598,N_285,N_2597);
or U7599 (N_7599,N_794,N_1739);
nand U7600 (N_7600,N_3537,N_1344);
or U7601 (N_7601,N_2598,N_4906);
or U7602 (N_7602,N_2542,N_1649);
or U7603 (N_7603,N_475,N_1761);
or U7604 (N_7604,N_2292,N_2834);
or U7605 (N_7605,N_2748,N_883);
nand U7606 (N_7606,N_2011,N_251);
nand U7607 (N_7607,N_1808,N_1130);
nor U7608 (N_7608,N_1137,N_173);
and U7609 (N_7609,N_411,N_2646);
nor U7610 (N_7610,N_1183,N_3706);
nand U7611 (N_7611,N_3862,N_1601);
or U7612 (N_7612,N_4876,N_1596);
and U7613 (N_7613,N_3247,N_3690);
or U7614 (N_7614,N_1599,N_2516);
nand U7615 (N_7615,N_1512,N_2242);
or U7616 (N_7616,N_1108,N_757);
nor U7617 (N_7617,N_384,N_3689);
nand U7618 (N_7618,N_2734,N_1415);
nor U7619 (N_7619,N_1052,N_2004);
and U7620 (N_7620,N_4842,N_4501);
nand U7621 (N_7621,N_3900,N_4085);
or U7622 (N_7622,N_1052,N_1579);
and U7623 (N_7623,N_3606,N_1412);
nor U7624 (N_7624,N_2622,N_4126);
xor U7625 (N_7625,N_2086,N_358);
or U7626 (N_7626,N_542,N_4081);
or U7627 (N_7627,N_537,N_3417);
or U7628 (N_7628,N_1725,N_623);
nand U7629 (N_7629,N_1598,N_4790);
or U7630 (N_7630,N_1092,N_691);
nor U7631 (N_7631,N_1043,N_2571);
or U7632 (N_7632,N_4198,N_680);
and U7633 (N_7633,N_3811,N_764);
nand U7634 (N_7634,N_4710,N_3853);
or U7635 (N_7635,N_2631,N_2956);
or U7636 (N_7636,N_1145,N_2584);
nor U7637 (N_7637,N_4597,N_175);
or U7638 (N_7638,N_2839,N_1142);
and U7639 (N_7639,N_2529,N_3355);
xnor U7640 (N_7640,N_1136,N_2700);
and U7641 (N_7641,N_226,N_487);
or U7642 (N_7642,N_2062,N_1636);
nand U7643 (N_7643,N_762,N_692);
and U7644 (N_7644,N_2851,N_2611);
nor U7645 (N_7645,N_1408,N_519);
nand U7646 (N_7646,N_2592,N_4777);
nand U7647 (N_7647,N_4468,N_28);
or U7648 (N_7648,N_323,N_1851);
or U7649 (N_7649,N_3545,N_4098);
nor U7650 (N_7650,N_4384,N_1962);
nand U7651 (N_7651,N_4007,N_3199);
nor U7652 (N_7652,N_4976,N_286);
nor U7653 (N_7653,N_1353,N_418);
and U7654 (N_7654,N_1044,N_754);
and U7655 (N_7655,N_1182,N_2933);
xor U7656 (N_7656,N_727,N_2013);
xnor U7657 (N_7657,N_2679,N_285);
or U7658 (N_7658,N_4163,N_2231);
xnor U7659 (N_7659,N_2311,N_1471);
or U7660 (N_7660,N_485,N_1738);
nand U7661 (N_7661,N_1240,N_1550);
nor U7662 (N_7662,N_1302,N_3481);
nand U7663 (N_7663,N_3621,N_3229);
and U7664 (N_7664,N_2643,N_4151);
and U7665 (N_7665,N_2057,N_4034);
xnor U7666 (N_7666,N_2380,N_131);
nor U7667 (N_7667,N_4507,N_2859);
nor U7668 (N_7668,N_1051,N_832);
nand U7669 (N_7669,N_2576,N_4660);
nor U7670 (N_7670,N_4258,N_1510);
nor U7671 (N_7671,N_3705,N_1584);
or U7672 (N_7672,N_390,N_397);
nand U7673 (N_7673,N_310,N_4914);
xor U7674 (N_7674,N_433,N_916);
or U7675 (N_7675,N_1476,N_923);
nor U7676 (N_7676,N_1019,N_3322);
and U7677 (N_7677,N_480,N_1342);
or U7678 (N_7678,N_4297,N_3046);
nor U7679 (N_7679,N_1779,N_2142);
nand U7680 (N_7680,N_3289,N_3812);
nor U7681 (N_7681,N_3685,N_1007);
xnor U7682 (N_7682,N_1573,N_3598);
nand U7683 (N_7683,N_1788,N_3582);
nor U7684 (N_7684,N_2044,N_2834);
or U7685 (N_7685,N_2856,N_1558);
nand U7686 (N_7686,N_4143,N_4809);
nand U7687 (N_7687,N_2166,N_2604);
nand U7688 (N_7688,N_439,N_550);
nand U7689 (N_7689,N_3063,N_36);
and U7690 (N_7690,N_4475,N_4059);
and U7691 (N_7691,N_4045,N_1097);
nor U7692 (N_7692,N_1001,N_1280);
or U7693 (N_7693,N_2654,N_1466);
or U7694 (N_7694,N_4105,N_794);
and U7695 (N_7695,N_2630,N_2724);
and U7696 (N_7696,N_3268,N_4564);
and U7697 (N_7697,N_2706,N_4143);
nand U7698 (N_7698,N_144,N_1885);
nand U7699 (N_7699,N_4874,N_685);
nand U7700 (N_7700,N_1125,N_3936);
or U7701 (N_7701,N_2735,N_1736);
or U7702 (N_7702,N_1210,N_3865);
and U7703 (N_7703,N_4798,N_873);
or U7704 (N_7704,N_892,N_2100);
nor U7705 (N_7705,N_4949,N_1957);
xnor U7706 (N_7706,N_1216,N_1259);
or U7707 (N_7707,N_622,N_3627);
and U7708 (N_7708,N_2670,N_38);
and U7709 (N_7709,N_2379,N_2200);
nor U7710 (N_7710,N_1536,N_1075);
nand U7711 (N_7711,N_87,N_3911);
nand U7712 (N_7712,N_929,N_3395);
nor U7713 (N_7713,N_1974,N_1417);
or U7714 (N_7714,N_1467,N_4188);
and U7715 (N_7715,N_2495,N_4301);
nand U7716 (N_7716,N_334,N_4375);
nand U7717 (N_7717,N_1663,N_2325);
nor U7718 (N_7718,N_2224,N_2500);
nor U7719 (N_7719,N_4538,N_1951);
and U7720 (N_7720,N_3689,N_1195);
and U7721 (N_7721,N_2318,N_3821);
nand U7722 (N_7722,N_950,N_4509);
and U7723 (N_7723,N_38,N_434);
xnor U7724 (N_7724,N_165,N_3965);
nand U7725 (N_7725,N_4974,N_2304);
nand U7726 (N_7726,N_2452,N_1283);
nor U7727 (N_7727,N_478,N_1903);
or U7728 (N_7728,N_604,N_4635);
nor U7729 (N_7729,N_4239,N_20);
or U7730 (N_7730,N_1807,N_1110);
nand U7731 (N_7731,N_2041,N_1353);
nor U7732 (N_7732,N_615,N_313);
nor U7733 (N_7733,N_3259,N_760);
or U7734 (N_7734,N_3011,N_2428);
nor U7735 (N_7735,N_1879,N_3757);
and U7736 (N_7736,N_540,N_499);
nand U7737 (N_7737,N_3196,N_1232);
and U7738 (N_7738,N_2900,N_1252);
nand U7739 (N_7739,N_3655,N_1565);
xnor U7740 (N_7740,N_3687,N_4053);
nand U7741 (N_7741,N_2426,N_2855);
and U7742 (N_7742,N_2641,N_803);
and U7743 (N_7743,N_1230,N_4643);
nor U7744 (N_7744,N_4819,N_3916);
nand U7745 (N_7745,N_1602,N_1403);
and U7746 (N_7746,N_1221,N_4490);
and U7747 (N_7747,N_1245,N_3570);
nor U7748 (N_7748,N_2097,N_3404);
nor U7749 (N_7749,N_2295,N_1329);
nand U7750 (N_7750,N_4554,N_4714);
and U7751 (N_7751,N_428,N_2293);
or U7752 (N_7752,N_4738,N_2492);
or U7753 (N_7753,N_39,N_231);
nor U7754 (N_7754,N_3746,N_1921);
or U7755 (N_7755,N_1873,N_1264);
nor U7756 (N_7756,N_744,N_2885);
and U7757 (N_7757,N_1008,N_4317);
or U7758 (N_7758,N_1989,N_2377);
nor U7759 (N_7759,N_3773,N_3357);
and U7760 (N_7760,N_1979,N_422);
nand U7761 (N_7761,N_3734,N_1011);
or U7762 (N_7762,N_4462,N_2725);
xnor U7763 (N_7763,N_1944,N_4304);
and U7764 (N_7764,N_869,N_987);
or U7765 (N_7765,N_304,N_2944);
or U7766 (N_7766,N_2391,N_2191);
and U7767 (N_7767,N_1343,N_3448);
xor U7768 (N_7768,N_2823,N_3412);
nor U7769 (N_7769,N_4681,N_3310);
nor U7770 (N_7770,N_1244,N_4709);
or U7771 (N_7771,N_3046,N_3132);
nand U7772 (N_7772,N_632,N_2729);
or U7773 (N_7773,N_427,N_149);
nor U7774 (N_7774,N_2355,N_897);
and U7775 (N_7775,N_1854,N_3160);
nor U7776 (N_7776,N_1115,N_1950);
or U7777 (N_7777,N_2902,N_753);
nor U7778 (N_7778,N_653,N_4088);
nor U7779 (N_7779,N_2304,N_3419);
and U7780 (N_7780,N_2348,N_3555);
nor U7781 (N_7781,N_3752,N_446);
nand U7782 (N_7782,N_4992,N_2411);
nand U7783 (N_7783,N_1157,N_3640);
nand U7784 (N_7784,N_1949,N_3830);
and U7785 (N_7785,N_2895,N_2153);
or U7786 (N_7786,N_2021,N_2081);
or U7787 (N_7787,N_2552,N_4558);
and U7788 (N_7788,N_1233,N_4862);
or U7789 (N_7789,N_90,N_400);
nor U7790 (N_7790,N_850,N_4850);
nand U7791 (N_7791,N_4555,N_3238);
and U7792 (N_7792,N_603,N_3513);
and U7793 (N_7793,N_3621,N_3120);
and U7794 (N_7794,N_3216,N_1286);
and U7795 (N_7795,N_277,N_3192);
or U7796 (N_7796,N_1183,N_2423);
nand U7797 (N_7797,N_627,N_3136);
xnor U7798 (N_7798,N_3654,N_4193);
nor U7799 (N_7799,N_4166,N_1103);
nand U7800 (N_7800,N_4614,N_72);
nor U7801 (N_7801,N_3903,N_3647);
xnor U7802 (N_7802,N_318,N_4882);
or U7803 (N_7803,N_670,N_4765);
nand U7804 (N_7804,N_2523,N_4550);
nand U7805 (N_7805,N_3142,N_2346);
xor U7806 (N_7806,N_1268,N_989);
and U7807 (N_7807,N_2880,N_4963);
nand U7808 (N_7808,N_3742,N_419);
or U7809 (N_7809,N_2445,N_1595);
nand U7810 (N_7810,N_1985,N_3804);
xnor U7811 (N_7811,N_2506,N_893);
or U7812 (N_7812,N_791,N_2303);
or U7813 (N_7813,N_4812,N_1428);
nand U7814 (N_7814,N_3153,N_2281);
nand U7815 (N_7815,N_449,N_4438);
nor U7816 (N_7816,N_2746,N_619);
nor U7817 (N_7817,N_1296,N_4524);
nor U7818 (N_7818,N_2353,N_3869);
nand U7819 (N_7819,N_2012,N_231);
or U7820 (N_7820,N_4064,N_4297);
nor U7821 (N_7821,N_152,N_75);
xnor U7822 (N_7822,N_3746,N_1891);
nor U7823 (N_7823,N_4711,N_2415);
or U7824 (N_7824,N_1417,N_442);
or U7825 (N_7825,N_1879,N_1149);
or U7826 (N_7826,N_4666,N_2640);
nand U7827 (N_7827,N_653,N_4397);
xnor U7828 (N_7828,N_170,N_2048);
nor U7829 (N_7829,N_4364,N_4268);
nor U7830 (N_7830,N_3296,N_85);
or U7831 (N_7831,N_3338,N_3898);
nor U7832 (N_7832,N_4517,N_2085);
nor U7833 (N_7833,N_3650,N_2551);
and U7834 (N_7834,N_4255,N_3730);
nand U7835 (N_7835,N_3887,N_2960);
or U7836 (N_7836,N_1508,N_82);
nand U7837 (N_7837,N_4576,N_2903);
and U7838 (N_7838,N_1138,N_234);
or U7839 (N_7839,N_964,N_2904);
nand U7840 (N_7840,N_2564,N_175);
nor U7841 (N_7841,N_1838,N_2129);
nor U7842 (N_7842,N_4667,N_312);
nor U7843 (N_7843,N_197,N_3291);
nor U7844 (N_7844,N_1751,N_1315);
or U7845 (N_7845,N_1635,N_603);
nand U7846 (N_7846,N_1237,N_1681);
nor U7847 (N_7847,N_4457,N_2057);
and U7848 (N_7848,N_4459,N_789);
and U7849 (N_7849,N_3996,N_4395);
or U7850 (N_7850,N_196,N_2994);
and U7851 (N_7851,N_4075,N_3026);
or U7852 (N_7852,N_4015,N_2277);
and U7853 (N_7853,N_3548,N_1225);
nand U7854 (N_7854,N_3886,N_662);
and U7855 (N_7855,N_3259,N_3917);
and U7856 (N_7856,N_514,N_3371);
and U7857 (N_7857,N_2882,N_1483);
and U7858 (N_7858,N_1633,N_2732);
nor U7859 (N_7859,N_2140,N_3449);
nor U7860 (N_7860,N_4894,N_4035);
and U7861 (N_7861,N_4688,N_2933);
nand U7862 (N_7862,N_4690,N_3038);
xor U7863 (N_7863,N_258,N_923);
and U7864 (N_7864,N_4133,N_4532);
nand U7865 (N_7865,N_4835,N_4603);
and U7866 (N_7866,N_2133,N_3582);
nor U7867 (N_7867,N_2256,N_1240);
and U7868 (N_7868,N_3136,N_2744);
nor U7869 (N_7869,N_948,N_1076);
nor U7870 (N_7870,N_4423,N_701);
nor U7871 (N_7871,N_1825,N_3113);
or U7872 (N_7872,N_432,N_465);
or U7873 (N_7873,N_4356,N_1543);
nor U7874 (N_7874,N_3364,N_790);
nor U7875 (N_7875,N_241,N_538);
or U7876 (N_7876,N_1162,N_2771);
nor U7877 (N_7877,N_3952,N_465);
and U7878 (N_7878,N_3654,N_472);
nand U7879 (N_7879,N_2305,N_2634);
and U7880 (N_7880,N_4253,N_765);
nor U7881 (N_7881,N_735,N_4521);
nor U7882 (N_7882,N_2907,N_3729);
or U7883 (N_7883,N_1373,N_2922);
or U7884 (N_7884,N_1203,N_1754);
nor U7885 (N_7885,N_3594,N_4504);
or U7886 (N_7886,N_3481,N_2479);
nand U7887 (N_7887,N_266,N_966);
nor U7888 (N_7888,N_2969,N_1609);
and U7889 (N_7889,N_484,N_192);
or U7890 (N_7890,N_4786,N_1174);
and U7891 (N_7891,N_935,N_540);
or U7892 (N_7892,N_25,N_3209);
nor U7893 (N_7893,N_2264,N_2621);
nand U7894 (N_7894,N_1764,N_4335);
or U7895 (N_7895,N_1227,N_1739);
xnor U7896 (N_7896,N_3700,N_1841);
nor U7897 (N_7897,N_4375,N_1631);
nor U7898 (N_7898,N_3970,N_230);
xor U7899 (N_7899,N_3649,N_3559);
nor U7900 (N_7900,N_1928,N_92);
or U7901 (N_7901,N_3723,N_4161);
or U7902 (N_7902,N_1728,N_1693);
or U7903 (N_7903,N_1294,N_151);
nor U7904 (N_7904,N_2278,N_4057);
nor U7905 (N_7905,N_231,N_4560);
xnor U7906 (N_7906,N_3356,N_1776);
nand U7907 (N_7907,N_3785,N_3421);
nor U7908 (N_7908,N_1335,N_4076);
and U7909 (N_7909,N_4423,N_4659);
nor U7910 (N_7910,N_4322,N_617);
or U7911 (N_7911,N_1751,N_304);
and U7912 (N_7912,N_2931,N_2322);
nor U7913 (N_7913,N_4961,N_968);
and U7914 (N_7914,N_2846,N_7);
or U7915 (N_7915,N_4540,N_4468);
nand U7916 (N_7916,N_4575,N_468);
or U7917 (N_7917,N_4793,N_2229);
xor U7918 (N_7918,N_1591,N_2654);
nor U7919 (N_7919,N_1149,N_17);
or U7920 (N_7920,N_4330,N_2770);
nor U7921 (N_7921,N_4249,N_2122);
nor U7922 (N_7922,N_2738,N_3937);
or U7923 (N_7923,N_2325,N_2429);
and U7924 (N_7924,N_2694,N_4482);
or U7925 (N_7925,N_1787,N_2361);
xor U7926 (N_7926,N_980,N_3537);
or U7927 (N_7927,N_654,N_2019);
or U7928 (N_7928,N_2175,N_2229);
and U7929 (N_7929,N_1169,N_2935);
or U7930 (N_7930,N_602,N_4905);
or U7931 (N_7931,N_660,N_738);
xor U7932 (N_7932,N_1859,N_3590);
nand U7933 (N_7933,N_4743,N_3819);
or U7934 (N_7934,N_2550,N_2641);
or U7935 (N_7935,N_3889,N_495);
nand U7936 (N_7936,N_562,N_73);
or U7937 (N_7937,N_562,N_2171);
nor U7938 (N_7938,N_2792,N_3163);
xnor U7939 (N_7939,N_482,N_2406);
nor U7940 (N_7940,N_3219,N_1802);
nand U7941 (N_7941,N_1283,N_2143);
or U7942 (N_7942,N_1973,N_55);
nor U7943 (N_7943,N_1406,N_1654);
xor U7944 (N_7944,N_678,N_4714);
nor U7945 (N_7945,N_4283,N_1115);
nand U7946 (N_7946,N_2887,N_4406);
nand U7947 (N_7947,N_509,N_137);
and U7948 (N_7948,N_2029,N_2437);
xor U7949 (N_7949,N_4575,N_3780);
and U7950 (N_7950,N_4616,N_1864);
nand U7951 (N_7951,N_4262,N_4919);
nand U7952 (N_7952,N_1508,N_4491);
nor U7953 (N_7953,N_1221,N_579);
nand U7954 (N_7954,N_1099,N_4938);
nand U7955 (N_7955,N_3334,N_4555);
nand U7956 (N_7956,N_1709,N_1901);
or U7957 (N_7957,N_3946,N_2580);
and U7958 (N_7958,N_4320,N_3346);
and U7959 (N_7959,N_1707,N_4979);
or U7960 (N_7960,N_2810,N_2007);
and U7961 (N_7961,N_4686,N_4042);
and U7962 (N_7962,N_614,N_595);
or U7963 (N_7963,N_2968,N_4370);
or U7964 (N_7964,N_2205,N_1696);
nand U7965 (N_7965,N_3095,N_2170);
or U7966 (N_7966,N_1638,N_675);
xnor U7967 (N_7967,N_3649,N_720);
and U7968 (N_7968,N_431,N_307);
and U7969 (N_7969,N_1111,N_1717);
or U7970 (N_7970,N_4750,N_3061);
or U7971 (N_7971,N_4688,N_832);
or U7972 (N_7972,N_2766,N_1787);
nand U7973 (N_7973,N_3394,N_1872);
or U7974 (N_7974,N_2543,N_1274);
or U7975 (N_7975,N_4719,N_1122);
xor U7976 (N_7976,N_4285,N_2819);
and U7977 (N_7977,N_2136,N_1744);
xor U7978 (N_7978,N_4011,N_1973);
or U7979 (N_7979,N_2222,N_2225);
nor U7980 (N_7980,N_4157,N_2032);
xnor U7981 (N_7981,N_1324,N_4553);
or U7982 (N_7982,N_4272,N_2888);
nand U7983 (N_7983,N_3935,N_2402);
nand U7984 (N_7984,N_3051,N_1013);
nor U7985 (N_7985,N_507,N_1102);
nor U7986 (N_7986,N_4974,N_3268);
nor U7987 (N_7987,N_2649,N_2514);
or U7988 (N_7988,N_4331,N_1878);
xor U7989 (N_7989,N_2923,N_2857);
and U7990 (N_7990,N_1958,N_3260);
or U7991 (N_7991,N_3164,N_4623);
xor U7992 (N_7992,N_871,N_1379);
or U7993 (N_7993,N_48,N_4682);
xor U7994 (N_7994,N_2442,N_2997);
or U7995 (N_7995,N_2522,N_3754);
xor U7996 (N_7996,N_2198,N_402);
nor U7997 (N_7997,N_6,N_3472);
and U7998 (N_7998,N_2556,N_1987);
and U7999 (N_7999,N_1664,N_1706);
nand U8000 (N_8000,N_1871,N_4684);
nand U8001 (N_8001,N_2585,N_2311);
nor U8002 (N_8002,N_3192,N_4783);
or U8003 (N_8003,N_4998,N_499);
nor U8004 (N_8004,N_1553,N_3300);
or U8005 (N_8005,N_103,N_997);
and U8006 (N_8006,N_2892,N_620);
or U8007 (N_8007,N_1140,N_3541);
nor U8008 (N_8008,N_4404,N_619);
and U8009 (N_8009,N_2116,N_1967);
nand U8010 (N_8010,N_2180,N_236);
and U8011 (N_8011,N_2247,N_4809);
xor U8012 (N_8012,N_3313,N_1085);
nand U8013 (N_8013,N_1180,N_2024);
nand U8014 (N_8014,N_4205,N_1493);
xor U8015 (N_8015,N_3518,N_3731);
and U8016 (N_8016,N_4223,N_4634);
and U8017 (N_8017,N_4621,N_260);
or U8018 (N_8018,N_3464,N_4507);
and U8019 (N_8019,N_282,N_1900);
and U8020 (N_8020,N_1338,N_2362);
nand U8021 (N_8021,N_1993,N_4525);
or U8022 (N_8022,N_2054,N_3968);
and U8023 (N_8023,N_3570,N_2339);
nand U8024 (N_8024,N_865,N_2810);
and U8025 (N_8025,N_3206,N_721);
or U8026 (N_8026,N_4541,N_1366);
and U8027 (N_8027,N_2248,N_2546);
nand U8028 (N_8028,N_360,N_358);
and U8029 (N_8029,N_2161,N_4333);
xor U8030 (N_8030,N_3120,N_4435);
and U8031 (N_8031,N_1756,N_2358);
or U8032 (N_8032,N_1684,N_2924);
and U8033 (N_8033,N_2097,N_2176);
nor U8034 (N_8034,N_4410,N_2731);
and U8035 (N_8035,N_4065,N_737);
or U8036 (N_8036,N_3247,N_178);
and U8037 (N_8037,N_1267,N_1536);
and U8038 (N_8038,N_112,N_1455);
and U8039 (N_8039,N_3723,N_131);
or U8040 (N_8040,N_2966,N_1526);
nand U8041 (N_8041,N_3819,N_3473);
xor U8042 (N_8042,N_4837,N_2692);
nor U8043 (N_8043,N_3197,N_1874);
and U8044 (N_8044,N_2611,N_1488);
nand U8045 (N_8045,N_1493,N_3076);
nand U8046 (N_8046,N_1318,N_1458);
nor U8047 (N_8047,N_258,N_2068);
or U8048 (N_8048,N_547,N_736);
nand U8049 (N_8049,N_3440,N_216);
nor U8050 (N_8050,N_1810,N_4226);
and U8051 (N_8051,N_195,N_3789);
or U8052 (N_8052,N_1513,N_4223);
xor U8053 (N_8053,N_1542,N_3811);
nor U8054 (N_8054,N_3925,N_1312);
nor U8055 (N_8055,N_2178,N_445);
nor U8056 (N_8056,N_3797,N_4743);
and U8057 (N_8057,N_3947,N_1056);
nand U8058 (N_8058,N_3717,N_4051);
or U8059 (N_8059,N_2642,N_4273);
nand U8060 (N_8060,N_1486,N_338);
xnor U8061 (N_8061,N_1990,N_4110);
xor U8062 (N_8062,N_2907,N_4680);
or U8063 (N_8063,N_4271,N_3364);
nand U8064 (N_8064,N_3586,N_2419);
nor U8065 (N_8065,N_1754,N_128);
nor U8066 (N_8066,N_1659,N_4700);
or U8067 (N_8067,N_3075,N_1767);
or U8068 (N_8068,N_20,N_2882);
xor U8069 (N_8069,N_3457,N_4554);
nand U8070 (N_8070,N_2007,N_2023);
or U8071 (N_8071,N_3226,N_3422);
nand U8072 (N_8072,N_2427,N_3707);
and U8073 (N_8073,N_2455,N_4033);
and U8074 (N_8074,N_828,N_3929);
or U8075 (N_8075,N_155,N_1659);
or U8076 (N_8076,N_1501,N_874);
or U8077 (N_8077,N_4057,N_2602);
nand U8078 (N_8078,N_1712,N_3865);
xnor U8079 (N_8079,N_1348,N_4824);
and U8080 (N_8080,N_2444,N_3053);
and U8081 (N_8081,N_4528,N_2921);
nor U8082 (N_8082,N_4057,N_2699);
xor U8083 (N_8083,N_2569,N_3145);
and U8084 (N_8084,N_4099,N_209);
and U8085 (N_8085,N_624,N_3256);
or U8086 (N_8086,N_4203,N_2071);
or U8087 (N_8087,N_3895,N_1053);
nand U8088 (N_8088,N_2501,N_1871);
nor U8089 (N_8089,N_4900,N_798);
and U8090 (N_8090,N_4317,N_2612);
and U8091 (N_8091,N_2673,N_4034);
nand U8092 (N_8092,N_4511,N_1985);
and U8093 (N_8093,N_2914,N_502);
and U8094 (N_8094,N_2619,N_919);
or U8095 (N_8095,N_1851,N_3297);
or U8096 (N_8096,N_667,N_3441);
and U8097 (N_8097,N_4487,N_2004);
nor U8098 (N_8098,N_4537,N_761);
xnor U8099 (N_8099,N_1367,N_4463);
or U8100 (N_8100,N_428,N_3600);
nor U8101 (N_8101,N_675,N_4411);
or U8102 (N_8102,N_2642,N_1551);
xnor U8103 (N_8103,N_1887,N_4277);
or U8104 (N_8104,N_812,N_136);
and U8105 (N_8105,N_4075,N_1071);
nor U8106 (N_8106,N_1341,N_3172);
or U8107 (N_8107,N_715,N_1931);
and U8108 (N_8108,N_202,N_220);
or U8109 (N_8109,N_832,N_1593);
and U8110 (N_8110,N_1222,N_4911);
xnor U8111 (N_8111,N_4278,N_1500);
nand U8112 (N_8112,N_2369,N_2270);
xnor U8113 (N_8113,N_1960,N_4538);
nand U8114 (N_8114,N_1591,N_4970);
nand U8115 (N_8115,N_1675,N_3865);
xnor U8116 (N_8116,N_2892,N_4996);
or U8117 (N_8117,N_2830,N_3681);
or U8118 (N_8118,N_57,N_1569);
and U8119 (N_8119,N_2936,N_3216);
or U8120 (N_8120,N_1886,N_3370);
and U8121 (N_8121,N_4700,N_593);
nor U8122 (N_8122,N_2343,N_2203);
xnor U8123 (N_8123,N_2947,N_4062);
and U8124 (N_8124,N_376,N_4143);
and U8125 (N_8125,N_4760,N_2400);
nand U8126 (N_8126,N_2553,N_2914);
nor U8127 (N_8127,N_2699,N_2048);
or U8128 (N_8128,N_4602,N_523);
nand U8129 (N_8129,N_4095,N_3306);
or U8130 (N_8130,N_1903,N_1058);
or U8131 (N_8131,N_20,N_824);
and U8132 (N_8132,N_4276,N_264);
nor U8133 (N_8133,N_4216,N_1846);
and U8134 (N_8134,N_4165,N_2573);
and U8135 (N_8135,N_1243,N_77);
nor U8136 (N_8136,N_2098,N_500);
or U8137 (N_8137,N_4877,N_3409);
and U8138 (N_8138,N_4867,N_543);
nand U8139 (N_8139,N_1541,N_3414);
and U8140 (N_8140,N_2483,N_719);
xnor U8141 (N_8141,N_649,N_4223);
nand U8142 (N_8142,N_1623,N_900);
and U8143 (N_8143,N_553,N_1692);
or U8144 (N_8144,N_534,N_3357);
nand U8145 (N_8145,N_2477,N_1110);
or U8146 (N_8146,N_4830,N_1499);
and U8147 (N_8147,N_4622,N_3690);
and U8148 (N_8148,N_4372,N_1703);
nand U8149 (N_8149,N_371,N_3788);
and U8150 (N_8150,N_768,N_1125);
nand U8151 (N_8151,N_1307,N_3636);
nand U8152 (N_8152,N_4755,N_1069);
xnor U8153 (N_8153,N_1017,N_1629);
nor U8154 (N_8154,N_4874,N_3161);
xnor U8155 (N_8155,N_1032,N_3053);
or U8156 (N_8156,N_2047,N_3707);
or U8157 (N_8157,N_2353,N_254);
nand U8158 (N_8158,N_1586,N_4740);
or U8159 (N_8159,N_3697,N_4288);
nand U8160 (N_8160,N_4359,N_2888);
and U8161 (N_8161,N_2597,N_521);
and U8162 (N_8162,N_2313,N_3300);
nor U8163 (N_8163,N_2006,N_2754);
nor U8164 (N_8164,N_3867,N_2906);
and U8165 (N_8165,N_1398,N_3840);
nand U8166 (N_8166,N_2821,N_4667);
and U8167 (N_8167,N_943,N_4596);
nand U8168 (N_8168,N_1056,N_469);
xnor U8169 (N_8169,N_3820,N_4006);
nor U8170 (N_8170,N_2597,N_3573);
or U8171 (N_8171,N_4836,N_2368);
and U8172 (N_8172,N_4426,N_3896);
and U8173 (N_8173,N_3520,N_90);
nand U8174 (N_8174,N_2277,N_4446);
xnor U8175 (N_8175,N_2226,N_3285);
and U8176 (N_8176,N_1276,N_1636);
and U8177 (N_8177,N_2496,N_1054);
nand U8178 (N_8178,N_2829,N_794);
and U8179 (N_8179,N_1659,N_2062);
nor U8180 (N_8180,N_4455,N_1315);
or U8181 (N_8181,N_838,N_1517);
nor U8182 (N_8182,N_884,N_115);
or U8183 (N_8183,N_2185,N_466);
nand U8184 (N_8184,N_2238,N_591);
or U8185 (N_8185,N_2097,N_1674);
xnor U8186 (N_8186,N_3811,N_1844);
or U8187 (N_8187,N_2565,N_1219);
or U8188 (N_8188,N_791,N_3024);
nor U8189 (N_8189,N_1792,N_2162);
nand U8190 (N_8190,N_1763,N_3733);
or U8191 (N_8191,N_801,N_4365);
or U8192 (N_8192,N_3243,N_1289);
nor U8193 (N_8193,N_4182,N_262);
and U8194 (N_8194,N_3095,N_2300);
xnor U8195 (N_8195,N_4536,N_3789);
or U8196 (N_8196,N_3779,N_3910);
nor U8197 (N_8197,N_375,N_3765);
or U8198 (N_8198,N_549,N_909);
and U8199 (N_8199,N_2143,N_3503);
nand U8200 (N_8200,N_3789,N_1988);
and U8201 (N_8201,N_4854,N_4480);
nand U8202 (N_8202,N_1323,N_4954);
or U8203 (N_8203,N_230,N_1046);
and U8204 (N_8204,N_2325,N_3738);
xor U8205 (N_8205,N_4533,N_871);
and U8206 (N_8206,N_4792,N_4958);
nand U8207 (N_8207,N_381,N_225);
nor U8208 (N_8208,N_1589,N_3006);
nand U8209 (N_8209,N_1038,N_4638);
and U8210 (N_8210,N_2270,N_1752);
or U8211 (N_8211,N_822,N_407);
or U8212 (N_8212,N_1164,N_1178);
and U8213 (N_8213,N_1914,N_1976);
nor U8214 (N_8214,N_1396,N_4582);
nor U8215 (N_8215,N_1477,N_3912);
and U8216 (N_8216,N_1535,N_4638);
or U8217 (N_8217,N_331,N_4061);
nand U8218 (N_8218,N_686,N_4114);
and U8219 (N_8219,N_2803,N_242);
nor U8220 (N_8220,N_2175,N_4525);
xor U8221 (N_8221,N_4101,N_2459);
nor U8222 (N_8222,N_3525,N_1079);
or U8223 (N_8223,N_2088,N_2388);
and U8224 (N_8224,N_1271,N_2867);
nand U8225 (N_8225,N_1515,N_2320);
nor U8226 (N_8226,N_1855,N_1758);
nor U8227 (N_8227,N_3272,N_4512);
or U8228 (N_8228,N_1903,N_3415);
and U8229 (N_8229,N_1004,N_3073);
and U8230 (N_8230,N_4726,N_4970);
and U8231 (N_8231,N_239,N_3209);
or U8232 (N_8232,N_3114,N_1894);
or U8233 (N_8233,N_4237,N_2983);
nor U8234 (N_8234,N_2279,N_573);
nand U8235 (N_8235,N_1867,N_2508);
or U8236 (N_8236,N_1788,N_4944);
and U8237 (N_8237,N_217,N_2434);
nand U8238 (N_8238,N_4223,N_1151);
or U8239 (N_8239,N_4675,N_2006);
or U8240 (N_8240,N_4730,N_3538);
or U8241 (N_8241,N_2547,N_2087);
and U8242 (N_8242,N_3720,N_617);
or U8243 (N_8243,N_2713,N_4371);
or U8244 (N_8244,N_4806,N_2908);
and U8245 (N_8245,N_1023,N_1187);
xnor U8246 (N_8246,N_3057,N_4718);
nor U8247 (N_8247,N_333,N_1791);
or U8248 (N_8248,N_1152,N_4444);
nand U8249 (N_8249,N_2607,N_614);
xnor U8250 (N_8250,N_2656,N_3008);
nand U8251 (N_8251,N_4133,N_4972);
nand U8252 (N_8252,N_228,N_1142);
xnor U8253 (N_8253,N_1281,N_2826);
nand U8254 (N_8254,N_1490,N_94);
and U8255 (N_8255,N_685,N_2784);
or U8256 (N_8256,N_4452,N_4058);
nand U8257 (N_8257,N_4806,N_1758);
nor U8258 (N_8258,N_2223,N_2692);
or U8259 (N_8259,N_4316,N_594);
or U8260 (N_8260,N_3485,N_3005);
or U8261 (N_8261,N_3624,N_3277);
nand U8262 (N_8262,N_1879,N_1038);
and U8263 (N_8263,N_1801,N_2670);
xor U8264 (N_8264,N_187,N_144);
or U8265 (N_8265,N_3815,N_1732);
and U8266 (N_8266,N_143,N_1984);
or U8267 (N_8267,N_4190,N_1168);
xor U8268 (N_8268,N_319,N_3893);
nand U8269 (N_8269,N_1583,N_2064);
or U8270 (N_8270,N_2058,N_3070);
nor U8271 (N_8271,N_2498,N_4050);
or U8272 (N_8272,N_428,N_4717);
nand U8273 (N_8273,N_1277,N_1042);
xor U8274 (N_8274,N_187,N_1538);
or U8275 (N_8275,N_230,N_3022);
or U8276 (N_8276,N_946,N_4154);
nand U8277 (N_8277,N_1320,N_1797);
nand U8278 (N_8278,N_4933,N_765);
or U8279 (N_8279,N_2490,N_2154);
or U8280 (N_8280,N_2155,N_3835);
and U8281 (N_8281,N_4655,N_1158);
nor U8282 (N_8282,N_2050,N_601);
nor U8283 (N_8283,N_932,N_207);
nand U8284 (N_8284,N_576,N_2983);
nor U8285 (N_8285,N_959,N_4580);
nand U8286 (N_8286,N_3966,N_4849);
or U8287 (N_8287,N_772,N_3352);
and U8288 (N_8288,N_2557,N_4148);
nand U8289 (N_8289,N_1993,N_2351);
xnor U8290 (N_8290,N_3864,N_388);
nor U8291 (N_8291,N_1338,N_1859);
and U8292 (N_8292,N_281,N_1649);
xor U8293 (N_8293,N_1816,N_859);
or U8294 (N_8294,N_1936,N_4492);
or U8295 (N_8295,N_2114,N_1831);
nor U8296 (N_8296,N_348,N_14);
or U8297 (N_8297,N_653,N_3253);
xnor U8298 (N_8298,N_3738,N_4122);
nand U8299 (N_8299,N_1570,N_437);
and U8300 (N_8300,N_179,N_2778);
or U8301 (N_8301,N_3634,N_1454);
or U8302 (N_8302,N_3852,N_4650);
nand U8303 (N_8303,N_128,N_2827);
and U8304 (N_8304,N_3507,N_4809);
nand U8305 (N_8305,N_1938,N_3720);
xor U8306 (N_8306,N_4283,N_931);
nor U8307 (N_8307,N_1773,N_789);
and U8308 (N_8308,N_3524,N_41);
and U8309 (N_8309,N_384,N_4236);
or U8310 (N_8310,N_3906,N_1926);
nor U8311 (N_8311,N_4746,N_2676);
and U8312 (N_8312,N_2335,N_4479);
nand U8313 (N_8313,N_4627,N_4155);
or U8314 (N_8314,N_2094,N_4529);
or U8315 (N_8315,N_2767,N_3263);
or U8316 (N_8316,N_863,N_3280);
and U8317 (N_8317,N_2910,N_2390);
nand U8318 (N_8318,N_3214,N_1758);
or U8319 (N_8319,N_4892,N_3256);
and U8320 (N_8320,N_1745,N_3817);
or U8321 (N_8321,N_3166,N_3786);
and U8322 (N_8322,N_2555,N_166);
nor U8323 (N_8323,N_4722,N_835);
or U8324 (N_8324,N_168,N_2468);
and U8325 (N_8325,N_1310,N_2848);
nor U8326 (N_8326,N_3768,N_2254);
nand U8327 (N_8327,N_1200,N_4854);
nand U8328 (N_8328,N_1031,N_3923);
nand U8329 (N_8329,N_4352,N_3180);
and U8330 (N_8330,N_2539,N_2085);
and U8331 (N_8331,N_3253,N_3051);
and U8332 (N_8332,N_1673,N_3744);
nor U8333 (N_8333,N_4499,N_4325);
and U8334 (N_8334,N_2173,N_4947);
nand U8335 (N_8335,N_3460,N_1967);
or U8336 (N_8336,N_474,N_2530);
or U8337 (N_8337,N_4254,N_2404);
nor U8338 (N_8338,N_3998,N_1920);
or U8339 (N_8339,N_4344,N_2531);
and U8340 (N_8340,N_1802,N_409);
nor U8341 (N_8341,N_4562,N_2985);
nor U8342 (N_8342,N_1037,N_4254);
or U8343 (N_8343,N_579,N_2898);
nand U8344 (N_8344,N_3206,N_953);
nor U8345 (N_8345,N_2064,N_542);
or U8346 (N_8346,N_3638,N_3838);
xor U8347 (N_8347,N_3028,N_4943);
nand U8348 (N_8348,N_1813,N_454);
nand U8349 (N_8349,N_4917,N_3450);
nor U8350 (N_8350,N_2526,N_3179);
nor U8351 (N_8351,N_1688,N_206);
nand U8352 (N_8352,N_1188,N_4649);
xnor U8353 (N_8353,N_704,N_325);
xnor U8354 (N_8354,N_4020,N_703);
nand U8355 (N_8355,N_3739,N_502);
or U8356 (N_8356,N_3266,N_1618);
nand U8357 (N_8357,N_4446,N_3709);
nand U8358 (N_8358,N_2500,N_505);
or U8359 (N_8359,N_4723,N_3997);
or U8360 (N_8360,N_1677,N_647);
and U8361 (N_8361,N_4101,N_3911);
nand U8362 (N_8362,N_2585,N_815);
nor U8363 (N_8363,N_1222,N_4924);
and U8364 (N_8364,N_33,N_2860);
or U8365 (N_8365,N_44,N_75);
nand U8366 (N_8366,N_4792,N_4225);
nand U8367 (N_8367,N_838,N_2318);
nand U8368 (N_8368,N_855,N_2331);
nor U8369 (N_8369,N_2654,N_4749);
or U8370 (N_8370,N_2207,N_1291);
nor U8371 (N_8371,N_629,N_2550);
xor U8372 (N_8372,N_2830,N_98);
xor U8373 (N_8373,N_509,N_1994);
or U8374 (N_8374,N_810,N_4483);
nor U8375 (N_8375,N_1308,N_3170);
or U8376 (N_8376,N_843,N_4547);
nand U8377 (N_8377,N_3524,N_357);
xnor U8378 (N_8378,N_2395,N_2495);
nand U8379 (N_8379,N_3097,N_4896);
and U8380 (N_8380,N_3216,N_1614);
and U8381 (N_8381,N_4560,N_3249);
nand U8382 (N_8382,N_2517,N_1980);
and U8383 (N_8383,N_4091,N_1008);
or U8384 (N_8384,N_2211,N_4304);
or U8385 (N_8385,N_664,N_1932);
nand U8386 (N_8386,N_4436,N_3831);
nor U8387 (N_8387,N_4232,N_2334);
or U8388 (N_8388,N_2068,N_2761);
or U8389 (N_8389,N_328,N_1669);
nand U8390 (N_8390,N_3580,N_3009);
or U8391 (N_8391,N_538,N_2478);
and U8392 (N_8392,N_999,N_4726);
nand U8393 (N_8393,N_3087,N_686);
and U8394 (N_8394,N_2350,N_2477);
and U8395 (N_8395,N_1097,N_449);
or U8396 (N_8396,N_3051,N_625);
nor U8397 (N_8397,N_1022,N_993);
and U8398 (N_8398,N_4276,N_130);
nand U8399 (N_8399,N_3802,N_2951);
and U8400 (N_8400,N_3330,N_2982);
xor U8401 (N_8401,N_446,N_2660);
xnor U8402 (N_8402,N_2596,N_4333);
nand U8403 (N_8403,N_1383,N_1006);
or U8404 (N_8404,N_3728,N_565);
nor U8405 (N_8405,N_1928,N_2445);
or U8406 (N_8406,N_3831,N_1510);
and U8407 (N_8407,N_1410,N_2976);
and U8408 (N_8408,N_3909,N_2561);
nor U8409 (N_8409,N_2675,N_3177);
nor U8410 (N_8410,N_2698,N_528);
nor U8411 (N_8411,N_2147,N_4171);
nand U8412 (N_8412,N_2307,N_2545);
nor U8413 (N_8413,N_3856,N_1944);
nand U8414 (N_8414,N_1374,N_997);
xor U8415 (N_8415,N_1035,N_1169);
or U8416 (N_8416,N_2101,N_2710);
or U8417 (N_8417,N_4808,N_4653);
nor U8418 (N_8418,N_2035,N_4503);
or U8419 (N_8419,N_3418,N_91);
or U8420 (N_8420,N_1353,N_1764);
or U8421 (N_8421,N_3911,N_326);
nor U8422 (N_8422,N_984,N_3771);
nand U8423 (N_8423,N_2656,N_4069);
nand U8424 (N_8424,N_102,N_3180);
nor U8425 (N_8425,N_357,N_3103);
and U8426 (N_8426,N_4274,N_4670);
and U8427 (N_8427,N_2382,N_2872);
and U8428 (N_8428,N_3740,N_3528);
and U8429 (N_8429,N_2518,N_4414);
or U8430 (N_8430,N_3465,N_2280);
and U8431 (N_8431,N_1012,N_442);
and U8432 (N_8432,N_1960,N_1186);
xnor U8433 (N_8433,N_1003,N_2737);
or U8434 (N_8434,N_3237,N_3477);
nor U8435 (N_8435,N_2262,N_1063);
xor U8436 (N_8436,N_3839,N_2230);
nor U8437 (N_8437,N_1683,N_2998);
or U8438 (N_8438,N_4668,N_2563);
xnor U8439 (N_8439,N_2472,N_1302);
and U8440 (N_8440,N_542,N_834);
nor U8441 (N_8441,N_4621,N_452);
or U8442 (N_8442,N_150,N_3649);
nor U8443 (N_8443,N_4686,N_4192);
or U8444 (N_8444,N_4544,N_426);
nand U8445 (N_8445,N_747,N_2996);
nor U8446 (N_8446,N_4126,N_4379);
nor U8447 (N_8447,N_4827,N_4829);
xor U8448 (N_8448,N_4590,N_3633);
nand U8449 (N_8449,N_380,N_3489);
nor U8450 (N_8450,N_1625,N_800);
nand U8451 (N_8451,N_4849,N_1211);
nand U8452 (N_8452,N_3962,N_2601);
nand U8453 (N_8453,N_2758,N_2333);
or U8454 (N_8454,N_3232,N_694);
nand U8455 (N_8455,N_72,N_1620);
nor U8456 (N_8456,N_247,N_2579);
or U8457 (N_8457,N_3384,N_4627);
and U8458 (N_8458,N_142,N_1693);
and U8459 (N_8459,N_284,N_3881);
nor U8460 (N_8460,N_3924,N_658);
nand U8461 (N_8461,N_1544,N_3606);
and U8462 (N_8462,N_336,N_1839);
or U8463 (N_8463,N_3590,N_3283);
nor U8464 (N_8464,N_428,N_2065);
nand U8465 (N_8465,N_1044,N_4343);
or U8466 (N_8466,N_377,N_1731);
and U8467 (N_8467,N_1270,N_4541);
or U8468 (N_8468,N_1521,N_4081);
or U8469 (N_8469,N_135,N_2359);
nand U8470 (N_8470,N_3173,N_293);
and U8471 (N_8471,N_4621,N_4065);
nor U8472 (N_8472,N_1888,N_178);
xor U8473 (N_8473,N_4713,N_3040);
and U8474 (N_8474,N_2708,N_2425);
xnor U8475 (N_8475,N_3106,N_903);
and U8476 (N_8476,N_408,N_2070);
nor U8477 (N_8477,N_2036,N_4324);
nor U8478 (N_8478,N_1624,N_1463);
and U8479 (N_8479,N_1611,N_3861);
nand U8480 (N_8480,N_4061,N_4396);
nand U8481 (N_8481,N_3446,N_344);
and U8482 (N_8482,N_3503,N_4265);
nand U8483 (N_8483,N_390,N_1552);
and U8484 (N_8484,N_3273,N_2382);
nor U8485 (N_8485,N_4723,N_177);
nand U8486 (N_8486,N_4006,N_4033);
and U8487 (N_8487,N_4286,N_2730);
and U8488 (N_8488,N_3747,N_985);
or U8489 (N_8489,N_4952,N_1533);
nand U8490 (N_8490,N_2008,N_703);
nand U8491 (N_8491,N_3539,N_1912);
xor U8492 (N_8492,N_1450,N_1654);
nor U8493 (N_8493,N_449,N_1263);
nand U8494 (N_8494,N_1040,N_2753);
nand U8495 (N_8495,N_355,N_4888);
nand U8496 (N_8496,N_2552,N_3238);
nor U8497 (N_8497,N_2508,N_4993);
nand U8498 (N_8498,N_2833,N_3036);
nor U8499 (N_8499,N_908,N_3426);
nor U8500 (N_8500,N_408,N_1127);
xor U8501 (N_8501,N_89,N_1043);
nand U8502 (N_8502,N_4603,N_638);
or U8503 (N_8503,N_567,N_332);
nand U8504 (N_8504,N_3894,N_2152);
and U8505 (N_8505,N_3973,N_3473);
and U8506 (N_8506,N_2550,N_4673);
nand U8507 (N_8507,N_4886,N_4096);
or U8508 (N_8508,N_4613,N_1678);
nand U8509 (N_8509,N_803,N_4861);
nand U8510 (N_8510,N_1133,N_2307);
and U8511 (N_8511,N_4502,N_3894);
nor U8512 (N_8512,N_2920,N_3110);
nand U8513 (N_8513,N_2004,N_1995);
nand U8514 (N_8514,N_3910,N_4042);
and U8515 (N_8515,N_351,N_3384);
xor U8516 (N_8516,N_4785,N_4295);
or U8517 (N_8517,N_584,N_902);
and U8518 (N_8518,N_1115,N_3140);
nor U8519 (N_8519,N_4080,N_1960);
and U8520 (N_8520,N_4028,N_4932);
nand U8521 (N_8521,N_4827,N_1830);
nor U8522 (N_8522,N_3558,N_1814);
nand U8523 (N_8523,N_3586,N_3739);
xnor U8524 (N_8524,N_3395,N_3565);
or U8525 (N_8525,N_3300,N_4768);
nand U8526 (N_8526,N_827,N_4370);
or U8527 (N_8527,N_1421,N_1350);
nand U8528 (N_8528,N_2532,N_2221);
and U8529 (N_8529,N_3442,N_1181);
nor U8530 (N_8530,N_455,N_1886);
and U8531 (N_8531,N_3231,N_1560);
nor U8532 (N_8532,N_4455,N_2183);
xor U8533 (N_8533,N_4317,N_3585);
nand U8534 (N_8534,N_1778,N_3492);
and U8535 (N_8535,N_325,N_2922);
nand U8536 (N_8536,N_1613,N_3643);
and U8537 (N_8537,N_2183,N_400);
nand U8538 (N_8538,N_4853,N_1706);
xor U8539 (N_8539,N_1087,N_1337);
nand U8540 (N_8540,N_2732,N_1188);
nor U8541 (N_8541,N_2404,N_4138);
nor U8542 (N_8542,N_4138,N_4783);
nand U8543 (N_8543,N_2805,N_1994);
nor U8544 (N_8544,N_2768,N_4565);
or U8545 (N_8545,N_206,N_1710);
or U8546 (N_8546,N_1079,N_3741);
nor U8547 (N_8547,N_2189,N_4349);
and U8548 (N_8548,N_2031,N_4814);
nor U8549 (N_8549,N_3011,N_4570);
or U8550 (N_8550,N_2743,N_4430);
nand U8551 (N_8551,N_2807,N_2696);
or U8552 (N_8552,N_1028,N_691);
or U8553 (N_8553,N_2778,N_3802);
or U8554 (N_8554,N_2128,N_3299);
nor U8555 (N_8555,N_2319,N_2847);
nand U8556 (N_8556,N_4480,N_195);
nand U8557 (N_8557,N_608,N_3970);
nand U8558 (N_8558,N_3038,N_4875);
or U8559 (N_8559,N_4255,N_2034);
and U8560 (N_8560,N_3459,N_3969);
or U8561 (N_8561,N_4664,N_167);
nand U8562 (N_8562,N_2745,N_2151);
nor U8563 (N_8563,N_2713,N_733);
nand U8564 (N_8564,N_1703,N_3746);
and U8565 (N_8565,N_1094,N_996);
and U8566 (N_8566,N_4234,N_4549);
and U8567 (N_8567,N_2550,N_4246);
and U8568 (N_8568,N_3642,N_1665);
and U8569 (N_8569,N_2761,N_1668);
or U8570 (N_8570,N_870,N_2570);
nand U8571 (N_8571,N_4491,N_4927);
and U8572 (N_8572,N_1942,N_1581);
or U8573 (N_8573,N_1170,N_3570);
or U8574 (N_8574,N_226,N_585);
and U8575 (N_8575,N_2651,N_2461);
or U8576 (N_8576,N_990,N_750);
xnor U8577 (N_8577,N_745,N_4261);
nand U8578 (N_8578,N_155,N_3575);
and U8579 (N_8579,N_4647,N_3638);
and U8580 (N_8580,N_249,N_4104);
nand U8581 (N_8581,N_2219,N_4677);
nor U8582 (N_8582,N_4261,N_1414);
or U8583 (N_8583,N_4868,N_4612);
and U8584 (N_8584,N_1392,N_3626);
xor U8585 (N_8585,N_4186,N_2945);
or U8586 (N_8586,N_4120,N_3862);
or U8587 (N_8587,N_3248,N_2428);
and U8588 (N_8588,N_290,N_4923);
nor U8589 (N_8589,N_1647,N_3825);
and U8590 (N_8590,N_2927,N_2930);
nand U8591 (N_8591,N_396,N_1598);
nand U8592 (N_8592,N_4706,N_2240);
nor U8593 (N_8593,N_1031,N_716);
nor U8594 (N_8594,N_43,N_1276);
nor U8595 (N_8595,N_4738,N_4065);
or U8596 (N_8596,N_4946,N_1365);
and U8597 (N_8597,N_2548,N_1066);
and U8598 (N_8598,N_1207,N_3109);
xor U8599 (N_8599,N_3185,N_4297);
xnor U8600 (N_8600,N_4456,N_3935);
or U8601 (N_8601,N_4093,N_1072);
and U8602 (N_8602,N_1289,N_3656);
or U8603 (N_8603,N_3042,N_3633);
nand U8604 (N_8604,N_715,N_3566);
nor U8605 (N_8605,N_181,N_4676);
nand U8606 (N_8606,N_1210,N_37);
nand U8607 (N_8607,N_4631,N_1136);
or U8608 (N_8608,N_4269,N_3249);
and U8609 (N_8609,N_2704,N_2085);
nor U8610 (N_8610,N_3164,N_1538);
or U8611 (N_8611,N_336,N_3381);
and U8612 (N_8612,N_2832,N_2172);
xor U8613 (N_8613,N_2856,N_2503);
and U8614 (N_8614,N_3527,N_3246);
and U8615 (N_8615,N_1211,N_2417);
nand U8616 (N_8616,N_443,N_1983);
nand U8617 (N_8617,N_335,N_2093);
or U8618 (N_8618,N_3086,N_62);
nor U8619 (N_8619,N_3107,N_4487);
nand U8620 (N_8620,N_1452,N_3089);
nand U8621 (N_8621,N_3169,N_2703);
or U8622 (N_8622,N_4222,N_2176);
xnor U8623 (N_8623,N_1307,N_1284);
or U8624 (N_8624,N_4415,N_3995);
nor U8625 (N_8625,N_672,N_1536);
and U8626 (N_8626,N_3855,N_4585);
or U8627 (N_8627,N_435,N_2919);
nor U8628 (N_8628,N_283,N_50);
nor U8629 (N_8629,N_2397,N_451);
xnor U8630 (N_8630,N_250,N_1584);
nand U8631 (N_8631,N_343,N_2602);
nor U8632 (N_8632,N_3409,N_661);
and U8633 (N_8633,N_895,N_2077);
and U8634 (N_8634,N_2793,N_2805);
and U8635 (N_8635,N_3878,N_4675);
or U8636 (N_8636,N_2834,N_461);
or U8637 (N_8637,N_4000,N_996);
nor U8638 (N_8638,N_804,N_4252);
xnor U8639 (N_8639,N_201,N_4781);
or U8640 (N_8640,N_1351,N_4469);
nor U8641 (N_8641,N_379,N_1955);
and U8642 (N_8642,N_4530,N_4870);
nand U8643 (N_8643,N_1130,N_4163);
nor U8644 (N_8644,N_3794,N_4271);
nor U8645 (N_8645,N_472,N_205);
and U8646 (N_8646,N_737,N_1611);
and U8647 (N_8647,N_1941,N_1749);
nor U8648 (N_8648,N_684,N_2280);
and U8649 (N_8649,N_1809,N_658);
or U8650 (N_8650,N_492,N_1003);
nor U8651 (N_8651,N_434,N_3951);
and U8652 (N_8652,N_3788,N_3696);
nor U8653 (N_8653,N_4449,N_4693);
and U8654 (N_8654,N_300,N_2920);
and U8655 (N_8655,N_1601,N_589);
nand U8656 (N_8656,N_4628,N_4633);
nor U8657 (N_8657,N_671,N_2298);
nor U8658 (N_8658,N_4876,N_1535);
nand U8659 (N_8659,N_2164,N_1444);
nor U8660 (N_8660,N_4251,N_4704);
nand U8661 (N_8661,N_529,N_3265);
nand U8662 (N_8662,N_3144,N_1769);
nor U8663 (N_8663,N_3182,N_4577);
xnor U8664 (N_8664,N_2584,N_2803);
nand U8665 (N_8665,N_434,N_4448);
or U8666 (N_8666,N_4189,N_4736);
and U8667 (N_8667,N_3383,N_2503);
and U8668 (N_8668,N_295,N_4987);
nand U8669 (N_8669,N_1715,N_2990);
xor U8670 (N_8670,N_2208,N_2505);
and U8671 (N_8671,N_155,N_3719);
nor U8672 (N_8672,N_2274,N_4245);
nor U8673 (N_8673,N_3037,N_833);
or U8674 (N_8674,N_1152,N_3736);
or U8675 (N_8675,N_4162,N_2240);
nor U8676 (N_8676,N_1126,N_2793);
xor U8677 (N_8677,N_97,N_3124);
or U8678 (N_8678,N_1071,N_7);
nand U8679 (N_8679,N_1150,N_4296);
and U8680 (N_8680,N_4950,N_3901);
nand U8681 (N_8681,N_2258,N_2867);
nor U8682 (N_8682,N_1818,N_4252);
nor U8683 (N_8683,N_2149,N_199);
nand U8684 (N_8684,N_225,N_4676);
or U8685 (N_8685,N_1645,N_1004);
nor U8686 (N_8686,N_4935,N_545);
nand U8687 (N_8687,N_3923,N_2461);
and U8688 (N_8688,N_3938,N_2353);
or U8689 (N_8689,N_1701,N_2691);
nand U8690 (N_8690,N_1633,N_223);
nor U8691 (N_8691,N_3264,N_1446);
and U8692 (N_8692,N_2762,N_722);
and U8693 (N_8693,N_3326,N_1901);
and U8694 (N_8694,N_191,N_560);
and U8695 (N_8695,N_4651,N_1709);
nand U8696 (N_8696,N_2759,N_4684);
and U8697 (N_8697,N_4717,N_1408);
and U8698 (N_8698,N_4730,N_2556);
and U8699 (N_8699,N_2025,N_2745);
nand U8700 (N_8700,N_3618,N_3616);
nor U8701 (N_8701,N_2241,N_4095);
nand U8702 (N_8702,N_1265,N_478);
nor U8703 (N_8703,N_1079,N_3201);
nor U8704 (N_8704,N_2243,N_2598);
and U8705 (N_8705,N_4102,N_2957);
nand U8706 (N_8706,N_1995,N_4651);
and U8707 (N_8707,N_288,N_3549);
or U8708 (N_8708,N_3921,N_3556);
and U8709 (N_8709,N_4609,N_825);
nand U8710 (N_8710,N_938,N_1924);
and U8711 (N_8711,N_1673,N_3809);
nand U8712 (N_8712,N_3642,N_566);
or U8713 (N_8713,N_2963,N_1187);
nand U8714 (N_8714,N_4651,N_3446);
and U8715 (N_8715,N_877,N_3020);
or U8716 (N_8716,N_4417,N_374);
nand U8717 (N_8717,N_117,N_3942);
or U8718 (N_8718,N_3534,N_3802);
and U8719 (N_8719,N_4542,N_4080);
xnor U8720 (N_8720,N_1050,N_4225);
nand U8721 (N_8721,N_1340,N_482);
nor U8722 (N_8722,N_2701,N_3263);
xnor U8723 (N_8723,N_4846,N_2207);
nor U8724 (N_8724,N_3934,N_3753);
nor U8725 (N_8725,N_1490,N_4082);
and U8726 (N_8726,N_157,N_162);
or U8727 (N_8727,N_2221,N_1462);
or U8728 (N_8728,N_300,N_2082);
and U8729 (N_8729,N_1197,N_3693);
or U8730 (N_8730,N_3045,N_592);
or U8731 (N_8731,N_4298,N_3733);
xor U8732 (N_8732,N_1669,N_4257);
or U8733 (N_8733,N_179,N_4388);
nor U8734 (N_8734,N_1520,N_231);
and U8735 (N_8735,N_2259,N_3589);
xnor U8736 (N_8736,N_2551,N_2390);
and U8737 (N_8737,N_2717,N_712);
nor U8738 (N_8738,N_3513,N_2112);
nor U8739 (N_8739,N_3948,N_2778);
or U8740 (N_8740,N_4077,N_536);
or U8741 (N_8741,N_4925,N_740);
nand U8742 (N_8742,N_4490,N_217);
and U8743 (N_8743,N_3968,N_14);
nand U8744 (N_8744,N_3938,N_4121);
nand U8745 (N_8745,N_1945,N_3897);
or U8746 (N_8746,N_3314,N_4213);
nor U8747 (N_8747,N_522,N_1489);
and U8748 (N_8748,N_2856,N_1533);
and U8749 (N_8749,N_4313,N_70);
or U8750 (N_8750,N_2647,N_4959);
and U8751 (N_8751,N_332,N_1164);
or U8752 (N_8752,N_170,N_4736);
and U8753 (N_8753,N_4837,N_4014);
or U8754 (N_8754,N_570,N_1110);
and U8755 (N_8755,N_1272,N_4662);
and U8756 (N_8756,N_3244,N_2939);
nor U8757 (N_8757,N_4733,N_1183);
nand U8758 (N_8758,N_2265,N_531);
nor U8759 (N_8759,N_1009,N_3062);
or U8760 (N_8760,N_4481,N_880);
nand U8761 (N_8761,N_4300,N_2942);
or U8762 (N_8762,N_2359,N_4691);
xor U8763 (N_8763,N_3117,N_4824);
and U8764 (N_8764,N_284,N_3998);
nand U8765 (N_8765,N_2990,N_1503);
nand U8766 (N_8766,N_989,N_1085);
and U8767 (N_8767,N_1205,N_730);
nor U8768 (N_8768,N_650,N_3768);
and U8769 (N_8769,N_4066,N_661);
nand U8770 (N_8770,N_3756,N_2359);
nand U8771 (N_8771,N_3465,N_3428);
or U8772 (N_8772,N_2845,N_3382);
nand U8773 (N_8773,N_2331,N_1203);
nand U8774 (N_8774,N_362,N_764);
or U8775 (N_8775,N_4047,N_861);
nor U8776 (N_8776,N_463,N_2337);
and U8777 (N_8777,N_433,N_4839);
nand U8778 (N_8778,N_871,N_3915);
or U8779 (N_8779,N_4327,N_4799);
nand U8780 (N_8780,N_3344,N_4147);
and U8781 (N_8781,N_2074,N_1171);
nor U8782 (N_8782,N_3766,N_3707);
xnor U8783 (N_8783,N_2428,N_163);
and U8784 (N_8784,N_3712,N_3514);
nor U8785 (N_8785,N_1808,N_3433);
and U8786 (N_8786,N_2673,N_2969);
and U8787 (N_8787,N_1763,N_1611);
xor U8788 (N_8788,N_565,N_2848);
and U8789 (N_8789,N_4336,N_2156);
nor U8790 (N_8790,N_505,N_4770);
nand U8791 (N_8791,N_2934,N_4420);
xnor U8792 (N_8792,N_3005,N_1542);
nand U8793 (N_8793,N_4770,N_4339);
nor U8794 (N_8794,N_4430,N_3814);
xnor U8795 (N_8795,N_3340,N_4833);
xnor U8796 (N_8796,N_1834,N_3774);
nor U8797 (N_8797,N_4904,N_3827);
xor U8798 (N_8798,N_2233,N_4244);
nand U8799 (N_8799,N_1872,N_4021);
xor U8800 (N_8800,N_365,N_1915);
or U8801 (N_8801,N_374,N_280);
nand U8802 (N_8802,N_1601,N_3458);
nand U8803 (N_8803,N_3679,N_2485);
nand U8804 (N_8804,N_153,N_1511);
nor U8805 (N_8805,N_1924,N_2514);
or U8806 (N_8806,N_1142,N_1813);
or U8807 (N_8807,N_1888,N_4988);
nor U8808 (N_8808,N_1278,N_4650);
nand U8809 (N_8809,N_471,N_2562);
nand U8810 (N_8810,N_1418,N_277);
or U8811 (N_8811,N_4692,N_2953);
nor U8812 (N_8812,N_747,N_2146);
and U8813 (N_8813,N_695,N_4515);
nor U8814 (N_8814,N_1449,N_4187);
or U8815 (N_8815,N_672,N_4437);
and U8816 (N_8816,N_4468,N_1890);
nor U8817 (N_8817,N_2974,N_4607);
or U8818 (N_8818,N_4479,N_2146);
and U8819 (N_8819,N_1200,N_3928);
or U8820 (N_8820,N_1986,N_2840);
and U8821 (N_8821,N_1732,N_1656);
or U8822 (N_8822,N_4059,N_877);
xnor U8823 (N_8823,N_4186,N_295);
and U8824 (N_8824,N_4882,N_4390);
or U8825 (N_8825,N_2755,N_103);
nor U8826 (N_8826,N_1819,N_2311);
nand U8827 (N_8827,N_551,N_3663);
or U8828 (N_8828,N_3037,N_4498);
or U8829 (N_8829,N_3358,N_2073);
or U8830 (N_8830,N_1393,N_3045);
and U8831 (N_8831,N_830,N_1400);
nor U8832 (N_8832,N_272,N_1746);
or U8833 (N_8833,N_4693,N_3839);
and U8834 (N_8834,N_17,N_4355);
or U8835 (N_8835,N_4055,N_4456);
and U8836 (N_8836,N_4803,N_4420);
and U8837 (N_8837,N_4635,N_3365);
nor U8838 (N_8838,N_426,N_1835);
nor U8839 (N_8839,N_1776,N_4604);
nor U8840 (N_8840,N_1574,N_4374);
nor U8841 (N_8841,N_2080,N_2990);
nand U8842 (N_8842,N_1137,N_2388);
xor U8843 (N_8843,N_180,N_2546);
nand U8844 (N_8844,N_3933,N_716);
and U8845 (N_8845,N_4847,N_3181);
nor U8846 (N_8846,N_2599,N_839);
xnor U8847 (N_8847,N_3249,N_1437);
and U8848 (N_8848,N_3491,N_3918);
and U8849 (N_8849,N_1103,N_2635);
nand U8850 (N_8850,N_2153,N_1757);
nor U8851 (N_8851,N_3068,N_1050);
and U8852 (N_8852,N_1488,N_2680);
or U8853 (N_8853,N_3684,N_3171);
nor U8854 (N_8854,N_4399,N_2192);
and U8855 (N_8855,N_1047,N_1953);
nor U8856 (N_8856,N_1716,N_3677);
nor U8857 (N_8857,N_1703,N_4989);
or U8858 (N_8858,N_4605,N_2584);
nand U8859 (N_8859,N_2700,N_18);
or U8860 (N_8860,N_110,N_2378);
or U8861 (N_8861,N_967,N_2365);
and U8862 (N_8862,N_3749,N_844);
nand U8863 (N_8863,N_4614,N_3994);
or U8864 (N_8864,N_354,N_403);
nand U8865 (N_8865,N_4709,N_493);
nand U8866 (N_8866,N_1494,N_4957);
nand U8867 (N_8867,N_3933,N_1103);
or U8868 (N_8868,N_774,N_3402);
or U8869 (N_8869,N_4554,N_1088);
or U8870 (N_8870,N_1143,N_2475);
nand U8871 (N_8871,N_1324,N_3326);
and U8872 (N_8872,N_2241,N_1723);
xor U8873 (N_8873,N_2069,N_1090);
nand U8874 (N_8874,N_1386,N_605);
or U8875 (N_8875,N_181,N_4026);
xor U8876 (N_8876,N_4541,N_3778);
nor U8877 (N_8877,N_2671,N_2666);
and U8878 (N_8878,N_4396,N_4355);
nand U8879 (N_8879,N_1324,N_3091);
nand U8880 (N_8880,N_2124,N_2947);
nand U8881 (N_8881,N_2501,N_9);
nand U8882 (N_8882,N_3846,N_1856);
and U8883 (N_8883,N_2883,N_4910);
or U8884 (N_8884,N_116,N_2794);
nor U8885 (N_8885,N_4589,N_4376);
and U8886 (N_8886,N_3465,N_251);
or U8887 (N_8887,N_4106,N_773);
or U8888 (N_8888,N_232,N_3802);
and U8889 (N_8889,N_112,N_4351);
or U8890 (N_8890,N_4840,N_13);
nand U8891 (N_8891,N_1915,N_230);
or U8892 (N_8892,N_3877,N_3968);
and U8893 (N_8893,N_3631,N_2335);
and U8894 (N_8894,N_3026,N_3471);
nor U8895 (N_8895,N_355,N_2473);
or U8896 (N_8896,N_3817,N_4177);
xnor U8897 (N_8897,N_536,N_934);
nor U8898 (N_8898,N_318,N_915);
nor U8899 (N_8899,N_4008,N_766);
nor U8900 (N_8900,N_2509,N_4139);
or U8901 (N_8901,N_980,N_4148);
nand U8902 (N_8902,N_4592,N_3330);
nor U8903 (N_8903,N_4775,N_4400);
or U8904 (N_8904,N_2615,N_1901);
nand U8905 (N_8905,N_1838,N_2153);
nor U8906 (N_8906,N_4114,N_1416);
or U8907 (N_8907,N_3578,N_4943);
xor U8908 (N_8908,N_3760,N_3974);
nand U8909 (N_8909,N_2006,N_398);
and U8910 (N_8910,N_666,N_4438);
nor U8911 (N_8911,N_3224,N_2476);
nor U8912 (N_8912,N_2103,N_1498);
or U8913 (N_8913,N_3375,N_4995);
or U8914 (N_8914,N_3942,N_4322);
nand U8915 (N_8915,N_1504,N_1192);
or U8916 (N_8916,N_4258,N_1903);
xnor U8917 (N_8917,N_4885,N_1891);
nor U8918 (N_8918,N_3061,N_905);
nor U8919 (N_8919,N_216,N_2929);
or U8920 (N_8920,N_153,N_3677);
nor U8921 (N_8921,N_1260,N_452);
and U8922 (N_8922,N_939,N_3096);
nand U8923 (N_8923,N_204,N_4954);
or U8924 (N_8924,N_4301,N_1144);
nand U8925 (N_8925,N_4457,N_4592);
xnor U8926 (N_8926,N_919,N_3274);
or U8927 (N_8927,N_2373,N_609);
nor U8928 (N_8928,N_4076,N_2563);
nand U8929 (N_8929,N_4217,N_987);
nand U8930 (N_8930,N_3196,N_781);
xnor U8931 (N_8931,N_4274,N_1773);
or U8932 (N_8932,N_350,N_1596);
and U8933 (N_8933,N_3375,N_4014);
and U8934 (N_8934,N_340,N_4434);
or U8935 (N_8935,N_1648,N_2122);
nor U8936 (N_8936,N_2670,N_3159);
xnor U8937 (N_8937,N_1249,N_725);
nand U8938 (N_8938,N_3652,N_4683);
or U8939 (N_8939,N_258,N_3731);
and U8940 (N_8940,N_2223,N_969);
nor U8941 (N_8941,N_1997,N_1932);
or U8942 (N_8942,N_4708,N_4063);
nor U8943 (N_8943,N_1069,N_4058);
nor U8944 (N_8944,N_1931,N_1953);
nor U8945 (N_8945,N_35,N_3452);
xnor U8946 (N_8946,N_303,N_4517);
or U8947 (N_8947,N_44,N_1842);
nand U8948 (N_8948,N_3944,N_104);
nor U8949 (N_8949,N_1860,N_4236);
nand U8950 (N_8950,N_1596,N_4020);
nor U8951 (N_8951,N_1214,N_2036);
or U8952 (N_8952,N_2015,N_2273);
nand U8953 (N_8953,N_4903,N_2070);
nand U8954 (N_8954,N_4368,N_4972);
and U8955 (N_8955,N_1623,N_3655);
or U8956 (N_8956,N_40,N_3504);
nor U8957 (N_8957,N_4146,N_4957);
or U8958 (N_8958,N_1168,N_631);
and U8959 (N_8959,N_2828,N_1016);
and U8960 (N_8960,N_3493,N_2416);
nor U8961 (N_8961,N_3925,N_1159);
and U8962 (N_8962,N_3041,N_3675);
nor U8963 (N_8963,N_3156,N_4393);
nand U8964 (N_8964,N_2357,N_2982);
nor U8965 (N_8965,N_724,N_1060);
and U8966 (N_8966,N_255,N_4711);
or U8967 (N_8967,N_4690,N_610);
nand U8968 (N_8968,N_2032,N_1556);
nor U8969 (N_8969,N_4486,N_1457);
and U8970 (N_8970,N_140,N_4057);
xnor U8971 (N_8971,N_742,N_2981);
or U8972 (N_8972,N_4520,N_4084);
and U8973 (N_8973,N_4278,N_1094);
nand U8974 (N_8974,N_4484,N_746);
xnor U8975 (N_8975,N_409,N_2532);
nor U8976 (N_8976,N_647,N_2274);
nand U8977 (N_8977,N_1157,N_3896);
nor U8978 (N_8978,N_586,N_1356);
nor U8979 (N_8979,N_1521,N_4895);
nand U8980 (N_8980,N_3173,N_2235);
nand U8981 (N_8981,N_1945,N_230);
nand U8982 (N_8982,N_2009,N_2654);
or U8983 (N_8983,N_3634,N_2767);
and U8984 (N_8984,N_821,N_1300);
or U8985 (N_8985,N_230,N_3518);
and U8986 (N_8986,N_1185,N_4234);
or U8987 (N_8987,N_4850,N_861);
nand U8988 (N_8988,N_912,N_4156);
and U8989 (N_8989,N_1955,N_1449);
or U8990 (N_8990,N_2008,N_1612);
or U8991 (N_8991,N_1693,N_2450);
nor U8992 (N_8992,N_1640,N_4077);
nor U8993 (N_8993,N_181,N_3868);
and U8994 (N_8994,N_4640,N_2814);
or U8995 (N_8995,N_255,N_1465);
nor U8996 (N_8996,N_2137,N_4104);
or U8997 (N_8997,N_4884,N_1270);
nand U8998 (N_8998,N_1447,N_3186);
nand U8999 (N_8999,N_3416,N_1658);
nor U9000 (N_9000,N_882,N_764);
nand U9001 (N_9001,N_820,N_4186);
or U9002 (N_9002,N_3246,N_2540);
and U9003 (N_9003,N_574,N_1400);
nand U9004 (N_9004,N_205,N_4013);
nor U9005 (N_9005,N_228,N_1774);
nor U9006 (N_9006,N_445,N_4678);
and U9007 (N_9007,N_3520,N_3869);
or U9008 (N_9008,N_4424,N_567);
nor U9009 (N_9009,N_2051,N_1176);
and U9010 (N_9010,N_2940,N_1257);
nor U9011 (N_9011,N_4438,N_2894);
and U9012 (N_9012,N_2086,N_1283);
xor U9013 (N_9013,N_2320,N_497);
nand U9014 (N_9014,N_1596,N_3721);
and U9015 (N_9015,N_3379,N_1551);
and U9016 (N_9016,N_618,N_2676);
or U9017 (N_9017,N_1303,N_1925);
or U9018 (N_9018,N_1191,N_270);
and U9019 (N_9019,N_4460,N_1544);
nand U9020 (N_9020,N_1314,N_4640);
xor U9021 (N_9021,N_4181,N_1780);
or U9022 (N_9022,N_4741,N_384);
nand U9023 (N_9023,N_3215,N_1330);
nor U9024 (N_9024,N_551,N_77);
nor U9025 (N_9025,N_4226,N_4344);
nor U9026 (N_9026,N_4417,N_1424);
nor U9027 (N_9027,N_460,N_990);
nand U9028 (N_9028,N_4959,N_3306);
or U9029 (N_9029,N_521,N_3370);
and U9030 (N_9030,N_2659,N_395);
and U9031 (N_9031,N_1303,N_1339);
nor U9032 (N_9032,N_1928,N_3624);
and U9033 (N_9033,N_3,N_1788);
xnor U9034 (N_9034,N_3667,N_2277);
or U9035 (N_9035,N_2483,N_1945);
nor U9036 (N_9036,N_658,N_1855);
and U9037 (N_9037,N_2248,N_3625);
and U9038 (N_9038,N_614,N_1089);
or U9039 (N_9039,N_753,N_4911);
and U9040 (N_9040,N_3131,N_2484);
or U9041 (N_9041,N_67,N_1654);
nor U9042 (N_9042,N_4510,N_4063);
nor U9043 (N_9043,N_3505,N_226);
nor U9044 (N_9044,N_4118,N_1636);
xnor U9045 (N_9045,N_1394,N_632);
or U9046 (N_9046,N_4217,N_3736);
nor U9047 (N_9047,N_2019,N_1398);
xor U9048 (N_9048,N_65,N_2229);
nand U9049 (N_9049,N_2057,N_1718);
or U9050 (N_9050,N_1278,N_1847);
and U9051 (N_9051,N_3450,N_2933);
nand U9052 (N_9052,N_2908,N_4094);
nand U9053 (N_9053,N_1449,N_1110);
nand U9054 (N_9054,N_2953,N_4816);
xnor U9055 (N_9055,N_806,N_335);
xor U9056 (N_9056,N_4805,N_4347);
nand U9057 (N_9057,N_4187,N_2814);
nor U9058 (N_9058,N_543,N_919);
or U9059 (N_9059,N_1176,N_1403);
and U9060 (N_9060,N_4196,N_4756);
and U9061 (N_9061,N_4364,N_208);
nor U9062 (N_9062,N_4925,N_661);
nand U9063 (N_9063,N_1323,N_3884);
xor U9064 (N_9064,N_4292,N_3357);
nand U9065 (N_9065,N_2700,N_3866);
or U9066 (N_9066,N_4733,N_3360);
or U9067 (N_9067,N_1044,N_2828);
nand U9068 (N_9068,N_4732,N_3085);
nand U9069 (N_9069,N_163,N_1530);
nand U9070 (N_9070,N_3004,N_3017);
nor U9071 (N_9071,N_3314,N_2664);
and U9072 (N_9072,N_3814,N_2448);
xnor U9073 (N_9073,N_2741,N_3762);
xnor U9074 (N_9074,N_2834,N_303);
nor U9075 (N_9075,N_3499,N_3954);
and U9076 (N_9076,N_3969,N_4088);
nand U9077 (N_9077,N_923,N_3842);
and U9078 (N_9078,N_4718,N_80);
nand U9079 (N_9079,N_1172,N_3067);
or U9080 (N_9080,N_1753,N_1973);
nor U9081 (N_9081,N_4863,N_4914);
and U9082 (N_9082,N_3791,N_2005);
nor U9083 (N_9083,N_4062,N_4181);
nand U9084 (N_9084,N_3113,N_1198);
and U9085 (N_9085,N_189,N_242);
or U9086 (N_9086,N_372,N_4679);
nor U9087 (N_9087,N_4232,N_4478);
and U9088 (N_9088,N_1602,N_4794);
nand U9089 (N_9089,N_4866,N_2803);
and U9090 (N_9090,N_4752,N_127);
nand U9091 (N_9091,N_3931,N_4974);
and U9092 (N_9092,N_341,N_1480);
and U9093 (N_9093,N_1250,N_2490);
nor U9094 (N_9094,N_3533,N_2554);
nor U9095 (N_9095,N_3115,N_1849);
nor U9096 (N_9096,N_1795,N_2966);
or U9097 (N_9097,N_2046,N_2841);
nand U9098 (N_9098,N_2557,N_4851);
nand U9099 (N_9099,N_2848,N_2842);
nor U9100 (N_9100,N_4523,N_1008);
nor U9101 (N_9101,N_1711,N_519);
and U9102 (N_9102,N_2177,N_2230);
xnor U9103 (N_9103,N_4633,N_1814);
nand U9104 (N_9104,N_2477,N_4047);
or U9105 (N_9105,N_674,N_1860);
xor U9106 (N_9106,N_4024,N_4669);
and U9107 (N_9107,N_2651,N_4485);
nand U9108 (N_9108,N_2192,N_1134);
xor U9109 (N_9109,N_3675,N_4056);
nand U9110 (N_9110,N_1484,N_4642);
nand U9111 (N_9111,N_2716,N_2921);
nor U9112 (N_9112,N_1949,N_83);
nor U9113 (N_9113,N_54,N_3920);
nand U9114 (N_9114,N_1400,N_795);
nor U9115 (N_9115,N_172,N_4200);
nor U9116 (N_9116,N_3684,N_4165);
or U9117 (N_9117,N_1495,N_2654);
nor U9118 (N_9118,N_982,N_4779);
and U9119 (N_9119,N_1711,N_654);
and U9120 (N_9120,N_2690,N_2462);
nor U9121 (N_9121,N_2281,N_546);
or U9122 (N_9122,N_2682,N_642);
or U9123 (N_9123,N_4212,N_1965);
xnor U9124 (N_9124,N_495,N_3952);
and U9125 (N_9125,N_4507,N_688);
or U9126 (N_9126,N_2606,N_338);
or U9127 (N_9127,N_1993,N_2066);
nand U9128 (N_9128,N_116,N_4001);
xor U9129 (N_9129,N_3897,N_2788);
or U9130 (N_9130,N_2627,N_1349);
nand U9131 (N_9131,N_3793,N_2933);
xor U9132 (N_9132,N_4436,N_4404);
or U9133 (N_9133,N_4364,N_3438);
nor U9134 (N_9134,N_1464,N_6);
nor U9135 (N_9135,N_3585,N_1678);
or U9136 (N_9136,N_915,N_3535);
or U9137 (N_9137,N_1546,N_4386);
and U9138 (N_9138,N_4074,N_412);
and U9139 (N_9139,N_3115,N_3197);
and U9140 (N_9140,N_2254,N_659);
nand U9141 (N_9141,N_1356,N_2238);
nor U9142 (N_9142,N_1915,N_4331);
nor U9143 (N_9143,N_4963,N_1603);
nand U9144 (N_9144,N_1899,N_240);
nand U9145 (N_9145,N_2936,N_4531);
nor U9146 (N_9146,N_1194,N_4625);
nand U9147 (N_9147,N_694,N_2568);
or U9148 (N_9148,N_1016,N_3187);
and U9149 (N_9149,N_495,N_3110);
or U9150 (N_9150,N_912,N_630);
nor U9151 (N_9151,N_482,N_3700);
nand U9152 (N_9152,N_2135,N_1279);
nand U9153 (N_9153,N_2905,N_3026);
or U9154 (N_9154,N_1083,N_1584);
nand U9155 (N_9155,N_4381,N_2877);
nand U9156 (N_9156,N_951,N_3358);
nand U9157 (N_9157,N_2107,N_1012);
and U9158 (N_9158,N_4744,N_410);
or U9159 (N_9159,N_4452,N_1520);
and U9160 (N_9160,N_940,N_2798);
nor U9161 (N_9161,N_3880,N_2123);
or U9162 (N_9162,N_3525,N_3700);
and U9163 (N_9163,N_500,N_2647);
nand U9164 (N_9164,N_3770,N_469);
nor U9165 (N_9165,N_248,N_2617);
or U9166 (N_9166,N_492,N_2208);
nand U9167 (N_9167,N_1695,N_1766);
or U9168 (N_9168,N_481,N_3406);
nor U9169 (N_9169,N_1141,N_1055);
nor U9170 (N_9170,N_3208,N_1727);
nor U9171 (N_9171,N_2859,N_1862);
xnor U9172 (N_9172,N_3594,N_3902);
nor U9173 (N_9173,N_4866,N_2095);
xor U9174 (N_9174,N_2955,N_922);
nor U9175 (N_9175,N_706,N_4758);
nor U9176 (N_9176,N_641,N_4866);
nand U9177 (N_9177,N_2016,N_2877);
and U9178 (N_9178,N_3358,N_1536);
nand U9179 (N_9179,N_3592,N_1832);
and U9180 (N_9180,N_4203,N_4611);
xor U9181 (N_9181,N_4921,N_2586);
nor U9182 (N_9182,N_3704,N_2610);
xnor U9183 (N_9183,N_3020,N_99);
and U9184 (N_9184,N_4033,N_3859);
nand U9185 (N_9185,N_1079,N_4015);
and U9186 (N_9186,N_3568,N_2775);
nor U9187 (N_9187,N_3256,N_356);
or U9188 (N_9188,N_2650,N_1251);
nand U9189 (N_9189,N_2052,N_3364);
nand U9190 (N_9190,N_2155,N_4081);
or U9191 (N_9191,N_434,N_4827);
nor U9192 (N_9192,N_1247,N_4689);
or U9193 (N_9193,N_2613,N_4801);
xnor U9194 (N_9194,N_2943,N_156);
xnor U9195 (N_9195,N_2038,N_278);
and U9196 (N_9196,N_3732,N_3037);
nand U9197 (N_9197,N_1885,N_4293);
or U9198 (N_9198,N_894,N_3712);
or U9199 (N_9199,N_2108,N_3809);
nor U9200 (N_9200,N_3701,N_3737);
xor U9201 (N_9201,N_2821,N_2690);
nand U9202 (N_9202,N_4128,N_3841);
xor U9203 (N_9203,N_2335,N_4292);
nand U9204 (N_9204,N_313,N_467);
nand U9205 (N_9205,N_1285,N_45);
nand U9206 (N_9206,N_1758,N_2782);
xor U9207 (N_9207,N_2273,N_3915);
or U9208 (N_9208,N_3516,N_4036);
or U9209 (N_9209,N_2128,N_823);
nand U9210 (N_9210,N_500,N_2480);
nand U9211 (N_9211,N_48,N_2141);
xor U9212 (N_9212,N_1329,N_1606);
nand U9213 (N_9213,N_470,N_369);
xor U9214 (N_9214,N_4251,N_2608);
nor U9215 (N_9215,N_3664,N_2106);
or U9216 (N_9216,N_4577,N_566);
and U9217 (N_9217,N_4442,N_3405);
and U9218 (N_9218,N_3191,N_4816);
nand U9219 (N_9219,N_2374,N_1398);
xnor U9220 (N_9220,N_851,N_4024);
nand U9221 (N_9221,N_3719,N_3860);
and U9222 (N_9222,N_2095,N_3349);
and U9223 (N_9223,N_249,N_1974);
nand U9224 (N_9224,N_730,N_2168);
or U9225 (N_9225,N_369,N_2463);
and U9226 (N_9226,N_770,N_2880);
nand U9227 (N_9227,N_4799,N_4157);
nand U9228 (N_9228,N_4088,N_3672);
nor U9229 (N_9229,N_3680,N_533);
and U9230 (N_9230,N_3239,N_4363);
nor U9231 (N_9231,N_2593,N_2367);
or U9232 (N_9232,N_4422,N_1756);
nor U9233 (N_9233,N_2552,N_3728);
xnor U9234 (N_9234,N_2631,N_2630);
nand U9235 (N_9235,N_3409,N_4958);
xor U9236 (N_9236,N_1703,N_1405);
nand U9237 (N_9237,N_1195,N_4706);
or U9238 (N_9238,N_1594,N_1950);
nor U9239 (N_9239,N_1936,N_2936);
or U9240 (N_9240,N_4551,N_1767);
and U9241 (N_9241,N_1034,N_1505);
and U9242 (N_9242,N_2187,N_13);
and U9243 (N_9243,N_1658,N_4032);
xnor U9244 (N_9244,N_2511,N_4276);
or U9245 (N_9245,N_3779,N_354);
and U9246 (N_9246,N_799,N_4065);
xor U9247 (N_9247,N_3677,N_953);
xnor U9248 (N_9248,N_4012,N_1817);
or U9249 (N_9249,N_1852,N_1781);
nand U9250 (N_9250,N_4821,N_2735);
nor U9251 (N_9251,N_3117,N_4227);
or U9252 (N_9252,N_3957,N_14);
nand U9253 (N_9253,N_3438,N_1054);
nand U9254 (N_9254,N_81,N_1822);
nand U9255 (N_9255,N_3280,N_1257);
nor U9256 (N_9256,N_3745,N_2743);
and U9257 (N_9257,N_160,N_588);
nor U9258 (N_9258,N_2736,N_3193);
nand U9259 (N_9259,N_3921,N_732);
nor U9260 (N_9260,N_3706,N_2598);
and U9261 (N_9261,N_2709,N_3105);
and U9262 (N_9262,N_2817,N_1753);
or U9263 (N_9263,N_4509,N_1799);
or U9264 (N_9264,N_655,N_779);
nor U9265 (N_9265,N_806,N_2412);
nand U9266 (N_9266,N_2892,N_2935);
and U9267 (N_9267,N_935,N_2547);
or U9268 (N_9268,N_3717,N_4341);
nor U9269 (N_9269,N_1078,N_922);
xnor U9270 (N_9270,N_2621,N_920);
xnor U9271 (N_9271,N_257,N_2622);
or U9272 (N_9272,N_3571,N_2301);
nor U9273 (N_9273,N_3582,N_2782);
and U9274 (N_9274,N_2974,N_2188);
and U9275 (N_9275,N_3207,N_336);
or U9276 (N_9276,N_4854,N_4332);
nor U9277 (N_9277,N_578,N_1476);
nor U9278 (N_9278,N_4609,N_3723);
nor U9279 (N_9279,N_235,N_89);
xnor U9280 (N_9280,N_4755,N_3407);
xnor U9281 (N_9281,N_293,N_2574);
nand U9282 (N_9282,N_3091,N_1218);
nand U9283 (N_9283,N_4482,N_1276);
nand U9284 (N_9284,N_3288,N_119);
nand U9285 (N_9285,N_3713,N_524);
nor U9286 (N_9286,N_2219,N_4472);
and U9287 (N_9287,N_1398,N_2266);
and U9288 (N_9288,N_798,N_1290);
or U9289 (N_9289,N_2265,N_4118);
and U9290 (N_9290,N_4381,N_1626);
nand U9291 (N_9291,N_3085,N_1639);
nor U9292 (N_9292,N_1481,N_247);
or U9293 (N_9293,N_1699,N_1657);
nand U9294 (N_9294,N_3414,N_1893);
nor U9295 (N_9295,N_4754,N_1668);
and U9296 (N_9296,N_403,N_1507);
nand U9297 (N_9297,N_910,N_1692);
xnor U9298 (N_9298,N_688,N_2099);
nand U9299 (N_9299,N_1827,N_3453);
xnor U9300 (N_9300,N_2007,N_1938);
nand U9301 (N_9301,N_2364,N_4533);
nand U9302 (N_9302,N_3290,N_4475);
nand U9303 (N_9303,N_2260,N_1194);
and U9304 (N_9304,N_2150,N_3704);
nand U9305 (N_9305,N_838,N_1741);
xor U9306 (N_9306,N_3712,N_3776);
nand U9307 (N_9307,N_4263,N_3873);
nand U9308 (N_9308,N_4060,N_4044);
nand U9309 (N_9309,N_670,N_3595);
xnor U9310 (N_9310,N_3173,N_1618);
xor U9311 (N_9311,N_4059,N_4090);
nand U9312 (N_9312,N_741,N_2892);
and U9313 (N_9313,N_449,N_1409);
nand U9314 (N_9314,N_482,N_298);
and U9315 (N_9315,N_894,N_2129);
or U9316 (N_9316,N_1811,N_1125);
and U9317 (N_9317,N_975,N_3569);
and U9318 (N_9318,N_100,N_1549);
or U9319 (N_9319,N_2274,N_2355);
xor U9320 (N_9320,N_3305,N_2158);
and U9321 (N_9321,N_500,N_4986);
and U9322 (N_9322,N_2759,N_1031);
or U9323 (N_9323,N_2969,N_999);
nand U9324 (N_9324,N_2483,N_2843);
nor U9325 (N_9325,N_2435,N_905);
and U9326 (N_9326,N_4721,N_227);
or U9327 (N_9327,N_3107,N_1719);
nor U9328 (N_9328,N_3605,N_2139);
nor U9329 (N_9329,N_789,N_259);
nand U9330 (N_9330,N_1659,N_2039);
or U9331 (N_9331,N_1120,N_252);
nor U9332 (N_9332,N_1415,N_3302);
xnor U9333 (N_9333,N_218,N_3502);
nand U9334 (N_9334,N_2741,N_3133);
and U9335 (N_9335,N_3569,N_1558);
xor U9336 (N_9336,N_209,N_106);
nand U9337 (N_9337,N_181,N_3834);
or U9338 (N_9338,N_1400,N_4259);
and U9339 (N_9339,N_2910,N_1863);
and U9340 (N_9340,N_3551,N_4003);
nand U9341 (N_9341,N_3274,N_3621);
nand U9342 (N_9342,N_2083,N_4216);
or U9343 (N_9343,N_3448,N_4492);
and U9344 (N_9344,N_226,N_3046);
nor U9345 (N_9345,N_1975,N_1123);
or U9346 (N_9346,N_2091,N_3992);
nor U9347 (N_9347,N_2181,N_68);
nor U9348 (N_9348,N_3149,N_2962);
and U9349 (N_9349,N_438,N_4137);
nand U9350 (N_9350,N_4111,N_3106);
nand U9351 (N_9351,N_2605,N_2877);
nor U9352 (N_9352,N_732,N_1783);
nand U9353 (N_9353,N_279,N_2219);
nor U9354 (N_9354,N_2284,N_3009);
nor U9355 (N_9355,N_3656,N_575);
nor U9356 (N_9356,N_611,N_3564);
and U9357 (N_9357,N_4386,N_2986);
nand U9358 (N_9358,N_1226,N_957);
or U9359 (N_9359,N_511,N_4730);
nand U9360 (N_9360,N_4521,N_987);
and U9361 (N_9361,N_859,N_2016);
nand U9362 (N_9362,N_4010,N_1155);
or U9363 (N_9363,N_991,N_3781);
nor U9364 (N_9364,N_3762,N_4586);
nor U9365 (N_9365,N_2615,N_1260);
nand U9366 (N_9366,N_1692,N_3473);
nor U9367 (N_9367,N_4777,N_3211);
nand U9368 (N_9368,N_2710,N_4510);
or U9369 (N_9369,N_3912,N_2288);
or U9370 (N_9370,N_3677,N_629);
nor U9371 (N_9371,N_594,N_2023);
or U9372 (N_9372,N_1589,N_3236);
nor U9373 (N_9373,N_153,N_27);
nand U9374 (N_9374,N_4656,N_2367);
nand U9375 (N_9375,N_4349,N_2993);
or U9376 (N_9376,N_4209,N_1272);
nor U9377 (N_9377,N_4,N_455);
or U9378 (N_9378,N_2831,N_851);
and U9379 (N_9379,N_1422,N_960);
nor U9380 (N_9380,N_2484,N_4295);
nor U9381 (N_9381,N_4457,N_2746);
or U9382 (N_9382,N_1150,N_2273);
and U9383 (N_9383,N_810,N_1302);
nand U9384 (N_9384,N_516,N_403);
nand U9385 (N_9385,N_1483,N_1229);
or U9386 (N_9386,N_1071,N_3824);
nand U9387 (N_9387,N_4114,N_3390);
nand U9388 (N_9388,N_4082,N_2946);
nand U9389 (N_9389,N_4184,N_4211);
nor U9390 (N_9390,N_1955,N_2848);
and U9391 (N_9391,N_4310,N_4487);
and U9392 (N_9392,N_2059,N_1551);
and U9393 (N_9393,N_4938,N_2976);
or U9394 (N_9394,N_94,N_3583);
nand U9395 (N_9395,N_3449,N_4769);
or U9396 (N_9396,N_4059,N_2049);
and U9397 (N_9397,N_918,N_1255);
or U9398 (N_9398,N_1558,N_1560);
nand U9399 (N_9399,N_3480,N_3772);
nor U9400 (N_9400,N_4005,N_802);
or U9401 (N_9401,N_4355,N_3911);
or U9402 (N_9402,N_454,N_606);
and U9403 (N_9403,N_2329,N_813);
nor U9404 (N_9404,N_1491,N_1225);
nor U9405 (N_9405,N_4222,N_3721);
nand U9406 (N_9406,N_4566,N_233);
nand U9407 (N_9407,N_2312,N_4146);
or U9408 (N_9408,N_899,N_4980);
or U9409 (N_9409,N_2391,N_4272);
and U9410 (N_9410,N_3073,N_3307);
nor U9411 (N_9411,N_1510,N_3569);
or U9412 (N_9412,N_2286,N_3189);
or U9413 (N_9413,N_4943,N_4011);
or U9414 (N_9414,N_1168,N_469);
nand U9415 (N_9415,N_2518,N_1829);
nor U9416 (N_9416,N_4350,N_1334);
or U9417 (N_9417,N_1101,N_2223);
nand U9418 (N_9418,N_4187,N_1592);
nor U9419 (N_9419,N_1052,N_90);
and U9420 (N_9420,N_1029,N_3206);
or U9421 (N_9421,N_1317,N_906);
or U9422 (N_9422,N_3554,N_60);
nor U9423 (N_9423,N_1927,N_2671);
and U9424 (N_9424,N_2180,N_2862);
nor U9425 (N_9425,N_3710,N_426);
nand U9426 (N_9426,N_4214,N_3351);
and U9427 (N_9427,N_4338,N_1579);
nor U9428 (N_9428,N_918,N_4846);
and U9429 (N_9429,N_2306,N_2539);
nor U9430 (N_9430,N_3152,N_2916);
nand U9431 (N_9431,N_2487,N_2048);
xnor U9432 (N_9432,N_1280,N_4167);
nor U9433 (N_9433,N_3673,N_1914);
or U9434 (N_9434,N_2820,N_1172);
and U9435 (N_9435,N_4455,N_3581);
nor U9436 (N_9436,N_4804,N_1580);
xnor U9437 (N_9437,N_4714,N_1996);
and U9438 (N_9438,N_3430,N_3385);
nor U9439 (N_9439,N_4768,N_4219);
nor U9440 (N_9440,N_4733,N_1943);
nor U9441 (N_9441,N_2291,N_1451);
nor U9442 (N_9442,N_4788,N_4164);
nor U9443 (N_9443,N_1152,N_3819);
nand U9444 (N_9444,N_610,N_3247);
and U9445 (N_9445,N_4698,N_179);
nor U9446 (N_9446,N_4645,N_2864);
nand U9447 (N_9447,N_4098,N_1442);
and U9448 (N_9448,N_3700,N_73);
nand U9449 (N_9449,N_2195,N_4114);
nor U9450 (N_9450,N_1296,N_2054);
and U9451 (N_9451,N_2724,N_4739);
or U9452 (N_9452,N_2993,N_4535);
or U9453 (N_9453,N_2893,N_4114);
xor U9454 (N_9454,N_387,N_2853);
nand U9455 (N_9455,N_1422,N_1914);
and U9456 (N_9456,N_4505,N_3475);
nand U9457 (N_9457,N_4621,N_1005);
nand U9458 (N_9458,N_4831,N_2629);
or U9459 (N_9459,N_545,N_2470);
nor U9460 (N_9460,N_4140,N_1176);
and U9461 (N_9461,N_632,N_3268);
or U9462 (N_9462,N_1836,N_4219);
nand U9463 (N_9463,N_854,N_3539);
nand U9464 (N_9464,N_3487,N_2573);
and U9465 (N_9465,N_1189,N_2821);
and U9466 (N_9466,N_4933,N_287);
nor U9467 (N_9467,N_2866,N_3329);
nand U9468 (N_9468,N_2183,N_1928);
nor U9469 (N_9469,N_2784,N_2089);
nand U9470 (N_9470,N_152,N_395);
or U9471 (N_9471,N_1400,N_859);
nor U9472 (N_9472,N_464,N_771);
or U9473 (N_9473,N_509,N_1837);
and U9474 (N_9474,N_3293,N_562);
nor U9475 (N_9475,N_1706,N_4667);
and U9476 (N_9476,N_1634,N_1803);
nor U9477 (N_9477,N_4100,N_282);
nand U9478 (N_9478,N_2669,N_4012);
and U9479 (N_9479,N_3782,N_1878);
nor U9480 (N_9480,N_749,N_4366);
and U9481 (N_9481,N_27,N_1844);
nand U9482 (N_9482,N_1678,N_3847);
and U9483 (N_9483,N_711,N_110);
or U9484 (N_9484,N_1419,N_3827);
xnor U9485 (N_9485,N_1205,N_1089);
nand U9486 (N_9486,N_1578,N_2537);
nor U9487 (N_9487,N_2967,N_2957);
nor U9488 (N_9488,N_2887,N_3086);
and U9489 (N_9489,N_614,N_4968);
nand U9490 (N_9490,N_1072,N_2135);
or U9491 (N_9491,N_1852,N_997);
and U9492 (N_9492,N_421,N_4002);
nor U9493 (N_9493,N_4300,N_2463);
nand U9494 (N_9494,N_360,N_1741);
nand U9495 (N_9495,N_2451,N_2931);
nand U9496 (N_9496,N_2299,N_2129);
or U9497 (N_9497,N_586,N_1551);
nand U9498 (N_9498,N_2021,N_1492);
nand U9499 (N_9499,N_3603,N_4515);
nor U9500 (N_9500,N_3794,N_4120);
nand U9501 (N_9501,N_4180,N_2501);
or U9502 (N_9502,N_1161,N_251);
or U9503 (N_9503,N_4855,N_1929);
and U9504 (N_9504,N_1064,N_4620);
nand U9505 (N_9505,N_1403,N_2731);
and U9506 (N_9506,N_4594,N_1172);
or U9507 (N_9507,N_2112,N_4155);
nand U9508 (N_9508,N_3463,N_3769);
nand U9509 (N_9509,N_1501,N_3123);
and U9510 (N_9510,N_726,N_3690);
and U9511 (N_9511,N_4256,N_4426);
or U9512 (N_9512,N_2337,N_1682);
nor U9513 (N_9513,N_88,N_114);
nor U9514 (N_9514,N_2496,N_4813);
nor U9515 (N_9515,N_2967,N_2816);
nor U9516 (N_9516,N_2247,N_4588);
and U9517 (N_9517,N_1966,N_4968);
and U9518 (N_9518,N_4168,N_1010);
or U9519 (N_9519,N_2333,N_3019);
nand U9520 (N_9520,N_144,N_2328);
or U9521 (N_9521,N_3704,N_318);
and U9522 (N_9522,N_2873,N_2539);
and U9523 (N_9523,N_2829,N_2667);
or U9524 (N_9524,N_1992,N_1667);
nand U9525 (N_9525,N_2973,N_1400);
and U9526 (N_9526,N_1778,N_2456);
xor U9527 (N_9527,N_4709,N_68);
nand U9528 (N_9528,N_2741,N_2483);
or U9529 (N_9529,N_2546,N_2655);
and U9530 (N_9530,N_876,N_4862);
nand U9531 (N_9531,N_111,N_1365);
or U9532 (N_9532,N_543,N_2764);
nand U9533 (N_9533,N_3445,N_2294);
nor U9534 (N_9534,N_2784,N_2328);
or U9535 (N_9535,N_1937,N_746);
and U9536 (N_9536,N_4242,N_446);
nor U9537 (N_9537,N_1153,N_3259);
or U9538 (N_9538,N_4397,N_1952);
and U9539 (N_9539,N_3263,N_1527);
and U9540 (N_9540,N_1802,N_1609);
and U9541 (N_9541,N_2916,N_1959);
nand U9542 (N_9542,N_3628,N_4789);
or U9543 (N_9543,N_2224,N_908);
and U9544 (N_9544,N_1457,N_2873);
nor U9545 (N_9545,N_2203,N_4659);
and U9546 (N_9546,N_1425,N_4796);
and U9547 (N_9547,N_2115,N_1619);
xnor U9548 (N_9548,N_4631,N_953);
or U9549 (N_9549,N_2983,N_1664);
or U9550 (N_9550,N_4279,N_4923);
or U9551 (N_9551,N_3672,N_4906);
xor U9552 (N_9552,N_2888,N_1324);
and U9553 (N_9553,N_1703,N_718);
and U9554 (N_9554,N_2348,N_1218);
nand U9555 (N_9555,N_2195,N_2090);
or U9556 (N_9556,N_4956,N_2097);
nor U9557 (N_9557,N_2649,N_2996);
and U9558 (N_9558,N_2927,N_337);
nor U9559 (N_9559,N_1524,N_3319);
and U9560 (N_9560,N_1580,N_3088);
nand U9561 (N_9561,N_4288,N_811);
nand U9562 (N_9562,N_3637,N_1653);
xnor U9563 (N_9563,N_4557,N_2044);
or U9564 (N_9564,N_1285,N_4796);
nand U9565 (N_9565,N_1993,N_2589);
or U9566 (N_9566,N_275,N_542);
nor U9567 (N_9567,N_2475,N_354);
nor U9568 (N_9568,N_610,N_4086);
or U9569 (N_9569,N_1987,N_1231);
nor U9570 (N_9570,N_769,N_1470);
nor U9571 (N_9571,N_2062,N_885);
or U9572 (N_9572,N_4036,N_2267);
nor U9573 (N_9573,N_2262,N_2985);
and U9574 (N_9574,N_1706,N_1511);
nand U9575 (N_9575,N_2547,N_2392);
xnor U9576 (N_9576,N_1124,N_1034);
nor U9577 (N_9577,N_4202,N_1428);
and U9578 (N_9578,N_3422,N_1360);
or U9579 (N_9579,N_35,N_3778);
nor U9580 (N_9580,N_2190,N_876);
nand U9581 (N_9581,N_3391,N_2284);
or U9582 (N_9582,N_2021,N_4864);
nand U9583 (N_9583,N_4295,N_2400);
or U9584 (N_9584,N_629,N_2431);
nand U9585 (N_9585,N_2644,N_2339);
and U9586 (N_9586,N_2695,N_4788);
and U9587 (N_9587,N_1377,N_4623);
nand U9588 (N_9588,N_2720,N_3525);
nor U9589 (N_9589,N_1574,N_241);
nand U9590 (N_9590,N_1853,N_2243);
nand U9591 (N_9591,N_2142,N_4736);
and U9592 (N_9592,N_1037,N_1151);
nor U9593 (N_9593,N_3585,N_411);
and U9594 (N_9594,N_1814,N_3779);
nand U9595 (N_9595,N_2243,N_2052);
or U9596 (N_9596,N_1943,N_4462);
and U9597 (N_9597,N_1682,N_4692);
nand U9598 (N_9598,N_4664,N_3075);
nor U9599 (N_9599,N_1937,N_2080);
and U9600 (N_9600,N_3201,N_1326);
and U9601 (N_9601,N_512,N_3715);
nor U9602 (N_9602,N_4081,N_4402);
nor U9603 (N_9603,N_4217,N_4650);
xor U9604 (N_9604,N_2379,N_4914);
and U9605 (N_9605,N_370,N_2864);
xor U9606 (N_9606,N_2421,N_363);
and U9607 (N_9607,N_1511,N_1204);
and U9608 (N_9608,N_3723,N_2216);
or U9609 (N_9609,N_1043,N_2727);
or U9610 (N_9610,N_2237,N_2616);
or U9611 (N_9611,N_1311,N_131);
nor U9612 (N_9612,N_3934,N_4258);
nor U9613 (N_9613,N_3198,N_4438);
and U9614 (N_9614,N_2484,N_4601);
nand U9615 (N_9615,N_4558,N_990);
nand U9616 (N_9616,N_4192,N_4280);
nor U9617 (N_9617,N_2500,N_6);
nor U9618 (N_9618,N_4471,N_3844);
nand U9619 (N_9619,N_2975,N_995);
nand U9620 (N_9620,N_62,N_885);
and U9621 (N_9621,N_3599,N_2763);
and U9622 (N_9622,N_910,N_3478);
nor U9623 (N_9623,N_1199,N_2199);
and U9624 (N_9624,N_2576,N_3758);
xor U9625 (N_9625,N_1592,N_3014);
and U9626 (N_9626,N_2461,N_4036);
nand U9627 (N_9627,N_1646,N_1043);
nor U9628 (N_9628,N_2315,N_565);
nand U9629 (N_9629,N_2212,N_349);
nand U9630 (N_9630,N_4111,N_988);
nand U9631 (N_9631,N_2504,N_3347);
xnor U9632 (N_9632,N_214,N_4639);
nor U9633 (N_9633,N_4120,N_2515);
and U9634 (N_9634,N_2069,N_2107);
nand U9635 (N_9635,N_3625,N_487);
and U9636 (N_9636,N_3663,N_2789);
nand U9637 (N_9637,N_2245,N_4498);
and U9638 (N_9638,N_2923,N_2396);
or U9639 (N_9639,N_4627,N_2595);
nor U9640 (N_9640,N_1570,N_1452);
nand U9641 (N_9641,N_1371,N_739);
nor U9642 (N_9642,N_611,N_1957);
nand U9643 (N_9643,N_4174,N_3511);
or U9644 (N_9644,N_2548,N_1111);
nand U9645 (N_9645,N_4168,N_3920);
xor U9646 (N_9646,N_4929,N_3997);
or U9647 (N_9647,N_134,N_3670);
or U9648 (N_9648,N_953,N_1190);
nand U9649 (N_9649,N_1529,N_1102);
or U9650 (N_9650,N_621,N_2268);
nor U9651 (N_9651,N_2705,N_3793);
nor U9652 (N_9652,N_2355,N_4657);
xor U9653 (N_9653,N_1083,N_937);
nor U9654 (N_9654,N_4532,N_2566);
xnor U9655 (N_9655,N_2628,N_3529);
nand U9656 (N_9656,N_2417,N_2819);
or U9657 (N_9657,N_152,N_1197);
or U9658 (N_9658,N_98,N_496);
nand U9659 (N_9659,N_1083,N_2936);
and U9660 (N_9660,N_2543,N_4248);
or U9661 (N_9661,N_3995,N_1246);
nor U9662 (N_9662,N_2288,N_4080);
and U9663 (N_9663,N_3694,N_2382);
xnor U9664 (N_9664,N_3188,N_1773);
or U9665 (N_9665,N_2739,N_3138);
and U9666 (N_9666,N_55,N_773);
and U9667 (N_9667,N_4553,N_3392);
and U9668 (N_9668,N_504,N_3328);
and U9669 (N_9669,N_3011,N_3402);
nand U9670 (N_9670,N_2425,N_871);
xor U9671 (N_9671,N_1277,N_4656);
or U9672 (N_9672,N_3291,N_1518);
or U9673 (N_9673,N_3331,N_882);
nor U9674 (N_9674,N_2620,N_481);
xnor U9675 (N_9675,N_1034,N_3277);
xor U9676 (N_9676,N_1662,N_398);
and U9677 (N_9677,N_145,N_1598);
and U9678 (N_9678,N_2239,N_226);
nor U9679 (N_9679,N_1818,N_843);
and U9680 (N_9680,N_2111,N_3899);
or U9681 (N_9681,N_862,N_2350);
nand U9682 (N_9682,N_4302,N_4975);
nand U9683 (N_9683,N_1713,N_1878);
nand U9684 (N_9684,N_1716,N_604);
nor U9685 (N_9685,N_4514,N_710);
and U9686 (N_9686,N_1994,N_4327);
and U9687 (N_9687,N_3720,N_2480);
or U9688 (N_9688,N_1090,N_2092);
nand U9689 (N_9689,N_3688,N_2188);
or U9690 (N_9690,N_2994,N_2873);
nor U9691 (N_9691,N_4473,N_291);
and U9692 (N_9692,N_4722,N_3095);
nor U9693 (N_9693,N_4621,N_3271);
xnor U9694 (N_9694,N_4832,N_1079);
nand U9695 (N_9695,N_818,N_2428);
and U9696 (N_9696,N_3284,N_1634);
nor U9697 (N_9697,N_2520,N_4094);
nand U9698 (N_9698,N_898,N_2329);
nand U9699 (N_9699,N_3510,N_4711);
nor U9700 (N_9700,N_2996,N_1739);
nand U9701 (N_9701,N_1709,N_2138);
and U9702 (N_9702,N_3130,N_731);
or U9703 (N_9703,N_4208,N_3099);
or U9704 (N_9704,N_3578,N_1478);
xor U9705 (N_9705,N_4443,N_1374);
or U9706 (N_9706,N_264,N_1179);
and U9707 (N_9707,N_4073,N_3217);
or U9708 (N_9708,N_438,N_784);
nand U9709 (N_9709,N_3477,N_4037);
or U9710 (N_9710,N_2624,N_1189);
xnor U9711 (N_9711,N_273,N_2806);
or U9712 (N_9712,N_1848,N_215);
and U9713 (N_9713,N_4515,N_1219);
and U9714 (N_9714,N_3119,N_930);
and U9715 (N_9715,N_2968,N_1346);
and U9716 (N_9716,N_2488,N_1245);
and U9717 (N_9717,N_250,N_2848);
or U9718 (N_9718,N_4247,N_20);
nor U9719 (N_9719,N_4230,N_1274);
or U9720 (N_9720,N_4107,N_1217);
and U9721 (N_9721,N_2938,N_4376);
and U9722 (N_9722,N_2012,N_869);
nor U9723 (N_9723,N_655,N_3965);
and U9724 (N_9724,N_3656,N_224);
and U9725 (N_9725,N_2134,N_188);
nor U9726 (N_9726,N_4437,N_317);
or U9727 (N_9727,N_530,N_2942);
nor U9728 (N_9728,N_2607,N_1435);
nand U9729 (N_9729,N_4080,N_3021);
or U9730 (N_9730,N_3428,N_2675);
nand U9731 (N_9731,N_2989,N_1171);
nor U9732 (N_9732,N_1219,N_2394);
nand U9733 (N_9733,N_2852,N_3668);
nand U9734 (N_9734,N_1694,N_309);
xor U9735 (N_9735,N_1121,N_4473);
nand U9736 (N_9736,N_2043,N_737);
nand U9737 (N_9737,N_2161,N_256);
and U9738 (N_9738,N_4578,N_3453);
nand U9739 (N_9739,N_4022,N_4441);
nor U9740 (N_9740,N_1582,N_926);
nor U9741 (N_9741,N_2961,N_1152);
and U9742 (N_9742,N_3429,N_3878);
nor U9743 (N_9743,N_3791,N_4267);
and U9744 (N_9744,N_2718,N_2377);
and U9745 (N_9745,N_932,N_1011);
or U9746 (N_9746,N_915,N_1080);
xnor U9747 (N_9747,N_178,N_1688);
xnor U9748 (N_9748,N_1627,N_19);
and U9749 (N_9749,N_3660,N_778);
and U9750 (N_9750,N_4127,N_1249);
or U9751 (N_9751,N_300,N_3306);
or U9752 (N_9752,N_4368,N_2880);
xnor U9753 (N_9753,N_312,N_1460);
nor U9754 (N_9754,N_2736,N_1380);
or U9755 (N_9755,N_2742,N_3255);
xor U9756 (N_9756,N_3365,N_3080);
xor U9757 (N_9757,N_4134,N_2453);
and U9758 (N_9758,N_3823,N_3817);
nand U9759 (N_9759,N_3769,N_1185);
or U9760 (N_9760,N_751,N_5);
nor U9761 (N_9761,N_2570,N_742);
and U9762 (N_9762,N_4174,N_2032);
or U9763 (N_9763,N_4990,N_543);
nor U9764 (N_9764,N_4520,N_1301);
nand U9765 (N_9765,N_648,N_3352);
or U9766 (N_9766,N_797,N_928);
nand U9767 (N_9767,N_344,N_188);
and U9768 (N_9768,N_2742,N_2312);
nor U9769 (N_9769,N_1446,N_1980);
and U9770 (N_9770,N_2121,N_4209);
xnor U9771 (N_9771,N_1359,N_94);
or U9772 (N_9772,N_1198,N_1110);
nand U9773 (N_9773,N_3269,N_23);
nor U9774 (N_9774,N_4629,N_4210);
nand U9775 (N_9775,N_3644,N_498);
nand U9776 (N_9776,N_4832,N_2756);
nand U9777 (N_9777,N_1222,N_3277);
and U9778 (N_9778,N_2914,N_1135);
or U9779 (N_9779,N_1471,N_4857);
nand U9780 (N_9780,N_4940,N_2484);
and U9781 (N_9781,N_2292,N_691);
xor U9782 (N_9782,N_719,N_1196);
or U9783 (N_9783,N_3977,N_4365);
nor U9784 (N_9784,N_4838,N_1839);
nor U9785 (N_9785,N_4966,N_4893);
nor U9786 (N_9786,N_681,N_3893);
and U9787 (N_9787,N_4305,N_196);
nand U9788 (N_9788,N_3771,N_4801);
or U9789 (N_9789,N_4674,N_2323);
nor U9790 (N_9790,N_1415,N_3931);
and U9791 (N_9791,N_3632,N_1000);
nand U9792 (N_9792,N_2654,N_3875);
nor U9793 (N_9793,N_4664,N_2357);
nand U9794 (N_9794,N_2239,N_4928);
nand U9795 (N_9795,N_3237,N_3918);
nor U9796 (N_9796,N_3993,N_3562);
and U9797 (N_9797,N_1715,N_517);
nand U9798 (N_9798,N_3700,N_4162);
and U9799 (N_9799,N_49,N_4411);
xor U9800 (N_9800,N_468,N_3929);
and U9801 (N_9801,N_4534,N_3747);
or U9802 (N_9802,N_3813,N_2475);
nand U9803 (N_9803,N_3470,N_1931);
xnor U9804 (N_9804,N_3690,N_3346);
and U9805 (N_9805,N_3075,N_3693);
nor U9806 (N_9806,N_25,N_3486);
or U9807 (N_9807,N_1489,N_1259);
nand U9808 (N_9808,N_4074,N_3919);
or U9809 (N_9809,N_4126,N_4909);
nand U9810 (N_9810,N_1030,N_2638);
nor U9811 (N_9811,N_3654,N_1552);
nor U9812 (N_9812,N_3228,N_4314);
xor U9813 (N_9813,N_3281,N_2489);
nor U9814 (N_9814,N_1038,N_4576);
nand U9815 (N_9815,N_365,N_1608);
nand U9816 (N_9816,N_431,N_388);
xnor U9817 (N_9817,N_3290,N_2319);
and U9818 (N_9818,N_969,N_4636);
nor U9819 (N_9819,N_1470,N_1381);
or U9820 (N_9820,N_3646,N_3406);
nand U9821 (N_9821,N_3522,N_4476);
nand U9822 (N_9822,N_4751,N_1053);
nand U9823 (N_9823,N_3064,N_1110);
and U9824 (N_9824,N_40,N_3875);
xor U9825 (N_9825,N_2893,N_1410);
nor U9826 (N_9826,N_2817,N_4853);
nand U9827 (N_9827,N_2546,N_290);
or U9828 (N_9828,N_4734,N_955);
nor U9829 (N_9829,N_263,N_1473);
nor U9830 (N_9830,N_1675,N_4554);
or U9831 (N_9831,N_4753,N_2726);
or U9832 (N_9832,N_2436,N_3003);
or U9833 (N_9833,N_2206,N_1067);
nor U9834 (N_9834,N_2370,N_2724);
and U9835 (N_9835,N_2311,N_2061);
nor U9836 (N_9836,N_1002,N_3368);
or U9837 (N_9837,N_97,N_3789);
or U9838 (N_9838,N_1517,N_2216);
or U9839 (N_9839,N_712,N_3101);
nor U9840 (N_9840,N_4233,N_4830);
nor U9841 (N_9841,N_4111,N_2968);
or U9842 (N_9842,N_4240,N_499);
and U9843 (N_9843,N_2290,N_3491);
and U9844 (N_9844,N_4491,N_2721);
xnor U9845 (N_9845,N_3814,N_3412);
nand U9846 (N_9846,N_4580,N_4033);
or U9847 (N_9847,N_1713,N_1511);
nor U9848 (N_9848,N_3710,N_658);
or U9849 (N_9849,N_966,N_4417);
nand U9850 (N_9850,N_1103,N_3290);
and U9851 (N_9851,N_3860,N_4305);
or U9852 (N_9852,N_2784,N_3894);
nor U9853 (N_9853,N_1093,N_4116);
nand U9854 (N_9854,N_233,N_3106);
and U9855 (N_9855,N_3119,N_4628);
nand U9856 (N_9856,N_4160,N_805);
and U9857 (N_9857,N_1233,N_3993);
or U9858 (N_9858,N_1804,N_951);
nor U9859 (N_9859,N_3431,N_1106);
nor U9860 (N_9860,N_806,N_4909);
and U9861 (N_9861,N_1586,N_813);
and U9862 (N_9862,N_1710,N_4729);
nor U9863 (N_9863,N_209,N_4482);
or U9864 (N_9864,N_192,N_1657);
xor U9865 (N_9865,N_667,N_4334);
and U9866 (N_9866,N_1183,N_2991);
nor U9867 (N_9867,N_2959,N_253);
nand U9868 (N_9868,N_1159,N_810);
nand U9869 (N_9869,N_4065,N_723);
xnor U9870 (N_9870,N_378,N_3595);
or U9871 (N_9871,N_353,N_837);
or U9872 (N_9872,N_4950,N_2149);
or U9873 (N_9873,N_2812,N_965);
nor U9874 (N_9874,N_3252,N_2716);
or U9875 (N_9875,N_1289,N_244);
nand U9876 (N_9876,N_1862,N_1795);
nand U9877 (N_9877,N_893,N_539);
nor U9878 (N_9878,N_1725,N_3248);
and U9879 (N_9879,N_1603,N_3409);
or U9880 (N_9880,N_4336,N_4871);
nand U9881 (N_9881,N_3884,N_2354);
nor U9882 (N_9882,N_234,N_2304);
xor U9883 (N_9883,N_2543,N_1310);
or U9884 (N_9884,N_3753,N_3547);
or U9885 (N_9885,N_4709,N_4982);
and U9886 (N_9886,N_4596,N_1799);
xnor U9887 (N_9887,N_3828,N_85);
or U9888 (N_9888,N_2244,N_2760);
and U9889 (N_9889,N_1628,N_4898);
or U9890 (N_9890,N_5,N_2138);
nor U9891 (N_9891,N_2018,N_1399);
nor U9892 (N_9892,N_2396,N_2557);
or U9893 (N_9893,N_656,N_2515);
nor U9894 (N_9894,N_880,N_916);
xnor U9895 (N_9895,N_2351,N_415);
nand U9896 (N_9896,N_3765,N_3146);
nor U9897 (N_9897,N_3139,N_2533);
nand U9898 (N_9898,N_3362,N_2456);
and U9899 (N_9899,N_42,N_1978);
nor U9900 (N_9900,N_3722,N_1245);
and U9901 (N_9901,N_2215,N_111);
nand U9902 (N_9902,N_7,N_191);
nand U9903 (N_9903,N_88,N_2430);
and U9904 (N_9904,N_1258,N_958);
nor U9905 (N_9905,N_1513,N_4982);
or U9906 (N_9906,N_1350,N_1876);
and U9907 (N_9907,N_3546,N_2896);
or U9908 (N_9908,N_2823,N_3218);
and U9909 (N_9909,N_4892,N_2267);
nand U9910 (N_9910,N_1893,N_4852);
nand U9911 (N_9911,N_4905,N_1935);
nor U9912 (N_9912,N_1348,N_1613);
xor U9913 (N_9913,N_2318,N_2178);
or U9914 (N_9914,N_2330,N_4297);
nand U9915 (N_9915,N_4297,N_2780);
nor U9916 (N_9916,N_4983,N_358);
and U9917 (N_9917,N_470,N_1841);
or U9918 (N_9918,N_2876,N_2327);
and U9919 (N_9919,N_874,N_1855);
and U9920 (N_9920,N_300,N_3201);
nand U9921 (N_9921,N_3874,N_247);
xor U9922 (N_9922,N_4888,N_4530);
and U9923 (N_9923,N_4054,N_1936);
xnor U9924 (N_9924,N_1201,N_1667);
and U9925 (N_9925,N_1521,N_4985);
and U9926 (N_9926,N_3974,N_1441);
or U9927 (N_9927,N_2240,N_3545);
nor U9928 (N_9928,N_3404,N_2756);
nor U9929 (N_9929,N_3825,N_3744);
xor U9930 (N_9930,N_2685,N_4649);
or U9931 (N_9931,N_1932,N_2949);
nor U9932 (N_9932,N_2680,N_366);
nand U9933 (N_9933,N_4654,N_113);
nor U9934 (N_9934,N_1680,N_2244);
and U9935 (N_9935,N_3218,N_1260);
or U9936 (N_9936,N_851,N_4053);
nor U9937 (N_9937,N_649,N_4480);
nand U9938 (N_9938,N_3344,N_1948);
xor U9939 (N_9939,N_90,N_4071);
and U9940 (N_9940,N_4033,N_3083);
nand U9941 (N_9941,N_3733,N_9);
nand U9942 (N_9942,N_3190,N_4860);
nor U9943 (N_9943,N_531,N_3026);
and U9944 (N_9944,N_3807,N_1843);
nand U9945 (N_9945,N_2591,N_4574);
nor U9946 (N_9946,N_1024,N_2825);
or U9947 (N_9947,N_2137,N_3059);
nand U9948 (N_9948,N_1140,N_3218);
nand U9949 (N_9949,N_1296,N_4423);
xor U9950 (N_9950,N_977,N_812);
and U9951 (N_9951,N_399,N_1592);
or U9952 (N_9952,N_2503,N_1099);
nor U9953 (N_9953,N_4826,N_1291);
xnor U9954 (N_9954,N_4640,N_2901);
or U9955 (N_9955,N_2431,N_747);
and U9956 (N_9956,N_264,N_220);
or U9957 (N_9957,N_4048,N_536);
or U9958 (N_9958,N_4044,N_3477);
and U9959 (N_9959,N_4498,N_777);
or U9960 (N_9960,N_4293,N_3905);
nand U9961 (N_9961,N_4676,N_2362);
or U9962 (N_9962,N_2095,N_3755);
nor U9963 (N_9963,N_2977,N_2293);
and U9964 (N_9964,N_2817,N_557);
and U9965 (N_9965,N_383,N_2104);
nor U9966 (N_9966,N_2295,N_13);
nand U9967 (N_9967,N_716,N_101);
and U9968 (N_9968,N_4223,N_2736);
or U9969 (N_9969,N_4399,N_1317);
xor U9970 (N_9970,N_420,N_2807);
nor U9971 (N_9971,N_4662,N_4917);
or U9972 (N_9972,N_166,N_3794);
nor U9973 (N_9973,N_2083,N_1382);
or U9974 (N_9974,N_111,N_774);
and U9975 (N_9975,N_4836,N_938);
nor U9976 (N_9976,N_1532,N_761);
nor U9977 (N_9977,N_342,N_4007);
nor U9978 (N_9978,N_3053,N_1097);
nand U9979 (N_9979,N_2247,N_3768);
and U9980 (N_9980,N_1037,N_4748);
and U9981 (N_9981,N_4536,N_2005);
nand U9982 (N_9982,N_4002,N_411);
nand U9983 (N_9983,N_786,N_4262);
or U9984 (N_9984,N_1176,N_3307);
nand U9985 (N_9985,N_4209,N_1924);
or U9986 (N_9986,N_2411,N_2846);
or U9987 (N_9987,N_2848,N_1163);
or U9988 (N_9988,N_17,N_3092);
nand U9989 (N_9989,N_4215,N_665);
and U9990 (N_9990,N_1711,N_2597);
and U9991 (N_9991,N_2387,N_148);
nor U9992 (N_9992,N_117,N_4721);
and U9993 (N_9993,N_2521,N_2105);
xor U9994 (N_9994,N_4809,N_3429);
and U9995 (N_9995,N_278,N_2639);
and U9996 (N_9996,N_486,N_3838);
nor U9997 (N_9997,N_4692,N_631);
or U9998 (N_9998,N_4839,N_2637);
nor U9999 (N_9999,N_2735,N_4900);
or U10000 (N_10000,N_6114,N_8889);
or U10001 (N_10001,N_6367,N_8414);
nand U10002 (N_10002,N_9642,N_9942);
and U10003 (N_10003,N_5642,N_9992);
or U10004 (N_10004,N_6081,N_5422);
xor U10005 (N_10005,N_9384,N_7512);
nor U10006 (N_10006,N_9711,N_7455);
nand U10007 (N_10007,N_5322,N_6262);
nand U10008 (N_10008,N_5460,N_7283);
or U10009 (N_10009,N_7821,N_6406);
and U10010 (N_10010,N_9926,N_5574);
nor U10011 (N_10011,N_9034,N_6239);
nor U10012 (N_10012,N_6767,N_5597);
or U10013 (N_10013,N_7612,N_7861);
and U10014 (N_10014,N_9988,N_9090);
nor U10015 (N_10015,N_8278,N_5491);
and U10016 (N_10016,N_9420,N_6445);
and U10017 (N_10017,N_8736,N_8345);
nand U10018 (N_10018,N_8806,N_5655);
and U10019 (N_10019,N_8125,N_8769);
xnor U10020 (N_10020,N_9506,N_5571);
and U10021 (N_10021,N_5798,N_8646);
and U10022 (N_10022,N_6893,N_8279);
and U10023 (N_10023,N_6671,N_5237);
nor U10024 (N_10024,N_8775,N_6645);
or U10025 (N_10025,N_9855,N_7272);
nor U10026 (N_10026,N_6333,N_8255);
or U10027 (N_10027,N_5507,N_7242);
nand U10028 (N_10028,N_7531,N_7252);
nand U10029 (N_10029,N_8175,N_8836);
or U10030 (N_10030,N_9691,N_5921);
or U10031 (N_10031,N_7948,N_8997);
nor U10032 (N_10032,N_8390,N_6039);
xnor U10033 (N_10033,N_9836,N_5898);
nand U10034 (N_10034,N_6998,N_9229);
or U10035 (N_10035,N_7057,N_5693);
xor U10036 (N_10036,N_9455,N_8027);
or U10037 (N_10037,N_7785,N_9225);
and U10038 (N_10038,N_8469,N_8969);
and U10039 (N_10039,N_5011,N_9805);
or U10040 (N_10040,N_9631,N_6506);
nor U10041 (N_10041,N_8398,N_6533);
or U10042 (N_10042,N_9155,N_5689);
xnor U10043 (N_10043,N_8701,N_6644);
and U10044 (N_10044,N_6425,N_8638);
nor U10045 (N_10045,N_6672,N_9152);
nand U10046 (N_10046,N_5244,N_7894);
and U10047 (N_10047,N_6088,N_8204);
nand U10048 (N_10048,N_5379,N_6718);
nand U10049 (N_10049,N_8802,N_7820);
nand U10050 (N_10050,N_6844,N_6670);
and U10051 (N_10051,N_7402,N_5695);
nand U10052 (N_10052,N_6054,N_7227);
or U10053 (N_10053,N_6261,N_6525);
nor U10054 (N_10054,N_6236,N_9796);
nor U10055 (N_10055,N_8239,N_9877);
nand U10056 (N_10056,N_9434,N_6488);
nand U10057 (N_10057,N_8168,N_8086);
and U10058 (N_10058,N_9228,N_6611);
and U10059 (N_10059,N_7139,N_7117);
xor U10060 (N_10060,N_5313,N_8309);
and U10061 (N_10061,N_8515,N_7831);
nor U10062 (N_10062,N_9703,N_5954);
nor U10063 (N_10063,N_9361,N_9615);
and U10064 (N_10064,N_8322,N_8604);
and U10065 (N_10065,N_8008,N_9098);
and U10066 (N_10066,N_7822,N_5189);
nand U10067 (N_10067,N_6568,N_6772);
or U10068 (N_10068,N_5418,N_6908);
or U10069 (N_10069,N_9078,N_5537);
or U10070 (N_10070,N_8334,N_7191);
and U10071 (N_10071,N_9782,N_9413);
nor U10072 (N_10072,N_7603,N_8349);
nor U10073 (N_10073,N_7463,N_8828);
nand U10074 (N_10074,N_9274,N_8792);
nor U10075 (N_10075,N_8302,N_6309);
or U10076 (N_10076,N_7849,N_6117);
nor U10077 (N_10077,N_5601,N_5468);
or U10078 (N_10078,N_9114,N_5360);
xor U10079 (N_10079,N_9151,N_8963);
nand U10080 (N_10080,N_8379,N_8776);
xnor U10081 (N_10081,N_9680,N_7717);
nor U10082 (N_10082,N_6785,N_8602);
xor U10083 (N_10083,N_5339,N_6135);
nor U10084 (N_10084,N_8020,N_7507);
nand U10085 (N_10085,N_6770,N_7571);
nand U10086 (N_10086,N_6062,N_9529);
nor U10087 (N_10087,N_5531,N_9170);
nor U10088 (N_10088,N_6963,N_8090);
nand U10089 (N_10089,N_5253,N_7696);
and U10090 (N_10090,N_8825,N_5449);
nand U10091 (N_10091,N_8863,N_7311);
nand U10092 (N_10092,N_9661,N_7949);
nor U10093 (N_10093,N_9684,N_5439);
xnor U10094 (N_10094,N_7200,N_6268);
or U10095 (N_10095,N_6561,N_9614);
and U10096 (N_10096,N_6842,N_5606);
and U10097 (N_10097,N_7780,N_9427);
or U10098 (N_10098,N_9545,N_8760);
or U10099 (N_10099,N_6192,N_6880);
nand U10100 (N_10100,N_6359,N_9653);
nor U10101 (N_10101,N_5045,N_9858);
xor U10102 (N_10102,N_8171,N_9867);
or U10103 (N_10103,N_6314,N_5669);
nand U10104 (N_10104,N_9321,N_9804);
xor U10105 (N_10105,N_6873,N_6447);
or U10106 (N_10106,N_6678,N_7560);
nand U10107 (N_10107,N_7941,N_7210);
or U10108 (N_10108,N_8260,N_9008);
nor U10109 (N_10109,N_9356,N_8912);
xor U10110 (N_10110,N_7414,N_6846);
xor U10111 (N_10111,N_8669,N_9281);
nand U10112 (N_10112,N_6265,N_8527);
nor U10113 (N_10113,N_5716,N_6702);
nor U10114 (N_10114,N_8870,N_9770);
nor U10115 (N_10115,N_8440,N_5917);
nor U10116 (N_10116,N_8552,N_6771);
nor U10117 (N_10117,N_5535,N_6895);
and U10118 (N_10118,N_6101,N_6625);
or U10119 (N_10119,N_8630,N_9419);
nor U10120 (N_10120,N_5272,N_8299);
xnor U10121 (N_10121,N_8980,N_8206);
nand U10122 (N_10122,N_7582,N_9999);
and U10123 (N_10123,N_8610,N_9310);
and U10124 (N_10124,N_8780,N_7224);
xnor U10125 (N_10125,N_9421,N_7115);
nor U10126 (N_10126,N_9983,N_6321);
nor U10127 (N_10127,N_7538,N_9298);
nor U10128 (N_10128,N_9442,N_7352);
xnor U10129 (N_10129,N_8730,N_8851);
and U10130 (N_10130,N_7336,N_7979);
nor U10131 (N_10131,N_7593,N_8782);
and U10132 (N_10132,N_8950,N_7077);
nand U10133 (N_10133,N_8317,N_9575);
or U10134 (N_10134,N_7319,N_6038);
nor U10135 (N_10135,N_5826,N_9479);
nand U10136 (N_10136,N_8094,N_7845);
or U10137 (N_10137,N_7756,N_5594);
nor U10138 (N_10138,N_7288,N_5931);
nor U10139 (N_10139,N_7028,N_6177);
xnor U10140 (N_10140,N_9380,N_9996);
and U10141 (N_10141,N_7905,N_7680);
nor U10142 (N_10142,N_9168,N_6685);
and U10143 (N_10143,N_5152,N_5024);
nand U10144 (N_10144,N_7164,N_9120);
and U10145 (N_10145,N_8964,N_8289);
nor U10146 (N_10146,N_8209,N_9888);
nand U10147 (N_10147,N_7720,N_9276);
xor U10148 (N_10148,N_9700,N_8453);
nor U10149 (N_10149,N_7497,N_7240);
and U10150 (N_10150,N_6807,N_8346);
nor U10151 (N_10151,N_9487,N_6696);
nor U10152 (N_10152,N_6097,N_5678);
nor U10153 (N_10153,N_6171,N_5065);
nor U10154 (N_10154,N_6869,N_5544);
nor U10155 (N_10155,N_9613,N_9252);
and U10156 (N_10156,N_6441,N_7241);
or U10157 (N_10157,N_8535,N_5703);
nand U10158 (N_10158,N_9000,N_7471);
nand U10159 (N_10159,N_6566,N_9594);
xor U10160 (N_10160,N_9205,N_8261);
or U10161 (N_10161,N_9169,N_7765);
xnor U10162 (N_10162,N_7809,N_9390);
nand U10163 (N_10163,N_8884,N_9404);
nand U10164 (N_10164,N_6835,N_8170);
and U10165 (N_10165,N_6460,N_6461);
or U10166 (N_10166,N_8575,N_9895);
nor U10167 (N_10167,N_9671,N_6667);
or U10168 (N_10168,N_6371,N_5769);
and U10169 (N_10169,N_5876,N_8650);
nand U10170 (N_10170,N_5635,N_9226);
or U10171 (N_10171,N_8338,N_9446);
nand U10172 (N_10172,N_8690,N_5393);
or U10173 (N_10173,N_5150,N_6626);
and U10174 (N_10174,N_5151,N_9569);
nand U10175 (N_10175,N_7098,N_6986);
nand U10176 (N_10176,N_7536,N_9727);
and U10177 (N_10177,N_6312,N_7082);
nor U10178 (N_10178,N_5881,N_5082);
and U10179 (N_10179,N_5293,N_7842);
nand U10180 (N_10180,N_8468,N_5160);
nor U10181 (N_10181,N_8273,N_7031);
nand U10182 (N_10182,N_6762,N_9737);
or U10183 (N_10183,N_5569,N_9182);
nor U10184 (N_10184,N_6436,N_6059);
nand U10185 (N_10185,N_5793,N_9813);
and U10186 (N_10186,N_5196,N_6692);
nor U10187 (N_10187,N_9944,N_8499);
or U10188 (N_10188,N_8378,N_8374);
nand U10189 (N_10189,N_9341,N_8558);
or U10190 (N_10190,N_6044,N_5178);
nand U10191 (N_10191,N_9324,N_5839);
nand U10192 (N_10192,N_6002,N_8968);
and U10193 (N_10193,N_5552,N_9918);
or U10194 (N_10194,N_5651,N_9773);
and U10195 (N_10195,N_9962,N_8428);
nand U10196 (N_10196,N_9577,N_9852);
nand U10197 (N_10197,N_7744,N_6623);
and U10198 (N_10198,N_9932,N_6402);
nand U10199 (N_10199,N_8739,N_8693);
nand U10200 (N_10200,N_7564,N_6683);
or U10201 (N_10201,N_7903,N_7770);
nor U10202 (N_10202,N_7273,N_7673);
or U10203 (N_10203,N_7931,N_9022);
or U10204 (N_10204,N_7214,N_6180);
or U10205 (N_10205,N_6643,N_7549);
nand U10206 (N_10206,N_7403,N_9993);
xnor U10207 (N_10207,N_5381,N_7938);
nand U10208 (N_10208,N_7628,N_8924);
nor U10209 (N_10209,N_5009,N_8114);
nand U10210 (N_10210,N_6875,N_9269);
nor U10211 (N_10211,N_5128,N_5423);
or U10212 (N_10212,N_8077,N_7394);
or U10213 (N_10213,N_5472,N_8603);
or U10214 (N_10214,N_7937,N_8894);
or U10215 (N_10215,N_6581,N_7529);
and U10216 (N_10216,N_7685,N_8612);
and U10217 (N_10217,N_8465,N_6348);
or U10218 (N_10218,N_7278,N_6489);
xor U10219 (N_10219,N_8305,N_8708);
nand U10220 (N_10220,N_7623,N_7189);
nand U10221 (N_10221,N_5999,N_8905);
nand U10222 (N_10222,N_8256,N_9722);
or U10223 (N_10223,N_5484,N_9534);
or U10224 (N_10224,N_6279,N_8557);
nor U10225 (N_10225,N_8581,N_8495);
nor U10226 (N_10226,N_6907,N_5820);
nor U10227 (N_10227,N_9611,N_7990);
nand U10228 (N_10228,N_9785,N_7650);
and U10229 (N_10229,N_9550,N_5825);
nor U10230 (N_10230,N_7943,N_9904);
and U10231 (N_10231,N_9872,N_8972);
xnor U10232 (N_10232,N_8052,N_9809);
or U10233 (N_10233,N_6629,N_9917);
xor U10234 (N_10234,N_5577,N_6464);
and U10235 (N_10235,N_8272,N_9103);
or U10236 (N_10236,N_9043,N_5366);
and U10237 (N_10237,N_8003,N_8173);
or U10238 (N_10238,N_5673,N_6700);
xnor U10239 (N_10239,N_6664,N_9842);
or U10240 (N_10240,N_9862,N_6400);
nor U10241 (N_10241,N_5210,N_6947);
and U10242 (N_10242,N_9827,N_6377);
or U10243 (N_10243,N_8647,N_5390);
nand U10244 (N_10244,N_6127,N_5315);
or U10245 (N_10245,N_5721,N_5890);
nand U10246 (N_10246,N_8526,N_6077);
nor U10247 (N_10247,N_6887,N_9081);
nor U10248 (N_10248,N_5020,N_7957);
or U10249 (N_10249,N_6537,N_7970);
nor U10250 (N_10250,N_8424,N_7936);
and U10251 (N_10251,N_7800,N_7426);
nand U10252 (N_10252,N_8534,N_9835);
xnor U10253 (N_10253,N_8885,N_8834);
or U10254 (N_10254,N_8692,N_8136);
nand U10255 (N_10255,N_9641,N_7178);
nand U10256 (N_10256,N_5772,N_5333);
nand U10257 (N_10257,N_5075,N_7841);
nand U10258 (N_10258,N_6426,N_6946);
or U10259 (N_10259,N_7651,N_7611);
and U10260 (N_10260,N_5136,N_6933);
xor U10261 (N_10261,N_9967,N_7149);
nor U10262 (N_10262,N_7901,N_9542);
nor U10263 (N_10263,N_5149,N_5628);
nand U10264 (N_10264,N_8085,N_7889);
nand U10265 (N_10265,N_9712,N_8662);
nor U10266 (N_10266,N_6641,N_6648);
nand U10267 (N_10267,N_5907,N_5170);
and U10268 (N_10268,N_8039,N_6805);
nand U10269 (N_10269,N_8127,N_5164);
nand U10270 (N_10270,N_9985,N_6480);
and U10271 (N_10271,N_6450,N_6572);
or U10272 (N_10272,N_5522,N_7425);
nand U10273 (N_10273,N_5636,N_6379);
and U10274 (N_10274,N_8799,N_9672);
or U10275 (N_10275,N_9297,N_8771);
and U10276 (N_10276,N_7345,N_6316);
or U10277 (N_10277,N_6288,N_9316);
and U10278 (N_10278,N_7550,N_8936);
nand U10279 (N_10279,N_7368,N_9431);
or U10280 (N_10280,N_7775,N_6134);
nand U10281 (N_10281,N_7776,N_8995);
or U10282 (N_10282,N_5966,N_5733);
nand U10283 (N_10283,N_9174,N_9202);
or U10284 (N_10284,N_9301,N_5123);
nor U10285 (N_10285,N_5148,N_6756);
nand U10286 (N_10286,N_7328,N_6949);
and U10287 (N_10287,N_5300,N_6118);
and U10288 (N_10288,N_9216,N_8507);
nor U10289 (N_10289,N_9167,N_5791);
nor U10290 (N_10290,N_6226,N_8831);
or U10291 (N_10291,N_7927,N_9923);
nor U10292 (N_10292,N_6191,N_5956);
nor U10293 (N_10293,N_9503,N_7334);
or U10294 (N_10294,N_7642,N_6677);
and U10295 (N_10295,N_6405,N_8986);
nor U10296 (N_10296,N_9949,N_8759);
nand U10297 (N_10297,N_9497,N_6124);
nand U10298 (N_10298,N_5982,N_9035);
xor U10299 (N_10299,N_8627,N_5514);
and U10300 (N_10300,N_8767,N_5250);
nor U10301 (N_10301,N_5974,N_8586);
nand U10302 (N_10302,N_6746,N_6380);
nand U10303 (N_10303,N_7589,N_8975);
and U10304 (N_10304,N_9473,N_9148);
and U10305 (N_10305,N_9368,N_6952);
and U10306 (N_10306,N_9335,N_7600);
nor U10307 (N_10307,N_7857,N_5550);
or U10308 (N_10308,N_5835,N_9500);
and U10309 (N_10309,N_9769,N_6126);
nand U10310 (N_10310,N_8128,N_9732);
nand U10311 (N_10311,N_5896,N_8354);
nor U10312 (N_10312,N_8977,N_7411);
xor U10313 (N_10313,N_7689,N_9760);
or U10314 (N_10314,N_5183,N_8725);
nor U10315 (N_10315,N_5072,N_7653);
or U10316 (N_10316,N_6597,N_9571);
and U10317 (N_10317,N_7478,N_9398);
or U10318 (N_10318,N_5770,N_9012);
or U10319 (N_10319,N_5489,N_8313);
nor U10320 (N_10320,N_9747,N_5645);
and U10321 (N_10321,N_5041,N_8853);
xor U10322 (N_10322,N_8304,N_5586);
and U10323 (N_10323,N_9441,N_6219);
and U10324 (N_10324,N_7535,N_7338);
nand U10325 (N_10325,N_6529,N_5370);
or U10326 (N_10326,N_6215,N_7473);
nand U10327 (N_10327,N_7062,N_8595);
or U10328 (N_10328,N_9898,N_7452);
nor U10329 (N_10329,N_6853,N_7634);
or U10330 (N_10330,N_8382,N_8318);
and U10331 (N_10331,N_8350,N_7525);
and U10332 (N_10332,N_9319,N_6631);
nand U10333 (N_10333,N_8518,N_8504);
or U10334 (N_10334,N_5749,N_7147);
or U10335 (N_10335,N_5022,N_9919);
or U10336 (N_10336,N_5199,N_8658);
nor U10337 (N_10337,N_5412,N_6128);
or U10338 (N_10338,N_6153,N_9171);
and U10339 (N_10339,N_8655,N_8904);
or U10340 (N_10340,N_6094,N_7299);
xor U10341 (N_10341,N_7724,N_9041);
nand U10342 (N_10342,N_7044,N_9403);
xor U10343 (N_10343,N_9338,N_5480);
and U10344 (N_10344,N_8031,N_5130);
or U10345 (N_10345,N_9303,N_5702);
nand U10346 (N_10346,N_8930,N_6502);
nand U10347 (N_10347,N_5388,N_6123);
nand U10348 (N_10348,N_9055,N_5098);
xor U10349 (N_10349,N_9652,N_6145);
and U10350 (N_10350,N_9519,N_7312);
nor U10351 (N_10351,N_7699,N_5868);
and U10352 (N_10352,N_6711,N_7469);
nand U10353 (N_10353,N_8796,N_6722);
nor U10354 (N_10354,N_5071,N_6747);
and U10355 (N_10355,N_6372,N_5394);
nand U10356 (N_10356,N_7706,N_5052);
or U10357 (N_10357,N_6200,N_6512);
nand U10358 (N_10358,N_7774,N_8666);
or U10359 (N_10359,N_8190,N_8893);
xnor U10360 (N_10360,N_7517,N_8282);
or U10361 (N_10361,N_6090,N_6847);
nand U10362 (N_10362,N_8861,N_7930);
or U10363 (N_10363,N_5105,N_5371);
nand U10364 (N_10364,N_9211,N_6340);
or U10365 (N_10365,N_6198,N_8177);
and U10366 (N_10366,N_7193,N_5346);
nor U10367 (N_10367,N_6043,N_6858);
and U10368 (N_10368,N_6110,N_9411);
and U10369 (N_10369,N_5943,N_7423);
nand U10370 (N_10370,N_9578,N_6286);
nor U10371 (N_10371,N_7045,N_7122);
nand U10372 (N_10372,N_9030,N_9708);
nor U10373 (N_10373,N_9027,N_9444);
nor U10374 (N_10374,N_7350,N_5368);
nand U10375 (N_10375,N_8793,N_9891);
and U10376 (N_10376,N_9663,N_9296);
or U10377 (N_10377,N_6428,N_9137);
or U10378 (N_10378,N_5551,N_8989);
and U10379 (N_10379,N_7382,N_8340);
nor U10380 (N_10380,N_9802,N_5103);
nand U10381 (N_10381,N_7050,N_9948);
or U10382 (N_10382,N_8048,N_5997);
or U10383 (N_10383,N_7808,N_5975);
or U10384 (N_10384,N_7356,N_8813);
nor U10385 (N_10385,N_6891,N_8211);
and U10386 (N_10386,N_7834,N_6015);
nor U10387 (N_10387,N_7435,N_7144);
or U10388 (N_10388,N_5362,N_8142);
or U10389 (N_10389,N_6632,N_5915);
nand U10390 (N_10390,N_8914,N_5297);
or U10391 (N_10391,N_5725,N_8290);
or U10392 (N_10392,N_5837,N_7992);
or U10393 (N_10393,N_6270,N_6374);
nor U10394 (N_10394,N_9566,N_5078);
nor U10395 (N_10395,N_7461,N_5374);
nand U10396 (N_10396,N_5989,N_8899);
xor U10397 (N_10397,N_7998,N_9378);
and U10398 (N_10398,N_7054,N_5765);
nor U10399 (N_10399,N_7534,N_7935);
nand U10400 (N_10400,N_6248,N_6291);
or U10401 (N_10401,N_8033,N_8179);
nand U10402 (N_10402,N_5990,N_7121);
and U10403 (N_10403,N_9123,N_6105);
and U10404 (N_10404,N_6560,N_8888);
or U10405 (N_10405,N_9655,N_5444);
nand U10406 (N_10406,N_9619,N_9394);
and U10407 (N_10407,N_5181,N_5802);
and U10408 (N_10408,N_5838,N_9336);
nand U10409 (N_10409,N_5467,N_6652);
or U10410 (N_10410,N_6125,N_5572);
nand U10411 (N_10411,N_8006,N_9306);
nor U10412 (N_10412,N_9754,N_8865);
nand U10413 (N_10413,N_6948,N_7939);
and U10414 (N_10414,N_9510,N_7914);
and U10415 (N_10415,N_5220,N_5013);
and U10416 (N_10416,N_7856,N_5967);
or U10417 (N_10417,N_8448,N_9789);
nor U10418 (N_10418,N_9465,N_8176);
nor U10419 (N_10419,N_5545,N_5100);
nand U10420 (N_10420,N_9406,N_7391);
xnor U10421 (N_10421,N_9443,N_5163);
nor U10422 (N_10422,N_5364,N_5515);
xnor U10423 (N_10423,N_8234,N_7295);
and U10424 (N_10424,N_9219,N_6010);
nand U10425 (N_10425,N_6619,N_9963);
or U10426 (N_10426,N_7485,N_7103);
nand U10427 (N_10427,N_9957,N_5165);
and U10428 (N_10428,N_9612,N_6705);
xnor U10429 (N_10429,N_9593,N_8554);
nand U10430 (N_10430,N_6578,N_5897);
or U10431 (N_10431,N_5027,N_5146);
nor U10432 (N_10432,N_9902,N_7095);
and U10433 (N_10433,N_9920,N_6555);
nand U10434 (N_10434,N_9248,N_6956);
nor U10435 (N_10435,N_8860,N_6527);
or U10436 (N_10436,N_6073,N_5532);
nor U10437 (N_10437,N_7047,N_9812);
or U10438 (N_10438,N_6828,N_6591);
xnor U10439 (N_10439,N_5326,N_6544);
nor U10440 (N_10440,N_5275,N_9127);
nor U10441 (N_10441,N_5910,N_7844);
and U10442 (N_10442,N_8482,N_5980);
or U10443 (N_10443,N_5466,N_7137);
or U10444 (N_10444,N_7397,N_8103);
nand U10445 (N_10445,N_9292,N_7329);
and U10446 (N_10446,N_9975,N_9721);
xnor U10447 (N_10447,N_8611,N_5824);
xnor U10448 (N_10448,N_7942,N_5026);
or U10449 (N_10449,N_9834,N_7041);
nor U10450 (N_10450,N_9866,N_6491);
or U10451 (N_10451,N_8629,N_5707);
xor U10452 (N_10452,N_8976,N_5805);
nand U10453 (N_10453,N_9504,N_5406);
xor U10454 (N_10454,N_9665,N_5332);
xnor U10455 (N_10455,N_8714,N_8410);
or U10456 (N_10456,N_6188,N_8472);
nand U10457 (N_10457,N_8752,N_8119);
and U10458 (N_10458,N_8425,N_9340);
and U10459 (N_10459,N_9807,N_7037);
and U10460 (N_10460,N_8874,N_7313);
nand U10461 (N_10461,N_7799,N_5887);
nor U10462 (N_10462,N_7038,N_6453);
nor U10463 (N_10463,N_9971,N_5252);
nand U10464 (N_10464,N_6350,N_6583);
and U10465 (N_10465,N_7718,N_9230);
and U10466 (N_10466,N_5036,N_6539);
or U10467 (N_10467,N_9313,N_6334);
or U10468 (N_10468,N_8212,N_5950);
xor U10469 (N_10469,N_6325,N_8113);
and U10470 (N_10470,N_7399,N_8798);
nor U10471 (N_10471,N_6909,N_7255);
nand U10472 (N_10472,N_9913,N_9283);
nor U10473 (N_10473,N_6837,N_9318);
nand U10474 (N_10474,N_5946,N_6076);
and U10475 (N_10475,N_7663,N_9689);
or U10476 (N_10476,N_5134,N_7183);
nand U10477 (N_10477,N_8707,N_8058);
nand U10478 (N_10478,N_9131,N_9644);
nand U10479 (N_10479,N_7275,N_5007);
xor U10480 (N_10480,N_9110,N_6695);
nor U10481 (N_10481,N_8392,N_9587);
and U10482 (N_10482,N_7987,N_6413);
or U10483 (N_10483,N_6342,N_7872);
or U10484 (N_10484,N_6384,N_8291);
and U10485 (N_10485,N_5383,N_7173);
nand U10486 (N_10486,N_8065,N_5619);
nand U10487 (N_10487,N_8651,N_7972);
and U10488 (N_10488,N_6690,N_6423);
and U10489 (N_10489,N_8901,N_6034);
nand U10490 (N_10490,N_6704,N_6944);
xnor U10491 (N_10491,N_6363,N_5867);
nor U10492 (N_10492,N_6150,N_7766);
nor U10493 (N_10493,N_6030,N_9024);
nand U10494 (N_10494,N_5631,N_6037);
or U10495 (N_10495,N_5386,N_5548);
and U10496 (N_10496,N_9931,N_5743);
and U10497 (N_10497,N_7684,N_9477);
and U10498 (N_10498,N_7969,N_7755);
nand U10499 (N_10499,N_6993,N_6792);
nand U10500 (N_10500,N_6758,N_9549);
and U10501 (N_10501,N_6531,N_9498);
nand U10502 (N_10502,N_6144,N_7180);
nor U10503 (N_10503,N_8892,N_7616);
xor U10504 (N_10504,N_8697,N_5169);
and U10505 (N_10505,N_6019,N_8040);
nor U10506 (N_10506,N_8089,N_7917);
xor U10507 (N_10507,N_9476,N_5992);
xor U10508 (N_10508,N_5447,N_5546);
nand U10509 (N_10509,N_9555,N_6614);
nor U10510 (N_10510,N_6295,N_6440);
xor U10511 (N_10511,N_9753,N_8722);
and U10512 (N_10512,N_7035,N_7817);
xor U10513 (N_10513,N_5983,N_8164);
nor U10514 (N_10514,N_5140,N_8947);
nor U10515 (N_10515,N_7661,N_6618);
and U10516 (N_10516,N_8862,N_6033);
and U10517 (N_10517,N_5538,N_5477);
nand U10518 (N_10518,N_9004,N_9126);
and U10519 (N_10519,N_8606,N_6504);
and U10520 (N_10520,N_8622,N_6913);
or U10521 (N_10521,N_6027,N_7540);
nand U10522 (N_10522,N_6404,N_6175);
or U10523 (N_10523,N_8116,N_7881);
or U10524 (N_10524,N_6760,N_7645);
xnor U10525 (N_10525,N_5351,N_9134);
nand U10526 (N_10526,N_7036,N_7552);
and U10527 (N_10527,N_9149,N_7168);
xnor U10528 (N_10528,N_8510,N_8918);
nor U10529 (N_10529,N_6341,N_8092);
or U10530 (N_10530,N_5675,N_7043);
nor U10531 (N_10531,N_7209,N_9883);
xnor U10532 (N_10532,N_9977,N_9639);
xor U10533 (N_10533,N_6203,N_9193);
nor U10534 (N_10534,N_9270,N_8568);
or U10535 (N_10535,N_8956,N_9188);
and U10536 (N_10536,N_9871,N_5690);
xor U10537 (N_10537,N_8498,N_6308);
or U10538 (N_10538,N_5399,N_5937);
nand U10539 (N_10539,N_8230,N_7456);
or U10540 (N_10540,N_7353,N_9466);
and U10541 (N_10541,N_6416,N_5303);
nor U10542 (N_10542,N_6048,N_6103);
or U10543 (N_10543,N_9738,N_6032);
and U10544 (N_10544,N_5508,N_6600);
or U10545 (N_10545,N_7530,N_7480);
nand U10546 (N_10546,N_8395,N_6471);
and U10547 (N_10547,N_9943,N_8357);
or U10548 (N_10548,N_6920,N_8954);
and U10549 (N_10549,N_9670,N_8270);
or U10550 (N_10550,N_9414,N_8998);
or U10551 (N_10551,N_5880,N_9096);
or U10552 (N_10552,N_9181,N_9668);
nor U10553 (N_10553,N_9065,N_6222);
and U10554 (N_10554,N_6483,N_7988);
or U10555 (N_10555,N_9713,N_6719);
xor U10556 (N_10556,N_5435,N_9750);
or U10557 (N_10557,N_6082,N_6885);
or U10558 (N_10558,N_5384,N_5575);
and U10559 (N_10559,N_6894,N_8750);
or U10560 (N_10560,N_6451,N_8531);
or U10561 (N_10561,N_9304,N_5789);
xor U10562 (N_10562,N_8503,N_8803);
nand U10563 (N_10563,N_5495,N_8188);
or U10564 (N_10564,N_7464,N_9720);
and U10565 (N_10565,N_6759,N_6638);
or U10566 (N_10566,N_9927,N_8895);
nand U10567 (N_10567,N_5207,N_5778);
and U10568 (N_10568,N_8900,N_6443);
nand U10569 (N_10569,N_8247,N_6630);
or U10570 (N_10570,N_5595,N_7816);
xnor U10571 (N_10571,N_9574,N_6006);
nor U10572 (N_10572,N_5347,N_5091);
or U10573 (N_10573,N_9660,N_7639);
nor U10574 (N_10574,N_5832,N_9115);
or U10575 (N_10575,N_8208,N_5664);
nand U10576 (N_10576,N_5948,N_9635);
and U10577 (N_10577,N_5227,N_5391);
nand U10578 (N_10578,N_6358,N_7308);
and U10579 (N_10579,N_5236,N_8073);
or U10580 (N_10580,N_7398,N_5358);
or U10581 (N_10581,N_9261,N_8541);
and U10582 (N_10582,N_7358,N_9308);
nor U10583 (N_10583,N_9496,N_8162);
and U10584 (N_10584,N_6823,N_7741);
and U10585 (N_10585,N_5836,N_9348);
or U10586 (N_10586,N_5557,N_6878);
nand U10587 (N_10587,N_8081,N_8361);
or U10588 (N_10588,N_5884,N_6780);
nor U10589 (N_10589,N_7270,N_9490);
nor U10590 (N_10590,N_8841,N_8511);
nor U10591 (N_10591,N_8698,N_6565);
xor U10592 (N_10592,N_6868,N_9818);
and U10593 (N_10593,N_7479,N_5885);
nor U10594 (N_10594,N_5436,N_9705);
xor U10595 (N_10595,N_7567,N_5913);
or U10596 (N_10596,N_5099,N_7204);
nor U10597 (N_10597,N_5774,N_7871);
nor U10598 (N_10598,N_6872,N_7418);
xnor U10599 (N_10599,N_6636,N_7379);
or U10600 (N_10600,N_5963,N_9586);
or U10601 (N_10601,N_9630,N_6906);
or U10602 (N_10602,N_8580,N_5790);
and U10603 (N_10603,N_6803,N_7813);
or U10604 (N_10604,N_5785,N_6959);
and U10605 (N_10605,N_5108,N_6433);
nand U10606 (N_10606,N_6115,N_9268);
nand U10607 (N_10607,N_5739,N_7052);
and U10608 (N_10608,N_6294,N_9197);
and U10609 (N_10609,N_6310,N_8307);
and U10610 (N_10610,N_7725,N_6796);
nand U10611 (N_10611,N_5563,N_9887);
xnor U10612 (N_10612,N_6850,N_9099);
and U10613 (N_10613,N_8011,N_5767);
and U10614 (N_10614,N_8949,N_6257);
or U10615 (N_10615,N_9023,N_5747);
or U10616 (N_10616,N_6376,N_8002);
nand U10617 (N_10617,N_7421,N_8644);
or U10618 (N_10618,N_7120,N_7453);
nand U10619 (N_10619,N_9777,N_7437);
or U10620 (N_10620,N_7400,N_7460);
and U10621 (N_10621,N_8107,N_8087);
and U10622 (N_10622,N_8288,N_8161);
nor U10623 (N_10623,N_7928,N_9145);
nor U10624 (N_10624,N_7683,N_5660);
or U10625 (N_10625,N_5705,N_5102);
nand U10626 (N_10626,N_7226,N_8564);
or U10627 (N_10627,N_9050,N_7501);
or U10628 (N_10628,N_9102,N_9486);
nand U10629 (N_10629,N_6370,N_8044);
or U10630 (N_10630,N_6201,N_8845);
or U10631 (N_10631,N_6212,N_7784);
nor U10632 (N_10632,N_7487,N_8263);
and U10633 (N_10633,N_9288,N_5902);
nor U10634 (N_10634,N_6463,N_5014);
or U10635 (N_10635,N_6929,N_8559);
and U10636 (N_10636,N_8470,N_6352);
or U10637 (N_10637,N_7363,N_7907);
or U10638 (N_10638,N_8399,N_6486);
or U10639 (N_10639,N_8156,N_8858);
nand U10640 (N_10640,N_7341,N_8483);
nand U10641 (N_10641,N_5206,N_6674);
nor U10642 (N_10642,N_6691,N_8365);
nand U10643 (N_10643,N_8372,N_7627);
nand U10644 (N_10644,N_7910,N_7443);
and U10645 (N_10645,N_5922,N_6111);
xnor U10646 (N_10646,N_5679,N_5302);
nand U10647 (N_10647,N_8032,N_9787);
nand U10648 (N_10648,N_9860,N_5081);
xor U10649 (N_10649,N_8054,N_8015);
nor U10650 (N_10650,N_6981,N_7865);
nand U10651 (N_10651,N_8567,N_8939);
or U10652 (N_10652,N_7804,N_5061);
nand U10653 (N_10653,N_9793,N_8454);
nor U10654 (N_10654,N_7073,N_5620);
nor U10655 (N_10655,N_9839,N_9909);
or U10656 (N_10656,N_9189,N_9535);
and U10657 (N_10657,N_8922,N_8336);
nand U10658 (N_10658,N_6680,N_8833);
and U10659 (N_10659,N_6501,N_5173);
nand U10660 (N_10660,N_8458,N_8220);
and U10661 (N_10661,N_7503,N_8367);
or U10662 (N_10662,N_7626,N_7326);
nand U10663 (N_10663,N_5414,N_5018);
xnor U10664 (N_10664,N_9259,N_8958);
nand U10665 (N_10665,N_8943,N_7575);
nand U10666 (N_10666,N_5086,N_6132);
nand U10667 (N_10667,N_9725,N_6167);
nand U10668 (N_10668,N_9964,N_9258);
and U10669 (N_10669,N_8484,N_5540);
nand U10670 (N_10670,N_7013,N_8800);
xnor U10671 (N_10671,N_9560,N_6739);
xor U10672 (N_10672,N_9426,N_8388);
or U10673 (N_10673,N_5638,N_9666);
and U10674 (N_10674,N_7649,N_9850);
or U10675 (N_10675,N_7475,N_9869);
and U10676 (N_10676,N_5715,N_9204);
or U10677 (N_10677,N_9138,N_8520);
and U10678 (N_10678,N_7511,N_7387);
nand U10679 (N_10679,N_9597,N_7873);
nand U10680 (N_10680,N_9989,N_9646);
and U10681 (N_10681,N_6068,N_6179);
or U10682 (N_10682,N_5849,N_9121);
or U10683 (N_10683,N_7974,N_7778);
or U10684 (N_10684,N_9798,N_7946);
or U10685 (N_10685,N_9016,N_6156);
and U10686 (N_10686,N_8331,N_7823);
nor U10687 (N_10687,N_5201,N_7012);
or U10688 (N_10688,N_8859,N_8815);
nand U10689 (N_10689,N_8101,N_8443);
nor U10690 (N_10690,N_5779,N_6801);
nand U10691 (N_10691,N_5677,N_8434);
nor U10692 (N_10692,N_5166,N_9714);
nor U10693 (N_10693,N_8878,N_7408);
nand U10694 (N_10694,N_8284,N_7558);
nor U10695 (N_10695,N_6154,N_9676);
and U10696 (N_10696,N_6980,N_5464);
or U10697 (N_10697,N_6496,N_7030);
xnor U10698 (N_10698,N_7547,N_6896);
nor U10699 (N_10699,N_7848,N_5336);
xnor U10700 (N_10700,N_5698,N_8952);
or U10701 (N_10701,N_8005,N_7459);
nand U10702 (N_10702,N_7257,N_7569);
nand U10703 (N_10703,N_5727,N_7991);
and U10704 (N_10704,N_8642,N_5794);
or U10705 (N_10705,N_7314,N_5908);
nand U10706 (N_10706,N_5787,N_6883);
nor U10707 (N_10707,N_5734,N_9354);
or U10708 (N_10708,N_5592,N_5800);
or U10709 (N_10709,N_7025,N_5259);
nand U10710 (N_10710,N_8460,N_5389);
or U10711 (N_10711,N_6515,N_7591);
and U10712 (N_10712,N_8778,N_9744);
and U10713 (N_10713,N_5258,N_8225);
nand U10714 (N_10714,N_9241,N_8413);
nand U10715 (N_10715,N_5046,N_7419);
or U10716 (N_10716,N_5006,N_7735);
nand U10717 (N_10717,N_9514,N_9930);
and U10718 (N_10718,N_7108,N_8358);
xor U10719 (N_10719,N_5987,N_5474);
and U10720 (N_10720,N_5205,N_6892);
or U10721 (N_10721,N_9565,N_8838);
xor U10722 (N_10722,N_8529,N_8069);
or U10723 (N_10723,N_7968,N_7710);
nor U10724 (N_10724,N_6616,N_6378);
nor U10725 (N_10725,N_8830,N_5962);
nor U10726 (N_10726,N_8213,N_5854);
or U10727 (N_10727,N_9290,N_8896);
nand U10728 (N_10728,N_9453,N_6777);
or U10729 (N_10729,N_5615,N_9637);
xnor U10730 (N_10730,N_7428,N_8231);
nor U10731 (N_10731,N_5017,N_8618);
and U10732 (N_10732,N_9075,N_7597);
or U10733 (N_10733,N_9408,N_9781);
nand U10734 (N_10734,N_6456,N_9522);
xnor U10735 (N_10735,N_8764,N_7742);
and U10736 (N_10736,N_7232,N_7631);
nor U10737 (N_10737,N_7143,N_8934);
nor U10738 (N_10738,N_8232,N_7114);
nor U10739 (N_10739,N_6987,N_8186);
nand U10740 (N_10740,N_9623,N_8017);
nand U10741 (N_10741,N_9130,N_7715);
and U10742 (N_10742,N_6978,N_5930);
nand U10743 (N_10743,N_5891,N_9645);
or U10744 (N_10744,N_5209,N_7693);
or U10745 (N_10745,N_6732,N_6173);
nand U10746 (N_10746,N_7965,N_8241);
nand U10747 (N_10747,N_9783,N_5775);
or U10748 (N_10748,N_7151,N_7213);
and U10749 (N_10749,N_7258,N_7339);
or U10750 (N_10750,N_5417,N_9831);
nand U10751 (N_10751,N_9589,N_7899);
nand U10752 (N_10752,N_7934,N_6001);
nand U10753 (N_10753,N_7094,N_7267);
or U10754 (N_10754,N_8391,N_8632);
or U10755 (N_10755,N_5019,N_7205);
and U10756 (N_10756,N_7837,N_6141);
nor U10757 (N_10757,N_6914,N_8636);
or U10758 (N_10758,N_8192,N_5356);
or U10759 (N_10759,N_8362,N_8789);
xnor U10760 (N_10760,N_5198,N_9071);
and U10761 (N_10761,N_5329,N_9209);
xnor U10762 (N_10762,N_5057,N_5858);
or U10763 (N_10763,N_7148,N_7282);
xor U10764 (N_10764,N_9876,N_9245);
nor U10765 (N_10765,N_5583,N_9762);
nor U10766 (N_10766,N_9854,N_9579);
or U10767 (N_10767,N_5053,N_8463);
nand U10768 (N_10768,N_8246,N_9328);
and U10769 (N_10769,N_7883,N_7633);
or U10770 (N_10770,N_6833,N_5043);
nand U10771 (N_10771,N_5613,N_7434);
nand U10772 (N_10772,N_7602,N_8166);
nand U10773 (N_10773,N_5877,N_7365);
nor U10774 (N_10774,N_8000,N_9031);
and U10775 (N_10775,N_9820,N_5899);
and U10776 (N_10776,N_6347,N_6588);
nand U10777 (N_10777,N_5947,N_5093);
nand U10778 (N_10778,N_8821,N_5564);
nor U10779 (N_10779,N_8210,N_8446);
nor U10780 (N_10780,N_9701,N_6481);
and U10781 (N_10781,N_5708,N_7483);
nor U10782 (N_10782,N_8826,N_6324);
xor U10783 (N_10783,N_5429,N_7019);
or U10784 (N_10784,N_7732,N_5518);
xor U10785 (N_10785,N_9799,N_9936);
and U10786 (N_10786,N_7113,N_8088);
nand U10787 (N_10787,N_8222,N_6932);
nor U10788 (N_10788,N_8047,N_8363);
or U10789 (N_10789,N_7445,N_8721);
nor U10790 (N_10790,N_5728,N_8133);
and U10791 (N_10791,N_6707,N_9585);
nand U10792 (N_10792,N_5382,N_6882);
nor U10793 (N_10793,N_6970,N_6148);
or U10794 (N_10794,N_5203,N_6196);
or U10795 (N_10795,N_8699,N_7430);
xor U10796 (N_10796,N_6227,N_7736);
xor U10797 (N_10797,N_9464,N_5010);
nand U10798 (N_10798,N_6681,N_8734);
and U10799 (N_10799,N_6036,N_5612);
or U10800 (N_10800,N_6752,N_6795);
and U10801 (N_10801,N_6553,N_6710);
nand U10802 (N_10802,N_7730,N_6615);
nor U10803 (N_10803,N_7230,N_6296);
nand U10804 (N_10804,N_7932,N_6589);
xor U10805 (N_10805,N_5050,N_7954);
or U10806 (N_10806,N_5295,N_8794);
or U10807 (N_10807,N_7690,N_6439);
nand U10808 (N_10808,N_7208,N_7220);
nor U10809 (N_10809,N_7034,N_9108);
nand U10810 (N_10810,N_5005,N_7973);
nand U10811 (N_10811,N_8064,N_6160);
nand U10812 (N_10812,N_5961,N_8181);
nand U10813 (N_10813,N_5355,N_6449);
nand U10814 (N_10814,N_5330,N_6113);
nand U10815 (N_10815,N_8928,N_9360);
and U10816 (N_10816,N_5582,N_8566);
nor U10817 (N_10817,N_7177,N_5556);
nor U10818 (N_10818,N_5895,N_9568);
and U10819 (N_10819,N_8201,N_6509);
nand U10820 (N_10820,N_9588,N_7758);
or U10821 (N_10821,N_9771,N_8041);
or U10822 (N_10822,N_6992,N_9199);
nor U10823 (N_10823,N_5892,N_8070);
and U10824 (N_10824,N_7513,N_6183);
nor U10825 (N_10825,N_8386,N_9890);
or U10826 (N_10826,N_5589,N_8328);
xor U10827 (N_10827,N_6493,N_9385);
and U10828 (N_10828,N_9235,N_6716);
nor U10829 (N_10829,N_5457,N_8295);
or U10830 (N_10830,N_7022,N_9692);
nand U10831 (N_10831,N_7559,N_8748);
xor U10832 (N_10832,N_5200,N_9352);
and U10833 (N_10833,N_6210,N_9604);
nand U10834 (N_10834,N_8663,N_5424);
xor U10835 (N_10835,N_8745,N_9749);
or U10836 (N_10836,N_6635,N_8808);
or U10837 (N_10837,N_7796,N_8123);
xor U10838 (N_10838,N_9778,N_8303);
nand U10839 (N_10839,N_8496,N_9563);
nor U10840 (N_10840,N_7640,N_8719);
nand U10841 (N_10841,N_5861,N_8251);
and U10842 (N_10842,N_5257,N_6810);
xor U10843 (N_10843,N_5062,N_8917);
nand U10844 (N_10844,N_7893,N_8513);
and U10845 (N_10845,N_7118,N_8716);
nand U10846 (N_10846,N_9609,N_7862);
nor U10847 (N_10847,N_7373,N_8193);
and U10848 (N_10848,N_6437,N_8550);
nor U10849 (N_10849,N_8660,N_8276);
or U10850 (N_10850,N_6706,N_6238);
and U10851 (N_10851,N_6564,N_5426);
nand U10852 (N_10852,N_7604,N_8323);
nand U10853 (N_10853,N_6311,N_5590);
nand U10854 (N_10854,N_5519,N_5331);
nand U10855 (N_10855,N_5344,N_8971);
or U10856 (N_10856,N_7064,N_5630);
or U10857 (N_10857,N_8674,N_9667);
nand U10858 (N_10858,N_5037,N_7153);
and U10859 (N_10859,N_6283,N_7196);
and U10860 (N_10860,N_8664,N_5314);
nand U10861 (N_10861,N_7201,N_5215);
or U10862 (N_10862,N_9469,N_9758);
xnor U10863 (N_10863,N_6231,N_8140);
or U10864 (N_10864,N_5661,N_6519);
xor U10865 (N_10865,N_9657,N_7017);
nand U10866 (N_10866,N_8151,N_5247);
and U10867 (N_10867,N_8754,N_8593);
or U10868 (N_10868,N_9353,N_7068);
or U10869 (N_10869,N_9140,N_5754);
and U10870 (N_10870,N_5398,N_6438);
or U10871 (N_10871,N_6943,N_6202);
nor U10872 (N_10872,N_6745,N_9885);
and U10873 (N_10873,N_5847,N_5924);
and U10874 (N_10874,N_9906,N_8829);
and U10875 (N_10875,N_8111,N_9287);
or U10876 (N_10876,N_6557,N_5752);
and U10877 (N_10877,N_6620,N_5000);
and U10878 (N_10878,N_6014,N_5706);
or U10879 (N_10879,N_7665,N_5274);
xor U10880 (N_10880,N_5534,N_9133);
xor U10881 (N_10881,N_5030,N_8620);
and U10882 (N_10882,N_9200,N_7076);
xnor U10883 (N_10883,N_9648,N_8837);
or U10884 (N_10884,N_9719,N_7056);
or U10885 (N_10885,N_8880,N_7409);
nor U10886 (N_10886,N_9364,N_7268);
nor U10887 (N_10887,N_6302,N_7099);
or U10888 (N_10888,N_5283,N_6816);
and U10889 (N_10889,N_9755,N_5353);
and U10890 (N_10890,N_9495,N_7746);
xor U10891 (N_10891,N_9673,N_6213);
and U10892 (N_10892,N_6763,N_7854);
and U10893 (N_10893,N_5811,N_8777);
nor U10894 (N_10894,N_5299,N_7083);
and U10895 (N_10895,N_7337,N_7859);
or U10896 (N_10896,N_7502,N_8824);
nor U10897 (N_10897,N_8371,N_6181);
xor U10898 (N_10898,N_9581,N_6187);
or U10899 (N_10899,N_9201,N_5576);
nand U10900 (N_10900,N_9329,N_8763);
xor U10901 (N_10901,N_8668,N_7726);
and U10902 (N_10902,N_7199,N_7285);
and U10903 (N_10903,N_6806,N_5973);
nand U10904 (N_10904,N_8978,N_8624);
nand U10905 (N_10905,N_9966,N_5485);
nor U10906 (N_10906,N_8180,N_5001);
nor U10907 (N_10907,N_8816,N_8906);
nor U10908 (N_10908,N_6092,N_9695);
and U10909 (N_10909,N_9622,N_5421);
or U10910 (N_10910,N_5969,N_7924);
nor U10911 (N_10911,N_6275,N_6934);
nor U10912 (N_10912,N_6052,N_9584);
nand U10913 (N_10913,N_6817,N_9617);
nand U10914 (N_10914,N_9649,N_5354);
xnor U10915 (N_10915,N_7779,N_7745);
nand U10916 (N_10916,N_5505,N_7950);
and U10917 (N_10917,N_8732,N_5883);
nand U10918 (N_10918,N_9074,N_9709);
and U10919 (N_10919,N_8056,N_8628);
nand U10920 (N_10920,N_6856,N_5936);
nand U10921 (N_10921,N_6389,N_6356);
or U10922 (N_10922,N_6787,N_9236);
or U10923 (N_10923,N_6604,N_8417);
and U10924 (N_10924,N_7999,N_8359);
and U10925 (N_10925,N_9247,N_7847);
or U10926 (N_10926,N_7005,N_8987);
nor U10927 (N_10927,N_9129,N_7436);
or U10928 (N_10928,N_9210,N_6108);
nand U10929 (N_10929,N_7986,N_8265);
nand U10930 (N_10930,N_7727,N_6608);
or U10931 (N_10931,N_5919,N_9315);
and U10932 (N_10932,N_8174,N_9032);
and U10933 (N_10933,N_9806,N_7666);
or U10934 (N_10934,N_8437,N_5316);
and U10935 (N_10935,N_5490,N_6116);
nor U10936 (N_10936,N_8751,N_8135);
and U10937 (N_10937,N_9960,N_9728);
nor U10938 (N_10938,N_8869,N_6064);
and U10939 (N_10939,N_5668,N_7106);
and U10940 (N_10940,N_9819,N_9605);
nand U10941 (N_10941,N_7444,N_9454);
nand U10942 (N_10942,N_5012,N_6357);
or U10943 (N_10943,N_9857,N_6830);
and U10944 (N_10944,N_9325,N_5517);
nor U10945 (N_10945,N_5307,N_6186);
or U10946 (N_10946,N_9302,N_9305);
xor U10947 (N_10947,N_7051,N_9814);
nand U10948 (N_10948,N_5542,N_7011);
or U10949 (N_10949,N_8704,N_5187);
nor U10950 (N_10950,N_9621,N_9432);
nand U10951 (N_10951,N_9718,N_6579);
nand U10952 (N_10952,N_5523,N_7598);
nor U10953 (N_10953,N_8562,N_5591);
nor U10954 (N_10954,N_8765,N_6109);
nand U10955 (N_10955,N_5218,N_9447);
nand U10956 (N_10956,N_7171,N_5828);
and U10957 (N_10957,N_7852,N_8143);
and U10958 (N_10958,N_7592,N_7422);
or U10959 (N_10959,N_5232,N_7159);
or U10960 (N_10960,N_6637,N_7747);
and U10961 (N_10961,N_9196,N_6046);
or U10962 (N_10962,N_6593,N_6514);
and U10963 (N_10963,N_7496,N_9307);
or U10964 (N_10964,N_8012,N_9856);
or U10965 (N_10965,N_5610,N_6303);
nor U10966 (N_10966,N_8298,N_9616);
nand U10967 (N_10967,N_6412,N_6022);
nand U10968 (N_10968,N_5223,N_9582);
nand U10969 (N_10969,N_5711,N_9377);
or U10970 (N_10970,N_6075,N_5410);
nand U10971 (N_10971,N_9933,N_5039);
nand U10972 (N_10972,N_6985,N_5821);
nand U10973 (N_10973,N_8756,N_8426);
nor U10974 (N_10974,N_6429,N_7686);
xor U10975 (N_10975,N_9889,N_6786);
nor U10976 (N_10976,N_7532,N_8249);
or U10977 (N_10977,N_7740,N_7279);
xor U10978 (N_10978,N_8749,N_8281);
nand U10979 (N_10979,N_6382,N_5428);
and U10980 (N_10980,N_7853,N_9069);
nand U10981 (N_10981,N_7585,N_7089);
and U10982 (N_10982,N_5132,N_8038);
and U10983 (N_10983,N_5185,N_9387);
nand U10984 (N_10984,N_6871,N_7309);
nand U10985 (N_10985,N_6865,N_5087);
or U10986 (N_10986,N_6339,N_9471);
or U10987 (N_10987,N_8957,N_7281);
nor U10988 (N_10988,N_9533,N_8106);
nor U10989 (N_10989,N_7280,N_8561);
nor U10990 (N_10990,N_9972,N_8105);
nor U10991 (N_10991,N_8050,N_8046);
and U10992 (N_10992,N_5872,N_7947);
nor U10993 (N_10993,N_7882,N_5304);
nand U10994 (N_10994,N_8075,N_7063);
and U10995 (N_10995,N_9539,N_6713);
and U10996 (N_10996,N_8696,N_6964);
nor U10997 (N_10997,N_6193,N_8080);
nand U10998 (N_10998,N_6864,N_7545);
or U10999 (N_10999,N_5741,N_9003);
nor U11000 (N_11000,N_9485,N_9445);
nand U11001 (N_11001,N_9790,N_7620);
nand U11002 (N_11002,N_5806,N_5759);
nor U11003 (N_11003,N_6194,N_7472);
and U11004 (N_11004,N_7524,N_8582);
or U11005 (N_11005,N_5372,N_9690);
nor U11006 (N_11006,N_5873,N_7021);
xnor U11007 (N_11007,N_7110,N_7792);
and U11008 (N_11008,N_5599,N_8715);
or U11009 (N_11009,N_9402,N_5945);
or U11010 (N_11010,N_6398,N_9810);
nor U11011 (N_11011,N_7192,N_8030);
and U11012 (N_11012,N_8920,N_7360);
or U11013 (N_11013,N_7832,N_6102);
nor U11014 (N_11014,N_8848,N_8598);
nand U11015 (N_11015,N_6605,N_8522);
nand U11016 (N_11016,N_9878,N_7298);
and U11017 (N_11017,N_9607,N_6053);
or U11018 (N_11018,N_6112,N_5095);
xnor U11019 (N_11019,N_9132,N_5976);
or U11020 (N_11020,N_9417,N_6421);
nand U11021 (N_11021,N_8329,N_9797);
and U11022 (N_11022,N_9399,N_8467);
nand U11023 (N_11023,N_9811,N_7643);
nor U11024 (N_11024,N_5003,N_5446);
and U11025 (N_11025,N_9788,N_8227);
xnor U11026 (N_11026,N_5396,N_8130);
nor U11027 (N_11027,N_7376,N_6467);
or U11028 (N_11028,N_6249,N_8615);
nand U11029 (N_11029,N_8055,N_9528);
and U11030 (N_11030,N_7953,N_6383);
nor U11031 (N_11031,N_9389,N_6988);
nand U11032 (N_11032,N_6031,N_7676);
and U11033 (N_11033,N_5499,N_5451);
or U11034 (N_11034,N_8319,N_8583);
or U11035 (N_11035,N_7836,N_6162);
and U11036 (N_11036,N_6427,N_8051);
nor U11037 (N_11037,N_7406,N_8421);
nor U11038 (N_11038,N_6414,N_7080);
nor U11039 (N_11039,N_6924,N_7315);
nor U11040 (N_11040,N_5106,N_5217);
nor U11041 (N_11041,N_6241,N_6741);
and U11042 (N_11042,N_6923,N_7573);
or U11043 (N_11043,N_5585,N_9240);
or U11044 (N_11044,N_9880,N_8607);
nor U11045 (N_11045,N_5498,N_9848);
nor U11046 (N_11046,N_6245,N_8146);
or U11047 (N_11047,N_9015,N_6170);
or U11048 (N_11048,N_5055,N_8910);
nand U11049 (N_11049,N_5044,N_9119);
nor U11050 (N_11050,N_7964,N_9047);
nand U11051 (N_11051,N_5455,N_9675);
or U11052 (N_11052,N_5500,N_8405);
nand U11053 (N_11053,N_7719,N_6698);
and U11054 (N_11054,N_5404,N_6318);
nand U11055 (N_11055,N_8864,N_8788);
or U11056 (N_11056,N_6163,N_6042);
nor U11057 (N_11057,N_5048,N_7234);
and U11058 (N_11058,N_5337,N_5768);
or U11059 (N_11059,N_5157,N_5555);
or U11060 (N_11060,N_7003,N_5262);
nor U11061 (N_11061,N_5833,N_9864);
nand U11062 (N_11062,N_9491,N_8840);
nor U11063 (N_11063,N_8597,N_7868);
nand U11064 (N_11064,N_6018,N_5874);
nand U11065 (N_11065,N_7060,N_7124);
and U11066 (N_11066,N_9516,N_8021);
nor U11067 (N_11067,N_7833,N_7828);
nand U11068 (N_11068,N_5926,N_6084);
and U11069 (N_11069,N_7644,N_5623);
and U11070 (N_11070,N_7897,N_9687);
nor U11071 (N_11071,N_6930,N_9634);
nor U11072 (N_11072,N_6159,N_5138);
nand U11073 (N_11073,N_6267,N_7291);
xnor U11074 (N_11074,N_6774,N_6079);
nand U11075 (N_11075,N_9523,N_5144);
nor U11076 (N_11076,N_9543,N_5993);
or U11077 (N_11077,N_5637,N_5473);
nand U11078 (N_11078,N_5780,N_7286);
nor U11079 (N_11079,N_6734,N_7184);
or U11080 (N_11080,N_8720,N_7014);
nand U11081 (N_11081,N_5680,N_7239);
nand U11082 (N_11082,N_8953,N_8908);
or U11083 (N_11083,N_8955,N_7129);
and U11084 (N_11084,N_6392,N_6765);
nand U11085 (N_11085,N_9538,N_8407);
xnor U11086 (N_11086,N_9656,N_7876);
nor U11087 (N_11087,N_8762,N_8091);
and U11088 (N_11088,N_8587,N_5090);
nor U11089 (N_11089,N_9007,N_6931);
nand U11090 (N_11090,N_5909,N_6809);
nand U11091 (N_11091,N_8571,N_9610);
and U11092 (N_11092,N_8347,N_6216);
nor U11093 (N_11093,N_8242,N_5665);
or U11094 (N_11094,N_7251,N_7372);
xor U11095 (N_11095,N_9073,N_6911);
and U11096 (N_11096,N_7504,N_6601);
or U11097 (N_11097,N_8199,N_6857);
and U11098 (N_11098,N_7167,N_9739);
and U11099 (N_11099,N_5320,N_8262);
xor U11100 (N_11100,N_7781,N_5291);
and U11101 (N_11101,N_6693,N_9057);
or U11102 (N_11102,N_9295,N_6554);
nand U11103 (N_11103,N_7923,N_7024);
nor U11104 (N_11104,N_8590,N_9044);
nor U11105 (N_11105,N_7528,N_6954);
nand U11106 (N_11106,N_6281,N_7093);
or U11107 (N_11107,N_9664,N_5234);
nor U11108 (N_11108,N_7884,N_7565);
xnor U11109 (N_11109,N_8072,N_6961);
and U11110 (N_11110,N_5114,N_5696);
xor U11111 (N_11111,N_7556,N_8530);
and U11112 (N_11112,N_5663,N_6396);
nor U11113 (N_11113,N_9829,N_5965);
nor U11114 (N_11114,N_9468,N_5342);
or U11115 (N_11115,N_5408,N_7677);
nor U11116 (N_11116,N_7654,N_8022);
and U11117 (N_11117,N_7219,N_6814);
or U11118 (N_11118,N_6462,N_5385);
or U11119 (N_11119,N_9493,N_8264);
nand U11120 (N_11120,N_6478,N_9320);
xor U11121 (N_11121,N_7348,N_5070);
and U11122 (N_11122,N_8671,N_6548);
or U11123 (N_11123,N_7136,N_9536);
nand U11124 (N_11124,N_5433,N_6399);
nor U11125 (N_11125,N_9144,N_7112);
and U11126 (N_11126,N_7484,N_9740);
or U11127 (N_11127,N_6142,N_9892);
nor U11128 (N_11128,N_8219,N_9331);
or U11129 (N_11129,N_8274,N_5452);
nor U11130 (N_11130,N_6235,N_8292);
and U11131 (N_11131,N_6550,N_7141);
nor U11132 (N_11132,N_6259,N_8684);
and U11133 (N_11133,N_6285,N_5228);
xor U11134 (N_11134,N_7514,N_6255);
or U11135 (N_11135,N_5647,N_9489);
nor U11136 (N_11136,N_5762,N_5788);
nor U11137 (N_11137,N_8599,N_8768);
xor U11138 (N_11138,N_7142,N_5155);
and U11139 (N_11139,N_8480,N_9452);
nor U11140 (N_11140,N_7317,N_9821);
xor U11141 (N_11141,N_7566,N_7074);
or U11142 (N_11142,N_6130,N_5803);
or U11143 (N_11143,N_7581,N_7102);
and U11144 (N_11144,N_9945,N_7451);
nand U11145 (N_11145,N_5238,N_6784);
nand U11146 (N_11146,N_5799,N_7401);
and U11147 (N_11147,N_5245,N_7359);
nor U11148 (N_11148,N_6395,N_5497);
or U11149 (N_11149,N_5319,N_9254);
nor U11150 (N_11150,N_8153,N_5288);
nor U11151 (N_11151,N_7671,N_8351);
and U11152 (N_11152,N_6282,N_7697);
and U11153 (N_11153,N_7636,N_5292);
nand U11154 (N_11154,N_5413,N_6517);
and U11155 (N_11155,N_5176,N_9658);
nor U11156 (N_11156,N_6065,N_9488);
xnor U11157 (N_11157,N_9743,N_9178);
or U11158 (N_11158,N_6477,N_9751);
and U11159 (N_11159,N_7827,N_7271);
and U11160 (N_11160,N_6609,N_8416);
nand U11161 (N_11161,N_7231,N_9618);
or U11162 (N_11162,N_9086,N_8248);
nand U11163 (N_11163,N_6976,N_7235);
nand U11164 (N_11164,N_7132,N_9659);
nor U11165 (N_11165,N_6137,N_7170);
and U11166 (N_11166,N_6107,N_6613);
or U11167 (N_11167,N_7812,N_6328);
or U11168 (N_11168,N_7407,N_5691);
nor U11169 (N_11169,N_6206,N_5682);
nor U11170 (N_11170,N_5520,N_7335);
or U11171 (N_11171,N_6633,N_5646);
nor U11172 (N_11172,N_7874,N_6345);
xor U11173 (N_11173,N_6974,N_9910);
and U11174 (N_11174,N_7548,N_6021);
nand U11175 (N_11175,N_5174,N_7303);
nor U11176 (N_11176,N_9590,N_9309);
nand U11177 (N_11177,N_8315,N_5688);
and U11178 (N_11178,N_9091,N_5934);
nor U11179 (N_11179,N_9499,N_6789);
nor U11180 (N_11180,N_5266,N_7072);
nor U11181 (N_11181,N_8018,N_8457);
and U11182 (N_11182,N_6329,N_7276);
nand U11183 (N_11183,N_8330,N_7481);
nor U11184 (N_11184,N_5659,N_8645);
and U11185 (N_11185,N_5614,N_6822);
nand U11186 (N_11186,N_6272,N_5296);
nand U11187 (N_11187,N_5939,N_8695);
nor U11188 (N_11188,N_5782,N_6599);
xnor U11189 (N_11189,N_7647,N_7539);
nor U11190 (N_11190,N_7956,N_5279);
nand U11191 (N_11191,N_9077,N_7610);
or U11192 (N_11192,N_5409,N_7632);
nor U11193 (N_11193,N_7737,N_6945);
nand U11194 (N_11194,N_7490,N_9363);
or U11195 (N_11195,N_8592,N_8563);
or U11196 (N_11196,N_7301,N_8981);
or U11197 (N_11197,N_9505,N_5501);
or U11198 (N_11198,N_8962,N_5334);
nand U11199 (N_11199,N_9291,N_5920);
nor U11200 (N_11200,N_6417,N_5034);
nor U11201 (N_11201,N_9879,N_7367);
nor U11202 (N_11202,N_6505,N_6240);
nand U11203 (N_11203,N_9774,N_7026);
nand U11204 (N_11204,N_7819,N_6292);
or U11205 (N_11205,N_8037,N_6190);
nand U11206 (N_11206,N_5960,N_7971);
xnor U11207 (N_11207,N_9264,N_8617);
nand U11208 (N_11208,N_7658,N_5083);
nor U11209 (N_11209,N_8649,N_6168);
nor U11210 (N_11210,N_6926,N_8341);
or U11211 (N_11211,N_5276,N_7551);
xnor U11212 (N_11212,N_5142,N_8855);
and U11213 (N_11213,N_8122,N_6975);
nor U11214 (N_11214,N_5543,N_7462);
or U11215 (N_11215,N_8476,N_8891);
xor U11216 (N_11216,N_5042,N_8406);
nor U11217 (N_11217,N_7904,N_5801);
nand U11218 (N_11218,N_6250,N_5402);
nand U11219 (N_11219,N_9636,N_8847);
nor U11220 (N_11220,N_5084,N_7863);
and U11221 (N_11221,N_5761,N_6829);
nor U11222 (N_11222,N_6781,N_8548);
and U11223 (N_11223,N_7892,N_5970);
xor U11224 (N_11224,N_8283,N_6473);
or U11225 (N_11225,N_6408,N_8710);
and U11226 (N_11226,N_8844,N_5306);
or U11227 (N_11227,N_7449,N_6149);
nand U11228 (N_11228,N_7840,N_9893);
or U11229 (N_11229,N_7152,N_9286);
nand U11230 (N_11230,N_8189,N_9147);
or U11231 (N_11231,N_7978,N_5265);
nand U11232 (N_11232,N_7659,N_6832);
nor U11233 (N_11233,N_5879,N_7860);
xnor U11234 (N_11234,N_9969,N_6394);
and U11235 (N_11235,N_7522,N_9213);
nand U11236 (N_11236,N_7704,N_7249);
xnor U11237 (N_11237,N_7858,N_9186);
or U11238 (N_11238,N_6955,N_7248);
and U11239 (N_11239,N_9154,N_9342);
or U11240 (N_11240,N_9763,N_5968);
xnor U11241 (N_11241,N_7165,N_9172);
or U11242 (N_11242,N_8381,N_6375);
nor U11243 (N_11243,N_9547,N_7789);
or U11244 (N_11244,N_5529,N_8221);
xnor U11245 (N_11245,N_6251,N_6263);
nand U11246 (N_11246,N_8294,N_9815);
or U11247 (N_11247,N_9344,N_6232);
or U11248 (N_11248,N_8783,N_7160);
nor U11249 (N_11249,N_5431,N_6793);
nand U11250 (N_11250,N_5524,N_7306);
and U11251 (N_11251,N_9391,N_7431);
nand U11252 (N_11252,N_5724,N_8095);
nor U11253 (N_11253,N_8689,N_5025);
nand U11254 (N_11254,N_6845,N_5998);
nor U11255 (N_11255,N_5671,N_5167);
or U11256 (N_11256,N_5483,N_5654);
and U11257 (N_11257,N_8108,N_8609);
and U11258 (N_11258,N_8326,N_7499);
nand U11259 (N_11259,N_9280,N_8713);
or U11260 (N_11260,N_6518,N_7870);
nand U11261 (N_11261,N_9629,N_8461);
and U11262 (N_11262,N_7027,N_9028);
and U11263 (N_11263,N_5871,N_7975);
nor U11264 (N_11264,N_9990,N_7588);
or U11265 (N_11265,N_8195,N_6757);
xnor U11266 (N_11266,N_9934,N_9164);
and U11267 (N_11267,N_9011,N_8100);
nor U11268 (N_11268,N_9185,N_7510);
or U11269 (N_11269,N_5942,N_9548);
nand U11270 (N_11270,N_5731,N_6089);
or U11271 (N_11271,N_6540,N_7635);
nor U11272 (N_11272,N_6526,N_9724);
nor U11273 (N_11273,N_7752,N_5860);
or U11274 (N_11274,N_7701,N_5916);
or U11275 (N_11275,N_5154,N_6764);
and U11276 (N_11276,N_5568,N_9084);
nand U11277 (N_11277,N_6686,N_6576);
and U11278 (N_11278,N_5378,N_7521);
and U11279 (N_11279,N_8271,N_9863);
nand U11280 (N_11280,N_5667,N_8787);
nor U11281 (N_11281,N_6790,N_7786);
nand U11282 (N_11282,N_9233,N_8353);
or U11283 (N_11283,N_8913,N_8746);
xor U11284 (N_11284,N_5212,N_6901);
and U11285 (N_11285,N_8335,N_9257);
nor U11286 (N_11286,N_9014,N_7416);
or U11287 (N_11287,N_7212,N_8286);
xor U11288 (N_11288,N_6266,N_6881);
nor U11289 (N_11289,N_7158,N_9669);
nor U11290 (N_11290,N_7161,N_6773);
nor U11291 (N_11291,N_5124,N_9080);
nor U11292 (N_11292,N_5504,N_8723);
or U11293 (N_11293,N_7890,N_6650);
and U11294 (N_11294,N_9165,N_8724);
nand U11295 (N_11295,N_5193,N_7850);
or U11296 (N_11296,N_6653,N_6979);
nand U11297 (N_11297,N_6778,N_7637);
nor U11298 (N_11298,N_6813,N_6234);
nand U11299 (N_11299,N_5527,N_7029);
and U11300 (N_11300,N_5726,N_5719);
and U11301 (N_11301,N_9021,N_7966);
or U11302 (N_11302,N_9092,N_9358);
nor U11303 (N_11303,N_5904,N_7793);
or U11304 (N_11304,N_8228,N_7294);
nor U11305 (N_11305,N_7287,N_9741);
nand U11306 (N_11306,N_9250,N_9602);
or U11307 (N_11307,N_7835,N_5536);
nor U11308 (N_11308,N_7450,N_9958);
or U11309 (N_11309,N_5650,N_9118);
nand U11310 (N_11310,N_6499,N_5666);
nand U11311 (N_11311,N_5607,N_9449);
or U11312 (N_11312,N_7682,N_6164);
xnor U11313 (N_11313,N_6751,N_5729);
or U11314 (N_11314,N_8393,N_6008);
nor U11315 (N_11315,N_6510,N_8451);
and U11316 (N_11316,N_8025,N_7769);
nand U11317 (N_11317,N_9674,N_8418);
nor U11318 (N_11318,N_7392,N_8200);
or U11319 (N_11319,N_5085,N_7615);
nand U11320 (N_11320,N_7498,N_8352);
or U11321 (N_11321,N_5440,N_7994);
or U11322 (N_11322,N_6420,N_6808);
nor U11323 (N_11323,N_8938,N_6199);
and U11324 (N_11324,N_9010,N_5927);
and U11325 (N_11325,N_9373,N_8223);
and U11326 (N_11326,N_5603,N_9459);
or U11327 (N_11327,N_8287,N_5289);
nand U11328 (N_11328,N_5955,N_9765);
or U11329 (N_11329,N_6968,N_5158);
or U11330 (N_11330,N_5617,N_8819);
or U11331 (N_11331,N_8532,N_7223);
nand U11332 (N_11332,N_9053,N_7563);
nor U11333 (N_11333,N_7355,N_5756);
and U11334 (N_11334,N_9961,N_6639);
or U11335 (N_11335,N_6221,N_6898);
nand U11336 (N_11336,N_8691,N_7371);
nand U11337 (N_11337,N_7662,N_6996);
nand U11338 (N_11338,N_5023,N_6804);
nor U11339 (N_11339,N_8774,N_9438);
nand U11340 (N_11340,N_5143,N_5777);
and U11341 (N_11341,N_5882,N_7688);
nand U11342 (N_11342,N_7384,N_5579);
nand U11343 (N_11343,N_6574,N_5092);
nand U11344 (N_11344,N_6476,N_6331);
nor U11345 (N_11345,N_6960,N_5345);
nor U11346 (N_11346,N_5807,N_6482);
nand U11347 (N_11347,N_5121,N_8118);
nor U11348 (N_11348,N_8677,N_9766);
nor U11349 (N_11349,N_8497,N_8594);
nor U11350 (N_11350,N_9251,N_9508);
nor U11351 (N_11351,N_9101,N_7067);
or U11352 (N_11352,N_7333,N_9125);
xnor U11353 (N_11353,N_6799,N_5903);
nor U11354 (N_11354,N_5808,N_9775);
and U11355 (N_11355,N_5131,N_5445);
nand U11356 (N_11356,N_9483,N_6995);
nor U11357 (N_11357,N_7016,N_8553);
nand U11358 (N_11358,N_5732,N_9729);
and U11359 (N_11359,N_5940,N_6182);
nor U11360 (N_11360,N_9156,N_8389);
and U11361 (N_11361,N_8925,N_7386);
nor U11362 (N_11362,N_5763,N_7675);
and U11363 (N_11363,N_9206,N_7933);
nor U11364 (N_11364,N_5463,N_7918);
xnor U11365 (N_11365,N_7738,N_6688);
nor U11366 (N_11366,N_5147,N_8712);
nor U11367 (N_11367,N_6516,N_5834);
nand U11368 (N_11368,N_5229,N_6524);
and U11369 (N_11369,N_7070,N_7705);
nand U11370 (N_11370,N_6448,N_9433);
and U11371 (N_11371,N_7794,N_6000);
xnor U11372 (N_11372,N_9776,N_9374);
xnor U11373 (N_11373,N_9952,N_5054);
nand U11374 (N_11374,N_5730,N_6020);
or U11375 (N_11375,N_8944,N_8409);
nand U11376 (N_11376,N_9643,N_5195);
and U11377 (N_11377,N_9511,N_5361);
xnor U11378 (N_11378,N_9400,N_7700);
or U11379 (N_11379,N_9089,N_7508);
nand U11380 (N_11380,N_5676,N_5327);
or U11381 (N_11381,N_6225,N_7330);
nand U11382 (N_11382,N_9779,N_6158);
and U11383 (N_11383,N_7006,N_5139);
or U11384 (N_11384,N_9275,N_6607);
nand U11385 (N_11385,N_7613,N_6538);
or U11386 (N_11386,N_7188,N_7388);
and U11387 (N_11387,N_8060,N_9830);
nor U11388 (N_11388,N_6269,N_6990);
xor U11389 (N_11389,N_5454,N_7783);
xor U11390 (N_11390,N_6521,N_5935);
and U11391 (N_11391,N_5561,N_5710);
and U11392 (N_11392,N_7754,N_6754);
nor U11393 (N_11393,N_8579,N_8661);
xnor U11394 (N_11394,N_7482,N_9845);
nand U11395 (N_11395,N_5588,N_8506);
nand U11396 (N_11396,N_8574,N_8741);
nand U11397 (N_11397,N_9093,N_7561);
and U11398 (N_11398,N_9576,N_8112);
xor U11399 (N_11399,N_8680,N_7292);
nand U11400 (N_11400,N_7261,N_6821);
and U11401 (N_11401,N_5736,N_8979);
and U11402 (N_11402,N_6155,N_8974);
nand U11403 (N_11403,N_5753,N_5182);
or U11404 (N_11404,N_7186,N_7594);
and U11405 (N_11405,N_9710,N_8215);
nor U11406 (N_11406,N_5261,N_9561);
nand U11407 (N_11407,N_6951,N_7568);
xor U11408 (N_11408,N_7713,N_7259);
nand U11409 (N_11409,N_6085,N_7125);
or U11410 (N_11410,N_8447,N_5179);
or U11411 (N_11411,N_7216,N_5401);
nor U11412 (N_11412,N_8311,N_8996);
nand U11413 (N_11413,N_8656,N_6391);
xor U11414 (N_11414,N_9440,N_9238);
or U11415 (N_11415,N_5626,N_9376);
nand U11416 (N_11416,N_9062,N_8804);
nor U11417 (N_11417,N_5219,N_9986);
and U11418 (N_11418,N_9651,N_5031);
or U11419 (N_11419,N_6470,N_9851);
nor U11420 (N_11420,N_9780,N_6783);
xor U11421 (N_11421,N_8761,N_7427);
or U11422 (N_11422,N_8321,N_7369);
or U11423 (N_11423,N_9861,N_8797);
or U11424 (N_11424,N_7269,N_9841);
and U11425 (N_11425,N_8415,N_8297);
or U11426 (N_11426,N_7195,N_7579);
nand U11427 (N_11427,N_7381,N_8028);
and U11428 (N_11428,N_8608,N_5033);
or U11429 (N_11429,N_7300,N_8702);
or U11430 (N_11430,N_7716,N_6185);
and U11431 (N_11431,N_9051,N_9143);
and U11432 (N_11432,N_7290,N_8867);
nand U11433 (N_11433,N_7007,N_9795);
or U11434 (N_11434,N_7759,N_8441);
and U11435 (N_11435,N_7722,N_8474);
nand U11436 (N_11436,N_8542,N_6313);
nand U11437 (N_11437,N_7116,N_6146);
nor U11438 (N_11438,N_8633,N_6397);
nor U11439 (N_11439,N_9183,N_9939);
or U11440 (N_11440,N_8576,N_7433);
and U11441 (N_11441,N_7574,N_5080);
nand U11442 (N_11442,N_5503,N_5119);
or U11443 (N_11443,N_5771,N_6479);
or U11444 (N_11444,N_8325,N_5470);
and U11445 (N_11445,N_5496,N_9217);
and U11446 (N_11446,N_7349,N_9212);
nor U11447 (N_11447,N_8435,N_5277);
nor U11448 (N_11448,N_7617,N_9859);
nor U11449 (N_11449,N_7256,N_5827);
xnor U11450 (N_11450,N_6086,N_6454);
or U11451 (N_11451,N_9242,N_9456);
or U11452 (N_11452,N_6900,N_7791);
nor U11453 (N_11453,N_8790,N_9061);
nor U11454 (N_11454,N_7157,N_6330);
and U11455 (N_11455,N_7440,N_8886);
and U11456 (N_11456,N_8556,N_8948);
nand U11457 (N_11457,N_5469,N_8420);
and U11458 (N_11458,N_7457,N_6256);
nor U11459 (N_11459,N_9875,N_5222);
nor U11460 (N_11460,N_9214,N_6942);
xor U11461 (N_11461,N_8240,N_8376);
xor U11462 (N_11462,N_7107,N_5141);
nand U11463 (N_11463,N_8832,N_9317);
nand U11464 (N_11464,N_9767,N_7879);
nor U11465 (N_11465,N_8951,N_6495);
or U11466 (N_11466,N_8364,N_7891);
or U11467 (N_11467,N_6761,N_7801);
nor U11468 (N_11468,N_6520,N_7537);
nor U11469 (N_11469,N_8296,N_9113);
or U11470 (N_11470,N_6172,N_5290);
or U11471 (N_11471,N_5305,N_6743);
nor U11472 (N_11472,N_9401,N_9208);
nand U11473 (N_11473,N_5984,N_6028);
or U11474 (N_11474,N_6848,N_8942);
and U11475 (N_11475,N_8310,N_7109);
xor U11476 (N_11476,N_7619,N_9620);
nand U11477 (N_11477,N_9025,N_7130);
nor U11478 (N_11478,N_5488,N_5925);
and U11479 (N_11479,N_8818,N_8423);
nand U11480 (N_11480,N_5294,N_8098);
xor U11481 (N_11481,N_6432,N_9262);
or U11482 (N_11482,N_8466,N_5118);
nand U11483 (N_11483,N_9955,N_5704);
or U11484 (N_11484,N_9334,N_5251);
and U11485 (N_11485,N_5269,N_6442);
xor U11486 (N_11486,N_7814,N_9823);
and U11487 (N_11487,N_7679,N_9005);
and U11488 (N_11488,N_6299,N_5900);
and U11489 (N_11489,N_5471,N_5958);
and U11490 (N_11490,N_9136,N_5783);
nor U11491 (N_11491,N_5325,N_6523);
nand U11492 (N_11492,N_8703,N_5991);
nand U11493 (N_11493,N_5744,N_6922);
or U11494 (N_11494,N_7648,N_6839);
nand U11495 (N_11495,N_6485,N_9150);
and U11496 (N_11496,N_7245,N_9255);
nor U11497 (N_11497,N_7962,N_8450);
or U11498 (N_11498,N_6886,N_5686);
nor U11499 (N_11499,N_8570,N_8907);
or U11500 (N_11500,N_9106,N_6903);
nand U11501 (N_11501,N_8524,N_7246);
xnor U11502 (N_11502,N_5377,N_9037);
or U11503 (N_11503,N_9717,N_9865);
and U11504 (N_11504,N_6305,N_7596);
nand U11505 (N_11505,N_5658,N_5375);
and U11506 (N_11506,N_8823,N_8679);
nor U11507 (N_11507,N_5649,N_8339);
xnor U11508 (N_11508,N_6274,N_6009);
or U11509 (N_11509,N_6577,N_5889);
nor U11510 (N_11510,N_9840,N_8412);
or U11511 (N_11511,N_9370,N_8449);
or U11512 (N_11512,N_6326,N_9570);
or U11513 (N_11513,N_7477,N_6244);
nor U11514 (N_11514,N_7385,N_9678);
and U11515 (N_11515,N_5231,N_5509);
nor U11516 (N_11516,N_6446,N_7912);
nor U11517 (N_11517,N_6592,N_8029);
and U11518 (N_11518,N_8547,N_9244);
nor U11519 (N_11519,N_7657,N_5804);
and U11520 (N_11520,N_7806,N_7091);
or U11521 (N_11521,N_8145,N_5094);
nand U11522 (N_11522,N_8540,N_7040);
nor U11523 (N_11523,N_9482,N_6726);
and U11524 (N_11524,N_7748,N_8293);
nor U11525 (N_11525,N_7324,N_8729);
nand U11526 (N_11526,N_5797,N_7429);
or U11527 (N_11527,N_9808,N_8735);
nor U11528 (N_11528,N_5737,N_5249);
nand U11529 (N_11529,N_9686,N_6838);
or U11530 (N_11530,N_5308,N_6099);
or U11531 (N_11531,N_6344,N_5979);
and U11532 (N_11532,N_6689,N_9731);
and U11533 (N_11533,N_5786,N_7305);
and U11534 (N_11534,N_8152,N_9109);
nor U11535 (N_11535,N_8301,N_8013);
nor U11536 (N_11536,N_9256,N_6569);
or U11537 (N_11537,N_5478,N_8805);
nor U11538 (N_11538,N_8673,N_9696);
or U11539 (N_11539,N_9357,N_5208);
or U11540 (N_11540,N_9551,N_9817);
and U11541 (N_11541,N_8687,N_7721);
nor U11542 (N_11542,N_7438,N_7377);
nand U11543 (N_11543,N_8967,N_9450);
nand U11544 (N_11544,N_7788,N_7323);
and U11545 (N_11545,N_9564,N_9925);
nand U11546 (N_11546,N_6748,N_7607);
nor U11547 (N_11547,N_9347,N_8757);
and U11548 (N_11548,N_6936,N_6530);
nand U11549 (N_11549,N_5175,N_5748);
nor U11550 (N_11550,N_9980,N_6056);
and U11551 (N_11551,N_8104,N_6012);
or U11552 (N_11552,N_7896,N_6368);
and U11553 (N_11553,N_6811,N_8194);
or U11554 (N_11554,N_5064,N_7084);
or U11555 (N_11555,N_9513,N_8452);
or U11556 (N_11556,N_6989,N_8872);
xnor U11557 (N_11557,N_8747,N_6617);
and U11558 (N_11558,N_7830,N_6697);
nand U11559 (N_11559,N_6723,N_5701);
nand U11560 (N_11560,N_7888,N_9606);
or U11561 (N_11561,N_5713,N_7698);
xnor U11562 (N_11562,N_9685,N_5233);
nor U11563 (N_11563,N_6415,N_5271);
or U11564 (N_11564,N_7753,N_9484);
or U11565 (N_11565,N_7729,N_6715);
nand U11566 (N_11566,N_9580,N_7667);
nand U11567 (N_11567,N_7250,N_7442);
nor U11568 (N_11568,N_6621,N_9105);
and U11569 (N_11569,N_5822,N_9343);
nand U11570 (N_11570,N_7506,N_6280);
and U11571 (N_11571,N_5267,N_6278);
or U11572 (N_11572,N_6487,N_5343);
and U11573 (N_11573,N_6469,N_8890);
nor U11574 (N_11574,N_5021,N_9886);
or U11575 (N_11575,N_8132,N_8933);
or U11576 (N_11576,N_5323,N_6863);
or U11577 (N_11577,N_9624,N_5395);
nor U11578 (N_11578,N_5397,N_5988);
or U11579 (N_11579,N_6925,N_5978);
xnor U11580 (N_11580,N_8016,N_5177);
or U11581 (N_11581,N_8849,N_9733);
and U11582 (N_11582,N_9627,N_7458);
or U11583 (N_11583,N_8549,N_8373);
nor U11584 (N_11584,N_5760,N_6876);
nor U11585 (N_11585,N_7618,N_7763);
and U11586 (N_11586,N_9524,N_5723);
and U11587 (N_11587,N_5938,N_9017);
or U11588 (N_11588,N_9951,N_8810);
nand U11589 (N_11589,N_8269,N_9405);
and U11590 (N_11590,N_6874,N_8758);
or U11591 (N_11591,N_6559,N_6093);
or U11592 (N_11592,N_8019,N_8641);
xnor U11593 (N_11593,N_9540,N_9801);
and U11594 (N_11594,N_6836,N_8578);
and U11595 (N_11595,N_5416,N_6800);
xor U11596 (N_11596,N_7182,N_9480);
nand U11597 (N_11597,N_9337,N_8477);
nand U11598 (N_11598,N_9312,N_6070);
nor U11599 (N_11599,N_8784,N_5906);
nor U11600 (N_11600,N_7059,N_5341);
nand U11601 (N_11601,N_8149,N_8408);
or U11602 (N_11602,N_6497,N_8640);
or U11603 (N_11603,N_5194,N_6161);
nand U11604 (N_11604,N_5605,N_8965);
nand U11605 (N_11605,N_9682,N_5784);
or U11606 (N_11606,N_8356,N_8097);
nand U11607 (N_11607,N_8544,N_5644);
nor U11608 (N_11608,N_6750,N_9745);
or U11609 (N_11609,N_8902,N_7354);
nand U11610 (N_11610,N_8486,N_9063);
nand U11611 (N_11611,N_7572,N_6051);
or U11612 (N_11612,N_6366,N_6224);
or U11613 (N_11613,N_6023,N_5101);
xor U11614 (N_11614,N_9847,N_5656);
nor U11615 (N_11615,N_6815,N_6628);
nor U11616 (N_11616,N_7215,N_6586);
nor U11617 (N_11617,N_6915,N_9111);
and U11618 (N_11618,N_6071,N_5122);
nand U11619 (N_11619,N_8868,N_9600);
and U11620 (N_11620,N_5959,N_5816);
nor U11621 (N_11621,N_8516,N_5475);
xor U11622 (N_11622,N_7955,N_8945);
or U11623 (N_11623,N_7678,N_8994);
and U11624 (N_11624,N_5750,N_8591);
xor U11625 (N_11625,N_5172,N_6937);
nand U11626 (N_11626,N_6602,N_5683);
and U11627 (N_11627,N_5742,N_8184);
nand U11628 (N_11628,N_5857,N_9253);
or U11629 (N_11629,N_5681,N_5109);
nor U11630 (N_11630,N_5461,N_5116);
nor U11631 (N_11631,N_8937,N_5365);
and U11632 (N_11632,N_9416,N_5949);
nand U11633 (N_11633,N_9825,N_7818);
nor U11634 (N_11634,N_5002,N_6494);
or U11635 (N_11635,N_5110,N_9520);
nand U11636 (N_11636,N_7846,N_8300);
nor U11637 (N_11637,N_9849,N_9463);
nand U11638 (N_11638,N_6646,N_8369);
nand U11639 (N_11639,N_9215,N_5995);
nand U11640 (N_11640,N_5047,N_5869);
or U11641 (N_11641,N_9911,N_8519);
nor U11642 (N_11642,N_5202,N_9553);
nor U11643 (N_11643,N_6584,N_7131);
xnor U11644 (N_11644,N_7601,N_9279);
and U11645 (N_11645,N_6091,N_9956);
nor U11646 (N_11646,N_8916,N_8990);
and U11647 (N_11647,N_6035,N_7413);
nand U11648 (N_11648,N_5225,N_8093);
nor U11649 (N_11649,N_9192,N_7155);
or U11650 (N_11650,N_6729,N_5581);
nand U11651 (N_11651,N_8536,N_5420);
nor U11652 (N_11652,N_8589,N_8254);
nand U11653 (N_11653,N_5263,N_9365);
nor U11654 (N_11654,N_5624,N_8445);
and U11655 (N_11655,N_6237,N_6862);
or U11656 (N_11656,N_9128,N_5056);
or U11657 (N_11657,N_8665,N_6252);
or U11658 (N_11658,N_9198,N_6534);
nor U11659 (N_11659,N_7225,N_9786);
nand U11660 (N_11660,N_8625,N_8876);
nor U11661 (N_11661,N_6958,N_7135);
nand U11662 (N_11662,N_7707,N_9979);
xnor U11663 (N_11663,N_7614,N_7920);
nor U11664 (N_11664,N_5240,N_9650);
xnor U11665 (N_11665,N_7922,N_5870);
nand U11666 (N_11666,N_9333,N_8700);
nor U11667 (N_11667,N_7656,N_7018);
and U11668 (N_11668,N_7389,N_6972);
nor U11669 (N_11669,N_7505,N_7578);
or U11670 (N_11670,N_8216,N_6714);
nor U11671 (N_11671,N_5533,N_6418);
xor U11672 (N_11672,N_8384,N_9914);
and U11673 (N_11673,N_5640,N_5192);
and U11674 (N_11674,N_9822,N_8694);
and U11675 (N_11675,N_9742,N_6317);
and U11676 (N_11676,N_5687,N_6074);
or U11677 (N_11677,N_5443,N_7237);
xnor U11678 (N_11678,N_8551,N_7802);
nand U11679 (N_11679,N_8545,N_7163);
nand U11680 (N_11680,N_7867,N_7175);
xor U11681 (N_11681,N_7069,N_7010);
nor U11682 (N_11682,N_9573,N_8285);
nor U11683 (N_11683,N_5184,N_6666);
or U11684 (N_11684,N_9894,N_5235);
nand U11685 (N_11685,N_5792,N_8178);
nor U11686 (N_11686,N_6005,N_5112);
nand U11687 (N_11687,N_5738,N_7002);
and U11688 (N_11688,N_7674,N_6727);
nand U11689 (N_11689,N_8537,N_6725);
and U11690 (N_11690,N_9289,N_9625);
or U11691 (N_11691,N_5850,N_9870);
or U11692 (N_11692,N_9688,N_6119);
nand U11693 (N_11693,N_9608,N_6003);
and U11694 (N_11694,N_8811,N_6258);
nand U11695 (N_11695,N_5254,N_9273);
or U11696 (N_11696,N_6013,N_8814);
or U11697 (N_11697,N_9899,N_8678);
nand U11698 (N_11698,N_9761,N_5076);
xor U11699 (N_11699,N_6289,N_9599);
nand U11700 (N_11700,N_7154,N_8059);
or U11701 (N_11701,N_9314,N_8682);
nand U11702 (N_11702,N_8355,N_6712);
nand U11703 (N_11703,N_5405,N_9900);
nand U11704 (N_11704,N_6041,N_6802);
nand U11705 (N_11705,N_6087,N_9723);
xnor U11706 (N_11706,N_6831,N_5159);
nor U11707 (N_11707,N_9697,N_7071);
and U11708 (N_11708,N_8523,N_7342);
nor U11709 (N_11709,N_7646,N_7370);
or U11710 (N_11710,N_7081,N_6542);
nand U11711 (N_11711,N_7960,N_7925);
and U11712 (N_11712,N_9959,N_9897);
and U11713 (N_11713,N_6994,N_8165);
and U11714 (N_11714,N_5104,N_7039);
and U11715 (N_11715,N_6230,N_8820);
or U11716 (N_11716,N_5311,N_9282);
nand U11717 (N_11717,N_9381,N_5616);
or U11718 (N_11718,N_6151,N_5812);
nand U11719 (N_11719,N_9087,N_6381);
nor U11720 (N_11720,N_9559,N_7734);
and U11721 (N_11721,N_6627,N_9518);
xor U11722 (N_11722,N_7346,N_8652);
xor U11723 (N_11723,N_8560,N_6304);
and U11724 (N_11724,N_8657,N_8042);
or U11725 (N_11725,N_9397,N_6668);
nand U11726 (N_11726,N_9187,N_5851);
and U11727 (N_11727,N_5632,N_6362);
nand U11728 (N_11728,N_9067,N_8929);
nand U11729 (N_11729,N_7695,N_6888);
nand U11730 (N_11730,N_7325,N_9359);
or U11731 (N_11731,N_8268,N_7162);
or U11732 (N_11732,N_7331,N_6861);
and U11733 (N_11733,N_9161,N_8717);
nand U11734 (N_11734,N_7877,N_7383);
nor U11735 (N_11735,N_7533,N_7523);
and U11736 (N_11736,N_8572,N_9873);
nor U11737 (N_11737,N_5718,N_9679);
nor U11738 (N_11738,N_9407,N_7760);
and U11739 (N_11739,N_7777,N_8521);
nor U11740 (N_11740,N_5494,N_6129);
xnor U11741 (N_11741,N_9982,N_6247);
nand U11742 (N_11742,N_5700,N_6140);
or U11743 (N_11743,N_5264,N_8167);
nor U11744 (N_11744,N_7878,N_9159);
nand U11745 (N_11745,N_8344,N_6902);
and U11746 (N_11746,N_9392,N_7415);
and U11747 (N_11747,N_8218,N_6364);
nand U11748 (N_11748,N_9905,N_7474);
and U11749 (N_11749,N_7491,N_5952);
and U11750 (N_11750,N_8781,N_7952);
or U11751 (N_11751,N_7222,N_8332);
xnor U11752 (N_11752,N_9532,N_7622);
and U11753 (N_11753,N_8185,N_8626);
and U11754 (N_11754,N_6825,N_9046);
or U11755 (N_11755,N_8187,N_7075);
or U11756 (N_11756,N_6870,N_7126);
and U11757 (N_11757,N_5126,N_5674);
nand U11758 (N_11758,N_5539,N_8172);
nand U11759 (N_11759,N_7289,N_6679);
or U11760 (N_11760,N_5079,N_8197);
nor U11761 (N_11761,N_8812,N_5893);
or U11762 (N_11762,N_9704,N_5662);
or U11763 (N_11763,N_5298,N_8585);
nand U11764 (N_11764,N_8683,N_9953);
and U11765 (N_11765,N_6642,N_8327);
nor U11766 (N_11766,N_7053,N_8400);
and U11767 (N_11767,N_9562,N_7886);
nor U11768 (N_11768,N_7128,N_7810);
and U11769 (N_11769,N_5853,N_5115);
or U11770 (N_11770,N_5197,N_7486);
and U11771 (N_11771,N_5566,N_8546);
and U11772 (N_11772,N_5831,N_5562);
and U11773 (N_11773,N_9300,N_8471);
and U11774 (N_11774,N_6490,N_7803);
nand U11775 (N_11775,N_6541,N_9941);
nand U11776 (N_11776,N_8182,N_6139);
nand U11777 (N_11777,N_8074,N_6025);
nand U11778 (N_11778,N_5817,N_6189);
and U11779 (N_11779,N_8601,N_8785);
xor U11780 (N_11780,N_6260,N_6818);
xnor U11781 (N_11781,N_7247,N_6624);
and U11782 (N_11782,N_7166,N_7621);
and U11783 (N_11783,N_9097,N_9726);
and U11784 (N_11784,N_9928,N_5430);
or U11785 (N_11785,N_5239,N_7586);
nor U11786 (N_11786,N_6336,N_6852);
nand U11787 (N_11787,N_5097,N_5781);
nor U11788 (N_11788,N_5621,N_7798);
xnor U11789 (N_11789,N_9628,N_7140);
and U11790 (N_11790,N_6634,N_9567);
nor U11791 (N_11791,N_7750,N_7562);
nor U11792 (N_11792,N_7509,N_9396);
nor U11793 (N_11793,N_8850,N_7609);
and U11794 (N_11794,N_9284,N_9502);
xor U11795 (N_11795,N_6143,N_6024);
nor U11796 (N_11796,N_5161,N_8169);
xor U11797 (N_11797,N_5643,N_7584);
nand U11798 (N_11798,N_5751,N_7839);
nor U11799 (N_11799,N_7652,N_5609);
nand U11800 (N_11800,N_6939,N_9746);
and U11801 (N_11801,N_5442,N_9736);
or U11802 (N_11802,N_6253,N_8616);
and U11803 (N_11803,N_8514,N_9094);
nand U11804 (N_11804,N_5776,N_7088);
or U11805 (N_11805,N_9222,N_9083);
nand U11806 (N_11806,N_5513,N_7996);
or U11807 (N_11807,N_9141,N_6917);
nor U11808 (N_11808,N_8079,N_6484);
nor U11809 (N_11809,N_8898,N_7172);
or U11810 (N_11810,N_5004,N_7266);
nand U11811 (N_11811,N_6066,N_7494);
nor U11812 (N_11812,N_7824,N_6859);
and U11813 (N_11813,N_7101,N_5317);
and U11814 (N_11814,N_9976,N_7104);
nor U11815 (N_11815,N_9907,N_9223);
xnor U11816 (N_11816,N_8926,N_5029);
and U11817 (N_11817,N_8822,N_7238);
nand U11818 (N_11818,N_8429,N_7375);
nor U11819 (N_11819,N_7599,N_5190);
xor U11820 (N_11820,N_6730,N_9422);
or U11821 (N_11821,N_5268,N_6050);
xor U11822 (N_11822,N_9759,N_9844);
xnor U11823 (N_11823,N_7702,N_5066);
nand U11824 (N_11824,N_8473,N_5618);
or U11825 (N_11825,N_5270,N_7908);
or U11826 (N_11826,N_8877,N_5573);
and U11827 (N_11827,N_7773,N_6197);
nor U11828 (N_11828,N_5411,N_9056);
nor U11829 (N_11829,N_6434,N_7708);
or U11830 (N_11830,N_8487,N_9968);
or U11831 (N_11831,N_9592,N_6899);
and U11832 (N_11832,N_7518,N_6444);
nand U11833 (N_11833,N_9371,N_7495);
or U11834 (N_11834,N_9882,N_6169);
or U11835 (N_11835,N_8320,N_8258);
and U11836 (N_11836,N_5845,N_5549);
nand U11837 (N_11837,N_8203,N_9938);
or U11838 (N_11838,N_9339,N_5846);
nand U11839 (N_11839,N_9884,N_7004);
and U11840 (N_11840,N_6080,N_9437);
and U11841 (N_11841,N_6459,N_7097);
nor U11842 (N_11842,N_5280,N_9076);
nand U11843 (N_11843,N_5844,N_7541);
nor U11844 (N_11844,N_9552,N_6558);
and U11845 (N_11845,N_8062,N_9272);
nor U11846 (N_11846,N_7263,N_6708);
or U11847 (N_11847,N_8444,N_6841);
and U11848 (N_11848,N_9379,N_9757);
or U11849 (N_11849,N_7123,N_9756);
and U11850 (N_11850,N_9991,N_8442);
nand U11851 (N_11851,N_9267,N_6928);
and U11852 (N_11852,N_7898,N_6724);
nand U11853 (N_11853,N_8489,N_8043);
and U11854 (N_11854,N_6498,N_6779);
or U11855 (N_11855,N_8459,N_8827);
or U11856 (N_11856,N_9070,N_6122);
and U11857 (N_11857,N_6063,N_7023);
or U11858 (N_11858,N_9929,N_5863);
and U11859 (N_11859,N_5652,N_7919);
and U11860 (N_11860,N_6927,N_6207);
nor U11861 (N_11861,N_7468,N_9940);
nand U11862 (N_11862,N_5596,N_8431);
or U11863 (N_11863,N_5810,N_9706);
nor U11864 (N_11864,N_9546,N_5717);
xnor U11865 (N_11865,N_5758,N_5241);
xnor U11866 (N_11866,N_9526,N_6430);
xnor U11867 (N_11867,N_6452,N_7179);
and U11868 (N_11868,N_6673,N_6435);
nand U11869 (N_11869,N_7669,N_7174);
and U11870 (N_11870,N_5367,N_8479);
nand U11871 (N_11871,N_9803,N_9467);
or U11872 (N_11872,N_9707,N_7790);
and U11873 (N_11873,N_9326,N_7583);
nand U11874 (N_11874,N_5685,N_8067);
nand U11875 (N_11875,N_5321,N_8935);
nand U11876 (N_11876,N_9294,N_8817);
or U11877 (N_11877,N_8375,N_8940);
xor U11878 (N_11878,N_8004,N_8035);
and U11879 (N_11879,N_7902,N_9066);
nor U11880 (N_11880,N_6612,N_5224);
or U11881 (N_11881,N_6424,N_5578);
or U11882 (N_11882,N_8394,N_8370);
xor U11883 (N_11883,N_7344,N_8596);
nand U11884 (N_11884,N_8881,N_5415);
nand U11885 (N_11885,N_8992,N_9355);
nand U11886 (N_11886,N_9915,N_5186);
and U11887 (N_11887,N_5813,N_8637);
nor U11888 (N_11888,N_9285,N_5815);
or U11889 (N_11889,N_7085,N_5453);
and U11890 (N_11890,N_5554,N_9681);
xnor U11891 (N_11891,N_7079,N_9632);
nand U11892 (N_11892,N_9995,N_9322);
nand U11893 (N_11893,N_6323,N_6567);
nor U11894 (N_11894,N_9039,N_6208);
or U11895 (N_11895,N_7218,N_9195);
xor U11896 (N_11896,N_7887,N_5699);
nor U11897 (N_11897,N_9153,N_5348);
or U11898 (N_11898,N_6669,N_5278);
and U11899 (N_11899,N_9640,N_5049);
nand U11900 (N_11900,N_7145,N_6165);
or U11901 (N_11901,N_6866,N_5648);
and U11902 (N_11902,N_7772,N_6997);
nor U11903 (N_11903,N_7320,N_7692);
nor U11904 (N_11904,N_5309,N_9662);
and U11905 (N_11905,N_6152,N_9946);
xor U11906 (N_11906,N_5427,N_6004);
nand U11907 (N_11907,N_8502,N_8742);
or U11908 (N_11908,N_7061,N_6916);
nand U11909 (N_11909,N_7374,N_8253);
xor U11910 (N_11910,N_9227,N_7997);
or U11911 (N_11911,N_7515,N_7733);
and U11912 (N_11912,N_8053,N_6503);
and U11913 (N_11913,N_7260,N_9987);
nand U11914 (N_11914,N_8071,N_5328);
or U11915 (N_11915,N_6322,N_5248);
or U11916 (N_11916,N_7424,N_5972);
nor U11917 (N_11917,N_8348,N_5458);
or U11918 (N_11918,N_7712,N_6594);
nand U11919 (N_11919,N_7906,N_8709);
and U11920 (N_11920,N_6919,N_5120);
nand U11921 (N_11921,N_6950,N_9026);
nor U11922 (N_11922,N_8843,N_7236);
nor U11923 (N_11923,N_8036,N_5407);
nor U11924 (N_11924,N_9998,N_7519);
or U11925 (N_11925,N_7254,N_6573);
and U11926 (N_11926,N_8879,N_9853);
or U11927 (N_11927,N_6549,N_7641);
nand U11928 (N_11928,N_7767,N_6775);
xnor U11929 (N_11929,N_9583,N_9846);
nand U11930 (N_11930,N_6228,N_5145);
or U11931 (N_11931,N_8024,N_8207);
and U11932 (N_11932,N_8654,N_8932);
nor U11933 (N_11933,N_5073,N_7194);
nand U11934 (N_11934,N_7203,N_6465);
xnor U11935 (N_11935,N_5387,N_5273);
nand U11936 (N_11936,N_7380,N_8007);
or U11937 (N_11937,N_5481,N_7554);
nor U11938 (N_11938,N_6728,N_9448);
nor U11939 (N_11939,N_9095,N_6290);
xnor U11940 (N_11940,N_7577,N_7265);
and U11941 (N_11941,N_5191,N_8857);
or U11942 (N_11942,N_5875,N_7492);
or U11943 (N_11943,N_9896,N_9752);
nand U11944 (N_11944,N_8686,N_8377);
nor U11945 (N_11945,N_7092,N_7228);
and U11946 (N_11946,N_8436,N_9521);
nand U11947 (N_11947,N_7361,N_9002);
and U11948 (N_11948,N_8245,N_8543);
nand U11949 (N_11949,N_5284,N_8875);
xor U11950 (N_11950,N_5918,N_5153);
nor U11951 (N_11951,N_8163,N_9512);
nor U11952 (N_11952,N_7446,N_9557);
nand U11953 (N_11953,N_7557,N_9045);
xnor U11954 (N_11954,N_6131,N_6659);
nand U11955 (N_11955,N_6297,N_9052);
xor U11956 (N_11956,N_5487,N_7655);
nand U11957 (N_11957,N_8614,N_8873);
and U11958 (N_11958,N_5286,N_6884);
nand U11959 (N_11959,N_6178,N_9515);
nand U11960 (N_11960,N_7929,N_6016);
or U11961 (N_11961,N_8455,N_8160);
and U11962 (N_11962,N_9243,N_5722);
nor U11963 (N_11963,N_8706,N_7838);
and U11964 (N_11964,N_8733,N_5672);
nand U11965 (N_11965,N_6640,N_7595);
nor U11966 (N_11966,N_9424,N_9033);
and U11967 (N_11967,N_7981,N_6849);
nor U11968 (N_11968,N_9160,N_5932);
nor U11969 (N_11969,N_8726,N_5380);
or U11970 (N_11970,N_9478,N_8941);
xnor U11971 (N_11971,N_8432,N_5634);
xor U11972 (N_11972,N_5074,N_7866);
nor U11973 (N_11973,N_6788,N_9088);
or U11974 (N_11974,N_8333,N_5180);
nand U11975 (N_11975,N_5482,N_6794);
nand U11976 (N_11976,N_7393,N_8539);
or U11977 (N_11977,N_8866,N_9530);
nor U11978 (N_11978,N_6327,N_8045);
nor U11979 (N_11979,N_6293,N_8205);
nand U11980 (N_11980,N_6388,N_7977);
or U11981 (N_11981,N_6532,N_9984);
xor U11982 (N_11982,N_5127,N_6475);
or U11983 (N_11983,N_7396,N_8387);
or U11984 (N_11984,N_8229,N_8233);
nor U11985 (N_11985,N_7211,N_5450);
nand U11986 (N_11986,N_6742,N_6563);
nor U11987 (N_11987,N_7864,N_6782);
or U11988 (N_11988,N_6897,N_5392);
and U11989 (N_11989,N_9194,N_6912);
or U11990 (N_11990,N_7138,N_9974);
nand U11991 (N_11991,N_7316,N_9124);
or U11992 (N_11992,N_8259,N_5996);
and U11993 (N_11993,N_8144,N_7322);
and U11994 (N_11994,N_9139,N_9383);
or U11995 (N_11995,N_7687,N_6973);
or U11996 (N_11996,N_6999,N_6543);
and U11997 (N_11997,N_9085,N_9001);
nand U11998 (N_11998,N_9218,N_7880);
nor U11999 (N_11999,N_8014,N_6078);
nor U12000 (N_12000,N_9462,N_8961);
nand U12001 (N_12001,N_9833,N_9677);
nand U12002 (N_12002,N_9994,N_9112);
xnor U12003 (N_12003,N_6466,N_6060);
nor U12004 (N_12004,N_5629,N_8419);
xnor U12005 (N_12005,N_6953,N_6665);
or U12006 (N_12006,N_8801,N_5622);
nor U12007 (N_12007,N_7797,N_9207);
nand U12008 (N_12008,N_6966,N_6721);
and U12009 (N_12009,N_7915,N_6468);
nand U12010 (N_12010,N_8475,N_9525);
and U12011 (N_12011,N_6941,N_8565);
and U12012 (N_12012,N_9824,N_7940);
and U12013 (N_12013,N_9366,N_8110);
or U12014 (N_12014,N_8852,N_6661);
xor U12015 (N_12015,N_9950,N_7297);
nand U12016 (N_12016,N_5567,N_9184);
nor U12017 (N_12017,N_5243,N_9458);
or U12018 (N_12018,N_5246,N_9122);
or U12019 (N_12019,N_5923,N_9176);
nand U12020 (N_12020,N_5425,N_7605);
nor U12021 (N_12021,N_6606,N_9507);
and U12022 (N_12022,N_6242,N_8226);
nand U12023 (N_12023,N_7467,N_9981);
or U12024 (N_12024,N_6387,N_6353);
or U12025 (N_12025,N_7111,N_8183);
xor U12026 (N_12026,N_7378,N_6709);
nand U12027 (N_12027,N_9474,N_5859);
nand U12028 (N_12028,N_8150,N_8517);
nand U12029 (N_12029,N_9082,N_6768);
or U12030 (N_12030,N_6889,N_8117);
and U12031 (N_12031,N_9224,N_8856);
or U12032 (N_12032,N_8383,N_8198);
nand U12033 (N_12033,N_5111,N_8023);
nor U12034 (N_12034,N_9698,N_7587);
xor U12035 (N_12035,N_7000,N_8488);
and U12036 (N_12036,N_7187,N_8773);
nand U12037 (N_12037,N_5541,N_8839);
and U12038 (N_12038,N_7362,N_6720);
nor U12039 (N_12039,N_8481,N_9367);
nand U12040 (N_12040,N_9412,N_9278);
or U12041 (N_12041,N_8277,N_7913);
and U12042 (N_12042,N_5168,N_8525);
or U12043 (N_12043,N_6058,N_9922);
nand U12044 (N_12044,N_5281,N_7340);
nor U12045 (N_12045,N_8235,N_8505);
xor U12046 (N_12046,N_5310,N_9177);
and U12047 (N_12047,N_7728,N_7447);
and U12048 (N_12048,N_9735,N_5476);
nand U12049 (N_12049,N_7829,N_9009);
nor U12050 (N_12050,N_8921,N_7751);
or U12051 (N_12051,N_5994,N_6300);
nor U12052 (N_12052,N_5865,N_5755);
xnor U12053 (N_12053,N_8685,N_8770);
or U12054 (N_12054,N_9382,N_7959);
nor U12055 (N_12055,N_7015,N_6422);
xor U12056 (N_12056,N_9647,N_7916);
and U12057 (N_12057,N_6834,N_7410);
nor U12058 (N_12058,N_8738,N_5069);
and U12059 (N_12059,N_8422,N_6596);
xnor U12060 (N_12060,N_5301,N_8946);
nor U12061 (N_12061,N_8533,N_6663);
nor U12062 (N_12062,N_5547,N_6687);
and U12063 (N_12063,N_6147,N_7580);
or U12064 (N_12064,N_9058,N_9832);
nor U12065 (N_12065,N_7395,N_8478);
nand U12066 (N_12066,N_5137,N_7851);
nand U12067 (N_12067,N_5971,N_8882);
nand U12068 (N_12068,N_6369,N_7032);
or U12069 (N_12069,N_5600,N_7169);
nand U12070 (N_12070,N_5823,N_8138);
or U12071 (N_12071,N_5855,N_5627);
nor U12072 (N_12072,N_9038,N_6603);
and U12073 (N_12073,N_5842,N_5502);
nor U12074 (N_12074,N_7150,N_9558);
nand U12075 (N_12075,N_8766,N_7190);
and U12076 (N_12076,N_6867,N_8728);
or U12077 (N_12077,N_8396,N_6276);
nor U12078 (N_12078,N_5059,N_7390);
nand U12079 (N_12079,N_9048,N_7343);
or U12080 (N_12080,N_6890,N_5040);
nand U12081 (N_12081,N_6791,N_5856);
nand U12082 (N_12082,N_9232,N_6284);
nor U12083 (N_12083,N_8439,N_6343);
nand U12084 (N_12084,N_6287,N_7984);
nor U12085 (N_12085,N_6271,N_5510);
nand U12086 (N_12086,N_6827,N_7347);
or U12087 (N_12087,N_8635,N_7293);
nor U12088 (N_12088,N_6136,N_7439);
nand U12089 (N_12089,N_9346,N_9059);
nand U12090 (N_12090,N_6657,N_9874);
or U12091 (N_12091,N_9393,N_9029);
and U12092 (N_12092,N_6656,N_8807);
xnor U12093 (N_12093,N_6595,N_5862);
nand U12094 (N_12094,N_6740,N_8084);
or U12095 (N_12095,N_6393,N_8243);
nor U12096 (N_12096,N_5530,N_9868);
nor U12097 (N_12097,N_5670,N_6307);
nor U12098 (N_12098,N_7629,N_6214);
and U12099 (N_12099,N_8134,N_8337);
or U12100 (N_12100,N_7448,N_6246);
and U12101 (N_12101,N_9013,N_5911);
and U12102 (N_12102,N_9006,N_6431);
nand U12103 (N_12103,N_7364,N_5403);
nand U12104 (N_12104,N_7843,N_5912);
nor U12105 (N_12105,N_5400,N_8809);
and U12106 (N_12106,N_6095,N_7357);
and U12107 (N_12107,N_9572,N_5888);
and U12108 (N_12108,N_8141,N_6204);
nor U12109 (N_12109,N_7961,N_7826);
nor U12110 (N_12110,N_8672,N_6338);
nor U12111 (N_12111,N_6571,N_8923);
xnor U12112 (N_12112,N_8403,N_8982);
and U12113 (N_12113,N_9730,N_8159);
and U12114 (N_12114,N_6360,N_6840);
nor U12115 (N_12115,N_8919,N_7526);
nor U12116 (N_12116,N_6797,N_5171);
and U12117 (N_12117,N_6744,N_7302);
xor U12118 (N_12118,N_8427,N_8931);
nand U12119 (N_12119,N_9277,N_7181);
nand U12120 (N_12120,N_7100,N_9601);
xnor U12121 (N_12121,N_6401,N_8991);
and U12122 (N_12122,N_9036,N_9937);
nand U12123 (N_12123,N_5944,N_8740);
nor U12124 (N_12124,N_7318,N_5125);
or U12125 (N_12125,N_5060,N_5512);
nor U12126 (N_12126,N_6176,N_9425);
nand U12127 (N_12127,N_7664,N_8257);
and U12128 (N_12128,N_8528,N_8343);
xor U12129 (N_12129,N_9430,N_5357);
or U12130 (N_12130,N_8224,N_5639);
nor U12131 (N_12131,N_7768,N_8508);
and U12132 (N_12132,N_9234,N_8057);
xnor U12133 (N_12133,N_9531,N_6991);
and U12134 (N_12134,N_6737,N_8275);
and U12135 (N_12135,N_8368,N_6585);
nand U12136 (N_12136,N_7087,N_6133);
or U12137 (N_12137,N_6717,N_8137);
nand U12138 (N_12138,N_5977,N_6798);
and U12139 (N_12139,N_6910,N_9019);
nor U12140 (N_12140,N_5528,N_6301);
nor U12141 (N_12141,N_7711,N_8538);
or U12142 (N_12142,N_9837,N_9350);
or U12143 (N_12143,N_5459,N_8049);
or U12144 (N_12144,N_6682,N_6045);
nand U12145 (N_12145,N_6026,N_5216);
nand U12146 (N_12146,N_6703,N_8063);
nor U12147 (N_12147,N_8883,N_6500);
or U12148 (N_12148,N_8214,N_7049);
nor U12149 (N_12149,N_6508,N_8139);
or U12150 (N_12150,N_6390,N_9772);
nor U12151 (N_12151,N_7875,N_8490);
nand U12152 (N_12152,N_9973,N_5894);
nor U12153 (N_12153,N_9901,N_7058);
nand U12154 (N_12154,N_8314,N_9693);
or U12155 (N_12155,N_5986,N_7404);
nand U12156 (N_12156,N_6904,N_9107);
or U12157 (N_12157,N_8667,N_6029);
or U12158 (N_12158,N_8494,N_8010);
or U12159 (N_12159,N_7321,N_8306);
nand U12160 (N_12160,N_6610,N_9410);
or U12161 (N_12161,N_6319,N_7277);
nor U12162 (N_12162,N_8623,N_6855);
and U12163 (N_12163,N_8026,N_5438);
nand U12164 (N_12164,N_8462,N_5230);
nand U12165 (N_12165,N_8115,N_6658);
nand U12166 (N_12166,N_5135,N_7921);
nor U12167 (N_12167,N_8316,N_7127);
or U12168 (N_12168,N_9100,N_8854);
xor U12169 (N_12169,N_5864,N_7544);
nor U12170 (N_12170,N_9415,N_5506);
and U12171 (N_12171,N_9260,N_7958);
or U12172 (N_12172,N_6776,N_6753);
or U12173 (N_12173,N_6580,N_8430);
nand U12174 (N_12174,N_5985,N_6570);
xor U12175 (N_12175,N_9916,N_7454);
nand U12176 (N_12176,N_8653,N_7253);
and U12177 (N_12177,N_9166,N_8631);
and U12178 (N_12178,N_9935,N_9596);
or U12179 (N_12179,N_7066,N_9293);
nand U12180 (N_12180,N_9472,N_6049);
nand U12181 (N_12181,N_6984,N_8147);
and U12182 (N_12182,N_9492,N_5602);
and U12183 (N_12183,N_9517,N_7638);
nand U12184 (N_12184,N_9715,N_5941);
xnor U12185 (N_12185,N_5560,N_5766);
and U12186 (N_12186,N_9190,N_9843);
xnor U12187 (N_12187,N_7606,N_5107);
xor U12188 (N_12188,N_9439,N_7995);
nand U12189 (N_12189,N_5242,N_8744);
and U12190 (N_12190,N_7980,N_6556);
or U12191 (N_12191,N_6229,N_8613);
and U12192 (N_12192,N_6174,N_9395);
and U12193 (N_12193,N_8555,N_5318);
or U12194 (N_12194,N_5486,N_8659);
nand U12195 (N_12195,N_8083,N_9903);
nand U12196 (N_12196,N_7156,N_9220);
nand U12197 (N_12197,N_6492,N_7660);
nand U12198 (N_12198,N_5558,N_7476);
nand U12199 (N_12199,N_7926,N_9764);
or U12200 (N_12200,N_8846,N_9633);
and U12201 (N_12201,N_6098,N_8109);
nand U12202 (N_12202,N_9117,N_9018);
and U12203 (N_12203,N_7488,N_5133);
nand U12204 (N_12204,N_9409,N_8491);
and U12205 (N_12205,N_8078,N_8124);
or U12206 (N_12206,N_7811,N_9180);
nand U12207 (N_12207,N_6166,N_5905);
and U12208 (N_12208,N_8842,N_5570);
nand U12209 (N_12209,N_9509,N_8577);
nor U12210 (N_12210,N_6738,N_7198);
and U12211 (N_12211,N_5058,N_9460);
nor U12212 (N_12212,N_8984,N_5525);
xor U12213 (N_12213,N_9598,N_9716);
or U12214 (N_12214,N_9470,N_6660);
and U12215 (N_12215,N_7207,N_9908);
nand U12216 (N_12216,N_8985,N_5063);
and U12217 (N_12217,N_8835,N_8121);
xor U12218 (N_12218,N_7630,N_7470);
nor U12219 (N_12219,N_8731,N_7489);
or U12220 (N_12220,N_8999,N_8973);
and U12221 (N_12221,N_5830,N_6662);
or U12222 (N_12222,N_9791,N_6507);
nand U12223 (N_12223,N_6335,N_6971);
and U12224 (N_12224,N_9369,N_9068);
and U12225 (N_12225,N_9060,N_6157);
or U12226 (N_12226,N_5709,N_9158);
and U12227 (N_12227,N_8250,N_5657);
nand U12228 (N_12228,N_6407,N_7412);
or U12229 (N_12229,N_6017,N_6104);
or U12230 (N_12230,N_5282,N_9924);
nand U12231 (N_12231,N_6649,N_8404);
and U12232 (N_12232,N_6458,N_6455);
or U12233 (N_12233,N_7542,N_5363);
nand U12234 (N_12234,N_9654,N_7761);
or U12235 (N_12235,N_6511,N_5795);
nor U12236 (N_12236,N_7570,N_6472);
nor U12237 (N_12237,N_6575,N_6528);
nor U12238 (N_12238,N_8034,N_6860);
or U12239 (N_12239,N_7555,N_6731);
nand U12240 (N_12240,N_8061,N_5312);
and U12241 (N_12241,N_6320,N_9694);
and U12242 (N_12242,N_6654,N_9064);
and U12243 (N_12243,N_5796,N_8126);
or U12244 (N_12244,N_9203,N_8456);
nor U12245 (N_12245,N_7815,N_5516);
and U12246 (N_12246,N_6047,N_7590);
and U12247 (N_12247,N_7307,N_8485);
and U12248 (N_12248,N_9265,N_7500);
xnor U12249 (N_12249,N_8915,N_7493);
xor U12250 (N_12250,N_8584,N_5213);
nand U12251 (N_12251,N_7176,N_6209);
or U12252 (N_12252,N_8779,N_5511);
nand U12253 (N_12253,N_5448,N_7096);
or U12254 (N_12254,N_5565,N_5928);
xor U12255 (N_12255,N_7625,N_8600);
or U12256 (N_12256,N_5843,N_6824);
xnor U12257 (N_12257,N_7274,N_8438);
xnor U12258 (N_12258,N_9816,N_5964);
nor U12259 (N_12259,N_6138,N_9146);
nor U12260 (N_12260,N_7909,N_9423);
xnor U12261 (N_12261,N_8619,N_8573);
or U12262 (N_12262,N_8342,N_5641);
nand U12263 (N_12263,N_9330,N_6766);
or U12264 (N_12264,N_8670,N_7787);
or U12265 (N_12265,N_6411,N_9072);
or U12266 (N_12266,N_8385,N_7967);
and U12267 (N_12267,N_5604,N_6195);
nor U12268 (N_12268,N_6749,N_9997);
nand U12269 (N_12269,N_5841,N_6918);
nor U12270 (N_12270,N_7020,N_6877);
xor U12271 (N_12271,N_9978,N_8500);
nor U12272 (N_12272,N_6273,N_7762);
nor U12273 (N_12273,N_5015,N_9246);
and U12274 (N_12274,N_6100,N_5953);
or U12275 (N_12275,N_5493,N_9554);
or U12276 (N_12276,N_7119,N_5598);
nor U12277 (N_12277,N_7703,N_6755);
nor U12278 (N_12278,N_8959,N_9327);
and U12279 (N_12279,N_9699,N_9231);
nor U12280 (N_12280,N_5951,N_9162);
and U12281 (N_12281,N_6306,N_6938);
nand U12282 (N_12282,N_6218,N_6879);
and U12283 (N_12283,N_8280,N_5256);
and U12284 (N_12284,N_5028,N_5255);
xnor U12285 (N_12285,N_5349,N_7310);
nand U12286 (N_12286,N_9591,N_9173);
nor U12287 (N_12287,N_7983,N_7366);
or U12288 (N_12288,N_5735,N_9020);
nand U12289 (N_12289,N_7624,N_9451);
nor U12290 (N_12290,N_9541,N_6067);
and U12291 (N_12291,N_5608,N_5773);
nand U12292 (N_12292,N_8569,N_5162);
nand U12293 (N_12293,N_6332,N_8157);
nand U12294 (N_12294,N_6676,N_5848);
nand U12295 (N_12295,N_6854,N_6651);
nor U12296 (N_12296,N_6843,N_8312);
nand U12297 (N_12297,N_6254,N_8102);
and U12298 (N_12298,N_7739,N_8786);
xnor U12299 (N_12299,N_6121,N_5188);
nor U12300 (N_12300,N_6547,N_8676);
and U12301 (N_12301,N_8238,N_6354);
xnor U12302 (N_12302,N_9800,N_8753);
or U12303 (N_12303,N_6277,N_9299);
nand U12304 (N_12304,N_5068,N_8993);
nand U12305 (N_12305,N_7963,N_6812);
or U12306 (N_12306,N_6675,N_8068);
and U12307 (N_12307,N_5757,N_8966);
xor U12308 (N_12308,N_7185,N_9603);
xor U12309 (N_12309,N_7146,N_9104);
or U12310 (N_12310,N_5373,N_7749);
xor U12311 (N_12311,N_6977,N_6061);
or U12312 (N_12312,N_6735,N_8131);
and U12313 (N_12313,N_5096,N_6535);
or U12314 (N_12314,N_9556,N_5035);
nand U12315 (N_12315,N_5714,N_8158);
nor U12316 (N_12316,N_8202,N_6701);
nand U12317 (N_12317,N_9595,N_8711);
nand U12318 (N_12318,N_9734,N_7048);
and U12319 (N_12319,N_7795,N_5746);
nand U12320 (N_12320,N_7233,N_6220);
and U12321 (N_12321,N_8648,N_8464);
nand U12322 (N_12322,N_7055,N_8360);
or U12323 (N_12323,N_6522,N_8639);
and U12324 (N_12324,N_6365,N_7543);
nor U12325 (N_12325,N_5465,N_5697);
nor U12326 (N_12326,N_6647,N_5633);
nor U12327 (N_12327,N_9970,N_5492);
xnor U12328 (N_12328,N_7825,N_5434);
nand U12329 (N_12329,N_8927,N_7911);
nor U12330 (N_12330,N_7982,N_9239);
nand U12331 (N_12331,N_5287,N_5335);
xnor U12332 (N_12332,N_7782,N_5653);
xor U12333 (N_12333,N_9362,N_9142);
nor U12334 (N_12334,N_7244,N_5369);
nand U12335 (N_12335,N_8129,N_7670);
nand U12336 (N_12336,N_5038,N_7516);
nor U12337 (N_12337,N_6223,N_9311);
nor U12338 (N_12338,N_5878,N_5587);
or U12339 (N_12339,N_9175,N_6184);
nand U12340 (N_12340,N_9135,N_5559);
or U12341 (N_12341,N_5338,N_7046);
nand U12342 (N_12342,N_9372,N_9375);
nor U12343 (N_12343,N_5376,N_9544);
nor U12344 (N_12344,N_8588,N_5957);
nand U12345 (N_12345,N_5712,N_5809);
nor U12346 (N_12346,N_7243,N_8911);
xor U12347 (N_12347,N_9461,N_6962);
or U12348 (N_12348,N_9179,N_5129);
nor U12349 (N_12349,N_7221,N_5088);
nand U12350 (N_12350,N_9191,N_8411);
and U12351 (N_12351,N_9221,N_7090);
or U12352 (N_12352,N_5226,N_5914);
nand U12353 (N_12353,N_7743,N_6957);
nand U12354 (N_12354,N_9079,N_6513);
or U12355 (N_12355,N_6699,N_5260);
nand U12356 (N_12356,N_6769,N_5720);
and U12357 (N_12357,N_7197,N_8120);
nor U12358 (N_12358,N_8001,N_7262);
and U12359 (N_12359,N_5580,N_6940);
xnor U12360 (N_12360,N_6552,N_9040);
nor U12361 (N_12361,N_6622,N_9049);
or U12362 (N_12362,N_7807,N_5611);
nor U12363 (N_12363,N_5156,N_6582);
nand U12364 (N_12364,N_8970,N_5032);
nor U12365 (N_12365,N_8643,N_7764);
xor U12366 (N_12366,N_8743,N_5432);
nand U12367 (N_12367,N_8252,N_6590);
nand U12368 (N_12368,N_8795,N_5077);
xnor U12369 (N_12369,N_8897,N_9702);
xnor U12370 (N_12370,N_5117,N_9054);
nor U12371 (N_12371,N_8675,N_5553);
and U12372 (N_12372,N_9912,N_8903);
nand U12373 (N_12373,N_7945,N_9921);
xor U12374 (N_12374,N_6819,N_6106);
and U12375 (N_12375,N_6598,N_7731);
nor U12376 (N_12376,N_6545,N_7989);
and U12377 (N_12377,N_9163,N_9157);
nor U12378 (N_12378,N_5852,N_8727);
or U12379 (N_12379,N_6403,N_6298);
nand U12380 (N_12380,N_5221,N_9428);
xor U12381 (N_12381,N_5886,N_5113);
nor U12382 (N_12382,N_6967,N_5684);
nand U12383 (N_12383,N_9388,N_6536);
nor U12384 (N_12384,N_7576,N_6351);
nor U12385 (N_12385,N_8397,N_6820);
or U12386 (N_12386,N_6337,N_8236);
and U12387 (N_12387,N_6120,N_7009);
and U12388 (N_12388,N_8988,N_7417);
or U12389 (N_12389,N_5818,N_9947);
and U12390 (N_12390,N_7217,N_6982);
and U12391 (N_12391,N_9537,N_6826);
and U12392 (N_12392,N_7757,N_7042);
nor U12393 (N_12393,N_6983,N_8096);
nor U12394 (N_12394,N_7206,N_8082);
nand U12395 (N_12395,N_9237,N_6386);
or U12396 (N_12396,N_7304,N_6736);
nand U12397 (N_12397,N_6007,N_9349);
nor U12398 (N_12398,N_8983,N_6072);
xnor U12399 (N_12399,N_9042,N_9638);
and U12400 (N_12400,N_8871,N_7332);
or U12401 (N_12401,N_7001,N_8755);
nand U12402 (N_12402,N_7855,N_5419);
xor U12403 (N_12403,N_5008,N_7134);
or U12404 (N_12404,N_5462,N_9351);
or U12405 (N_12405,N_7202,N_7723);
nor U12406 (N_12406,N_7133,N_7900);
and U12407 (N_12407,N_8308,N_7405);
nand U12408 (N_12408,N_9792,N_6851);
or U12409 (N_12409,N_5285,N_5067);
and U12410 (N_12410,N_7441,N_7668);
nor U12411 (N_12411,N_9826,N_8509);
xor U12412 (N_12412,N_6562,N_5350);
and U12413 (N_12413,N_9116,N_7420);
nand U12414 (N_12414,N_8681,N_9271);
nand U12415 (N_12415,N_7351,N_9475);
or U12416 (N_12416,N_7672,N_9626);
nor U12417 (N_12417,N_8621,N_5584);
nand U12418 (N_12418,N_5866,N_8266);
nor U12419 (N_12419,N_5694,N_8324);
nor U12420 (N_12420,N_8380,N_6419);
and U12421 (N_12421,N_8148,N_9683);
nor U12422 (N_12422,N_9828,N_5479);
nor U12423 (N_12423,N_7608,N_6733);
nand U12424 (N_12424,N_8076,N_9323);
or U12425 (N_12425,N_6315,N_8196);
nand U12426 (N_12426,N_9345,N_9965);
or U12427 (N_12427,N_5016,N_5840);
nor U12428 (N_12428,N_7078,N_7432);
nand U12429 (N_12429,N_6410,N_8501);
nand U12430 (N_12430,N_8909,N_6587);
nor U12431 (N_12431,N_6040,N_6205);
or U12432 (N_12432,N_5214,N_6655);
nor U12433 (N_12433,N_8402,N_5359);
and U12434 (N_12434,N_5352,N_7527);
nor U12435 (N_12435,N_8493,N_5814);
xor U12436 (N_12436,N_5456,N_8772);
or U12437 (N_12437,N_8433,N_6457);
or U12438 (N_12438,N_5981,N_6233);
xnor U12439 (N_12439,N_9429,N_7885);
nand U12440 (N_12440,N_7546,N_6546);
nor U12441 (N_12441,N_6355,N_6217);
nor U12442 (N_12442,N_9386,N_6921);
and U12443 (N_12443,N_7709,N_9954);
or U12444 (N_12444,N_9527,N_8267);
nand U12445 (N_12445,N_6935,N_9838);
nor U12446 (N_12446,N_9457,N_8791);
or U12447 (N_12447,N_5740,N_9435);
nand U12448 (N_12448,N_5204,N_7771);
or U12449 (N_12449,N_9263,N_6474);
xnor U12450 (N_12450,N_7805,N_5593);
and U12451 (N_12451,N_7264,N_9332);
or U12452 (N_12452,N_6349,N_5437);
and U12453 (N_12453,N_8737,N_7520);
or U12454 (N_12454,N_8705,N_6373);
nand U12455 (N_12455,N_7993,N_6096);
and U12456 (N_12456,N_8154,N_7869);
and U12457 (N_12457,N_8099,N_7229);
or U12458 (N_12458,N_8492,N_7691);
or U12459 (N_12459,N_5929,N_7976);
and U12460 (N_12460,N_8718,N_5521);
nor U12461 (N_12461,N_6346,N_5764);
nor U12462 (N_12462,N_5745,N_5340);
nand U12463 (N_12463,N_9794,N_8634);
nand U12464 (N_12464,N_7465,N_6361);
or U12465 (N_12465,N_9784,N_5625);
xor U12466 (N_12466,N_6211,N_6011);
nor U12467 (N_12467,N_7466,N_7694);
nor U12468 (N_12468,N_8960,N_5901);
and U12469 (N_12469,N_5051,N_9494);
and U12470 (N_12470,N_6057,N_5089);
nand U12471 (N_12471,N_6684,N_5829);
xnor U12472 (N_12472,N_8605,N_7284);
nor U12473 (N_12473,N_6969,N_8244);
or U12474 (N_12474,N_8887,N_8366);
nor U12475 (N_12475,N_7681,N_5819);
nor U12476 (N_12476,N_9481,N_6409);
or U12477 (N_12477,N_7065,N_5211);
and U12478 (N_12478,N_6694,N_5441);
xor U12479 (N_12479,N_6069,N_7296);
nor U12480 (N_12480,N_6551,N_8401);
or U12481 (N_12481,N_5692,N_5526);
and U12482 (N_12482,N_7008,N_7086);
or U12483 (N_12483,N_6083,N_9881);
and U12484 (N_12484,N_7553,N_9748);
or U12485 (N_12485,N_8066,N_9436);
or U12486 (N_12486,N_7944,N_7951);
xnor U12487 (N_12487,N_6243,N_9266);
and U12488 (N_12488,N_9249,N_8217);
nand U12489 (N_12489,N_8512,N_6965);
nor U12490 (N_12490,N_7327,N_9768);
nand U12491 (N_12491,N_7714,N_9501);
xor U12492 (N_12492,N_8191,N_5324);
nand U12493 (N_12493,N_8155,N_7895);
or U12494 (N_12494,N_6905,N_7985);
nand U12495 (N_12495,N_9418,N_8688);
nand U12496 (N_12496,N_6264,N_7105);
nor U12497 (N_12497,N_7033,N_8009);
nor U12498 (N_12498,N_6385,N_8237);
and U12499 (N_12499,N_6055,N_5933);
or U12500 (N_12500,N_8612,N_8655);
xnor U12501 (N_12501,N_9665,N_5895);
or U12502 (N_12502,N_8745,N_6016);
nor U12503 (N_12503,N_5486,N_7331);
or U12504 (N_12504,N_9000,N_7208);
nor U12505 (N_12505,N_9010,N_9517);
nand U12506 (N_12506,N_9471,N_8806);
nor U12507 (N_12507,N_7582,N_9818);
nor U12508 (N_12508,N_6859,N_9336);
xnor U12509 (N_12509,N_8720,N_6962);
nor U12510 (N_12510,N_5827,N_7429);
nor U12511 (N_12511,N_5415,N_5331);
nor U12512 (N_12512,N_9650,N_5669);
nand U12513 (N_12513,N_8232,N_7540);
nor U12514 (N_12514,N_8006,N_8764);
and U12515 (N_12515,N_7927,N_5895);
nor U12516 (N_12516,N_8190,N_7190);
nor U12517 (N_12517,N_6060,N_8789);
nor U12518 (N_12518,N_8009,N_6105);
and U12519 (N_12519,N_5143,N_9587);
or U12520 (N_12520,N_7473,N_8414);
nor U12521 (N_12521,N_5731,N_9284);
nand U12522 (N_12522,N_5202,N_7959);
or U12523 (N_12523,N_9748,N_7793);
nand U12524 (N_12524,N_8433,N_5805);
and U12525 (N_12525,N_6429,N_9132);
nand U12526 (N_12526,N_5365,N_7314);
nand U12527 (N_12527,N_8386,N_7968);
and U12528 (N_12528,N_8898,N_8944);
nand U12529 (N_12529,N_7320,N_8617);
nor U12530 (N_12530,N_7459,N_7710);
nor U12531 (N_12531,N_7711,N_5808);
nor U12532 (N_12532,N_7739,N_8669);
nand U12533 (N_12533,N_9522,N_6248);
and U12534 (N_12534,N_8805,N_9738);
nor U12535 (N_12535,N_9305,N_5243);
nand U12536 (N_12536,N_7086,N_8851);
and U12537 (N_12537,N_9977,N_5728);
nand U12538 (N_12538,N_6363,N_7507);
nand U12539 (N_12539,N_9870,N_8518);
nand U12540 (N_12540,N_9273,N_8655);
and U12541 (N_12541,N_9509,N_8328);
xor U12542 (N_12542,N_9671,N_8643);
or U12543 (N_12543,N_5698,N_7085);
nor U12544 (N_12544,N_8679,N_8601);
nor U12545 (N_12545,N_6294,N_7068);
or U12546 (N_12546,N_7894,N_5325);
nor U12547 (N_12547,N_7618,N_5678);
or U12548 (N_12548,N_7807,N_6755);
nor U12549 (N_12549,N_6795,N_9400);
and U12550 (N_12550,N_8995,N_7012);
nand U12551 (N_12551,N_8776,N_8202);
and U12552 (N_12552,N_8987,N_9972);
nor U12553 (N_12553,N_8539,N_7927);
nand U12554 (N_12554,N_8162,N_9738);
nand U12555 (N_12555,N_7886,N_9852);
nor U12556 (N_12556,N_6487,N_8020);
nand U12557 (N_12557,N_5464,N_8422);
xnor U12558 (N_12558,N_5137,N_8996);
nand U12559 (N_12559,N_8528,N_9639);
and U12560 (N_12560,N_5171,N_6273);
or U12561 (N_12561,N_5723,N_5255);
or U12562 (N_12562,N_7356,N_7284);
or U12563 (N_12563,N_8067,N_7065);
or U12564 (N_12564,N_6657,N_7987);
or U12565 (N_12565,N_6392,N_7138);
xnor U12566 (N_12566,N_5823,N_9222);
nand U12567 (N_12567,N_6952,N_7556);
nand U12568 (N_12568,N_5935,N_8879);
xnor U12569 (N_12569,N_9831,N_6592);
nor U12570 (N_12570,N_8353,N_5400);
xnor U12571 (N_12571,N_6154,N_9837);
xnor U12572 (N_12572,N_7244,N_6692);
nor U12573 (N_12573,N_8207,N_9694);
nand U12574 (N_12574,N_5434,N_6109);
nor U12575 (N_12575,N_5889,N_7867);
or U12576 (N_12576,N_7046,N_9774);
xnor U12577 (N_12577,N_6627,N_6875);
nor U12578 (N_12578,N_9010,N_8561);
and U12579 (N_12579,N_9166,N_6748);
nor U12580 (N_12580,N_7396,N_7559);
nand U12581 (N_12581,N_8390,N_6512);
and U12582 (N_12582,N_9458,N_5770);
nor U12583 (N_12583,N_9040,N_9027);
or U12584 (N_12584,N_8127,N_8493);
and U12585 (N_12585,N_9696,N_7769);
nor U12586 (N_12586,N_6452,N_6674);
nand U12587 (N_12587,N_9773,N_5783);
xor U12588 (N_12588,N_8041,N_6390);
nand U12589 (N_12589,N_6478,N_7196);
xor U12590 (N_12590,N_5974,N_9884);
nor U12591 (N_12591,N_8379,N_8507);
nand U12592 (N_12592,N_5593,N_6956);
nor U12593 (N_12593,N_9922,N_5359);
and U12594 (N_12594,N_7383,N_6495);
and U12595 (N_12595,N_9620,N_5552);
and U12596 (N_12596,N_7241,N_8153);
nor U12597 (N_12597,N_7765,N_7377);
xor U12598 (N_12598,N_9875,N_6659);
and U12599 (N_12599,N_6948,N_8378);
or U12600 (N_12600,N_5733,N_8099);
or U12601 (N_12601,N_9917,N_8675);
xor U12602 (N_12602,N_7690,N_7316);
nor U12603 (N_12603,N_8459,N_8084);
nand U12604 (N_12604,N_5669,N_8580);
xor U12605 (N_12605,N_6889,N_7860);
nand U12606 (N_12606,N_6308,N_5786);
nand U12607 (N_12607,N_6634,N_9771);
xnor U12608 (N_12608,N_6604,N_7515);
nand U12609 (N_12609,N_7740,N_6108);
nor U12610 (N_12610,N_8536,N_8167);
nand U12611 (N_12611,N_6184,N_9774);
nor U12612 (N_12612,N_5874,N_8679);
xor U12613 (N_12613,N_7137,N_7722);
and U12614 (N_12614,N_9315,N_8684);
nor U12615 (N_12615,N_5673,N_8849);
nor U12616 (N_12616,N_6520,N_7541);
nand U12617 (N_12617,N_6029,N_5506);
xor U12618 (N_12618,N_9864,N_8050);
and U12619 (N_12619,N_8146,N_8299);
nand U12620 (N_12620,N_7402,N_9209);
nand U12621 (N_12621,N_7529,N_7393);
nor U12622 (N_12622,N_7809,N_9734);
and U12623 (N_12623,N_9230,N_9447);
or U12624 (N_12624,N_8756,N_5634);
xnor U12625 (N_12625,N_6627,N_6107);
nor U12626 (N_12626,N_5831,N_7901);
and U12627 (N_12627,N_8546,N_8790);
or U12628 (N_12628,N_8511,N_9314);
or U12629 (N_12629,N_5835,N_9008);
and U12630 (N_12630,N_5500,N_8765);
xnor U12631 (N_12631,N_8029,N_7707);
nand U12632 (N_12632,N_8590,N_8683);
or U12633 (N_12633,N_5581,N_7003);
nand U12634 (N_12634,N_8563,N_5308);
or U12635 (N_12635,N_9606,N_9027);
xor U12636 (N_12636,N_7050,N_5410);
or U12637 (N_12637,N_5092,N_9839);
xnor U12638 (N_12638,N_7853,N_9792);
or U12639 (N_12639,N_8508,N_6440);
and U12640 (N_12640,N_8933,N_8875);
and U12641 (N_12641,N_5683,N_7510);
nand U12642 (N_12642,N_6565,N_7445);
nand U12643 (N_12643,N_6248,N_8195);
or U12644 (N_12644,N_9103,N_9606);
xor U12645 (N_12645,N_9425,N_9096);
and U12646 (N_12646,N_5643,N_6494);
nor U12647 (N_12647,N_8350,N_5324);
and U12648 (N_12648,N_8103,N_7932);
and U12649 (N_12649,N_8415,N_5931);
or U12650 (N_12650,N_8904,N_7507);
and U12651 (N_12651,N_7523,N_8916);
and U12652 (N_12652,N_5789,N_8459);
and U12653 (N_12653,N_9987,N_7666);
nand U12654 (N_12654,N_6364,N_9557);
nand U12655 (N_12655,N_7301,N_8632);
or U12656 (N_12656,N_6582,N_7635);
nand U12657 (N_12657,N_5104,N_8605);
and U12658 (N_12658,N_8916,N_9169);
or U12659 (N_12659,N_7258,N_8846);
and U12660 (N_12660,N_8054,N_7801);
or U12661 (N_12661,N_6108,N_5703);
or U12662 (N_12662,N_5895,N_5932);
nor U12663 (N_12663,N_7870,N_7685);
or U12664 (N_12664,N_7529,N_8764);
and U12665 (N_12665,N_5855,N_5743);
and U12666 (N_12666,N_5053,N_7274);
xor U12667 (N_12667,N_8296,N_6482);
nand U12668 (N_12668,N_9840,N_6691);
nor U12669 (N_12669,N_9186,N_7920);
nor U12670 (N_12670,N_6369,N_9415);
nand U12671 (N_12671,N_9768,N_5537);
nand U12672 (N_12672,N_5039,N_9988);
nor U12673 (N_12673,N_5628,N_8272);
nand U12674 (N_12674,N_6678,N_6917);
or U12675 (N_12675,N_8421,N_5511);
and U12676 (N_12676,N_9571,N_6751);
nor U12677 (N_12677,N_8735,N_6918);
nor U12678 (N_12678,N_5423,N_7388);
nand U12679 (N_12679,N_7047,N_8232);
and U12680 (N_12680,N_6175,N_5252);
nor U12681 (N_12681,N_9018,N_8818);
and U12682 (N_12682,N_6524,N_5130);
nand U12683 (N_12683,N_6720,N_8202);
and U12684 (N_12684,N_6483,N_5479);
or U12685 (N_12685,N_9580,N_7227);
nor U12686 (N_12686,N_6923,N_6867);
nand U12687 (N_12687,N_8692,N_6487);
nor U12688 (N_12688,N_8206,N_8865);
or U12689 (N_12689,N_7783,N_8180);
or U12690 (N_12690,N_5732,N_5392);
nor U12691 (N_12691,N_5080,N_8897);
nand U12692 (N_12692,N_9560,N_6557);
or U12693 (N_12693,N_8975,N_6013);
or U12694 (N_12694,N_8642,N_6842);
or U12695 (N_12695,N_5589,N_5875);
xor U12696 (N_12696,N_8980,N_6073);
nor U12697 (N_12697,N_9064,N_9994);
nand U12698 (N_12698,N_9100,N_6450);
or U12699 (N_12699,N_6462,N_5314);
and U12700 (N_12700,N_5483,N_6834);
or U12701 (N_12701,N_5212,N_5095);
or U12702 (N_12702,N_5024,N_9459);
or U12703 (N_12703,N_9291,N_9948);
and U12704 (N_12704,N_9697,N_7413);
nor U12705 (N_12705,N_9843,N_9910);
or U12706 (N_12706,N_8510,N_5798);
or U12707 (N_12707,N_7352,N_8152);
or U12708 (N_12708,N_8819,N_5334);
or U12709 (N_12709,N_8953,N_8696);
nor U12710 (N_12710,N_9985,N_6687);
and U12711 (N_12711,N_8781,N_8135);
or U12712 (N_12712,N_6476,N_7318);
nor U12713 (N_12713,N_8481,N_6676);
xor U12714 (N_12714,N_5447,N_5056);
nand U12715 (N_12715,N_7028,N_7113);
nand U12716 (N_12716,N_8882,N_9867);
nor U12717 (N_12717,N_8313,N_6752);
or U12718 (N_12718,N_8789,N_5060);
and U12719 (N_12719,N_5883,N_7145);
or U12720 (N_12720,N_9541,N_8062);
nand U12721 (N_12721,N_5731,N_5922);
xor U12722 (N_12722,N_8900,N_7906);
nand U12723 (N_12723,N_9405,N_6681);
nor U12724 (N_12724,N_6472,N_9151);
nor U12725 (N_12725,N_7885,N_6499);
nor U12726 (N_12726,N_9127,N_6623);
and U12727 (N_12727,N_7662,N_9316);
nor U12728 (N_12728,N_7971,N_6864);
or U12729 (N_12729,N_9079,N_6448);
or U12730 (N_12730,N_5627,N_9905);
and U12731 (N_12731,N_8225,N_8993);
or U12732 (N_12732,N_8936,N_7007);
nor U12733 (N_12733,N_8237,N_6160);
or U12734 (N_12734,N_7771,N_8135);
and U12735 (N_12735,N_8887,N_7556);
nand U12736 (N_12736,N_8672,N_6164);
and U12737 (N_12737,N_7042,N_7481);
xnor U12738 (N_12738,N_7458,N_9519);
or U12739 (N_12739,N_5122,N_6224);
and U12740 (N_12740,N_9066,N_6339);
nand U12741 (N_12741,N_6280,N_8069);
or U12742 (N_12742,N_6214,N_7574);
nor U12743 (N_12743,N_8041,N_5538);
or U12744 (N_12744,N_8513,N_8507);
and U12745 (N_12745,N_7584,N_7531);
nor U12746 (N_12746,N_6770,N_5987);
nand U12747 (N_12747,N_6311,N_9413);
or U12748 (N_12748,N_7734,N_8385);
nand U12749 (N_12749,N_7168,N_8834);
or U12750 (N_12750,N_6422,N_6557);
nor U12751 (N_12751,N_9880,N_9153);
nand U12752 (N_12752,N_9373,N_6326);
xnor U12753 (N_12753,N_6289,N_6066);
or U12754 (N_12754,N_8280,N_7910);
and U12755 (N_12755,N_7096,N_5018);
and U12756 (N_12756,N_5613,N_8891);
nand U12757 (N_12757,N_7649,N_8535);
and U12758 (N_12758,N_5144,N_9562);
nor U12759 (N_12759,N_7487,N_6610);
nor U12760 (N_12760,N_8125,N_5176);
xor U12761 (N_12761,N_8782,N_9698);
nand U12762 (N_12762,N_7257,N_7316);
xor U12763 (N_12763,N_7962,N_7919);
xnor U12764 (N_12764,N_6509,N_9330);
and U12765 (N_12765,N_5563,N_6143);
nor U12766 (N_12766,N_9076,N_6818);
or U12767 (N_12767,N_8866,N_9927);
or U12768 (N_12768,N_6216,N_7444);
nor U12769 (N_12769,N_8820,N_7182);
nor U12770 (N_12770,N_7291,N_7164);
xnor U12771 (N_12771,N_6115,N_8296);
or U12772 (N_12772,N_5696,N_7220);
nand U12773 (N_12773,N_5357,N_6298);
nor U12774 (N_12774,N_6477,N_7953);
and U12775 (N_12775,N_5188,N_9016);
or U12776 (N_12776,N_6130,N_6478);
nand U12777 (N_12777,N_7624,N_9850);
and U12778 (N_12778,N_5965,N_5998);
or U12779 (N_12779,N_6244,N_9814);
nor U12780 (N_12780,N_9426,N_6496);
or U12781 (N_12781,N_6559,N_8971);
or U12782 (N_12782,N_7337,N_8573);
and U12783 (N_12783,N_9980,N_7313);
or U12784 (N_12784,N_8233,N_8843);
xor U12785 (N_12785,N_9765,N_5973);
xor U12786 (N_12786,N_9838,N_9577);
or U12787 (N_12787,N_7901,N_5625);
nand U12788 (N_12788,N_7994,N_9397);
or U12789 (N_12789,N_8412,N_8707);
nand U12790 (N_12790,N_8844,N_8410);
nand U12791 (N_12791,N_5038,N_6632);
nor U12792 (N_12792,N_9960,N_5332);
or U12793 (N_12793,N_6652,N_6523);
or U12794 (N_12794,N_5480,N_6353);
nand U12795 (N_12795,N_8836,N_6508);
nor U12796 (N_12796,N_5126,N_9905);
nand U12797 (N_12797,N_9264,N_8825);
nor U12798 (N_12798,N_8864,N_9694);
nor U12799 (N_12799,N_5854,N_7012);
and U12800 (N_12800,N_5046,N_5653);
nand U12801 (N_12801,N_5444,N_9040);
and U12802 (N_12802,N_5429,N_5054);
nor U12803 (N_12803,N_9570,N_6534);
xnor U12804 (N_12804,N_8726,N_8163);
and U12805 (N_12805,N_9582,N_5137);
nor U12806 (N_12806,N_9377,N_8893);
or U12807 (N_12807,N_7731,N_6001);
or U12808 (N_12808,N_5350,N_9467);
nor U12809 (N_12809,N_8466,N_9130);
nand U12810 (N_12810,N_8491,N_9717);
nand U12811 (N_12811,N_8177,N_7494);
or U12812 (N_12812,N_5117,N_6346);
nand U12813 (N_12813,N_5404,N_5687);
and U12814 (N_12814,N_8800,N_9255);
nor U12815 (N_12815,N_9091,N_9457);
nand U12816 (N_12816,N_6917,N_5146);
nand U12817 (N_12817,N_8223,N_5745);
nand U12818 (N_12818,N_8482,N_9280);
nand U12819 (N_12819,N_7954,N_5653);
and U12820 (N_12820,N_6573,N_5267);
nor U12821 (N_12821,N_6310,N_7079);
nor U12822 (N_12822,N_7402,N_6030);
and U12823 (N_12823,N_6667,N_5734);
nor U12824 (N_12824,N_6731,N_6127);
and U12825 (N_12825,N_7099,N_6212);
nor U12826 (N_12826,N_8444,N_8392);
xnor U12827 (N_12827,N_5514,N_6165);
and U12828 (N_12828,N_6834,N_8577);
nand U12829 (N_12829,N_6696,N_5947);
xor U12830 (N_12830,N_6266,N_8226);
nor U12831 (N_12831,N_5461,N_7136);
nand U12832 (N_12832,N_5380,N_5725);
nor U12833 (N_12833,N_5096,N_7768);
nor U12834 (N_12834,N_6386,N_5094);
xnor U12835 (N_12835,N_5189,N_5214);
nand U12836 (N_12836,N_6486,N_9377);
nand U12837 (N_12837,N_9452,N_5884);
nand U12838 (N_12838,N_8334,N_8632);
and U12839 (N_12839,N_8679,N_8672);
nand U12840 (N_12840,N_5668,N_9607);
or U12841 (N_12841,N_6941,N_5677);
nand U12842 (N_12842,N_9471,N_7758);
or U12843 (N_12843,N_8764,N_8600);
xnor U12844 (N_12844,N_5255,N_8465);
nor U12845 (N_12845,N_5786,N_5171);
nor U12846 (N_12846,N_7846,N_5882);
nor U12847 (N_12847,N_6312,N_7782);
nor U12848 (N_12848,N_7157,N_7523);
and U12849 (N_12849,N_6508,N_8941);
xor U12850 (N_12850,N_7925,N_9389);
nand U12851 (N_12851,N_5154,N_6038);
nor U12852 (N_12852,N_6543,N_6231);
or U12853 (N_12853,N_6239,N_9855);
or U12854 (N_12854,N_8790,N_6658);
and U12855 (N_12855,N_8891,N_7276);
xnor U12856 (N_12856,N_7831,N_5194);
xor U12857 (N_12857,N_9949,N_5497);
nand U12858 (N_12858,N_8473,N_5948);
or U12859 (N_12859,N_9218,N_8256);
nor U12860 (N_12860,N_5239,N_6004);
nand U12861 (N_12861,N_7029,N_9144);
nand U12862 (N_12862,N_9370,N_5203);
nor U12863 (N_12863,N_7990,N_5845);
or U12864 (N_12864,N_6620,N_8796);
nand U12865 (N_12865,N_8055,N_5035);
or U12866 (N_12866,N_6219,N_7962);
nand U12867 (N_12867,N_9403,N_8216);
nor U12868 (N_12868,N_8927,N_7866);
nand U12869 (N_12869,N_5591,N_9396);
and U12870 (N_12870,N_7395,N_5909);
nor U12871 (N_12871,N_9067,N_8840);
nand U12872 (N_12872,N_5760,N_5126);
or U12873 (N_12873,N_6020,N_8022);
nor U12874 (N_12874,N_9252,N_6737);
or U12875 (N_12875,N_5363,N_7131);
or U12876 (N_12876,N_9526,N_8576);
nand U12877 (N_12877,N_7625,N_5221);
xor U12878 (N_12878,N_5665,N_9675);
nor U12879 (N_12879,N_5667,N_5715);
or U12880 (N_12880,N_5211,N_5554);
and U12881 (N_12881,N_5316,N_5487);
nand U12882 (N_12882,N_5246,N_8880);
and U12883 (N_12883,N_9476,N_8174);
nor U12884 (N_12884,N_9262,N_8156);
or U12885 (N_12885,N_7537,N_9698);
nor U12886 (N_12886,N_7067,N_9376);
or U12887 (N_12887,N_9101,N_8674);
nand U12888 (N_12888,N_9217,N_5530);
xor U12889 (N_12889,N_9052,N_7769);
nor U12890 (N_12890,N_6458,N_8609);
nand U12891 (N_12891,N_5017,N_7755);
and U12892 (N_12892,N_6340,N_5617);
nor U12893 (N_12893,N_8715,N_7445);
or U12894 (N_12894,N_8276,N_8093);
nand U12895 (N_12895,N_8341,N_5155);
nor U12896 (N_12896,N_6045,N_6835);
or U12897 (N_12897,N_8521,N_7732);
and U12898 (N_12898,N_8065,N_8880);
or U12899 (N_12899,N_5214,N_8837);
nand U12900 (N_12900,N_5195,N_7379);
nor U12901 (N_12901,N_9137,N_9022);
nor U12902 (N_12902,N_5263,N_6317);
nor U12903 (N_12903,N_9742,N_9228);
nand U12904 (N_12904,N_6843,N_8714);
and U12905 (N_12905,N_6490,N_5714);
and U12906 (N_12906,N_6619,N_8226);
nand U12907 (N_12907,N_5838,N_7175);
and U12908 (N_12908,N_9229,N_9538);
or U12909 (N_12909,N_5050,N_9493);
xnor U12910 (N_12910,N_6240,N_7299);
nor U12911 (N_12911,N_7871,N_6503);
and U12912 (N_12912,N_9718,N_8623);
xor U12913 (N_12913,N_6899,N_9316);
nand U12914 (N_12914,N_5286,N_8483);
nor U12915 (N_12915,N_7051,N_5134);
nor U12916 (N_12916,N_7679,N_7296);
nand U12917 (N_12917,N_9321,N_9890);
nand U12918 (N_12918,N_5657,N_8492);
or U12919 (N_12919,N_8309,N_9798);
nor U12920 (N_12920,N_6416,N_9293);
or U12921 (N_12921,N_6376,N_8119);
and U12922 (N_12922,N_9269,N_6215);
and U12923 (N_12923,N_5848,N_6248);
nor U12924 (N_12924,N_5789,N_7659);
and U12925 (N_12925,N_8746,N_6568);
nand U12926 (N_12926,N_5888,N_7666);
nor U12927 (N_12927,N_6204,N_5533);
nor U12928 (N_12928,N_6655,N_5587);
and U12929 (N_12929,N_9459,N_6150);
nor U12930 (N_12930,N_8316,N_9101);
nor U12931 (N_12931,N_6111,N_7449);
or U12932 (N_12932,N_5742,N_7431);
or U12933 (N_12933,N_9412,N_5111);
and U12934 (N_12934,N_9695,N_5510);
or U12935 (N_12935,N_6903,N_7732);
nor U12936 (N_12936,N_8397,N_5768);
nor U12937 (N_12937,N_8934,N_9478);
or U12938 (N_12938,N_9652,N_9241);
and U12939 (N_12939,N_7695,N_9394);
and U12940 (N_12940,N_9999,N_7400);
or U12941 (N_12941,N_9966,N_6858);
nor U12942 (N_12942,N_5211,N_5025);
or U12943 (N_12943,N_5388,N_8029);
and U12944 (N_12944,N_7785,N_5064);
nand U12945 (N_12945,N_9535,N_6074);
and U12946 (N_12946,N_9608,N_8374);
xor U12947 (N_12947,N_6339,N_8234);
nand U12948 (N_12948,N_6051,N_7525);
or U12949 (N_12949,N_8089,N_9769);
and U12950 (N_12950,N_8914,N_5120);
nor U12951 (N_12951,N_9139,N_8201);
xnor U12952 (N_12952,N_5172,N_5706);
xor U12953 (N_12953,N_5527,N_5380);
and U12954 (N_12954,N_8920,N_6710);
or U12955 (N_12955,N_8374,N_8167);
nand U12956 (N_12956,N_5621,N_7456);
nor U12957 (N_12957,N_8060,N_8236);
or U12958 (N_12958,N_9538,N_9010);
and U12959 (N_12959,N_7223,N_8539);
nand U12960 (N_12960,N_6066,N_5698);
nand U12961 (N_12961,N_5739,N_5214);
nor U12962 (N_12962,N_7634,N_5072);
xor U12963 (N_12963,N_9275,N_8282);
nand U12964 (N_12964,N_7997,N_7582);
and U12965 (N_12965,N_9242,N_5300);
nor U12966 (N_12966,N_6115,N_6470);
nand U12967 (N_12967,N_7488,N_7542);
nand U12968 (N_12968,N_6722,N_8988);
or U12969 (N_12969,N_8219,N_9338);
or U12970 (N_12970,N_8480,N_8440);
or U12971 (N_12971,N_9746,N_6245);
xor U12972 (N_12972,N_6802,N_5483);
or U12973 (N_12973,N_6122,N_5051);
and U12974 (N_12974,N_5305,N_9383);
nand U12975 (N_12975,N_5109,N_9693);
or U12976 (N_12976,N_9028,N_6546);
and U12977 (N_12977,N_8652,N_9560);
and U12978 (N_12978,N_6718,N_8138);
or U12979 (N_12979,N_6657,N_8693);
and U12980 (N_12980,N_7496,N_5089);
nand U12981 (N_12981,N_7250,N_7675);
nand U12982 (N_12982,N_5428,N_5088);
nor U12983 (N_12983,N_8556,N_6254);
nand U12984 (N_12984,N_6670,N_7676);
xor U12985 (N_12985,N_5290,N_8659);
and U12986 (N_12986,N_7937,N_6709);
nor U12987 (N_12987,N_9416,N_8316);
nand U12988 (N_12988,N_5757,N_9800);
nand U12989 (N_12989,N_7687,N_5271);
or U12990 (N_12990,N_7971,N_9294);
nor U12991 (N_12991,N_8990,N_9919);
nor U12992 (N_12992,N_9521,N_8408);
xor U12993 (N_12993,N_7376,N_9062);
and U12994 (N_12994,N_6810,N_9880);
or U12995 (N_12995,N_8113,N_8873);
nor U12996 (N_12996,N_7246,N_5842);
nor U12997 (N_12997,N_7783,N_8578);
nor U12998 (N_12998,N_6800,N_7097);
or U12999 (N_12999,N_7165,N_7759);
or U13000 (N_13000,N_8465,N_9893);
nor U13001 (N_13001,N_6618,N_7745);
and U13002 (N_13002,N_5852,N_5783);
or U13003 (N_13003,N_9566,N_5632);
and U13004 (N_13004,N_5244,N_7603);
or U13005 (N_13005,N_6187,N_7503);
nand U13006 (N_13006,N_6199,N_6862);
or U13007 (N_13007,N_6398,N_8656);
xor U13008 (N_13008,N_7626,N_6905);
or U13009 (N_13009,N_9359,N_9332);
xor U13010 (N_13010,N_7442,N_8524);
xor U13011 (N_13011,N_6598,N_6079);
xor U13012 (N_13012,N_7704,N_9011);
and U13013 (N_13013,N_6044,N_7935);
nand U13014 (N_13014,N_9513,N_8306);
nor U13015 (N_13015,N_8139,N_6181);
nand U13016 (N_13016,N_6427,N_8355);
or U13017 (N_13017,N_9692,N_7416);
nor U13018 (N_13018,N_9316,N_9549);
or U13019 (N_13019,N_6960,N_9153);
and U13020 (N_13020,N_5868,N_8446);
or U13021 (N_13021,N_6988,N_9529);
and U13022 (N_13022,N_5378,N_8094);
or U13023 (N_13023,N_9513,N_7981);
nor U13024 (N_13024,N_8154,N_9583);
nand U13025 (N_13025,N_5739,N_8818);
and U13026 (N_13026,N_7073,N_7824);
xor U13027 (N_13027,N_8722,N_9648);
and U13028 (N_13028,N_7960,N_5164);
xor U13029 (N_13029,N_7858,N_9946);
or U13030 (N_13030,N_5876,N_8122);
nor U13031 (N_13031,N_7197,N_5414);
or U13032 (N_13032,N_6490,N_8722);
and U13033 (N_13033,N_7189,N_6828);
nor U13034 (N_13034,N_6939,N_5950);
and U13035 (N_13035,N_7712,N_8133);
xnor U13036 (N_13036,N_8600,N_5925);
nand U13037 (N_13037,N_6378,N_6896);
nand U13038 (N_13038,N_5557,N_6997);
or U13039 (N_13039,N_7955,N_9649);
nor U13040 (N_13040,N_7071,N_6785);
nor U13041 (N_13041,N_7673,N_9663);
nand U13042 (N_13042,N_5947,N_8605);
xnor U13043 (N_13043,N_7043,N_9636);
nor U13044 (N_13044,N_7929,N_5462);
or U13045 (N_13045,N_7195,N_5978);
and U13046 (N_13046,N_7968,N_8934);
nor U13047 (N_13047,N_6805,N_6715);
xor U13048 (N_13048,N_7841,N_7081);
nor U13049 (N_13049,N_9899,N_5629);
and U13050 (N_13050,N_8828,N_7910);
or U13051 (N_13051,N_9578,N_7027);
or U13052 (N_13052,N_5771,N_9070);
or U13053 (N_13053,N_6137,N_6642);
or U13054 (N_13054,N_7412,N_5390);
nand U13055 (N_13055,N_8416,N_6937);
or U13056 (N_13056,N_7036,N_9935);
or U13057 (N_13057,N_7733,N_6837);
xor U13058 (N_13058,N_8695,N_6776);
or U13059 (N_13059,N_9943,N_9921);
and U13060 (N_13060,N_7542,N_8332);
nand U13061 (N_13061,N_6379,N_6327);
nand U13062 (N_13062,N_9443,N_5905);
nor U13063 (N_13063,N_7699,N_7785);
and U13064 (N_13064,N_7930,N_5876);
xnor U13065 (N_13065,N_5014,N_5758);
xor U13066 (N_13066,N_9815,N_7144);
and U13067 (N_13067,N_6194,N_5657);
nor U13068 (N_13068,N_5348,N_5879);
nand U13069 (N_13069,N_7344,N_7534);
or U13070 (N_13070,N_8575,N_5344);
nor U13071 (N_13071,N_6061,N_8058);
or U13072 (N_13072,N_7649,N_8719);
xor U13073 (N_13073,N_6912,N_6294);
nor U13074 (N_13074,N_8630,N_6910);
nand U13075 (N_13075,N_9707,N_5298);
or U13076 (N_13076,N_7149,N_8202);
nor U13077 (N_13077,N_9717,N_5153);
or U13078 (N_13078,N_5833,N_6224);
nor U13079 (N_13079,N_5457,N_7446);
nor U13080 (N_13080,N_9245,N_6315);
nand U13081 (N_13081,N_7183,N_5786);
nand U13082 (N_13082,N_6344,N_9839);
and U13083 (N_13083,N_9803,N_6674);
nand U13084 (N_13084,N_9265,N_5834);
and U13085 (N_13085,N_7301,N_5692);
and U13086 (N_13086,N_7502,N_7755);
and U13087 (N_13087,N_5901,N_9807);
nor U13088 (N_13088,N_5238,N_7623);
xor U13089 (N_13089,N_5482,N_7773);
nor U13090 (N_13090,N_8706,N_9445);
xor U13091 (N_13091,N_6262,N_8203);
nor U13092 (N_13092,N_7911,N_9520);
nor U13093 (N_13093,N_7012,N_9152);
or U13094 (N_13094,N_9827,N_8656);
or U13095 (N_13095,N_7553,N_8450);
and U13096 (N_13096,N_6178,N_5699);
and U13097 (N_13097,N_6302,N_9918);
and U13098 (N_13098,N_5871,N_6535);
or U13099 (N_13099,N_6790,N_5647);
and U13100 (N_13100,N_6174,N_8329);
or U13101 (N_13101,N_7811,N_9328);
nand U13102 (N_13102,N_5023,N_5667);
nor U13103 (N_13103,N_6876,N_8910);
or U13104 (N_13104,N_6814,N_9381);
nand U13105 (N_13105,N_8785,N_7678);
and U13106 (N_13106,N_5202,N_9392);
nand U13107 (N_13107,N_9562,N_9049);
nand U13108 (N_13108,N_8678,N_6113);
and U13109 (N_13109,N_6778,N_6235);
or U13110 (N_13110,N_9186,N_5270);
xor U13111 (N_13111,N_9424,N_8308);
nand U13112 (N_13112,N_7241,N_5311);
and U13113 (N_13113,N_5948,N_5742);
xor U13114 (N_13114,N_6349,N_6882);
nor U13115 (N_13115,N_9430,N_5037);
xor U13116 (N_13116,N_6419,N_6370);
nand U13117 (N_13117,N_5229,N_5777);
nand U13118 (N_13118,N_8412,N_9152);
nor U13119 (N_13119,N_5229,N_6918);
nor U13120 (N_13120,N_5256,N_9082);
nand U13121 (N_13121,N_6435,N_5487);
and U13122 (N_13122,N_5406,N_7464);
xnor U13123 (N_13123,N_5283,N_8700);
nand U13124 (N_13124,N_8003,N_6489);
nor U13125 (N_13125,N_5334,N_9395);
nand U13126 (N_13126,N_7607,N_5147);
or U13127 (N_13127,N_7683,N_5594);
nor U13128 (N_13128,N_6009,N_6192);
and U13129 (N_13129,N_9590,N_5426);
nor U13130 (N_13130,N_9493,N_8995);
nand U13131 (N_13131,N_5433,N_5542);
and U13132 (N_13132,N_7588,N_8269);
nor U13133 (N_13133,N_9384,N_9113);
nand U13134 (N_13134,N_5909,N_6810);
and U13135 (N_13135,N_9902,N_8506);
nand U13136 (N_13136,N_5622,N_5058);
and U13137 (N_13137,N_9720,N_5761);
and U13138 (N_13138,N_7652,N_9162);
or U13139 (N_13139,N_7548,N_7054);
or U13140 (N_13140,N_6879,N_7157);
nor U13141 (N_13141,N_8272,N_8947);
nor U13142 (N_13142,N_7666,N_7751);
nand U13143 (N_13143,N_5558,N_7021);
nor U13144 (N_13144,N_7850,N_8981);
and U13145 (N_13145,N_7439,N_6744);
nand U13146 (N_13146,N_9512,N_7839);
nand U13147 (N_13147,N_5225,N_7135);
nand U13148 (N_13148,N_9605,N_7031);
nor U13149 (N_13149,N_9400,N_7083);
or U13150 (N_13150,N_8286,N_8949);
and U13151 (N_13151,N_8339,N_8419);
or U13152 (N_13152,N_8203,N_7372);
xor U13153 (N_13153,N_6721,N_9903);
or U13154 (N_13154,N_7894,N_8012);
nand U13155 (N_13155,N_7345,N_9452);
or U13156 (N_13156,N_9309,N_7334);
nand U13157 (N_13157,N_9545,N_9923);
xor U13158 (N_13158,N_6499,N_7071);
nand U13159 (N_13159,N_7126,N_8930);
xnor U13160 (N_13160,N_6776,N_6957);
nor U13161 (N_13161,N_9981,N_5398);
xnor U13162 (N_13162,N_6208,N_8289);
xnor U13163 (N_13163,N_7022,N_9603);
or U13164 (N_13164,N_5534,N_6600);
xor U13165 (N_13165,N_5389,N_8485);
and U13166 (N_13166,N_8011,N_6156);
and U13167 (N_13167,N_7508,N_5179);
nand U13168 (N_13168,N_8945,N_8600);
nand U13169 (N_13169,N_9427,N_7217);
nand U13170 (N_13170,N_8270,N_8036);
xnor U13171 (N_13171,N_7183,N_7382);
nor U13172 (N_13172,N_7149,N_8621);
and U13173 (N_13173,N_8452,N_9822);
nand U13174 (N_13174,N_8942,N_7154);
and U13175 (N_13175,N_6490,N_9679);
or U13176 (N_13176,N_9454,N_5556);
nand U13177 (N_13177,N_9971,N_7906);
nor U13178 (N_13178,N_5574,N_7811);
nor U13179 (N_13179,N_7133,N_7817);
nor U13180 (N_13180,N_6697,N_5274);
nor U13181 (N_13181,N_9329,N_5649);
and U13182 (N_13182,N_8119,N_8662);
nor U13183 (N_13183,N_8730,N_7424);
nand U13184 (N_13184,N_6172,N_6653);
or U13185 (N_13185,N_7425,N_7568);
or U13186 (N_13186,N_6312,N_6515);
nand U13187 (N_13187,N_7485,N_6799);
or U13188 (N_13188,N_8489,N_5147);
and U13189 (N_13189,N_5845,N_7898);
nand U13190 (N_13190,N_8993,N_9821);
or U13191 (N_13191,N_6317,N_7780);
xor U13192 (N_13192,N_7711,N_6119);
or U13193 (N_13193,N_8330,N_5352);
and U13194 (N_13194,N_9614,N_5304);
nand U13195 (N_13195,N_5606,N_5300);
or U13196 (N_13196,N_8512,N_6660);
and U13197 (N_13197,N_7200,N_6611);
nand U13198 (N_13198,N_9556,N_7853);
nand U13199 (N_13199,N_8695,N_7741);
or U13200 (N_13200,N_7568,N_7537);
nand U13201 (N_13201,N_6914,N_6080);
nand U13202 (N_13202,N_7128,N_5000);
xnor U13203 (N_13203,N_6040,N_9638);
or U13204 (N_13204,N_8337,N_9908);
nor U13205 (N_13205,N_7638,N_7489);
nand U13206 (N_13206,N_9796,N_6920);
xnor U13207 (N_13207,N_8044,N_5481);
or U13208 (N_13208,N_5716,N_6473);
or U13209 (N_13209,N_6114,N_6195);
xnor U13210 (N_13210,N_6794,N_5043);
or U13211 (N_13211,N_7523,N_7166);
nand U13212 (N_13212,N_7585,N_8650);
and U13213 (N_13213,N_9414,N_7044);
or U13214 (N_13214,N_5616,N_7308);
and U13215 (N_13215,N_8853,N_6955);
and U13216 (N_13216,N_7386,N_6116);
nor U13217 (N_13217,N_9742,N_7228);
nor U13218 (N_13218,N_7052,N_9858);
and U13219 (N_13219,N_9232,N_5866);
nand U13220 (N_13220,N_5545,N_7891);
and U13221 (N_13221,N_9149,N_7683);
and U13222 (N_13222,N_6250,N_9440);
or U13223 (N_13223,N_7475,N_8395);
xnor U13224 (N_13224,N_7060,N_7751);
nor U13225 (N_13225,N_7488,N_5996);
nor U13226 (N_13226,N_9086,N_6752);
or U13227 (N_13227,N_8241,N_8685);
and U13228 (N_13228,N_5724,N_7405);
and U13229 (N_13229,N_7154,N_9401);
and U13230 (N_13230,N_5382,N_6416);
or U13231 (N_13231,N_8332,N_5875);
nor U13232 (N_13232,N_8835,N_5789);
and U13233 (N_13233,N_6571,N_6187);
nor U13234 (N_13234,N_5479,N_9388);
and U13235 (N_13235,N_7498,N_8646);
or U13236 (N_13236,N_5258,N_9928);
xor U13237 (N_13237,N_8900,N_9693);
and U13238 (N_13238,N_7461,N_7109);
and U13239 (N_13239,N_6953,N_8203);
nand U13240 (N_13240,N_9034,N_7324);
or U13241 (N_13241,N_9152,N_8194);
and U13242 (N_13242,N_9068,N_7357);
xor U13243 (N_13243,N_9687,N_7612);
or U13244 (N_13244,N_7032,N_9522);
nand U13245 (N_13245,N_9931,N_6042);
or U13246 (N_13246,N_7336,N_7396);
nand U13247 (N_13247,N_6026,N_5489);
xnor U13248 (N_13248,N_5038,N_5800);
or U13249 (N_13249,N_6595,N_8715);
xor U13250 (N_13250,N_8400,N_5933);
nor U13251 (N_13251,N_8213,N_7383);
or U13252 (N_13252,N_9563,N_5451);
nand U13253 (N_13253,N_6478,N_6622);
nor U13254 (N_13254,N_5192,N_5371);
nor U13255 (N_13255,N_9409,N_6729);
nor U13256 (N_13256,N_6645,N_7289);
and U13257 (N_13257,N_6335,N_6480);
or U13258 (N_13258,N_5813,N_5067);
nand U13259 (N_13259,N_7136,N_5705);
or U13260 (N_13260,N_9418,N_9098);
nor U13261 (N_13261,N_7269,N_6913);
nand U13262 (N_13262,N_5259,N_6030);
nor U13263 (N_13263,N_6342,N_9940);
or U13264 (N_13264,N_5040,N_8122);
and U13265 (N_13265,N_5681,N_8056);
or U13266 (N_13266,N_7258,N_9599);
nand U13267 (N_13267,N_6853,N_9050);
nand U13268 (N_13268,N_7917,N_9690);
and U13269 (N_13269,N_6367,N_9588);
or U13270 (N_13270,N_6915,N_6327);
nor U13271 (N_13271,N_9370,N_7169);
nor U13272 (N_13272,N_6199,N_5570);
nand U13273 (N_13273,N_5582,N_6631);
nand U13274 (N_13274,N_7831,N_8005);
nand U13275 (N_13275,N_5225,N_7051);
and U13276 (N_13276,N_9516,N_5730);
nand U13277 (N_13277,N_8892,N_9276);
and U13278 (N_13278,N_9235,N_7718);
and U13279 (N_13279,N_7324,N_8540);
and U13280 (N_13280,N_6179,N_9219);
xor U13281 (N_13281,N_6691,N_7649);
and U13282 (N_13282,N_9280,N_6313);
and U13283 (N_13283,N_7429,N_5700);
or U13284 (N_13284,N_9982,N_5723);
nor U13285 (N_13285,N_6065,N_8430);
and U13286 (N_13286,N_9572,N_7012);
and U13287 (N_13287,N_6896,N_9746);
nand U13288 (N_13288,N_7288,N_8381);
nand U13289 (N_13289,N_7969,N_7627);
and U13290 (N_13290,N_9715,N_9331);
or U13291 (N_13291,N_6822,N_8569);
and U13292 (N_13292,N_8346,N_8050);
and U13293 (N_13293,N_9145,N_9652);
or U13294 (N_13294,N_6411,N_8737);
xnor U13295 (N_13295,N_6413,N_9615);
or U13296 (N_13296,N_8367,N_5296);
xor U13297 (N_13297,N_6840,N_6891);
or U13298 (N_13298,N_5628,N_8313);
nand U13299 (N_13299,N_8241,N_5425);
nand U13300 (N_13300,N_9173,N_9545);
nand U13301 (N_13301,N_9687,N_5110);
and U13302 (N_13302,N_8368,N_7805);
xnor U13303 (N_13303,N_8876,N_6036);
nor U13304 (N_13304,N_5216,N_5391);
and U13305 (N_13305,N_9093,N_9955);
xnor U13306 (N_13306,N_7565,N_7456);
nor U13307 (N_13307,N_7600,N_5748);
or U13308 (N_13308,N_8128,N_9577);
xnor U13309 (N_13309,N_6904,N_6460);
nor U13310 (N_13310,N_6910,N_6005);
nor U13311 (N_13311,N_8774,N_9603);
nand U13312 (N_13312,N_7017,N_6666);
nor U13313 (N_13313,N_9410,N_5250);
and U13314 (N_13314,N_8021,N_8318);
or U13315 (N_13315,N_9501,N_9470);
nand U13316 (N_13316,N_9826,N_8447);
nor U13317 (N_13317,N_9614,N_5216);
or U13318 (N_13318,N_9881,N_9183);
nor U13319 (N_13319,N_5775,N_6601);
nand U13320 (N_13320,N_5122,N_8669);
and U13321 (N_13321,N_9421,N_7732);
or U13322 (N_13322,N_8829,N_7687);
nor U13323 (N_13323,N_8835,N_6597);
and U13324 (N_13324,N_9564,N_5403);
or U13325 (N_13325,N_8549,N_7584);
nor U13326 (N_13326,N_8080,N_9329);
and U13327 (N_13327,N_6353,N_5497);
nand U13328 (N_13328,N_7307,N_5687);
and U13329 (N_13329,N_7396,N_8272);
nor U13330 (N_13330,N_9849,N_6852);
xnor U13331 (N_13331,N_6287,N_7624);
nor U13332 (N_13332,N_5391,N_9715);
or U13333 (N_13333,N_5774,N_8229);
or U13334 (N_13334,N_5282,N_9394);
xor U13335 (N_13335,N_5959,N_7410);
nor U13336 (N_13336,N_8058,N_7707);
and U13337 (N_13337,N_7352,N_9650);
and U13338 (N_13338,N_8281,N_9020);
nand U13339 (N_13339,N_5904,N_6836);
nand U13340 (N_13340,N_9596,N_8210);
and U13341 (N_13341,N_7866,N_7290);
nand U13342 (N_13342,N_9612,N_6417);
xnor U13343 (N_13343,N_8501,N_8320);
nand U13344 (N_13344,N_8676,N_9729);
nor U13345 (N_13345,N_6759,N_8400);
nor U13346 (N_13346,N_5199,N_5661);
and U13347 (N_13347,N_8680,N_5652);
and U13348 (N_13348,N_7188,N_9947);
and U13349 (N_13349,N_6081,N_8021);
nor U13350 (N_13350,N_7836,N_7285);
or U13351 (N_13351,N_8556,N_8348);
or U13352 (N_13352,N_6779,N_8554);
or U13353 (N_13353,N_5111,N_5369);
and U13354 (N_13354,N_8361,N_8992);
nor U13355 (N_13355,N_5055,N_9276);
or U13356 (N_13356,N_9118,N_6601);
nor U13357 (N_13357,N_6407,N_5077);
nand U13358 (N_13358,N_8341,N_5338);
or U13359 (N_13359,N_5889,N_5190);
nand U13360 (N_13360,N_7597,N_8600);
nor U13361 (N_13361,N_9775,N_8435);
and U13362 (N_13362,N_7311,N_6660);
and U13363 (N_13363,N_7566,N_9176);
xor U13364 (N_13364,N_8629,N_7063);
or U13365 (N_13365,N_6086,N_6604);
nand U13366 (N_13366,N_6681,N_5485);
xnor U13367 (N_13367,N_9632,N_7882);
or U13368 (N_13368,N_6630,N_8009);
or U13369 (N_13369,N_9683,N_7934);
or U13370 (N_13370,N_5296,N_5727);
and U13371 (N_13371,N_8156,N_5773);
nand U13372 (N_13372,N_6125,N_5653);
nand U13373 (N_13373,N_6136,N_8885);
nand U13374 (N_13374,N_6533,N_7063);
and U13375 (N_13375,N_9094,N_5426);
nand U13376 (N_13376,N_9502,N_6052);
or U13377 (N_13377,N_5209,N_5771);
or U13378 (N_13378,N_5178,N_5056);
or U13379 (N_13379,N_7529,N_7251);
xnor U13380 (N_13380,N_9232,N_6097);
nor U13381 (N_13381,N_7001,N_8608);
nand U13382 (N_13382,N_7947,N_6616);
or U13383 (N_13383,N_6562,N_5737);
and U13384 (N_13384,N_6508,N_9535);
nand U13385 (N_13385,N_7918,N_8016);
nand U13386 (N_13386,N_5831,N_9491);
or U13387 (N_13387,N_7238,N_8980);
nor U13388 (N_13388,N_9217,N_9320);
nor U13389 (N_13389,N_9430,N_7369);
xor U13390 (N_13390,N_8604,N_7494);
nor U13391 (N_13391,N_5507,N_6651);
nand U13392 (N_13392,N_6599,N_6225);
and U13393 (N_13393,N_7456,N_9666);
or U13394 (N_13394,N_8067,N_9335);
nand U13395 (N_13395,N_9197,N_9890);
nor U13396 (N_13396,N_8593,N_6665);
or U13397 (N_13397,N_8198,N_8605);
xor U13398 (N_13398,N_9550,N_7772);
or U13399 (N_13399,N_9451,N_7884);
or U13400 (N_13400,N_9049,N_8919);
or U13401 (N_13401,N_8394,N_6538);
and U13402 (N_13402,N_9584,N_8149);
or U13403 (N_13403,N_6310,N_7178);
nor U13404 (N_13404,N_5996,N_6002);
nor U13405 (N_13405,N_7303,N_6027);
nor U13406 (N_13406,N_7374,N_6097);
xnor U13407 (N_13407,N_8628,N_8946);
nand U13408 (N_13408,N_7448,N_7896);
nor U13409 (N_13409,N_8815,N_6757);
nand U13410 (N_13410,N_9545,N_7229);
nor U13411 (N_13411,N_9468,N_5928);
nor U13412 (N_13412,N_8574,N_5581);
xor U13413 (N_13413,N_9679,N_8638);
or U13414 (N_13414,N_9062,N_9757);
or U13415 (N_13415,N_5480,N_7537);
and U13416 (N_13416,N_7669,N_6346);
nor U13417 (N_13417,N_8861,N_5346);
or U13418 (N_13418,N_7737,N_7975);
or U13419 (N_13419,N_8749,N_5332);
nor U13420 (N_13420,N_7903,N_9104);
nor U13421 (N_13421,N_9258,N_8530);
or U13422 (N_13422,N_7387,N_5210);
or U13423 (N_13423,N_5189,N_6803);
nand U13424 (N_13424,N_8214,N_7078);
and U13425 (N_13425,N_8733,N_6336);
and U13426 (N_13426,N_7301,N_6228);
xor U13427 (N_13427,N_7609,N_9979);
nand U13428 (N_13428,N_5857,N_5568);
nor U13429 (N_13429,N_7792,N_7973);
and U13430 (N_13430,N_6148,N_8637);
nand U13431 (N_13431,N_8805,N_9105);
and U13432 (N_13432,N_5702,N_7884);
and U13433 (N_13433,N_8580,N_6250);
nand U13434 (N_13434,N_7232,N_6484);
and U13435 (N_13435,N_5069,N_6206);
nor U13436 (N_13436,N_6177,N_6610);
nand U13437 (N_13437,N_7454,N_8954);
and U13438 (N_13438,N_8385,N_9734);
nor U13439 (N_13439,N_8076,N_7636);
and U13440 (N_13440,N_8815,N_7210);
nand U13441 (N_13441,N_8366,N_5598);
and U13442 (N_13442,N_8837,N_9189);
or U13443 (N_13443,N_6005,N_6107);
nor U13444 (N_13444,N_8653,N_5175);
nand U13445 (N_13445,N_7835,N_6225);
or U13446 (N_13446,N_6849,N_6206);
nand U13447 (N_13447,N_7431,N_5044);
and U13448 (N_13448,N_9533,N_9809);
xnor U13449 (N_13449,N_7099,N_9703);
xor U13450 (N_13450,N_8013,N_9677);
xnor U13451 (N_13451,N_5992,N_5223);
xor U13452 (N_13452,N_6551,N_6427);
or U13453 (N_13453,N_8482,N_5844);
and U13454 (N_13454,N_9219,N_6457);
nor U13455 (N_13455,N_6657,N_9295);
nor U13456 (N_13456,N_8538,N_8348);
and U13457 (N_13457,N_5532,N_7287);
xnor U13458 (N_13458,N_8984,N_9111);
or U13459 (N_13459,N_6108,N_6465);
nor U13460 (N_13460,N_8491,N_7640);
nor U13461 (N_13461,N_7895,N_8306);
xor U13462 (N_13462,N_9132,N_7011);
and U13463 (N_13463,N_8857,N_8896);
or U13464 (N_13464,N_6196,N_6083);
nor U13465 (N_13465,N_8074,N_5887);
nor U13466 (N_13466,N_9997,N_9020);
or U13467 (N_13467,N_6436,N_6561);
nor U13468 (N_13468,N_6379,N_5299);
and U13469 (N_13469,N_9238,N_8314);
nand U13470 (N_13470,N_6082,N_6262);
and U13471 (N_13471,N_7056,N_5396);
or U13472 (N_13472,N_5086,N_9401);
nand U13473 (N_13473,N_9679,N_9166);
and U13474 (N_13474,N_8820,N_6571);
nor U13475 (N_13475,N_5655,N_9558);
and U13476 (N_13476,N_9768,N_6732);
and U13477 (N_13477,N_6260,N_7004);
or U13478 (N_13478,N_5783,N_8083);
or U13479 (N_13479,N_7462,N_6218);
or U13480 (N_13480,N_7968,N_8249);
nor U13481 (N_13481,N_8455,N_8608);
or U13482 (N_13482,N_6095,N_8770);
or U13483 (N_13483,N_6811,N_6658);
or U13484 (N_13484,N_7266,N_9208);
and U13485 (N_13485,N_6030,N_8497);
or U13486 (N_13486,N_6919,N_7466);
or U13487 (N_13487,N_8590,N_9501);
and U13488 (N_13488,N_5749,N_5380);
nor U13489 (N_13489,N_7851,N_6544);
and U13490 (N_13490,N_5130,N_5853);
nand U13491 (N_13491,N_6463,N_9038);
or U13492 (N_13492,N_5019,N_7617);
nand U13493 (N_13493,N_7075,N_9493);
nor U13494 (N_13494,N_6177,N_8622);
nand U13495 (N_13495,N_6521,N_9718);
nor U13496 (N_13496,N_6986,N_9041);
nand U13497 (N_13497,N_9776,N_7394);
nand U13498 (N_13498,N_8651,N_8604);
nor U13499 (N_13499,N_5418,N_7062);
or U13500 (N_13500,N_7613,N_5734);
nor U13501 (N_13501,N_7527,N_9899);
xnor U13502 (N_13502,N_6109,N_9629);
and U13503 (N_13503,N_5308,N_8931);
nor U13504 (N_13504,N_5233,N_9040);
xor U13505 (N_13505,N_7143,N_7368);
or U13506 (N_13506,N_9212,N_5695);
nor U13507 (N_13507,N_8845,N_8267);
nand U13508 (N_13508,N_9177,N_6954);
nor U13509 (N_13509,N_7272,N_5802);
and U13510 (N_13510,N_5894,N_8649);
nand U13511 (N_13511,N_8375,N_5624);
nand U13512 (N_13512,N_6836,N_5963);
nand U13513 (N_13513,N_9085,N_7405);
xor U13514 (N_13514,N_5899,N_8731);
and U13515 (N_13515,N_5379,N_7703);
or U13516 (N_13516,N_6196,N_6158);
or U13517 (N_13517,N_9836,N_8315);
and U13518 (N_13518,N_9686,N_8080);
nand U13519 (N_13519,N_6654,N_7577);
or U13520 (N_13520,N_8094,N_5657);
or U13521 (N_13521,N_9183,N_5963);
or U13522 (N_13522,N_5042,N_6950);
and U13523 (N_13523,N_9842,N_8762);
or U13524 (N_13524,N_5476,N_9004);
nand U13525 (N_13525,N_5881,N_7741);
nor U13526 (N_13526,N_7009,N_8882);
and U13527 (N_13527,N_7305,N_9560);
or U13528 (N_13528,N_9010,N_7977);
nand U13529 (N_13529,N_7039,N_5908);
or U13530 (N_13530,N_5689,N_7410);
nor U13531 (N_13531,N_5161,N_6385);
nor U13532 (N_13532,N_9330,N_8619);
nor U13533 (N_13533,N_6240,N_8978);
nand U13534 (N_13534,N_8451,N_5945);
nor U13535 (N_13535,N_5366,N_5308);
nand U13536 (N_13536,N_5113,N_9115);
and U13537 (N_13537,N_7137,N_5474);
or U13538 (N_13538,N_9275,N_7234);
or U13539 (N_13539,N_5041,N_7569);
nor U13540 (N_13540,N_7510,N_8179);
nand U13541 (N_13541,N_5892,N_6920);
and U13542 (N_13542,N_7611,N_7357);
nand U13543 (N_13543,N_7802,N_7793);
xor U13544 (N_13544,N_7499,N_5734);
nand U13545 (N_13545,N_5064,N_5990);
nand U13546 (N_13546,N_5787,N_6013);
nand U13547 (N_13547,N_5973,N_9955);
nor U13548 (N_13548,N_7851,N_7254);
or U13549 (N_13549,N_7975,N_9078);
nand U13550 (N_13550,N_6902,N_9225);
nand U13551 (N_13551,N_8456,N_8826);
or U13552 (N_13552,N_7083,N_8847);
nor U13553 (N_13553,N_7300,N_9759);
or U13554 (N_13554,N_5203,N_8118);
xor U13555 (N_13555,N_9193,N_9593);
or U13556 (N_13556,N_6915,N_8300);
and U13557 (N_13557,N_5121,N_7647);
nand U13558 (N_13558,N_7783,N_9456);
and U13559 (N_13559,N_5103,N_7523);
or U13560 (N_13560,N_7670,N_8191);
nor U13561 (N_13561,N_6816,N_8377);
nor U13562 (N_13562,N_5411,N_5574);
nor U13563 (N_13563,N_6140,N_7667);
nand U13564 (N_13564,N_5635,N_5334);
or U13565 (N_13565,N_9948,N_9675);
and U13566 (N_13566,N_5589,N_5909);
xor U13567 (N_13567,N_8619,N_5572);
nor U13568 (N_13568,N_9379,N_5045);
nor U13569 (N_13569,N_7965,N_8788);
nor U13570 (N_13570,N_5970,N_5563);
and U13571 (N_13571,N_6188,N_5072);
and U13572 (N_13572,N_9732,N_6400);
or U13573 (N_13573,N_7382,N_7489);
nor U13574 (N_13574,N_7140,N_5479);
or U13575 (N_13575,N_5976,N_6320);
nor U13576 (N_13576,N_6764,N_9632);
and U13577 (N_13577,N_7026,N_7849);
nor U13578 (N_13578,N_5194,N_8783);
nand U13579 (N_13579,N_6198,N_5376);
or U13580 (N_13580,N_9212,N_8303);
nor U13581 (N_13581,N_7905,N_7259);
nor U13582 (N_13582,N_9995,N_7457);
and U13583 (N_13583,N_9541,N_5616);
nor U13584 (N_13584,N_7500,N_8864);
or U13585 (N_13585,N_5526,N_6864);
or U13586 (N_13586,N_8535,N_6011);
nor U13587 (N_13587,N_5815,N_8429);
and U13588 (N_13588,N_9337,N_8445);
nand U13589 (N_13589,N_7514,N_8011);
nand U13590 (N_13590,N_8732,N_8284);
nand U13591 (N_13591,N_9324,N_8574);
nand U13592 (N_13592,N_5547,N_7130);
nor U13593 (N_13593,N_5262,N_7417);
nand U13594 (N_13594,N_7341,N_8512);
nor U13595 (N_13595,N_9768,N_7848);
nand U13596 (N_13596,N_6719,N_5835);
nor U13597 (N_13597,N_6903,N_6196);
or U13598 (N_13598,N_5284,N_5573);
xnor U13599 (N_13599,N_7018,N_9379);
and U13600 (N_13600,N_6422,N_9444);
nor U13601 (N_13601,N_5644,N_6522);
nand U13602 (N_13602,N_7329,N_5780);
xnor U13603 (N_13603,N_6174,N_6273);
nor U13604 (N_13604,N_7112,N_8732);
nor U13605 (N_13605,N_5179,N_6540);
xnor U13606 (N_13606,N_5726,N_7095);
or U13607 (N_13607,N_9197,N_6013);
or U13608 (N_13608,N_9743,N_8745);
nand U13609 (N_13609,N_7123,N_9239);
or U13610 (N_13610,N_8142,N_8202);
and U13611 (N_13611,N_5452,N_6197);
nor U13612 (N_13612,N_5944,N_9253);
nor U13613 (N_13613,N_8441,N_9820);
nor U13614 (N_13614,N_6450,N_6987);
or U13615 (N_13615,N_7890,N_8384);
xnor U13616 (N_13616,N_8691,N_7026);
or U13617 (N_13617,N_5637,N_9852);
nor U13618 (N_13618,N_8478,N_9445);
nand U13619 (N_13619,N_7120,N_9718);
or U13620 (N_13620,N_9527,N_9154);
nor U13621 (N_13621,N_8013,N_5181);
and U13622 (N_13622,N_5700,N_9917);
nor U13623 (N_13623,N_7921,N_6245);
or U13624 (N_13624,N_8105,N_8665);
nor U13625 (N_13625,N_7949,N_7719);
nor U13626 (N_13626,N_8770,N_6325);
xnor U13627 (N_13627,N_6840,N_8041);
or U13628 (N_13628,N_9761,N_5564);
and U13629 (N_13629,N_8115,N_5419);
and U13630 (N_13630,N_8475,N_5749);
nor U13631 (N_13631,N_9799,N_5802);
and U13632 (N_13632,N_5683,N_8852);
or U13633 (N_13633,N_9553,N_7440);
and U13634 (N_13634,N_5005,N_7127);
and U13635 (N_13635,N_8663,N_8038);
or U13636 (N_13636,N_9694,N_7641);
and U13637 (N_13637,N_8218,N_7481);
or U13638 (N_13638,N_5486,N_8654);
nand U13639 (N_13639,N_7559,N_8254);
and U13640 (N_13640,N_8585,N_6218);
and U13641 (N_13641,N_5699,N_8071);
and U13642 (N_13642,N_6138,N_5099);
xnor U13643 (N_13643,N_5896,N_8575);
or U13644 (N_13644,N_6122,N_6178);
and U13645 (N_13645,N_9931,N_8989);
nand U13646 (N_13646,N_5131,N_8736);
nor U13647 (N_13647,N_8497,N_5200);
and U13648 (N_13648,N_9768,N_9191);
and U13649 (N_13649,N_9719,N_6166);
nor U13650 (N_13650,N_8011,N_5213);
and U13651 (N_13651,N_5888,N_6234);
nor U13652 (N_13652,N_6061,N_7018);
and U13653 (N_13653,N_8207,N_5893);
nand U13654 (N_13654,N_9143,N_9158);
or U13655 (N_13655,N_6808,N_9751);
nor U13656 (N_13656,N_9164,N_9116);
or U13657 (N_13657,N_5165,N_9124);
nand U13658 (N_13658,N_7549,N_8054);
or U13659 (N_13659,N_9325,N_6351);
and U13660 (N_13660,N_8071,N_7484);
xnor U13661 (N_13661,N_9385,N_6737);
and U13662 (N_13662,N_9129,N_6927);
or U13663 (N_13663,N_7847,N_5012);
nand U13664 (N_13664,N_7626,N_9832);
and U13665 (N_13665,N_7460,N_5068);
nor U13666 (N_13666,N_6356,N_5381);
and U13667 (N_13667,N_5374,N_6999);
or U13668 (N_13668,N_5990,N_5633);
and U13669 (N_13669,N_5092,N_8348);
nor U13670 (N_13670,N_5105,N_7603);
or U13671 (N_13671,N_5541,N_8136);
nor U13672 (N_13672,N_7521,N_7894);
nor U13673 (N_13673,N_9030,N_9406);
nor U13674 (N_13674,N_9493,N_8665);
or U13675 (N_13675,N_6723,N_8260);
xor U13676 (N_13676,N_9264,N_6701);
and U13677 (N_13677,N_5760,N_8584);
or U13678 (N_13678,N_6395,N_9699);
xor U13679 (N_13679,N_9418,N_8550);
nor U13680 (N_13680,N_5568,N_8751);
or U13681 (N_13681,N_5896,N_6361);
nor U13682 (N_13682,N_5912,N_9441);
and U13683 (N_13683,N_9758,N_6304);
nor U13684 (N_13684,N_5918,N_6405);
or U13685 (N_13685,N_6189,N_9891);
nand U13686 (N_13686,N_5171,N_9030);
or U13687 (N_13687,N_5492,N_8453);
and U13688 (N_13688,N_5758,N_9819);
or U13689 (N_13689,N_7411,N_7172);
and U13690 (N_13690,N_8050,N_8429);
and U13691 (N_13691,N_8202,N_5885);
or U13692 (N_13692,N_5753,N_8168);
or U13693 (N_13693,N_8706,N_5433);
or U13694 (N_13694,N_6879,N_7507);
nand U13695 (N_13695,N_8335,N_8138);
and U13696 (N_13696,N_8944,N_8083);
nor U13697 (N_13697,N_9943,N_5927);
or U13698 (N_13698,N_7105,N_8640);
xnor U13699 (N_13699,N_9359,N_6525);
xnor U13700 (N_13700,N_6853,N_7336);
nand U13701 (N_13701,N_8883,N_8151);
or U13702 (N_13702,N_7557,N_9858);
xor U13703 (N_13703,N_8562,N_8760);
and U13704 (N_13704,N_7717,N_8112);
nand U13705 (N_13705,N_5728,N_5646);
nor U13706 (N_13706,N_7126,N_7218);
nor U13707 (N_13707,N_9896,N_7804);
or U13708 (N_13708,N_8320,N_6842);
and U13709 (N_13709,N_8417,N_8978);
xor U13710 (N_13710,N_7000,N_5356);
or U13711 (N_13711,N_6119,N_9987);
or U13712 (N_13712,N_9261,N_9422);
or U13713 (N_13713,N_7461,N_9966);
nor U13714 (N_13714,N_6451,N_7356);
and U13715 (N_13715,N_6511,N_7994);
xor U13716 (N_13716,N_7652,N_9994);
and U13717 (N_13717,N_7634,N_7694);
nand U13718 (N_13718,N_5859,N_7488);
nand U13719 (N_13719,N_5308,N_6139);
xnor U13720 (N_13720,N_7093,N_6185);
and U13721 (N_13721,N_5137,N_7246);
or U13722 (N_13722,N_9485,N_5582);
nor U13723 (N_13723,N_7276,N_9189);
nand U13724 (N_13724,N_5700,N_6408);
and U13725 (N_13725,N_7311,N_5961);
nor U13726 (N_13726,N_8750,N_8208);
and U13727 (N_13727,N_8924,N_5262);
nand U13728 (N_13728,N_8205,N_7860);
nand U13729 (N_13729,N_8260,N_5256);
or U13730 (N_13730,N_9013,N_6118);
nand U13731 (N_13731,N_7331,N_5176);
xor U13732 (N_13732,N_6587,N_6057);
nor U13733 (N_13733,N_5395,N_7161);
and U13734 (N_13734,N_5436,N_5973);
nor U13735 (N_13735,N_6984,N_7847);
and U13736 (N_13736,N_9492,N_6568);
or U13737 (N_13737,N_8308,N_8554);
or U13738 (N_13738,N_7138,N_5760);
nor U13739 (N_13739,N_7136,N_5431);
nand U13740 (N_13740,N_6191,N_7175);
nor U13741 (N_13741,N_6259,N_5288);
and U13742 (N_13742,N_8762,N_6841);
nand U13743 (N_13743,N_5847,N_8208);
and U13744 (N_13744,N_8900,N_6626);
and U13745 (N_13745,N_5637,N_8002);
or U13746 (N_13746,N_5178,N_6899);
nand U13747 (N_13747,N_5254,N_6048);
and U13748 (N_13748,N_6686,N_6165);
and U13749 (N_13749,N_5271,N_5739);
nand U13750 (N_13750,N_6920,N_7913);
and U13751 (N_13751,N_7129,N_5365);
xnor U13752 (N_13752,N_8788,N_8768);
and U13753 (N_13753,N_7405,N_5898);
and U13754 (N_13754,N_9934,N_5680);
xnor U13755 (N_13755,N_8784,N_9476);
nand U13756 (N_13756,N_5469,N_8030);
or U13757 (N_13757,N_8322,N_6590);
xor U13758 (N_13758,N_7415,N_8808);
or U13759 (N_13759,N_5255,N_9237);
nor U13760 (N_13760,N_9438,N_6136);
or U13761 (N_13761,N_6794,N_8254);
or U13762 (N_13762,N_8991,N_9774);
and U13763 (N_13763,N_6998,N_8990);
nand U13764 (N_13764,N_6275,N_5871);
nand U13765 (N_13765,N_9218,N_9629);
or U13766 (N_13766,N_8432,N_7597);
and U13767 (N_13767,N_6094,N_9154);
nand U13768 (N_13768,N_6939,N_8450);
nand U13769 (N_13769,N_6511,N_5065);
or U13770 (N_13770,N_5883,N_9073);
nand U13771 (N_13771,N_7970,N_8844);
nor U13772 (N_13772,N_6922,N_5492);
or U13773 (N_13773,N_5976,N_7223);
xnor U13774 (N_13774,N_8640,N_5359);
and U13775 (N_13775,N_6672,N_7084);
or U13776 (N_13776,N_5957,N_9807);
or U13777 (N_13777,N_8062,N_7854);
nor U13778 (N_13778,N_8619,N_9235);
nor U13779 (N_13779,N_8797,N_7131);
and U13780 (N_13780,N_7820,N_6075);
and U13781 (N_13781,N_7830,N_6710);
nand U13782 (N_13782,N_9198,N_9580);
and U13783 (N_13783,N_5860,N_7992);
or U13784 (N_13784,N_5682,N_9079);
nor U13785 (N_13785,N_9457,N_5639);
nand U13786 (N_13786,N_6101,N_8158);
and U13787 (N_13787,N_9240,N_6861);
nand U13788 (N_13788,N_7709,N_6853);
and U13789 (N_13789,N_5377,N_7858);
or U13790 (N_13790,N_9313,N_6280);
and U13791 (N_13791,N_6888,N_9513);
and U13792 (N_13792,N_5447,N_8831);
nor U13793 (N_13793,N_7518,N_8095);
and U13794 (N_13794,N_8987,N_7695);
and U13795 (N_13795,N_6086,N_5968);
and U13796 (N_13796,N_7217,N_7018);
nand U13797 (N_13797,N_7536,N_8755);
xor U13798 (N_13798,N_5450,N_8769);
and U13799 (N_13799,N_7248,N_8132);
and U13800 (N_13800,N_6384,N_6629);
nand U13801 (N_13801,N_8886,N_7859);
or U13802 (N_13802,N_6058,N_8264);
xor U13803 (N_13803,N_9845,N_5786);
and U13804 (N_13804,N_8088,N_5902);
nand U13805 (N_13805,N_9808,N_6998);
or U13806 (N_13806,N_5042,N_6996);
nand U13807 (N_13807,N_7140,N_5115);
and U13808 (N_13808,N_8884,N_9401);
nor U13809 (N_13809,N_9663,N_5295);
or U13810 (N_13810,N_8937,N_9171);
nor U13811 (N_13811,N_7362,N_8583);
xor U13812 (N_13812,N_9453,N_8225);
nand U13813 (N_13813,N_5319,N_8495);
nor U13814 (N_13814,N_5784,N_9130);
and U13815 (N_13815,N_8350,N_7636);
or U13816 (N_13816,N_6455,N_8204);
or U13817 (N_13817,N_8812,N_5671);
or U13818 (N_13818,N_7368,N_5473);
or U13819 (N_13819,N_6612,N_9412);
nor U13820 (N_13820,N_8354,N_9127);
or U13821 (N_13821,N_9772,N_5644);
and U13822 (N_13822,N_5637,N_9150);
nand U13823 (N_13823,N_6990,N_9554);
and U13824 (N_13824,N_5618,N_5317);
or U13825 (N_13825,N_5479,N_5667);
and U13826 (N_13826,N_8375,N_7117);
or U13827 (N_13827,N_8490,N_5479);
and U13828 (N_13828,N_6301,N_8225);
nand U13829 (N_13829,N_8169,N_5813);
nor U13830 (N_13830,N_6709,N_5029);
nand U13831 (N_13831,N_5810,N_8091);
and U13832 (N_13832,N_8130,N_7624);
nand U13833 (N_13833,N_8338,N_8384);
and U13834 (N_13834,N_7380,N_6270);
xnor U13835 (N_13835,N_8906,N_6040);
and U13836 (N_13836,N_8126,N_7944);
nor U13837 (N_13837,N_9251,N_9889);
or U13838 (N_13838,N_5855,N_9824);
nor U13839 (N_13839,N_5617,N_7510);
nand U13840 (N_13840,N_5776,N_9531);
nand U13841 (N_13841,N_5170,N_8581);
or U13842 (N_13842,N_8295,N_6701);
and U13843 (N_13843,N_7368,N_8530);
or U13844 (N_13844,N_6682,N_7460);
or U13845 (N_13845,N_7371,N_6925);
and U13846 (N_13846,N_7816,N_8391);
or U13847 (N_13847,N_5404,N_5463);
xnor U13848 (N_13848,N_6276,N_6253);
nand U13849 (N_13849,N_8103,N_8203);
or U13850 (N_13850,N_8691,N_6712);
and U13851 (N_13851,N_7497,N_9382);
or U13852 (N_13852,N_5596,N_7425);
nand U13853 (N_13853,N_9630,N_9572);
or U13854 (N_13854,N_8420,N_8922);
xor U13855 (N_13855,N_8016,N_5583);
nand U13856 (N_13856,N_9367,N_6177);
or U13857 (N_13857,N_5094,N_6402);
or U13858 (N_13858,N_8120,N_8625);
nand U13859 (N_13859,N_5235,N_5452);
nor U13860 (N_13860,N_7912,N_6544);
xor U13861 (N_13861,N_5295,N_8024);
nand U13862 (N_13862,N_9848,N_8592);
nor U13863 (N_13863,N_9357,N_8486);
nor U13864 (N_13864,N_8118,N_9633);
or U13865 (N_13865,N_6146,N_5646);
nor U13866 (N_13866,N_6448,N_5835);
or U13867 (N_13867,N_9374,N_6682);
or U13868 (N_13868,N_5325,N_6510);
nor U13869 (N_13869,N_5612,N_7873);
xor U13870 (N_13870,N_9368,N_5125);
or U13871 (N_13871,N_5034,N_7684);
and U13872 (N_13872,N_7519,N_9498);
nand U13873 (N_13873,N_7923,N_9838);
nand U13874 (N_13874,N_6922,N_6300);
or U13875 (N_13875,N_6562,N_7808);
nor U13876 (N_13876,N_5019,N_5259);
nor U13877 (N_13877,N_6983,N_5725);
nand U13878 (N_13878,N_6751,N_9790);
nand U13879 (N_13879,N_6480,N_5415);
or U13880 (N_13880,N_5016,N_5913);
or U13881 (N_13881,N_7313,N_7099);
nand U13882 (N_13882,N_5344,N_6382);
nor U13883 (N_13883,N_5483,N_6796);
xor U13884 (N_13884,N_6778,N_9316);
or U13885 (N_13885,N_8997,N_9633);
and U13886 (N_13886,N_7832,N_9188);
or U13887 (N_13887,N_6266,N_6667);
or U13888 (N_13888,N_8741,N_9280);
nand U13889 (N_13889,N_9063,N_7414);
and U13890 (N_13890,N_9027,N_8461);
and U13891 (N_13891,N_8109,N_8698);
nor U13892 (N_13892,N_6000,N_5185);
or U13893 (N_13893,N_7291,N_9922);
nor U13894 (N_13894,N_6274,N_9010);
and U13895 (N_13895,N_9429,N_8318);
or U13896 (N_13896,N_9157,N_8336);
nand U13897 (N_13897,N_9537,N_7670);
or U13898 (N_13898,N_6875,N_6589);
xnor U13899 (N_13899,N_6644,N_8936);
or U13900 (N_13900,N_6023,N_7005);
nand U13901 (N_13901,N_7819,N_7148);
nand U13902 (N_13902,N_6058,N_9878);
and U13903 (N_13903,N_8853,N_8307);
xnor U13904 (N_13904,N_9223,N_5770);
and U13905 (N_13905,N_8826,N_8226);
xor U13906 (N_13906,N_8694,N_6954);
or U13907 (N_13907,N_8202,N_7459);
and U13908 (N_13908,N_6617,N_6892);
nor U13909 (N_13909,N_7879,N_7585);
nor U13910 (N_13910,N_8962,N_5652);
or U13911 (N_13911,N_6447,N_6992);
and U13912 (N_13912,N_5796,N_8319);
and U13913 (N_13913,N_8752,N_5827);
nand U13914 (N_13914,N_9445,N_5350);
and U13915 (N_13915,N_6997,N_7113);
nand U13916 (N_13916,N_5734,N_9172);
nand U13917 (N_13917,N_6976,N_6753);
or U13918 (N_13918,N_7737,N_5033);
nor U13919 (N_13919,N_9550,N_9000);
or U13920 (N_13920,N_7411,N_5389);
or U13921 (N_13921,N_8130,N_6571);
or U13922 (N_13922,N_9971,N_9171);
nand U13923 (N_13923,N_6141,N_7257);
or U13924 (N_13924,N_7121,N_7998);
nand U13925 (N_13925,N_8686,N_9230);
or U13926 (N_13926,N_8977,N_9156);
or U13927 (N_13927,N_5851,N_5022);
and U13928 (N_13928,N_9537,N_8127);
nand U13929 (N_13929,N_6938,N_5580);
nand U13930 (N_13930,N_8642,N_9916);
and U13931 (N_13931,N_9910,N_8794);
xnor U13932 (N_13932,N_9481,N_5012);
and U13933 (N_13933,N_9940,N_5453);
or U13934 (N_13934,N_7947,N_7114);
nand U13935 (N_13935,N_6409,N_6496);
or U13936 (N_13936,N_6396,N_9800);
and U13937 (N_13937,N_9590,N_5314);
nand U13938 (N_13938,N_7569,N_6613);
or U13939 (N_13939,N_7647,N_7190);
and U13940 (N_13940,N_5803,N_7098);
and U13941 (N_13941,N_6977,N_7991);
and U13942 (N_13942,N_5997,N_5173);
or U13943 (N_13943,N_9826,N_6025);
and U13944 (N_13944,N_6626,N_8534);
and U13945 (N_13945,N_7415,N_7992);
and U13946 (N_13946,N_5922,N_6357);
nor U13947 (N_13947,N_9784,N_6008);
nand U13948 (N_13948,N_7516,N_5883);
and U13949 (N_13949,N_9228,N_9701);
nand U13950 (N_13950,N_6416,N_5077);
xor U13951 (N_13951,N_9649,N_5757);
and U13952 (N_13952,N_8118,N_9665);
and U13953 (N_13953,N_5093,N_6125);
xnor U13954 (N_13954,N_9174,N_5444);
nor U13955 (N_13955,N_5790,N_8345);
or U13956 (N_13956,N_9116,N_7207);
or U13957 (N_13957,N_7028,N_5565);
nor U13958 (N_13958,N_6726,N_5708);
nand U13959 (N_13959,N_8881,N_6909);
nor U13960 (N_13960,N_9909,N_7062);
nand U13961 (N_13961,N_7770,N_5535);
and U13962 (N_13962,N_5659,N_8310);
nor U13963 (N_13963,N_7114,N_8329);
nor U13964 (N_13964,N_7697,N_6529);
nor U13965 (N_13965,N_9503,N_6209);
nand U13966 (N_13966,N_9312,N_6727);
nand U13967 (N_13967,N_8327,N_9365);
nand U13968 (N_13968,N_9168,N_7294);
or U13969 (N_13969,N_7717,N_6089);
and U13970 (N_13970,N_6528,N_6376);
xor U13971 (N_13971,N_6806,N_5249);
nor U13972 (N_13972,N_5972,N_5290);
or U13973 (N_13973,N_6053,N_7527);
nand U13974 (N_13974,N_5612,N_7563);
and U13975 (N_13975,N_5640,N_6662);
xnor U13976 (N_13976,N_5434,N_7043);
nand U13977 (N_13977,N_7590,N_8169);
nand U13978 (N_13978,N_5950,N_6874);
or U13979 (N_13979,N_7859,N_7961);
and U13980 (N_13980,N_9225,N_5817);
or U13981 (N_13981,N_5633,N_9664);
or U13982 (N_13982,N_6350,N_9458);
nand U13983 (N_13983,N_9545,N_8137);
and U13984 (N_13984,N_5240,N_5086);
nor U13985 (N_13985,N_6556,N_7664);
and U13986 (N_13986,N_5422,N_9863);
nor U13987 (N_13987,N_5276,N_7502);
nand U13988 (N_13988,N_6349,N_9898);
nor U13989 (N_13989,N_9494,N_7844);
nand U13990 (N_13990,N_9485,N_7829);
and U13991 (N_13991,N_8718,N_7986);
xnor U13992 (N_13992,N_9586,N_6779);
and U13993 (N_13993,N_5546,N_7365);
nor U13994 (N_13994,N_7697,N_8634);
nor U13995 (N_13995,N_8831,N_6474);
or U13996 (N_13996,N_8540,N_5625);
or U13997 (N_13997,N_6673,N_9345);
and U13998 (N_13998,N_9316,N_5957);
xnor U13999 (N_13999,N_5874,N_5388);
or U14000 (N_14000,N_8128,N_7060);
and U14001 (N_14001,N_7116,N_5789);
nand U14002 (N_14002,N_9088,N_9245);
and U14003 (N_14003,N_6036,N_5610);
nand U14004 (N_14004,N_5955,N_8965);
or U14005 (N_14005,N_6949,N_6730);
nand U14006 (N_14006,N_5260,N_9386);
nor U14007 (N_14007,N_7249,N_8052);
nand U14008 (N_14008,N_5398,N_5331);
nor U14009 (N_14009,N_6195,N_7878);
nor U14010 (N_14010,N_9666,N_8963);
nand U14011 (N_14011,N_6668,N_7052);
or U14012 (N_14012,N_7753,N_6131);
nand U14013 (N_14013,N_8457,N_6042);
and U14014 (N_14014,N_8566,N_6527);
nor U14015 (N_14015,N_5689,N_6256);
nor U14016 (N_14016,N_9868,N_8810);
nor U14017 (N_14017,N_5821,N_6640);
and U14018 (N_14018,N_8085,N_7481);
or U14019 (N_14019,N_7619,N_8501);
xor U14020 (N_14020,N_9062,N_5090);
or U14021 (N_14021,N_5096,N_6162);
nand U14022 (N_14022,N_7432,N_6935);
or U14023 (N_14023,N_6739,N_9295);
xor U14024 (N_14024,N_6403,N_6604);
and U14025 (N_14025,N_7231,N_9752);
and U14026 (N_14026,N_7415,N_6164);
nor U14027 (N_14027,N_7303,N_5626);
or U14028 (N_14028,N_9910,N_6742);
and U14029 (N_14029,N_9168,N_9891);
and U14030 (N_14030,N_9634,N_8420);
and U14031 (N_14031,N_7082,N_7004);
and U14032 (N_14032,N_6754,N_8831);
nor U14033 (N_14033,N_5528,N_7056);
nand U14034 (N_14034,N_8691,N_9769);
and U14035 (N_14035,N_6507,N_5132);
nand U14036 (N_14036,N_9002,N_6784);
or U14037 (N_14037,N_8807,N_7075);
nor U14038 (N_14038,N_7585,N_7839);
nor U14039 (N_14039,N_5022,N_9264);
or U14040 (N_14040,N_7688,N_5780);
nand U14041 (N_14041,N_5280,N_9552);
nand U14042 (N_14042,N_7996,N_6546);
xor U14043 (N_14043,N_6188,N_8092);
xor U14044 (N_14044,N_9546,N_7564);
nor U14045 (N_14045,N_8492,N_8351);
nand U14046 (N_14046,N_6153,N_9856);
and U14047 (N_14047,N_9105,N_8120);
or U14048 (N_14048,N_9749,N_8038);
nor U14049 (N_14049,N_9379,N_5574);
nand U14050 (N_14050,N_6119,N_5184);
nand U14051 (N_14051,N_6451,N_6907);
nand U14052 (N_14052,N_9693,N_6670);
nor U14053 (N_14053,N_9114,N_8706);
nor U14054 (N_14054,N_6753,N_5994);
and U14055 (N_14055,N_7861,N_7213);
nor U14056 (N_14056,N_6567,N_9297);
or U14057 (N_14057,N_9132,N_9490);
and U14058 (N_14058,N_6297,N_5413);
or U14059 (N_14059,N_7580,N_9494);
nand U14060 (N_14060,N_6797,N_8614);
nand U14061 (N_14061,N_6097,N_7172);
xnor U14062 (N_14062,N_7246,N_6959);
or U14063 (N_14063,N_9292,N_7006);
or U14064 (N_14064,N_9113,N_7500);
or U14065 (N_14065,N_8313,N_7340);
or U14066 (N_14066,N_6947,N_9097);
and U14067 (N_14067,N_8208,N_6185);
and U14068 (N_14068,N_7178,N_7110);
or U14069 (N_14069,N_7553,N_5961);
xnor U14070 (N_14070,N_7174,N_6307);
or U14071 (N_14071,N_7416,N_5455);
nand U14072 (N_14072,N_6290,N_8590);
nor U14073 (N_14073,N_6497,N_5110);
and U14074 (N_14074,N_8867,N_9759);
nand U14075 (N_14075,N_8112,N_8239);
xor U14076 (N_14076,N_6472,N_9840);
nand U14077 (N_14077,N_5128,N_7539);
xor U14078 (N_14078,N_5581,N_7975);
nor U14079 (N_14079,N_5338,N_9773);
nor U14080 (N_14080,N_9907,N_7231);
nor U14081 (N_14081,N_5723,N_8797);
and U14082 (N_14082,N_8519,N_7679);
nand U14083 (N_14083,N_6181,N_9938);
xor U14084 (N_14084,N_7835,N_7137);
nor U14085 (N_14085,N_7222,N_7479);
or U14086 (N_14086,N_5022,N_6592);
nor U14087 (N_14087,N_8327,N_8188);
nor U14088 (N_14088,N_5374,N_5695);
nand U14089 (N_14089,N_9824,N_7339);
and U14090 (N_14090,N_9250,N_6820);
xnor U14091 (N_14091,N_5065,N_9010);
or U14092 (N_14092,N_5532,N_8329);
nor U14093 (N_14093,N_5320,N_8493);
or U14094 (N_14094,N_6827,N_8629);
nand U14095 (N_14095,N_7249,N_8677);
xnor U14096 (N_14096,N_5625,N_5358);
nor U14097 (N_14097,N_7988,N_8285);
and U14098 (N_14098,N_7926,N_8024);
and U14099 (N_14099,N_8108,N_5493);
nor U14100 (N_14100,N_9343,N_9745);
nand U14101 (N_14101,N_6425,N_7766);
nor U14102 (N_14102,N_9794,N_5421);
nor U14103 (N_14103,N_8637,N_6466);
or U14104 (N_14104,N_6516,N_9244);
nor U14105 (N_14105,N_7223,N_6619);
nor U14106 (N_14106,N_8676,N_5353);
nor U14107 (N_14107,N_5310,N_9704);
nand U14108 (N_14108,N_5077,N_8575);
or U14109 (N_14109,N_7114,N_6567);
nor U14110 (N_14110,N_6550,N_7088);
or U14111 (N_14111,N_7044,N_8507);
nand U14112 (N_14112,N_7863,N_8837);
nand U14113 (N_14113,N_5114,N_9265);
nand U14114 (N_14114,N_8105,N_7943);
and U14115 (N_14115,N_6052,N_9402);
nor U14116 (N_14116,N_8874,N_9643);
nor U14117 (N_14117,N_5927,N_9573);
or U14118 (N_14118,N_5312,N_8782);
and U14119 (N_14119,N_5967,N_6274);
nor U14120 (N_14120,N_8380,N_5162);
nand U14121 (N_14121,N_6248,N_5538);
or U14122 (N_14122,N_7131,N_5192);
or U14123 (N_14123,N_5798,N_9461);
and U14124 (N_14124,N_7361,N_7639);
or U14125 (N_14125,N_7681,N_6274);
nor U14126 (N_14126,N_5322,N_5956);
or U14127 (N_14127,N_5007,N_8950);
nand U14128 (N_14128,N_5090,N_9510);
and U14129 (N_14129,N_9663,N_7679);
or U14130 (N_14130,N_9716,N_5915);
xnor U14131 (N_14131,N_7597,N_9488);
and U14132 (N_14132,N_7495,N_9864);
nor U14133 (N_14133,N_6775,N_5722);
and U14134 (N_14134,N_9104,N_7237);
nor U14135 (N_14135,N_8199,N_5073);
or U14136 (N_14136,N_8918,N_9838);
xor U14137 (N_14137,N_6821,N_8545);
and U14138 (N_14138,N_7454,N_7074);
and U14139 (N_14139,N_9035,N_9365);
xor U14140 (N_14140,N_9986,N_5514);
nand U14141 (N_14141,N_9409,N_7319);
and U14142 (N_14142,N_7964,N_7592);
xnor U14143 (N_14143,N_6455,N_9480);
nor U14144 (N_14144,N_9814,N_7626);
nand U14145 (N_14145,N_8522,N_6926);
xnor U14146 (N_14146,N_5619,N_8144);
or U14147 (N_14147,N_5091,N_8371);
and U14148 (N_14148,N_5552,N_6248);
and U14149 (N_14149,N_9299,N_9867);
and U14150 (N_14150,N_9702,N_9972);
nand U14151 (N_14151,N_8984,N_6216);
and U14152 (N_14152,N_9184,N_7731);
and U14153 (N_14153,N_7325,N_7718);
nand U14154 (N_14154,N_5693,N_7178);
xor U14155 (N_14155,N_7899,N_6571);
nor U14156 (N_14156,N_8233,N_7351);
nor U14157 (N_14157,N_7131,N_8057);
or U14158 (N_14158,N_7277,N_9068);
or U14159 (N_14159,N_9160,N_8156);
and U14160 (N_14160,N_8868,N_8473);
and U14161 (N_14161,N_9709,N_9109);
nand U14162 (N_14162,N_7379,N_8454);
or U14163 (N_14163,N_8149,N_8325);
nand U14164 (N_14164,N_5768,N_6934);
nand U14165 (N_14165,N_6354,N_8660);
and U14166 (N_14166,N_6626,N_9061);
xnor U14167 (N_14167,N_7173,N_5476);
nor U14168 (N_14168,N_6569,N_5432);
nand U14169 (N_14169,N_8813,N_7953);
nor U14170 (N_14170,N_8135,N_6303);
xnor U14171 (N_14171,N_7620,N_5229);
xnor U14172 (N_14172,N_7874,N_9622);
and U14173 (N_14173,N_6951,N_5660);
nor U14174 (N_14174,N_5887,N_8539);
xor U14175 (N_14175,N_5489,N_9146);
or U14176 (N_14176,N_8783,N_7222);
nand U14177 (N_14177,N_6919,N_6303);
and U14178 (N_14178,N_8095,N_8126);
or U14179 (N_14179,N_9481,N_9656);
nand U14180 (N_14180,N_9254,N_9763);
and U14181 (N_14181,N_9823,N_6118);
or U14182 (N_14182,N_5210,N_6467);
nand U14183 (N_14183,N_6686,N_9000);
and U14184 (N_14184,N_9572,N_5270);
nand U14185 (N_14185,N_5310,N_5647);
or U14186 (N_14186,N_8485,N_8352);
or U14187 (N_14187,N_7542,N_7996);
nor U14188 (N_14188,N_5948,N_6700);
xnor U14189 (N_14189,N_7313,N_6206);
and U14190 (N_14190,N_8635,N_5012);
nor U14191 (N_14191,N_6499,N_6373);
or U14192 (N_14192,N_8590,N_9082);
or U14193 (N_14193,N_9639,N_7939);
or U14194 (N_14194,N_6528,N_5092);
xnor U14195 (N_14195,N_6480,N_9161);
or U14196 (N_14196,N_5298,N_6390);
nand U14197 (N_14197,N_7004,N_9415);
and U14198 (N_14198,N_6412,N_5873);
nor U14199 (N_14199,N_5185,N_6887);
xnor U14200 (N_14200,N_8809,N_9721);
xnor U14201 (N_14201,N_5865,N_8673);
or U14202 (N_14202,N_7378,N_6161);
nor U14203 (N_14203,N_7884,N_7011);
and U14204 (N_14204,N_7485,N_7099);
and U14205 (N_14205,N_5872,N_7329);
or U14206 (N_14206,N_8127,N_9998);
nor U14207 (N_14207,N_6226,N_8996);
nor U14208 (N_14208,N_7914,N_8193);
nand U14209 (N_14209,N_7934,N_8229);
or U14210 (N_14210,N_7059,N_6293);
or U14211 (N_14211,N_7575,N_8867);
nand U14212 (N_14212,N_6125,N_7572);
or U14213 (N_14213,N_9485,N_7433);
nand U14214 (N_14214,N_9839,N_9899);
or U14215 (N_14215,N_8947,N_7383);
and U14216 (N_14216,N_9080,N_8526);
xnor U14217 (N_14217,N_8468,N_8026);
nand U14218 (N_14218,N_7308,N_8014);
xor U14219 (N_14219,N_8786,N_8915);
and U14220 (N_14220,N_6607,N_9229);
or U14221 (N_14221,N_8108,N_9403);
or U14222 (N_14222,N_9014,N_9548);
and U14223 (N_14223,N_6171,N_6098);
nand U14224 (N_14224,N_6604,N_7256);
nand U14225 (N_14225,N_7450,N_5755);
nor U14226 (N_14226,N_6573,N_7820);
nor U14227 (N_14227,N_7114,N_9030);
nand U14228 (N_14228,N_8931,N_8248);
and U14229 (N_14229,N_8002,N_7249);
nor U14230 (N_14230,N_8317,N_6482);
and U14231 (N_14231,N_8379,N_9721);
or U14232 (N_14232,N_5587,N_6474);
xor U14233 (N_14233,N_8993,N_8779);
or U14234 (N_14234,N_8977,N_6452);
or U14235 (N_14235,N_7631,N_8946);
nand U14236 (N_14236,N_5650,N_9380);
and U14237 (N_14237,N_8274,N_6950);
nor U14238 (N_14238,N_6520,N_9119);
xnor U14239 (N_14239,N_7763,N_5658);
and U14240 (N_14240,N_7994,N_7877);
nor U14241 (N_14241,N_9995,N_9182);
nor U14242 (N_14242,N_9477,N_6057);
nand U14243 (N_14243,N_8200,N_8887);
nor U14244 (N_14244,N_5869,N_7993);
or U14245 (N_14245,N_5463,N_6593);
nor U14246 (N_14246,N_5276,N_7170);
xnor U14247 (N_14247,N_7927,N_6036);
or U14248 (N_14248,N_7923,N_9573);
or U14249 (N_14249,N_6146,N_7650);
or U14250 (N_14250,N_6977,N_6988);
or U14251 (N_14251,N_9411,N_8489);
nor U14252 (N_14252,N_9452,N_5856);
xor U14253 (N_14253,N_6615,N_8388);
nand U14254 (N_14254,N_8167,N_5876);
nor U14255 (N_14255,N_8331,N_9277);
nand U14256 (N_14256,N_5960,N_6841);
nand U14257 (N_14257,N_8457,N_8760);
or U14258 (N_14258,N_6073,N_8614);
nor U14259 (N_14259,N_8821,N_8068);
nor U14260 (N_14260,N_7021,N_6188);
and U14261 (N_14261,N_5956,N_5323);
nand U14262 (N_14262,N_9553,N_5105);
xor U14263 (N_14263,N_6926,N_7414);
nand U14264 (N_14264,N_5035,N_6484);
nand U14265 (N_14265,N_9904,N_8432);
nand U14266 (N_14266,N_7576,N_7054);
and U14267 (N_14267,N_5782,N_9644);
or U14268 (N_14268,N_9400,N_8649);
nor U14269 (N_14269,N_5946,N_7851);
nor U14270 (N_14270,N_7002,N_6788);
xnor U14271 (N_14271,N_7532,N_9331);
and U14272 (N_14272,N_8114,N_6679);
and U14273 (N_14273,N_7220,N_6798);
and U14274 (N_14274,N_9606,N_8025);
nor U14275 (N_14275,N_8861,N_6420);
nor U14276 (N_14276,N_7416,N_5145);
nand U14277 (N_14277,N_8658,N_7807);
nor U14278 (N_14278,N_6596,N_6730);
nand U14279 (N_14279,N_7691,N_9989);
nand U14280 (N_14280,N_5662,N_9028);
or U14281 (N_14281,N_5524,N_7983);
nor U14282 (N_14282,N_9432,N_9171);
and U14283 (N_14283,N_9569,N_5479);
or U14284 (N_14284,N_7730,N_8224);
nor U14285 (N_14285,N_9042,N_5022);
xnor U14286 (N_14286,N_6393,N_8868);
nor U14287 (N_14287,N_7792,N_8840);
xnor U14288 (N_14288,N_9906,N_9130);
xor U14289 (N_14289,N_8866,N_8489);
and U14290 (N_14290,N_7760,N_5599);
or U14291 (N_14291,N_6383,N_8045);
nand U14292 (N_14292,N_6319,N_7139);
and U14293 (N_14293,N_6176,N_6080);
or U14294 (N_14294,N_5336,N_9987);
nand U14295 (N_14295,N_7884,N_8587);
and U14296 (N_14296,N_9556,N_9438);
xor U14297 (N_14297,N_5952,N_7019);
or U14298 (N_14298,N_5874,N_8623);
nand U14299 (N_14299,N_5248,N_7156);
xnor U14300 (N_14300,N_9674,N_9602);
or U14301 (N_14301,N_6930,N_8506);
nor U14302 (N_14302,N_7033,N_6871);
nor U14303 (N_14303,N_8992,N_9039);
and U14304 (N_14304,N_7420,N_5395);
or U14305 (N_14305,N_7208,N_5816);
or U14306 (N_14306,N_9769,N_7750);
and U14307 (N_14307,N_9838,N_8858);
nor U14308 (N_14308,N_5942,N_5215);
or U14309 (N_14309,N_5196,N_7824);
nor U14310 (N_14310,N_9233,N_5558);
or U14311 (N_14311,N_5462,N_8952);
xnor U14312 (N_14312,N_6061,N_9139);
or U14313 (N_14313,N_6011,N_5132);
and U14314 (N_14314,N_5775,N_9166);
nor U14315 (N_14315,N_9487,N_9521);
nand U14316 (N_14316,N_7241,N_8939);
nand U14317 (N_14317,N_7665,N_5418);
nor U14318 (N_14318,N_9406,N_8819);
nand U14319 (N_14319,N_5377,N_7667);
nor U14320 (N_14320,N_9248,N_7005);
and U14321 (N_14321,N_6094,N_6542);
or U14322 (N_14322,N_5956,N_5234);
nand U14323 (N_14323,N_8570,N_7717);
and U14324 (N_14324,N_5425,N_6438);
and U14325 (N_14325,N_6346,N_6956);
nor U14326 (N_14326,N_5341,N_5911);
nand U14327 (N_14327,N_5886,N_8226);
xnor U14328 (N_14328,N_6205,N_7969);
and U14329 (N_14329,N_8411,N_6773);
nor U14330 (N_14330,N_9024,N_6566);
nor U14331 (N_14331,N_9144,N_8857);
or U14332 (N_14332,N_9100,N_5092);
nand U14333 (N_14333,N_6245,N_8052);
nand U14334 (N_14334,N_9596,N_7860);
and U14335 (N_14335,N_6108,N_7255);
nor U14336 (N_14336,N_5387,N_8380);
and U14337 (N_14337,N_7445,N_5124);
and U14338 (N_14338,N_5179,N_6715);
nand U14339 (N_14339,N_8222,N_5437);
nor U14340 (N_14340,N_6569,N_9545);
and U14341 (N_14341,N_6428,N_8351);
nor U14342 (N_14342,N_6680,N_5523);
and U14343 (N_14343,N_9084,N_7029);
xnor U14344 (N_14344,N_7039,N_5181);
nand U14345 (N_14345,N_6343,N_5768);
nand U14346 (N_14346,N_8860,N_6938);
nand U14347 (N_14347,N_6027,N_5162);
xor U14348 (N_14348,N_6449,N_8433);
xor U14349 (N_14349,N_9057,N_8977);
xor U14350 (N_14350,N_6992,N_9471);
xor U14351 (N_14351,N_8232,N_7093);
or U14352 (N_14352,N_6315,N_5802);
nor U14353 (N_14353,N_7116,N_7229);
nor U14354 (N_14354,N_7828,N_7391);
and U14355 (N_14355,N_9247,N_7637);
nand U14356 (N_14356,N_8782,N_7592);
and U14357 (N_14357,N_9993,N_7772);
or U14358 (N_14358,N_9864,N_7168);
or U14359 (N_14359,N_8689,N_9591);
or U14360 (N_14360,N_9278,N_5460);
or U14361 (N_14361,N_5245,N_7435);
nor U14362 (N_14362,N_5838,N_5885);
nand U14363 (N_14363,N_9682,N_7680);
or U14364 (N_14364,N_8791,N_9183);
xnor U14365 (N_14365,N_8344,N_5082);
and U14366 (N_14366,N_9379,N_8854);
nand U14367 (N_14367,N_7722,N_7535);
or U14368 (N_14368,N_6984,N_5834);
or U14369 (N_14369,N_5522,N_9234);
and U14370 (N_14370,N_7366,N_5982);
nand U14371 (N_14371,N_9125,N_8541);
or U14372 (N_14372,N_7519,N_7616);
nand U14373 (N_14373,N_5299,N_8125);
nand U14374 (N_14374,N_9988,N_8110);
nand U14375 (N_14375,N_8622,N_7666);
nand U14376 (N_14376,N_7707,N_9492);
and U14377 (N_14377,N_8800,N_7908);
nand U14378 (N_14378,N_7139,N_9467);
and U14379 (N_14379,N_6612,N_5662);
nand U14380 (N_14380,N_7291,N_5772);
nand U14381 (N_14381,N_5824,N_5852);
nor U14382 (N_14382,N_8242,N_6103);
nand U14383 (N_14383,N_9591,N_9427);
xor U14384 (N_14384,N_6871,N_8247);
and U14385 (N_14385,N_7516,N_6490);
and U14386 (N_14386,N_9971,N_9193);
and U14387 (N_14387,N_5043,N_6252);
nand U14388 (N_14388,N_8469,N_5698);
or U14389 (N_14389,N_5969,N_9187);
and U14390 (N_14390,N_5038,N_5550);
and U14391 (N_14391,N_8009,N_6125);
nand U14392 (N_14392,N_7346,N_8705);
or U14393 (N_14393,N_8370,N_8371);
and U14394 (N_14394,N_7223,N_5680);
or U14395 (N_14395,N_8290,N_6874);
nand U14396 (N_14396,N_9172,N_5522);
xnor U14397 (N_14397,N_5461,N_6991);
or U14398 (N_14398,N_6870,N_8110);
and U14399 (N_14399,N_8931,N_8515);
nor U14400 (N_14400,N_9681,N_9796);
or U14401 (N_14401,N_7142,N_5528);
nor U14402 (N_14402,N_6674,N_7004);
nor U14403 (N_14403,N_6529,N_7166);
xnor U14404 (N_14404,N_9118,N_9498);
nor U14405 (N_14405,N_8102,N_8358);
nor U14406 (N_14406,N_8463,N_9747);
and U14407 (N_14407,N_5218,N_6004);
nand U14408 (N_14408,N_9281,N_9335);
nor U14409 (N_14409,N_8681,N_6475);
and U14410 (N_14410,N_9697,N_9194);
and U14411 (N_14411,N_5234,N_9222);
and U14412 (N_14412,N_5412,N_8579);
xor U14413 (N_14413,N_6448,N_5894);
nand U14414 (N_14414,N_7995,N_8964);
nor U14415 (N_14415,N_6776,N_5225);
nor U14416 (N_14416,N_7880,N_7222);
nand U14417 (N_14417,N_7540,N_6119);
nor U14418 (N_14418,N_7439,N_5575);
and U14419 (N_14419,N_7662,N_9893);
or U14420 (N_14420,N_6136,N_8092);
nand U14421 (N_14421,N_6185,N_6274);
xor U14422 (N_14422,N_8223,N_9473);
or U14423 (N_14423,N_7705,N_8990);
nor U14424 (N_14424,N_8051,N_6896);
nand U14425 (N_14425,N_8754,N_8278);
nand U14426 (N_14426,N_8962,N_6514);
nor U14427 (N_14427,N_5724,N_5262);
or U14428 (N_14428,N_9105,N_8116);
and U14429 (N_14429,N_9782,N_9752);
and U14430 (N_14430,N_7520,N_5516);
nor U14431 (N_14431,N_9180,N_9109);
xnor U14432 (N_14432,N_7529,N_7639);
nor U14433 (N_14433,N_7021,N_5044);
nand U14434 (N_14434,N_5934,N_5470);
nand U14435 (N_14435,N_6290,N_7039);
and U14436 (N_14436,N_5641,N_5582);
and U14437 (N_14437,N_8289,N_7094);
nor U14438 (N_14438,N_7851,N_6126);
and U14439 (N_14439,N_5204,N_8187);
or U14440 (N_14440,N_5602,N_9619);
nor U14441 (N_14441,N_6957,N_7700);
and U14442 (N_14442,N_8144,N_5839);
or U14443 (N_14443,N_8946,N_8496);
nor U14444 (N_14444,N_5792,N_7441);
nand U14445 (N_14445,N_7272,N_9734);
and U14446 (N_14446,N_8442,N_6568);
or U14447 (N_14447,N_8831,N_6434);
and U14448 (N_14448,N_7690,N_7638);
nand U14449 (N_14449,N_6272,N_5984);
nand U14450 (N_14450,N_5289,N_6029);
nor U14451 (N_14451,N_9353,N_8259);
nor U14452 (N_14452,N_6713,N_8005);
nand U14453 (N_14453,N_5941,N_8813);
or U14454 (N_14454,N_7607,N_8101);
nor U14455 (N_14455,N_8051,N_5660);
or U14456 (N_14456,N_9823,N_8196);
nor U14457 (N_14457,N_7916,N_8032);
and U14458 (N_14458,N_5095,N_8375);
nand U14459 (N_14459,N_9793,N_7084);
and U14460 (N_14460,N_5003,N_6513);
and U14461 (N_14461,N_8695,N_7013);
and U14462 (N_14462,N_7372,N_6567);
and U14463 (N_14463,N_6442,N_9810);
and U14464 (N_14464,N_9913,N_6053);
and U14465 (N_14465,N_5245,N_9960);
nand U14466 (N_14466,N_8195,N_6782);
and U14467 (N_14467,N_6878,N_8959);
nor U14468 (N_14468,N_7161,N_5537);
nor U14469 (N_14469,N_6326,N_6353);
or U14470 (N_14470,N_7614,N_7232);
nor U14471 (N_14471,N_5055,N_8509);
and U14472 (N_14472,N_5777,N_8852);
and U14473 (N_14473,N_8545,N_5853);
nor U14474 (N_14474,N_9575,N_5930);
or U14475 (N_14475,N_6715,N_7411);
nor U14476 (N_14476,N_6402,N_9438);
or U14477 (N_14477,N_6135,N_7849);
nor U14478 (N_14478,N_5706,N_9710);
nor U14479 (N_14479,N_9711,N_9849);
and U14480 (N_14480,N_5125,N_7679);
nand U14481 (N_14481,N_5548,N_7202);
nor U14482 (N_14482,N_6757,N_5903);
nor U14483 (N_14483,N_7169,N_9864);
xor U14484 (N_14484,N_5106,N_6710);
and U14485 (N_14485,N_7226,N_6447);
nor U14486 (N_14486,N_5053,N_7159);
nand U14487 (N_14487,N_9781,N_5462);
nand U14488 (N_14488,N_8073,N_7160);
xor U14489 (N_14489,N_7657,N_5091);
nor U14490 (N_14490,N_9762,N_6010);
and U14491 (N_14491,N_9208,N_7612);
nor U14492 (N_14492,N_5638,N_8082);
nand U14493 (N_14493,N_9670,N_7107);
xor U14494 (N_14494,N_6833,N_8803);
xnor U14495 (N_14495,N_8005,N_5055);
and U14496 (N_14496,N_7244,N_6134);
and U14497 (N_14497,N_6815,N_8893);
nor U14498 (N_14498,N_7378,N_8702);
xor U14499 (N_14499,N_8848,N_9982);
nor U14500 (N_14500,N_5324,N_6036);
nand U14501 (N_14501,N_8398,N_8199);
or U14502 (N_14502,N_8292,N_7556);
and U14503 (N_14503,N_7435,N_9254);
nand U14504 (N_14504,N_8071,N_7991);
or U14505 (N_14505,N_8640,N_6544);
nand U14506 (N_14506,N_5187,N_5400);
nor U14507 (N_14507,N_9417,N_8909);
or U14508 (N_14508,N_8747,N_6666);
nand U14509 (N_14509,N_9949,N_7487);
nand U14510 (N_14510,N_9728,N_6161);
or U14511 (N_14511,N_6949,N_5582);
nand U14512 (N_14512,N_5302,N_7615);
nand U14513 (N_14513,N_9350,N_6780);
and U14514 (N_14514,N_6190,N_9801);
or U14515 (N_14515,N_9086,N_8178);
or U14516 (N_14516,N_6467,N_5008);
nand U14517 (N_14517,N_8933,N_9756);
nor U14518 (N_14518,N_5998,N_9219);
or U14519 (N_14519,N_6374,N_6965);
nor U14520 (N_14520,N_7652,N_9067);
or U14521 (N_14521,N_7451,N_9064);
and U14522 (N_14522,N_7175,N_6358);
and U14523 (N_14523,N_8133,N_8622);
xnor U14524 (N_14524,N_6723,N_7979);
and U14525 (N_14525,N_6164,N_6431);
and U14526 (N_14526,N_6701,N_6962);
or U14527 (N_14527,N_5940,N_7333);
nand U14528 (N_14528,N_5274,N_8866);
and U14529 (N_14529,N_7187,N_6596);
nand U14530 (N_14530,N_8186,N_8662);
nand U14531 (N_14531,N_6723,N_6693);
nand U14532 (N_14532,N_6185,N_7535);
nand U14533 (N_14533,N_6597,N_5514);
and U14534 (N_14534,N_7378,N_9750);
nand U14535 (N_14535,N_5143,N_8329);
nor U14536 (N_14536,N_5129,N_5637);
and U14537 (N_14537,N_9128,N_9986);
nor U14538 (N_14538,N_9990,N_7349);
nor U14539 (N_14539,N_6414,N_9189);
nor U14540 (N_14540,N_7212,N_5043);
nor U14541 (N_14541,N_8429,N_5935);
or U14542 (N_14542,N_6196,N_7960);
nor U14543 (N_14543,N_7887,N_9122);
or U14544 (N_14544,N_5276,N_7149);
nor U14545 (N_14545,N_8437,N_6838);
xor U14546 (N_14546,N_8099,N_9599);
or U14547 (N_14547,N_6725,N_6238);
or U14548 (N_14548,N_9981,N_8005);
and U14549 (N_14549,N_6944,N_5687);
and U14550 (N_14550,N_6027,N_6445);
and U14551 (N_14551,N_8260,N_7620);
and U14552 (N_14552,N_6957,N_7203);
xor U14553 (N_14553,N_5632,N_8902);
xor U14554 (N_14554,N_6888,N_7084);
or U14555 (N_14555,N_8488,N_8485);
and U14556 (N_14556,N_8313,N_9295);
nand U14557 (N_14557,N_5922,N_9832);
and U14558 (N_14558,N_9936,N_7717);
and U14559 (N_14559,N_6679,N_5046);
nand U14560 (N_14560,N_7050,N_5406);
and U14561 (N_14561,N_8297,N_7270);
xnor U14562 (N_14562,N_7808,N_5700);
nor U14563 (N_14563,N_7531,N_6958);
and U14564 (N_14564,N_5026,N_8271);
nand U14565 (N_14565,N_8573,N_9302);
nand U14566 (N_14566,N_7777,N_5446);
nor U14567 (N_14567,N_5548,N_9925);
or U14568 (N_14568,N_5329,N_9301);
or U14569 (N_14569,N_5409,N_8080);
nor U14570 (N_14570,N_5958,N_8766);
or U14571 (N_14571,N_5857,N_8975);
or U14572 (N_14572,N_5089,N_9046);
and U14573 (N_14573,N_9738,N_7360);
and U14574 (N_14574,N_9661,N_7568);
nand U14575 (N_14575,N_8626,N_9992);
nand U14576 (N_14576,N_5239,N_6649);
or U14577 (N_14577,N_8126,N_6412);
and U14578 (N_14578,N_9348,N_7548);
nor U14579 (N_14579,N_7916,N_7398);
xnor U14580 (N_14580,N_8020,N_8474);
and U14581 (N_14581,N_8107,N_5686);
nand U14582 (N_14582,N_6514,N_6282);
nand U14583 (N_14583,N_8047,N_5675);
nand U14584 (N_14584,N_9718,N_9254);
nor U14585 (N_14585,N_6175,N_8756);
nor U14586 (N_14586,N_6342,N_7396);
nor U14587 (N_14587,N_6759,N_5226);
or U14588 (N_14588,N_6766,N_8395);
nor U14589 (N_14589,N_5388,N_9558);
nor U14590 (N_14590,N_9618,N_5159);
or U14591 (N_14591,N_5920,N_6082);
or U14592 (N_14592,N_9737,N_8064);
or U14593 (N_14593,N_5053,N_6392);
and U14594 (N_14594,N_8231,N_9176);
and U14595 (N_14595,N_8870,N_5054);
nand U14596 (N_14596,N_7479,N_7545);
nor U14597 (N_14597,N_9108,N_5946);
nand U14598 (N_14598,N_8904,N_5546);
and U14599 (N_14599,N_7694,N_6002);
and U14600 (N_14600,N_6325,N_5398);
nand U14601 (N_14601,N_8312,N_5948);
xnor U14602 (N_14602,N_5849,N_7346);
or U14603 (N_14603,N_6213,N_5712);
xor U14604 (N_14604,N_8256,N_9519);
and U14605 (N_14605,N_5337,N_5533);
and U14606 (N_14606,N_7053,N_8607);
and U14607 (N_14607,N_7472,N_9970);
and U14608 (N_14608,N_7897,N_9421);
nand U14609 (N_14609,N_5821,N_8812);
nor U14610 (N_14610,N_5721,N_7422);
and U14611 (N_14611,N_8169,N_7785);
and U14612 (N_14612,N_5255,N_7581);
nand U14613 (N_14613,N_7039,N_8044);
nand U14614 (N_14614,N_9376,N_8275);
and U14615 (N_14615,N_9549,N_6336);
and U14616 (N_14616,N_6420,N_7796);
or U14617 (N_14617,N_6861,N_5116);
xnor U14618 (N_14618,N_8327,N_9596);
nand U14619 (N_14619,N_7894,N_7480);
or U14620 (N_14620,N_5938,N_7457);
xnor U14621 (N_14621,N_7046,N_8193);
nand U14622 (N_14622,N_5964,N_6452);
and U14623 (N_14623,N_5002,N_8255);
and U14624 (N_14624,N_7520,N_6691);
and U14625 (N_14625,N_7498,N_9076);
xor U14626 (N_14626,N_6215,N_8646);
xnor U14627 (N_14627,N_7845,N_9804);
xnor U14628 (N_14628,N_9944,N_7235);
or U14629 (N_14629,N_7818,N_7688);
nor U14630 (N_14630,N_7628,N_6656);
or U14631 (N_14631,N_8828,N_5615);
nand U14632 (N_14632,N_6031,N_7483);
nand U14633 (N_14633,N_5625,N_6982);
and U14634 (N_14634,N_5441,N_5676);
nand U14635 (N_14635,N_5715,N_5465);
and U14636 (N_14636,N_5029,N_8193);
nand U14637 (N_14637,N_6462,N_7921);
nor U14638 (N_14638,N_6539,N_5874);
and U14639 (N_14639,N_5113,N_7111);
and U14640 (N_14640,N_9864,N_6240);
nor U14641 (N_14641,N_5232,N_8530);
nor U14642 (N_14642,N_9949,N_8567);
xor U14643 (N_14643,N_6581,N_6077);
nor U14644 (N_14644,N_8641,N_9011);
and U14645 (N_14645,N_8763,N_8205);
nor U14646 (N_14646,N_9020,N_6145);
xnor U14647 (N_14647,N_6628,N_7974);
nor U14648 (N_14648,N_7093,N_8162);
and U14649 (N_14649,N_5848,N_8513);
nand U14650 (N_14650,N_9838,N_8154);
nor U14651 (N_14651,N_5042,N_8912);
nor U14652 (N_14652,N_7477,N_7417);
nand U14653 (N_14653,N_6669,N_5630);
nor U14654 (N_14654,N_5690,N_8632);
nor U14655 (N_14655,N_5349,N_8504);
and U14656 (N_14656,N_7966,N_5961);
or U14657 (N_14657,N_8468,N_7390);
nand U14658 (N_14658,N_6179,N_9651);
nand U14659 (N_14659,N_6980,N_7854);
nand U14660 (N_14660,N_6861,N_9045);
or U14661 (N_14661,N_5161,N_7612);
nor U14662 (N_14662,N_8347,N_6055);
xnor U14663 (N_14663,N_6136,N_9155);
or U14664 (N_14664,N_8540,N_7065);
nor U14665 (N_14665,N_8558,N_9481);
nor U14666 (N_14666,N_5411,N_7072);
or U14667 (N_14667,N_8659,N_6830);
or U14668 (N_14668,N_7613,N_9967);
nor U14669 (N_14669,N_5412,N_5369);
nor U14670 (N_14670,N_6018,N_6556);
or U14671 (N_14671,N_8906,N_9211);
nand U14672 (N_14672,N_9462,N_8427);
and U14673 (N_14673,N_9000,N_9894);
and U14674 (N_14674,N_9947,N_9324);
or U14675 (N_14675,N_7538,N_6161);
nand U14676 (N_14676,N_9438,N_9589);
xor U14677 (N_14677,N_9631,N_8749);
and U14678 (N_14678,N_5588,N_8991);
nand U14679 (N_14679,N_7278,N_9101);
nor U14680 (N_14680,N_9046,N_9559);
xnor U14681 (N_14681,N_5887,N_9406);
or U14682 (N_14682,N_6133,N_5496);
nand U14683 (N_14683,N_8304,N_5661);
nor U14684 (N_14684,N_8074,N_7948);
and U14685 (N_14685,N_6100,N_6688);
nand U14686 (N_14686,N_5279,N_8195);
and U14687 (N_14687,N_8869,N_6667);
xor U14688 (N_14688,N_9785,N_8840);
and U14689 (N_14689,N_7242,N_9463);
nand U14690 (N_14690,N_5422,N_8655);
or U14691 (N_14691,N_7669,N_5071);
nand U14692 (N_14692,N_8245,N_5159);
or U14693 (N_14693,N_7053,N_6197);
nor U14694 (N_14694,N_5182,N_9103);
or U14695 (N_14695,N_7392,N_5077);
and U14696 (N_14696,N_5116,N_6691);
or U14697 (N_14697,N_5278,N_8804);
or U14698 (N_14698,N_7896,N_9987);
nand U14699 (N_14699,N_9644,N_7257);
and U14700 (N_14700,N_5155,N_9494);
and U14701 (N_14701,N_7155,N_9530);
nor U14702 (N_14702,N_5902,N_8457);
and U14703 (N_14703,N_5074,N_9869);
nor U14704 (N_14704,N_7082,N_7319);
xor U14705 (N_14705,N_7464,N_7516);
nor U14706 (N_14706,N_5861,N_7024);
nand U14707 (N_14707,N_8405,N_9871);
and U14708 (N_14708,N_5215,N_8250);
and U14709 (N_14709,N_9410,N_9512);
and U14710 (N_14710,N_9793,N_6918);
nor U14711 (N_14711,N_9862,N_7574);
and U14712 (N_14712,N_6724,N_8871);
nor U14713 (N_14713,N_9523,N_6145);
and U14714 (N_14714,N_9506,N_5866);
or U14715 (N_14715,N_5496,N_6292);
and U14716 (N_14716,N_7482,N_7214);
nand U14717 (N_14717,N_7735,N_7501);
or U14718 (N_14718,N_5759,N_7627);
nand U14719 (N_14719,N_7921,N_6007);
xnor U14720 (N_14720,N_7494,N_5539);
or U14721 (N_14721,N_9928,N_9129);
and U14722 (N_14722,N_7652,N_6407);
and U14723 (N_14723,N_7681,N_6528);
nand U14724 (N_14724,N_5546,N_6229);
xnor U14725 (N_14725,N_7461,N_9979);
and U14726 (N_14726,N_6068,N_7547);
and U14727 (N_14727,N_9674,N_5771);
or U14728 (N_14728,N_7234,N_6634);
nand U14729 (N_14729,N_7983,N_7390);
nand U14730 (N_14730,N_5896,N_7090);
or U14731 (N_14731,N_6711,N_6033);
and U14732 (N_14732,N_7649,N_8887);
and U14733 (N_14733,N_6373,N_8367);
nand U14734 (N_14734,N_7528,N_9331);
and U14735 (N_14735,N_8893,N_6563);
nand U14736 (N_14736,N_5311,N_5002);
nor U14737 (N_14737,N_7112,N_5117);
nand U14738 (N_14738,N_5557,N_9380);
and U14739 (N_14739,N_5641,N_6355);
nor U14740 (N_14740,N_6336,N_5886);
nor U14741 (N_14741,N_5860,N_8286);
or U14742 (N_14742,N_6940,N_8956);
or U14743 (N_14743,N_6070,N_8226);
nand U14744 (N_14744,N_9223,N_7976);
and U14745 (N_14745,N_7423,N_5697);
or U14746 (N_14746,N_6518,N_5553);
or U14747 (N_14747,N_7850,N_6699);
and U14748 (N_14748,N_5151,N_9106);
nand U14749 (N_14749,N_5324,N_5639);
and U14750 (N_14750,N_6636,N_7247);
nand U14751 (N_14751,N_9102,N_7706);
and U14752 (N_14752,N_8940,N_8871);
nor U14753 (N_14753,N_6158,N_9855);
and U14754 (N_14754,N_6568,N_8098);
nor U14755 (N_14755,N_5738,N_6547);
or U14756 (N_14756,N_7530,N_7782);
or U14757 (N_14757,N_5477,N_7680);
nor U14758 (N_14758,N_7860,N_6290);
nor U14759 (N_14759,N_9641,N_5844);
or U14760 (N_14760,N_7430,N_9336);
or U14761 (N_14761,N_6599,N_7128);
xnor U14762 (N_14762,N_5947,N_8798);
or U14763 (N_14763,N_7966,N_7490);
and U14764 (N_14764,N_8050,N_5887);
and U14765 (N_14765,N_7444,N_5415);
nand U14766 (N_14766,N_5242,N_9701);
nor U14767 (N_14767,N_8212,N_6447);
xor U14768 (N_14768,N_7034,N_7043);
nor U14769 (N_14769,N_7585,N_5919);
xnor U14770 (N_14770,N_5551,N_9928);
or U14771 (N_14771,N_9483,N_9819);
nor U14772 (N_14772,N_6440,N_9344);
xnor U14773 (N_14773,N_5039,N_7669);
nand U14774 (N_14774,N_6098,N_6214);
nand U14775 (N_14775,N_5084,N_7409);
or U14776 (N_14776,N_5562,N_9306);
xor U14777 (N_14777,N_5431,N_6898);
and U14778 (N_14778,N_8080,N_5502);
or U14779 (N_14779,N_7272,N_8238);
or U14780 (N_14780,N_6526,N_6993);
or U14781 (N_14781,N_8589,N_9947);
nand U14782 (N_14782,N_5194,N_6689);
or U14783 (N_14783,N_7594,N_7968);
nor U14784 (N_14784,N_7916,N_9345);
nand U14785 (N_14785,N_6090,N_8880);
nand U14786 (N_14786,N_8494,N_5476);
and U14787 (N_14787,N_7139,N_6435);
or U14788 (N_14788,N_5318,N_7522);
or U14789 (N_14789,N_5764,N_5051);
nor U14790 (N_14790,N_9271,N_9376);
nand U14791 (N_14791,N_7168,N_7461);
nor U14792 (N_14792,N_6307,N_9812);
or U14793 (N_14793,N_9628,N_5201);
or U14794 (N_14794,N_5606,N_8269);
nand U14795 (N_14795,N_6305,N_5065);
or U14796 (N_14796,N_9290,N_6874);
and U14797 (N_14797,N_9499,N_6368);
nand U14798 (N_14798,N_9361,N_5184);
or U14799 (N_14799,N_5146,N_9602);
nor U14800 (N_14800,N_7140,N_8195);
nor U14801 (N_14801,N_9668,N_5828);
nor U14802 (N_14802,N_9437,N_7815);
nand U14803 (N_14803,N_9957,N_6911);
and U14804 (N_14804,N_6810,N_5711);
and U14805 (N_14805,N_8515,N_6992);
nor U14806 (N_14806,N_6956,N_6516);
nand U14807 (N_14807,N_9906,N_5670);
nand U14808 (N_14808,N_6070,N_9001);
nor U14809 (N_14809,N_7611,N_5983);
or U14810 (N_14810,N_6292,N_7572);
or U14811 (N_14811,N_8131,N_8803);
nor U14812 (N_14812,N_6240,N_7157);
nand U14813 (N_14813,N_8392,N_6850);
or U14814 (N_14814,N_5385,N_7875);
nand U14815 (N_14815,N_5264,N_5740);
xnor U14816 (N_14816,N_9276,N_6097);
nand U14817 (N_14817,N_6114,N_5851);
nor U14818 (N_14818,N_8189,N_6350);
nor U14819 (N_14819,N_8420,N_8548);
nand U14820 (N_14820,N_8267,N_6739);
or U14821 (N_14821,N_9535,N_8824);
and U14822 (N_14822,N_6085,N_9020);
or U14823 (N_14823,N_5090,N_5430);
nor U14824 (N_14824,N_6871,N_5531);
nor U14825 (N_14825,N_9491,N_8959);
and U14826 (N_14826,N_5430,N_9553);
and U14827 (N_14827,N_8580,N_7299);
xor U14828 (N_14828,N_9037,N_6882);
xor U14829 (N_14829,N_6772,N_6882);
or U14830 (N_14830,N_7017,N_9839);
and U14831 (N_14831,N_7287,N_9561);
nand U14832 (N_14832,N_5509,N_8587);
nor U14833 (N_14833,N_5897,N_9898);
and U14834 (N_14834,N_7913,N_7370);
or U14835 (N_14835,N_6344,N_9732);
or U14836 (N_14836,N_8869,N_5831);
nand U14837 (N_14837,N_5382,N_7790);
and U14838 (N_14838,N_8219,N_9082);
nand U14839 (N_14839,N_6489,N_6063);
nor U14840 (N_14840,N_6058,N_5525);
nand U14841 (N_14841,N_8198,N_8756);
nor U14842 (N_14842,N_6475,N_6664);
or U14843 (N_14843,N_7591,N_6016);
or U14844 (N_14844,N_5317,N_8777);
and U14845 (N_14845,N_7510,N_8565);
or U14846 (N_14846,N_8086,N_7468);
nor U14847 (N_14847,N_5522,N_6390);
nand U14848 (N_14848,N_8656,N_6281);
nor U14849 (N_14849,N_9537,N_5901);
xor U14850 (N_14850,N_5227,N_8898);
and U14851 (N_14851,N_8377,N_6059);
nor U14852 (N_14852,N_7925,N_5312);
nor U14853 (N_14853,N_5225,N_9328);
or U14854 (N_14854,N_8396,N_6661);
nor U14855 (N_14855,N_8480,N_6514);
nor U14856 (N_14856,N_7180,N_7236);
xnor U14857 (N_14857,N_6876,N_9366);
nor U14858 (N_14858,N_6631,N_5726);
xor U14859 (N_14859,N_5900,N_8294);
or U14860 (N_14860,N_5301,N_6464);
nand U14861 (N_14861,N_7705,N_7553);
nand U14862 (N_14862,N_5408,N_5204);
or U14863 (N_14863,N_5832,N_7110);
and U14864 (N_14864,N_6050,N_6275);
and U14865 (N_14865,N_5849,N_5028);
or U14866 (N_14866,N_6552,N_6521);
nand U14867 (N_14867,N_6647,N_5726);
or U14868 (N_14868,N_5114,N_9895);
or U14869 (N_14869,N_9305,N_7881);
nand U14870 (N_14870,N_6677,N_9173);
nand U14871 (N_14871,N_8445,N_6502);
nand U14872 (N_14872,N_6524,N_7513);
nor U14873 (N_14873,N_9513,N_6499);
nand U14874 (N_14874,N_6112,N_8538);
and U14875 (N_14875,N_9527,N_5648);
and U14876 (N_14876,N_8241,N_6048);
and U14877 (N_14877,N_9389,N_8062);
and U14878 (N_14878,N_7946,N_7712);
and U14879 (N_14879,N_6211,N_8741);
nor U14880 (N_14880,N_6940,N_9607);
xor U14881 (N_14881,N_7772,N_9738);
nand U14882 (N_14882,N_9611,N_8677);
nand U14883 (N_14883,N_9697,N_9599);
nand U14884 (N_14884,N_5022,N_6908);
xor U14885 (N_14885,N_5757,N_7258);
xor U14886 (N_14886,N_6775,N_8154);
nand U14887 (N_14887,N_8776,N_7118);
xor U14888 (N_14888,N_7376,N_6067);
or U14889 (N_14889,N_6823,N_8446);
and U14890 (N_14890,N_9845,N_7063);
and U14891 (N_14891,N_9561,N_9909);
or U14892 (N_14892,N_7311,N_8464);
nor U14893 (N_14893,N_7849,N_7703);
nand U14894 (N_14894,N_7323,N_6290);
or U14895 (N_14895,N_9900,N_9274);
xor U14896 (N_14896,N_6487,N_9713);
and U14897 (N_14897,N_5176,N_9969);
nor U14898 (N_14898,N_5825,N_5540);
and U14899 (N_14899,N_9460,N_8167);
nand U14900 (N_14900,N_7027,N_9573);
and U14901 (N_14901,N_6124,N_8323);
or U14902 (N_14902,N_6864,N_6330);
and U14903 (N_14903,N_7991,N_5992);
and U14904 (N_14904,N_9541,N_8177);
xnor U14905 (N_14905,N_5663,N_7552);
nand U14906 (N_14906,N_9596,N_7717);
nor U14907 (N_14907,N_9585,N_5758);
xor U14908 (N_14908,N_5224,N_5661);
and U14909 (N_14909,N_7567,N_7695);
nand U14910 (N_14910,N_8860,N_8116);
or U14911 (N_14911,N_6582,N_7482);
nand U14912 (N_14912,N_6401,N_8224);
and U14913 (N_14913,N_6420,N_7146);
nor U14914 (N_14914,N_7828,N_7135);
or U14915 (N_14915,N_6134,N_8380);
or U14916 (N_14916,N_8149,N_7873);
nor U14917 (N_14917,N_8890,N_8196);
nand U14918 (N_14918,N_9612,N_9097);
nor U14919 (N_14919,N_6162,N_5871);
xnor U14920 (N_14920,N_8895,N_8923);
and U14921 (N_14921,N_9615,N_5268);
and U14922 (N_14922,N_9636,N_5059);
and U14923 (N_14923,N_6956,N_6978);
nand U14924 (N_14924,N_5273,N_6961);
nand U14925 (N_14925,N_7019,N_7864);
nand U14926 (N_14926,N_8001,N_8852);
nor U14927 (N_14927,N_6035,N_8781);
and U14928 (N_14928,N_5603,N_6092);
or U14929 (N_14929,N_7637,N_7650);
or U14930 (N_14930,N_9240,N_8756);
xor U14931 (N_14931,N_5085,N_6756);
or U14932 (N_14932,N_5169,N_8753);
and U14933 (N_14933,N_5757,N_7552);
nor U14934 (N_14934,N_6735,N_5051);
and U14935 (N_14935,N_5920,N_7833);
nand U14936 (N_14936,N_5214,N_6070);
and U14937 (N_14937,N_8482,N_7915);
nand U14938 (N_14938,N_5380,N_5993);
and U14939 (N_14939,N_7768,N_7328);
nand U14940 (N_14940,N_8695,N_5531);
and U14941 (N_14941,N_6114,N_8488);
or U14942 (N_14942,N_9033,N_9364);
or U14943 (N_14943,N_8698,N_8541);
nand U14944 (N_14944,N_5613,N_9492);
nor U14945 (N_14945,N_6810,N_5002);
and U14946 (N_14946,N_7582,N_6447);
and U14947 (N_14947,N_6787,N_5355);
nor U14948 (N_14948,N_9697,N_9386);
xnor U14949 (N_14949,N_7567,N_7552);
or U14950 (N_14950,N_8677,N_9055);
and U14951 (N_14951,N_7538,N_9635);
nor U14952 (N_14952,N_7681,N_8509);
xor U14953 (N_14953,N_8127,N_8436);
and U14954 (N_14954,N_9340,N_9593);
nand U14955 (N_14955,N_6474,N_8684);
and U14956 (N_14956,N_5153,N_5852);
nand U14957 (N_14957,N_8081,N_6829);
nor U14958 (N_14958,N_5814,N_9393);
or U14959 (N_14959,N_6584,N_9677);
and U14960 (N_14960,N_6494,N_5576);
or U14961 (N_14961,N_8390,N_8451);
nor U14962 (N_14962,N_6006,N_8685);
xor U14963 (N_14963,N_9912,N_9485);
or U14964 (N_14964,N_6537,N_5790);
and U14965 (N_14965,N_7870,N_7681);
nand U14966 (N_14966,N_7587,N_8151);
and U14967 (N_14967,N_9088,N_5579);
nand U14968 (N_14968,N_9813,N_5942);
or U14969 (N_14969,N_6181,N_5053);
or U14970 (N_14970,N_5414,N_5622);
and U14971 (N_14971,N_7296,N_6264);
or U14972 (N_14972,N_6941,N_9630);
nand U14973 (N_14973,N_8078,N_6369);
nand U14974 (N_14974,N_8725,N_5794);
nand U14975 (N_14975,N_5008,N_7791);
nand U14976 (N_14976,N_8355,N_8837);
or U14977 (N_14977,N_6614,N_5078);
nor U14978 (N_14978,N_5348,N_5370);
or U14979 (N_14979,N_7976,N_7692);
and U14980 (N_14980,N_5470,N_5161);
or U14981 (N_14981,N_7094,N_8053);
or U14982 (N_14982,N_6922,N_9068);
and U14983 (N_14983,N_5676,N_6468);
xnor U14984 (N_14984,N_6461,N_9377);
nor U14985 (N_14985,N_5077,N_8671);
xnor U14986 (N_14986,N_8821,N_6780);
or U14987 (N_14987,N_6537,N_8505);
nand U14988 (N_14988,N_5438,N_5408);
or U14989 (N_14989,N_9916,N_9861);
nor U14990 (N_14990,N_7303,N_6714);
or U14991 (N_14991,N_9887,N_7058);
nor U14992 (N_14992,N_6567,N_9291);
and U14993 (N_14993,N_9549,N_5892);
nand U14994 (N_14994,N_6635,N_9565);
nor U14995 (N_14995,N_7778,N_9240);
xnor U14996 (N_14996,N_9654,N_8194);
nand U14997 (N_14997,N_9156,N_5941);
nand U14998 (N_14998,N_6143,N_9940);
nor U14999 (N_14999,N_8218,N_5105);
and U15000 (N_15000,N_13428,N_10746);
or U15001 (N_15001,N_10769,N_14887);
nand U15002 (N_15002,N_14534,N_12045);
and U15003 (N_15003,N_13090,N_12129);
nand U15004 (N_15004,N_13681,N_14413);
nor U15005 (N_15005,N_10911,N_13599);
nor U15006 (N_15006,N_10389,N_14407);
xnor U15007 (N_15007,N_13429,N_12611);
nor U15008 (N_15008,N_14997,N_10284);
nand U15009 (N_15009,N_11497,N_12671);
xnor U15010 (N_15010,N_12016,N_12894);
or U15011 (N_15011,N_12314,N_13733);
nand U15012 (N_15012,N_13687,N_14859);
or U15013 (N_15013,N_13401,N_10337);
nand U15014 (N_15014,N_12091,N_11176);
and U15015 (N_15015,N_13947,N_10042);
and U15016 (N_15016,N_13528,N_10381);
nand U15017 (N_15017,N_12086,N_11329);
nor U15018 (N_15018,N_10397,N_12307);
nor U15019 (N_15019,N_13637,N_10522);
or U15020 (N_15020,N_12521,N_12906);
or U15021 (N_15021,N_12678,N_14619);
nand U15022 (N_15022,N_12940,N_12143);
nand U15023 (N_15023,N_13778,N_12490);
nand U15024 (N_15024,N_12549,N_12784);
or U15025 (N_15025,N_11663,N_12869);
nand U15026 (N_15026,N_12547,N_11340);
nand U15027 (N_15027,N_10182,N_10120);
or U15028 (N_15028,N_13828,N_14272);
xor U15029 (N_15029,N_12475,N_12529);
xor U15030 (N_15030,N_13409,N_11810);
nand U15031 (N_15031,N_11233,N_10311);
or U15032 (N_15032,N_10817,N_11991);
nand U15033 (N_15033,N_14021,N_13595);
nor U15034 (N_15034,N_13743,N_10516);
or U15035 (N_15035,N_13500,N_14654);
xnor U15036 (N_15036,N_13193,N_10652);
and U15037 (N_15037,N_13965,N_14628);
nand U15038 (N_15038,N_10904,N_12881);
nand U15039 (N_15039,N_10637,N_11613);
xnor U15040 (N_15040,N_11175,N_13502);
xnor U15041 (N_15041,N_11589,N_13818);
nor U15042 (N_15042,N_10358,N_10479);
and U15043 (N_15043,N_12087,N_12638);
nor U15044 (N_15044,N_10335,N_10260);
nor U15045 (N_15045,N_12964,N_11461);
xor U15046 (N_15046,N_11580,N_14632);
nand U15047 (N_15047,N_10588,N_12172);
nor U15048 (N_15048,N_13136,N_14872);
nand U15049 (N_15049,N_14219,N_13508);
or U15050 (N_15050,N_14816,N_12453);
or U15051 (N_15051,N_13648,N_14792);
or U15052 (N_15052,N_10357,N_14122);
xnor U15053 (N_15053,N_13601,N_14095);
xor U15054 (N_15054,N_13945,N_13123);
nand U15055 (N_15055,N_11996,N_11983);
nand U15056 (N_15056,N_12102,N_10642);
xor U15057 (N_15057,N_12957,N_10520);
nor U15058 (N_15058,N_11487,N_13179);
or U15059 (N_15059,N_14115,N_13115);
nand U15060 (N_15060,N_14360,N_10569);
nand U15061 (N_15061,N_12867,N_14811);
or U15062 (N_15062,N_13685,N_11404);
nand U15063 (N_15063,N_10749,N_13373);
and U15064 (N_15064,N_14314,N_12511);
nor U15065 (N_15065,N_10411,N_10849);
nand U15066 (N_15066,N_13762,N_14941);
and U15067 (N_15067,N_11002,N_14414);
or U15068 (N_15068,N_13151,N_11909);
xnor U15069 (N_15069,N_11857,N_13354);
xnor U15070 (N_15070,N_12442,N_11345);
nand U15071 (N_15071,N_10062,N_11185);
and U15072 (N_15072,N_13333,N_14500);
nand U15073 (N_15073,N_10709,N_10139);
and U15074 (N_15074,N_13911,N_13886);
nand U15075 (N_15075,N_12724,N_12455);
nor U15076 (N_15076,N_14329,N_14452);
or U15077 (N_15077,N_13114,N_14768);
and U15078 (N_15078,N_14305,N_14819);
nand U15079 (N_15079,N_10860,N_11736);
or U15080 (N_15080,N_12734,N_10681);
nor U15081 (N_15081,N_12268,N_13993);
nor U15082 (N_15082,N_11808,N_14116);
and U15083 (N_15083,N_10835,N_11799);
nand U15084 (N_15084,N_10744,N_12259);
and U15085 (N_15085,N_10005,N_13348);
xor U15086 (N_15086,N_10007,N_12066);
and U15087 (N_15087,N_14156,N_10159);
or U15088 (N_15088,N_10444,N_12236);
and U15089 (N_15089,N_10067,N_11207);
or U15090 (N_15090,N_13990,N_10981);
or U15091 (N_15091,N_14922,N_13150);
or U15092 (N_15092,N_14847,N_11761);
nand U15093 (N_15093,N_10465,N_13269);
and U15094 (N_15094,N_14126,N_12341);
nand U15095 (N_15095,N_14641,N_12757);
nand U15096 (N_15096,N_11769,N_14580);
nor U15097 (N_15097,N_13244,N_11555);
or U15098 (N_15098,N_12523,N_11143);
or U15099 (N_15099,N_12979,N_14627);
and U15100 (N_15100,N_11014,N_14103);
xnor U15101 (N_15101,N_10099,N_13312);
nand U15102 (N_15102,N_14213,N_12030);
nand U15103 (N_15103,N_11858,N_10288);
and U15104 (N_15104,N_10793,N_14386);
or U15105 (N_15105,N_12868,N_10676);
or U15106 (N_15106,N_11362,N_14513);
xnor U15107 (N_15107,N_14027,N_14001);
or U15108 (N_15108,N_10096,N_13506);
xnor U15109 (N_15109,N_10338,N_14633);
nand U15110 (N_15110,N_14173,N_12099);
nor U15111 (N_15111,N_10447,N_13768);
nand U15112 (N_15112,N_12194,N_14446);
and U15113 (N_15113,N_10997,N_11814);
nor U15114 (N_15114,N_11147,N_11048);
nor U15115 (N_15115,N_12753,N_12234);
and U15116 (N_15116,N_13520,N_12324);
nand U15117 (N_15117,N_10626,N_13544);
nor U15118 (N_15118,N_10100,N_11079);
nand U15119 (N_15119,N_12269,N_11480);
and U15120 (N_15120,N_12127,N_10719);
or U15121 (N_15121,N_13960,N_11010);
and U15122 (N_15122,N_10897,N_10307);
xnor U15123 (N_15123,N_14221,N_11964);
nand U15124 (N_15124,N_10540,N_12850);
nor U15125 (N_15125,N_14114,N_13198);
nand U15126 (N_15126,N_11894,N_10234);
or U15127 (N_15127,N_13356,N_11112);
or U15128 (N_15128,N_13570,N_13636);
and U15129 (N_15129,N_14226,N_14032);
nor U15130 (N_15130,N_14992,N_13522);
nand U15131 (N_15131,N_11144,N_13660);
nand U15132 (N_15132,N_11256,N_12592);
xor U15133 (N_15133,N_12833,N_14042);
or U15134 (N_15134,N_12758,N_12261);
or U15135 (N_15135,N_12243,N_14083);
and U15136 (N_15136,N_10106,N_11790);
nor U15137 (N_15137,N_12928,N_13596);
xor U15138 (N_15138,N_11101,N_14248);
and U15139 (N_15139,N_11383,N_11561);
nand U15140 (N_15140,N_12262,N_12913);
xor U15141 (N_15141,N_14434,N_14472);
nand U15142 (N_15142,N_14635,N_14063);
nor U15143 (N_15143,N_12403,N_10842);
and U15144 (N_15144,N_11444,N_13635);
or U15145 (N_15145,N_11392,N_10325);
and U15146 (N_15146,N_12827,N_11577);
nor U15147 (N_15147,N_14172,N_13930);
nor U15148 (N_15148,N_10323,N_13718);
nand U15149 (N_15149,N_14821,N_10063);
nand U15150 (N_15150,N_12154,N_11693);
and U15151 (N_15151,N_10261,N_14842);
and U15152 (N_15152,N_12935,N_14369);
xor U15153 (N_15153,N_12445,N_12700);
and U15154 (N_15154,N_13547,N_14899);
xnor U15155 (N_15155,N_14312,N_10259);
nand U15156 (N_15156,N_14445,N_11998);
or U15157 (N_15157,N_13414,N_11262);
nand U15158 (N_15158,N_13017,N_13974);
and U15159 (N_15159,N_11355,N_12610);
and U15160 (N_15160,N_14541,N_10901);
nor U15161 (N_15161,N_11850,N_13604);
nor U15162 (N_15162,N_12842,N_11700);
nor U15163 (N_15163,N_11091,N_11372);
nand U15164 (N_15164,N_10002,N_12205);
xor U15165 (N_15165,N_11007,N_14080);
or U15166 (N_15166,N_14603,N_13292);
nor U15167 (N_15167,N_13258,N_11085);
xor U15168 (N_15168,N_11518,N_13479);
or U15169 (N_15169,N_12464,N_14300);
or U15170 (N_15170,N_10346,N_10299);
nor U15171 (N_15171,N_12369,N_11695);
nor U15172 (N_15172,N_10995,N_11968);
or U15173 (N_15173,N_14400,N_10797);
or U15174 (N_15174,N_12480,N_12681);
nor U15175 (N_15175,N_13232,N_11221);
nand U15176 (N_15176,N_11039,N_12658);
and U15177 (N_15177,N_12804,N_12003);
nand U15178 (N_15178,N_11942,N_11706);
or U15179 (N_15179,N_12690,N_10424);
or U15180 (N_15180,N_14709,N_13709);
and U15181 (N_15181,N_11180,N_10623);
and U15182 (N_15182,N_11327,N_12704);
and U15183 (N_15183,N_11364,N_13240);
or U15184 (N_15184,N_11645,N_11703);
and U15185 (N_15185,N_14136,N_12532);
nand U15186 (N_15186,N_10718,N_11911);
and U15187 (N_15187,N_12508,N_13282);
and U15188 (N_15188,N_14542,N_14128);
nand U15189 (N_15189,N_13840,N_13933);
nor U15190 (N_15190,N_10431,N_14134);
nor U15191 (N_15191,N_11644,N_14878);
nor U15192 (N_15192,N_12315,N_11542);
or U15193 (N_15193,N_14165,N_12162);
nand U15194 (N_15194,N_14223,N_13235);
or U15195 (N_15195,N_14530,N_10295);
nand U15196 (N_15196,N_10858,N_11801);
nor U15197 (N_15197,N_10929,N_10183);
nor U15198 (N_15198,N_13915,N_11688);
or U15199 (N_15199,N_11873,N_12503);
or U15200 (N_15200,N_11431,N_14455);
nor U15201 (N_15201,N_14191,N_10846);
or U15202 (N_15202,N_10024,N_11666);
or U15203 (N_15203,N_12527,N_13940);
nand U15204 (N_15204,N_10443,N_10170);
xnor U15205 (N_15205,N_14443,N_10954);
nor U15206 (N_15206,N_11677,N_14787);
nand U15207 (N_15207,N_13003,N_14484);
nor U15208 (N_15208,N_14293,N_12374);
nor U15209 (N_15209,N_11659,N_13287);
or U15210 (N_15210,N_13777,N_11713);
nor U15211 (N_15211,N_14592,N_13626);
and U15212 (N_15212,N_10300,N_11300);
nor U15213 (N_15213,N_14320,N_11776);
or U15214 (N_15214,N_11435,N_11584);
nand U15215 (N_15215,N_14815,N_11220);
and U15216 (N_15216,N_10494,N_10272);
nand U15217 (N_15217,N_11490,N_10659);
or U15218 (N_15218,N_12620,N_12947);
nor U15219 (N_15219,N_11935,N_13438);
nor U15220 (N_15220,N_14757,N_12103);
nor U15221 (N_15221,N_10376,N_13227);
nor U15222 (N_15222,N_13028,N_14192);
and U15223 (N_15223,N_13968,N_12082);
xor U15224 (N_15224,N_14038,N_12021);
xor U15225 (N_15225,N_13723,N_10871);
nand U15226 (N_15226,N_11832,N_10463);
or U15227 (N_15227,N_12150,N_14323);
nand U15228 (N_15228,N_12586,N_12722);
xnor U15229 (N_15229,N_11152,N_13276);
nand U15230 (N_15230,N_11162,N_14206);
and U15231 (N_15231,N_12557,N_11075);
and U15232 (N_15232,N_10016,N_11793);
nand U15233 (N_15233,N_10931,N_14169);
or U15234 (N_15234,N_14625,N_10332);
nand U15235 (N_15235,N_14236,N_12889);
nor U15236 (N_15236,N_13309,N_11575);
or U15237 (N_15237,N_14267,N_13592);
nand U15238 (N_15238,N_12924,N_10976);
nand U15239 (N_15239,N_14715,N_10693);
nor U15240 (N_15240,N_13259,N_12751);
or U15241 (N_15241,N_12594,N_11378);
or U15242 (N_15242,N_10449,N_10552);
xor U15243 (N_15243,N_12017,N_13856);
nor U15244 (N_15244,N_12248,N_14108);
or U15245 (N_15245,N_14729,N_14341);
nand U15246 (N_15246,N_12591,N_11042);
or U15247 (N_15247,N_14913,N_11377);
or U15248 (N_15248,N_10070,N_10894);
nand U15249 (N_15249,N_14000,N_10989);
nand U15250 (N_15250,N_10783,N_12944);
nand U15251 (N_15251,N_12798,N_10815);
nor U15252 (N_15252,N_10700,N_14177);
xnor U15253 (N_15253,N_14880,N_14692);
nor U15254 (N_15254,N_14297,N_12651);
or U15255 (N_15255,N_11366,N_11533);
nor U15256 (N_15256,N_12201,N_13187);
or U15257 (N_15257,N_10476,N_11811);
or U15258 (N_15258,N_13884,N_12417);
and U15259 (N_15259,N_13490,N_10194);
nor U15260 (N_15260,N_13204,N_12578);
nor U15261 (N_15261,N_14196,N_14767);
nor U15262 (N_15262,N_12258,N_10390);
nand U15263 (N_15263,N_10575,N_13266);
or U15264 (N_15264,N_11953,N_12545);
or U15265 (N_15265,N_11111,N_14486);
nor U15266 (N_15266,N_13427,N_13530);
nor U15267 (N_15267,N_13682,N_10730);
nor U15268 (N_15268,N_13816,N_12520);
or U15269 (N_15269,N_14858,N_13526);
and U15270 (N_15270,N_10727,N_11643);
or U15271 (N_15271,N_14102,N_14144);
xor U15272 (N_15272,N_14433,N_12037);
nor U15273 (N_15273,N_14860,N_11986);
xnor U15274 (N_15274,N_13537,N_14660);
and U15275 (N_15275,N_13398,N_10916);
xor U15276 (N_15276,N_10184,N_12141);
and U15277 (N_15277,N_14884,N_11123);
or U15278 (N_15278,N_11549,N_14519);
nor U15279 (N_15279,N_13847,N_11463);
and U15280 (N_15280,N_12956,N_10314);
nand U15281 (N_15281,N_13999,N_11158);
or U15282 (N_15282,N_12712,N_14317);
and U15283 (N_15283,N_12117,N_11865);
and U15284 (N_15284,N_11192,N_13486);
nand U15285 (N_15285,N_13832,N_10496);
nor U15286 (N_15286,N_14402,N_10172);
and U15287 (N_15287,N_12849,N_14886);
or U15288 (N_15288,N_11900,N_10638);
nor U15289 (N_15289,N_14578,N_14769);
nor U15290 (N_15290,N_10178,N_12422);
nor U15291 (N_15291,N_10636,N_11815);
nand U15292 (N_15292,N_14178,N_11563);
nand U15293 (N_15293,N_11129,N_11166);
and U15294 (N_15294,N_11806,N_10956);
xnor U15295 (N_15295,N_12534,N_11177);
and U15296 (N_15296,N_10662,N_13317);
nor U15297 (N_15297,N_14539,N_11318);
or U15298 (N_15298,N_14867,N_14969);
xor U15299 (N_15299,N_12145,N_12107);
nand U15300 (N_15300,N_12797,N_12996);
or U15301 (N_15301,N_14962,N_13914);
nor U15302 (N_15302,N_11100,N_14024);
nand U15303 (N_15303,N_14735,N_12937);
and U15304 (N_15304,N_13168,N_10750);
and U15305 (N_15305,N_10869,N_13834);
or U15306 (N_15306,N_10065,N_14512);
or U15307 (N_15307,N_12413,N_13955);
nand U15308 (N_15308,N_13837,N_12308);
nor U15309 (N_15309,N_11619,N_12392);
nor U15310 (N_15310,N_12619,N_11062);
nand U15311 (N_15311,N_11989,N_11015);
or U15312 (N_15312,N_11024,N_13802);
nand U15313 (N_15313,N_13656,N_11985);
nand U15314 (N_15314,N_14075,N_12014);
nand U15315 (N_15315,N_10045,N_10125);
nand U15316 (N_15316,N_14785,N_13923);
or U15317 (N_15317,N_10830,N_13581);
nand U15318 (N_15318,N_12961,N_13699);
nand U15319 (N_15319,N_11181,N_13800);
nand U15320 (N_15320,N_11813,N_11514);
nor U15321 (N_15321,N_10190,N_10874);
nor U15322 (N_15322,N_13824,N_11981);
nor U15323 (N_15323,N_10220,N_13518);
and U15324 (N_15324,N_13814,N_10383);
and U15325 (N_15325,N_11705,N_14575);
nand U15326 (N_15326,N_13891,N_14154);
or U15327 (N_15327,N_10786,N_14371);
nand U15328 (N_15328,N_12977,N_10036);
xnor U15329 (N_15329,N_12531,N_12760);
xor U15330 (N_15330,N_11474,N_12049);
and U15331 (N_15331,N_12763,N_14378);
nand U15332 (N_15332,N_11750,N_11076);
or U15333 (N_15333,N_13476,N_10561);
or U15334 (N_15334,N_13880,N_14170);
nand U15335 (N_15335,N_13070,N_13543);
or U15336 (N_15336,N_14664,N_14299);
nor U15337 (N_15337,N_11852,N_12285);
nand U15338 (N_15338,N_11585,N_12930);
or U15339 (N_15339,N_14220,N_11733);
nor U15340 (N_15340,N_10484,N_11120);
or U15341 (N_15341,N_14492,N_13576);
and U15342 (N_15342,N_11336,N_10084);
nand U15343 (N_15343,N_14079,N_12284);
nor U15344 (N_15344,N_14559,N_14622);
nor U15345 (N_15345,N_12096,N_11478);
or U15346 (N_15346,N_10453,N_14797);
or U15347 (N_15347,N_10739,N_10115);
nor U15348 (N_15348,N_10047,N_12186);
or U15349 (N_15349,N_13843,N_11970);
nand U15350 (N_15350,N_10820,N_13841);
nand U15351 (N_15351,N_14753,N_12782);
and U15352 (N_15352,N_11264,N_11106);
or U15353 (N_15353,N_12231,N_11895);
or U15354 (N_15354,N_13691,N_11684);
nand U15355 (N_15355,N_10359,N_13836);
nand U15356 (N_15356,N_10278,N_14645);
nor U15357 (N_15357,N_11127,N_10102);
nand U15358 (N_15358,N_14451,N_12479);
and U15359 (N_15359,N_13644,N_12837);
or U15360 (N_15360,N_13774,N_14623);
nor U15361 (N_15361,N_14538,N_10832);
nor U15362 (N_15362,N_14590,N_14249);
nor U15363 (N_15363,N_10882,N_13206);
nand U15364 (N_15364,N_11893,N_13555);
xor U15365 (N_15365,N_11548,N_10661);
or U15366 (N_15366,N_13689,N_11247);
nand U15367 (N_15367,N_13735,N_10663);
nand U15368 (N_15368,N_12768,N_12904);
and U15369 (N_15369,N_11373,N_14958);
nor U15370 (N_15370,N_14780,N_13741);
nand U15371 (N_15371,N_12943,N_14523);
nor U15372 (N_15372,N_11962,N_12239);
nor U15373 (N_15373,N_14171,N_13618);
and U15374 (N_15374,N_10111,N_14487);
nand U15375 (N_15375,N_14460,N_11060);
nor U15376 (N_15376,N_13922,N_12174);
or U15377 (N_15377,N_12701,N_11477);
and U15378 (N_15378,N_10581,N_10862);
nand U15379 (N_15379,N_12474,N_14980);
nor U15380 (N_15380,N_14588,N_12783);
or U15381 (N_15381,N_11482,N_10094);
nor U15382 (N_15382,N_12735,N_14928);
nor U15383 (N_15383,N_12719,N_10924);
nand U15384 (N_15384,N_13052,N_10231);
nor U15385 (N_15385,N_14937,N_12655);
xor U15386 (N_15386,N_14703,N_12555);
nor U15387 (N_15387,N_11056,N_11839);
nor U15388 (N_15388,N_13853,N_13089);
nand U15389 (N_15389,N_13598,N_11923);
nand U15390 (N_15390,N_10728,N_10428);
nand U15391 (N_15391,N_11363,N_13747);
and U15392 (N_15392,N_11065,N_14309);
and U15393 (N_15393,N_13374,N_11414);
nor U15394 (N_15394,N_11438,N_12368);
xnor U15395 (N_15395,N_11571,N_10748);
nor U15396 (N_15396,N_14574,N_14339);
xnor U15397 (N_15397,N_13190,N_11406);
and U15398 (N_15398,N_11907,N_10705);
and U15399 (N_15399,N_13305,N_11036);
and U15400 (N_15400,N_14977,N_14311);
or U15401 (N_15401,N_12978,N_11034);
nand U15402 (N_15402,N_14130,N_13324);
or U15403 (N_15403,N_13377,N_11081);
and U15404 (N_15404,N_10725,N_12663);
and U15405 (N_15405,N_11673,N_14676);
nand U15406 (N_15406,N_13865,N_13858);
nand U15407 (N_15407,N_12641,N_13446);
nand U15408 (N_15408,N_12486,N_11702);
nand U15409 (N_15409,N_13402,N_13810);
nor U15410 (N_15410,N_14274,N_14728);
nand U15411 (N_15411,N_11652,N_11339);
nor U15412 (N_15412,N_11789,N_14826);
nand U15413 (N_15413,N_11540,N_14450);
nand U15414 (N_15414,N_13166,N_11317);
nand U15415 (N_15415,N_11308,N_10157);
xnor U15416 (N_15416,N_12942,N_11605);
nand U15417 (N_15417,N_14188,N_14076);
or U15418 (N_15418,N_11301,N_12232);
nand U15419 (N_15419,N_11441,N_12384);
or U15420 (N_15420,N_14241,N_14935);
nor U15421 (N_15421,N_14074,N_11053);
nand U15422 (N_15422,N_13261,N_10187);
and U15423 (N_15423,N_12057,N_14256);
or U15424 (N_15424,N_10292,N_10457);
xnor U15425 (N_15425,N_11583,N_13307);
nor U15426 (N_15426,N_11795,N_10483);
nor U15427 (N_15427,N_10150,N_10471);
nand U15428 (N_15428,N_14184,N_14747);
or U15429 (N_15429,N_13091,N_11190);
xor U15430 (N_15430,N_12908,N_10205);
or U15431 (N_15431,N_14214,N_12170);
or U15432 (N_15432,N_11578,N_10472);
or U15433 (N_15433,N_13285,N_13254);
nand U15434 (N_15434,N_14572,N_13803);
nor U15435 (N_15435,N_10991,N_10826);
nor U15436 (N_15436,N_10630,N_13044);
nand U15437 (N_15437,N_13917,N_12482);
nor U15438 (N_15438,N_14945,N_14278);
and U15439 (N_15439,N_13162,N_11523);
nand U15440 (N_15440,N_13291,N_10501);
nand U15441 (N_15441,N_11669,N_11350);
nor U15442 (N_15442,N_10229,N_12350);
and U15443 (N_15443,N_14036,N_12795);
xor U15444 (N_15444,N_13642,N_10848);
nor U15445 (N_15445,N_12807,N_12874);
and U15446 (N_15446,N_10928,N_11326);
and U15447 (N_15447,N_11494,N_14324);
nor U15448 (N_15448,N_10072,N_13364);
nand U15449 (N_15449,N_11905,N_11504);
nand U15450 (N_15450,N_14630,N_13846);
and U15451 (N_15451,N_10854,N_14097);
and U15452 (N_15452,N_12607,N_11498);
nand U15453 (N_15453,N_11739,N_13729);
nand U15454 (N_15454,N_13465,N_12402);
and U15455 (N_15455,N_11073,N_14589);
and U15456 (N_15456,N_11754,N_14604);
nor U15457 (N_15457,N_12054,N_13049);
and U15458 (N_15458,N_11816,N_10404);
and U15459 (N_15459,N_12033,N_10083);
nor U15460 (N_15460,N_14783,N_13451);
xor U15461 (N_15461,N_12927,N_12685);
nand U15462 (N_15462,N_13455,N_13624);
and U15463 (N_15463,N_12856,N_14412);
and U15464 (N_15464,N_14639,N_11965);
or U15465 (N_15465,N_10140,N_11236);
or U15466 (N_15466,N_13929,N_11689);
and U15467 (N_15467,N_10915,N_12321);
nor U15468 (N_15468,N_13420,N_12726);
nor U15469 (N_15469,N_14012,N_14976);
or U15470 (N_15470,N_11631,N_13861);
nor U15471 (N_15471,N_11940,N_11579);
xor U15472 (N_15472,N_10114,N_14504);
or U15473 (N_15473,N_12838,N_14333);
nor U15474 (N_15474,N_12395,N_13724);
nor U15475 (N_15475,N_14495,N_10382);
and U15476 (N_15476,N_13279,N_13625);
xor U15477 (N_15477,N_14587,N_13630);
xnor U15478 (N_15478,N_14596,N_12061);
or U15479 (N_15479,N_10736,N_13772);
nand U15480 (N_15480,N_10087,N_10054);
and U15481 (N_15481,N_11245,N_11788);
nor U15482 (N_15482,N_10910,N_14035);
xor U15483 (N_15483,N_11067,N_10526);
nor U15484 (N_15484,N_13584,N_11777);
nor U15485 (N_15485,N_12467,N_12898);
or U15486 (N_15486,N_12713,N_13804);
nor U15487 (N_15487,N_10865,N_11222);
or U15488 (N_15488,N_11187,N_11827);
or U15489 (N_15489,N_11086,N_13726);
and U15490 (N_15490,N_12036,N_14798);
nor U15491 (N_15491,N_14059,N_10201);
and U15492 (N_15492,N_13120,N_12432);
xor U15493 (N_15493,N_11417,N_14268);
or U15494 (N_15494,N_11128,N_14907);
xnor U15495 (N_15495,N_10840,N_13807);
nor U15496 (N_15496,N_14135,N_13953);
nand U15497 (N_15497,N_10448,N_11179);
nor U15498 (N_15498,N_13361,N_12767);
nor U15499 (N_15499,N_10035,N_13692);
nand U15500 (N_15500,N_11202,N_13342);
and U15501 (N_15501,N_14934,N_11698);
nor U15502 (N_15502,N_13615,N_11430);
nand U15503 (N_15503,N_12624,N_10755);
and U15504 (N_15504,N_11945,N_14337);
nor U15505 (N_15505,N_13525,N_14258);
nor U15506 (N_15506,N_14218,N_13640);
or U15507 (N_15507,N_10870,N_13501);
and U15508 (N_15508,N_12222,N_11337);
nor U15509 (N_15509,N_14621,N_10658);
nor U15510 (N_15510,N_13739,N_11615);
nor U15511 (N_15511,N_10564,N_10691);
nor U15512 (N_15512,N_14540,N_11718);
xnor U15513 (N_15513,N_14914,N_14494);
and U15514 (N_15514,N_12195,N_14073);
nor U15515 (N_15515,N_11607,N_11822);
and U15516 (N_15516,N_11493,N_13157);
nand U15517 (N_15517,N_13434,N_10450);
xor U15518 (N_15518,N_13881,N_11590);
xnor U15519 (N_15519,N_13972,N_10161);
or U15520 (N_15520,N_11775,N_13766);
nor U15521 (N_15521,N_13565,N_12404);
nor U15522 (N_15522,N_13738,N_13613);
xnor U15523 (N_15523,N_12144,N_14933);
and U15524 (N_15524,N_13458,N_10060);
and U15525 (N_15525,N_12267,N_10608);
or U15526 (N_15526,N_11069,N_12998);
xnor U15527 (N_15527,N_12414,N_13875);
nor U15528 (N_15528,N_12139,N_13897);
and U15529 (N_15529,N_14854,N_13603);
and U15530 (N_15530,N_14802,N_12932);
and U15531 (N_15531,N_12007,N_13606);
xor U15532 (N_15532,N_12829,N_10364);
and U15533 (N_15533,N_12675,N_13484);
and U15534 (N_15534,N_11009,N_13622);
or U15535 (N_15535,N_11604,N_14975);
nand U15536 (N_15536,N_10713,N_12640);
xnor U15537 (N_15537,N_10554,N_14570);
nor U15538 (N_15538,N_14485,N_12771);
xor U15539 (N_15539,N_10572,N_13431);
and U15540 (N_15540,N_13505,N_10765);
or U15541 (N_15541,N_11840,N_13054);
and U15542 (N_15542,N_12759,N_12864);
nand U15543 (N_15543,N_11521,N_10212);
or U15544 (N_15544,N_14019,N_14929);
nor U15545 (N_15545,N_10688,N_13132);
or U15546 (N_15546,N_13888,N_11159);
and U15547 (N_15547,N_14704,N_14924);
nand U15548 (N_15548,N_10410,N_14834);
nor U15549 (N_15549,N_12509,N_10961);
nand U15550 (N_15550,N_12695,N_14824);
or U15551 (N_15551,N_13013,N_12809);
or U15552 (N_15552,N_13016,N_12202);
xor U15553 (N_15553,N_13012,N_11765);
nand U15554 (N_15554,N_11074,N_13869);
nor U15555 (N_15555,N_10394,N_11138);
or U15556 (N_15556,N_10009,N_10971);
and U15557 (N_15557,N_14522,N_11359);
nand U15558 (N_15558,N_14727,N_14959);
xnor U15559 (N_15559,N_10920,N_11136);
nor U15560 (N_15560,N_12953,N_14003);
or U15561 (N_15561,N_13108,N_14529);
nand U15562 (N_15562,N_12020,N_10669);
or U15563 (N_15563,N_10014,N_14751);
or U15564 (N_15564,N_12365,N_10982);
or U15565 (N_15565,N_11116,N_11535);
and U15566 (N_15566,N_14991,N_14612);
nand U15567 (N_15567,N_11785,N_11019);
nand U15568 (N_15568,N_14380,N_14548);
nor U15569 (N_15569,N_14475,N_13820);
nand U15570 (N_15570,N_13478,N_12176);
or U15571 (N_15571,N_14970,N_11454);
and U15572 (N_15572,N_10506,N_13055);
nand U15573 (N_15573,N_11194,N_11934);
nor U15574 (N_15574,N_14967,N_10167);
or U15575 (N_15575,N_11021,N_14391);
nand U15576 (N_15576,N_11341,N_10964);
nand U15577 (N_15577,N_10019,N_12083);
nor U15578 (N_15578,N_13098,N_12839);
nand U15579 (N_15579,N_10055,N_14424);
and U15580 (N_15580,N_13352,N_11562);
or U15581 (N_15581,N_10702,N_13664);
and U15582 (N_15582,N_11824,N_10290);
or U15583 (N_15583,N_13293,N_13189);
nand U15584 (N_15584,N_12791,N_13073);
and U15585 (N_15585,N_14536,N_10135);
or U15586 (N_15586,N_12821,N_11520);
nor U15587 (N_15587,N_11551,N_13201);
nand U15588 (N_15588,N_12301,N_13080);
and U15589 (N_15589,N_10972,N_13202);
nand U15590 (N_15590,N_13696,N_11331);
nand U15591 (N_15591,N_12461,N_11206);
and U15592 (N_15592,N_10377,N_12994);
nor U15593 (N_15593,N_14197,N_10156);
and U15594 (N_15594,N_12185,N_10493);
nand U15595 (N_15595,N_14840,N_12562);
or U15596 (N_15596,N_10811,N_14366);
or U15597 (N_15597,N_11741,N_12601);
xor U15598 (N_15598,N_12031,N_13347);
nor U15599 (N_15599,N_13253,N_14215);
and U15600 (N_15600,N_10855,N_14498);
xor U15601 (N_15601,N_11199,N_10647);
or U15602 (N_15602,N_12570,N_10959);
and U15603 (N_15603,N_11465,N_11939);
and U15604 (N_15604,N_11980,N_10185);
and U15605 (N_15605,N_13864,N_10442);
nor U15606 (N_15606,N_10085,N_14152);
or U15607 (N_15607,N_12811,N_14644);
nand U15608 (N_15608,N_14245,N_10729);
nand U15609 (N_15609,N_11918,N_14688);
xnor U15610 (N_15610,N_13734,N_11307);
nor U15611 (N_15611,N_14493,N_13335);
nor U15612 (N_15612,N_10142,N_12596);
nand U15613 (N_15613,N_11967,N_11955);
or U15614 (N_15614,N_10697,N_11637);
nand U15615 (N_15615,N_14874,N_13763);
or U15616 (N_15616,N_13112,N_14072);
nor U15617 (N_15617,N_11011,N_14225);
or U15618 (N_15618,N_13288,N_11216);
xor U15619 (N_15619,N_12071,N_14653);
xor U15620 (N_15620,N_13862,N_13755);
and U15621 (N_15621,N_12313,N_12788);
or U15622 (N_15622,N_11188,N_12317);
xor U15623 (N_15623,N_13872,N_14789);
nor U15624 (N_15624,N_11272,N_11505);
nand U15625 (N_15625,N_11415,N_14850);
nor U15626 (N_15626,N_10703,N_11835);
and U15627 (N_15627,N_10145,N_10204);
nor U15628 (N_15628,N_11608,N_11038);
and U15629 (N_15629,N_11146,N_10475);
or U15630 (N_15630,N_14813,N_12843);
or U15631 (N_15631,N_11712,N_12235);
or U15632 (N_15632,N_14543,N_12130);
and U15633 (N_15633,N_10550,N_10197);
or U15634 (N_15634,N_11211,N_10827);
or U15635 (N_15635,N_10488,N_14346);
and U15636 (N_15636,N_10504,N_14974);
and U15637 (N_15637,N_10628,N_14748);
and U15638 (N_15638,N_13384,N_10402);
and U15639 (N_15639,N_11358,N_14061);
or U15640 (N_15640,N_14940,N_10934);
and U15641 (N_15641,N_12832,N_13882);
and U15642 (N_15642,N_11325,N_11779);
nor U15643 (N_15643,N_14466,N_10490);
nor U15644 (N_15644,N_13238,N_11897);
or U15645 (N_15645,N_13719,N_12697);
nor U15646 (N_15646,N_10137,N_11035);
nor U15647 (N_15647,N_13638,N_10547);
and U15648 (N_15648,N_13663,N_11083);
or U15649 (N_15649,N_11771,N_12500);
xor U15650 (N_15650,N_11890,N_13967);
or U15651 (N_15651,N_11248,N_14004);
or U15652 (N_15652,N_12941,N_13809);
and U15653 (N_15653,N_14442,N_13243);
nor U15654 (N_15654,N_12214,N_13472);
nand U15655 (N_15655,N_14362,N_12175);
and U15656 (N_15656,N_12627,N_13318);
or U15657 (N_15657,N_12346,N_10246);
nor U15658 (N_15658,N_13776,N_11045);
or U15659 (N_15659,N_12633,N_12242);
or U15660 (N_15660,N_10451,N_12090);
or U15661 (N_15661,N_11390,N_13503);
and U15662 (N_15662,N_10644,N_12471);
nand U15663 (N_15663,N_10088,N_14605);
or U15664 (N_15664,N_12566,N_14952);
or U15665 (N_15665,N_12484,N_14185);
and U15666 (N_15666,N_10975,N_14138);
nand U15667 (N_15667,N_14803,N_10574);
or U15668 (N_15668,N_13694,N_14301);
xnor U15669 (N_15669,N_13524,N_12128);
xor U15670 (N_15670,N_10782,N_14893);
nor U15671 (N_15671,N_12420,N_11315);
xnor U15672 (N_15672,N_10925,N_14438);
and U15673 (N_15673,N_12292,N_14836);
nand U15674 (N_15674,N_11837,N_12347);
nand U15675 (N_15675,N_10505,N_10646);
and U15676 (N_15676,N_13935,N_11943);
nand U15677 (N_15677,N_12976,N_13556);
xnor U15678 (N_15678,N_14954,N_13903);
nand U15679 (N_15679,N_13445,N_14488);
or U15680 (N_15680,N_12389,N_13946);
nor U15681 (N_15681,N_11132,N_11834);
nor U15682 (N_15682,N_13097,N_13873);
nand U15683 (N_15683,N_13975,N_12830);
or U15684 (N_15684,N_11049,N_14009);
nand U15685 (N_15685,N_10257,N_10876);
nor U15686 (N_15686,N_12206,N_11794);
and U15687 (N_15687,N_11961,N_11087);
nand U15688 (N_15688,N_13651,N_10202);
and U15689 (N_15689,N_11472,N_12761);
or U15690 (N_15690,N_10710,N_12394);
nand U15691 (N_15691,N_13519,N_10199);
nor U15692 (N_15692,N_10879,N_11559);
or U15693 (N_15693,N_13184,N_10527);
nand U15694 (N_15694,N_13585,N_14989);
nor U15695 (N_15695,N_12564,N_10885);
nor U15696 (N_15696,N_13753,N_12255);
and U15697 (N_15697,N_13683,N_12524);
nor U15698 (N_15698,N_12501,N_12728);
xor U15699 (N_15699,N_13633,N_12951);
or U15700 (N_15700,N_11913,N_14014);
nor U15701 (N_15701,N_14711,N_10734);
or U15702 (N_15702,N_13916,N_11592);
nor U15703 (N_15703,N_13498,N_13621);
and U15704 (N_15704,N_11628,N_12851);
nor U15705 (N_15705,N_13079,N_13062);
nor U15706 (N_15706,N_11028,N_13989);
nand U15707 (N_15707,N_14626,N_12421);
nand U15708 (N_15708,N_11032,N_10824);
or U15709 (N_15709,N_10320,N_14374);
nor U15710 (N_15710,N_14765,N_12497);
nand U15711 (N_15711,N_12755,N_13218);
xnor U15712 (N_15712,N_11255,N_13363);
nand U15713 (N_15713,N_12826,N_13612);
or U15714 (N_15714,N_12358,N_13107);
nor U15715 (N_15715,N_11947,N_11522);
or U15716 (N_15716,N_11936,N_12866);
nand U15717 (N_15717,N_13155,N_13283);
and U15718 (N_15718,N_14981,N_11982);
nand U15719 (N_15719,N_12148,N_13966);
nor U15720 (N_15720,N_14071,N_14425);
nand U15721 (N_15721,N_10939,N_12900);
and U15722 (N_15722,N_12733,N_13433);
or U15723 (N_15723,N_14983,N_11241);
xor U15724 (N_15724,N_11883,N_10279);
nor U15725 (N_15725,N_10792,N_10984);
or U15726 (N_15726,N_12519,N_14761);
nand U15727 (N_15727,N_11587,N_12329);
nand U15728 (N_15728,N_14545,N_14919);
nor U15729 (N_15729,N_12647,N_13758);
or U15730 (N_15730,N_12665,N_14401);
nor U15731 (N_15731,N_11033,N_13617);
nor U15732 (N_15732,N_12011,N_10436);
nand U15733 (N_15733,N_10671,N_10429);
and U15734 (N_15734,N_12773,N_10640);
and U15735 (N_15735,N_11552,N_12548);
xor U15736 (N_15736,N_12561,N_12397);
nor U15737 (N_15737,N_10845,N_12418);
and U15738 (N_15738,N_11606,N_14395);
nor U15739 (N_15739,N_11809,N_12559);
and U15740 (N_15740,N_12462,N_11738);
and U15741 (N_15741,N_10834,N_11526);
or U15742 (N_15742,N_13004,N_11405);
nor U15743 (N_15743,N_11670,N_11416);
or U15744 (N_15744,N_10687,N_11999);
nor U15745 (N_15745,N_13793,N_13593);
and U15746 (N_15746,N_14732,N_14408);
or U15747 (N_15747,N_13550,N_12459);
nand U15748 (N_15748,N_12111,N_11117);
nand U15749 (N_15749,N_11979,N_14106);
or U15750 (N_15750,N_12664,N_11773);
and U15751 (N_15751,N_12122,N_11259);
or U15752 (N_15752,N_10254,N_10001);
or U15753 (N_15753,N_13646,N_10967);
or U15754 (N_15754,N_14775,N_13529);
nor U15755 (N_15755,N_12042,N_14088);
and U15756 (N_15756,N_11124,N_11830);
or U15757 (N_15757,N_14687,N_11952);
or U15758 (N_15758,N_12101,N_12750);
nand U15759 (N_15759,N_14505,N_10580);
or U15760 (N_15760,N_10666,N_11203);
or U15761 (N_15761,N_11838,N_12512);
nand U15762 (N_15762,N_11080,N_10542);
nor U15763 (N_15763,N_10452,N_10033);
and U15764 (N_15764,N_10586,N_10942);
and U15765 (N_15765,N_14658,N_14533);
or U15766 (N_15766,N_13801,N_13867);
nand U15767 (N_15767,N_13489,N_14026);
nor U15768 (N_15768,N_12730,N_10612);
or U15769 (N_15769,N_13769,N_14743);
nor U15770 (N_15770,N_14479,N_13815);
or U15771 (N_15771,N_13540,N_11055);
or U15772 (N_15772,N_11365,N_10406);
or U15773 (N_15773,N_14799,N_12211);
nand U15774 (N_15774,N_10305,N_10208);
nand U15775 (N_15775,N_12720,N_14280);
or U15776 (N_15776,N_11742,N_12598);
xnor U15777 (N_15777,N_12550,N_11110);
nor U15778 (N_15778,N_14276,N_14355);
nand U15779 (N_15779,N_13851,N_11064);
or U15780 (N_15780,N_11845,N_12863);
or U15781 (N_15781,N_10026,N_11061);
nor U15782 (N_15782,N_10076,N_12469);
and U15783 (N_15783,N_13000,N_11544);
nand U15784 (N_15784,N_12970,N_13313);
and U15785 (N_15785,N_10225,N_11948);
or U15786 (N_15786,N_10957,N_13591);
and U15787 (N_15787,N_11856,N_13181);
nand U15788 (N_15788,N_13199,N_13432);
or U15789 (N_15789,N_14938,N_10951);
nor U15790 (N_15790,N_13667,N_10021);
or U15791 (N_15791,N_13678,N_12081);
nand U15792 (N_15792,N_12064,N_13560);
nand U15793 (N_15793,N_14866,N_14212);
nor U15794 (N_15794,N_14851,N_10643);
or U15795 (N_15795,N_14168,N_10819);
nor U15796 (N_15796,N_11333,N_13388);
nand U15797 (N_15797,N_12390,N_12776);
xor U15798 (N_15798,N_10103,N_12896);
nand U15799 (N_15799,N_12051,N_11987);
xor U15800 (N_15800,N_11721,N_14978);
or U15801 (N_15801,N_13460,N_14372);
or U15802 (N_15802,N_12410,N_11319);
nor U15803 (N_15803,N_12583,N_13951);
nand U15804 (N_15804,N_14388,N_11859);
nor U15805 (N_15805,N_14340,N_10795);
or U15806 (N_15806,N_12920,N_14028);
nand U15807 (N_15807,N_14571,N_11624);
nand U15808 (N_15808,N_14861,N_14682);
nor U15809 (N_15809,N_14064,N_13210);
and U15810 (N_15810,N_13539,N_14648);
nand U15811 (N_15811,N_14689,N_13608);
nor U15812 (N_15812,N_11593,N_13453);
xnor U15813 (N_15813,N_14697,N_12067);
nand U15814 (N_15814,N_13693,N_11030);
or U15815 (N_15815,N_13284,N_11426);
and U15816 (N_15816,N_10711,N_10482);
nor U15817 (N_15817,N_11594,N_12425);
and U15818 (N_15818,N_13255,N_12180);
nand U15819 (N_15819,N_11413,N_12657);
nand U15820 (N_15820,N_11235,N_11418);
and U15821 (N_15821,N_12954,N_14927);
xnor U15822 (N_15822,N_14120,N_14582);
and U15823 (N_15823,N_11610,N_14602);
and U15824 (N_15824,N_12637,N_13871);
or U15825 (N_15825,N_11285,N_13789);
and U15826 (N_15826,N_10238,N_10618);
and U15827 (N_15827,N_10413,N_13126);
nand U15828 (N_15828,N_14232,N_12428);
xnor U15829 (N_15829,N_10531,N_11975);
or U15830 (N_15830,N_14678,N_10682);
nand U15831 (N_15831,N_11334,N_13614);
nand U15832 (N_15832,N_12073,N_10003);
and U15833 (N_15833,N_14207,N_11941);
or U15834 (N_15834,N_13779,N_12808);
nand U15835 (N_15835,N_13898,N_10888);
xnor U15836 (N_15836,N_11450,N_11541);
and U15837 (N_15837,N_14591,N_14930);
or U15838 (N_15838,N_13751,N_12636);
nand U15839 (N_15839,N_12539,N_10222);
nor U15840 (N_15840,N_13297,N_12485);
nand U15841 (N_15841,N_10441,N_10716);
nor U15842 (N_15842,N_13488,N_12609);
nand U15843 (N_15843,N_11862,N_12745);
xor U15844 (N_15844,N_12716,N_10203);
and U15845 (N_15845,N_13298,N_14755);
xnor U15846 (N_15846,N_11708,N_11547);
or U15847 (N_15847,N_10006,N_12575);
and U15848 (N_15848,N_12960,N_10985);
and U15849 (N_15849,N_12063,N_13991);
or U15850 (N_15850,N_12648,N_12965);
nor U15851 (N_15851,N_13437,N_11844);
nor U15852 (N_15852,N_14295,N_10392);
xor U15853 (N_15853,N_13554,N_11763);
or U15854 (N_15854,N_12834,N_11745);
and U15855 (N_15855,N_13260,N_11000);
or U15856 (N_15856,N_14511,N_11892);
xnor U15857 (N_15857,N_13538,N_13326);
nand U15858 (N_15858,N_14502,N_13175);
nand U15859 (N_15859,N_11025,N_13934);
and U15860 (N_15860,N_12567,N_12041);
nor U15861 (N_15861,N_11680,N_14674);
nor U15862 (N_15862,N_10768,N_11178);
and U15863 (N_15863,N_10685,N_13938);
or U15864 (N_15864,N_11658,N_14865);
or U15865 (N_15865,N_11507,N_10535);
xnor U15866 (N_15866,N_12424,N_10708);
or U15867 (N_15867,N_10511,N_10952);
nor U15868 (N_15868,N_12370,N_12613);
nor U15869 (N_15869,N_11407,N_12025);
or U15870 (N_15870,N_14086,N_14149);
and U15871 (N_15871,N_13826,N_11495);
nand U15872 (N_15872,N_10438,N_11956);
nand U15873 (N_15873,N_14030,N_11697);
nand U15874 (N_15874,N_11978,N_10706);
xor U15875 (N_15875,N_10566,N_10751);
nor U15876 (N_15876,N_12948,N_13075);
nor U15877 (N_15877,N_11230,N_14283);
and U15878 (N_15878,N_11774,N_10326);
xor U15879 (N_15879,N_11261,N_14045);
nand U15880 (N_15880,N_14099,N_13095);
or U15881 (N_15881,N_14145,N_10151);
nor U15882 (N_15882,N_13499,N_10240);
nor U15883 (N_15883,N_12891,N_14269);
xor U15884 (N_15884,N_13690,N_11927);
xnor U15885 (N_15885,N_12729,N_10822);
nand U15886 (N_15886,N_13732,N_10491);
and U15887 (N_15887,N_12399,N_11660);
nand U15888 (N_15888,N_14342,N_12731);
nand U15889 (N_15889,N_12212,N_14465);
or U15890 (N_15890,N_13513,N_14067);
xor U15891 (N_15891,N_13715,N_13746);
nor U15892 (N_15892,N_12670,N_11885);
and U15893 (N_15893,N_10348,N_13280);
and U15894 (N_15894,N_13406,N_13467);
nand U15895 (N_15895,N_11099,N_11841);
nand U15896 (N_15896,N_12777,N_11440);
or U15897 (N_15897,N_10095,N_10043);
or U15898 (N_15898,N_10650,N_11280);
or U15899 (N_15899,N_14742,N_14749);
xnor U15900 (N_15900,N_14895,N_13448);
nor U15901 (N_15901,N_12652,N_14563);
and U15902 (N_15902,N_13811,N_12668);
xnor U15903 (N_15903,N_10621,N_10470);
xor U15904 (N_15904,N_12325,N_12914);
and U15905 (N_15905,N_10629,N_12587);
and U15906 (N_15906,N_13926,N_14812);
and U15907 (N_15907,N_10969,N_14982);
nand U15908 (N_15908,N_12226,N_13979);
nor U15909 (N_15909,N_13493,N_13586);
xor U15910 (N_15910,N_12406,N_10507);
nand U15911 (N_15911,N_12157,N_14351);
xnor U15912 (N_15912,N_12882,N_10274);
and U15913 (N_15913,N_13575,N_11411);
or U15914 (N_15914,N_14259,N_10570);
nor U15915 (N_15915,N_11113,N_12472);
or U15916 (N_15916,N_14565,N_11924);
xnor U15917 (N_15917,N_14235,N_12643);
nor U15918 (N_15918,N_10360,N_12888);
xnor U15919 (N_15919,N_11385,N_13808);
and U15920 (N_15920,N_14525,N_12605);
and U15921 (N_15921,N_13362,N_14526);
and U15922 (N_15922,N_10767,N_14915);
and U15923 (N_15923,N_13343,N_11434);
nand U15924 (N_15924,N_14186,N_12448);
nand U15925 (N_15925,N_10678,N_10268);
nor U15926 (N_15926,N_10425,N_13127);
and U15927 (N_15927,N_11393,N_14005);
and U15928 (N_15928,N_11068,N_13470);
and U15929 (N_15929,N_11151,N_12385);
and U15930 (N_15930,N_12702,N_13410);
nor U15931 (N_15931,N_13509,N_10434);
nor U15932 (N_15932,N_13890,N_12688);
nand U15933 (N_15933,N_11517,N_14318);
nor U15934 (N_15934,N_13582,N_14679);
nor U15935 (N_15935,N_11225,N_11446);
xnor U15936 (N_15936,N_11442,N_10432);
or U15937 (N_15937,N_12094,N_10833);
nor U15938 (N_15938,N_11933,N_11994);
nor U15939 (N_15939,N_13386,N_14509);
or U15940 (N_15940,N_14471,N_10302);
and U15941 (N_15941,N_13963,N_10594);
and U15942 (N_15942,N_10027,N_10801);
nor U15943 (N_15943,N_13959,N_12553);
nand U15944 (N_15944,N_14949,N_10241);
nand U15945 (N_15945,N_10122,N_10000);
nand U15946 (N_15946,N_13063,N_10524);
and U15947 (N_15947,N_11908,N_13587);
and U15948 (N_15948,N_12493,N_14017);
and U15949 (N_15949,N_14161,N_12715);
and U15950 (N_15950,N_10480,N_13077);
nand U15951 (N_15951,N_13020,N_10741);
xnor U15952 (N_15952,N_12166,N_12216);
and U15953 (N_15953,N_13750,N_10174);
and U15954 (N_15954,N_14411,N_13397);
or U15955 (N_15955,N_11877,N_11565);
nand U15956 (N_15956,N_12056,N_10224);
or U15957 (N_15957,N_12775,N_14175);
or U15958 (N_15958,N_13909,N_12560);
or U15959 (N_15959,N_10478,N_11330);
and U15960 (N_15960,N_11369,N_11029);
nor U15961 (N_15961,N_10081,N_14650);
nor U15962 (N_15962,N_13588,N_11473);
nand U15963 (N_15963,N_12921,N_12433);
and U15964 (N_15964,N_13262,N_12585);
or U15965 (N_15965,N_11114,N_10181);
nor U15966 (N_15966,N_10930,N_14956);
or U15967 (N_15967,N_13985,N_12263);
nand U15968 (N_15968,N_10707,N_10753);
nand U15969 (N_15969,N_13605,N_13220);
and U15970 (N_15970,N_14375,N_13459);
nor U15971 (N_15971,N_14354,N_14501);
or U15972 (N_15972,N_11108,N_13874);
or U15973 (N_15973,N_13275,N_14011);
nor U15974 (N_15974,N_13619,N_10330);
or U15975 (N_15975,N_10074,N_11298);
or U15976 (N_15976,N_10657,N_10466);
nor U15977 (N_15977,N_10788,N_13759);
or U15978 (N_15978,N_11167,N_11229);
nor U15979 (N_15979,N_14569,N_14552);
nor U15980 (N_15980,N_10113,N_12931);
nor U15981 (N_15981,N_11534,N_14422);
nor U15982 (N_15982,N_11499,N_10266);
nor U15983 (N_15983,N_10439,N_12714);
xor U15984 (N_15984,N_10077,N_10474);
xnor U15985 (N_15985,N_11462,N_12053);
nor U15986 (N_15986,N_10189,N_12488);
xnor U15987 (N_15987,N_11251,N_14763);
nor U15988 (N_15988,N_12740,N_13019);
and U15989 (N_15989,N_10029,N_12893);
nor U15990 (N_15990,N_14925,N_14593);
and U15991 (N_15991,N_13389,N_14584);
nand U15992 (N_15992,N_13970,N_13887);
nor U15993 (N_15993,N_12322,N_12902);
nand U15994 (N_15994,N_14764,N_13106);
or U15995 (N_15995,N_12085,N_13393);
or U15996 (N_15996,N_13245,N_12528);
nor U15997 (N_15997,N_14174,N_11784);
nand U15998 (N_15998,N_13146,N_12848);
nor U15999 (N_15999,N_12793,N_10902);
nor U16000 (N_16000,N_14467,N_13430);
nor U16001 (N_16001,N_12219,N_12069);
nand U16002 (N_16002,N_13566,N_14912);
and U16003 (N_16003,N_14334,N_10576);
and U16004 (N_16004,N_13103,N_11254);
xnor U16005 (N_16005,N_12140,N_10602);
nand U16006 (N_16006,N_10866,N_14015);
nor U16007 (N_16007,N_12372,N_10887);
and U16008 (N_16008,N_10313,N_10356);
nor U16009 (N_16009,N_10296,N_11052);
xor U16010 (N_16010,N_11598,N_11460);
nand U16011 (N_16011,N_13021,N_13767);
nor U16012 (N_16012,N_11791,N_12095);
or U16013 (N_16013,N_13711,N_10992);
or U16014 (N_16014,N_12000,N_12373);
or U16015 (N_16015,N_13831,N_13242);
and U16016 (N_16016,N_13385,N_14151);
or U16017 (N_16017,N_12617,N_10403);
or U16018 (N_16018,N_13421,N_12916);
nand U16019 (N_16019,N_14008,N_12359);
nand U16020 (N_16020,N_10273,N_10587);
and U16021 (N_16021,N_10460,N_12077);
or U16022 (N_16022,N_12408,N_13294);
nor U16023 (N_16023,N_10617,N_13208);
nand U16024 (N_16024,N_12831,N_11884);
nand U16025 (N_16025,N_12249,N_12551);
or U16026 (N_16026,N_14998,N_14985);
or U16027 (N_16027,N_10909,N_13058);
nand U16028 (N_16028,N_13230,N_12023);
nor U16029 (N_16029,N_13299,N_11269);
and U16030 (N_16030,N_13558,N_11276);
or U16031 (N_16031,N_13203,N_11273);
nand U16032 (N_16032,N_10784,N_10400);
and U16033 (N_16033,N_14917,N_11012);
nand U16034 (N_16034,N_10131,N_12669);
and U16035 (N_16035,N_10154,N_14405);
nor U16036 (N_16036,N_10464,N_13191);
or U16037 (N_16037,N_11966,N_11286);
nand U16038 (N_16038,N_11448,N_10766);
and U16039 (N_16039,N_13885,N_12055);
and U16040 (N_16040,N_13957,N_14208);
nor U16041 (N_16041,N_10541,N_10092);
or U16042 (N_16042,N_11260,N_10068);
nor U16043 (N_16043,N_14430,N_12764);
nor U16044 (N_16044,N_10395,N_12810);
nor U16045 (N_16045,N_13607,N_11503);
xor U16046 (N_16046,N_12538,N_11977);
nand U16047 (N_16047,N_10673,N_10794);
nor U16048 (N_16048,N_10408,N_11277);
nor U16049 (N_16049,N_11831,N_10373);
nor U16050 (N_16050,N_14410,N_13662);
nor U16051 (N_16051,N_11546,N_11722);
and U16052 (N_16052,N_14598,N_14243);
and U16053 (N_16053,N_13906,N_11676);
or U16054 (N_16054,N_14266,N_10679);
nand U16055 (N_16055,N_12079,N_14831);
nand U16056 (N_16056,N_10075,N_13295);
and U16057 (N_16057,N_13426,N_13234);
nand U16058 (N_16058,N_11299,N_10169);
or U16059 (N_16059,N_14547,N_13948);
nor U16060 (N_16060,N_12741,N_12870);
or U16061 (N_16061,N_12541,N_12183);
nor U16062 (N_16062,N_12919,N_11704);
nor U16063 (N_16063,N_13048,N_12723);
nand U16064 (N_16064,N_12985,N_14646);
and U16065 (N_16065,N_12200,N_10044);
nor U16066 (N_16066,N_13024,N_14665);
nor U16067 (N_16067,N_14096,N_14478);
and U16068 (N_16068,N_13404,N_11072);
and U16069 (N_16069,N_12470,N_11743);
and U16070 (N_16070,N_14550,N_12161);
xor U16071 (N_16071,N_11043,N_11869);
nand U16072 (N_16072,N_10219,N_10512);
xor U16073 (N_16073,N_12241,N_10251);
or U16074 (N_16074,N_14609,N_10974);
xnor U16075 (N_16075,N_14806,N_13748);
nor U16076 (N_16076,N_14048,N_12852);
or U16077 (N_16077,N_10312,N_11174);
xnor U16078 (N_16078,N_12097,N_13219);
nand U16079 (N_16079,N_11570,N_10343);
nor U16080 (N_16080,N_13798,N_12173);
nor U16081 (N_16081,N_14111,N_14308);
or U16082 (N_16082,N_12126,N_10605);
nor U16083 (N_16083,N_13781,N_11682);
nand U16084 (N_16084,N_10633,N_14698);
or U16085 (N_16085,N_11650,N_13647);
or U16086 (N_16086,N_12709,N_11107);
nor U16087 (N_16087,N_13268,N_14966);
nor U16088 (N_16088,N_14222,N_11529);
and U16089 (N_16089,N_12612,N_12213);
nor U16090 (N_16090,N_12646,N_13119);
xnor U16091 (N_16091,N_11780,N_12812);
or U16092 (N_16092,N_13169,N_13380);
and U16093 (N_16093,N_10712,N_13271);
nand U16094 (N_16094,N_11524,N_13892);
nand U16095 (N_16095,N_13344,N_11335);
and U16096 (N_16096,N_11133,N_10370);
and U16097 (N_16097,N_12386,N_13848);
nand U16098 (N_16098,N_13737,N_11798);
nand U16099 (N_16099,N_10041,N_11204);
nand U16100 (N_16100,N_11787,N_11037);
nor U16101 (N_16101,N_11917,N_11716);
nor U16102 (N_16102,N_12012,N_10473);
or U16103 (N_16103,N_14620,N_10369);
nor U16104 (N_16104,N_10955,N_12275);
xnor U16105 (N_16105,N_13928,N_13236);
nand U16106 (N_16106,N_11851,N_14090);
xor U16107 (N_16107,N_11786,N_10763);
nand U16108 (N_16108,N_14343,N_10281);
or U16109 (N_16109,N_10053,N_12339);
nand U16110 (N_16110,N_12084,N_10919);
nor U16111 (N_16111,N_13355,N_12933);
xnor U16112 (N_16112,N_10614,N_12434);
or U16113 (N_16113,N_10258,N_11288);
or U16114 (N_16114,N_11352,N_12656);
and U16115 (N_16115,N_14693,N_10590);
or U16116 (N_16116,N_13712,N_12993);
and U16117 (N_16117,N_13341,N_10195);
nand U16118 (N_16118,N_14508,N_14642);
or U16119 (N_16119,N_14399,N_10694);
and U16120 (N_16120,N_14349,N_13270);
or U16121 (N_16121,N_14409,N_13217);
or U16122 (N_16122,N_12331,N_14659);
nor U16123 (N_16123,N_10252,N_10993);
and U16124 (N_16124,N_14608,N_11197);
nor U16125 (N_16125,N_14972,N_10467);
nor U16126 (N_16126,N_12240,N_10287);
nor U16127 (N_16127,N_13918,N_14796);
or U16128 (N_16128,N_13721,N_13447);
nor U16129 (N_16129,N_11802,N_11723);
nor U16130 (N_16130,N_13144,N_11635);
and U16131 (N_16131,N_13590,N_12836);
nand U16132 (N_16132,N_14772,N_10264);
nand U16133 (N_16133,N_14118,N_13659);
nand U16134 (N_16134,N_14483,N_11614);
or U16135 (N_16135,N_14058,N_12496);
nand U16136 (N_16136,N_14224,N_11854);
and U16137 (N_16137,N_14868,N_12456);
or U16138 (N_16138,N_11047,N_12251);
or U16139 (N_16139,N_12192,N_13919);
or U16140 (N_16140,N_14756,N_10789);
nor U16141 (N_16141,N_14896,N_14795);
nor U16142 (N_16142,N_10987,N_13153);
nor U16143 (N_16143,N_11567,N_13346);
and U16144 (N_16144,N_12706,N_14801);
nand U16145 (N_16145,N_13001,N_11006);
xor U16146 (N_16146,N_12621,N_11903);
nor U16147 (N_16147,N_11672,N_14367);
or U16148 (N_16148,N_12209,N_11711);
nor U16149 (N_16149,N_10726,N_10624);
xor U16150 (N_16150,N_10485,N_11582);
and U16151 (N_16151,N_12674,N_13109);
nand U16152 (N_16152,N_14158,N_14322);
and U16153 (N_16153,N_10196,N_14327);
or U16154 (N_16154,N_12043,N_12348);
or U16155 (N_16155,N_14085,N_12171);
and U16156 (N_16156,N_13331,N_10010);
nand U16157 (N_16157,N_14685,N_11226);
and U16158 (N_16158,N_12573,N_10558);
or U16159 (N_16159,N_14364,N_13349);
nor U16160 (N_16160,N_12963,N_14315);
nand U16161 (N_16161,N_14926,N_11279);
xor U16162 (N_16162,N_14143,N_12958);
xnor U16163 (N_16163,N_12680,N_12294);
xnor U16164 (N_16164,N_11103,N_12283);
or U16165 (N_16165,N_12100,N_12959);
nand U16166 (N_16166,N_10818,N_12558);
nor U16167 (N_16167,N_12046,N_13439);
nor U16168 (N_16168,N_11904,N_11915);
nand U16169 (N_16169,N_12739,N_11849);
nor U16170 (N_16170,N_10355,N_14020);
and U16171 (N_16171,N_11044,N_11880);
and U16172 (N_16172,N_11200,N_14250);
and U16173 (N_16173,N_11679,N_10105);
nor U16174 (N_16174,N_14263,N_10012);
nor U16175 (N_16175,N_10737,N_11387);
nor U16176 (N_16176,N_13038,N_14473);
or U16177 (N_16177,N_14879,N_13311);
nor U16178 (N_16178,N_13997,N_13850);
nand U16179 (N_16179,N_10218,N_13548);
and U16180 (N_16180,N_13652,N_11217);
nand U16181 (N_16181,N_11574,N_12489);
nor U16182 (N_16182,N_12300,N_10898);
and U16183 (N_16183,N_14336,N_13611);
or U16184 (N_16184,N_13786,N_10935);
or U16185 (N_16185,N_11767,N_13392);
nor U16186 (N_16186,N_12135,N_14556);
nor U16187 (N_16187,N_11724,N_12593);
and U16188 (N_16188,N_13572,N_11902);
nand U16189 (N_16189,N_12686,N_11354);
nand U16190 (N_16190,N_10427,N_14431);
or U16191 (N_16191,N_14393,N_14025);
nor U16192 (N_16192,N_14507,N_14716);
xnor U16193 (N_16193,N_14694,N_14013);
and U16194 (N_16194,N_10701,N_12098);
or U16195 (N_16195,N_10953,N_10593);
or U16196 (N_16196,N_10613,N_10089);
nor U16197 (N_16197,N_12604,N_11306);
nor U16198 (N_16198,N_14754,N_10426);
nand U16199 (N_16199,N_11648,N_10601);
and U16200 (N_16200,N_10419,N_10960);
xor U16201 (N_16201,N_14723,N_10046);
and U16202 (N_16202,N_13159,N_11140);
and U16203 (N_16203,N_11375,N_14909);
or U16204 (N_16204,N_13316,N_10668);
xnor U16205 (N_16205,N_13756,N_10509);
or U16206 (N_16206,N_14900,N_10521);
nor U16207 (N_16207,N_14166,N_11818);
and U16208 (N_16208,N_12155,N_11205);
nand U16209 (N_16209,N_14968,N_14562);
nand U16210 (N_16210,N_13163,N_13794);
and U16211 (N_16211,N_13221,N_10469);
or U16212 (N_16212,N_12316,N_13278);
and U16213 (N_16213,N_13713,N_11094);
xnor U16214 (N_16214,N_10655,N_12504);
nor U16215 (N_16215,N_13795,N_12163);
nand U16216 (N_16216,N_12537,N_12457);
or U16217 (N_16217,N_14830,N_11651);
and U16218 (N_16218,N_10446,N_10056);
nor U16219 (N_16219,N_13481,N_12120);
nor U16220 (N_16220,N_14461,N_11963);
nor U16221 (N_16221,N_13485,N_14610);
nor U16222 (N_16222,N_14663,N_10256);
nand U16223 (N_16223,N_13765,N_13461);
or U16224 (N_16224,N_12579,N_11717);
nand U16225 (N_16225,N_11984,N_10393);
and U16226 (N_16226,N_13609,N_11756);
and U16227 (N_16227,N_11348,N_10747);
nand U16228 (N_16228,N_12309,N_14195);
or U16229 (N_16229,N_13839,N_10579);
nor U16230 (N_16230,N_13610,N_12871);
and U16231 (N_16231,N_14809,N_10649);
or U16232 (N_16232,N_13549,N_10764);
nand U16233 (N_16233,N_12207,N_12802);
or U16234 (N_16234,N_11611,N_10277);
or U16235 (N_16235,N_13931,N_10121);
nor U16236 (N_16236,N_14712,N_10486);
or U16237 (N_16237,N_14657,N_13441);
nand U16238 (N_16238,N_13161,N_13056);
nor U16239 (N_16239,N_10416,N_12847);
nand U16240 (N_16240,N_13121,N_13267);
or U16241 (N_16241,N_13559,N_12119);
nand U16242 (N_16242,N_10136,N_12008);
nor U16243 (N_16243,N_12966,N_14098);
and U16244 (N_16244,N_10321,N_11752);
and U16245 (N_16245,N_10422,N_13704);
nor U16246 (N_16246,N_11231,N_13239);
and U16247 (N_16247,N_11077,N_14931);
nor U16248 (N_16248,N_12694,N_12001);
nand U16249 (N_16249,N_10806,N_11484);
nor U16250 (N_16250,N_10059,N_13770);
and U16251 (N_16251,N_12502,N_12679);
xnor U16252 (N_16252,N_11958,N_13124);
nor U16253 (N_16253,N_14722,N_12569);
and U16254 (N_16254,N_10843,N_11737);
and U16255 (N_16255,N_11382,N_12544);
nor U16256 (N_16256,N_14406,N_10625);
nand U16257 (N_16257,N_11338,N_11796);
or U16258 (N_16258,N_11312,N_13844);
xnor U16259 (N_16259,N_11932,N_11237);
nand U16260 (N_16260,N_12683,N_12841);
nor U16261 (N_16261,N_13483,N_10235);
or U16262 (N_16262,N_10745,N_12599);
xor U16263 (N_16263,N_14680,N_12533);
and U16264 (N_16264,N_10609,N_10914);
nor U16265 (N_16265,N_10409,N_12884);
or U16266 (N_16266,N_11453,N_13215);
and U16267 (N_16267,N_11602,N_12274);
nor U16268 (N_16268,N_14068,N_12223);
nand U16269 (N_16269,N_12273,N_10875);
nand U16270 (N_16270,N_12452,N_10672);
or U16271 (N_16271,N_10525,N_14018);
or U16272 (N_16272,N_10347,N_10162);
nand U16273 (N_16273,N_14176,N_12632);
nand U16274 (N_16274,N_12747,N_12530);
nand U16275 (N_16275,N_11685,N_12492);
and U16276 (N_16276,N_14576,N_14984);
or U16277 (N_16277,N_14383,N_10778);
nor U16278 (N_16278,N_14482,N_11412);
nor U16279 (N_16279,N_10684,N_11408);
and U16280 (N_16280,N_11051,N_13228);
or U16281 (N_16281,N_14426,N_12256);
or U16282 (N_16282,N_14690,N_14706);
and U16283 (N_16283,N_10723,N_13176);
and U16284 (N_16284,N_12330,N_13551);
nor U16285 (N_16285,N_13670,N_14828);
and U16286 (N_16286,N_13736,N_10606);
or U16287 (N_16287,N_11646,N_11655);
xor U16288 (N_16288,N_10699,N_10127);
nand U16289 (N_16289,N_13129,N_11182);
nor U16290 (N_16290,N_13477,N_14979);
or U16291 (N_16291,N_13705,N_13629);
and U16292 (N_16292,N_10686,N_10837);
and U16293 (N_16293,N_14387,N_14294);
nor U16294 (N_16294,N_10872,N_11879);
nand U16295 (N_16295,N_13757,N_12416);
and U16296 (N_16296,N_12877,N_14210);
and U16297 (N_16297,N_13037,N_13521);
and U16298 (N_16298,N_12344,N_13300);
and U16299 (N_16299,N_11828,N_14781);
xor U16300 (N_16300,N_11059,N_10807);
nand U16301 (N_16301,N_10420,N_12905);
or U16302 (N_16302,N_12518,N_11876);
nand U16303 (N_16303,N_14774,N_11800);
nand U16304 (N_16304,N_13925,N_11612);
nand U16305 (N_16305,N_13223,N_10353);
nor U16306 (N_16306,N_12995,N_11920);
and U16307 (N_16307,N_13419,N_14109);
and U16308 (N_16308,N_14281,N_11855);
or U16309 (N_16309,N_13568,N_11988);
or U16310 (N_16310,N_14056,N_14988);
nand U16311 (N_16311,N_13504,N_12070);
nor U16312 (N_16312,N_12840,N_12506);
or U16313 (N_16313,N_13140,N_12732);
nand U16314 (N_16314,N_13994,N_11667);
nor U16315 (N_16315,N_10144,N_10091);
and U16316 (N_16316,N_13949,N_13510);
and U16317 (N_16317,N_10350,N_14291);
nand U16318 (N_16318,N_12108,N_14155);
xnor U16319 (N_16319,N_14908,N_13552);
and U16320 (N_16320,N_11396,N_10941);
or U16321 (N_16321,N_10008,N_10386);
or U16322 (N_16322,N_14242,N_11437);
nand U16323 (N_16323,N_12654,N_11227);
or U16324 (N_16324,N_12376,N_12412);
nor U16325 (N_16325,N_10039,N_13250);
and U16326 (N_16326,N_11423,N_13902);
nand U16327 (N_16327,N_11825,N_12134);
nand U16328 (N_16328,N_10149,N_10980);
and U16329 (N_16329,N_12526,N_14891);
xor U16330 (N_16330,N_14549,N_12858);
or U16331 (N_16331,N_11616,N_13015);
or U16332 (N_16332,N_10785,N_11620);
or U16333 (N_16333,N_10635,N_13330);
and U16334 (N_16334,N_13988,N_10539);
or U16335 (N_16335,N_14216,N_13396);
nand U16336 (N_16336,N_12487,N_12915);
nand U16337 (N_16337,N_11447,N_11153);
and U16338 (N_16338,N_10130,N_12514);
xnor U16339 (N_16339,N_11819,N_13131);
and U16340 (N_16340,N_14050,N_11668);
nor U16341 (N_16341,N_11004,N_13092);
nand U16342 (N_16342,N_13791,N_13562);
or U16343 (N_16343,N_13357,N_12189);
nor U16344 (N_16344,N_14555,N_11296);
and U16345 (N_16345,N_14745,N_13399);
xnor U16346 (N_16346,N_13405,N_14607);
nor U16347 (N_16347,N_12233,N_14365);
nand U16348 (N_16348,N_13207,N_13156);
and U16349 (N_16349,N_13365,N_10518);
and U16350 (N_16350,N_12078,N_13082);
nor U16351 (N_16351,N_14518,N_14857);
nor U16352 (N_16352,N_14303,N_11432);
nand U16353 (N_16353,N_14686,N_11995);
or U16354 (N_16354,N_12006,N_10810);
nand U16355 (N_16355,N_14237,N_12215);
nor U16356 (N_16356,N_14823,N_10921);
or U16357 (N_16357,N_10248,N_12574);
nor U16358 (N_16358,N_13145,N_12984);
nor U16359 (N_16359,N_11538,N_13391);
and U16360 (N_16360,N_13725,N_13413);
or U16361 (N_16361,N_12692,N_14837);
nor U16362 (N_16362,N_10050,N_12401);
nand U16363 (N_16363,N_10610,N_12182);
and U16364 (N_16364,N_11829,N_11361);
or U16365 (N_16365,N_13754,N_11525);
or U16366 (N_16366,N_12952,N_13578);
nand U16367 (N_16367,N_12556,N_11782);
nor U16368 (N_16368,N_14771,N_12980);
nand U16369 (N_16369,N_12483,N_11536);
or U16370 (N_16370,N_11748,N_14253);
or U16371 (N_16371,N_12019,N_14527);
and U16372 (N_16372,N_13627,N_14428);
nor U16373 (N_16373,N_11757,N_14435);
and U16374 (N_16374,N_13883,N_11316);
nor U16375 (N_16375,N_11268,N_12010);
nor U16376 (N_16376,N_10177,N_11888);
nor U16377 (N_16377,N_10831,N_10632);
or U16378 (N_16378,N_10631,N_12845);
or U16379 (N_16379,N_10040,N_14702);
and U16380 (N_16380,N_10168,N_13827);
and U16381 (N_16381,N_13248,N_12572);
and U16382 (N_16382,N_14617,N_12676);
nor U16383 (N_16383,N_12407,N_14564);
nand U16384 (N_16384,N_14275,N_13623);
and U16385 (N_16385,N_12451,N_14396);
nand U16386 (N_16386,N_12026,N_11710);
and U16387 (N_16387,N_13981,N_14046);
nor U16388 (N_16388,N_11755,N_11803);
and U16389 (N_16389,N_13650,N_13273);
nand U16390 (N_16390,N_14499,N_10148);
nor U16391 (N_16391,N_11089,N_14898);
and U16392 (N_16392,N_10048,N_13177);
nand U16393 (N_16393,N_11486,N_12009);
or U16394 (N_16394,N_13057,N_13138);
and U16395 (N_16395,N_11186,N_12297);
nand U16396 (N_16396,N_13553,N_12516);
and U16397 (N_16397,N_11657,N_13784);
and U16398 (N_16398,N_12477,N_13322);
and U16399 (N_16399,N_10173,N_11603);
and U16400 (N_16400,N_14287,N_10082);
or U16401 (N_16401,N_10227,N_13367);
or U16402 (N_16402,N_14532,N_12290);
and U16403 (N_16403,N_11539,N_14429);
and U16404 (N_16404,N_11912,N_14601);
or U16405 (N_16405,N_11720,N_14838);
nor U16406 (N_16406,N_11872,N_12929);
and U16407 (N_16407,N_11224,N_13195);
xnor U16408 (N_16408,N_10803,N_14010);
or U16409 (N_16409,N_10086,N_11258);
or U16410 (N_16410,N_11134,N_13564);
nor U16411 (N_16411,N_10762,N_11906);
nand U16412 (N_16412,N_13408,N_10627);
nand U16413 (N_16413,N_11531,N_14398);
nor U16414 (N_16414,N_13921,N_10423);
and U16415 (N_16415,N_10317,N_13122);
nor U16416 (N_16416,N_10455,N_12287);
and U16417 (N_16417,N_12286,N_11609);
nor U16418 (N_16418,N_11374,N_14647);
and U16419 (N_16419,N_13849,N_13571);
or U16420 (N_16420,N_10861,N_13072);
nand U16421 (N_16421,N_14420,N_14916);
nor U16422 (N_16422,N_11322,N_13982);
and U16423 (N_16423,N_10759,N_13130);
xnor U16424 (N_16424,N_12328,N_14888);
or U16425 (N_16425,N_11455,N_11910);
and U16426 (N_16426,N_14150,N_13205);
or U16427 (N_16427,N_13895,N_10328);
nor U16428 (N_16428,N_11436,N_14852);
and U16429 (N_16429,N_12463,N_12703);
and U16430 (N_16430,N_10804,N_14065);
xnor U16431 (N_16431,N_12018,N_11403);
and U16432 (N_16432,N_11759,N_12792);
nor U16433 (N_16433,N_14368,N_10232);
nand U16434 (N_16434,N_14147,N_12790);
xor U16435 (N_16435,N_10543,N_12887);
nand U16436 (N_16436,N_14853,N_12221);
and U16437 (N_16437,N_13045,N_12873);
or U16438 (N_16438,N_10945,N_13060);
nor U16439 (N_16439,N_11990,N_11554);
and U16440 (N_16440,N_14055,N_13231);
or U16441 (N_16441,N_12391,N_13473);
nand U16442 (N_16442,N_14855,N_12693);
nor U16443 (N_16443,N_12781,N_13491);
or U16444 (N_16444,N_10940,N_10513);
xnor U16445 (N_16445,N_13961,N_12278);
xor U16446 (N_16446,N_14943,N_14304);
nand U16447 (N_16447,N_12999,N_13321);
nor U16448 (N_16448,N_13783,N_12178);
and U16449 (N_16449,N_13744,N_10589);
nand U16450 (N_16450,N_10322,N_11218);
nand U16451 (N_16451,N_13301,N_14700);
xor U16452 (N_16452,N_12440,N_13154);
nor U16453 (N_16453,N_14029,N_12333);
and U16454 (N_16454,N_10743,N_12649);
nand U16455 (N_16455,N_13378,N_10270);
nand U16456 (N_16456,N_14131,N_11214);
nor U16457 (N_16457,N_10396,N_13474);
and U16458 (N_16458,N_11501,N_10567);
nand U16459 (N_16459,N_14117,N_12616);
and U16460 (N_16460,N_14777,N_11483);
nor U16461 (N_16461,N_10933,N_10303);
and U16462 (N_16462,N_10456,N_10677);
and U16463 (N_16463,N_14282,N_14885);
or U16464 (N_16464,N_13002,N_14480);
xnor U16465 (N_16465,N_13971,N_13714);
nand U16466 (N_16466,N_14766,N_12169);
and U16467 (N_16467,N_13031,N_13790);
nor U16468 (N_16468,N_10695,N_13541);
and U16469 (N_16469,N_13010,N_10563);
xor U16470 (N_16470,N_10733,N_13517);
or U16471 (N_16471,N_12717,N_13379);
nand U16472 (N_16472,N_14681,N_12481);
nor U16473 (N_16473,N_10622,N_11419);
or U16474 (N_16474,N_10233,N_10329);
nor U16475 (N_16475,N_10878,N_12766);
and U16476 (N_16476,N_13009,N_12899);
and U16477 (N_16477,N_12203,N_10814);
nor U16478 (N_16478,N_13535,N_13135);
or U16479 (N_16479,N_13825,N_13817);
and U16480 (N_16480,N_10134,N_14705);
nor U16481 (N_16481,N_13602,N_11591);
nand U16482 (N_16482,N_11957,N_13212);
nand U16483 (N_16483,N_12264,N_13879);
or U16484 (N_16484,N_10049,N_11459);
nand U16485 (N_16485,N_11451,N_14082);
nor U16486 (N_16486,N_11130,N_10037);
xor U16487 (N_16487,N_14127,N_11376);
nor U16488 (N_16488,N_10604,N_13167);
or U16489 (N_16489,N_10798,N_14023);
nor U16490 (N_16490,N_12814,N_10979);
nor U16491 (N_16491,N_14289,N_12946);
or U16492 (N_16492,N_11896,N_11938);
nand U16493 (N_16493,N_12744,N_10477);
and U16494 (N_16494,N_14491,N_12968);
nand U16495 (N_16495,N_13907,N_10109);
or U16496 (N_16496,N_13657,N_13904);
or U16497 (N_16497,N_13034,N_12672);
xor U16498 (N_16498,N_14906,N_14091);
or U16499 (N_16499,N_11726,N_10293);
or U16500 (N_16500,N_11433,N_10124);
and U16501 (N_16501,N_10497,N_14961);
nand U16502 (N_16502,N_13165,N_11281);
nor U16503 (N_16503,N_12435,N_10461);
or U16504 (N_16504,N_13450,N_10851);
nand U16505 (N_16505,N_14776,N_12853);
and U16506 (N_16506,N_14695,N_10193);
nor U16507 (N_16507,N_13859,N_11018);
xnor U16508 (N_16508,N_10544,N_14092);
nor U16509 (N_16509,N_10670,N_12918);
nand U16510 (N_16510,N_14561,N_14615);
nor U16511 (N_16511,N_12002,N_11257);
xor U16512 (N_16512,N_12156,N_11171);
xor U16513 (N_16513,N_13327,N_14385);
nor U16514 (N_16514,N_13716,N_12320);
nor U16515 (N_16515,N_13920,N_13977);
or U16516 (N_16516,N_10275,N_10079);
or U16517 (N_16517,N_10454,N_14246);
nor U16518 (N_16518,N_10304,N_12800);
or U16519 (N_16519,N_13360,N_10228);
nor U16520 (N_16520,N_12938,N_13494);
and U16521 (N_16521,N_13641,N_10890);
xor U16522 (N_16522,N_13424,N_13133);
nand U16523 (N_16523,N_14077,N_10031);
xnor U16524 (N_16524,N_11249,N_14910);
nor U16525 (N_16525,N_11267,N_12825);
nand U16526 (N_16526,N_13958,N_11265);
or U16527 (N_16527,N_13631,N_12415);
xnor U16528 (N_16528,N_13076,N_12950);
and U16529 (N_16529,N_14528,N_14882);
nor U16530 (N_16530,N_13924,N_12110);
and U16531 (N_16531,N_13561,N_12303);
nor U16532 (N_16532,N_10595,N_10721);
and U16533 (N_16533,N_14668,N_14187);
nor U16534 (N_16534,N_11654,N_14129);
xor U16535 (N_16535,N_13533,N_11778);
nand U16536 (N_16536,N_12595,N_11864);
nor U16537 (N_16537,N_14066,N_14788);
nand U16538 (N_16538,N_14229,N_10362);
xor U16539 (N_16539,N_11874,N_11891);
nor U16540 (N_16540,N_12230,N_10179);
or U16541 (N_16541,N_13014,N_14577);
and U16542 (N_16542,N_12121,N_13209);
nand U16543 (N_16543,N_10816,N_12565);
nand U16544 (N_16544,N_13083,N_10236);
or U16545 (N_16545,N_10696,N_12381);
nand U16546 (N_16546,N_10405,N_13290);
and U16547 (N_16547,N_14474,N_11633);
or U16548 (N_16548,N_14255,N_13545);
or U16549 (N_16549,N_12104,N_13482);
or U16550 (N_16550,N_12817,N_10823);
and U16551 (N_16551,N_10880,N_10615);
and U16552 (N_16552,N_12282,N_12436);
and U16553 (N_16553,N_10499,N_14113);
and U16554 (N_16554,N_13939,N_13546);
and U16555 (N_16555,N_11232,N_13942);
nor U16556 (N_16556,N_10962,N_14752);
nand U16557 (N_16557,N_12819,N_11641);
or U16558 (N_16558,N_14579,N_14119);
nand U16559 (N_16559,N_14203,N_11661);
nand U16560 (N_16560,N_12159,N_13854);
nor U16561 (N_16561,N_12343,N_14724);
nand U16562 (N_16562,N_11398,N_14233);
and U16563 (N_16563,N_12910,N_10459);
or U16564 (N_16564,N_14440,N_11821);
nand U16565 (N_16565,N_12352,N_10886);
nand U16566 (N_16566,N_14257,N_10596);
nand U16567 (N_16567,N_13403,N_11458);
and U16568 (N_16568,N_12247,N_10838);
xor U16569 (N_16569,N_12319,N_11126);
and U16570 (N_16570,N_13149,N_12280);
and U16571 (N_16571,N_12746,N_14918);
nor U16572 (N_16572,N_10245,N_11866);
and U16573 (N_16573,N_11090,N_12754);
and U16574 (N_16574,N_14284,N_12039);
xor U16575 (N_16575,N_13773,N_11553);
nand U16576 (N_16576,N_12065,N_14376);
nand U16577 (N_16577,N_12427,N_14070);
nand U16578 (N_16578,N_13583,N_11095);
and U16579 (N_16579,N_10847,N_13589);
or U16580 (N_16580,N_13695,N_10051);
nor U16581 (N_16581,N_11550,N_12917);
nor U16582 (N_16582,N_12886,N_12614);
and U16583 (N_16583,N_14902,N_13328);
or U16584 (N_16584,N_10495,N_11488);
or U16585 (N_16585,N_10648,N_10138);
or U16586 (N_16586,N_12975,N_11054);
or U16587 (N_16587,N_10057,N_14441);
nor U16588 (N_16588,N_13196,N_11783);
nand U16589 (N_16589,N_11427,N_14403);
nand U16590 (N_16590,N_12217,N_12517);
nand U16591 (N_16591,N_13047,N_11762);
or U16592 (N_16592,N_10468,N_12749);
or U16593 (N_16593,N_10508,N_10994);
nand U16594 (N_16594,N_14503,N_12270);
and U16595 (N_16595,N_11156,N_12684);
and U16596 (N_16596,N_11115,N_12522);
and U16597 (N_16597,N_10949,N_14911);
xor U16598 (N_16598,N_10800,N_12563);
and U16599 (N_16599,N_14290,N_14313);
nor U16600 (N_16600,N_10061,N_12304);
and U16601 (N_16601,N_13495,N_10207);
nor U16602 (N_16602,N_11527,N_13418);
or U16603 (N_16603,N_10771,N_13878);
xor U16604 (N_16604,N_10881,N_14894);
and U16605 (N_16605,N_14347,N_13454);
nor U16606 (N_16606,N_12438,N_13978);
or U16607 (N_16607,N_14779,N_12363);
nand U16608 (N_16608,N_10118,N_14613);
nor U16609 (N_16609,N_11293,N_14636);
xnor U16610 (N_16610,N_14960,N_11532);
nand U16611 (N_16611,N_11734,N_13443);
nor U16612 (N_16612,N_12131,N_13071);
and U16613 (N_16613,N_12257,N_11421);
and U16614 (N_16614,N_12945,N_14350);
and U16615 (N_16615,N_12865,N_11343);
nor U16616 (N_16616,N_14995,N_10906);
xor U16617 (N_16617,N_10160,N_12114);
or U16618 (N_16618,N_14439,N_13067);
nor U16619 (N_16619,N_13941,N_12293);
nor U16620 (N_16620,N_14358,N_14510);
nor U16621 (N_16621,N_12364,N_10557);
xor U16622 (N_16622,N_11569,N_13901);
and U16623 (N_16623,N_11781,N_11008);
or U16624 (N_16624,N_10582,N_14953);
nor U16625 (N_16625,N_12986,N_12340);
and U16626 (N_16626,N_14137,N_10345);
nand U16627 (N_16627,N_14614,N_12088);
or U16628 (N_16628,N_10839,N_11386);
nor U16629 (N_16629,N_12050,N_11804);
or U16630 (N_16630,N_12577,N_14477);
xnor U16631 (N_16631,N_14481,N_14054);
xor U16632 (N_16632,N_14377,N_14204);
nand U16633 (N_16633,N_13183,N_14252);
and U16634 (N_16634,N_13799,N_12860);
and U16635 (N_16635,N_12822,N_14849);
nand U16636 (N_16636,N_11471,N_13241);
or U16637 (N_16637,N_13113,N_12327);
nand U16638 (N_16638,N_11303,N_12644);
nand U16639 (N_16639,N_11557,N_10022);
nor U16640 (N_16640,N_10309,N_12311);
and U16641 (N_16641,N_14903,N_11309);
nor U16642 (N_16642,N_10922,N_14084);
nand U16643 (N_16643,N_13842,N_13304);
nand U16644 (N_16644,N_11160,N_14254);
and U16645 (N_16645,N_10553,N_10825);
xnor U16646 (N_16646,N_13634,N_12738);
or U16647 (N_16647,N_13796,N_10966);
xnor U16648 (N_16648,N_10255,N_11157);
xnor U16649 (N_16649,N_13654,N_10064);
and U16650 (N_16650,N_13319,N_11357);
nand U16651 (N_16651,N_10538,N_13675);
nand U16652 (N_16652,N_14069,N_10664);
or U16653 (N_16653,N_14586,N_10171);
nand U16654 (N_16654,N_11046,N_13830);
and U16655 (N_16655,N_12623,N_12737);
nor U16656 (N_16656,N_13645,N_12379);
nand U16657 (N_16657,N_12279,N_13148);
nor U16658 (N_16658,N_14163,N_11508);
xnor U16659 (N_16659,N_14202,N_11148);
or U16660 (N_16660,N_14100,N_13007);
or U16661 (N_16661,N_13340,N_12444);
and U16662 (N_16662,N_14273,N_14183);
nor U16663 (N_16663,N_12229,N_12338);
nand U16664 (N_16664,N_12498,N_13411);
nor U16665 (N_16665,N_13036,N_14845);
xnor U16666 (N_16666,N_11492,N_14209);
or U16667 (N_16667,N_12642,N_11428);
nor U16668 (N_16668,N_13111,N_10799);
nor U16669 (N_16669,N_10324,N_12334);
nor U16670 (N_16670,N_12380,N_12885);
nand U16671 (N_16671,N_11394,N_10536);
nor U16672 (N_16672,N_11500,N_12727);
or U16673 (N_16673,N_11195,N_12677);
nand U16674 (N_16674,N_13118,N_12708);
xnor U16675 (N_16675,N_11714,N_14261);
nor U16676 (N_16676,N_10597,N_13497);
and U16677 (N_16677,N_10690,N_14251);
nand U16678 (N_16678,N_14817,N_14205);
and U16679 (N_16679,N_12218,N_12967);
and U16680 (N_16680,N_12925,N_11749);
or U16681 (N_16681,N_14987,N_13400);
and U16682 (N_16682,N_13788,N_10551);
and U16683 (N_16683,N_11931,N_11401);
nand U16684 (N_16684,N_11496,N_12875);
nor U16685 (N_16685,N_12423,N_10537);
nor U16686 (N_16686,N_14672,N_12296);
nand U16687 (N_16687,N_12004,N_12844);
nand U16688 (N_16688,N_13860,N_13995);
nand U16689 (N_16689,N_12058,N_14352);
nor U16690 (N_16690,N_14675,N_13087);
and U16691 (N_16691,N_10385,N_12936);
nand U16692 (N_16692,N_13137,N_10549);
xnor U16693 (N_16693,N_12357,N_12260);
nor U16694 (N_16694,N_13351,N_13852);
nor U16695 (N_16695,N_13061,N_12903);
nand U16696 (N_16696,N_11342,N_13274);
xnor U16697 (N_16697,N_12158,N_10791);
or U16698 (N_16698,N_12437,N_12803);
nand U16699 (N_16699,N_10133,N_10301);
nor U16700 (N_16700,N_12846,N_13986);
nand U16701 (N_16701,N_10371,N_12926);
nand U16702 (N_16702,N_12901,N_13819);
nand U16703 (N_16703,N_14948,N_12699);
xnor U16704 (N_16704,N_13286,N_14818);
nand U16705 (N_16705,N_11656,N_10280);
nor U16706 (N_16706,N_14760,N_14717);
and U16707 (N_16707,N_10780,N_12813);
nor U16708 (N_16708,N_11973,N_14662);
nor U16709 (N_16709,N_12160,N_13900);
nand U16710 (N_16710,N_11847,N_13976);
and U16711 (N_16711,N_13745,N_10689);
or U16712 (N_16712,N_10584,N_10948);
xnor U16713 (N_16713,N_11929,N_13665);
or U16714 (N_16714,N_13440,N_11537);
and U16715 (N_16715,N_12288,N_14514);
or U16716 (N_16716,N_12038,N_10361);
nand U16717 (N_16717,N_11882,N_12281);
and U16718 (N_16718,N_12028,N_11729);
or U16719 (N_16719,N_13224,N_14667);
or U16720 (N_16720,N_14734,N_13464);
nor U16721 (N_16721,N_14677,N_12507);
nor U16722 (N_16722,N_10665,N_11922);
or U16723 (N_16723,N_10339,N_10724);
and U16724 (N_16724,N_14950,N_10414);
and U16725 (N_16725,N_11506,N_10903);
xnor U16726 (N_16726,N_13628,N_12164);
nand U16727 (N_16727,N_12245,N_12382);
or U16728 (N_16728,N_14286,N_11513);
nand U16729 (N_16729,N_14356,N_13673);
nor U16730 (N_16730,N_10598,N_11914);
xor U16731 (N_16731,N_12897,N_11730);
or U16732 (N_16732,N_13100,N_10853);
nor U16733 (N_16733,N_14234,N_10378);
nor U16734 (N_16734,N_11031,N_13376);
nor U16735 (N_16735,N_11284,N_11860);
xnor U16736 (N_16736,N_14296,N_11263);
and U16737 (N_16737,N_11228,N_13046);
nand U16738 (N_16738,N_12335,N_10388);
nand U16739 (N_16739,N_12794,N_11332);
and U16740 (N_16740,N_11183,N_13289);
nor U16741 (N_16741,N_11201,N_14007);
xor U16742 (N_16742,N_10375,N_10492);
or U16743 (N_16743,N_11324,N_14353);
and U16744 (N_16744,N_10917,N_13178);
xor U16745 (N_16745,N_10616,N_14244);
xnor U16746 (N_16746,N_14794,N_11699);
xnor U16747 (N_16747,N_14330,N_10836);
nor U16748 (N_16748,N_11219,N_11395);
or U16749 (N_16749,N_14310,N_13353);
nor U16750 (N_16750,N_14332,N_11950);
nand U16751 (N_16751,N_13035,N_13078);
and U16752 (N_16752,N_14741,N_13523);
xnor U16753 (N_16753,N_14640,N_11725);
nand U16754 (N_16754,N_11275,N_13390);
and U16755 (N_16755,N_11093,N_12510);
nand U16756 (N_16756,N_13085,N_13369);
nand U16757 (N_16757,N_12271,N_10654);
xnor U16758 (N_16758,N_10116,N_12265);
and U16759 (N_16759,N_10308,N_11198);
xnor U16760 (N_16760,N_12989,N_11135);
or U16761 (N_16761,N_13345,N_10970);
and U16762 (N_16762,N_12405,N_14469);
nor U16763 (N_16763,N_10216,N_13229);
nand U16764 (N_16764,N_12710,N_13728);
nand U16765 (N_16765,N_12460,N_10440);
or U16766 (N_16766,N_11588,N_12393);
and U16767 (N_16767,N_14348,N_11066);
nand U16768 (N_16768,N_14839,N_13822);
nand U16769 (N_16769,N_13125,N_10365);
or U16770 (N_16770,N_10772,N_11715);
nor U16771 (N_16771,N_14338,N_12590);
and U16772 (N_16772,N_14489,N_14844);
nor U16773 (N_16773,N_14848,N_13812);
nor U16774 (N_16774,N_12535,N_11568);
nor U16775 (N_16775,N_11843,N_10387);
nand U16776 (N_16776,N_13896,N_11639);
and U16777 (N_16777,N_14656,N_11141);
nor U16778 (N_16778,N_13821,N_12725);
and U16779 (N_16779,N_12377,N_10583);
or U16780 (N_16780,N_13102,N_12911);
or U16781 (N_16781,N_12326,N_10319);
nand U16782 (N_16782,N_11210,N_11172);
nand U16783 (N_16783,N_14581,N_11320);
or U16784 (N_16784,N_14634,N_14394);
nand U16785 (N_16785,N_10310,N_10132);
and U16786 (N_16786,N_12349,N_14016);
nand U16787 (N_16787,N_13932,N_11846);
nand U16788 (N_16788,N_11429,N_12752);
and U16789 (N_16789,N_14277,N_13252);
xor U16790 (N_16790,N_14404,N_10289);
nor U16791 (N_16791,N_10578,N_12124);
and U16792 (N_16792,N_10351,N_12167);
or U16793 (N_16793,N_12059,N_14094);
xnor U16794 (N_16794,N_13147,N_12711);
nand U16795 (N_16795,N_14521,N_11691);
nor U16796 (N_16796,N_10458,N_14599);
and U16797 (N_16797,N_12495,N_13117);
nand U16798 (N_16798,N_11997,N_14920);
nand U16799 (N_16799,N_13577,N_13005);
xor U16800 (N_16800,N_14710,N_10937);
nor U16801 (N_16801,N_13702,N_12151);
and U16802 (N_16802,N_12298,N_14189);
and U16803 (N_16803,N_12125,N_13180);
nor U16804 (N_16804,N_10656,N_14033);
or U16805 (N_16805,N_14384,N_10977);
or U16806 (N_16806,N_10249,N_13536);
or U16807 (N_16807,N_10907,N_12772);
nor U16808 (N_16808,N_13480,N_14190);
nor U16809 (N_16809,N_13567,N_14993);
and U16810 (N_16810,N_10363,N_13674);
or U16811 (N_16811,N_11191,N_12048);
nor U16812 (N_16812,N_10032,N_12366);
nor U16813 (N_16813,N_13158,N_14139);
nor U16814 (N_16814,N_14708,N_12152);
nand U16815 (N_16815,N_12855,N_12742);
or U16816 (N_16816,N_10653,N_14392);
and U16817 (N_16817,N_10215,N_13394);
nor U16818 (N_16818,N_14649,N_11937);
or U16819 (N_16819,N_10683,N_11674);
or U16820 (N_16820,N_10334,N_11173);
nor U16821 (N_16821,N_12992,N_12625);
and U16822 (N_16822,N_11168,N_14921);
or U16823 (N_16823,N_11683,N_10221);
nand U16824 (N_16824,N_12962,N_10211);
nor U16825 (N_16825,N_12815,N_14087);
or U16826 (N_16826,N_11887,N_10857);
nor U16827 (N_16827,N_10030,N_13222);
nor U16828 (N_16828,N_14124,N_10548);
nand U16829 (N_16829,N_10282,N_12305);
nor U16830 (N_16830,N_10731,N_14881);
nand U16831 (N_16831,N_14357,N_14583);
nand U16832 (N_16832,N_10418,N_14790);
nand U16833 (N_16833,N_11070,N_14427);
or U16834 (N_16834,N_11707,N_10944);
or U16835 (N_16835,N_13749,N_12705);
or U16836 (N_16836,N_10675,N_12361);
or U16837 (N_16837,N_12371,N_12147);
and U16838 (N_16838,N_10223,N_10294);
or U16839 (N_16839,N_10146,N_14043);
and U16840 (N_16840,N_14081,N_10722);
and U16841 (N_16841,N_11102,N_13964);
nor U16842 (N_16842,N_13160,N_13334);
and U16843 (N_16843,N_12204,N_13658);
nor U16844 (N_16844,N_10796,N_10926);
or U16845 (N_16845,N_14638,N_13173);
or U16846 (N_16846,N_11479,N_12289);
or U16847 (N_16847,N_12208,N_10884);
nand U16848 (N_16848,N_14800,N_14560);
and U16849 (N_16849,N_12362,N_12820);
or U16850 (N_16850,N_10517,N_11071);
or U16851 (N_16851,N_10163,N_14432);
and U16852 (N_16852,N_12052,N_12047);
xor U16853 (N_16853,N_11491,N_13557);
nand U16854 (N_16854,N_10946,N_12022);
and U16855 (N_16855,N_13579,N_10752);
or U16856 (N_16856,N_14524,N_11082);
or U16857 (N_16857,N_13469,N_14316);
nand U16858 (N_16858,N_14260,N_11121);
nor U16859 (N_16859,N_14737,N_10900);
nor U16860 (N_16860,N_10756,N_11623);
nand U16861 (N_16861,N_11634,N_12252);
xnor U16862 (N_16862,N_13412,N_10152);
nand U16863 (N_16863,N_14892,N_13669);
and U16864 (N_16864,N_12027,N_11595);
and U16865 (N_16865,N_10591,N_12388);
nor U16866 (N_16866,N_13025,N_11861);
or U16867 (N_16867,N_12922,N_12805);
nand U16868 (N_16868,N_11104,N_10379);
nor U16869 (N_16869,N_10829,N_12013);
nand U16870 (N_16870,N_12237,N_13033);
or U16871 (N_16871,N_11016,N_14230);
nand U16872 (N_16872,N_11728,N_13870);
xor U16873 (N_16873,N_12582,N_11466);
nand U16874 (N_16874,N_12246,N_12137);
and U16875 (N_16875,N_12872,N_11878);
or U16876 (N_16876,N_11449,N_10430);
and U16877 (N_16877,N_12116,N_13256);
xnor U16878 (N_16878,N_11926,N_14247);
xor U16879 (N_16879,N_10297,N_13780);
nand U16880 (N_16880,N_12628,N_11746);
or U16881 (N_16881,N_12743,N_13442);
nand U16882 (N_16882,N_11470,N_11600);
nor U16883 (N_16883,N_11243,N_13128);
and U16884 (N_16884,N_11696,N_13194);
and U16885 (N_16885,N_14307,N_14370);
nor U16886 (N_16886,N_10098,N_12323);
or U16887 (N_16887,N_10873,N_11630);
or U16888 (N_16888,N_14725,N_11573);
or U16889 (N_16889,N_11271,N_12571);
or U16890 (N_16890,N_11125,N_10927);
and U16891 (N_16891,N_11314,N_11766);
xnor U16892 (N_16892,N_13174,N_13649);
nor U16893 (N_16893,N_12536,N_14585);
nor U16894 (N_16894,N_12673,N_11826);
nand U16895 (N_16895,N_13563,N_10052);
nor U16896 (N_16896,N_13671,N_13170);
xor U16897 (N_16897,N_11391,N_13188);
xor U16898 (N_16898,N_12603,N_11502);
nand U16899 (N_16899,N_11919,N_10333);
xnor U16900 (N_16900,N_10230,N_14684);
or U16901 (N_16901,N_13030,N_11747);
and U16902 (N_16902,N_14345,N_12430);
and U16903 (N_16903,N_13068,N_13101);
and U16904 (N_16904,N_14022,N_12981);
nand U16905 (N_16905,N_10011,N_11443);
nand U16906 (N_16906,N_10018,N_14506);
or U16907 (N_16907,N_12299,N_11621);
nor U16908 (N_16908,N_13730,N_14164);
nor U16909 (N_16909,N_14037,N_12650);
and U16910 (N_16910,N_13573,N_14568);
nand U16911 (N_16911,N_12458,N_10147);
nor U16912 (N_16912,N_12113,N_12972);
and U16913 (N_16913,N_13051,N_13040);
xor U16914 (N_16914,N_12336,N_11863);
xor U16915 (N_16915,N_14616,N_12515);
nand U16916 (N_16916,N_12580,N_14279);
nand U16917 (N_16917,N_13889,N_13383);
nor U16918 (N_16918,N_13164,N_13332);
nor U16919 (N_16919,N_11397,N_13247);
nand U16920 (N_16920,N_14955,N_13338);
or U16921 (N_16921,N_10936,N_11239);
or U16922 (N_16922,N_11510,N_14947);
nand U16923 (N_16923,N_14875,N_11558);
and U16924 (N_16924,N_13775,N_10107);
and U16925 (N_16925,N_11149,N_11468);
nor U16926 (N_16926,N_14141,N_14182);
xor U16927 (N_16927,N_10892,N_11469);
nor U16928 (N_16928,N_14444,N_13027);
and U16929 (N_16929,N_11969,N_11599);
or U16930 (N_16930,N_13370,N_10267);
nor U16931 (N_16931,N_11792,N_11797);
xor U16932 (N_16932,N_10391,N_11380);
xor U16933 (N_16933,N_14990,N_14573);
nand U16934 (N_16934,N_10023,N_10069);
and U16935 (N_16935,N_13679,N_14986);
or U16936 (N_16936,N_14321,N_10895);
nor U16937 (N_16937,N_11294,N_11367);
nand U16938 (N_16938,N_13857,N_11057);
nor U16939 (N_16939,N_12306,N_14463);
xor U16940 (N_16940,N_12721,N_14292);
or U16941 (N_16941,N_11311,N_10996);
nand U16942 (N_16942,N_11509,N_10180);
and U16943 (N_16943,N_11109,N_11601);
nand U16944 (N_16944,N_14470,N_14051);
and U16945 (N_16945,N_14436,N_11234);
nor U16946 (N_16946,N_12778,N_13094);
nand U16947 (N_16947,N_12387,N_13835);
and U16948 (N_16948,N_13668,N_12089);
and U16949 (N_16949,N_12682,N_13050);
nand U16950 (N_16950,N_10119,N_10253);
and U16951 (N_16951,N_10698,N_14994);
xnor U16952 (N_16952,N_11425,N_12971);
and U16953 (N_16953,N_12312,N_13782);
nand U16954 (N_16954,N_13023,N_13701);
or U16955 (N_16955,N_13065,N_12115);
xnor U16956 (N_16956,N_14825,N_12639);
and U16957 (N_16957,N_10607,N_10889);
nor U16958 (N_16958,N_14758,N_13954);
nand U16959 (N_16959,N_11328,N_11627);
or U16960 (N_16960,N_10108,N_10533);
nor U16961 (N_16961,N_11512,N_12588);
nand U16962 (N_16962,N_10805,N_14211);
and U16963 (N_16963,N_14567,N_14041);
xor U16964 (N_16964,N_10812,N_13616);
nand U16965 (N_16965,N_12146,N_14397);
and U16966 (N_16966,N_13096,N_11671);
and U16967 (N_16967,N_11626,N_13813);
and U16968 (N_16968,N_12074,N_12857);
xor U16969 (N_16969,N_12769,N_13105);
and U16970 (N_16970,N_11960,N_12828);
or U16971 (N_16971,N_12801,N_12499);
nand U16972 (N_16972,N_12608,N_13368);
nor U16973 (N_16973,N_14331,N_13984);
nor U16974 (N_16974,N_10667,N_14932);
or U16975 (N_16975,N_13272,N_12687);
and U16976 (N_16976,N_12876,N_12396);
nand U16977 (N_16977,N_14468,N_12034);
nor U16978 (N_16978,N_10166,N_14720);
nor U16979 (N_16979,N_13893,N_10155);
or U16980 (N_16980,N_13717,N_12786);
and U16981 (N_16981,N_10983,N_10715);
nand U16982 (N_16982,N_12332,N_10093);
or U16983 (N_16983,N_12360,N_14719);
and U16984 (N_16984,N_14062,N_13838);
or U16985 (N_16985,N_10239,N_13069);
nand U16986 (N_16986,N_12190,N_14750);
nor U16987 (N_16987,N_12645,N_10209);
and U16988 (N_16988,N_10263,N_14517);
or U16989 (N_16989,N_14160,N_12835);
xnor U16990 (N_16990,N_10620,N_14101);
nor U16991 (N_16991,N_14437,N_13706);
or U16992 (N_16992,N_14936,N_14112);
or U16993 (N_16993,N_10988,N_11476);
and U16994 (N_16994,N_12149,N_10998);
and U16995 (N_16995,N_12659,N_14683);
nor U16996 (N_16996,N_14833,N_14618);
and U16997 (N_16997,N_12991,N_11384);
nand U16998 (N_16998,N_14739,N_13395);
nor U16999 (N_16999,N_12035,N_13877);
nand U17000 (N_17000,N_11297,N_10327);
and U17001 (N_17001,N_12449,N_14319);
or U17002 (N_17002,N_14923,N_10104);
nand U17003 (N_17003,N_10262,N_13320);
nand U17004 (N_17004,N_12468,N_12029);
xor U17005 (N_17005,N_14873,N_11515);
or U17006 (N_17006,N_12770,N_11753);
xor U17007 (N_17007,N_10773,N_12353);
nand U17008 (N_17008,N_10808,N_10770);
nand U17009 (N_17009,N_12179,N_14419);
nor U17010 (N_17010,N_10532,N_12093);
and U17011 (N_17011,N_11833,N_10714);
or U17012 (N_17012,N_14132,N_14328);
and U17013 (N_17013,N_13952,N_11867);
nand U17014 (N_17014,N_13752,N_11647);
nor U17015 (N_17015,N_11758,N_12653);
nor U17016 (N_17016,N_13216,N_10958);
nor U17017 (N_17017,N_14285,N_10828);
or U17018 (N_17018,N_10247,N_12635);
and U17019 (N_17019,N_13511,N_13620);
nor U17020 (N_17020,N_11992,N_11572);
xor U17021 (N_17021,N_11681,N_12142);
or U17022 (N_17022,N_14201,N_11928);
nor U17023 (N_17023,N_13466,N_14807);
xor U17024 (N_17024,N_13226,N_11664);
nor U17025 (N_17025,N_13899,N_10559);
nand U17026 (N_17026,N_12291,N_13265);
and U17027 (N_17027,N_12123,N_13249);
nand U17028 (N_17028,N_11270,N_11875);
nor U17029 (N_17029,N_12597,N_11976);
or U17030 (N_17030,N_10226,N_14699);
nor U17031 (N_17031,N_12473,N_11402);
nor U17032 (N_17032,N_10918,N_12513);
xor U17033 (N_17033,N_12823,N_10153);
and U17034 (N_17034,N_13382,N_13797);
nor U17035 (N_17035,N_11868,N_13110);
and U17036 (N_17036,N_13008,N_14566);
or U17037 (N_17037,N_12818,N_10515);
nor U17038 (N_17038,N_13366,N_12465);
nand U17039 (N_17039,N_10923,N_13764);
and U17040 (N_17040,N_13580,N_11242);
nand U17041 (N_17041,N_10066,N_12277);
nand U17042 (N_17042,N_10175,N_10844);
or U17043 (N_17043,N_14594,N_13296);
and U17044 (N_17044,N_11122,N_14239);
or U17045 (N_17045,N_11625,N_11050);
or U17046 (N_17046,N_10519,N_14105);
xnor U17047 (N_17047,N_11155,N_10433);
and U17048 (N_17048,N_10775,N_12806);
nand U17049 (N_17049,N_12660,N_13792);
and U17050 (N_17050,N_13569,N_14558);
or U17051 (N_17051,N_14448,N_11881);
or U17052 (N_17052,N_13787,N_13081);
and U17053 (N_17053,N_10198,N_12446);
nand U17054 (N_17054,N_14846,N_14496);
nand U17055 (N_17055,N_13064,N_11215);
nand U17056 (N_17056,N_14804,N_12949);
nor U17057 (N_17057,N_13708,N_10176);
or U17058 (N_17058,N_14942,N_12196);
nor U17059 (N_17059,N_10863,N_10117);
or U17060 (N_17060,N_13688,N_14271);
and U17061 (N_17061,N_14060,N_13325);
nand U17062 (N_17062,N_11772,N_10813);
and U17063 (N_17063,N_11744,N_10599);
nand U17064 (N_17064,N_12890,N_13597);
nand U17065 (N_17065,N_14670,N_10206);
nand U17066 (N_17066,N_11946,N_14516);
and U17067 (N_17067,N_10732,N_13246);
nor U17068 (N_17068,N_14381,N_13973);
or U17069 (N_17069,N_11564,N_13018);
and U17070 (N_17070,N_10534,N_10298);
nor U17071 (N_17071,N_12787,N_11768);
xnor U17072 (N_17072,N_14363,N_12138);
or U17073 (N_17073,N_12136,N_14199);
and U17074 (N_17074,N_14814,N_10908);
nand U17075 (N_17075,N_12197,N_13722);
nand U17076 (N_17076,N_10143,N_12907);
nand U17077 (N_17077,N_14344,N_10973);
and U17078 (N_17078,N_14829,N_10213);
and U17079 (N_17079,N_12581,N_12883);
nand U17080 (N_17080,N_14306,N_13600);
or U17081 (N_17081,N_10503,N_10528);
nand U17082 (N_17082,N_14361,N_11026);
and U17083 (N_17083,N_11353,N_10742);
or U17084 (N_17084,N_11150,N_14288);
or U17085 (N_17085,N_10192,N_11452);
or U17086 (N_17086,N_12630,N_10489);
and U17087 (N_17087,N_14390,N_11388);
or U17088 (N_17088,N_11959,N_12040);
or U17089 (N_17089,N_12354,N_14759);
nor U17090 (N_17090,N_11662,N_14643);
or U17091 (N_17091,N_11475,N_13022);
or U17092 (N_17092,N_13855,N_11951);
and U17093 (N_17093,N_10435,N_11751);
and U17094 (N_17094,N_11266,N_13655);
nand U17095 (N_17095,N_11088,N_14146);
or U17096 (N_17096,N_14637,N_10947);
nand U17097 (N_17097,N_13496,N_10754);
nor U17098 (N_17098,N_10932,N_10864);
or U17099 (N_17099,N_11848,N_11930);
nor U17100 (N_17100,N_10028,N_14157);
xnor U17101 (N_17101,N_13876,N_12244);
or U17102 (N_17102,N_11344,N_12779);
nor U17103 (N_17103,N_11165,N_12955);
nor U17104 (N_17104,N_13302,N_10316);
and U17105 (N_17105,N_13703,N_12443);
nor U17106 (N_17106,N_10342,N_10651);
xor U17107 (N_17107,N_14537,N_13314);
or U17108 (N_17108,N_10899,N_10758);
nor U17109 (N_17109,N_10735,N_14415);
xor U17110 (N_17110,N_10437,N_10128);
or U17111 (N_17111,N_13805,N_11456);
nand U17112 (N_17112,N_12796,N_10950);
nor U17113 (N_17113,N_13233,N_11886);
nor U17114 (N_17114,N_12153,N_11511);
nand U17115 (N_17115,N_11145,N_14835);
and U17116 (N_17116,N_10760,N_10905);
nand U17117 (N_17117,N_14652,N_11649);
or U17118 (N_17118,N_12774,N_12375);
or U17119 (N_17119,N_14786,N_14808);
or U17120 (N_17120,N_12228,N_11063);
or U17121 (N_17121,N_13707,N_10481);
nand U17122 (N_17122,N_10071,N_11731);
nor U17123 (N_17123,N_12540,N_14696);
and U17124 (N_17124,N_13913,N_13213);
nor U17125 (N_17125,N_14447,N_11530);
nand U17126 (N_17126,N_14691,N_10271);
and U17127 (N_17127,N_14262,N_13833);
nor U17128 (N_17128,N_12345,N_10777);
nor U17129 (N_17129,N_13653,N_10421);
nor U17130 (N_17130,N_11581,N_13417);
and U17131 (N_17131,N_13315,N_11807);
nor U17132 (N_17132,N_12554,N_14359);
nor U17133 (N_17133,N_14784,N_11223);
or U17134 (N_17134,N_10850,N_14827);
and U17135 (N_17135,N_12253,N_11812);
and U17136 (N_17136,N_12987,N_14520);
and U17137 (N_17137,N_14039,N_14047);
nor U17138 (N_17138,N_10186,N_10592);
nor U17139 (N_17139,N_14744,N_10276);
and U17140 (N_17140,N_13032,N_11516);
nor U17141 (N_17141,N_10191,N_13339);
or U17142 (N_17142,N_12220,N_11617);
or U17143 (N_17143,N_14731,N_11836);
nand U17144 (N_17144,N_11949,N_14515);
or U17145 (N_17145,N_10217,N_11586);
or U17146 (N_17146,N_10611,N_11313);
nor U17147 (N_17147,N_14053,N_12187);
nand U17148 (N_17148,N_10546,N_12634);
nand U17149 (N_17149,N_13171,N_14999);
xnor U17150 (N_17150,N_14701,N_10331);
nor U17151 (N_17151,N_10401,N_12667);
xor U17152 (N_17152,N_10340,N_13487);
nand U17153 (N_17153,N_11528,N_14148);
xor U17154 (N_17154,N_13956,N_12454);
nand U17155 (N_17155,N_11481,N_13594);
nor U17156 (N_17156,N_10407,N_14963);
nor U17157 (N_17157,N_10560,N_13866);
or U17158 (N_17158,N_14629,N_13507);
and U17159 (N_17159,N_10306,N_14651);
nand U17160 (N_17160,N_14421,N_10244);
and U17161 (N_17161,N_10372,N_12661);
or U17162 (N_17162,N_11842,N_10912);
nand U17163 (N_17163,N_12165,N_12177);
and U17164 (N_17164,N_10237,N_11022);
or U17165 (N_17165,N_11467,N_11295);
nand U17166 (N_17166,N_14736,N_14726);
or U17167 (N_17167,N_12024,N_11278);
nor U17168 (N_17168,N_10761,N_10013);
and U17169 (N_17169,N_10078,N_14820);
nor U17170 (N_17170,N_11464,N_10692);
and U17171 (N_17171,N_14939,N_11283);
or U17172 (N_17172,N_14373,N_14180);
xor U17173 (N_17173,N_14418,N_10986);
or U17174 (N_17174,N_14326,N_10110);
nand U17175 (N_17175,N_12411,N_14140);
nor U17176 (N_17176,N_12691,N_12478);
nor U17177 (N_17177,N_12181,N_12862);
nand U17178 (N_17178,N_12939,N_10634);
nand U17179 (N_17179,N_13152,N_12748);
or U17180 (N_17180,N_13444,N_12589);
and U17181 (N_17181,N_10034,N_12859);
nor U17182 (N_17182,N_14462,N_10781);
or U17183 (N_17183,N_12602,N_12106);
xor U17184 (N_17184,N_12696,N_13053);
or U17185 (N_17185,N_10913,N_11640);
nand U17186 (N_17186,N_13720,N_12342);
and U17187 (N_17187,N_13099,N_13980);
nor U17188 (N_17188,N_13303,N_11618);
xor U17189 (N_17189,N_10660,N_13358);
and U17190 (N_17190,N_14762,N_14302);
and U17191 (N_17191,N_14778,N_12439);
nor U17192 (N_17192,N_10555,N_14335);
or U17193 (N_17193,N_11993,N_14631);
and U17194 (N_17194,N_14782,N_10978);
nand U17195 (N_17195,N_13336,N_12015);
nand U17196 (N_17196,N_13043,N_11596);
nor U17197 (N_17197,N_13944,N_10250);
nand U17198 (N_17198,N_11323,N_11142);
or U17199 (N_17199,N_12973,N_12005);
nor U17200 (N_17200,N_12337,N_10336);
and U17201 (N_17201,N_12542,N_13742);
nor U17202 (N_17202,N_13435,N_14965);
nor U17203 (N_17203,N_10883,N_13416);
or U17204 (N_17204,N_12250,N_11379);
nand U17205 (N_17205,N_12356,N_11972);
and U17206 (N_17206,N_11287,N_14240);
nand U17207 (N_17207,N_11351,N_14133);
or U17208 (N_17208,N_10141,N_13039);
nor U17209 (N_17209,N_14904,N_11556);
or U17210 (N_17210,N_10188,N_14194);
or U17211 (N_17211,N_14856,N_14325);
nor U17212 (N_17212,N_13350,N_11764);
nand U17213 (N_17213,N_11282,N_14733);
nor U17214 (N_17214,N_10680,N_14002);
nor U17215 (N_17215,N_13643,N_10868);
or U17216 (N_17216,N_10354,N_13359);
nor U17217 (N_17217,N_11400,N_10790);
and U17218 (N_17218,N_14611,N_11820);
and U17219 (N_17219,N_13142,N_14714);
nand U17220 (N_17220,N_10774,N_12816);
xor U17221 (N_17221,N_11686,N_11457);
nand U17222 (N_17222,N_14740,N_10243);
nor U17223 (N_17223,N_12351,N_12615);
and U17224 (N_17224,N_10214,N_11719);
or U17225 (N_17225,N_12132,N_14270);
and U17226 (N_17226,N_14901,N_13029);
nor U17227 (N_17227,N_14713,N_12224);
and U17228 (N_17228,N_11690,N_11632);
or U17229 (N_17229,N_13257,N_11020);
nor U17230 (N_17230,N_10344,N_14718);
nor U17231 (N_17231,N_14876,N_12378);
and U17232 (N_17232,N_12450,N_11732);
and U17233 (N_17233,N_10286,N_12974);
nor U17234 (N_17234,N_14298,N_10210);
nor U17235 (N_17235,N_12191,N_12756);
nand U17236 (N_17236,N_11576,N_10852);
or U17237 (N_17237,N_12854,N_13006);
nand U17238 (N_17238,N_13468,N_11445);
or U17239 (N_17239,N_11097,N_10129);
nand U17240 (N_17240,N_10740,N_14600);
nand U17241 (N_17241,N_11003,N_11489);
or U17242 (N_17242,N_14673,N_13672);
nor U17243 (N_17243,N_14996,N_11889);
xor U17244 (N_17244,N_14883,N_11084);
or U17245 (N_17245,N_14389,N_11853);
nand U17246 (N_17246,N_13908,N_14423);
or U17247 (N_17247,N_12494,N_12075);
or U17248 (N_17248,N_14863,N_13185);
xnor U17249 (N_17249,N_11439,N_13987);
nor U17250 (N_17250,N_10415,N_12295);
and U17251 (N_17251,N_10004,N_14864);
or U17252 (N_17252,N_12466,N_10562);
nand U17253 (N_17253,N_11371,N_14159);
and U17254 (N_17254,N_10856,N_10891);
nand U17255 (N_17255,N_12072,N_11870);
or U17256 (N_17256,N_13905,N_14107);
and U17257 (N_17257,N_13436,N_14231);
and U17258 (N_17258,N_14661,N_10398);
and U17259 (N_17259,N_14707,N_11925);
nor U17260 (N_17260,N_12546,N_11629);
or U17261 (N_17261,N_12060,N_12880);
nor U17262 (N_17262,N_13462,N_11823);
nor U17263 (N_17263,N_13771,N_13415);
or U17264 (N_17264,N_10938,N_11017);
nand U17265 (N_17265,N_13950,N_14179);
or U17266 (N_17266,N_11410,N_14557);
and U17267 (N_17267,N_14531,N_11420);
and U17268 (N_17268,N_12505,N_14040);
and U17269 (N_17269,N_13387,N_14957);
nor U17270 (N_17270,N_12383,N_13471);
nand U17271 (N_17271,N_12584,N_12310);
or U17272 (N_17272,N_13337,N_13542);
nand U17273 (N_17273,N_12367,N_13066);
xnor U17274 (N_17274,N_11013,N_13310);
xnor U17275 (N_17275,N_14791,N_11543);
nor U17276 (N_17276,N_13074,N_13192);
or U17277 (N_17277,N_11349,N_12426);
nor U17278 (N_17278,N_14089,N_14497);
or U17279 (N_17279,N_10164,N_13306);
or U17280 (N_17280,N_14544,N_14721);
or U17281 (N_17281,N_14738,N_11131);
nand U17282 (N_17282,N_13927,N_10877);
and U17283 (N_17283,N_13829,N_12622);
nand U17284 (N_17284,N_14535,N_13532);
nor U17285 (N_17285,N_12707,N_14449);
nand U17286 (N_17286,N_11709,N_12631);
xor U17287 (N_17287,N_11161,N_13371);
xor U17288 (N_17288,N_14822,N_14553);
xor U17289 (N_17289,N_13992,N_10058);
xor U17290 (N_17290,N_12626,N_11687);
or U17291 (N_17291,N_13845,N_13041);
and U17292 (N_17292,N_10585,N_10514);
nor U17293 (N_17293,N_11291,N_11092);
and U17294 (N_17294,N_13996,N_12441);
or U17295 (N_17295,N_14006,N_10999);
or U17296 (N_17296,N_12780,N_10859);
nor U17297 (N_17297,N_12188,N_13936);
xor U17298 (N_17298,N_14200,N_13381);
nor U17299 (N_17299,N_12210,N_13457);
or U17300 (N_17300,N_11058,N_14123);
xor U17301 (N_17301,N_13308,N_13407);
or U17302 (N_17302,N_11921,N_12718);
nand U17303 (N_17303,N_14773,N_13422);
nand U17304 (N_17304,N_13740,N_11289);
or U17305 (N_17305,N_13104,N_12429);
or U17306 (N_17306,N_10341,N_14669);
nand U17307 (N_17307,N_10090,N_10738);
and U17308 (N_17308,N_11292,N_11105);
or U17309 (N_17309,N_12923,N_14655);
and U17310 (N_17310,N_13214,N_11694);
or U17311 (N_17311,N_14153,N_11916);
nand U17312 (N_17312,N_10821,N_12892);
or U17313 (N_17313,N_11304,N_11368);
xor U17314 (N_17314,N_12076,N_10025);
nand U17315 (N_17315,N_11974,N_10498);
or U17316 (N_17316,N_13186,N_12525);
and U17317 (N_17317,N_11944,N_10571);
or U17318 (N_17318,N_14746,N_10380);
and U17319 (N_17319,N_13425,N_14490);
nor U17320 (N_17320,N_12355,N_10577);
nor U17321 (N_17321,N_11184,N_11636);
or U17322 (N_17322,N_13677,N_13281);
nand U17323 (N_17323,N_13998,N_14217);
nor U17324 (N_17324,N_14862,N_14227);
nor U17325 (N_17325,N_11485,N_14464);
or U17326 (N_17326,N_13200,N_12227);
and U17327 (N_17327,N_14110,N_10158);
and U17328 (N_17328,N_11370,N_10565);
nor U17329 (N_17329,N_10200,N_10265);
nand U17330 (N_17330,N_14459,N_11208);
nor U17331 (N_17331,N_10545,N_14870);
nor U17332 (N_17332,N_13527,N_13806);
or U17333 (N_17333,N_13531,N_10291);
or U17334 (N_17334,N_14810,N_13141);
nor U17335 (N_17335,N_10349,N_11901);
nand U17336 (N_17336,N_12409,N_11321);
and U17337 (N_17337,N_11770,N_13731);
or U17338 (N_17338,N_10374,N_13666);
and U17339 (N_17339,N_14142,N_12909);
nand U17340 (N_17340,N_12662,N_10757);
nor U17341 (N_17341,N_13225,N_11638);
and U17342 (N_17342,N_11545,N_14973);
or U17343 (N_17343,N_14964,N_12431);
or U17344 (N_17344,N_14458,N_14666);
and U17345 (N_17345,N_12118,N_14265);
nand U17346 (N_17346,N_11005,N_13697);
nor U17347 (N_17347,N_14454,N_10704);
nor U17348 (N_17348,N_11597,N_10568);
and U17349 (N_17349,N_11169,N_12266);
nor U17350 (N_17350,N_10445,N_10510);
nand U17351 (N_17351,N_10269,N_11274);
nand U17352 (N_17352,N_12789,N_14871);
nand U17353 (N_17353,N_11665,N_10556);
nor U17354 (N_17354,N_10787,N_11346);
nand U17355 (N_17355,N_12184,N_14546);
or U17356 (N_17356,N_11347,N_11170);
and U17357 (N_17357,N_12568,N_14832);
or U17358 (N_17358,N_11389,N_11164);
or U17359 (N_17359,N_12934,N_13086);
and U17360 (N_17360,N_10366,N_10530);
nand U17361 (N_17361,N_11692,N_12044);
or U17362 (N_17362,N_13182,N_13264);
nor U17363 (N_17363,N_13492,N_12254);
and U17364 (N_17364,N_12276,N_10523);
nor U17365 (N_17365,N_11642,N_11163);
xnor U17366 (N_17366,N_13456,N_13761);
nor U17367 (N_17367,N_14125,N_14951);
nand U17368 (N_17368,N_10943,N_13084);
and U17369 (N_17369,N_11735,N_11740);
xnor U17370 (N_17370,N_11189,N_11310);
and U17371 (N_17371,N_13680,N_11040);
nor U17372 (N_17372,N_11305,N_10963);
nor U17373 (N_17373,N_14805,N_11701);
and U17374 (N_17374,N_12032,N_10809);
nand U17375 (N_17375,N_14606,N_10417);
or U17376 (N_17376,N_14052,N_13684);
nand U17377 (N_17377,N_10412,N_13197);
or U17378 (N_17378,N_11399,N_14049);
nand U17379 (N_17379,N_14416,N_14597);
nand U17380 (N_17380,N_13449,N_10487);
nand U17381 (N_17381,N_13172,N_11240);
nor U17382 (N_17382,N_13910,N_14624);
and U17383 (N_17383,N_14770,N_13143);
xnor U17384 (N_17384,N_11253,N_11899);
nand U17385 (N_17385,N_14382,N_12997);
nand U17386 (N_17386,N_14554,N_12689);
nor U17387 (N_17387,N_11675,N_12666);
and U17388 (N_17388,N_14198,N_10896);
nor U17389 (N_17389,N_13912,N_13375);
nand U17390 (N_17390,N_12318,N_11246);
or U17391 (N_17391,N_12272,N_13463);
and U17392 (N_17392,N_14121,N_12785);
nor U17393 (N_17393,N_14031,N_12225);
xor U17394 (N_17394,N_14457,N_11238);
or U17395 (N_17395,N_13211,N_13515);
or U17396 (N_17396,N_13514,N_10384);
xnor U17397 (N_17397,N_13088,N_11137);
nand U17398 (N_17398,N_12193,N_11805);
and U17399 (N_17399,N_14057,N_13093);
nand U17400 (N_17400,N_11653,N_14181);
and U17401 (N_17401,N_12168,N_10500);
nand U17402 (N_17402,N_12552,N_13116);
nor U17403 (N_17403,N_11898,N_13983);
and U17404 (N_17404,N_10619,N_11727);
and U17405 (N_17405,N_12878,N_12080);
or U17406 (N_17406,N_14093,N_12447);
nand U17407 (N_17407,N_11290,N_13760);
nor U17408 (N_17408,N_12302,N_11193);
nand U17409 (N_17409,N_14730,N_14843);
xnor U17410 (N_17410,N_10867,N_10315);
nand U17411 (N_17411,N_14167,N_12398);
and U17412 (N_17412,N_13423,N_10367);
nand U17413 (N_17413,N_10165,N_13698);
and U17414 (N_17414,N_12105,N_10802);
nand U17415 (N_17415,N_10779,N_14162);
and U17416 (N_17416,N_11360,N_13323);
nand U17417 (N_17417,N_12969,N_13475);
nand U17418 (N_17418,N_10285,N_10073);
or U17419 (N_17419,N_14889,N_13516);
nand U17420 (N_17420,N_11760,N_11139);
and U17421 (N_17421,N_13263,N_14417);
nor U17422 (N_17422,N_11356,N_13727);
or U17423 (N_17423,N_12895,N_13863);
xnor U17424 (N_17424,N_14551,N_12799);
or U17425 (N_17425,N_12824,N_13632);
nand U17426 (N_17426,N_11096,N_13237);
nand U17427 (N_17427,N_11971,N_14193);
nor U17428 (N_17428,N_12199,N_10968);
nor U17429 (N_17429,N_14228,N_14841);
nand U17430 (N_17430,N_11566,N_11252);
nor U17431 (N_17431,N_14869,N_12198);
xor U17432 (N_17432,N_12419,N_10017);
or U17433 (N_17433,N_10502,N_12762);
nand U17434 (N_17434,N_12988,N_10990);
or U17435 (N_17435,N_13639,N_10020);
and U17436 (N_17436,N_14238,N_14944);
or U17437 (N_17437,N_13969,N_10641);
and U17438 (N_17438,N_13962,N_12543);
nand U17439 (N_17439,N_13937,N_14453);
or U17440 (N_17440,N_10318,N_10352);
nand U17441 (N_17441,N_12576,N_11023);
or U17442 (N_17442,N_10101,N_11118);
nor U17443 (N_17443,N_12698,N_11519);
and U17444 (N_17444,N_14264,N_12982);
nor U17445 (N_17445,N_12765,N_14793);
and U17446 (N_17446,N_13011,N_10776);
xor U17447 (N_17447,N_10038,N_12629);
or U17448 (N_17448,N_12990,N_13372);
and U17449 (N_17449,N_14905,N_14379);
or U17450 (N_17450,N_13534,N_10080);
and U17451 (N_17451,N_14034,N_11409);
or U17452 (N_17452,N_11098,N_11250);
nand U17453 (N_17453,N_10242,N_10674);
nand U17454 (N_17454,N_10600,N_13134);
nor U17455 (N_17455,N_11209,N_10573);
or U17456 (N_17456,N_11213,N_13686);
nor U17457 (N_17457,N_11244,N_13329);
nand U17458 (N_17458,N_11027,N_12491);
nand U17459 (N_17459,N_10015,N_13277);
nor U17460 (N_17460,N_10717,N_14104);
nand U17461 (N_17461,N_14595,N_14890);
or U17462 (N_17462,N_12912,N_11422);
nor U17463 (N_17463,N_11001,N_12618);
xor U17464 (N_17464,N_14476,N_10112);
nand U17465 (N_17465,N_12092,N_13574);
nor U17466 (N_17466,N_12606,N_10283);
nand U17467 (N_17467,N_10368,N_12400);
or U17468 (N_17468,N_11041,N_13894);
and U17469 (N_17469,N_11817,N_12861);
nor U17470 (N_17470,N_14671,N_12112);
and U17471 (N_17471,N_13943,N_12736);
and U17472 (N_17472,N_13676,N_13026);
nand U17473 (N_17473,N_13452,N_10529);
nor U17474 (N_17474,N_14897,N_12133);
nor U17475 (N_17475,N_14971,N_12476);
and U17476 (N_17476,N_11622,N_11871);
nor U17477 (N_17477,N_11154,N_13823);
or U17478 (N_17478,N_10603,N_10639);
or U17479 (N_17479,N_12068,N_13785);
nand U17480 (N_17480,N_10893,N_13512);
xnor U17481 (N_17481,N_10720,N_11954);
nand U17482 (N_17482,N_10645,N_11381);
nand U17483 (N_17483,N_11119,N_11302);
and U17484 (N_17484,N_13710,N_14456);
nor U17485 (N_17485,N_11078,N_11212);
or U17486 (N_17486,N_12109,N_10123);
or U17487 (N_17487,N_14044,N_13059);
nand U17488 (N_17488,N_13042,N_13868);
nand U17489 (N_17489,N_11196,N_10841);
nand U17490 (N_17490,N_12879,N_11678);
or U17491 (N_17491,N_13139,N_13661);
nor U17492 (N_17492,N_13251,N_11424);
nor U17493 (N_17493,N_10126,N_13700);
and U17494 (N_17494,N_11560,N_12600);
xnor U17495 (N_17495,N_10399,N_14078);
or U17496 (N_17496,N_12983,N_10965);
nor U17497 (N_17497,N_12238,N_14946);
and U17498 (N_17498,N_10097,N_10462);
nand U17499 (N_17499,N_12062,N_14877);
and U17500 (N_17500,N_12051,N_13098);
or U17501 (N_17501,N_11119,N_13408);
and U17502 (N_17502,N_12105,N_14506);
xnor U17503 (N_17503,N_10228,N_12422);
nor U17504 (N_17504,N_13293,N_12213);
nor U17505 (N_17505,N_10015,N_13938);
xnor U17506 (N_17506,N_12586,N_12561);
nor U17507 (N_17507,N_14043,N_11952);
and U17508 (N_17508,N_13052,N_13520);
nor U17509 (N_17509,N_13709,N_12242);
and U17510 (N_17510,N_13940,N_10581);
nand U17511 (N_17511,N_11097,N_10044);
xor U17512 (N_17512,N_12814,N_10173);
or U17513 (N_17513,N_13226,N_14710);
nor U17514 (N_17514,N_11644,N_12226);
xnor U17515 (N_17515,N_11598,N_11875);
nand U17516 (N_17516,N_10528,N_13856);
or U17517 (N_17517,N_13152,N_12043);
xnor U17518 (N_17518,N_10835,N_14106);
and U17519 (N_17519,N_13431,N_11656);
nand U17520 (N_17520,N_11157,N_10975);
nand U17521 (N_17521,N_11696,N_12458);
and U17522 (N_17522,N_13437,N_14889);
or U17523 (N_17523,N_10246,N_11094);
or U17524 (N_17524,N_12580,N_11824);
nor U17525 (N_17525,N_14850,N_11622);
nor U17526 (N_17526,N_11445,N_11686);
nand U17527 (N_17527,N_10075,N_12010);
nand U17528 (N_17528,N_11790,N_11358);
and U17529 (N_17529,N_11223,N_11252);
and U17530 (N_17530,N_13650,N_11430);
or U17531 (N_17531,N_13153,N_13991);
and U17532 (N_17532,N_11000,N_12812);
and U17533 (N_17533,N_12213,N_13230);
nor U17534 (N_17534,N_13467,N_13959);
nor U17535 (N_17535,N_10163,N_11703);
or U17536 (N_17536,N_11595,N_11082);
nand U17537 (N_17537,N_14804,N_13706);
nand U17538 (N_17538,N_13235,N_13327);
nor U17539 (N_17539,N_11613,N_13395);
or U17540 (N_17540,N_14995,N_11260);
or U17541 (N_17541,N_14284,N_14844);
nand U17542 (N_17542,N_11605,N_14031);
nor U17543 (N_17543,N_11370,N_11646);
or U17544 (N_17544,N_11274,N_10915);
nand U17545 (N_17545,N_12812,N_10828);
nor U17546 (N_17546,N_10379,N_12389);
or U17547 (N_17547,N_10488,N_13899);
xor U17548 (N_17548,N_14015,N_14683);
and U17549 (N_17549,N_11698,N_13487);
and U17550 (N_17550,N_10561,N_12097);
or U17551 (N_17551,N_14108,N_14502);
or U17552 (N_17552,N_14864,N_12293);
nand U17553 (N_17553,N_12361,N_11615);
nor U17554 (N_17554,N_14473,N_14797);
or U17555 (N_17555,N_14916,N_11204);
or U17556 (N_17556,N_10522,N_11071);
and U17557 (N_17557,N_10902,N_11115);
nor U17558 (N_17558,N_14878,N_12346);
nor U17559 (N_17559,N_13461,N_14915);
or U17560 (N_17560,N_14455,N_12375);
and U17561 (N_17561,N_14555,N_10494);
nand U17562 (N_17562,N_10795,N_13681);
nand U17563 (N_17563,N_10659,N_12957);
nor U17564 (N_17564,N_14321,N_13015);
xnor U17565 (N_17565,N_11709,N_12265);
or U17566 (N_17566,N_11320,N_13155);
nor U17567 (N_17567,N_13138,N_12510);
nand U17568 (N_17568,N_10246,N_11701);
or U17569 (N_17569,N_10960,N_12386);
nand U17570 (N_17570,N_11774,N_10035);
nor U17571 (N_17571,N_11963,N_14929);
nand U17572 (N_17572,N_14514,N_10439);
or U17573 (N_17573,N_12647,N_11131);
nor U17574 (N_17574,N_14149,N_12165);
or U17575 (N_17575,N_13175,N_14501);
or U17576 (N_17576,N_12774,N_12149);
nand U17577 (N_17577,N_11061,N_12278);
xnor U17578 (N_17578,N_11207,N_11025);
nor U17579 (N_17579,N_14858,N_14412);
or U17580 (N_17580,N_12643,N_11388);
and U17581 (N_17581,N_10504,N_11687);
or U17582 (N_17582,N_14623,N_11650);
or U17583 (N_17583,N_11424,N_14129);
nand U17584 (N_17584,N_11642,N_12861);
xor U17585 (N_17585,N_10330,N_12208);
nand U17586 (N_17586,N_14907,N_11848);
nand U17587 (N_17587,N_10051,N_13912);
nand U17588 (N_17588,N_14175,N_14647);
nor U17589 (N_17589,N_12146,N_14769);
nand U17590 (N_17590,N_10661,N_14519);
xnor U17591 (N_17591,N_10366,N_14010);
nand U17592 (N_17592,N_14882,N_13342);
and U17593 (N_17593,N_12348,N_14771);
nor U17594 (N_17594,N_13303,N_12905);
nor U17595 (N_17595,N_13828,N_11801);
nor U17596 (N_17596,N_14905,N_12115);
nor U17597 (N_17597,N_14254,N_10929);
nor U17598 (N_17598,N_10332,N_13296);
and U17599 (N_17599,N_13894,N_14100);
nor U17600 (N_17600,N_10733,N_10249);
nor U17601 (N_17601,N_13505,N_14527);
or U17602 (N_17602,N_10205,N_10202);
nand U17603 (N_17603,N_13186,N_11008);
nor U17604 (N_17604,N_12691,N_13436);
or U17605 (N_17605,N_13381,N_12559);
and U17606 (N_17606,N_12782,N_12302);
nand U17607 (N_17607,N_13367,N_12009);
nor U17608 (N_17608,N_13168,N_14333);
nor U17609 (N_17609,N_14769,N_10079);
or U17610 (N_17610,N_10294,N_14912);
and U17611 (N_17611,N_11892,N_11742);
or U17612 (N_17612,N_10944,N_11633);
xor U17613 (N_17613,N_11829,N_14299);
and U17614 (N_17614,N_13246,N_14274);
and U17615 (N_17615,N_10105,N_12860);
nand U17616 (N_17616,N_11219,N_14166);
nor U17617 (N_17617,N_14662,N_14894);
nand U17618 (N_17618,N_14376,N_12568);
or U17619 (N_17619,N_10689,N_14670);
and U17620 (N_17620,N_14531,N_14052);
and U17621 (N_17621,N_12788,N_11559);
nor U17622 (N_17622,N_14265,N_11800);
and U17623 (N_17623,N_12382,N_11162);
xnor U17624 (N_17624,N_10309,N_11863);
nor U17625 (N_17625,N_14397,N_14975);
xnor U17626 (N_17626,N_13779,N_14423);
and U17627 (N_17627,N_13556,N_14875);
nand U17628 (N_17628,N_13415,N_14930);
nand U17629 (N_17629,N_12275,N_10280);
nand U17630 (N_17630,N_13584,N_14042);
and U17631 (N_17631,N_10862,N_14592);
nor U17632 (N_17632,N_10840,N_14215);
xnor U17633 (N_17633,N_13028,N_14978);
and U17634 (N_17634,N_10201,N_11864);
nor U17635 (N_17635,N_12906,N_10810);
or U17636 (N_17636,N_13024,N_13695);
or U17637 (N_17637,N_13427,N_12466);
xnor U17638 (N_17638,N_11204,N_11223);
or U17639 (N_17639,N_13052,N_13321);
and U17640 (N_17640,N_13189,N_11384);
nand U17641 (N_17641,N_11928,N_13587);
nor U17642 (N_17642,N_14686,N_14182);
nor U17643 (N_17643,N_12846,N_13810);
nand U17644 (N_17644,N_13679,N_11830);
nand U17645 (N_17645,N_10394,N_12899);
or U17646 (N_17646,N_12239,N_12162);
or U17647 (N_17647,N_14481,N_11508);
or U17648 (N_17648,N_12175,N_10367);
and U17649 (N_17649,N_14701,N_12020);
nor U17650 (N_17650,N_14695,N_14987);
nand U17651 (N_17651,N_13546,N_11638);
xor U17652 (N_17652,N_10074,N_11609);
nor U17653 (N_17653,N_13421,N_12410);
nor U17654 (N_17654,N_12747,N_12710);
or U17655 (N_17655,N_14494,N_10605);
or U17656 (N_17656,N_14174,N_11708);
nor U17657 (N_17657,N_14628,N_10742);
nor U17658 (N_17658,N_10889,N_11728);
or U17659 (N_17659,N_11124,N_11919);
xnor U17660 (N_17660,N_13519,N_12758);
or U17661 (N_17661,N_11447,N_12656);
nand U17662 (N_17662,N_13049,N_11152);
xor U17663 (N_17663,N_14875,N_10603);
nand U17664 (N_17664,N_13320,N_14726);
nand U17665 (N_17665,N_10622,N_12039);
nand U17666 (N_17666,N_12740,N_12949);
and U17667 (N_17667,N_12176,N_13958);
and U17668 (N_17668,N_14249,N_14656);
and U17669 (N_17669,N_11966,N_13007);
nand U17670 (N_17670,N_11296,N_11452);
and U17671 (N_17671,N_12378,N_11820);
xnor U17672 (N_17672,N_12072,N_14541);
xnor U17673 (N_17673,N_13093,N_10333);
and U17674 (N_17674,N_14851,N_10299);
and U17675 (N_17675,N_10783,N_14805);
and U17676 (N_17676,N_11245,N_12576);
or U17677 (N_17677,N_11308,N_13448);
xor U17678 (N_17678,N_10802,N_12655);
xnor U17679 (N_17679,N_10910,N_14323);
or U17680 (N_17680,N_13825,N_11594);
or U17681 (N_17681,N_10568,N_10027);
nand U17682 (N_17682,N_10197,N_10467);
nor U17683 (N_17683,N_12778,N_14430);
nor U17684 (N_17684,N_12926,N_12650);
nor U17685 (N_17685,N_13492,N_12137);
or U17686 (N_17686,N_13321,N_11042);
nor U17687 (N_17687,N_12399,N_13779);
nor U17688 (N_17688,N_10288,N_13845);
or U17689 (N_17689,N_11111,N_12119);
nand U17690 (N_17690,N_11376,N_11169);
or U17691 (N_17691,N_12532,N_10510);
xnor U17692 (N_17692,N_12033,N_12818);
and U17693 (N_17693,N_14612,N_14176);
nor U17694 (N_17694,N_14190,N_11163);
or U17695 (N_17695,N_12746,N_13809);
nor U17696 (N_17696,N_10579,N_14744);
nand U17697 (N_17697,N_11989,N_14878);
or U17698 (N_17698,N_11755,N_11899);
or U17699 (N_17699,N_11509,N_14109);
or U17700 (N_17700,N_13117,N_14106);
xor U17701 (N_17701,N_12035,N_11762);
and U17702 (N_17702,N_14322,N_13283);
nor U17703 (N_17703,N_14447,N_12636);
nand U17704 (N_17704,N_11194,N_13052);
or U17705 (N_17705,N_11814,N_10461);
nand U17706 (N_17706,N_12817,N_13249);
nor U17707 (N_17707,N_12737,N_13786);
and U17708 (N_17708,N_13025,N_13586);
xnor U17709 (N_17709,N_10360,N_13516);
nor U17710 (N_17710,N_10976,N_10015);
nand U17711 (N_17711,N_11269,N_11669);
nand U17712 (N_17712,N_12060,N_10541);
and U17713 (N_17713,N_11469,N_11588);
and U17714 (N_17714,N_12127,N_13185);
or U17715 (N_17715,N_12611,N_10527);
nor U17716 (N_17716,N_12318,N_11087);
or U17717 (N_17717,N_11004,N_10747);
or U17718 (N_17718,N_13204,N_13344);
and U17719 (N_17719,N_12824,N_13233);
or U17720 (N_17720,N_12460,N_12703);
xor U17721 (N_17721,N_10556,N_11087);
or U17722 (N_17722,N_13418,N_12385);
nand U17723 (N_17723,N_14131,N_12359);
or U17724 (N_17724,N_10446,N_14992);
and U17725 (N_17725,N_11787,N_12431);
or U17726 (N_17726,N_13368,N_14576);
or U17727 (N_17727,N_12558,N_10013);
nand U17728 (N_17728,N_14707,N_14784);
xnor U17729 (N_17729,N_12620,N_14562);
xor U17730 (N_17730,N_13343,N_11040);
or U17731 (N_17731,N_11176,N_11354);
and U17732 (N_17732,N_12035,N_13720);
and U17733 (N_17733,N_10964,N_14754);
nand U17734 (N_17734,N_14957,N_14396);
nor U17735 (N_17735,N_10211,N_11357);
nor U17736 (N_17736,N_11448,N_11832);
and U17737 (N_17737,N_12855,N_12636);
nand U17738 (N_17738,N_14564,N_11705);
xor U17739 (N_17739,N_10626,N_12329);
nand U17740 (N_17740,N_10905,N_14476);
nand U17741 (N_17741,N_11332,N_14592);
nor U17742 (N_17742,N_11598,N_13002);
nor U17743 (N_17743,N_13241,N_14654);
nand U17744 (N_17744,N_10325,N_11563);
nor U17745 (N_17745,N_13827,N_13318);
nor U17746 (N_17746,N_10556,N_11053);
or U17747 (N_17747,N_11758,N_13051);
or U17748 (N_17748,N_14381,N_12955);
nor U17749 (N_17749,N_12796,N_11403);
nand U17750 (N_17750,N_12234,N_14818);
and U17751 (N_17751,N_10497,N_13773);
xor U17752 (N_17752,N_12864,N_12866);
nor U17753 (N_17753,N_10559,N_12021);
or U17754 (N_17754,N_11745,N_14824);
and U17755 (N_17755,N_12369,N_13884);
or U17756 (N_17756,N_11976,N_13879);
xor U17757 (N_17757,N_13667,N_11708);
or U17758 (N_17758,N_14412,N_12296);
or U17759 (N_17759,N_12893,N_14337);
nor U17760 (N_17760,N_10519,N_12790);
xnor U17761 (N_17761,N_10183,N_10555);
xnor U17762 (N_17762,N_12679,N_11734);
and U17763 (N_17763,N_11676,N_10977);
and U17764 (N_17764,N_10037,N_14784);
or U17765 (N_17765,N_11115,N_13422);
and U17766 (N_17766,N_12127,N_12733);
or U17767 (N_17767,N_11281,N_10987);
or U17768 (N_17768,N_12698,N_13669);
nand U17769 (N_17769,N_14880,N_12363);
xnor U17770 (N_17770,N_14130,N_13275);
or U17771 (N_17771,N_10804,N_14905);
nand U17772 (N_17772,N_10497,N_14266);
nand U17773 (N_17773,N_14831,N_13876);
nand U17774 (N_17774,N_10738,N_13727);
nor U17775 (N_17775,N_10879,N_11958);
nor U17776 (N_17776,N_14224,N_12790);
nor U17777 (N_17777,N_11175,N_11254);
xor U17778 (N_17778,N_10243,N_11664);
nand U17779 (N_17779,N_10464,N_12108);
nand U17780 (N_17780,N_12320,N_11899);
nand U17781 (N_17781,N_13358,N_14479);
nand U17782 (N_17782,N_13937,N_13209);
or U17783 (N_17783,N_12207,N_12657);
xnor U17784 (N_17784,N_13386,N_14156);
nor U17785 (N_17785,N_11206,N_14309);
xor U17786 (N_17786,N_12168,N_14067);
and U17787 (N_17787,N_12304,N_12880);
nand U17788 (N_17788,N_12966,N_11190);
or U17789 (N_17789,N_11829,N_12983);
nand U17790 (N_17790,N_13493,N_11555);
and U17791 (N_17791,N_14051,N_11218);
and U17792 (N_17792,N_14214,N_10145);
or U17793 (N_17793,N_13013,N_11287);
or U17794 (N_17794,N_11422,N_11478);
nor U17795 (N_17795,N_10405,N_10565);
nand U17796 (N_17796,N_12054,N_13122);
nand U17797 (N_17797,N_10935,N_14704);
and U17798 (N_17798,N_10762,N_13099);
and U17799 (N_17799,N_13985,N_14061);
nand U17800 (N_17800,N_11395,N_11741);
nand U17801 (N_17801,N_10786,N_12679);
and U17802 (N_17802,N_14038,N_14669);
nor U17803 (N_17803,N_12673,N_10852);
nand U17804 (N_17804,N_11512,N_10055);
or U17805 (N_17805,N_14897,N_12211);
nor U17806 (N_17806,N_11991,N_12301);
xor U17807 (N_17807,N_10722,N_13661);
and U17808 (N_17808,N_12865,N_13672);
and U17809 (N_17809,N_11033,N_12994);
or U17810 (N_17810,N_10398,N_12994);
or U17811 (N_17811,N_12467,N_14583);
nand U17812 (N_17812,N_12697,N_13032);
nor U17813 (N_17813,N_14782,N_13510);
and U17814 (N_17814,N_14203,N_12057);
nand U17815 (N_17815,N_11818,N_10033);
and U17816 (N_17816,N_14299,N_13231);
nand U17817 (N_17817,N_14379,N_12769);
and U17818 (N_17818,N_13384,N_14455);
or U17819 (N_17819,N_10992,N_12988);
xor U17820 (N_17820,N_13116,N_10168);
or U17821 (N_17821,N_13668,N_12447);
and U17822 (N_17822,N_11249,N_11096);
or U17823 (N_17823,N_12845,N_14679);
xnor U17824 (N_17824,N_10219,N_14777);
or U17825 (N_17825,N_12348,N_13173);
nor U17826 (N_17826,N_11950,N_11923);
nand U17827 (N_17827,N_11878,N_14932);
or U17828 (N_17828,N_13458,N_13257);
nor U17829 (N_17829,N_12842,N_14373);
nor U17830 (N_17830,N_14589,N_13847);
nor U17831 (N_17831,N_14769,N_12502);
nand U17832 (N_17832,N_13950,N_10310);
nand U17833 (N_17833,N_13836,N_12696);
and U17834 (N_17834,N_13989,N_12382);
or U17835 (N_17835,N_13067,N_10402);
xnor U17836 (N_17836,N_11164,N_14299);
or U17837 (N_17837,N_12852,N_13056);
nor U17838 (N_17838,N_11082,N_12851);
xor U17839 (N_17839,N_12972,N_10769);
and U17840 (N_17840,N_11351,N_14807);
or U17841 (N_17841,N_13497,N_12562);
nor U17842 (N_17842,N_14551,N_13219);
nor U17843 (N_17843,N_13992,N_14851);
or U17844 (N_17844,N_11449,N_11990);
xnor U17845 (N_17845,N_10032,N_10213);
nor U17846 (N_17846,N_14392,N_10030);
or U17847 (N_17847,N_11754,N_13224);
nor U17848 (N_17848,N_10216,N_10365);
and U17849 (N_17849,N_14618,N_13737);
and U17850 (N_17850,N_13796,N_14635);
nor U17851 (N_17851,N_11597,N_13614);
or U17852 (N_17852,N_14056,N_12221);
xor U17853 (N_17853,N_10009,N_14943);
and U17854 (N_17854,N_14322,N_11710);
and U17855 (N_17855,N_14165,N_12690);
or U17856 (N_17856,N_14145,N_12036);
nand U17857 (N_17857,N_14648,N_10002);
or U17858 (N_17858,N_11603,N_13359);
nor U17859 (N_17859,N_13888,N_11408);
nand U17860 (N_17860,N_14643,N_11789);
nor U17861 (N_17861,N_13819,N_14740);
nand U17862 (N_17862,N_11877,N_10217);
xor U17863 (N_17863,N_12034,N_12412);
nor U17864 (N_17864,N_10071,N_14777);
or U17865 (N_17865,N_14525,N_12906);
xor U17866 (N_17866,N_14993,N_13782);
nor U17867 (N_17867,N_13786,N_14008);
nor U17868 (N_17868,N_14095,N_10734);
or U17869 (N_17869,N_13236,N_14963);
or U17870 (N_17870,N_11809,N_12258);
and U17871 (N_17871,N_12650,N_12954);
xor U17872 (N_17872,N_13309,N_10308);
nor U17873 (N_17873,N_13744,N_10860);
and U17874 (N_17874,N_10942,N_13347);
nand U17875 (N_17875,N_11549,N_14615);
nor U17876 (N_17876,N_12313,N_13909);
or U17877 (N_17877,N_10000,N_11158);
xnor U17878 (N_17878,N_14458,N_11471);
nand U17879 (N_17879,N_11576,N_12704);
nor U17880 (N_17880,N_10521,N_13978);
or U17881 (N_17881,N_10796,N_10983);
or U17882 (N_17882,N_11773,N_10629);
nor U17883 (N_17883,N_13905,N_11362);
and U17884 (N_17884,N_14386,N_13525);
and U17885 (N_17885,N_13592,N_12231);
xor U17886 (N_17886,N_14706,N_12082);
and U17887 (N_17887,N_14333,N_13190);
xnor U17888 (N_17888,N_11248,N_14359);
nand U17889 (N_17889,N_12585,N_13676);
nor U17890 (N_17890,N_10741,N_14990);
and U17891 (N_17891,N_12575,N_13002);
nor U17892 (N_17892,N_14173,N_13918);
or U17893 (N_17893,N_13503,N_14244);
xnor U17894 (N_17894,N_14577,N_12100);
or U17895 (N_17895,N_14818,N_10666);
nand U17896 (N_17896,N_12220,N_10820);
and U17897 (N_17897,N_13349,N_14032);
or U17898 (N_17898,N_10735,N_12863);
or U17899 (N_17899,N_14018,N_13436);
and U17900 (N_17900,N_14956,N_12651);
nor U17901 (N_17901,N_12289,N_14755);
or U17902 (N_17902,N_12628,N_11596);
nand U17903 (N_17903,N_13005,N_11082);
and U17904 (N_17904,N_12380,N_12164);
and U17905 (N_17905,N_13673,N_10776);
or U17906 (N_17906,N_13500,N_12340);
nand U17907 (N_17907,N_13612,N_10567);
and U17908 (N_17908,N_12432,N_11416);
nand U17909 (N_17909,N_13810,N_11960);
or U17910 (N_17910,N_13787,N_13123);
and U17911 (N_17911,N_10262,N_13138);
nor U17912 (N_17912,N_12198,N_11383);
nand U17913 (N_17913,N_13214,N_10609);
and U17914 (N_17914,N_11603,N_12455);
nor U17915 (N_17915,N_11917,N_12742);
xnor U17916 (N_17916,N_14069,N_10516);
nand U17917 (N_17917,N_14253,N_13387);
nor U17918 (N_17918,N_11207,N_12671);
and U17919 (N_17919,N_14375,N_12514);
nand U17920 (N_17920,N_14653,N_14285);
and U17921 (N_17921,N_11161,N_11052);
and U17922 (N_17922,N_13513,N_11787);
nand U17923 (N_17923,N_10817,N_13692);
nor U17924 (N_17924,N_13015,N_13986);
nor U17925 (N_17925,N_12944,N_13064);
nand U17926 (N_17926,N_11582,N_11581);
or U17927 (N_17927,N_13987,N_12600);
nand U17928 (N_17928,N_10782,N_14772);
xnor U17929 (N_17929,N_14429,N_11257);
nor U17930 (N_17930,N_10417,N_12806);
xor U17931 (N_17931,N_14140,N_10841);
or U17932 (N_17932,N_11779,N_10620);
or U17933 (N_17933,N_12618,N_12374);
nand U17934 (N_17934,N_10546,N_11319);
nand U17935 (N_17935,N_13058,N_13682);
nand U17936 (N_17936,N_13265,N_12993);
or U17937 (N_17937,N_13473,N_13506);
nor U17938 (N_17938,N_11717,N_13113);
nand U17939 (N_17939,N_12298,N_14909);
nor U17940 (N_17940,N_12500,N_11883);
nand U17941 (N_17941,N_13089,N_12920);
and U17942 (N_17942,N_12265,N_14164);
and U17943 (N_17943,N_12727,N_13168);
and U17944 (N_17944,N_10746,N_12678);
and U17945 (N_17945,N_13458,N_12664);
nand U17946 (N_17946,N_14590,N_11045);
nor U17947 (N_17947,N_13630,N_12430);
or U17948 (N_17948,N_10007,N_13671);
xnor U17949 (N_17949,N_13734,N_12580);
and U17950 (N_17950,N_11234,N_14315);
and U17951 (N_17951,N_10444,N_12291);
and U17952 (N_17952,N_14879,N_11574);
or U17953 (N_17953,N_11753,N_10012);
and U17954 (N_17954,N_12666,N_13065);
and U17955 (N_17955,N_12102,N_12258);
or U17956 (N_17956,N_11952,N_11534);
and U17957 (N_17957,N_13401,N_12316);
nor U17958 (N_17958,N_12446,N_11652);
or U17959 (N_17959,N_12471,N_10203);
and U17960 (N_17960,N_13887,N_10107);
nand U17961 (N_17961,N_11768,N_12422);
nand U17962 (N_17962,N_10828,N_12621);
and U17963 (N_17963,N_12820,N_11229);
and U17964 (N_17964,N_13799,N_13909);
and U17965 (N_17965,N_12072,N_12371);
or U17966 (N_17966,N_12772,N_12140);
xor U17967 (N_17967,N_14621,N_11618);
or U17968 (N_17968,N_14091,N_12581);
nor U17969 (N_17969,N_10560,N_13930);
nand U17970 (N_17970,N_10749,N_12480);
nor U17971 (N_17971,N_14130,N_10236);
and U17972 (N_17972,N_10164,N_12192);
nand U17973 (N_17973,N_12249,N_14029);
nor U17974 (N_17974,N_13550,N_10793);
xnor U17975 (N_17975,N_11553,N_12023);
or U17976 (N_17976,N_11811,N_14321);
nand U17977 (N_17977,N_14796,N_14798);
and U17978 (N_17978,N_13271,N_14180);
nand U17979 (N_17979,N_14211,N_14430);
or U17980 (N_17980,N_10881,N_10562);
and U17981 (N_17981,N_11454,N_13447);
nor U17982 (N_17982,N_10288,N_12462);
xor U17983 (N_17983,N_12893,N_11720);
nor U17984 (N_17984,N_14373,N_13179);
nand U17985 (N_17985,N_11158,N_13670);
and U17986 (N_17986,N_11436,N_12189);
nand U17987 (N_17987,N_10793,N_12286);
or U17988 (N_17988,N_12748,N_11688);
and U17989 (N_17989,N_11206,N_10379);
or U17990 (N_17990,N_12705,N_10954);
nand U17991 (N_17991,N_13500,N_11663);
xor U17992 (N_17992,N_13784,N_12749);
nor U17993 (N_17993,N_12785,N_12061);
nand U17994 (N_17994,N_12723,N_11867);
nor U17995 (N_17995,N_10516,N_14833);
nand U17996 (N_17996,N_11981,N_10274);
xor U17997 (N_17997,N_12361,N_12212);
nor U17998 (N_17998,N_14242,N_12708);
or U17999 (N_17999,N_14810,N_11674);
and U18000 (N_18000,N_10700,N_10653);
nand U18001 (N_18001,N_13998,N_12338);
and U18002 (N_18002,N_13372,N_11371);
or U18003 (N_18003,N_14505,N_12452);
nor U18004 (N_18004,N_14663,N_11600);
xor U18005 (N_18005,N_12851,N_14619);
xor U18006 (N_18006,N_14595,N_11304);
xor U18007 (N_18007,N_10010,N_13055);
nand U18008 (N_18008,N_11164,N_10342);
xnor U18009 (N_18009,N_10121,N_14491);
nor U18010 (N_18010,N_13753,N_14266);
nand U18011 (N_18011,N_12893,N_10334);
xor U18012 (N_18012,N_11245,N_11004);
and U18013 (N_18013,N_14709,N_11268);
nor U18014 (N_18014,N_11245,N_10804);
or U18015 (N_18015,N_11969,N_11611);
nand U18016 (N_18016,N_13349,N_14003);
nand U18017 (N_18017,N_11121,N_12193);
and U18018 (N_18018,N_12401,N_14635);
nand U18019 (N_18019,N_12771,N_14277);
and U18020 (N_18020,N_14242,N_11207);
and U18021 (N_18021,N_12452,N_10691);
or U18022 (N_18022,N_10130,N_12737);
nand U18023 (N_18023,N_14164,N_10554);
and U18024 (N_18024,N_12385,N_11143);
nor U18025 (N_18025,N_11634,N_13982);
and U18026 (N_18026,N_12040,N_14806);
nand U18027 (N_18027,N_14230,N_12903);
nor U18028 (N_18028,N_11039,N_11446);
or U18029 (N_18029,N_10740,N_11142);
nor U18030 (N_18030,N_14365,N_14272);
nand U18031 (N_18031,N_10097,N_10963);
nor U18032 (N_18032,N_13091,N_11341);
nand U18033 (N_18033,N_11310,N_10439);
and U18034 (N_18034,N_10128,N_11750);
xnor U18035 (N_18035,N_10495,N_12895);
nor U18036 (N_18036,N_10578,N_14037);
xor U18037 (N_18037,N_13029,N_10158);
xor U18038 (N_18038,N_10412,N_13327);
nor U18039 (N_18039,N_14071,N_10257);
nand U18040 (N_18040,N_14722,N_10227);
and U18041 (N_18041,N_10247,N_13699);
nor U18042 (N_18042,N_12571,N_14991);
and U18043 (N_18043,N_14195,N_11591);
or U18044 (N_18044,N_12032,N_11431);
nand U18045 (N_18045,N_12919,N_11847);
nor U18046 (N_18046,N_13271,N_11276);
or U18047 (N_18047,N_10048,N_14047);
or U18048 (N_18048,N_13977,N_12261);
nor U18049 (N_18049,N_13806,N_14670);
or U18050 (N_18050,N_11669,N_12113);
or U18051 (N_18051,N_11820,N_13362);
or U18052 (N_18052,N_12762,N_11854);
nor U18053 (N_18053,N_13035,N_12977);
nor U18054 (N_18054,N_14210,N_13703);
xor U18055 (N_18055,N_14661,N_12687);
and U18056 (N_18056,N_10949,N_13733);
nand U18057 (N_18057,N_14156,N_11800);
and U18058 (N_18058,N_12260,N_14123);
xor U18059 (N_18059,N_14666,N_11662);
nor U18060 (N_18060,N_13964,N_10120);
or U18061 (N_18061,N_12500,N_10214);
nand U18062 (N_18062,N_10455,N_11139);
nand U18063 (N_18063,N_12871,N_13774);
or U18064 (N_18064,N_14667,N_14085);
or U18065 (N_18065,N_12585,N_14636);
or U18066 (N_18066,N_13333,N_10285);
nand U18067 (N_18067,N_12542,N_14072);
nor U18068 (N_18068,N_14744,N_12790);
and U18069 (N_18069,N_11973,N_11559);
or U18070 (N_18070,N_11344,N_10456);
and U18071 (N_18071,N_14277,N_13283);
xnor U18072 (N_18072,N_11207,N_11564);
and U18073 (N_18073,N_12070,N_14407);
and U18074 (N_18074,N_13037,N_14719);
nor U18075 (N_18075,N_12309,N_14114);
nand U18076 (N_18076,N_11137,N_11368);
and U18077 (N_18077,N_14876,N_11219);
nand U18078 (N_18078,N_12041,N_12147);
nor U18079 (N_18079,N_14857,N_13061);
and U18080 (N_18080,N_11861,N_14587);
and U18081 (N_18081,N_11632,N_13303);
and U18082 (N_18082,N_12699,N_10477);
nor U18083 (N_18083,N_10426,N_12211);
or U18084 (N_18084,N_10171,N_14790);
nor U18085 (N_18085,N_13492,N_10100);
or U18086 (N_18086,N_12024,N_12615);
nor U18087 (N_18087,N_14974,N_11766);
and U18088 (N_18088,N_12769,N_10378);
xnor U18089 (N_18089,N_12845,N_14366);
and U18090 (N_18090,N_12162,N_10180);
nor U18091 (N_18091,N_11593,N_10020);
xor U18092 (N_18092,N_10222,N_12903);
nand U18093 (N_18093,N_14397,N_14527);
or U18094 (N_18094,N_13977,N_11347);
and U18095 (N_18095,N_13418,N_10291);
or U18096 (N_18096,N_12415,N_12850);
and U18097 (N_18097,N_14957,N_13600);
and U18098 (N_18098,N_11394,N_13738);
xnor U18099 (N_18099,N_11397,N_12631);
and U18100 (N_18100,N_12436,N_10015);
xor U18101 (N_18101,N_10494,N_13136);
nor U18102 (N_18102,N_12728,N_14924);
xnor U18103 (N_18103,N_12650,N_14720);
nand U18104 (N_18104,N_11528,N_11746);
xnor U18105 (N_18105,N_11550,N_12553);
nor U18106 (N_18106,N_14937,N_10261);
nand U18107 (N_18107,N_10630,N_12197);
nand U18108 (N_18108,N_14947,N_13626);
or U18109 (N_18109,N_13772,N_13693);
and U18110 (N_18110,N_14562,N_11894);
or U18111 (N_18111,N_14628,N_14724);
nand U18112 (N_18112,N_12127,N_13994);
and U18113 (N_18113,N_13736,N_12340);
or U18114 (N_18114,N_10052,N_12864);
and U18115 (N_18115,N_10151,N_13795);
and U18116 (N_18116,N_11659,N_11073);
nand U18117 (N_18117,N_12848,N_11927);
and U18118 (N_18118,N_10140,N_14469);
nor U18119 (N_18119,N_13508,N_14836);
and U18120 (N_18120,N_10579,N_14130);
and U18121 (N_18121,N_14020,N_13975);
or U18122 (N_18122,N_12871,N_14471);
and U18123 (N_18123,N_12445,N_13366);
nor U18124 (N_18124,N_12938,N_13173);
nor U18125 (N_18125,N_14835,N_12609);
or U18126 (N_18126,N_12098,N_12868);
nand U18127 (N_18127,N_13798,N_10345);
and U18128 (N_18128,N_13507,N_11892);
and U18129 (N_18129,N_10442,N_13112);
nand U18130 (N_18130,N_13521,N_12299);
nor U18131 (N_18131,N_14013,N_10335);
and U18132 (N_18132,N_14286,N_11525);
nor U18133 (N_18133,N_12131,N_11428);
nand U18134 (N_18134,N_11881,N_14054);
and U18135 (N_18135,N_10593,N_14198);
xor U18136 (N_18136,N_11269,N_14495);
nand U18137 (N_18137,N_14650,N_11550);
and U18138 (N_18138,N_11047,N_13528);
or U18139 (N_18139,N_10454,N_11642);
nand U18140 (N_18140,N_14717,N_11242);
xor U18141 (N_18141,N_13422,N_11016);
or U18142 (N_18142,N_13797,N_12735);
or U18143 (N_18143,N_14886,N_12127);
or U18144 (N_18144,N_13938,N_10696);
or U18145 (N_18145,N_13293,N_11959);
nor U18146 (N_18146,N_10559,N_12497);
and U18147 (N_18147,N_13410,N_11654);
nand U18148 (N_18148,N_14034,N_10669);
nand U18149 (N_18149,N_13841,N_14343);
nor U18150 (N_18150,N_13869,N_14788);
and U18151 (N_18151,N_10719,N_14973);
nor U18152 (N_18152,N_11209,N_11452);
or U18153 (N_18153,N_11017,N_13195);
nand U18154 (N_18154,N_12571,N_14762);
and U18155 (N_18155,N_12033,N_14291);
nor U18156 (N_18156,N_12469,N_12791);
nor U18157 (N_18157,N_13904,N_10342);
and U18158 (N_18158,N_13022,N_12507);
and U18159 (N_18159,N_12148,N_14010);
or U18160 (N_18160,N_12165,N_11692);
and U18161 (N_18161,N_10178,N_13597);
or U18162 (N_18162,N_14004,N_12005);
nand U18163 (N_18163,N_10630,N_10380);
nor U18164 (N_18164,N_11066,N_10474);
nor U18165 (N_18165,N_14212,N_13324);
xnor U18166 (N_18166,N_11041,N_11312);
and U18167 (N_18167,N_13375,N_12604);
and U18168 (N_18168,N_11165,N_13385);
or U18169 (N_18169,N_13514,N_11893);
or U18170 (N_18170,N_14380,N_10484);
nor U18171 (N_18171,N_13485,N_13908);
or U18172 (N_18172,N_10351,N_14590);
nand U18173 (N_18173,N_14634,N_11949);
xor U18174 (N_18174,N_11279,N_11230);
and U18175 (N_18175,N_14772,N_13190);
nand U18176 (N_18176,N_13389,N_10622);
and U18177 (N_18177,N_10112,N_14282);
and U18178 (N_18178,N_14463,N_14827);
and U18179 (N_18179,N_12607,N_14763);
and U18180 (N_18180,N_14334,N_13212);
nor U18181 (N_18181,N_14256,N_12741);
or U18182 (N_18182,N_10537,N_14633);
and U18183 (N_18183,N_11174,N_14764);
and U18184 (N_18184,N_12586,N_10199);
xor U18185 (N_18185,N_13874,N_14225);
and U18186 (N_18186,N_12704,N_11329);
and U18187 (N_18187,N_12727,N_14920);
xnor U18188 (N_18188,N_13317,N_14872);
nand U18189 (N_18189,N_13308,N_14431);
nand U18190 (N_18190,N_14268,N_12560);
nand U18191 (N_18191,N_13832,N_10343);
nand U18192 (N_18192,N_13307,N_14440);
nand U18193 (N_18193,N_10820,N_12323);
nor U18194 (N_18194,N_13452,N_12412);
nor U18195 (N_18195,N_10815,N_11810);
or U18196 (N_18196,N_10819,N_14153);
or U18197 (N_18197,N_12182,N_11084);
nor U18198 (N_18198,N_13185,N_12908);
nand U18199 (N_18199,N_10871,N_13061);
or U18200 (N_18200,N_13886,N_12163);
or U18201 (N_18201,N_10426,N_13805);
and U18202 (N_18202,N_10791,N_14568);
nand U18203 (N_18203,N_11828,N_12296);
xnor U18204 (N_18204,N_12345,N_13472);
nor U18205 (N_18205,N_10228,N_14045);
nand U18206 (N_18206,N_12366,N_11186);
nor U18207 (N_18207,N_11025,N_10777);
nor U18208 (N_18208,N_13206,N_14847);
nor U18209 (N_18209,N_12957,N_13706);
xor U18210 (N_18210,N_10441,N_13739);
and U18211 (N_18211,N_12629,N_10307);
nor U18212 (N_18212,N_12681,N_10737);
xnor U18213 (N_18213,N_12917,N_14112);
nand U18214 (N_18214,N_11513,N_10951);
or U18215 (N_18215,N_13651,N_14716);
nor U18216 (N_18216,N_10507,N_10686);
or U18217 (N_18217,N_10454,N_14197);
xor U18218 (N_18218,N_11580,N_12826);
and U18219 (N_18219,N_14008,N_10876);
nand U18220 (N_18220,N_12184,N_13708);
nand U18221 (N_18221,N_11280,N_14494);
or U18222 (N_18222,N_11199,N_14052);
nand U18223 (N_18223,N_13420,N_12945);
nor U18224 (N_18224,N_10951,N_11947);
nor U18225 (N_18225,N_14613,N_14215);
or U18226 (N_18226,N_11515,N_13668);
nor U18227 (N_18227,N_12941,N_10081);
or U18228 (N_18228,N_13344,N_11699);
xnor U18229 (N_18229,N_10784,N_14700);
nand U18230 (N_18230,N_14893,N_11454);
nand U18231 (N_18231,N_14775,N_11528);
and U18232 (N_18232,N_14930,N_14735);
or U18233 (N_18233,N_13554,N_12699);
or U18234 (N_18234,N_10744,N_12355);
nor U18235 (N_18235,N_14008,N_11296);
nand U18236 (N_18236,N_12089,N_12869);
or U18237 (N_18237,N_10958,N_13798);
and U18238 (N_18238,N_14757,N_13728);
nand U18239 (N_18239,N_12258,N_11444);
or U18240 (N_18240,N_12286,N_11839);
or U18241 (N_18241,N_13763,N_11576);
and U18242 (N_18242,N_12188,N_11158);
nand U18243 (N_18243,N_11950,N_12082);
xnor U18244 (N_18244,N_12698,N_11546);
or U18245 (N_18245,N_14370,N_10567);
and U18246 (N_18246,N_10435,N_13063);
or U18247 (N_18247,N_14999,N_13717);
and U18248 (N_18248,N_14138,N_12947);
nand U18249 (N_18249,N_14485,N_13772);
or U18250 (N_18250,N_13946,N_14789);
nor U18251 (N_18251,N_14517,N_13682);
nand U18252 (N_18252,N_12601,N_10135);
and U18253 (N_18253,N_13463,N_10077);
nor U18254 (N_18254,N_14260,N_14374);
and U18255 (N_18255,N_12161,N_13102);
nand U18256 (N_18256,N_11526,N_13049);
nand U18257 (N_18257,N_14772,N_14946);
nor U18258 (N_18258,N_13035,N_13687);
nor U18259 (N_18259,N_10078,N_12447);
nand U18260 (N_18260,N_13549,N_12798);
and U18261 (N_18261,N_11231,N_12483);
nand U18262 (N_18262,N_12615,N_14684);
and U18263 (N_18263,N_12649,N_10218);
or U18264 (N_18264,N_11530,N_10048);
nand U18265 (N_18265,N_10045,N_14072);
nand U18266 (N_18266,N_12505,N_10484);
and U18267 (N_18267,N_14785,N_13875);
and U18268 (N_18268,N_13172,N_12507);
xor U18269 (N_18269,N_14327,N_13060);
nand U18270 (N_18270,N_14810,N_13635);
nand U18271 (N_18271,N_12610,N_13298);
or U18272 (N_18272,N_10697,N_13556);
and U18273 (N_18273,N_13857,N_10989);
or U18274 (N_18274,N_11055,N_10188);
nor U18275 (N_18275,N_13218,N_14649);
or U18276 (N_18276,N_13274,N_10461);
or U18277 (N_18277,N_14170,N_13842);
xor U18278 (N_18278,N_10546,N_13928);
and U18279 (N_18279,N_14594,N_11561);
nor U18280 (N_18280,N_14383,N_13681);
nor U18281 (N_18281,N_12633,N_12842);
and U18282 (N_18282,N_11637,N_11677);
nand U18283 (N_18283,N_13084,N_10926);
or U18284 (N_18284,N_10247,N_11224);
or U18285 (N_18285,N_10201,N_11102);
and U18286 (N_18286,N_10113,N_13221);
and U18287 (N_18287,N_11187,N_10430);
nor U18288 (N_18288,N_12720,N_11132);
and U18289 (N_18289,N_13036,N_10379);
or U18290 (N_18290,N_13694,N_11401);
nor U18291 (N_18291,N_13978,N_14309);
and U18292 (N_18292,N_10243,N_10711);
or U18293 (N_18293,N_11642,N_14890);
nor U18294 (N_18294,N_11636,N_11628);
nand U18295 (N_18295,N_10541,N_11918);
nor U18296 (N_18296,N_12707,N_13995);
nor U18297 (N_18297,N_10094,N_13515);
nor U18298 (N_18298,N_12976,N_10311);
and U18299 (N_18299,N_12845,N_13525);
nor U18300 (N_18300,N_13689,N_11353);
nand U18301 (N_18301,N_14524,N_14318);
xnor U18302 (N_18302,N_11411,N_10141);
or U18303 (N_18303,N_12225,N_13859);
and U18304 (N_18304,N_11310,N_11477);
nand U18305 (N_18305,N_12492,N_10807);
xor U18306 (N_18306,N_12919,N_11269);
or U18307 (N_18307,N_11188,N_11957);
or U18308 (N_18308,N_11911,N_12598);
nor U18309 (N_18309,N_13470,N_10337);
nand U18310 (N_18310,N_10929,N_10173);
nand U18311 (N_18311,N_11242,N_11898);
nand U18312 (N_18312,N_12661,N_14917);
and U18313 (N_18313,N_11382,N_11558);
and U18314 (N_18314,N_13476,N_12387);
and U18315 (N_18315,N_11984,N_11948);
nor U18316 (N_18316,N_10426,N_14769);
nand U18317 (N_18317,N_12218,N_10746);
and U18318 (N_18318,N_10144,N_10487);
nor U18319 (N_18319,N_14628,N_13283);
and U18320 (N_18320,N_11094,N_13174);
xnor U18321 (N_18321,N_12225,N_14431);
and U18322 (N_18322,N_14301,N_11265);
xnor U18323 (N_18323,N_14455,N_12064);
nand U18324 (N_18324,N_14626,N_11695);
or U18325 (N_18325,N_10104,N_10749);
nand U18326 (N_18326,N_11526,N_10152);
or U18327 (N_18327,N_11850,N_14849);
xnor U18328 (N_18328,N_14490,N_10269);
or U18329 (N_18329,N_14419,N_13721);
or U18330 (N_18330,N_13758,N_10248);
nor U18331 (N_18331,N_11062,N_13147);
xnor U18332 (N_18332,N_11308,N_11490);
nand U18333 (N_18333,N_13359,N_14126);
nor U18334 (N_18334,N_11508,N_12350);
nand U18335 (N_18335,N_11194,N_11372);
and U18336 (N_18336,N_13908,N_13752);
nand U18337 (N_18337,N_11816,N_10032);
nor U18338 (N_18338,N_10827,N_13782);
or U18339 (N_18339,N_12456,N_14757);
nand U18340 (N_18340,N_10034,N_13924);
and U18341 (N_18341,N_14658,N_11425);
nor U18342 (N_18342,N_11461,N_10473);
xnor U18343 (N_18343,N_11766,N_13421);
and U18344 (N_18344,N_11728,N_13484);
xor U18345 (N_18345,N_14186,N_13246);
nor U18346 (N_18346,N_11548,N_14069);
nand U18347 (N_18347,N_13397,N_14991);
nor U18348 (N_18348,N_11863,N_12029);
and U18349 (N_18349,N_14437,N_13737);
or U18350 (N_18350,N_11043,N_11721);
nand U18351 (N_18351,N_12179,N_12212);
nand U18352 (N_18352,N_14586,N_11266);
or U18353 (N_18353,N_10641,N_11946);
or U18354 (N_18354,N_13301,N_10681);
nand U18355 (N_18355,N_14019,N_14368);
nor U18356 (N_18356,N_11665,N_14609);
nand U18357 (N_18357,N_14007,N_10313);
or U18358 (N_18358,N_13437,N_14861);
xor U18359 (N_18359,N_11442,N_11689);
xnor U18360 (N_18360,N_12836,N_11279);
or U18361 (N_18361,N_11686,N_11244);
and U18362 (N_18362,N_14219,N_12499);
xnor U18363 (N_18363,N_12695,N_13808);
or U18364 (N_18364,N_10760,N_14572);
or U18365 (N_18365,N_12469,N_14826);
nor U18366 (N_18366,N_13099,N_12271);
xnor U18367 (N_18367,N_10799,N_10026);
nand U18368 (N_18368,N_13294,N_12783);
nor U18369 (N_18369,N_10345,N_11057);
xor U18370 (N_18370,N_13464,N_14247);
xor U18371 (N_18371,N_12899,N_12960);
nand U18372 (N_18372,N_13026,N_12536);
nor U18373 (N_18373,N_14666,N_11587);
and U18374 (N_18374,N_11137,N_12298);
and U18375 (N_18375,N_13903,N_11930);
or U18376 (N_18376,N_14772,N_12956);
xor U18377 (N_18377,N_13961,N_10805);
or U18378 (N_18378,N_10684,N_11950);
nand U18379 (N_18379,N_14799,N_12262);
xor U18380 (N_18380,N_13584,N_11693);
nor U18381 (N_18381,N_14442,N_10471);
or U18382 (N_18382,N_12281,N_14367);
nand U18383 (N_18383,N_10260,N_11436);
and U18384 (N_18384,N_10571,N_12076);
or U18385 (N_18385,N_10941,N_10874);
nor U18386 (N_18386,N_10510,N_14914);
nor U18387 (N_18387,N_11890,N_13740);
nor U18388 (N_18388,N_12459,N_13635);
xnor U18389 (N_18389,N_13365,N_10871);
nor U18390 (N_18390,N_14407,N_11228);
nand U18391 (N_18391,N_12171,N_11227);
or U18392 (N_18392,N_12193,N_13843);
nor U18393 (N_18393,N_14954,N_14590);
nor U18394 (N_18394,N_10914,N_10057);
nor U18395 (N_18395,N_11957,N_11652);
and U18396 (N_18396,N_10904,N_10425);
xnor U18397 (N_18397,N_14075,N_14216);
nand U18398 (N_18398,N_11545,N_11151);
nand U18399 (N_18399,N_14899,N_11985);
or U18400 (N_18400,N_12968,N_13191);
nor U18401 (N_18401,N_12832,N_11682);
nor U18402 (N_18402,N_14395,N_11570);
and U18403 (N_18403,N_14256,N_10946);
nand U18404 (N_18404,N_12494,N_11851);
and U18405 (N_18405,N_14700,N_10059);
xnor U18406 (N_18406,N_12979,N_13770);
xnor U18407 (N_18407,N_11135,N_10269);
or U18408 (N_18408,N_10166,N_12068);
or U18409 (N_18409,N_10444,N_14012);
and U18410 (N_18410,N_10897,N_14614);
or U18411 (N_18411,N_14246,N_10863);
and U18412 (N_18412,N_14905,N_11483);
and U18413 (N_18413,N_12431,N_14757);
nor U18414 (N_18414,N_11617,N_12109);
nor U18415 (N_18415,N_11128,N_14467);
xor U18416 (N_18416,N_13361,N_10926);
xnor U18417 (N_18417,N_12727,N_11601);
or U18418 (N_18418,N_11829,N_14448);
and U18419 (N_18419,N_10682,N_10061);
and U18420 (N_18420,N_11215,N_11607);
xor U18421 (N_18421,N_10711,N_13986);
nor U18422 (N_18422,N_14161,N_10460);
nor U18423 (N_18423,N_11913,N_13861);
or U18424 (N_18424,N_14595,N_10013);
or U18425 (N_18425,N_10111,N_10939);
nand U18426 (N_18426,N_13893,N_13533);
or U18427 (N_18427,N_14382,N_12901);
or U18428 (N_18428,N_14794,N_10638);
nand U18429 (N_18429,N_14648,N_11424);
or U18430 (N_18430,N_11699,N_10132);
nand U18431 (N_18431,N_13267,N_14638);
or U18432 (N_18432,N_12717,N_14429);
or U18433 (N_18433,N_13193,N_12761);
or U18434 (N_18434,N_12313,N_13265);
nand U18435 (N_18435,N_14539,N_10361);
or U18436 (N_18436,N_12853,N_14234);
nand U18437 (N_18437,N_13555,N_10396);
or U18438 (N_18438,N_14788,N_14610);
and U18439 (N_18439,N_14548,N_12661);
or U18440 (N_18440,N_13252,N_13043);
nand U18441 (N_18441,N_14939,N_11368);
nor U18442 (N_18442,N_14569,N_13664);
and U18443 (N_18443,N_11405,N_10436);
and U18444 (N_18444,N_12128,N_12609);
or U18445 (N_18445,N_11232,N_12071);
and U18446 (N_18446,N_14341,N_10909);
nor U18447 (N_18447,N_10296,N_13106);
or U18448 (N_18448,N_13588,N_14588);
nand U18449 (N_18449,N_12451,N_14209);
nor U18450 (N_18450,N_12610,N_12686);
nor U18451 (N_18451,N_13366,N_14442);
and U18452 (N_18452,N_13977,N_13791);
and U18453 (N_18453,N_10322,N_13636);
nand U18454 (N_18454,N_12874,N_10315);
xnor U18455 (N_18455,N_10419,N_13437);
or U18456 (N_18456,N_10084,N_14062);
nor U18457 (N_18457,N_13193,N_10413);
and U18458 (N_18458,N_13544,N_13846);
nor U18459 (N_18459,N_13756,N_13413);
nand U18460 (N_18460,N_14457,N_12423);
nand U18461 (N_18461,N_11351,N_14021);
nor U18462 (N_18462,N_14422,N_13300);
nand U18463 (N_18463,N_12200,N_10080);
nand U18464 (N_18464,N_14040,N_13303);
and U18465 (N_18465,N_13766,N_10641);
nor U18466 (N_18466,N_10292,N_11542);
nand U18467 (N_18467,N_11643,N_14326);
nor U18468 (N_18468,N_11977,N_13888);
nor U18469 (N_18469,N_14134,N_12800);
or U18470 (N_18470,N_12233,N_14916);
nor U18471 (N_18471,N_12812,N_14523);
nand U18472 (N_18472,N_13613,N_10312);
nand U18473 (N_18473,N_10589,N_14563);
xnor U18474 (N_18474,N_10987,N_10135);
and U18475 (N_18475,N_13208,N_14925);
or U18476 (N_18476,N_10762,N_12646);
or U18477 (N_18477,N_11607,N_11946);
or U18478 (N_18478,N_11400,N_13002);
or U18479 (N_18479,N_10758,N_14601);
nor U18480 (N_18480,N_13745,N_14311);
nor U18481 (N_18481,N_13860,N_10919);
or U18482 (N_18482,N_13590,N_14117);
and U18483 (N_18483,N_14970,N_11369);
nand U18484 (N_18484,N_14388,N_13836);
and U18485 (N_18485,N_14084,N_10007);
and U18486 (N_18486,N_13950,N_14212);
or U18487 (N_18487,N_14491,N_12971);
and U18488 (N_18488,N_14386,N_14666);
and U18489 (N_18489,N_14757,N_14736);
nand U18490 (N_18490,N_12948,N_10480);
nand U18491 (N_18491,N_12504,N_12255);
or U18492 (N_18492,N_11270,N_14583);
xor U18493 (N_18493,N_10990,N_13582);
nor U18494 (N_18494,N_10740,N_12542);
or U18495 (N_18495,N_13269,N_11325);
and U18496 (N_18496,N_14553,N_11198);
nand U18497 (N_18497,N_14528,N_13539);
nand U18498 (N_18498,N_11075,N_10994);
or U18499 (N_18499,N_13145,N_13503);
nand U18500 (N_18500,N_11647,N_10445);
or U18501 (N_18501,N_13382,N_12056);
nor U18502 (N_18502,N_10867,N_12423);
nand U18503 (N_18503,N_11330,N_11942);
nor U18504 (N_18504,N_14299,N_13496);
xnor U18505 (N_18505,N_14587,N_11982);
nor U18506 (N_18506,N_11393,N_13838);
xor U18507 (N_18507,N_13020,N_14292);
and U18508 (N_18508,N_14915,N_12157);
nor U18509 (N_18509,N_11404,N_10827);
nor U18510 (N_18510,N_11336,N_13716);
nor U18511 (N_18511,N_13760,N_12135);
or U18512 (N_18512,N_13602,N_13604);
nor U18513 (N_18513,N_12210,N_12350);
and U18514 (N_18514,N_10943,N_13653);
or U18515 (N_18515,N_12698,N_10300);
xor U18516 (N_18516,N_11199,N_10772);
nand U18517 (N_18517,N_13144,N_14012);
and U18518 (N_18518,N_11755,N_13246);
nor U18519 (N_18519,N_13679,N_13516);
xor U18520 (N_18520,N_12468,N_13776);
and U18521 (N_18521,N_12256,N_13754);
or U18522 (N_18522,N_12277,N_14281);
or U18523 (N_18523,N_11098,N_12032);
and U18524 (N_18524,N_12972,N_11248);
or U18525 (N_18525,N_11812,N_10242);
or U18526 (N_18526,N_11446,N_12770);
nand U18527 (N_18527,N_14357,N_14830);
nor U18528 (N_18528,N_11757,N_14720);
nand U18529 (N_18529,N_12589,N_11907);
xor U18530 (N_18530,N_10901,N_14815);
xnor U18531 (N_18531,N_10091,N_12037);
and U18532 (N_18532,N_12878,N_11860);
xnor U18533 (N_18533,N_10695,N_10006);
nor U18534 (N_18534,N_10472,N_14243);
nand U18535 (N_18535,N_11893,N_12642);
or U18536 (N_18536,N_10524,N_14143);
and U18537 (N_18537,N_10806,N_10109);
xor U18538 (N_18538,N_12578,N_13360);
or U18539 (N_18539,N_12580,N_14994);
nor U18540 (N_18540,N_10623,N_10652);
or U18541 (N_18541,N_10603,N_12586);
nor U18542 (N_18542,N_14129,N_12937);
nand U18543 (N_18543,N_13957,N_10576);
or U18544 (N_18544,N_13273,N_13537);
and U18545 (N_18545,N_13899,N_11046);
and U18546 (N_18546,N_11641,N_12708);
and U18547 (N_18547,N_10131,N_13932);
and U18548 (N_18548,N_14412,N_11180);
nand U18549 (N_18549,N_13233,N_13208);
and U18550 (N_18550,N_12186,N_10242);
or U18551 (N_18551,N_11582,N_14564);
nor U18552 (N_18552,N_10724,N_10393);
or U18553 (N_18553,N_10692,N_11276);
and U18554 (N_18554,N_10402,N_12838);
nor U18555 (N_18555,N_12745,N_10710);
nand U18556 (N_18556,N_12972,N_11799);
nor U18557 (N_18557,N_13184,N_11340);
or U18558 (N_18558,N_12940,N_11504);
and U18559 (N_18559,N_10483,N_10271);
nand U18560 (N_18560,N_10324,N_10649);
and U18561 (N_18561,N_12503,N_11049);
nand U18562 (N_18562,N_14901,N_11691);
nand U18563 (N_18563,N_10380,N_13346);
nor U18564 (N_18564,N_11283,N_12911);
nor U18565 (N_18565,N_11932,N_10523);
nor U18566 (N_18566,N_11994,N_12132);
and U18567 (N_18567,N_13201,N_11624);
or U18568 (N_18568,N_14613,N_12519);
nor U18569 (N_18569,N_14122,N_11787);
and U18570 (N_18570,N_13854,N_13813);
nand U18571 (N_18571,N_11534,N_11028);
nand U18572 (N_18572,N_13043,N_14146);
and U18573 (N_18573,N_14269,N_10764);
and U18574 (N_18574,N_10225,N_11922);
or U18575 (N_18575,N_12998,N_12008);
xor U18576 (N_18576,N_14386,N_11561);
or U18577 (N_18577,N_11399,N_11313);
nor U18578 (N_18578,N_13539,N_11649);
nor U18579 (N_18579,N_13748,N_12872);
xnor U18580 (N_18580,N_12217,N_13221);
and U18581 (N_18581,N_11070,N_14850);
xnor U18582 (N_18582,N_12019,N_14068);
and U18583 (N_18583,N_13900,N_12918);
and U18584 (N_18584,N_11548,N_10537);
nor U18585 (N_18585,N_10209,N_12282);
nand U18586 (N_18586,N_10450,N_13620);
and U18587 (N_18587,N_11720,N_12096);
nor U18588 (N_18588,N_11823,N_13457);
nand U18589 (N_18589,N_11360,N_14390);
nor U18590 (N_18590,N_12945,N_14973);
nor U18591 (N_18591,N_13242,N_13574);
or U18592 (N_18592,N_14768,N_13957);
or U18593 (N_18593,N_14756,N_10523);
and U18594 (N_18594,N_10662,N_11897);
and U18595 (N_18595,N_12953,N_11698);
and U18596 (N_18596,N_10668,N_13417);
and U18597 (N_18597,N_14460,N_11611);
nand U18598 (N_18598,N_13083,N_12533);
nand U18599 (N_18599,N_14436,N_10331);
nand U18600 (N_18600,N_14609,N_13040);
nand U18601 (N_18601,N_13387,N_14512);
nor U18602 (N_18602,N_11168,N_12882);
nand U18603 (N_18603,N_12442,N_10123);
or U18604 (N_18604,N_11388,N_13887);
or U18605 (N_18605,N_11088,N_10514);
nor U18606 (N_18606,N_11913,N_11652);
and U18607 (N_18607,N_14173,N_12723);
nor U18608 (N_18608,N_13639,N_13762);
nand U18609 (N_18609,N_11997,N_12242);
or U18610 (N_18610,N_11209,N_10978);
nand U18611 (N_18611,N_13521,N_13847);
nor U18612 (N_18612,N_10129,N_11908);
nor U18613 (N_18613,N_11109,N_10867);
or U18614 (N_18614,N_14316,N_14422);
nand U18615 (N_18615,N_11472,N_12211);
and U18616 (N_18616,N_12972,N_10020);
and U18617 (N_18617,N_14390,N_10878);
nand U18618 (N_18618,N_10115,N_12558);
nand U18619 (N_18619,N_10659,N_10858);
nand U18620 (N_18620,N_10346,N_13847);
xor U18621 (N_18621,N_13607,N_11107);
or U18622 (N_18622,N_13026,N_12651);
nand U18623 (N_18623,N_12918,N_11665);
nand U18624 (N_18624,N_14271,N_14732);
nor U18625 (N_18625,N_13247,N_13709);
nand U18626 (N_18626,N_12989,N_11821);
and U18627 (N_18627,N_14360,N_13367);
and U18628 (N_18628,N_12609,N_13929);
or U18629 (N_18629,N_10311,N_12065);
and U18630 (N_18630,N_10676,N_10599);
nor U18631 (N_18631,N_11205,N_11841);
nand U18632 (N_18632,N_10761,N_12399);
nand U18633 (N_18633,N_13770,N_10326);
nor U18634 (N_18634,N_14174,N_14706);
nor U18635 (N_18635,N_13339,N_14708);
xnor U18636 (N_18636,N_11658,N_13926);
or U18637 (N_18637,N_13517,N_10049);
xor U18638 (N_18638,N_13708,N_10871);
or U18639 (N_18639,N_10437,N_10533);
nand U18640 (N_18640,N_12916,N_11087);
nand U18641 (N_18641,N_11579,N_14210);
or U18642 (N_18642,N_10572,N_11835);
xor U18643 (N_18643,N_12863,N_10208);
or U18644 (N_18644,N_12596,N_14247);
nand U18645 (N_18645,N_13192,N_14688);
nor U18646 (N_18646,N_11134,N_13755);
nand U18647 (N_18647,N_12431,N_10185);
and U18648 (N_18648,N_11270,N_14286);
or U18649 (N_18649,N_10642,N_10121);
nor U18650 (N_18650,N_14759,N_12277);
nor U18651 (N_18651,N_13452,N_12750);
nand U18652 (N_18652,N_12099,N_13002);
or U18653 (N_18653,N_10447,N_13388);
and U18654 (N_18654,N_10500,N_14891);
or U18655 (N_18655,N_12328,N_14916);
or U18656 (N_18656,N_11229,N_11913);
nand U18657 (N_18657,N_10368,N_11074);
nand U18658 (N_18658,N_13618,N_12003);
or U18659 (N_18659,N_13486,N_11115);
nor U18660 (N_18660,N_12727,N_12689);
nand U18661 (N_18661,N_11952,N_13982);
nor U18662 (N_18662,N_11301,N_14078);
or U18663 (N_18663,N_13003,N_13859);
and U18664 (N_18664,N_14282,N_14544);
nand U18665 (N_18665,N_12029,N_13737);
nand U18666 (N_18666,N_11473,N_10034);
nor U18667 (N_18667,N_10528,N_12136);
xnor U18668 (N_18668,N_10569,N_10784);
or U18669 (N_18669,N_10152,N_14963);
nand U18670 (N_18670,N_10984,N_13822);
xnor U18671 (N_18671,N_11944,N_12822);
or U18672 (N_18672,N_11974,N_11498);
or U18673 (N_18673,N_11402,N_12166);
nand U18674 (N_18674,N_13880,N_14579);
nand U18675 (N_18675,N_12548,N_12232);
or U18676 (N_18676,N_14047,N_10301);
xor U18677 (N_18677,N_12693,N_11758);
nand U18678 (N_18678,N_11835,N_11476);
and U18679 (N_18679,N_10896,N_12011);
or U18680 (N_18680,N_12453,N_10262);
and U18681 (N_18681,N_11523,N_10956);
and U18682 (N_18682,N_12437,N_12027);
and U18683 (N_18683,N_12222,N_14907);
or U18684 (N_18684,N_13014,N_13843);
or U18685 (N_18685,N_14434,N_11216);
nor U18686 (N_18686,N_11672,N_11417);
nand U18687 (N_18687,N_12455,N_10757);
and U18688 (N_18688,N_11527,N_13519);
and U18689 (N_18689,N_12514,N_11338);
nor U18690 (N_18690,N_12647,N_13837);
and U18691 (N_18691,N_13598,N_11102);
nand U18692 (N_18692,N_12297,N_12913);
and U18693 (N_18693,N_14634,N_10412);
nor U18694 (N_18694,N_12026,N_10782);
nand U18695 (N_18695,N_14473,N_11389);
nor U18696 (N_18696,N_14140,N_14500);
nor U18697 (N_18697,N_14222,N_12656);
xor U18698 (N_18698,N_13172,N_13296);
and U18699 (N_18699,N_11719,N_11809);
xnor U18700 (N_18700,N_12919,N_12513);
nor U18701 (N_18701,N_10941,N_12828);
nor U18702 (N_18702,N_14112,N_13134);
nand U18703 (N_18703,N_13868,N_12801);
or U18704 (N_18704,N_13951,N_14491);
xnor U18705 (N_18705,N_13150,N_12281);
and U18706 (N_18706,N_14321,N_11327);
or U18707 (N_18707,N_10658,N_12262);
or U18708 (N_18708,N_11301,N_14651);
and U18709 (N_18709,N_10258,N_13991);
or U18710 (N_18710,N_14129,N_13588);
nand U18711 (N_18711,N_14643,N_13722);
or U18712 (N_18712,N_14817,N_11847);
nor U18713 (N_18713,N_11545,N_10466);
or U18714 (N_18714,N_14546,N_11736);
nor U18715 (N_18715,N_10334,N_11095);
nor U18716 (N_18716,N_10436,N_12397);
xor U18717 (N_18717,N_11390,N_12715);
and U18718 (N_18718,N_13208,N_13569);
nor U18719 (N_18719,N_10669,N_11034);
nor U18720 (N_18720,N_11469,N_10118);
or U18721 (N_18721,N_12829,N_11221);
xor U18722 (N_18722,N_11853,N_11534);
or U18723 (N_18723,N_10955,N_11417);
or U18724 (N_18724,N_10930,N_13456);
nor U18725 (N_18725,N_10365,N_12822);
nor U18726 (N_18726,N_13125,N_10376);
nand U18727 (N_18727,N_13882,N_11774);
nor U18728 (N_18728,N_10738,N_13554);
or U18729 (N_18729,N_11305,N_14854);
xnor U18730 (N_18730,N_13967,N_11262);
nor U18731 (N_18731,N_12268,N_11918);
nor U18732 (N_18732,N_14674,N_14521);
nand U18733 (N_18733,N_10049,N_14608);
and U18734 (N_18734,N_13051,N_14769);
or U18735 (N_18735,N_12915,N_11908);
xor U18736 (N_18736,N_10540,N_13878);
or U18737 (N_18737,N_11085,N_11410);
nor U18738 (N_18738,N_10860,N_13642);
or U18739 (N_18739,N_10897,N_13577);
xnor U18740 (N_18740,N_13802,N_13816);
nor U18741 (N_18741,N_12071,N_13972);
and U18742 (N_18742,N_11604,N_13948);
nor U18743 (N_18743,N_14027,N_11478);
and U18744 (N_18744,N_10818,N_10229);
nor U18745 (N_18745,N_14543,N_13171);
and U18746 (N_18746,N_13955,N_14582);
nand U18747 (N_18747,N_10184,N_10448);
and U18748 (N_18748,N_13105,N_11829);
nor U18749 (N_18749,N_10223,N_14685);
or U18750 (N_18750,N_11769,N_10167);
and U18751 (N_18751,N_12200,N_12416);
nand U18752 (N_18752,N_10782,N_11733);
nor U18753 (N_18753,N_11736,N_12873);
or U18754 (N_18754,N_10854,N_10039);
and U18755 (N_18755,N_14139,N_11565);
nor U18756 (N_18756,N_10526,N_11567);
and U18757 (N_18757,N_12442,N_13441);
or U18758 (N_18758,N_11925,N_11241);
nand U18759 (N_18759,N_12539,N_14400);
and U18760 (N_18760,N_13325,N_11142);
nand U18761 (N_18761,N_11910,N_11983);
or U18762 (N_18762,N_11990,N_10433);
or U18763 (N_18763,N_13736,N_13708);
nand U18764 (N_18764,N_10981,N_11107);
xnor U18765 (N_18765,N_13294,N_11802);
nor U18766 (N_18766,N_10337,N_10671);
and U18767 (N_18767,N_11656,N_12372);
or U18768 (N_18768,N_13618,N_13597);
xor U18769 (N_18769,N_14722,N_13550);
nor U18770 (N_18770,N_10981,N_14870);
or U18771 (N_18771,N_12446,N_13041);
and U18772 (N_18772,N_10418,N_11382);
nand U18773 (N_18773,N_11794,N_13112);
nand U18774 (N_18774,N_11106,N_11064);
xor U18775 (N_18775,N_12705,N_13071);
or U18776 (N_18776,N_12716,N_13464);
and U18777 (N_18777,N_14656,N_13206);
nor U18778 (N_18778,N_13909,N_12598);
or U18779 (N_18779,N_12812,N_10079);
or U18780 (N_18780,N_12448,N_13261);
nand U18781 (N_18781,N_14069,N_12549);
or U18782 (N_18782,N_13465,N_10039);
and U18783 (N_18783,N_10876,N_10370);
nand U18784 (N_18784,N_14555,N_11978);
nand U18785 (N_18785,N_10572,N_12453);
and U18786 (N_18786,N_13038,N_11290);
and U18787 (N_18787,N_10299,N_14178);
or U18788 (N_18788,N_10752,N_11751);
nor U18789 (N_18789,N_10429,N_12355);
nor U18790 (N_18790,N_13075,N_10294);
nor U18791 (N_18791,N_13753,N_10504);
or U18792 (N_18792,N_12573,N_14292);
nand U18793 (N_18793,N_10041,N_11514);
nand U18794 (N_18794,N_12114,N_13142);
nor U18795 (N_18795,N_12296,N_12092);
nand U18796 (N_18796,N_12688,N_11593);
and U18797 (N_18797,N_12776,N_14609);
nor U18798 (N_18798,N_11244,N_12453);
xnor U18799 (N_18799,N_13359,N_11817);
nand U18800 (N_18800,N_12340,N_10646);
nor U18801 (N_18801,N_12344,N_13776);
and U18802 (N_18802,N_14757,N_12441);
nor U18803 (N_18803,N_14418,N_13915);
and U18804 (N_18804,N_10887,N_11175);
xnor U18805 (N_18805,N_12366,N_13318);
nor U18806 (N_18806,N_14700,N_14763);
nor U18807 (N_18807,N_13357,N_14149);
nor U18808 (N_18808,N_14544,N_10925);
nand U18809 (N_18809,N_12640,N_14910);
nor U18810 (N_18810,N_11998,N_12684);
or U18811 (N_18811,N_14780,N_11056);
or U18812 (N_18812,N_12891,N_13904);
nor U18813 (N_18813,N_13424,N_14024);
nor U18814 (N_18814,N_11427,N_10389);
or U18815 (N_18815,N_10200,N_14804);
or U18816 (N_18816,N_11420,N_14734);
nor U18817 (N_18817,N_13756,N_10142);
or U18818 (N_18818,N_10206,N_14683);
nor U18819 (N_18819,N_13166,N_14116);
nand U18820 (N_18820,N_10689,N_12805);
nor U18821 (N_18821,N_11277,N_11850);
and U18822 (N_18822,N_10228,N_13537);
nor U18823 (N_18823,N_11261,N_13544);
and U18824 (N_18824,N_12736,N_14904);
and U18825 (N_18825,N_12008,N_11261);
nor U18826 (N_18826,N_11695,N_13917);
xnor U18827 (N_18827,N_12197,N_13770);
or U18828 (N_18828,N_13501,N_14226);
nor U18829 (N_18829,N_10088,N_13616);
nand U18830 (N_18830,N_12206,N_14643);
nor U18831 (N_18831,N_11678,N_13013);
and U18832 (N_18832,N_11264,N_14383);
nand U18833 (N_18833,N_12972,N_14373);
nor U18834 (N_18834,N_13043,N_12313);
nor U18835 (N_18835,N_13196,N_13357);
nand U18836 (N_18836,N_14699,N_11636);
nor U18837 (N_18837,N_13301,N_12634);
nor U18838 (N_18838,N_11184,N_12734);
xor U18839 (N_18839,N_12126,N_10713);
nand U18840 (N_18840,N_12701,N_12845);
or U18841 (N_18841,N_10438,N_12734);
or U18842 (N_18842,N_13615,N_11408);
and U18843 (N_18843,N_10926,N_10869);
nand U18844 (N_18844,N_14970,N_12836);
nor U18845 (N_18845,N_11155,N_13772);
nand U18846 (N_18846,N_13771,N_14086);
or U18847 (N_18847,N_11602,N_13274);
and U18848 (N_18848,N_14105,N_13992);
nand U18849 (N_18849,N_14376,N_10013);
and U18850 (N_18850,N_11535,N_10079);
nor U18851 (N_18851,N_13849,N_12043);
nand U18852 (N_18852,N_11803,N_13078);
and U18853 (N_18853,N_10885,N_14042);
nand U18854 (N_18854,N_11587,N_12262);
and U18855 (N_18855,N_14226,N_12878);
or U18856 (N_18856,N_10449,N_11307);
nor U18857 (N_18857,N_11848,N_11090);
and U18858 (N_18858,N_12085,N_10683);
nor U18859 (N_18859,N_14178,N_11294);
nor U18860 (N_18860,N_12417,N_14693);
nand U18861 (N_18861,N_12315,N_13568);
and U18862 (N_18862,N_12619,N_10284);
xor U18863 (N_18863,N_13404,N_11745);
nor U18864 (N_18864,N_11292,N_11586);
xnor U18865 (N_18865,N_11592,N_11244);
or U18866 (N_18866,N_10591,N_11184);
or U18867 (N_18867,N_14225,N_13555);
nor U18868 (N_18868,N_12879,N_10682);
nand U18869 (N_18869,N_11552,N_14722);
nand U18870 (N_18870,N_12312,N_13568);
nor U18871 (N_18871,N_12504,N_13401);
xnor U18872 (N_18872,N_12969,N_12613);
or U18873 (N_18873,N_12005,N_14924);
nand U18874 (N_18874,N_11229,N_12505);
nor U18875 (N_18875,N_13319,N_12100);
nor U18876 (N_18876,N_10099,N_13138);
nor U18877 (N_18877,N_10761,N_12620);
xnor U18878 (N_18878,N_13096,N_11397);
nor U18879 (N_18879,N_11204,N_13344);
nand U18880 (N_18880,N_12997,N_13473);
nand U18881 (N_18881,N_12622,N_11076);
and U18882 (N_18882,N_11602,N_14911);
nor U18883 (N_18883,N_14263,N_12884);
nand U18884 (N_18884,N_11982,N_11866);
nand U18885 (N_18885,N_13819,N_11284);
and U18886 (N_18886,N_10714,N_11601);
xor U18887 (N_18887,N_11094,N_13017);
nor U18888 (N_18888,N_11907,N_11826);
or U18889 (N_18889,N_10440,N_11251);
nor U18890 (N_18890,N_11528,N_13801);
xor U18891 (N_18891,N_13108,N_10204);
nand U18892 (N_18892,N_10729,N_12198);
and U18893 (N_18893,N_10971,N_10305);
nor U18894 (N_18894,N_14421,N_13836);
xor U18895 (N_18895,N_10888,N_10457);
nand U18896 (N_18896,N_14715,N_13530);
nor U18897 (N_18897,N_14030,N_14181);
nor U18898 (N_18898,N_12587,N_12150);
nand U18899 (N_18899,N_10433,N_12135);
nor U18900 (N_18900,N_11992,N_10027);
nor U18901 (N_18901,N_11430,N_10642);
or U18902 (N_18902,N_14085,N_14155);
nand U18903 (N_18903,N_12724,N_10707);
xnor U18904 (N_18904,N_11730,N_11792);
and U18905 (N_18905,N_10249,N_11642);
xnor U18906 (N_18906,N_12901,N_10962);
or U18907 (N_18907,N_13564,N_13859);
nor U18908 (N_18908,N_11773,N_10979);
and U18909 (N_18909,N_14447,N_10064);
nor U18910 (N_18910,N_13662,N_13824);
and U18911 (N_18911,N_11120,N_14031);
xor U18912 (N_18912,N_11991,N_13176);
or U18913 (N_18913,N_13500,N_13017);
and U18914 (N_18914,N_14472,N_14611);
nor U18915 (N_18915,N_14765,N_10174);
or U18916 (N_18916,N_11506,N_12155);
nor U18917 (N_18917,N_14948,N_13319);
or U18918 (N_18918,N_13783,N_14373);
nand U18919 (N_18919,N_12146,N_12776);
or U18920 (N_18920,N_10318,N_13264);
and U18921 (N_18921,N_10750,N_13414);
or U18922 (N_18922,N_13363,N_12517);
or U18923 (N_18923,N_10001,N_14831);
xnor U18924 (N_18924,N_14168,N_11358);
nor U18925 (N_18925,N_13643,N_12984);
nand U18926 (N_18926,N_10956,N_11348);
nor U18927 (N_18927,N_12163,N_14734);
and U18928 (N_18928,N_10610,N_12958);
nor U18929 (N_18929,N_14682,N_13277);
nand U18930 (N_18930,N_11203,N_11585);
or U18931 (N_18931,N_13427,N_10159);
nand U18932 (N_18932,N_10961,N_11540);
or U18933 (N_18933,N_12259,N_10264);
or U18934 (N_18934,N_11993,N_10042);
nand U18935 (N_18935,N_13295,N_14829);
nor U18936 (N_18936,N_11006,N_12927);
xnor U18937 (N_18937,N_11605,N_10177);
or U18938 (N_18938,N_14176,N_11509);
nor U18939 (N_18939,N_13029,N_12993);
and U18940 (N_18940,N_10331,N_11006);
nand U18941 (N_18941,N_10627,N_13287);
nand U18942 (N_18942,N_10470,N_10813);
and U18943 (N_18943,N_14423,N_13455);
nor U18944 (N_18944,N_13224,N_14744);
nand U18945 (N_18945,N_13236,N_10289);
or U18946 (N_18946,N_13541,N_12930);
nand U18947 (N_18947,N_11311,N_10799);
or U18948 (N_18948,N_14029,N_11319);
nand U18949 (N_18949,N_10070,N_11534);
nand U18950 (N_18950,N_11729,N_11317);
xor U18951 (N_18951,N_12333,N_13456);
nand U18952 (N_18952,N_11650,N_13696);
and U18953 (N_18953,N_12212,N_13418);
and U18954 (N_18954,N_12431,N_13566);
and U18955 (N_18955,N_13490,N_12199);
nand U18956 (N_18956,N_10099,N_11815);
nor U18957 (N_18957,N_14422,N_10922);
nand U18958 (N_18958,N_10525,N_10682);
nand U18959 (N_18959,N_10536,N_12164);
xnor U18960 (N_18960,N_11327,N_14836);
and U18961 (N_18961,N_11985,N_10561);
nand U18962 (N_18962,N_13438,N_12753);
nand U18963 (N_18963,N_14633,N_11310);
nor U18964 (N_18964,N_14371,N_14044);
nor U18965 (N_18965,N_11609,N_14714);
nor U18966 (N_18966,N_12628,N_11266);
nor U18967 (N_18967,N_13655,N_14777);
or U18968 (N_18968,N_10309,N_10060);
and U18969 (N_18969,N_13399,N_13071);
and U18970 (N_18970,N_14215,N_14227);
and U18971 (N_18971,N_11810,N_14582);
and U18972 (N_18972,N_10217,N_11894);
or U18973 (N_18973,N_12420,N_11616);
or U18974 (N_18974,N_10450,N_11082);
nand U18975 (N_18975,N_10447,N_12856);
or U18976 (N_18976,N_14692,N_14634);
nand U18977 (N_18977,N_13949,N_12919);
and U18978 (N_18978,N_14656,N_11471);
and U18979 (N_18979,N_12036,N_12819);
or U18980 (N_18980,N_14303,N_11963);
xnor U18981 (N_18981,N_13165,N_13588);
nor U18982 (N_18982,N_14886,N_12594);
nand U18983 (N_18983,N_13240,N_14474);
nand U18984 (N_18984,N_12332,N_12857);
nor U18985 (N_18985,N_12964,N_12535);
nand U18986 (N_18986,N_14655,N_14948);
nand U18987 (N_18987,N_13432,N_11707);
or U18988 (N_18988,N_13455,N_13947);
nor U18989 (N_18989,N_13653,N_14056);
nor U18990 (N_18990,N_11056,N_11531);
nor U18991 (N_18991,N_14419,N_11064);
nor U18992 (N_18992,N_14904,N_11502);
nor U18993 (N_18993,N_10631,N_14907);
and U18994 (N_18994,N_14284,N_10484);
and U18995 (N_18995,N_13569,N_11626);
nand U18996 (N_18996,N_13056,N_10488);
xor U18997 (N_18997,N_13850,N_12416);
nand U18998 (N_18998,N_11009,N_10890);
nand U18999 (N_18999,N_14229,N_12899);
nor U19000 (N_19000,N_11542,N_12851);
or U19001 (N_19001,N_13216,N_14057);
nor U19002 (N_19002,N_12580,N_14105);
or U19003 (N_19003,N_14727,N_10192);
or U19004 (N_19004,N_11648,N_13322);
and U19005 (N_19005,N_10972,N_13189);
nand U19006 (N_19006,N_14950,N_10073);
xor U19007 (N_19007,N_12800,N_10225);
xnor U19008 (N_19008,N_12084,N_14477);
nand U19009 (N_19009,N_13303,N_11908);
nor U19010 (N_19010,N_13846,N_11197);
and U19011 (N_19011,N_14518,N_14115);
and U19012 (N_19012,N_14904,N_11244);
and U19013 (N_19013,N_11328,N_14334);
and U19014 (N_19014,N_14026,N_10221);
and U19015 (N_19015,N_13569,N_12584);
or U19016 (N_19016,N_14228,N_14552);
nand U19017 (N_19017,N_12202,N_13097);
and U19018 (N_19018,N_14004,N_13395);
or U19019 (N_19019,N_10861,N_14392);
or U19020 (N_19020,N_10530,N_11262);
and U19021 (N_19021,N_12563,N_10813);
xnor U19022 (N_19022,N_11423,N_11754);
and U19023 (N_19023,N_14553,N_10462);
nor U19024 (N_19024,N_11630,N_10464);
nor U19025 (N_19025,N_12913,N_14722);
xor U19026 (N_19026,N_14684,N_11521);
nand U19027 (N_19027,N_10264,N_10941);
and U19028 (N_19028,N_14603,N_12306);
and U19029 (N_19029,N_13247,N_13653);
nand U19030 (N_19030,N_14368,N_11935);
or U19031 (N_19031,N_14312,N_12831);
nand U19032 (N_19032,N_10741,N_14379);
and U19033 (N_19033,N_14481,N_10261);
and U19034 (N_19034,N_12380,N_13131);
nand U19035 (N_19035,N_14189,N_10237);
nand U19036 (N_19036,N_14071,N_13817);
and U19037 (N_19037,N_11457,N_13603);
nand U19038 (N_19038,N_13561,N_10846);
nor U19039 (N_19039,N_12722,N_13917);
or U19040 (N_19040,N_13451,N_14108);
nand U19041 (N_19041,N_11261,N_14023);
nor U19042 (N_19042,N_12131,N_12614);
or U19043 (N_19043,N_14139,N_14326);
or U19044 (N_19044,N_14844,N_10830);
or U19045 (N_19045,N_12176,N_13773);
nor U19046 (N_19046,N_14101,N_13027);
and U19047 (N_19047,N_11012,N_10495);
nor U19048 (N_19048,N_11030,N_10041);
nand U19049 (N_19049,N_13397,N_10119);
and U19050 (N_19050,N_13590,N_13848);
or U19051 (N_19051,N_10156,N_14316);
or U19052 (N_19052,N_13541,N_10305);
or U19053 (N_19053,N_12839,N_14440);
or U19054 (N_19054,N_13821,N_11022);
and U19055 (N_19055,N_12277,N_12330);
xnor U19056 (N_19056,N_10777,N_10824);
nand U19057 (N_19057,N_13057,N_10412);
and U19058 (N_19058,N_11143,N_14447);
or U19059 (N_19059,N_10726,N_13341);
and U19060 (N_19060,N_13138,N_13882);
and U19061 (N_19061,N_10258,N_13691);
nor U19062 (N_19062,N_13079,N_11752);
or U19063 (N_19063,N_10259,N_14494);
nor U19064 (N_19064,N_12402,N_14706);
and U19065 (N_19065,N_10314,N_10729);
nand U19066 (N_19066,N_11201,N_13787);
nand U19067 (N_19067,N_14511,N_13700);
nor U19068 (N_19068,N_10626,N_11867);
nor U19069 (N_19069,N_10056,N_13962);
nand U19070 (N_19070,N_14118,N_11901);
and U19071 (N_19071,N_10690,N_11484);
nand U19072 (N_19072,N_13297,N_14673);
or U19073 (N_19073,N_14827,N_14020);
nor U19074 (N_19074,N_11606,N_11836);
and U19075 (N_19075,N_12509,N_10695);
nor U19076 (N_19076,N_13418,N_13647);
nand U19077 (N_19077,N_13957,N_10116);
or U19078 (N_19078,N_11554,N_13462);
or U19079 (N_19079,N_10758,N_13758);
and U19080 (N_19080,N_11791,N_10480);
or U19081 (N_19081,N_14235,N_10019);
nand U19082 (N_19082,N_14233,N_11135);
nor U19083 (N_19083,N_13215,N_10737);
nor U19084 (N_19084,N_10732,N_14572);
nand U19085 (N_19085,N_10995,N_12157);
and U19086 (N_19086,N_14454,N_10765);
or U19087 (N_19087,N_12053,N_13925);
or U19088 (N_19088,N_11765,N_10036);
nand U19089 (N_19089,N_11200,N_14217);
or U19090 (N_19090,N_13018,N_10587);
or U19091 (N_19091,N_12128,N_12397);
nor U19092 (N_19092,N_10251,N_11357);
nand U19093 (N_19093,N_13323,N_10840);
or U19094 (N_19094,N_11888,N_11973);
or U19095 (N_19095,N_13926,N_14673);
or U19096 (N_19096,N_14056,N_11764);
xor U19097 (N_19097,N_11648,N_12083);
and U19098 (N_19098,N_12296,N_13045);
nor U19099 (N_19099,N_14406,N_13674);
or U19100 (N_19100,N_13848,N_11775);
nor U19101 (N_19101,N_14922,N_11185);
or U19102 (N_19102,N_12157,N_14726);
xor U19103 (N_19103,N_12634,N_13870);
nor U19104 (N_19104,N_10266,N_13704);
and U19105 (N_19105,N_12672,N_13781);
nor U19106 (N_19106,N_10209,N_12621);
nor U19107 (N_19107,N_10715,N_14279);
or U19108 (N_19108,N_11800,N_14322);
and U19109 (N_19109,N_10126,N_10791);
or U19110 (N_19110,N_10268,N_12943);
or U19111 (N_19111,N_10384,N_10445);
xor U19112 (N_19112,N_13752,N_13489);
nand U19113 (N_19113,N_13448,N_12546);
or U19114 (N_19114,N_14865,N_14551);
or U19115 (N_19115,N_10825,N_11505);
or U19116 (N_19116,N_13506,N_13647);
xnor U19117 (N_19117,N_13655,N_14379);
nor U19118 (N_19118,N_14833,N_11711);
nor U19119 (N_19119,N_10575,N_11375);
and U19120 (N_19120,N_12023,N_14689);
nor U19121 (N_19121,N_10942,N_10392);
and U19122 (N_19122,N_14441,N_13733);
nand U19123 (N_19123,N_12103,N_12342);
nor U19124 (N_19124,N_10240,N_13862);
nand U19125 (N_19125,N_10317,N_10195);
nand U19126 (N_19126,N_10320,N_12087);
nor U19127 (N_19127,N_10426,N_14709);
and U19128 (N_19128,N_10899,N_11917);
or U19129 (N_19129,N_10246,N_11712);
and U19130 (N_19130,N_13689,N_14218);
nand U19131 (N_19131,N_10661,N_10194);
or U19132 (N_19132,N_12372,N_12773);
nand U19133 (N_19133,N_10974,N_11101);
nor U19134 (N_19134,N_11152,N_10121);
or U19135 (N_19135,N_12014,N_14285);
nor U19136 (N_19136,N_11903,N_10308);
and U19137 (N_19137,N_10272,N_10982);
and U19138 (N_19138,N_13098,N_12171);
and U19139 (N_19139,N_14220,N_14345);
and U19140 (N_19140,N_10719,N_14376);
and U19141 (N_19141,N_14373,N_14007);
nand U19142 (N_19142,N_10282,N_13677);
nor U19143 (N_19143,N_12703,N_10744);
nand U19144 (N_19144,N_12339,N_12490);
xnor U19145 (N_19145,N_11976,N_13158);
nor U19146 (N_19146,N_14535,N_13662);
and U19147 (N_19147,N_14961,N_11853);
nand U19148 (N_19148,N_11444,N_11873);
and U19149 (N_19149,N_10533,N_12787);
and U19150 (N_19150,N_11731,N_11370);
nor U19151 (N_19151,N_14668,N_14285);
and U19152 (N_19152,N_12150,N_13178);
or U19153 (N_19153,N_14688,N_13654);
or U19154 (N_19154,N_12265,N_11198);
nor U19155 (N_19155,N_10989,N_14311);
and U19156 (N_19156,N_14366,N_11351);
xor U19157 (N_19157,N_11461,N_13333);
nand U19158 (N_19158,N_13188,N_12186);
nand U19159 (N_19159,N_13555,N_11993);
or U19160 (N_19160,N_10358,N_11047);
nor U19161 (N_19161,N_14137,N_12207);
nand U19162 (N_19162,N_14826,N_13027);
or U19163 (N_19163,N_14012,N_10456);
nand U19164 (N_19164,N_13663,N_11582);
nor U19165 (N_19165,N_14307,N_12581);
or U19166 (N_19166,N_14394,N_14094);
and U19167 (N_19167,N_13692,N_10723);
xor U19168 (N_19168,N_11775,N_10443);
or U19169 (N_19169,N_12610,N_12699);
or U19170 (N_19170,N_10944,N_10906);
nand U19171 (N_19171,N_12323,N_12012);
nor U19172 (N_19172,N_13727,N_12476);
or U19173 (N_19173,N_14213,N_12859);
nand U19174 (N_19174,N_13045,N_12840);
or U19175 (N_19175,N_14358,N_11428);
or U19176 (N_19176,N_11260,N_11393);
and U19177 (N_19177,N_11671,N_14076);
xnor U19178 (N_19178,N_11435,N_14127);
nand U19179 (N_19179,N_10767,N_14261);
nor U19180 (N_19180,N_11157,N_14946);
and U19181 (N_19181,N_10842,N_13833);
or U19182 (N_19182,N_12211,N_14356);
nor U19183 (N_19183,N_10055,N_13096);
nor U19184 (N_19184,N_13287,N_12215);
nor U19185 (N_19185,N_12160,N_13580);
and U19186 (N_19186,N_14372,N_12957);
nand U19187 (N_19187,N_12710,N_11206);
nor U19188 (N_19188,N_13380,N_10815);
and U19189 (N_19189,N_10525,N_11937);
xor U19190 (N_19190,N_11011,N_13305);
or U19191 (N_19191,N_10003,N_11621);
nor U19192 (N_19192,N_10296,N_12702);
and U19193 (N_19193,N_14991,N_14986);
xnor U19194 (N_19194,N_10582,N_12372);
or U19195 (N_19195,N_13253,N_12819);
nor U19196 (N_19196,N_11400,N_12996);
and U19197 (N_19197,N_11760,N_13318);
and U19198 (N_19198,N_13176,N_11249);
or U19199 (N_19199,N_11202,N_14269);
and U19200 (N_19200,N_12089,N_13282);
or U19201 (N_19201,N_14163,N_12274);
xor U19202 (N_19202,N_13023,N_12329);
xnor U19203 (N_19203,N_14062,N_14438);
or U19204 (N_19204,N_12932,N_10596);
nand U19205 (N_19205,N_10856,N_11294);
or U19206 (N_19206,N_14416,N_11769);
nand U19207 (N_19207,N_10335,N_10528);
nand U19208 (N_19208,N_13338,N_10596);
and U19209 (N_19209,N_10629,N_12004);
nand U19210 (N_19210,N_10685,N_14721);
nor U19211 (N_19211,N_14625,N_14992);
or U19212 (N_19212,N_10814,N_14901);
and U19213 (N_19213,N_10574,N_13715);
nand U19214 (N_19214,N_12185,N_11726);
nor U19215 (N_19215,N_14580,N_14424);
nor U19216 (N_19216,N_14577,N_14011);
nand U19217 (N_19217,N_12538,N_12902);
nor U19218 (N_19218,N_11834,N_10423);
nand U19219 (N_19219,N_13687,N_11684);
or U19220 (N_19220,N_12849,N_12405);
nand U19221 (N_19221,N_11614,N_13821);
nand U19222 (N_19222,N_11131,N_10752);
nand U19223 (N_19223,N_13081,N_10229);
or U19224 (N_19224,N_13691,N_14931);
nor U19225 (N_19225,N_11269,N_14451);
xor U19226 (N_19226,N_10507,N_10017);
xor U19227 (N_19227,N_14741,N_14296);
xnor U19228 (N_19228,N_12182,N_12356);
nor U19229 (N_19229,N_10094,N_13450);
and U19230 (N_19230,N_10535,N_12649);
nand U19231 (N_19231,N_12592,N_11538);
nand U19232 (N_19232,N_13513,N_12719);
nor U19233 (N_19233,N_13089,N_14867);
xnor U19234 (N_19234,N_12982,N_13644);
xor U19235 (N_19235,N_14717,N_11803);
and U19236 (N_19236,N_13972,N_10445);
nor U19237 (N_19237,N_12132,N_13742);
or U19238 (N_19238,N_11319,N_10886);
nor U19239 (N_19239,N_13357,N_11714);
nand U19240 (N_19240,N_11869,N_11682);
xnor U19241 (N_19241,N_11249,N_12645);
nor U19242 (N_19242,N_12484,N_14875);
nand U19243 (N_19243,N_13800,N_11059);
and U19244 (N_19244,N_10842,N_14159);
and U19245 (N_19245,N_14485,N_13106);
or U19246 (N_19246,N_12847,N_14428);
and U19247 (N_19247,N_13109,N_11132);
and U19248 (N_19248,N_12417,N_14938);
nand U19249 (N_19249,N_10920,N_11398);
or U19250 (N_19250,N_12724,N_12687);
nor U19251 (N_19251,N_13274,N_11355);
nand U19252 (N_19252,N_14177,N_11679);
nor U19253 (N_19253,N_12380,N_11247);
and U19254 (N_19254,N_12677,N_14998);
xnor U19255 (N_19255,N_11211,N_14095);
nand U19256 (N_19256,N_12389,N_13247);
or U19257 (N_19257,N_14769,N_11485);
and U19258 (N_19258,N_13942,N_13670);
or U19259 (N_19259,N_11250,N_12714);
nor U19260 (N_19260,N_11651,N_14113);
or U19261 (N_19261,N_14876,N_13394);
and U19262 (N_19262,N_12326,N_14877);
and U19263 (N_19263,N_11610,N_14627);
nand U19264 (N_19264,N_12356,N_10679);
xor U19265 (N_19265,N_12696,N_11558);
nand U19266 (N_19266,N_10272,N_14203);
nor U19267 (N_19267,N_12171,N_10291);
and U19268 (N_19268,N_10294,N_10072);
or U19269 (N_19269,N_11090,N_11093);
nor U19270 (N_19270,N_10550,N_11664);
nor U19271 (N_19271,N_10137,N_13059);
nand U19272 (N_19272,N_12238,N_11012);
or U19273 (N_19273,N_14750,N_13125);
nand U19274 (N_19274,N_14904,N_13995);
nand U19275 (N_19275,N_13169,N_10009);
and U19276 (N_19276,N_14254,N_12253);
and U19277 (N_19277,N_10415,N_11823);
nor U19278 (N_19278,N_14770,N_14805);
nand U19279 (N_19279,N_13228,N_13666);
and U19280 (N_19280,N_12480,N_10061);
and U19281 (N_19281,N_14305,N_13315);
and U19282 (N_19282,N_11918,N_11986);
or U19283 (N_19283,N_14546,N_13580);
or U19284 (N_19284,N_14185,N_11692);
or U19285 (N_19285,N_10686,N_13821);
nand U19286 (N_19286,N_12948,N_12095);
nand U19287 (N_19287,N_12377,N_14423);
nand U19288 (N_19288,N_10957,N_12439);
nand U19289 (N_19289,N_13138,N_14403);
and U19290 (N_19290,N_11846,N_14690);
nand U19291 (N_19291,N_10884,N_11539);
or U19292 (N_19292,N_11857,N_14954);
nor U19293 (N_19293,N_10715,N_11013);
and U19294 (N_19294,N_10734,N_13936);
or U19295 (N_19295,N_10213,N_13814);
and U19296 (N_19296,N_11600,N_12892);
nand U19297 (N_19297,N_12887,N_11142);
or U19298 (N_19298,N_13985,N_13821);
and U19299 (N_19299,N_12261,N_11688);
nor U19300 (N_19300,N_14718,N_11301);
xor U19301 (N_19301,N_14365,N_14752);
or U19302 (N_19302,N_14826,N_13998);
nor U19303 (N_19303,N_10258,N_14152);
nand U19304 (N_19304,N_13705,N_10372);
xnor U19305 (N_19305,N_14673,N_13168);
or U19306 (N_19306,N_12998,N_14019);
nand U19307 (N_19307,N_11188,N_14368);
nor U19308 (N_19308,N_12413,N_10023);
or U19309 (N_19309,N_11036,N_13838);
nand U19310 (N_19310,N_12692,N_13105);
or U19311 (N_19311,N_12478,N_14220);
or U19312 (N_19312,N_14841,N_11058);
and U19313 (N_19313,N_14041,N_12889);
nand U19314 (N_19314,N_14420,N_14373);
or U19315 (N_19315,N_13490,N_10522);
nand U19316 (N_19316,N_13543,N_12934);
nand U19317 (N_19317,N_14345,N_10735);
or U19318 (N_19318,N_10303,N_12534);
nand U19319 (N_19319,N_14315,N_11639);
nor U19320 (N_19320,N_10705,N_14608);
or U19321 (N_19321,N_12052,N_14198);
nor U19322 (N_19322,N_10578,N_14707);
nor U19323 (N_19323,N_13201,N_10644);
or U19324 (N_19324,N_13093,N_11199);
nor U19325 (N_19325,N_10587,N_13494);
nor U19326 (N_19326,N_13298,N_12450);
or U19327 (N_19327,N_10495,N_11442);
nor U19328 (N_19328,N_10304,N_10376);
nand U19329 (N_19329,N_11031,N_11164);
or U19330 (N_19330,N_10599,N_14032);
or U19331 (N_19331,N_10764,N_10385);
xor U19332 (N_19332,N_12862,N_12535);
xnor U19333 (N_19333,N_14007,N_13359);
xnor U19334 (N_19334,N_11783,N_10104);
xor U19335 (N_19335,N_10936,N_10965);
xnor U19336 (N_19336,N_13174,N_10338);
or U19337 (N_19337,N_10378,N_10274);
or U19338 (N_19338,N_13435,N_14275);
and U19339 (N_19339,N_10410,N_10207);
and U19340 (N_19340,N_14699,N_14257);
nor U19341 (N_19341,N_13038,N_10532);
and U19342 (N_19342,N_14403,N_13592);
nor U19343 (N_19343,N_13851,N_12878);
or U19344 (N_19344,N_11480,N_10201);
nand U19345 (N_19345,N_12224,N_13377);
nand U19346 (N_19346,N_10760,N_11112);
nor U19347 (N_19347,N_12731,N_13451);
xor U19348 (N_19348,N_10701,N_12890);
nor U19349 (N_19349,N_11076,N_14879);
xor U19350 (N_19350,N_12980,N_10758);
nand U19351 (N_19351,N_14376,N_12634);
nand U19352 (N_19352,N_12568,N_12597);
nor U19353 (N_19353,N_11006,N_10586);
nor U19354 (N_19354,N_13476,N_14082);
xnor U19355 (N_19355,N_14650,N_11708);
nand U19356 (N_19356,N_12169,N_12465);
and U19357 (N_19357,N_11176,N_13731);
nor U19358 (N_19358,N_11078,N_10697);
nand U19359 (N_19359,N_14489,N_12316);
nand U19360 (N_19360,N_11123,N_12887);
nor U19361 (N_19361,N_10625,N_13189);
nor U19362 (N_19362,N_14550,N_10156);
or U19363 (N_19363,N_10563,N_12935);
or U19364 (N_19364,N_14378,N_12804);
nor U19365 (N_19365,N_11640,N_14108);
and U19366 (N_19366,N_12302,N_10234);
nand U19367 (N_19367,N_14476,N_13176);
or U19368 (N_19368,N_11095,N_12235);
and U19369 (N_19369,N_12679,N_11900);
or U19370 (N_19370,N_12039,N_14371);
nor U19371 (N_19371,N_12554,N_11301);
nand U19372 (N_19372,N_12725,N_11188);
or U19373 (N_19373,N_12417,N_13590);
or U19374 (N_19374,N_12793,N_13432);
and U19375 (N_19375,N_12895,N_12864);
nand U19376 (N_19376,N_12756,N_10356);
nand U19377 (N_19377,N_12815,N_12324);
or U19378 (N_19378,N_10699,N_13638);
nand U19379 (N_19379,N_13045,N_10341);
xor U19380 (N_19380,N_11942,N_14808);
and U19381 (N_19381,N_13012,N_10374);
xnor U19382 (N_19382,N_14259,N_14173);
or U19383 (N_19383,N_14931,N_10398);
nand U19384 (N_19384,N_14896,N_14658);
or U19385 (N_19385,N_12374,N_14370);
or U19386 (N_19386,N_11480,N_13924);
xor U19387 (N_19387,N_13996,N_10660);
and U19388 (N_19388,N_12073,N_13652);
xor U19389 (N_19389,N_10007,N_12115);
and U19390 (N_19390,N_13330,N_10434);
or U19391 (N_19391,N_14687,N_14510);
or U19392 (N_19392,N_12253,N_14977);
xor U19393 (N_19393,N_10096,N_13871);
xnor U19394 (N_19394,N_10441,N_14742);
or U19395 (N_19395,N_11786,N_14509);
nor U19396 (N_19396,N_12560,N_10514);
or U19397 (N_19397,N_12072,N_10768);
xor U19398 (N_19398,N_11104,N_10599);
or U19399 (N_19399,N_12029,N_11574);
nand U19400 (N_19400,N_11204,N_13433);
xor U19401 (N_19401,N_13333,N_13336);
or U19402 (N_19402,N_10205,N_12699);
and U19403 (N_19403,N_14517,N_14381);
nand U19404 (N_19404,N_12649,N_14372);
nor U19405 (N_19405,N_10605,N_14777);
nand U19406 (N_19406,N_11763,N_11021);
nor U19407 (N_19407,N_11329,N_13294);
and U19408 (N_19408,N_12728,N_12914);
and U19409 (N_19409,N_12275,N_13194);
and U19410 (N_19410,N_10426,N_10430);
or U19411 (N_19411,N_12380,N_12073);
nor U19412 (N_19412,N_10235,N_10638);
nor U19413 (N_19413,N_11992,N_11132);
nor U19414 (N_19414,N_14132,N_14604);
and U19415 (N_19415,N_12646,N_12710);
or U19416 (N_19416,N_10973,N_14933);
and U19417 (N_19417,N_14531,N_14389);
and U19418 (N_19418,N_10283,N_13712);
or U19419 (N_19419,N_12819,N_14568);
or U19420 (N_19420,N_10658,N_11486);
nand U19421 (N_19421,N_11437,N_11956);
or U19422 (N_19422,N_14983,N_10475);
or U19423 (N_19423,N_14283,N_10934);
and U19424 (N_19424,N_14754,N_13243);
nor U19425 (N_19425,N_11981,N_12293);
or U19426 (N_19426,N_14014,N_13313);
xnor U19427 (N_19427,N_11767,N_12893);
nand U19428 (N_19428,N_13237,N_10764);
and U19429 (N_19429,N_12820,N_14268);
and U19430 (N_19430,N_14793,N_14920);
nor U19431 (N_19431,N_12167,N_12049);
or U19432 (N_19432,N_14321,N_12139);
and U19433 (N_19433,N_11968,N_12005);
or U19434 (N_19434,N_13134,N_11312);
or U19435 (N_19435,N_10195,N_14860);
and U19436 (N_19436,N_14192,N_10962);
or U19437 (N_19437,N_10150,N_14836);
or U19438 (N_19438,N_10735,N_10945);
nand U19439 (N_19439,N_14229,N_13024);
nand U19440 (N_19440,N_11666,N_13624);
nand U19441 (N_19441,N_10397,N_14288);
xnor U19442 (N_19442,N_13523,N_13907);
nand U19443 (N_19443,N_11091,N_12194);
or U19444 (N_19444,N_14434,N_14213);
and U19445 (N_19445,N_14965,N_10998);
nor U19446 (N_19446,N_13620,N_10703);
nor U19447 (N_19447,N_10025,N_11360);
and U19448 (N_19448,N_14241,N_13314);
or U19449 (N_19449,N_11099,N_12602);
or U19450 (N_19450,N_14237,N_11398);
nor U19451 (N_19451,N_10699,N_12389);
or U19452 (N_19452,N_11563,N_13323);
xnor U19453 (N_19453,N_10479,N_11736);
or U19454 (N_19454,N_14321,N_10676);
or U19455 (N_19455,N_13861,N_10586);
nor U19456 (N_19456,N_12985,N_12720);
nor U19457 (N_19457,N_11581,N_12089);
nand U19458 (N_19458,N_14096,N_14850);
nand U19459 (N_19459,N_10793,N_12859);
xor U19460 (N_19460,N_14798,N_11631);
nand U19461 (N_19461,N_12953,N_11668);
xor U19462 (N_19462,N_13663,N_13397);
nand U19463 (N_19463,N_10457,N_14830);
or U19464 (N_19464,N_12534,N_11125);
xnor U19465 (N_19465,N_12322,N_12932);
nand U19466 (N_19466,N_14897,N_14396);
or U19467 (N_19467,N_13153,N_14316);
xnor U19468 (N_19468,N_14645,N_12457);
and U19469 (N_19469,N_12012,N_14021);
or U19470 (N_19470,N_11535,N_13512);
xor U19471 (N_19471,N_13017,N_13842);
xnor U19472 (N_19472,N_10637,N_12930);
nor U19473 (N_19473,N_11179,N_14679);
nand U19474 (N_19474,N_11927,N_14444);
or U19475 (N_19475,N_10607,N_14980);
or U19476 (N_19476,N_13156,N_12734);
or U19477 (N_19477,N_12113,N_14452);
nand U19478 (N_19478,N_12743,N_10779);
xor U19479 (N_19479,N_12455,N_13964);
or U19480 (N_19480,N_13158,N_12670);
and U19481 (N_19481,N_11671,N_12400);
nand U19482 (N_19482,N_11869,N_13557);
nor U19483 (N_19483,N_10764,N_10693);
xnor U19484 (N_19484,N_10106,N_13533);
nand U19485 (N_19485,N_14586,N_13594);
nand U19486 (N_19486,N_11139,N_11807);
xor U19487 (N_19487,N_13800,N_13374);
nand U19488 (N_19488,N_13110,N_11289);
nand U19489 (N_19489,N_10420,N_13687);
or U19490 (N_19490,N_12444,N_11743);
and U19491 (N_19491,N_13276,N_13831);
nand U19492 (N_19492,N_14891,N_14072);
nor U19493 (N_19493,N_12729,N_14073);
or U19494 (N_19494,N_14149,N_12487);
nand U19495 (N_19495,N_13592,N_10256);
or U19496 (N_19496,N_13354,N_11136);
or U19497 (N_19497,N_12407,N_10277);
and U19498 (N_19498,N_12565,N_13740);
nor U19499 (N_19499,N_11660,N_14404);
nand U19500 (N_19500,N_14143,N_11424);
and U19501 (N_19501,N_13320,N_13365);
and U19502 (N_19502,N_14050,N_10806);
and U19503 (N_19503,N_11001,N_13418);
nor U19504 (N_19504,N_10478,N_10261);
and U19505 (N_19505,N_14846,N_10424);
nand U19506 (N_19506,N_13652,N_12449);
nand U19507 (N_19507,N_14506,N_12772);
nor U19508 (N_19508,N_14658,N_14871);
xnor U19509 (N_19509,N_14382,N_11459);
nor U19510 (N_19510,N_10916,N_11123);
nand U19511 (N_19511,N_14753,N_14625);
nand U19512 (N_19512,N_14628,N_11001);
and U19513 (N_19513,N_14963,N_12298);
nor U19514 (N_19514,N_10030,N_12206);
or U19515 (N_19515,N_14459,N_11351);
and U19516 (N_19516,N_11314,N_13481);
and U19517 (N_19517,N_13741,N_13187);
nor U19518 (N_19518,N_13910,N_12800);
nor U19519 (N_19519,N_11458,N_12269);
and U19520 (N_19520,N_13671,N_13804);
and U19521 (N_19521,N_11749,N_13079);
nor U19522 (N_19522,N_10728,N_14332);
nand U19523 (N_19523,N_11104,N_11749);
nand U19524 (N_19524,N_11859,N_11324);
nor U19525 (N_19525,N_11060,N_13459);
or U19526 (N_19526,N_13032,N_14717);
and U19527 (N_19527,N_10456,N_13499);
nor U19528 (N_19528,N_12619,N_10097);
nand U19529 (N_19529,N_14098,N_11546);
nand U19530 (N_19530,N_10091,N_14001);
and U19531 (N_19531,N_14395,N_10409);
xor U19532 (N_19532,N_10488,N_14108);
xor U19533 (N_19533,N_13807,N_14485);
or U19534 (N_19534,N_10339,N_11912);
nor U19535 (N_19535,N_12884,N_12689);
xor U19536 (N_19536,N_13158,N_11890);
nand U19537 (N_19537,N_10402,N_12726);
nor U19538 (N_19538,N_12022,N_13275);
or U19539 (N_19539,N_12531,N_14240);
nand U19540 (N_19540,N_14234,N_10413);
xnor U19541 (N_19541,N_10155,N_14776);
or U19542 (N_19542,N_13443,N_10650);
or U19543 (N_19543,N_14781,N_13426);
nor U19544 (N_19544,N_14942,N_10514);
and U19545 (N_19545,N_10777,N_12621);
xnor U19546 (N_19546,N_12349,N_11051);
or U19547 (N_19547,N_14485,N_12838);
and U19548 (N_19548,N_10476,N_11373);
nor U19549 (N_19549,N_14355,N_14260);
xor U19550 (N_19550,N_10634,N_10999);
or U19551 (N_19551,N_13967,N_10551);
or U19552 (N_19552,N_12647,N_13600);
and U19553 (N_19553,N_12094,N_13833);
nand U19554 (N_19554,N_12504,N_12929);
or U19555 (N_19555,N_14064,N_10629);
xnor U19556 (N_19556,N_13032,N_10300);
xor U19557 (N_19557,N_10848,N_14842);
nand U19558 (N_19558,N_12287,N_14286);
nor U19559 (N_19559,N_13729,N_10315);
nor U19560 (N_19560,N_12557,N_13623);
nor U19561 (N_19561,N_12615,N_10119);
or U19562 (N_19562,N_13803,N_13290);
nand U19563 (N_19563,N_10253,N_12746);
nand U19564 (N_19564,N_10891,N_10383);
nor U19565 (N_19565,N_11901,N_12792);
and U19566 (N_19566,N_13644,N_11560);
nor U19567 (N_19567,N_13254,N_11367);
and U19568 (N_19568,N_14305,N_13191);
nand U19569 (N_19569,N_10094,N_10051);
and U19570 (N_19570,N_12135,N_11598);
xnor U19571 (N_19571,N_10442,N_12444);
and U19572 (N_19572,N_11680,N_13295);
or U19573 (N_19573,N_11647,N_11436);
nor U19574 (N_19574,N_10411,N_12314);
and U19575 (N_19575,N_11708,N_12304);
or U19576 (N_19576,N_13158,N_13031);
nor U19577 (N_19577,N_11886,N_11612);
or U19578 (N_19578,N_14824,N_14905);
nor U19579 (N_19579,N_14730,N_13535);
and U19580 (N_19580,N_12803,N_11292);
nand U19581 (N_19581,N_13232,N_10548);
nand U19582 (N_19582,N_13467,N_14897);
xnor U19583 (N_19583,N_14859,N_14986);
xnor U19584 (N_19584,N_11884,N_14774);
nor U19585 (N_19585,N_12629,N_11625);
nand U19586 (N_19586,N_12833,N_11900);
nand U19587 (N_19587,N_13105,N_14688);
or U19588 (N_19588,N_10338,N_12640);
nor U19589 (N_19589,N_14294,N_11347);
nand U19590 (N_19590,N_12593,N_11474);
nand U19591 (N_19591,N_10665,N_12814);
and U19592 (N_19592,N_13058,N_14394);
and U19593 (N_19593,N_14873,N_12242);
nor U19594 (N_19594,N_12051,N_10575);
xor U19595 (N_19595,N_11260,N_14753);
nand U19596 (N_19596,N_12499,N_14838);
and U19597 (N_19597,N_11665,N_11514);
nor U19598 (N_19598,N_14956,N_14980);
nor U19599 (N_19599,N_13375,N_10557);
or U19600 (N_19600,N_13705,N_10058);
and U19601 (N_19601,N_11201,N_10643);
or U19602 (N_19602,N_14410,N_10956);
and U19603 (N_19603,N_11231,N_13854);
nand U19604 (N_19604,N_13034,N_13757);
and U19605 (N_19605,N_13470,N_12972);
nand U19606 (N_19606,N_11305,N_12965);
nand U19607 (N_19607,N_12590,N_14742);
and U19608 (N_19608,N_14093,N_14230);
or U19609 (N_19609,N_13044,N_13296);
xor U19610 (N_19610,N_12360,N_11609);
and U19611 (N_19611,N_11852,N_12360);
or U19612 (N_19612,N_13246,N_11355);
nand U19613 (N_19613,N_13938,N_12836);
nand U19614 (N_19614,N_14781,N_13895);
nand U19615 (N_19615,N_10157,N_12576);
xor U19616 (N_19616,N_10289,N_10838);
or U19617 (N_19617,N_11052,N_13615);
and U19618 (N_19618,N_14152,N_10265);
nor U19619 (N_19619,N_13469,N_13981);
nand U19620 (N_19620,N_11470,N_13796);
or U19621 (N_19621,N_12788,N_13281);
or U19622 (N_19622,N_13976,N_14952);
nor U19623 (N_19623,N_11653,N_13300);
and U19624 (N_19624,N_12864,N_10737);
nor U19625 (N_19625,N_12713,N_12281);
and U19626 (N_19626,N_14925,N_14738);
or U19627 (N_19627,N_11052,N_10995);
nor U19628 (N_19628,N_14403,N_10923);
xnor U19629 (N_19629,N_13450,N_11767);
nor U19630 (N_19630,N_12323,N_14125);
xor U19631 (N_19631,N_10405,N_11195);
nor U19632 (N_19632,N_13577,N_13041);
or U19633 (N_19633,N_10318,N_14042);
or U19634 (N_19634,N_13394,N_13377);
nand U19635 (N_19635,N_12525,N_10911);
or U19636 (N_19636,N_12197,N_14107);
and U19637 (N_19637,N_10574,N_14984);
or U19638 (N_19638,N_11406,N_12952);
and U19639 (N_19639,N_11121,N_10833);
nor U19640 (N_19640,N_13166,N_11880);
nand U19641 (N_19641,N_11962,N_14496);
nor U19642 (N_19642,N_12862,N_13816);
nor U19643 (N_19643,N_10385,N_12569);
nor U19644 (N_19644,N_13132,N_12489);
nand U19645 (N_19645,N_11340,N_11467);
nor U19646 (N_19646,N_11257,N_12305);
or U19647 (N_19647,N_11096,N_11236);
and U19648 (N_19648,N_11297,N_12339);
nor U19649 (N_19649,N_13586,N_13203);
or U19650 (N_19650,N_10373,N_13067);
or U19651 (N_19651,N_11885,N_10845);
nand U19652 (N_19652,N_12548,N_14511);
or U19653 (N_19653,N_13141,N_12883);
nand U19654 (N_19654,N_10269,N_13591);
and U19655 (N_19655,N_13597,N_12947);
or U19656 (N_19656,N_14454,N_10474);
and U19657 (N_19657,N_12511,N_13819);
nor U19658 (N_19658,N_13765,N_14930);
nand U19659 (N_19659,N_13719,N_10574);
or U19660 (N_19660,N_13000,N_10639);
xnor U19661 (N_19661,N_11468,N_12196);
nand U19662 (N_19662,N_11901,N_13750);
or U19663 (N_19663,N_13780,N_12833);
nand U19664 (N_19664,N_13386,N_13545);
and U19665 (N_19665,N_13690,N_13232);
nor U19666 (N_19666,N_14235,N_11628);
or U19667 (N_19667,N_14325,N_11508);
or U19668 (N_19668,N_11240,N_11927);
nor U19669 (N_19669,N_10393,N_12353);
or U19670 (N_19670,N_14350,N_11501);
or U19671 (N_19671,N_11256,N_12491);
nand U19672 (N_19672,N_14432,N_14158);
or U19673 (N_19673,N_13863,N_12253);
nor U19674 (N_19674,N_13667,N_11311);
or U19675 (N_19675,N_11787,N_10850);
or U19676 (N_19676,N_11871,N_10834);
nor U19677 (N_19677,N_14003,N_13147);
or U19678 (N_19678,N_12026,N_11260);
or U19679 (N_19679,N_10293,N_14856);
nor U19680 (N_19680,N_12064,N_10603);
nor U19681 (N_19681,N_12262,N_11315);
nor U19682 (N_19682,N_13240,N_12090);
nor U19683 (N_19683,N_14211,N_14325);
nand U19684 (N_19684,N_12907,N_10523);
and U19685 (N_19685,N_14216,N_11897);
nor U19686 (N_19686,N_12250,N_14178);
or U19687 (N_19687,N_10237,N_11743);
nor U19688 (N_19688,N_14890,N_12175);
nand U19689 (N_19689,N_11688,N_14146);
or U19690 (N_19690,N_11368,N_14754);
xnor U19691 (N_19691,N_13203,N_14263);
xor U19692 (N_19692,N_10061,N_12441);
and U19693 (N_19693,N_13838,N_13255);
nand U19694 (N_19694,N_11937,N_11302);
nor U19695 (N_19695,N_13889,N_14976);
and U19696 (N_19696,N_10549,N_13680);
or U19697 (N_19697,N_11927,N_13078);
and U19698 (N_19698,N_12582,N_10395);
nor U19699 (N_19699,N_12854,N_10599);
or U19700 (N_19700,N_10415,N_12881);
nor U19701 (N_19701,N_13727,N_11404);
nand U19702 (N_19702,N_10154,N_11523);
or U19703 (N_19703,N_13403,N_13796);
or U19704 (N_19704,N_11653,N_10493);
nand U19705 (N_19705,N_14673,N_13892);
or U19706 (N_19706,N_11770,N_12308);
or U19707 (N_19707,N_11564,N_12262);
nor U19708 (N_19708,N_12386,N_14081);
nand U19709 (N_19709,N_10358,N_10561);
nor U19710 (N_19710,N_14801,N_11893);
nand U19711 (N_19711,N_12346,N_11390);
or U19712 (N_19712,N_12567,N_10062);
nand U19713 (N_19713,N_14938,N_12350);
or U19714 (N_19714,N_10943,N_14523);
nor U19715 (N_19715,N_11777,N_13529);
nand U19716 (N_19716,N_12994,N_13839);
and U19717 (N_19717,N_13858,N_12067);
nor U19718 (N_19718,N_13973,N_11031);
nand U19719 (N_19719,N_11095,N_13306);
and U19720 (N_19720,N_10830,N_12710);
and U19721 (N_19721,N_13811,N_11485);
and U19722 (N_19722,N_10805,N_13142);
and U19723 (N_19723,N_10172,N_14908);
and U19724 (N_19724,N_12897,N_10741);
nand U19725 (N_19725,N_12156,N_13905);
and U19726 (N_19726,N_11598,N_13691);
or U19727 (N_19727,N_13134,N_11619);
nor U19728 (N_19728,N_14172,N_11576);
nor U19729 (N_19729,N_11369,N_11238);
nor U19730 (N_19730,N_13011,N_10779);
or U19731 (N_19731,N_10475,N_10396);
nand U19732 (N_19732,N_14438,N_10357);
nand U19733 (N_19733,N_12785,N_13471);
nor U19734 (N_19734,N_14488,N_10016);
and U19735 (N_19735,N_14617,N_10800);
nand U19736 (N_19736,N_10267,N_13706);
xnor U19737 (N_19737,N_14760,N_13518);
nand U19738 (N_19738,N_14690,N_12812);
nor U19739 (N_19739,N_10828,N_14716);
and U19740 (N_19740,N_12307,N_12811);
nand U19741 (N_19741,N_10739,N_11493);
nand U19742 (N_19742,N_11244,N_13548);
nand U19743 (N_19743,N_11637,N_11240);
nand U19744 (N_19744,N_13969,N_14014);
or U19745 (N_19745,N_13056,N_14279);
nand U19746 (N_19746,N_10132,N_10353);
nand U19747 (N_19747,N_11026,N_11221);
nand U19748 (N_19748,N_10605,N_14223);
nand U19749 (N_19749,N_11064,N_11523);
nor U19750 (N_19750,N_14378,N_12553);
nand U19751 (N_19751,N_12096,N_12476);
nor U19752 (N_19752,N_14846,N_13817);
xor U19753 (N_19753,N_14820,N_10244);
and U19754 (N_19754,N_10221,N_13122);
or U19755 (N_19755,N_11299,N_11810);
nand U19756 (N_19756,N_14318,N_10797);
and U19757 (N_19757,N_14755,N_13893);
xnor U19758 (N_19758,N_12396,N_12866);
or U19759 (N_19759,N_10724,N_10494);
xor U19760 (N_19760,N_14782,N_13298);
xnor U19761 (N_19761,N_11525,N_11057);
or U19762 (N_19762,N_12575,N_11698);
nor U19763 (N_19763,N_10069,N_10517);
nand U19764 (N_19764,N_10212,N_14468);
nand U19765 (N_19765,N_12516,N_11998);
or U19766 (N_19766,N_13727,N_12913);
nand U19767 (N_19767,N_13633,N_10196);
nand U19768 (N_19768,N_12798,N_11079);
xnor U19769 (N_19769,N_12087,N_11183);
nor U19770 (N_19770,N_11993,N_14123);
xnor U19771 (N_19771,N_11992,N_14392);
nor U19772 (N_19772,N_14183,N_12957);
and U19773 (N_19773,N_12988,N_13286);
nand U19774 (N_19774,N_10795,N_10880);
nand U19775 (N_19775,N_12487,N_14908);
nand U19776 (N_19776,N_12112,N_10103);
and U19777 (N_19777,N_12175,N_14244);
nor U19778 (N_19778,N_13541,N_11949);
or U19779 (N_19779,N_12245,N_14541);
nand U19780 (N_19780,N_13417,N_11395);
or U19781 (N_19781,N_14831,N_12076);
and U19782 (N_19782,N_12522,N_13843);
and U19783 (N_19783,N_14938,N_13868);
and U19784 (N_19784,N_10440,N_11860);
nand U19785 (N_19785,N_10020,N_11292);
nand U19786 (N_19786,N_13089,N_10636);
and U19787 (N_19787,N_10261,N_11355);
nand U19788 (N_19788,N_14567,N_10051);
nor U19789 (N_19789,N_14417,N_14692);
nor U19790 (N_19790,N_10013,N_13827);
or U19791 (N_19791,N_12465,N_14531);
and U19792 (N_19792,N_11987,N_10680);
and U19793 (N_19793,N_11887,N_14739);
or U19794 (N_19794,N_10583,N_14736);
nand U19795 (N_19795,N_12674,N_11980);
and U19796 (N_19796,N_11490,N_13512);
or U19797 (N_19797,N_14372,N_14413);
and U19798 (N_19798,N_14891,N_10163);
nand U19799 (N_19799,N_11642,N_11512);
nand U19800 (N_19800,N_12335,N_12853);
and U19801 (N_19801,N_13294,N_14187);
and U19802 (N_19802,N_13563,N_10205);
nand U19803 (N_19803,N_11870,N_10672);
nor U19804 (N_19804,N_11677,N_10167);
or U19805 (N_19805,N_10886,N_11628);
or U19806 (N_19806,N_11212,N_12611);
or U19807 (N_19807,N_12335,N_14666);
xnor U19808 (N_19808,N_13072,N_12659);
nor U19809 (N_19809,N_13953,N_10833);
and U19810 (N_19810,N_11229,N_10018);
nor U19811 (N_19811,N_11672,N_10874);
and U19812 (N_19812,N_12903,N_14103);
nand U19813 (N_19813,N_14723,N_11692);
nor U19814 (N_19814,N_11865,N_10756);
xor U19815 (N_19815,N_14172,N_13159);
nand U19816 (N_19816,N_10621,N_13338);
xor U19817 (N_19817,N_11504,N_11668);
nor U19818 (N_19818,N_14880,N_12987);
xor U19819 (N_19819,N_11364,N_13816);
and U19820 (N_19820,N_14151,N_13745);
and U19821 (N_19821,N_12319,N_12442);
xnor U19822 (N_19822,N_11687,N_13293);
or U19823 (N_19823,N_12162,N_11385);
xor U19824 (N_19824,N_12680,N_12839);
or U19825 (N_19825,N_13628,N_10136);
and U19826 (N_19826,N_11730,N_12015);
or U19827 (N_19827,N_13022,N_10871);
and U19828 (N_19828,N_14313,N_10397);
nand U19829 (N_19829,N_14847,N_11860);
nor U19830 (N_19830,N_12299,N_13801);
and U19831 (N_19831,N_14629,N_13308);
xnor U19832 (N_19832,N_11195,N_10105);
and U19833 (N_19833,N_11623,N_11013);
xor U19834 (N_19834,N_10672,N_12131);
and U19835 (N_19835,N_14420,N_10969);
or U19836 (N_19836,N_12390,N_12926);
and U19837 (N_19837,N_12405,N_14580);
nand U19838 (N_19838,N_10223,N_13465);
nand U19839 (N_19839,N_12915,N_13800);
or U19840 (N_19840,N_13120,N_13974);
xnor U19841 (N_19841,N_12718,N_12540);
xnor U19842 (N_19842,N_11492,N_13978);
or U19843 (N_19843,N_10768,N_14077);
and U19844 (N_19844,N_10424,N_12308);
or U19845 (N_19845,N_12090,N_13484);
or U19846 (N_19846,N_14442,N_11293);
nand U19847 (N_19847,N_13718,N_13006);
and U19848 (N_19848,N_10767,N_11953);
xor U19849 (N_19849,N_13507,N_12123);
nand U19850 (N_19850,N_10080,N_10582);
xor U19851 (N_19851,N_14830,N_11742);
nor U19852 (N_19852,N_10985,N_14038);
nand U19853 (N_19853,N_14732,N_13975);
or U19854 (N_19854,N_12630,N_10122);
and U19855 (N_19855,N_14083,N_13052);
nand U19856 (N_19856,N_13665,N_14279);
or U19857 (N_19857,N_10138,N_14752);
nor U19858 (N_19858,N_12383,N_13011);
nor U19859 (N_19859,N_12543,N_14945);
or U19860 (N_19860,N_12638,N_13951);
nand U19861 (N_19861,N_11099,N_14887);
nand U19862 (N_19862,N_13153,N_13921);
nand U19863 (N_19863,N_12399,N_13425);
nor U19864 (N_19864,N_11757,N_13325);
nand U19865 (N_19865,N_10081,N_10923);
nor U19866 (N_19866,N_13214,N_11241);
and U19867 (N_19867,N_12348,N_12615);
nand U19868 (N_19868,N_12699,N_14553);
xor U19869 (N_19869,N_14183,N_10835);
xnor U19870 (N_19870,N_10885,N_10299);
xor U19871 (N_19871,N_10727,N_12413);
xnor U19872 (N_19872,N_12148,N_10596);
nor U19873 (N_19873,N_10430,N_14091);
xor U19874 (N_19874,N_11358,N_10189);
nor U19875 (N_19875,N_13145,N_14388);
and U19876 (N_19876,N_13214,N_12285);
nor U19877 (N_19877,N_12326,N_11546);
nor U19878 (N_19878,N_13276,N_12128);
nor U19879 (N_19879,N_14411,N_10040);
nor U19880 (N_19880,N_13111,N_11930);
nor U19881 (N_19881,N_11734,N_13927);
or U19882 (N_19882,N_11075,N_11414);
or U19883 (N_19883,N_14929,N_10192);
nor U19884 (N_19884,N_10390,N_14373);
nor U19885 (N_19885,N_11534,N_11526);
nor U19886 (N_19886,N_14689,N_10758);
nor U19887 (N_19887,N_11800,N_14260);
nand U19888 (N_19888,N_14577,N_14621);
nand U19889 (N_19889,N_13337,N_13528);
xor U19890 (N_19890,N_12595,N_10354);
nor U19891 (N_19891,N_13573,N_13948);
or U19892 (N_19892,N_14518,N_12736);
and U19893 (N_19893,N_10404,N_10488);
nand U19894 (N_19894,N_10587,N_12206);
nand U19895 (N_19895,N_11361,N_14750);
nor U19896 (N_19896,N_10153,N_12679);
nor U19897 (N_19897,N_10261,N_14962);
nand U19898 (N_19898,N_14748,N_14058);
xnor U19899 (N_19899,N_11436,N_11057);
and U19900 (N_19900,N_13131,N_13035);
and U19901 (N_19901,N_13903,N_11542);
nand U19902 (N_19902,N_13250,N_12073);
and U19903 (N_19903,N_11604,N_12463);
and U19904 (N_19904,N_12374,N_13994);
nor U19905 (N_19905,N_10774,N_12659);
and U19906 (N_19906,N_10651,N_12473);
and U19907 (N_19907,N_13549,N_13696);
or U19908 (N_19908,N_12231,N_11246);
or U19909 (N_19909,N_12687,N_13721);
and U19910 (N_19910,N_14780,N_12917);
nor U19911 (N_19911,N_11843,N_11747);
or U19912 (N_19912,N_10737,N_14732);
nand U19913 (N_19913,N_10277,N_12554);
nand U19914 (N_19914,N_10585,N_13512);
nor U19915 (N_19915,N_10699,N_12715);
and U19916 (N_19916,N_14147,N_12056);
nor U19917 (N_19917,N_11064,N_11642);
or U19918 (N_19918,N_14574,N_10242);
nor U19919 (N_19919,N_13498,N_11091);
and U19920 (N_19920,N_11116,N_10839);
and U19921 (N_19921,N_12348,N_13045);
nand U19922 (N_19922,N_12277,N_14207);
nand U19923 (N_19923,N_13455,N_13697);
nor U19924 (N_19924,N_10315,N_13810);
nand U19925 (N_19925,N_12913,N_14521);
nor U19926 (N_19926,N_10796,N_10268);
and U19927 (N_19927,N_10703,N_14259);
nor U19928 (N_19928,N_14980,N_14458);
nor U19929 (N_19929,N_14307,N_14232);
or U19930 (N_19930,N_13624,N_12753);
and U19931 (N_19931,N_10741,N_10121);
nand U19932 (N_19932,N_10926,N_11796);
and U19933 (N_19933,N_13357,N_12939);
or U19934 (N_19934,N_10627,N_14297);
or U19935 (N_19935,N_11982,N_14308);
nand U19936 (N_19936,N_10174,N_14175);
nand U19937 (N_19937,N_10872,N_10879);
or U19938 (N_19938,N_12921,N_11464);
nor U19939 (N_19939,N_11084,N_12337);
nand U19940 (N_19940,N_12866,N_11412);
and U19941 (N_19941,N_12811,N_10687);
and U19942 (N_19942,N_10062,N_12135);
nor U19943 (N_19943,N_11987,N_14982);
or U19944 (N_19944,N_13438,N_11298);
nand U19945 (N_19945,N_11423,N_13178);
xnor U19946 (N_19946,N_11507,N_12659);
nor U19947 (N_19947,N_11521,N_10797);
nand U19948 (N_19948,N_11578,N_12790);
xor U19949 (N_19949,N_10426,N_12656);
and U19950 (N_19950,N_11278,N_14000);
and U19951 (N_19951,N_12809,N_12626);
nand U19952 (N_19952,N_13258,N_12439);
nand U19953 (N_19953,N_11191,N_12282);
nand U19954 (N_19954,N_14910,N_11750);
xor U19955 (N_19955,N_12752,N_11058);
or U19956 (N_19956,N_14935,N_10685);
nand U19957 (N_19957,N_13255,N_12392);
xor U19958 (N_19958,N_10082,N_11275);
nand U19959 (N_19959,N_10835,N_14849);
nor U19960 (N_19960,N_14924,N_13291);
and U19961 (N_19961,N_11075,N_13850);
or U19962 (N_19962,N_14320,N_14601);
and U19963 (N_19963,N_13808,N_13420);
and U19964 (N_19964,N_13422,N_13105);
and U19965 (N_19965,N_14770,N_12397);
nor U19966 (N_19966,N_14433,N_11443);
or U19967 (N_19967,N_10501,N_13856);
xnor U19968 (N_19968,N_14690,N_14578);
nor U19969 (N_19969,N_13836,N_11158);
xor U19970 (N_19970,N_11446,N_14022);
and U19971 (N_19971,N_12875,N_11312);
nand U19972 (N_19972,N_12219,N_11716);
nor U19973 (N_19973,N_14115,N_11367);
nor U19974 (N_19974,N_11400,N_13260);
nor U19975 (N_19975,N_13493,N_10920);
nand U19976 (N_19976,N_13233,N_11085);
or U19977 (N_19977,N_11969,N_12360);
nor U19978 (N_19978,N_11085,N_12746);
or U19979 (N_19979,N_11076,N_11796);
and U19980 (N_19980,N_14712,N_12423);
nor U19981 (N_19981,N_14224,N_10537);
xor U19982 (N_19982,N_10431,N_10838);
nand U19983 (N_19983,N_10669,N_12533);
nor U19984 (N_19984,N_12672,N_13941);
or U19985 (N_19985,N_14441,N_14359);
nor U19986 (N_19986,N_10065,N_13682);
or U19987 (N_19987,N_10716,N_11838);
and U19988 (N_19988,N_10637,N_14209);
xor U19989 (N_19989,N_14610,N_13835);
xnor U19990 (N_19990,N_14286,N_11444);
and U19991 (N_19991,N_14771,N_10013);
xor U19992 (N_19992,N_14499,N_10112);
nor U19993 (N_19993,N_10442,N_11495);
xnor U19994 (N_19994,N_14748,N_14280);
nand U19995 (N_19995,N_13715,N_13567);
and U19996 (N_19996,N_14929,N_11608);
nand U19997 (N_19997,N_14794,N_10103);
nand U19998 (N_19998,N_11392,N_10509);
xnor U19999 (N_19999,N_10648,N_10083);
nor U20000 (N_20000,N_15516,N_19927);
nand U20001 (N_20001,N_15770,N_19326);
and U20002 (N_20002,N_17696,N_15286);
or U20003 (N_20003,N_16563,N_18445);
nor U20004 (N_20004,N_18258,N_16586);
and U20005 (N_20005,N_18244,N_19521);
nor U20006 (N_20006,N_15031,N_18307);
or U20007 (N_20007,N_17316,N_16114);
and U20008 (N_20008,N_18289,N_17545);
or U20009 (N_20009,N_16316,N_15760);
xor U20010 (N_20010,N_17768,N_17770);
and U20011 (N_20011,N_15141,N_19695);
or U20012 (N_20012,N_15102,N_18196);
or U20013 (N_20013,N_17810,N_17113);
nand U20014 (N_20014,N_17098,N_16060);
or U20015 (N_20015,N_19812,N_19188);
nand U20016 (N_20016,N_18771,N_15407);
nor U20017 (N_20017,N_15841,N_19191);
and U20018 (N_20018,N_18931,N_16098);
xor U20019 (N_20019,N_18456,N_18750);
nand U20020 (N_20020,N_16153,N_16438);
nand U20021 (N_20021,N_17443,N_17022);
or U20022 (N_20022,N_15625,N_18953);
nand U20023 (N_20023,N_17230,N_15877);
nor U20024 (N_20024,N_16923,N_17073);
and U20025 (N_20025,N_15854,N_16799);
nor U20026 (N_20026,N_19793,N_19732);
or U20027 (N_20027,N_15299,N_17792);
nand U20028 (N_20028,N_19496,N_18490);
or U20029 (N_20029,N_19803,N_16411);
nand U20030 (N_20030,N_15883,N_18123);
and U20031 (N_20031,N_19038,N_17755);
nor U20032 (N_20032,N_17589,N_15732);
nand U20033 (N_20033,N_17165,N_17763);
nor U20034 (N_20034,N_17556,N_15641);
or U20035 (N_20035,N_16392,N_15472);
nand U20036 (N_20036,N_17050,N_18969);
or U20037 (N_20037,N_15055,N_16310);
nand U20038 (N_20038,N_17520,N_16531);
and U20039 (N_20039,N_19725,N_19042);
nor U20040 (N_20040,N_15067,N_15795);
nor U20041 (N_20041,N_15367,N_17823);
and U20042 (N_20042,N_17775,N_18359);
nand U20043 (N_20043,N_17424,N_17732);
nor U20044 (N_20044,N_17415,N_15348);
nand U20045 (N_20045,N_18089,N_19456);
and U20046 (N_20046,N_16115,N_17963);
and U20047 (N_20047,N_16755,N_18113);
or U20048 (N_20048,N_15354,N_17650);
nor U20049 (N_20049,N_19097,N_18042);
xor U20050 (N_20050,N_16610,N_17568);
or U20051 (N_20051,N_15408,N_17661);
nand U20052 (N_20052,N_15405,N_16713);
nand U20053 (N_20053,N_16108,N_16277);
nand U20054 (N_20054,N_16720,N_16619);
nor U20055 (N_20055,N_15894,N_16100);
and U20056 (N_20056,N_15713,N_15862);
and U20057 (N_20057,N_15647,N_17538);
nor U20058 (N_20058,N_15529,N_15123);
nand U20059 (N_20059,N_19316,N_18919);
or U20060 (N_20060,N_18486,N_15960);
and U20061 (N_20061,N_18461,N_17607);
and U20062 (N_20062,N_18728,N_19482);
or U20063 (N_20063,N_15621,N_15062);
or U20064 (N_20064,N_17311,N_16585);
xor U20065 (N_20065,N_15683,N_16640);
nor U20066 (N_20066,N_18471,N_19970);
nand U20067 (N_20067,N_17234,N_17903);
and U20068 (N_20068,N_19043,N_16184);
nand U20069 (N_20069,N_16395,N_17937);
xnor U20070 (N_20070,N_15701,N_17644);
and U20071 (N_20071,N_16746,N_17675);
nor U20072 (N_20072,N_17727,N_15169);
nand U20073 (N_20073,N_18335,N_18309);
nand U20074 (N_20074,N_18477,N_15613);
nand U20075 (N_20075,N_17793,N_18663);
nand U20076 (N_20076,N_15742,N_19268);
nand U20077 (N_20077,N_18357,N_15043);
nor U20078 (N_20078,N_19088,N_18971);
nor U20079 (N_20079,N_16293,N_16848);
and U20080 (N_20080,N_18773,N_18339);
and U20081 (N_20081,N_18669,N_15993);
and U20082 (N_20082,N_16227,N_17319);
xor U20083 (N_20083,N_18873,N_16988);
or U20084 (N_20084,N_15487,N_19397);
nand U20085 (N_20085,N_18866,N_17587);
nand U20086 (N_20086,N_17566,N_15360);
nand U20087 (N_20087,N_16786,N_15921);
nor U20088 (N_20088,N_17984,N_16462);
xnor U20089 (N_20089,N_17645,N_19443);
nor U20090 (N_20090,N_16377,N_17345);
xnor U20091 (N_20091,N_17181,N_17851);
or U20092 (N_20092,N_15422,N_15934);
or U20093 (N_20093,N_17772,N_18774);
or U20094 (N_20094,N_15281,N_18909);
xor U20095 (N_20095,N_16119,N_19834);
nand U20096 (N_20096,N_17571,N_19801);
nand U20097 (N_20097,N_16929,N_18813);
nand U20098 (N_20098,N_16215,N_18480);
and U20099 (N_20099,N_17553,N_15924);
or U20100 (N_20100,N_19848,N_19862);
nor U20101 (N_20101,N_17454,N_18615);
xnor U20102 (N_20102,N_17299,N_19486);
and U20103 (N_20103,N_18579,N_18758);
nor U20104 (N_20104,N_15144,N_16291);
and U20105 (N_20105,N_18393,N_15998);
and U20106 (N_20106,N_17972,N_15090);
nor U20107 (N_20107,N_17132,N_18641);
nand U20108 (N_20108,N_17776,N_19063);
nor U20109 (N_20109,N_18632,N_19284);
or U20110 (N_20110,N_19515,N_16123);
nor U20111 (N_20111,N_19250,N_18635);
and U20112 (N_20112,N_18325,N_17122);
and U20113 (N_20113,N_15492,N_15978);
and U20114 (N_20114,N_15497,N_15117);
and U20115 (N_20115,N_18047,N_16703);
nand U20116 (N_20116,N_18648,N_19671);
or U20117 (N_20117,N_15328,N_18779);
nand U20118 (N_20118,N_15139,N_17346);
nor U20119 (N_20119,N_17537,N_17910);
nor U20120 (N_20120,N_16389,N_18129);
nand U20121 (N_20121,N_17583,N_15650);
nand U20122 (N_20122,N_19347,N_16606);
or U20123 (N_20123,N_16443,N_15997);
or U20124 (N_20124,N_18831,N_17381);
or U20125 (N_20125,N_19401,N_15815);
nor U20126 (N_20126,N_16984,N_19736);
nand U20127 (N_20127,N_19608,N_17142);
or U20128 (N_20128,N_19594,N_15464);
and U20129 (N_20129,N_16396,N_18204);
nor U20130 (N_20130,N_15046,N_17664);
or U20131 (N_20131,N_15489,N_19052);
nand U20132 (N_20132,N_15794,N_15570);
nor U20133 (N_20133,N_15015,N_18988);
or U20134 (N_20134,N_15989,N_15975);
or U20135 (N_20135,N_19086,N_17210);
and U20136 (N_20136,N_16430,N_18961);
nand U20137 (N_20137,N_15509,N_17617);
and U20138 (N_20138,N_16325,N_16244);
nor U20139 (N_20139,N_17154,N_15298);
nor U20140 (N_20140,N_17268,N_16276);
nor U20141 (N_20141,N_17161,N_16948);
nor U20142 (N_20142,N_19916,N_15513);
nand U20143 (N_20143,N_15659,N_18535);
or U20144 (N_20144,N_15908,N_18804);
nand U20145 (N_20145,N_18941,N_18793);
or U20146 (N_20146,N_15124,N_17517);
nor U20147 (N_20147,N_18299,N_19035);
or U20148 (N_20148,N_16584,N_16925);
nor U20149 (N_20149,N_18139,N_16722);
nor U20150 (N_20150,N_16340,N_19391);
or U20151 (N_20151,N_18220,N_18508);
or U20152 (N_20152,N_19956,N_16598);
nand U20153 (N_20153,N_15684,N_18029);
or U20154 (N_20154,N_18968,N_18468);
nand U20155 (N_20155,N_16361,N_16618);
nor U20156 (N_20156,N_15536,N_16605);
nand U20157 (N_20157,N_19190,N_19855);
nor U20158 (N_20158,N_17817,N_16057);
and U20159 (N_20159,N_17205,N_16111);
or U20160 (N_20160,N_19788,N_19737);
nor U20161 (N_20161,N_15609,N_17215);
or U20162 (N_20162,N_15679,N_16835);
nand U20163 (N_20163,N_15576,N_19882);
nor U20164 (N_20164,N_16674,N_19340);
or U20165 (N_20165,N_15091,N_15358);
and U20166 (N_20166,N_17925,N_18956);
and U20167 (N_20167,N_15832,N_18489);
or U20168 (N_20168,N_18180,N_16024);
nor U20169 (N_20169,N_15869,N_15192);
and U20170 (N_20170,N_17484,N_16953);
nand U20171 (N_20171,N_16157,N_15109);
nand U20172 (N_20172,N_18562,N_15018);
nor U20173 (N_20173,N_15138,N_17973);
nor U20174 (N_20174,N_16936,N_15230);
nor U20175 (N_20175,N_16199,N_18484);
xnor U20176 (N_20176,N_15959,N_17873);
nor U20177 (N_20177,N_16066,N_19615);
nand U20178 (N_20178,N_17799,N_17407);
nor U20179 (N_20179,N_18483,N_19321);
or U20180 (N_20180,N_16302,N_16512);
xor U20181 (N_20181,N_16313,N_18937);
nand U20182 (N_20182,N_16080,N_15653);
nand U20183 (N_20183,N_16572,N_15001);
and U20184 (N_20184,N_18858,N_15886);
and U20185 (N_20185,N_18405,N_16678);
nor U20186 (N_20186,N_15700,N_15936);
or U20187 (N_20187,N_18412,N_19392);
nand U20188 (N_20188,N_18210,N_17889);
nor U20189 (N_20189,N_16632,N_18832);
and U20190 (N_20190,N_15637,N_18198);
and U20191 (N_20191,N_18580,N_16287);
or U20192 (N_20192,N_18695,N_15630);
xnor U20193 (N_20193,N_16207,N_19505);
or U20194 (N_20194,N_19081,N_15481);
or U20195 (N_20195,N_15948,N_16007);
nor U20196 (N_20196,N_19181,N_15041);
nand U20197 (N_20197,N_15480,N_19135);
and U20198 (N_20198,N_19382,N_17141);
and U20199 (N_20199,N_15498,N_19602);
nor U20200 (N_20200,N_16882,N_15147);
and U20201 (N_20201,N_15871,N_19715);
nor U20202 (N_20202,N_19674,N_18946);
or U20203 (N_20203,N_16687,N_19637);
nand U20204 (N_20204,N_19257,N_18955);
and U20205 (N_20205,N_17325,N_16910);
nand U20206 (N_20206,N_17597,N_16570);
or U20207 (N_20207,N_17365,N_17290);
and U20208 (N_20208,N_16349,N_17550);
or U20209 (N_20209,N_18698,N_16914);
and U20210 (N_20210,N_17264,N_18286);
xor U20211 (N_20211,N_16763,N_15163);
nor U20212 (N_20212,N_19807,N_17363);
or U20213 (N_20213,N_19977,N_18678);
nor U20214 (N_20214,N_17331,N_18559);
or U20215 (N_20215,N_18578,N_19403);
nand U20216 (N_20216,N_18671,N_19682);
nor U20217 (N_20217,N_15380,N_15897);
and U20218 (N_20218,N_18842,N_18326);
nor U20219 (N_20219,N_18132,N_19380);
and U20220 (N_20220,N_17766,N_18703);
nor U20221 (N_20221,N_17606,N_19213);
or U20222 (N_20222,N_19600,N_19858);
or U20223 (N_20223,N_17803,N_15825);
and U20224 (N_20224,N_16523,N_16874);
and U20225 (N_20225,N_15939,N_16224);
and U20226 (N_20226,N_17241,N_16436);
nand U20227 (N_20227,N_16802,N_19867);
nor U20228 (N_20228,N_15443,N_18538);
nand U20229 (N_20229,N_19751,N_18320);
nand U20230 (N_20230,N_18592,N_16771);
nand U20231 (N_20231,N_17988,N_18117);
nor U20232 (N_20232,N_19362,N_19293);
nand U20233 (N_20233,N_15577,N_15632);
nor U20234 (N_20234,N_19827,N_18531);
and U20235 (N_20235,N_17704,N_17414);
nand U20236 (N_20236,N_16429,N_15820);
or U20237 (N_20237,N_18203,N_17460);
or U20238 (N_20238,N_15127,N_15451);
nor U20239 (N_20239,N_16871,N_15342);
xnor U20240 (N_20240,N_17229,N_18500);
nand U20241 (N_20241,N_19123,N_18548);
and U20242 (N_20242,N_17062,N_16762);
and U20243 (N_20243,N_19092,N_16453);
and U20244 (N_20244,N_17099,N_16614);
and U20245 (N_20245,N_18388,N_17398);
nor U20246 (N_20246,N_15896,N_19149);
nand U20247 (N_20247,N_17863,N_15734);
or U20248 (N_20248,N_18452,N_17413);
xor U20249 (N_20249,N_18190,N_16040);
nand U20250 (N_20250,N_17052,N_18653);
xnor U20251 (N_20251,N_15793,N_17006);
xor U20252 (N_20252,N_16753,N_15827);
and U20253 (N_20253,N_16769,N_19694);
nor U20254 (N_20254,N_18834,N_17506);
nor U20255 (N_20255,N_15769,N_19872);
and U20256 (N_20256,N_15395,N_19624);
or U20257 (N_20257,N_19356,N_15914);
nand U20258 (N_20258,N_18084,N_15245);
nor U20259 (N_20259,N_15932,N_16768);
nand U20260 (N_20260,N_17942,N_19783);
xor U20261 (N_20261,N_16124,N_19782);
and U20262 (N_20262,N_15465,N_16707);
or U20263 (N_20263,N_17138,N_19084);
and U20264 (N_20264,N_16928,N_18802);
xnor U20265 (N_20265,N_16342,N_17720);
or U20266 (N_20266,N_19606,N_16601);
nand U20267 (N_20267,N_18905,N_15375);
nand U20268 (N_20268,N_18686,N_19335);
nor U20269 (N_20269,N_18867,N_18354);
and U20270 (N_20270,N_18826,N_16509);
or U20271 (N_20271,N_16859,N_18100);
or U20272 (N_20272,N_16938,N_15208);
or U20273 (N_20273,N_19417,N_19534);
nor U20274 (N_20274,N_17324,N_18718);
xnor U20275 (N_20275,N_16073,N_18967);
nor U20276 (N_20276,N_15437,N_18853);
nand U20277 (N_20277,N_19444,N_16685);
or U20278 (N_20278,N_19398,N_15910);
xnor U20279 (N_20279,N_16812,N_19144);
nand U20280 (N_20280,N_16943,N_17983);
or U20281 (N_20281,N_18680,N_17246);
nor U20282 (N_20282,N_19079,N_18994);
nand U20283 (N_20283,N_17193,N_16797);
and U20284 (N_20284,N_17280,N_15445);
nand U20285 (N_20285,N_15050,N_16472);
xnor U20286 (N_20286,N_16783,N_18249);
xnor U20287 (N_20287,N_17690,N_15634);
and U20288 (N_20288,N_19234,N_18332);
or U20289 (N_20289,N_18021,N_18202);
nor U20290 (N_20290,N_15707,N_17480);
xnor U20291 (N_20291,N_17105,N_16271);
nor U20292 (N_20292,N_18261,N_19050);
xor U20293 (N_20293,N_17883,N_18920);
and U20294 (N_20294,N_18275,N_17818);
or U20295 (N_20295,N_17080,N_15218);
or U20296 (N_20296,N_15204,N_18000);
nor U20297 (N_20297,N_18897,N_19543);
and U20298 (N_20298,N_15926,N_17308);
xnor U20299 (N_20299,N_16037,N_18270);
xnor U20300 (N_20300,N_18135,N_16103);
xnor U20301 (N_20301,N_15024,N_15476);
nand U20302 (N_20302,N_15963,N_15675);
and U20303 (N_20303,N_16908,N_18554);
nor U20304 (N_20304,N_17565,N_19044);
nand U20305 (N_20305,N_17301,N_17372);
or U20306 (N_20306,N_16044,N_19612);
and U20307 (N_20307,N_18241,N_15452);
and U20308 (N_20308,N_19108,N_17716);
nor U20309 (N_20309,N_15656,N_19780);
nor U20310 (N_20310,N_18928,N_17089);
nor U20311 (N_20311,N_18612,N_15321);
xor U20312 (N_20312,N_18990,N_19607);
or U20313 (N_20313,N_17876,N_18972);
and U20314 (N_20314,N_18345,N_19893);
or U20315 (N_20315,N_16331,N_16475);
and U20316 (N_20316,N_19437,N_19984);
nand U20317 (N_20317,N_16324,N_19013);
or U20318 (N_20318,N_17379,N_15237);
nand U20319 (N_20319,N_19911,N_15211);
and U20320 (N_20320,N_19476,N_17788);
or U20321 (N_20321,N_19436,N_18526);
nand U20322 (N_20322,N_16960,N_16834);
nand U20323 (N_20323,N_15273,N_19932);
xnor U20324 (N_20324,N_15602,N_15330);
xnor U20325 (N_20325,N_18647,N_15457);
or U20326 (N_20326,N_18308,N_17496);
or U20327 (N_20327,N_18255,N_18948);
and U20328 (N_20328,N_17189,N_15122);
xnor U20329 (N_20329,N_19313,N_16308);
xnor U20330 (N_20330,N_19021,N_19442);
and U20331 (N_20331,N_17457,N_17387);
nor U20332 (N_20332,N_17592,N_18626);
or U20333 (N_20333,N_16643,N_19345);
nor U20334 (N_20334,N_15698,N_18193);
nand U20335 (N_20335,N_17338,N_16195);
nor U20336 (N_20336,N_17020,N_17169);
or U20337 (N_20337,N_18938,N_19734);
nor U20338 (N_20338,N_16046,N_15682);
nand U20339 (N_20339,N_18589,N_19163);
nand U20340 (N_20340,N_16867,N_16997);
nor U20341 (N_20341,N_15677,N_19256);
and U20342 (N_20342,N_17834,N_15530);
nor U20343 (N_20343,N_16315,N_19950);
and U20344 (N_20344,N_18627,N_18583);
nand U20345 (N_20345,N_16375,N_15765);
nand U20346 (N_20346,N_16552,N_17312);
nor U20347 (N_20347,N_19273,N_15391);
or U20348 (N_20348,N_16930,N_16937);
and U20349 (N_20349,N_18852,N_17194);
and U20350 (N_20350,N_17527,N_16043);
and U20351 (N_20351,N_19167,N_19018);
and U20352 (N_20352,N_17039,N_16652);
nand U20353 (N_20353,N_18045,N_17015);
nand U20354 (N_20354,N_18374,N_19469);
xor U20355 (N_20355,N_16228,N_16955);
nor U20356 (N_20356,N_15154,N_15885);
xor U20357 (N_20357,N_16580,N_18720);
nor U20358 (N_20358,N_18701,N_18199);
nor U20359 (N_20359,N_16174,N_15935);
nor U20360 (N_20360,N_16992,N_15243);
nor U20361 (N_20361,N_15544,N_19104);
and U20362 (N_20362,N_15011,N_18808);
and U20363 (N_20363,N_16476,N_17888);
nand U20364 (N_20364,N_17995,N_17913);
nand U20365 (N_20365,N_19001,N_18913);
nand U20366 (N_20366,N_18574,N_19151);
or U20367 (N_20367,N_16279,N_17235);
nor U20368 (N_20368,N_18890,N_18982);
nor U20369 (N_20369,N_18713,N_15275);
or U20370 (N_20370,N_18654,N_19756);
nor U20371 (N_20371,N_17103,N_19841);
xnor U20372 (N_20372,N_17977,N_18534);
or U20373 (N_20373,N_17116,N_19741);
or U20374 (N_20374,N_19499,N_16017);
nand U20375 (N_20375,N_15241,N_18068);
and U20376 (N_20376,N_15953,N_19519);
or U20377 (N_20377,N_16106,N_19118);
nand U20378 (N_20378,N_17542,N_17611);
or U20379 (N_20379,N_18581,N_16983);
or U20380 (N_20380,N_17263,N_15103);
nand U20381 (N_20381,N_17777,N_15733);
and U20382 (N_20382,N_19473,N_17481);
or U20383 (N_20383,N_18302,N_16965);
nor U20384 (N_20384,N_17501,N_16417);
and U20385 (N_20385,N_19955,N_18874);
nor U20386 (N_20386,N_17886,N_17633);
and U20387 (N_20387,N_18106,N_19635);
or U20388 (N_20388,N_16508,N_15221);
nor U20389 (N_20389,N_15143,N_15327);
nor U20390 (N_20390,N_18185,N_17027);
or U20391 (N_20391,N_16716,N_18227);
xnor U20392 (N_20392,N_15592,N_15938);
nor U20393 (N_20393,N_17557,N_15767);
nor U20394 (N_20394,N_17710,N_15357);
and U20395 (N_20395,N_16084,N_17723);
and U20396 (N_20396,N_17416,N_17797);
nor U20397 (N_20397,N_18290,N_19604);
nand U20398 (N_20398,N_16721,N_16470);
xor U20399 (N_20399,N_15730,N_15416);
or U20400 (N_20400,N_15288,N_15586);
nand U20401 (N_20401,N_15119,N_19937);
nor U20402 (N_20402,N_18830,N_19998);
nor U20403 (N_20403,N_18136,N_15362);
or U20404 (N_20404,N_15979,N_19661);
or U20405 (N_20405,N_19148,N_19236);
xnor U20406 (N_20406,N_19419,N_15388);
and U20407 (N_20407,N_18823,N_16596);
nor U20408 (N_20408,N_15461,N_19838);
and U20409 (N_20409,N_17184,N_19854);
nand U20410 (N_20410,N_17249,N_15180);
or U20411 (N_20411,N_15879,N_16104);
nand U20412 (N_20412,N_17326,N_17750);
and U20413 (N_20413,N_17865,N_17148);
nand U20414 (N_20414,N_18514,N_17003);
nand U20415 (N_20415,N_15748,N_18043);
or U20416 (N_20416,N_18169,N_19287);
nand U20417 (N_20417,N_18032,N_18291);
nor U20418 (N_20418,N_17804,N_16458);
and U20419 (N_20419,N_15142,N_19590);
nand U20420 (N_20420,N_18434,N_18670);
and U20421 (N_20421,N_16649,N_16645);
and U20422 (N_20422,N_18310,N_19928);
or U20423 (N_20423,N_15235,N_19174);
or U20424 (N_20424,N_19690,N_17436);
or U20425 (N_20425,N_17997,N_19155);
and U20426 (N_20426,N_16258,N_18191);
or U20427 (N_20427,N_16588,N_16365);
nor U20428 (N_20428,N_15115,N_15397);
and U20429 (N_20429,N_18503,N_19040);
or U20430 (N_20430,N_19240,N_19225);
xor U20431 (N_20431,N_16845,N_18298);
nand U20432 (N_20432,N_18437,N_17315);
nor U20433 (N_20433,N_15696,N_19219);
nor U20434 (N_20434,N_15284,N_17602);
xnor U20435 (N_20435,N_15239,N_16934);
xor U20436 (N_20436,N_17030,N_19926);
nand U20437 (N_20437,N_16789,N_16319);
and U20438 (N_20438,N_16558,N_15655);
nand U20439 (N_20439,N_15216,N_19945);
nand U20440 (N_20440,N_19016,N_19312);
nand U20441 (N_20441,N_16127,N_15839);
or U20442 (N_20442,N_17614,N_18166);
nand U20443 (N_20443,N_19987,N_18116);
xor U20444 (N_20444,N_19860,N_17608);
nor U20445 (N_20445,N_16735,N_17117);
nor U20446 (N_20446,N_19479,N_16055);
and U20447 (N_20447,N_15073,N_16742);
or U20448 (N_20448,N_18597,N_16190);
nand U20449 (N_20449,N_19076,N_16001);
and U20450 (N_20450,N_19399,N_18271);
and U20451 (N_20451,N_18152,N_19260);
nor U20452 (N_20452,N_15468,N_17441);
and U20453 (N_20453,N_15944,N_16577);
or U20454 (N_20454,N_17064,N_17752);
or U20455 (N_20455,N_19210,N_19561);
and U20456 (N_20456,N_17479,N_16163);
nor U20457 (N_20457,N_18367,N_16469);
nand U20458 (N_20458,N_17273,N_16092);
nand U20459 (N_20459,N_15807,N_15096);
nand U20460 (N_20460,N_18738,N_15022);
or U20461 (N_20461,N_17699,N_19408);
or U20462 (N_20462,N_17172,N_19787);
or U20463 (N_20463,N_16749,N_17310);
nor U20464 (N_20464,N_18195,N_16917);
nand U20465 (N_20465,N_17366,N_17289);
nand U20466 (N_20466,N_17670,N_16274);
and U20467 (N_20467,N_19105,N_18712);
nor U20468 (N_20468,N_16264,N_16972);
nor U20469 (N_20469,N_19610,N_17756);
nor U20470 (N_20470,N_17483,N_18101);
nand U20471 (N_20471,N_18649,N_17652);
or U20472 (N_20472,N_15202,N_16376);
nand U20473 (N_20473,N_19949,N_17475);
nor U20474 (N_20474,N_18745,N_16465);
or U20475 (N_20475,N_18296,N_19343);
nor U20476 (N_20476,N_15318,N_16814);
or U20477 (N_20477,N_15300,N_18109);
nor U20478 (N_20478,N_19556,N_16857);
or U20479 (N_20479,N_16765,N_16906);
nor U20480 (N_20480,N_19462,N_19102);
nand U20481 (N_20481,N_16574,N_19548);
and U20482 (N_20482,N_15365,N_15850);
nand U20483 (N_20483,N_18172,N_19957);
or U20484 (N_20484,N_17114,N_19007);
or U20485 (N_20485,N_16963,N_19625);
and U20486 (N_20486,N_16909,N_16010);
or U20487 (N_20487,N_17966,N_19520);
nand U20488 (N_20488,N_15726,N_15227);
and U20489 (N_20489,N_19322,N_19455);
nand U20490 (N_20490,N_18668,N_19699);
nor U20491 (N_20491,N_18079,N_18533);
nand U20492 (N_20492,N_16201,N_19816);
nor U20493 (N_20493,N_16604,N_17223);
xor U20494 (N_20494,N_18173,N_19433);
or U20495 (N_20495,N_19415,N_15899);
xor U20496 (N_20496,N_18426,N_17048);
or U20497 (N_20497,N_18086,N_18833);
and U20498 (N_20498,N_18283,N_15833);
nor U20499 (N_20499,N_17385,N_16144);
nor U20500 (N_20500,N_16382,N_17397);
xnor U20501 (N_20501,N_15167,N_18383);
nor U20502 (N_20502,N_17642,N_19253);
nor U20503 (N_20503,N_17771,N_17708);
nand U20504 (N_20504,N_19239,N_17247);
or U20505 (N_20505,N_17250,N_17662);
and U20506 (N_20506,N_19306,N_15652);
nand U20507 (N_20507,N_19175,N_17049);
and U20508 (N_20508,N_18385,N_16218);
or U20509 (N_20509,N_15013,N_15704);
nor U20510 (N_20510,N_19824,N_15101);
xnor U20511 (N_20511,N_18229,N_15515);
nand U20512 (N_20512,N_19330,N_19572);
nor U20513 (N_20513,N_18070,N_19172);
nor U20514 (N_20514,N_19169,N_19748);
xor U20515 (N_20515,N_18506,N_19967);
nor U20516 (N_20516,N_15152,N_19506);
or U20517 (N_20517,N_15310,N_18104);
and U20518 (N_20518,N_18273,N_19669);
or U20519 (N_20519,N_19117,N_17898);
and U20520 (N_20520,N_16180,N_16792);
or U20521 (N_20521,N_15836,N_18693);
nand U20522 (N_20522,N_15785,N_17643);
nor U20523 (N_20523,N_18333,N_19651);
or U20524 (N_20524,N_17200,N_16099);
nor U20525 (N_20525,N_18545,N_18756);
and U20526 (N_20526,N_18734,N_17097);
nor U20527 (N_20527,N_15149,N_15116);
nand U20528 (N_20528,N_19712,N_16636);
nand U20529 (N_20529,N_16288,N_19541);
or U20530 (N_20530,N_16367,N_15941);
and U20531 (N_20531,N_18467,N_16327);
nor U20532 (N_20532,N_16975,N_19186);
and U20533 (N_20533,N_19184,N_16179);
nor U20534 (N_20534,N_15340,N_19898);
nand U20535 (N_20535,N_16050,N_19342);
or U20536 (N_20536,N_16656,N_15458);
or U20537 (N_20537,N_17962,N_15957);
and U20538 (N_20538,N_19871,N_17463);
nand U20539 (N_20539,N_17322,N_15068);
and U20540 (N_20540,N_18430,N_18942);
nor U20541 (N_20541,N_16782,N_19598);
and U20542 (N_20542,N_16303,N_17427);
and U20543 (N_20543,N_16217,N_18392);
or U20544 (N_20544,N_17522,N_19261);
and U20545 (N_20545,N_19731,N_15880);
or U20546 (N_20546,N_18504,N_15681);
and U20547 (N_20547,N_15564,N_18857);
and U20548 (N_20548,N_17769,N_17778);
nand U20549 (N_20549,N_17007,N_18519);
nand U20550 (N_20550,N_19776,N_18369);
and U20551 (N_20551,N_16504,N_16736);
nand U20552 (N_20552,N_15986,N_18167);
xnor U20553 (N_20553,N_18362,N_15561);
nor U20554 (N_20554,N_15629,N_17576);
nand U20555 (N_20555,N_18851,N_19297);
or U20556 (N_20556,N_16404,N_19822);
or U20557 (N_20557,N_15864,N_16881);
nor U20558 (N_20558,N_18730,N_16322);
xnor U20559 (N_20559,N_17647,N_19899);
xnor U20560 (N_20560,N_19564,N_19070);
nand U20561 (N_20561,N_18366,N_16280);
xnor U20562 (N_20562,N_19028,N_16565);
and U20563 (N_20563,N_15719,N_19868);
nand U20564 (N_20564,N_15473,N_17258);
nand U20565 (N_20565,N_18697,N_18398);
xnor U20566 (N_20566,N_15949,N_15995);
or U20567 (N_20567,N_17076,N_18634);
nand U20568 (N_20568,N_19930,N_17878);
nand U20569 (N_20569,N_15738,N_17107);
and U20570 (N_20570,N_19095,N_17430);
nor U20571 (N_20571,N_17836,N_17164);
and U20572 (N_20572,N_18930,N_17618);
or U20573 (N_20573,N_19923,N_16880);
nand U20574 (N_20574,N_15690,N_18660);
and U20575 (N_20575,N_15410,N_17761);
or U20576 (N_20576,N_17058,N_19537);
or U20577 (N_20577,N_18066,N_16440);
nor U20578 (N_20578,N_19048,N_17564);
or U20579 (N_20579,N_17108,N_16418);
or U20580 (N_20580,N_18895,N_16204);
nand U20581 (N_20581,N_19468,N_18762);
and U20582 (N_20582,N_17866,N_16499);
or U20583 (N_20583,N_15840,N_18814);
and U20584 (N_20584,N_17897,N_18093);
and U20585 (N_20585,N_19022,N_18420);
xnor U20586 (N_20586,N_19423,N_19791);
nand U20587 (N_20587,N_17738,N_17620);
and U20588 (N_20588,N_19536,N_15565);
nor U20589 (N_20589,N_16571,N_19067);
and U20590 (N_20590,N_19672,N_16833);
nor U20591 (N_20591,N_17271,N_16919);
or U20592 (N_20592,N_19634,N_16849);
nor U20593 (N_20593,N_16830,N_15373);
nor U20594 (N_20594,N_18102,N_18751);
nor U20595 (N_20595,N_18633,N_19975);
nor U20596 (N_20596,N_18124,N_16011);
or U20597 (N_20597,N_16904,N_16268);
nand U20598 (N_20598,N_19494,N_17505);
and U20599 (N_20599,N_16081,N_17439);
xnor U20600 (N_20600,N_18485,N_18735);
and U20601 (N_20601,N_17425,N_15579);
nor U20602 (N_20602,N_18729,N_15070);
nand U20603 (N_20603,N_17531,N_16415);
nor U20604 (N_20604,N_18950,N_16048);
nor U20605 (N_20605,N_18957,N_19716);
or U20606 (N_20606,N_18617,N_18372);
and U20607 (N_20607,N_19605,N_19470);
nor U20608 (N_20608,N_15114,N_16872);
nand U20609 (N_20609,N_16727,N_15988);
and U20610 (N_20610,N_19831,N_19996);
nor U20611 (N_20611,N_15984,N_19371);
or U20612 (N_20612,N_18860,N_18845);
nand U20613 (N_20613,N_17202,N_15210);
nand U20614 (N_20614,N_19243,N_17159);
or U20615 (N_20615,N_16068,N_19394);
or U20616 (N_20616,N_15242,N_18665);
nand U20617 (N_20617,N_19890,N_16478);
or U20618 (N_20618,N_15170,N_17368);
xnor U20619 (N_20619,N_19232,N_15254);
and U20620 (N_20620,N_18294,N_17572);
nor U20621 (N_20621,N_18546,N_15185);
nand U20622 (N_20622,N_17852,N_17954);
nor U20623 (N_20623,N_17621,N_18599);
xor U20624 (N_20624,N_15507,N_16850);
and U20625 (N_20625,N_15574,N_16189);
nand U20626 (N_20626,N_15039,N_15135);
or U20627 (N_20627,N_17570,N_19739);
nand U20628 (N_20628,N_15818,N_19222);
nand U20629 (N_20629,N_18947,N_19457);
or U20630 (N_20630,N_19015,N_15444);
and U20631 (N_20631,N_16594,N_16134);
xnor U20632 (N_20632,N_18246,N_18555);
and U20633 (N_20633,N_15728,N_17872);
or U20634 (N_20634,N_16852,N_19000);
xnor U20635 (N_20635,N_16739,N_16038);
and U20636 (N_20636,N_15292,N_18010);
nor U20637 (N_20637,N_17423,N_18158);
nand U20638 (N_20638,N_16416,N_15923);
nor U20639 (N_20639,N_16445,N_18142);
nor U20640 (N_20640,N_19185,N_17156);
nor U20641 (N_20641,N_16520,N_19933);
nand U20642 (N_20642,N_17624,N_16202);
nor U20643 (N_20643,N_17958,N_18740);
nand U20644 (N_20644,N_17106,N_15399);
and U20645 (N_20645,N_16627,N_17582);
and U20646 (N_20646,N_19584,N_16745);
and U20647 (N_20647,N_17981,N_19368);
nor U20648 (N_20648,N_15355,N_19289);
and U20649 (N_20649,N_18723,N_16661);
or U20650 (N_20650,N_16809,N_15434);
and U20651 (N_20651,N_15991,N_15190);
nor U20652 (N_20652,N_16079,N_18702);
nand U20653 (N_20653,N_15870,N_16628);
and U20654 (N_20654,N_16885,N_19863);
and U20655 (N_20655,N_15271,N_19447);
xor U20656 (N_20656,N_18775,N_18303);
nand U20657 (N_20657,N_19517,N_18908);
and U20658 (N_20658,N_19432,N_18386);
nand U20659 (N_20659,N_16326,N_19032);
or U20660 (N_20660,N_18561,N_16187);
xnor U20661 (N_20661,N_17227,N_17351);
and U20662 (N_20662,N_16272,N_19773);
and U20663 (N_20663,N_19781,N_15183);
or U20664 (N_20664,N_18573,N_15217);
and U20665 (N_20665,N_19504,N_19034);
and U20666 (N_20666,N_18277,N_19365);
nand U20667 (N_20667,N_16657,N_15909);
nor U20668 (N_20668,N_17980,N_17994);
nor U20669 (N_20669,N_18356,N_15627);
nor U20670 (N_20670,N_19227,N_15522);
nor U20671 (N_20671,N_15808,N_15386);
or U20672 (N_20672,N_16451,N_15197);
xor U20673 (N_20673,N_17839,N_16525);
and U20674 (N_20674,N_15234,N_17569);
xnor U20675 (N_20675,N_15466,N_16705);
or U20676 (N_20676,N_17856,N_15441);
or U20677 (N_20677,N_18030,N_15987);
nor U20678 (N_20678,N_15262,N_18799);
or U20679 (N_20679,N_16999,N_19103);
nor U20680 (N_20680,N_19768,N_17805);
xor U20681 (N_20681,N_19176,N_17525);
nand U20682 (N_20682,N_17253,N_18272);
nor U20683 (N_20683,N_18188,N_16901);
nand U20684 (N_20684,N_16087,N_16698);
xnor U20685 (N_20685,N_19477,N_16246);
xor U20686 (N_20686,N_15692,N_17472);
nand U20687 (N_20687,N_18714,N_17920);
or U20688 (N_20688,N_18827,N_18305);
nor U20689 (N_20689,N_16140,N_16352);
or U20690 (N_20690,N_15379,N_17199);
nand U20691 (N_20691,N_19439,N_19396);
nand U20692 (N_20692,N_19980,N_17567);
and U20693 (N_20693,N_17669,N_16947);
nor U20694 (N_20694,N_18675,N_18732);
xnor U20695 (N_20695,N_16651,N_16261);
nor U20696 (N_20696,N_16942,N_15922);
or U20697 (N_20697,N_17029,N_18935);
or U20698 (N_20698,N_17969,N_15058);
xnor U20699 (N_20699,N_17327,N_15314);
or U20700 (N_20700,N_19861,N_15477);
nand U20701 (N_20701,N_18351,N_17802);
nor U20702 (N_20702,N_18690,N_15585);
nand U20703 (N_20703,N_15065,N_18155);
nand U20704 (N_20704,N_18058,N_18110);
or U20705 (N_20705,N_16962,N_19936);
nand U20706 (N_20706,N_16492,N_19344);
nor U20707 (N_20707,N_19842,N_18803);
or U20708 (N_20708,N_16403,N_15343);
and U20709 (N_20709,N_19275,N_19636);
nor U20710 (N_20710,N_18811,N_16285);
and U20711 (N_20711,N_18007,N_18726);
nor U20712 (N_20712,N_16090,N_15928);
or U20713 (N_20713,N_16952,N_19675);
nand U20714 (N_20714,N_15580,N_19218);
and U20715 (N_20715,N_17780,N_18330);
nor U20716 (N_20716,N_17042,N_19940);
nor U20717 (N_20717,N_15136,N_17636);
and U20718 (N_20718,N_17613,N_19251);
xor U20719 (N_20719,N_16621,N_19885);
nand U20720 (N_20720,N_15431,N_19053);
xnor U20721 (N_20721,N_18789,N_16816);
nand U20722 (N_20722,N_18001,N_16958);
nor U20723 (N_20723,N_19372,N_16490);
and U20724 (N_20724,N_18311,N_18496);
and U20725 (N_20725,N_17170,N_15229);
nor U20726 (N_20726,N_19761,N_15370);
nand U20727 (N_20727,N_19024,N_16918);
nand U20728 (N_20728,N_17017,N_19799);
and U20729 (N_20729,N_15873,N_17512);
or U20730 (N_20730,N_15541,N_15250);
nand U20731 (N_20731,N_17298,N_18134);
or U20732 (N_20732,N_16198,N_15521);
and U20733 (N_20733,N_18088,N_16993);
nor U20734 (N_20734,N_18781,N_16634);
and U20735 (N_20735,N_17575,N_16171);
nand U20736 (N_20736,N_15456,N_18416);
nor U20737 (N_20737,N_19978,N_16803);
nand U20738 (N_20738,N_18539,N_17940);
or U20739 (N_20739,N_18904,N_19336);
nand U20740 (N_20740,N_16133,N_15891);
xor U20741 (N_20741,N_18510,N_15651);
nor U20742 (N_20742,N_15933,N_18444);
and U20743 (N_20743,N_15980,N_19346);
nand U20744 (N_20744,N_19789,N_16715);
xor U20745 (N_20745,N_16292,N_18914);
nor U20746 (N_20746,N_17731,N_16151);
or U20747 (N_20747,N_17014,N_19513);
nand U20748 (N_20748,N_17101,N_15323);
or U20749 (N_20749,N_15598,N_18417);
and U20750 (N_20750,N_15578,N_15902);
or U20751 (N_20751,N_17476,N_15471);
nor U20752 (N_20752,N_19179,N_15635);
xnor U20753 (N_20753,N_15778,N_17684);
nor U20754 (N_20754,N_19090,N_18604);
and U20755 (N_20755,N_17060,N_19351);
xor U20756 (N_20756,N_15589,N_17093);
nand U20757 (N_20757,N_15446,N_15848);
or U20758 (N_20758,N_17702,N_15768);
nand U20759 (N_20759,N_15857,N_16926);
xor U20760 (N_20760,N_16493,N_15731);
nor U20761 (N_20761,N_19701,N_19616);
or U20762 (N_20762,N_18411,N_19565);
xnor U20763 (N_20763,N_15259,N_17329);
xor U20764 (N_20764,N_19835,N_15925);
xor U20765 (N_20765,N_19058,N_16981);
or U20766 (N_20766,N_18404,N_19017);
nand U20767 (N_20767,N_17657,N_18019);
nor U20768 (N_20768,N_15415,N_18785);
nor U20769 (N_20769,N_18910,N_18023);
nor U20770 (N_20770,N_18376,N_19593);
xnor U20771 (N_20771,N_15020,N_18985);
xnor U20772 (N_20772,N_15037,N_17152);
nand U20773 (N_20773,N_18741,N_15337);
xor U20774 (N_20774,N_15547,N_19101);
nand U20775 (N_20775,N_16613,N_18005);
nand U20776 (N_20776,N_18828,N_18318);
nand U20777 (N_20777,N_16549,N_19083);
and U20778 (N_20778,N_18753,N_15236);
and U20779 (N_20779,N_19843,N_17133);
or U20780 (N_20780,N_17377,N_16245);
nor U20781 (N_20781,N_15905,N_19753);
or U20782 (N_20782,N_18078,N_16041);
and U20783 (N_20783,N_17631,N_19866);
or U20784 (N_20784,N_17487,N_16626);
and U20785 (N_20785,N_15572,N_18790);
nor U20786 (N_20786,N_16212,N_17411);
nor U20787 (N_20787,N_17964,N_15359);
nand U20788 (N_20788,N_16900,N_17764);
xor U20789 (N_20789,N_15829,N_16813);
nand U20790 (N_20790,N_16770,N_16065);
or U20791 (N_20791,N_18688,N_17100);
nor U20792 (N_20792,N_15326,N_19451);
or U20793 (N_20793,N_15605,N_18253);
nand U20794 (N_20794,N_16980,N_15086);
or U20795 (N_20795,N_19301,N_17595);
nor U20796 (N_20796,N_19145,N_17509);
or U20797 (N_20797,N_16014,N_16137);
nor U20798 (N_20798,N_18877,N_15004);
or U20799 (N_20799,N_19973,N_18077);
or U20800 (N_20800,N_17875,N_19375);
or U20801 (N_20801,N_17591,N_19259);
and U20802 (N_20802,N_19818,N_19770);
xor U20803 (N_20803,N_16329,N_18585);
nor U20804 (N_20804,N_17038,N_19579);
xor U20805 (N_20805,N_19650,N_18770);
xor U20806 (N_20806,N_18662,N_19318);
nor U20807 (N_20807,N_18168,N_17900);
nor U20808 (N_20808,N_18966,N_16130);
xor U20809 (N_20809,N_17471,N_19510);
or U20810 (N_20810,N_18183,N_19772);
and U20811 (N_20811,N_16869,N_17554);
nand U20812 (N_20812,N_17989,N_19904);
or U20813 (N_20813,N_15710,N_19112);
and U20814 (N_20814,N_19826,N_17513);
and U20815 (N_20815,N_19199,N_15523);
nand U20816 (N_20816,N_16945,N_19719);
or U20817 (N_20817,N_17588,N_17388);
nand U20818 (N_20818,N_19069,N_15931);
xnor U20819 (N_20819,N_19647,N_18264);
or U20820 (N_20820,N_19485,N_15674);
nor U20821 (N_20821,N_17283,N_17858);
nand U20822 (N_20822,N_16579,N_16561);
nor U20823 (N_20823,N_19767,N_16772);
nand U20824 (N_20824,N_19925,N_19976);
nand U20825 (N_20825,N_18457,N_17709);
nand U20826 (N_20826,N_17362,N_18062);
nand U20827 (N_20827,N_16252,N_19592);
xnor U20828 (N_20828,N_19653,N_17831);
nor U20829 (N_20829,N_18772,N_18044);
or U20830 (N_20830,N_15735,N_15779);
or U20831 (N_20831,N_18243,N_19809);
or U20832 (N_20832,N_16176,N_18973);
or U20833 (N_20833,N_15549,N_19883);
nor U20834 (N_20834,N_16473,N_19461);
nand U20835 (N_20835,N_17544,N_15723);
or U20836 (N_20836,N_19235,N_15133);
or U20837 (N_20837,N_19271,N_19296);
nand U20838 (N_20838,N_16582,N_19944);
or U20839 (N_20839,N_16355,N_18509);
nand U20840 (N_20840,N_18637,N_17270);
or U20841 (N_20841,N_19370,N_17011);
and U20842 (N_20842,N_17067,N_17526);
or U20843 (N_20843,N_19280,N_19501);
nor U20844 (N_20844,N_15519,N_16385);
nand U20845 (N_20845,N_15449,N_16078);
and U20846 (N_20846,N_16864,N_17139);
nand U20847 (N_20847,N_19990,N_19019);
nor U20848 (N_20848,N_19029,N_18849);
nand U20849 (N_20849,N_18118,N_19558);
and U20850 (N_20850,N_15228,N_19746);
nand U20851 (N_20851,N_18918,N_16146);
nand U20852 (N_20852,N_15194,N_19265);
or U20853 (N_20853,N_18609,N_16460);
xor U20854 (N_20854,N_15329,N_17749);
nand U20855 (N_20855,N_15595,N_18257);
nand U20856 (N_20856,N_15514,N_19237);
or U20857 (N_20857,N_15851,N_15644);
xor U20858 (N_20858,N_15312,N_17147);
or U20859 (N_20859,N_17257,N_16738);
and U20860 (N_20860,N_17658,N_17389);
nand U20861 (N_20861,N_18051,N_18237);
xor U20862 (N_20862,N_16503,N_17751);
and U20863 (N_20863,N_19655,N_16364);
or U20864 (N_20864,N_18226,N_18306);
nand U20865 (N_20865,N_18449,N_17516);
and U20866 (N_20866,N_18130,N_17518);
or U20867 (N_20867,N_17911,N_19611);
nand U20868 (N_20868,N_17124,N_19140);
nand U20869 (N_20869,N_19908,N_17978);
or U20870 (N_20870,N_19082,N_19300);
nand U20871 (N_20871,N_19742,N_19939);
nand U20872 (N_20872,N_15113,N_19248);
or U20873 (N_20873,N_18819,N_17849);
nor U20874 (N_20874,N_18760,N_19358);
or U20875 (N_20875,N_18898,N_19262);
nand U20876 (N_20876,N_16003,N_18959);
and U20877 (N_20877,N_16410,N_15913);
or U20878 (N_20878,N_15334,N_15104);
or U20879 (N_20879,N_17409,N_17168);
or U20880 (N_20880,N_15390,N_18162);
or U20881 (N_20881,N_15697,N_17666);
nor U20882 (N_20882,N_18218,N_15526);
nor U20883 (N_20883,N_16278,N_16861);
or U20884 (N_20884,N_16620,N_19683);
or U20885 (N_20885,N_15955,N_15074);
xnor U20886 (N_20886,N_17706,N_16236);
xnor U20887 (N_20887,N_15260,N_18882);
xnor U20888 (N_20888,N_15666,N_19727);
nand U20889 (N_20889,N_18493,N_15721);
and U20890 (N_20890,N_18742,N_15282);
and U20891 (N_20891,N_19664,N_17796);
xor U20892 (N_20892,N_19849,N_18418);
and U20893 (N_20893,N_17259,N_15542);
and U20894 (N_20894,N_16064,N_16791);
nor U20895 (N_20895,N_19231,N_18822);
nand U20896 (N_20896,N_18350,N_16711);
nor U20897 (N_20897,N_18122,N_17560);
nand U20898 (N_20898,N_18517,N_16684);
nor U20899 (N_20899,N_16615,N_17057);
nand U20900 (N_20900,N_19010,N_17417);
nor U20901 (N_20901,N_16447,N_17528);
and U20902 (N_20902,N_19652,N_16311);
or U20903 (N_20903,N_18235,N_17297);
and U20904 (N_20904,N_16967,N_17605);
or U20905 (N_20905,N_17012,N_16693);
nand U20906 (N_20906,N_15703,N_16281);
nor U20907 (N_20907,N_16359,N_16397);
or U20908 (N_20908,N_17671,N_16122);
nor U20909 (N_20909,N_17281,N_15276);
and U20910 (N_20910,N_16828,N_16823);
or U20911 (N_20911,N_16748,N_16009);
nand U20912 (N_20912,N_17126,N_15042);
and U20913 (N_20913,N_19684,N_16752);
or U20914 (N_20914,N_16131,N_15900);
and U20915 (N_20915,N_15423,N_18611);
or U20916 (N_20916,N_15056,N_17879);
or U20917 (N_20917,N_16455,N_16894);
nor U20918 (N_20918,N_17515,N_19800);
nand U20919 (N_20919,N_18040,N_17625);
or U20920 (N_20920,N_19638,N_16575);
nand U20921 (N_20921,N_18837,N_19471);
nor U20922 (N_20922,N_19728,N_19909);
nor U20923 (N_20923,N_17323,N_16307);
nand U20924 (N_20924,N_19162,N_16939);
nand U20925 (N_20925,N_18312,N_18542);
or U20926 (N_20926,N_18197,N_18371);
and U20927 (N_20927,N_18414,N_17140);
or U20928 (N_20928,N_18465,N_19563);
xnor U20929 (N_20929,N_17519,N_18645);
or U20930 (N_20930,N_16439,N_17681);
nor U20931 (N_20931,N_17715,N_15640);
and U20932 (N_20932,N_16856,N_17033);
xnor U20933 (N_20933,N_16784,N_19431);
nor U20934 (N_20934,N_15800,N_15660);
nor U20935 (N_20935,N_17214,N_17402);
or U20936 (N_20936,N_17581,N_19110);
or U20937 (N_20937,N_17123,N_17157);
or U20938 (N_20938,N_18681,N_17151);
or U20939 (N_20939,N_19660,N_16004);
or U20940 (N_20940,N_18454,N_18324);
and U20941 (N_20941,N_16021,N_16897);
nor U20942 (N_20942,N_18879,N_18962);
nand U20943 (N_20943,N_19743,N_19168);
xor U20944 (N_20944,N_18071,N_19808);
and U20945 (N_20945,N_17586,N_17844);
or U20946 (N_20946,N_19811,N_18676);
nand U20947 (N_20947,N_16994,N_18397);
and U20948 (N_20948,N_16328,N_15213);
and U20949 (N_20949,N_17540,N_16230);
nor U20950 (N_20950,N_17348,N_19769);
and U20951 (N_20951,N_17404,N_17174);
nand U20952 (N_20952,N_18287,N_15453);
and U20953 (N_20953,N_16629,N_17961);
and U20954 (N_20954,N_16441,N_19778);
and U20955 (N_20955,N_16390,N_16875);
and U20956 (N_20956,N_19677,N_18975);
nand U20957 (N_20957,N_17928,N_15027);
nor U20958 (N_20958,N_18974,N_16602);
or U20959 (N_20959,N_18146,N_19246);
and U20960 (N_20960,N_15076,N_19027);
nand U20961 (N_20961,N_16631,N_16826);
nand U20962 (N_20962,N_17508,N_15226);
or U20963 (N_20963,N_15335,N_15607);
and U20964 (N_20964,N_15968,N_16616);
or U20965 (N_20965,N_16027,N_19880);
or U20966 (N_20966,N_15853,N_17431);
or U20967 (N_20967,N_15994,N_15664);
nand U20968 (N_20968,N_15305,N_15688);
xnor U20969 (N_20969,N_19779,N_18125);
nand U20970 (N_20970,N_15562,N_16154);
nor U20971 (N_20971,N_16690,N_18248);
nand U20972 (N_20972,N_19020,N_16622);
or U20973 (N_20973,N_19993,N_15447);
nand U20974 (N_20974,N_16222,N_18316);
and U20975 (N_20975,N_18991,N_17736);
xnor U20976 (N_20976,N_18176,N_18655);
and U20977 (N_20977,N_17461,N_19644);
nor U20978 (N_20978,N_16428,N_19618);
nand U20979 (N_20979,N_19122,N_18978);
nor U20980 (N_20980,N_16855,N_18885);
and U20981 (N_20981,N_18119,N_16423);
nand U20982 (N_20982,N_17974,N_18902);
nand U20983 (N_20983,N_18638,N_17622);
and U20984 (N_20984,N_17646,N_19131);
nor U20985 (N_20985,N_16159,N_16317);
and U20986 (N_20986,N_15401,N_17473);
and U20987 (N_20987,N_17577,N_18475);
nor U20988 (N_20988,N_18451,N_15285);
xor U20989 (N_20989,N_18074,N_19484);
xor U20990 (N_20990,N_18900,N_17435);
nor U20991 (N_20991,N_19687,N_18281);
or U20992 (N_20992,N_16890,N_17857);
and U20993 (N_20993,N_18239,N_17683);
nand U20994 (N_20994,N_19325,N_18839);
or U20995 (N_20995,N_17688,N_18565);
and U20996 (N_20996,N_19966,N_19422);
nor U20997 (N_20997,N_19700,N_16343);
xnor U20998 (N_20998,N_17092,N_18147);
xnor U20999 (N_20999,N_16567,N_18797);
nand U21000 (N_21000,N_15512,N_17655);
or U21001 (N_21001,N_17725,N_16175);
nor U21002 (N_21002,N_17695,N_19157);
or U21003 (N_21003,N_17167,N_17111);
nor U21004 (N_21004,N_18709,N_16589);
or U21005 (N_21005,N_17562,N_17682);
nand U21006 (N_21006,N_15195,N_16895);
or U21007 (N_21007,N_18012,N_19954);
nor U21008 (N_21008,N_16026,N_16775);
or U21009 (N_21009,N_19852,N_18896);
nand U21010 (N_21010,N_16360,N_17807);
nand U21011 (N_21011,N_16107,N_16491);
nand U21012 (N_21012,N_16301,N_15752);
nand U21013 (N_21013,N_15246,N_16767);
nand U21014 (N_21014,N_16708,N_15372);
and U21015 (N_21015,N_15003,N_19679);
nor U21016 (N_21016,N_17221,N_19820);
nand U21017 (N_21017,N_19887,N_16502);
nor U21018 (N_21018,N_19377,N_15459);
nor U21019 (N_21019,N_16974,N_16670);
or U21020 (N_21020,N_19244,N_15389);
and U21021 (N_21021,N_16052,N_18692);
and U21022 (N_21022,N_19965,N_15026);
nand U21023 (N_21023,N_19552,N_16249);
and U21024 (N_21024,N_15118,N_19409);
nand U21025 (N_21025,N_15132,N_16239);
and U21026 (N_21026,N_17629,N_18881);
and U21027 (N_21027,N_19057,N_17192);
nor U21028 (N_21028,N_16744,N_19430);
and U21029 (N_21029,N_16891,N_15267);
or U21030 (N_21030,N_16555,N_17722);
nand U21031 (N_21031,N_18871,N_19488);
nor U21032 (N_21032,N_16012,N_18883);
nand U21033 (N_21033,N_17837,N_17219);
nor U21034 (N_21034,N_18699,N_19066);
or U21035 (N_21035,N_17743,N_17225);
or U21036 (N_21036,N_16663,N_18607);
or U21037 (N_21037,N_18263,N_17698);
or U21038 (N_21038,N_17349,N_17494);
nor U21039 (N_21039,N_19538,N_18981);
or U21040 (N_21040,N_16076,N_16524);
xnor U21041 (N_21041,N_17825,N_18232);
xor U21042 (N_21042,N_18221,N_16269);
nor U21043 (N_21043,N_16982,N_16940);
nor U21044 (N_21044,N_16235,N_15347);
nand U21045 (N_21045,N_15212,N_17668);
nor U21046 (N_21046,N_16843,N_16442);
nor U21047 (N_21047,N_15048,N_17628);
and U21048 (N_21048,N_17452,N_15244);
nor U21049 (N_21049,N_16858,N_16284);
or U21050 (N_21050,N_19763,N_17757);
nand U21051 (N_21051,N_15838,N_16211);
nand U21052 (N_21052,N_18402,N_19332);
and U21053 (N_21053,N_15559,N_17171);
nor U21054 (N_21054,N_17759,N_17503);
and U21055 (N_21055,N_19639,N_18952);
nand U21056 (N_21056,N_16916,N_18476);
nand U21057 (N_21057,N_16091,N_15740);
nor U21058 (N_21058,N_18880,N_17862);
and U21059 (N_21059,N_15099,N_19129);
nor U21060 (N_21060,N_17971,N_15614);
and U21061 (N_21061,N_15907,N_15709);
nand U21062 (N_21062,N_15846,N_16461);
nor U21063 (N_21063,N_19425,N_15364);
or U21064 (N_21064,N_16529,N_18396);
nand U21065 (N_21065,N_16838,N_15584);
or U21066 (N_21066,N_19467,N_16263);
nor U21067 (N_21067,N_16135,N_16924);
nand U21068 (N_21068,N_19143,N_17641);
or U21069 (N_21069,N_15534,N_19724);
nand U21070 (N_21070,N_19254,N_15826);
xor U21071 (N_21071,N_18979,N_18691);
or U21072 (N_21072,N_16806,N_16121);
and U21073 (N_21073,N_18976,N_18435);
nor U21074 (N_21074,N_18769,N_18447);
and U21075 (N_21075,N_17739,N_15266);
nor U21076 (N_21076,N_15159,N_19107);
and U21077 (N_21077,N_17498,N_15539);
and U21078 (N_21078,N_16370,N_17717);
nand U21079 (N_21079,N_16725,N_16020);
nand U21080 (N_21080,N_15591,N_15764);
nand U21081 (N_21081,N_17482,N_19744);
or U21082 (N_21082,N_17403,N_19481);
and U21083 (N_21083,N_16824,N_15587);
or U21084 (N_21084,N_16338,N_19304);
nor U21085 (N_21085,N_18175,N_17306);
nand U21086 (N_21086,N_17787,N_16051);
nor U21087 (N_21087,N_17357,N_18343);
nor U21088 (N_21088,N_18453,N_15424);
or U21089 (N_21089,N_16477,N_19755);
nor U21090 (N_21090,N_19367,N_18013);
or U21091 (N_21091,N_18868,N_17380);
and U21092 (N_21092,N_15428,N_16977);
and U21093 (N_21093,N_17860,N_18934);
or U21094 (N_21094,N_19291,N_18492);
or U21095 (N_21095,N_19740,N_16474);
nor U21096 (N_21096,N_15781,N_17228);
xor U21097 (N_21097,N_17703,N_17884);
and U21098 (N_21098,N_15178,N_17134);
or U21099 (N_21099,N_17504,N_15744);
nor U21100 (N_21100,N_16000,N_19338);
or U21101 (N_21101,N_16961,N_15265);
or U21102 (N_21102,N_19170,N_15188);
and U21103 (N_21103,N_19294,N_16932);
or U21104 (N_21104,N_19914,N_15371);
and U21105 (N_21105,N_16706,N_17485);
nand U21106 (N_21106,N_18075,N_17745);
or U21107 (N_21107,N_16724,N_19704);
nor U21108 (N_21108,N_16968,N_18657);
nor U21109 (N_21109,N_15759,N_15168);
or U21110 (N_21110,N_17638,N_15280);
nor U21111 (N_21111,N_16495,N_19361);
nor U21112 (N_21112,N_19586,N_17890);
nand U21113 (N_21113,N_17843,N_17393);
nor U21114 (N_21114,N_17619,N_18748);
nand U21115 (N_21115,N_19441,N_16216);
or U21116 (N_21116,N_15097,N_17991);
nor U21117 (N_21117,N_16062,N_17902);
or U21118 (N_21118,N_18052,N_15303);
nor U21119 (N_21119,N_17394,N_15385);
nor U21120 (N_21120,N_16289,N_19487);
nand U21121 (N_21121,N_15077,N_17341);
xnor U21122 (N_21122,N_18759,N_19678);
and U21123 (N_21123,N_16120,N_18111);
nor U21124 (N_21124,N_17811,N_18694);
xor U21125 (N_21125,N_15501,N_17287);
xnor U21126 (N_21126,N_18525,N_15269);
xor U21127 (N_21127,N_15956,N_18295);
and U21128 (N_21128,N_16732,N_15148);
or U21129 (N_21129,N_17529,N_16966);
xnor U21130 (N_21130,N_19546,N_16879);
nor U21131 (N_21131,N_19895,N_15490);
xor U21132 (N_21132,N_17534,N_18107);
nand U21133 (N_21133,N_16318,N_16054);
nor U21134 (N_21134,N_19535,N_16181);
nand U21135 (N_21135,N_16233,N_19378);
nand U21136 (N_21136,N_15008,N_16590);
and U21137 (N_21137,N_18795,N_16907);
nor U21138 (N_21138,N_15842,N_19238);
nor U21139 (N_21139,N_19319,N_17421);
or U21140 (N_21140,N_15705,N_16494);
nor U21141 (N_21141,N_17153,N_19307);
xor U21142 (N_21142,N_19139,N_15240);
nor U21143 (N_21143,N_18829,N_17918);
and U21144 (N_21144,N_16836,N_18838);
and U21145 (N_21145,N_18108,N_15722);
nor U21146 (N_21146,N_15983,N_19603);
and U21147 (N_21147,N_17965,N_17986);
nand U21148 (N_21148,N_17434,N_16379);
nand U21149 (N_21149,N_17502,N_19815);
nor U21150 (N_21150,N_19428,N_17679);
or U21151 (N_21151,N_17074,N_16862);
or U21152 (N_21152,N_17208,N_17917);
and U21153 (N_21153,N_18815,N_18642);
nor U21154 (N_21154,N_15790,N_16341);
nand U21155 (N_21155,N_17275,N_15661);
nand U21156 (N_21156,N_15691,N_19146);
and U21157 (N_21157,N_18606,N_19643);
nor U21158 (N_21158,N_15763,N_15289);
nand U21159 (N_21159,N_15895,N_15400);
xnor U21160 (N_21160,N_19255,N_15798);
nand U21161 (N_21161,N_16086,N_16094);
nor U21162 (N_21162,N_17993,N_16733);
nand U21163 (N_21163,N_18744,N_16182);
xor U21164 (N_21164,N_16511,N_19068);
nand U21165 (N_21165,N_16501,N_19317);
nand U21166 (N_21166,N_17774,N_19272);
or U21167 (N_21167,N_19766,N_18192);
nor U21168 (N_21168,N_19798,N_15203);
nor U21169 (N_21169,N_16424,N_16709);
xnor U21170 (N_21170,N_19152,N_15251);
xnor U21171 (N_21171,N_16431,N_19369);
or U21172 (N_21172,N_16097,N_17269);
nor U21173 (N_21173,N_15414,N_18687);
or U21174 (N_21174,N_18055,N_15843);
nand U21175 (N_21175,N_17733,N_15648);
nand U21176 (N_21176,N_15582,N_16912);
nand U21177 (N_21177,N_17047,N_18409);
xnor U21178 (N_21178,N_18923,N_17185);
nor U21179 (N_21179,N_17634,N_15505);
xnor U21180 (N_21180,N_15714,N_15409);
and U21181 (N_21181,N_18567,N_18313);
nand U21182 (N_21182,N_19749,N_17302);
or U21183 (N_21183,N_15754,N_15223);
nand U21184 (N_21184,N_15384,N_16393);
xor U21185 (N_21185,N_16654,N_18547);
xor U21186 (N_21186,N_17265,N_15435);
xnor U21187 (N_21187,N_16729,N_16196);
or U21188 (N_21188,N_18364,N_15258);
or U21189 (N_21189,N_18630,N_17626);
xnor U21190 (N_21190,N_19383,N_18365);
and U21191 (N_21191,N_17700,N_17459);
nor U21192 (N_21192,N_19384,N_18171);
and U21193 (N_21193,N_15867,N_19113);
or U21194 (N_21194,N_19648,N_19033);
nand U21195 (N_21195,N_16485,N_15916);
nor U21196 (N_21196,N_15366,N_19011);
and U21197 (N_21197,N_18757,N_16480);
or U21198 (N_21198,N_15583,N_18566);
and U21199 (N_21199,N_16205,N_17999);
or U21200 (N_21200,N_18347,N_18380);
xnor U21201 (N_21201,N_19226,N_17408);
and U21202 (N_21202,N_18274,N_18429);
nand U21203 (N_21203,N_15834,N_17450);
or U21204 (N_21204,N_15970,N_19134);
nor U21205 (N_21205,N_17127,N_18821);
or U21206 (N_21206,N_16356,N_19528);
nand U21207 (N_21207,N_16025,N_18940);
nand U21208 (N_21208,N_19988,N_16185);
or U21209 (N_21209,N_15753,N_15775);
nand U21210 (N_21210,N_18560,N_18749);
nand U21211 (N_21211,N_18658,N_18521);
nand U21212 (N_21212,N_16368,N_17639);
nand U21213 (N_21213,N_17291,N_16779);
and U21214 (N_21214,N_17742,N_17665);
or U21215 (N_21215,N_18761,N_15263);
nor U21216 (N_21216,N_15604,N_19363);
and U21217 (N_21217,N_19405,N_15772);
or U21218 (N_21218,N_18507,N_17551);
nor U21219 (N_21219,N_17748,N_15600);
nor U21220 (N_21220,N_15049,N_15990);
and U21221 (N_21221,N_19847,N_19879);
nand U21222 (N_21222,N_18225,N_19864);
nand U21223 (N_21223,N_18847,N_17701);
nor U21224 (N_21224,N_16063,N_18085);
nand U21225 (N_21225,N_18141,N_16372);
or U21226 (N_21226,N_17212,N_16760);
nor U21227 (N_21227,N_15919,N_18798);
or U21228 (N_21228,N_19036,N_16251);
and U21229 (N_21229,N_16544,N_19065);
nand U21230 (N_21230,N_19412,N_16564);
nor U21231 (N_21231,N_18297,N_16381);
or U21232 (N_21232,N_15992,N_16889);
xor U21233 (N_21233,N_16973,N_16132);
nand U21234 (N_21234,N_16583,N_17440);
or U21235 (N_21235,N_18153,N_19580);
nand U21236 (N_21236,N_18780,N_17707);
and U21237 (N_21237,N_18054,N_16630);
or U21238 (N_21238,N_19111,N_16056);
and U21239 (N_21239,N_15892,N_17492);
and U21240 (N_21240,N_17175,N_15092);
and U21241 (N_21241,N_16297,N_18541);
nand U21242 (N_21242,N_16082,N_18491);
or U21243 (N_21243,N_17536,N_19452);
nor U21244 (N_21244,N_17867,N_15619);
or U21245 (N_21245,N_17373,N_17859);
and U21246 (N_21246,N_15967,N_17830);
and U21247 (N_21247,N_15606,N_19116);
xnor U21248 (N_21248,N_19702,N_16344);
nor U21249 (N_21249,N_16518,N_17110);
nand U21250 (N_21250,N_16257,N_15429);
or U21251 (N_21251,N_18601,N_18478);
xor U21252 (N_21252,N_16898,N_18331);
or U21253 (N_21253,N_16560,N_17627);
xnor U21254 (N_21254,N_19100,N_18322);
or U21255 (N_21255,N_19642,N_17689);
and U21256 (N_21256,N_15985,N_16788);
nand U21257 (N_21257,N_18848,N_17240);
nor U21258 (N_21258,N_15403,N_16160);
or U21259 (N_21259,N_17714,N_19206);
and U21260 (N_21260,N_15596,N_17044);
nor U21261 (N_21261,N_15809,N_16243);
and U21262 (N_21262,N_15082,N_18673);
nand U21263 (N_21263,N_17352,N_15184);
nor U21264 (N_21264,N_15615,N_17068);
nand U21265 (N_21265,N_17612,N_19314);
and U21266 (N_21266,N_17673,N_18783);
and U21267 (N_21267,N_15040,N_18893);
or U21268 (N_21268,N_16177,N_18916);
nand U21269 (N_21269,N_16666,N_18327);
and U21270 (N_21270,N_19915,N_19942);
and U21271 (N_21271,N_15813,N_16496);
nor U21272 (N_21272,N_18915,N_19054);
or U21273 (N_21273,N_15270,N_17615);
or U21274 (N_21274,N_16541,N_18927);
xnor U21275 (N_21275,N_19480,N_15780);
and U21276 (N_21276,N_19888,N_18269);
or U21277 (N_21277,N_16751,N_17339);
nand U21278 (N_21278,N_18875,N_17996);
nand U21279 (N_21279,N_19374,N_18664);
nor U21280 (N_21280,N_17931,N_18394);
nand U21281 (N_21281,N_19979,N_19859);
or U21282 (N_21282,N_15081,N_16102);
xnor U21283 (N_21283,N_16053,N_17446);
or U21284 (N_21284,N_18529,N_19106);
nor U21285 (N_21285,N_17847,N_15972);
nor U21286 (N_21286,N_18382,N_16136);
xnor U21287 (N_21287,N_17278,N_19440);
and U21288 (N_21288,N_19349,N_15797);
nor U21289 (N_21289,N_17848,N_15059);
and U21290 (N_21290,N_17344,N_18140);
or U21291 (N_21291,N_18646,N_16519);
or U21292 (N_21292,N_15969,N_15387);
and U21293 (N_21293,N_19532,N_18513);
or U21294 (N_21294,N_16505,N_18917);
or U21295 (N_21295,N_15845,N_15153);
nand U21296 (N_21296,N_18844,N_19198);
nand U21297 (N_21297,N_18407,N_15974);
or U21298 (N_21298,N_18924,N_18659);
nor U21299 (N_21299,N_16597,N_17573);
nand U21300 (N_21300,N_17149,N_19889);
nand U21301 (N_21301,N_15847,N_18863);
or U21302 (N_21302,N_16671,N_17938);
nor U21303 (N_21303,N_16113,N_19857);
xnor U21304 (N_21304,N_16860,N_19154);
nand U21305 (N_21305,N_17256,N_19875);
or U21306 (N_21306,N_15494,N_15140);
nor U21307 (N_21307,N_17364,N_19270);
or U21308 (N_21308,N_16714,N_16740);
nor U21309 (N_21309,N_15193,N_15383);
or U21310 (N_21310,N_17486,N_15225);
nand U21311 (N_21311,N_19164,N_17785);
nand U21312 (N_21312,N_15171,N_18621);
nand U21313 (N_21313,N_16058,N_16047);
nor U21314 (N_21314,N_19522,N_15789);
nand U21315 (N_21315,N_18859,N_17077);
and U21316 (N_21316,N_17206,N_18200);
and U21317 (N_21317,N_15520,N_18046);
and U21318 (N_21318,N_17705,N_19750);
and U21319 (N_21319,N_15623,N_19943);
nand U21320 (N_21320,N_16013,N_16633);
or U21321 (N_21321,N_18498,N_15199);
and U21322 (N_21322,N_16006,N_16639);
or U21323 (N_21323,N_19161,N_18472);
nand U21324 (N_21324,N_18639,N_19575);
nand U21325 (N_21325,N_17255,N_16067);
nor U21326 (N_21326,N_18970,N_19518);
nor U21327 (N_21327,N_16667,N_15566);
xnor U21328 (N_21328,N_17821,N_15982);
xor U21329 (N_21329,N_19570,N_19046);
or U21330 (N_21330,N_15495,N_18410);
nand U21331 (N_21331,N_19795,N_18377);
nor U21332 (N_21332,N_17304,N_19009);
xor U21333 (N_21333,N_16109,N_15849);
nor U21334 (N_21334,N_16686,N_19355);
or U21335 (N_21335,N_17135,N_15356);
and U21336 (N_21336,N_16023,N_15893);
nand U21337 (N_21337,N_19568,N_16790);
xor U21338 (N_21338,N_18794,N_17767);
and U21339 (N_21339,N_16829,N_15463);
and U21340 (N_21340,N_18854,N_18894);
or U21341 (N_21341,N_15033,N_15256);
nor U21342 (N_21342,N_18072,N_17871);
nor U21343 (N_21343,N_15966,N_19128);
nor U21344 (N_21344,N_15264,N_17292);
nand U21345 (N_21345,N_18806,N_19931);
or U21346 (N_21346,N_18989,N_16801);
and U21347 (N_21347,N_17943,N_18603);
nor U21348 (N_21348,N_15352,N_16599);
nor U21349 (N_21349,N_16408,N_15737);
nand U21350 (N_21350,N_19676,N_17941);
or U21351 (N_21351,N_18523,N_19474);
and U21352 (N_21352,N_16173,N_16282);
and U21353 (N_21353,N_18906,N_17254);
nor U21354 (N_21354,N_19649,N_15643);
or U21355 (N_21355,N_15822,N_17084);
xnor U21356 (N_21356,N_16409,N_17574);
or U21357 (N_21357,N_19159,N_15404);
nor U21358 (N_21358,N_16625,N_17967);
nand U21359 (N_21359,N_17609,N_18424);
nor U21360 (N_21360,N_19379,N_15479);
and U21361 (N_21361,N_17458,N_17004);
nor U21362 (N_21362,N_19752,N_18958);
or U21363 (N_21363,N_17648,N_16902);
nor U21364 (N_21364,N_16225,N_19418);
or U21365 (N_21365,N_18128,N_19825);
nor U21366 (N_21366,N_18025,N_16780);
nor U21367 (N_21367,N_19514,N_15500);
and U21368 (N_21368,N_18421,N_16031);
and U21369 (N_21369,N_16481,N_19585);
and U21370 (N_21370,N_18963,N_18721);
or U21371 (N_21371,N_18964,N_16530);
nor U21372 (N_21372,N_19491,N_17947);
or U21373 (N_21373,N_15830,N_15368);
xnor U21374 (N_21374,N_18912,N_18640);
and U21375 (N_21375,N_15450,N_18443);
or U21376 (N_21376,N_16169,N_16688);
nand U21377 (N_21377,N_17061,N_15093);
xnor U21378 (N_21378,N_18288,N_19475);
and U21379 (N_21379,N_18038,N_18080);
nor U21380 (N_21380,N_15279,N_18752);
and U21381 (N_21381,N_17143,N_18170);
or U21382 (N_21382,N_17539,N_16432);
xor U21383 (N_21383,N_17433,N_18870);
nor U21384 (N_21384,N_17176,N_17104);
xnor U21385 (N_21385,N_18731,N_17237);
nand U21386 (N_21386,N_19207,N_17353);
and U21387 (N_21387,N_16336,N_18184);
nor U21388 (N_21388,N_16399,N_17355);
nand U21389 (N_21389,N_17356,N_19959);
nand U21390 (N_21390,N_19794,N_15608);
and U21391 (N_21391,N_17762,N_15525);
nand U21392 (N_21392,N_19026,N_18707);
nand U21393 (N_21393,N_18499,N_17809);
or U21394 (N_21394,N_18242,N_15488);
or U21395 (N_21395,N_17455,N_17102);
or U21396 (N_21396,N_19656,N_16294);
xor U21397 (N_21397,N_15784,N_19886);
xnor U21398 (N_21398,N_19402,N_19031);
or U21399 (N_21399,N_17451,N_17493);
and U21400 (N_21400,N_19080,N_18936);
and U21401 (N_21401,N_16758,N_17798);
nand U21402 (N_21402,N_15844,N_15175);
nand U21403 (N_21403,N_16747,N_18355);
nand U21404 (N_21404,N_17782,N_16976);
xor U21405 (N_21405,N_19183,N_18094);
and U21406 (N_21406,N_18095,N_15689);
or U21407 (N_21407,N_17590,N_18049);
and U21408 (N_21408,N_19997,N_19960);
nand U21409 (N_21409,N_19850,N_16827);
or U21410 (N_21410,N_17899,N_18387);
nor U21411 (N_21411,N_16658,N_16275);
and U21412 (N_21412,N_15567,N_17040);
or U21413 (N_21413,N_18843,N_17370);
xnor U21414 (N_21414,N_17746,N_15915);
or U21415 (N_21415,N_18992,N_15531);
nor U21416 (N_21416,N_16777,N_16911);
xnor U21417 (N_21417,N_19771,N_18081);
xnor U21418 (N_21418,N_19008,N_17136);
nor U21419 (N_21419,N_19673,N_16362);
xnor U21420 (N_21420,N_16270,N_18595);
nor U21421 (N_21421,N_16996,N_17180);
nand U21422 (N_21422,N_18650,N_15876);
nand U21423 (N_21423,N_19786,N_15325);
nand U21424 (N_21424,N_19211,N_15954);
nor U21425 (N_21425,N_15671,N_18901);
nor U21426 (N_21426,N_15810,N_17453);
and U21427 (N_21427,N_16648,N_17959);
nand U21428 (N_21428,N_16156,N_17422);
nand U21429 (N_21429,N_19697,N_15821);
and U21430 (N_21430,N_15257,N_17753);
nor U21431 (N_21431,N_17371,N_18182);
xor U21432 (N_21432,N_16095,N_18004);
and U21433 (N_21433,N_15556,N_17653);
and U21434 (N_21434,N_18754,N_18876);
nor U21435 (N_21435,N_19142,N_15290);
or U21436 (N_21436,N_16116,N_16241);
or U21437 (N_21437,N_19597,N_19133);
nand U21438 (N_21438,N_16008,N_17400);
and U21439 (N_21439,N_17693,N_18440);
or U21440 (N_21440,N_19717,N_19276);
or U21441 (N_21441,N_18131,N_17213);
and U21442 (N_21442,N_19216,N_18987);
and U21443 (N_21443,N_15080,N_15868);
and U21444 (N_21444,N_17096,N_19445);
or U21445 (N_21445,N_18233,N_17420);
xor U21446 (N_21446,N_18677,N_19454);
nor U21447 (N_21447,N_15532,N_19681);
nor U21448 (N_21448,N_19934,N_17640);
nor U21449 (N_21449,N_18725,N_18544);
or U21450 (N_21450,N_16692,N_17686);
and U21451 (N_21451,N_16607,N_18737);
nand U21452 (N_21452,N_16776,N_19894);
nor U21453 (N_21453,N_17419,N_16566);
nand U21454 (N_21454,N_19153,N_16538);
nand U21455 (N_21455,N_15977,N_16074);
and U21456 (N_21456,N_15920,N_19884);
and U21457 (N_21457,N_15307,N_18189);
nor U21458 (N_21458,N_19003,N_17786);
or U21459 (N_21459,N_15179,N_15699);
nor U21460 (N_21460,N_18208,N_16498);
or U21461 (N_21461,N_19400,N_19874);
nand U21462 (N_21462,N_15134,N_15593);
nor U21463 (N_21463,N_15811,N_19747);
or U21464 (N_21464,N_15448,N_15638);
or U21465 (N_21465,N_17896,N_16110);
or U21466 (N_21466,N_18747,N_18619);
xor U21467 (N_21467,N_16935,N_19951);
and U21468 (N_21468,N_19837,N_17095);
and U21469 (N_21469,N_17232,N_18536);
or U21470 (N_21470,N_16743,N_17616);
nand U21471 (N_21471,N_16964,N_19138);
or U21472 (N_21472,N_18602,N_16489);
nand U21473 (N_21473,N_19759,N_17718);
and U21474 (N_21474,N_16126,N_18679);
nor U21475 (N_21475,N_16796,N_16712);
and U21476 (N_21476,N_17374,N_16232);
xor U21477 (N_21477,N_16148,N_18053);
or U21478 (N_21478,N_19821,N_15942);
and U21479 (N_21479,N_15856,N_19464);
nand U21480 (N_21480,N_19891,N_19059);
and U21481 (N_21481,N_18878,N_18285);
xor U21482 (N_21482,N_15725,N_15047);
nand U21483 (N_21483,N_17318,N_15333);
nand U21484 (N_21484,N_19628,N_15198);
and U21485 (N_21485,N_16304,N_19792);
nand U21486 (N_21486,N_18636,N_16528);
or U21487 (N_21487,N_16178,N_16595);
or U21488 (N_21488,N_16305,N_15417);
nor U21489 (N_21489,N_15971,N_18391);
nor U21490 (N_21490,N_16545,N_19654);
nand U21491 (N_21491,N_19540,N_18090);
and U21492 (N_21492,N_16374,N_16540);
and U21493 (N_21493,N_16022,N_16016);
nand U21494 (N_21494,N_17183,N_15044);
xor U21495 (N_21495,N_19328,N_16283);
and U21496 (N_21496,N_16457,N_18861);
nor U21497 (N_21497,N_17236,N_17131);
nor U21498 (N_21498,N_16406,N_17912);
nand U21499 (N_21499,N_17087,N_19055);
nor U21500 (N_21500,N_16015,N_19547);
nor U21501 (N_21501,N_18120,N_16234);
or U21502 (N_21502,N_19735,N_15686);
nand U21503 (N_21503,N_19551,N_17711);
nand U21504 (N_21504,N_15427,N_19666);
nor U21505 (N_21505,N_15777,N_18048);
nor U21506 (N_21506,N_19393,N_19686);
or U21507 (N_21507,N_16844,N_19267);
and U21508 (N_21508,N_16818,N_17677);
or U21509 (N_21509,N_18651,N_17369);
xnor U21510 (N_21510,N_15051,N_18280);
nand U21511 (N_21511,N_17558,N_16841);
and U21512 (N_21512,N_16069,N_19527);
and U21513 (N_21513,N_17121,N_15181);
or U21514 (N_21514,N_19087,N_16611);
and U21515 (N_21515,N_19691,N_16951);
or U21516 (N_21516,N_18907,N_19587);
nand U21517 (N_21517,N_16077,N_17130);
nand U21518 (N_21518,N_18370,N_15344);
and U21519 (N_21519,N_15016,N_15636);
and U21520 (N_21520,N_17260,N_19426);
and U21521 (N_21521,N_16581,N_19404);
or U21522 (N_21522,N_15804,N_15252);
nor U21523 (N_21523,N_15667,N_16405);
nor U21524 (N_21524,N_16957,N_15546);
nand U21525 (N_21525,N_19282,N_18593);
nand U21526 (N_21526,N_19483,N_19233);
nand U21527 (N_21527,N_18479,N_18328);
or U21528 (N_21528,N_17901,N_17580);
and U21529 (N_21529,N_19446,N_16467);
and U21530 (N_21530,N_17929,N_18279);
nor U21531 (N_21531,N_17511,N_16547);
xnor U21532 (N_21532,N_17317,N_15336);
nand U21533 (N_21533,N_17747,N_19310);
and U21534 (N_21534,N_16337,N_19288);
nand U21535 (N_21535,N_19025,N_17806);
nor U21536 (N_21536,N_15749,N_17075);
nand U21537 (N_21537,N_18138,N_18733);
nor U21538 (N_21538,N_16837,N_17680);
nand U21539 (N_21539,N_16299,N_19508);
and U21540 (N_21540,N_16072,N_19049);
nand U21541 (N_21541,N_15189,N_15706);
nor U21542 (N_21542,N_18103,N_17307);
nand U21543 (N_21543,N_19071,N_17069);
nor U21544 (N_21544,N_19120,N_18855);
nand U21545 (N_21545,N_18977,N_17320);
or U21546 (N_21546,N_15060,N_18057);
nand U21547 (N_21547,N_19266,N_16170);
xnor U21548 (N_21548,N_17561,N_16096);
nand U21549 (N_21549,N_16209,N_15535);
nand U21550 (N_21550,N_17674,N_18031);
or U21551 (N_21551,N_19421,N_15486);
xnor U21552 (N_21552,N_19571,N_15762);
or U21553 (N_21553,N_19098,N_17632);
and U21554 (N_21554,N_15296,N_19745);
and U21555 (N_21555,N_17754,N_16158);
nor U21556 (N_21556,N_19817,N_19126);
nor U21557 (N_21557,N_18984,N_15543);
nand U21558 (N_21558,N_15338,N_16168);
or U21559 (N_21559,N_17850,N_19434);
and U21560 (N_21560,N_19897,N_16617);
nand U21561 (N_21561,N_18228,N_19329);
nand U21562 (N_21562,N_18704,N_18932);
and U21563 (N_21563,N_17112,N_19994);
nor U21564 (N_21564,N_19680,N_16172);
xor U21565 (N_21565,N_18522,N_16437);
nand U21566 (N_21566,N_15858,N_18996);
nor U21567 (N_21567,N_15433,N_18097);
or U21568 (N_21568,N_15121,N_18251);
xnor U21569 (N_21569,N_17412,N_17361);
nand U21570 (N_21570,N_18039,N_18442);
or U21571 (N_21571,N_15626,N_17975);
xnor U21572 (N_21572,N_16033,N_19047);
nor U21573 (N_21573,N_15773,N_15094);
or U21574 (N_21574,N_19839,N_19334);
and U21575 (N_21575,N_15973,N_15436);
and U21576 (N_21576,N_15537,N_16998);
nand U21577 (N_21577,N_19352,N_16737);
or U21578 (N_21578,N_17477,N_15952);
and U21579 (N_21579,N_19285,N_15301);
and U21580 (N_21580,N_19609,N_15311);
or U21581 (N_21581,N_15716,N_17464);
xor U21582 (N_21582,N_18428,N_15622);
and U21583 (N_21583,N_15165,N_16680);
and U21584 (N_21584,N_19709,N_15882);
nor U21585 (N_21585,N_18954,N_19195);
or U21586 (N_21586,N_17378,N_18587);
nor U21587 (N_21587,N_17781,N_15382);
and U21588 (N_21588,N_15155,N_19562);
nor U21589 (N_21589,N_18586,N_19156);
nand U21590 (N_21590,N_18614,N_16386);
nand U21591 (N_21591,N_18682,N_18315);
or U21592 (N_21592,N_16691,N_16522);
nand U21593 (N_21593,N_15107,N_16537);
nand U21594 (N_21594,N_19466,N_15528);
nand U21595 (N_21595,N_15750,N_15527);
and U21596 (N_21596,N_19177,N_15278);
and U21597 (N_21597,N_16774,N_15374);
xor U21598 (N_21598,N_16267,N_18564);
and U21599 (N_21599,N_19900,N_18778);
nand U21600 (N_21600,N_18850,N_15946);
xor U21601 (N_21601,N_16030,N_16145);
nand U21602 (N_21602,N_15421,N_18553);
xor U21603 (N_21603,N_19714,N_19333);
xnor U21604 (N_21604,N_19707,N_19764);
nor U21605 (N_21605,N_17987,N_16466);
nor U21606 (N_21606,N_19299,N_15918);
nor U21607 (N_21607,N_17956,N_16101);
nor U21608 (N_21608,N_16922,N_17816);
nand U21609 (N_21609,N_15553,N_18511);
and U21610 (N_21610,N_19390,N_19668);
and U21611 (N_21611,N_16647,N_18050);
and U21612 (N_21612,N_16832,N_18736);
nand U21613 (N_21613,N_18717,N_15503);
xor U21614 (N_21614,N_19387,N_17546);
nor U21615 (N_21615,N_19109,N_16223);
or U21616 (N_21616,N_16526,N_17218);
and U21617 (N_21617,N_15083,N_16854);
and U21618 (N_21618,N_19507,N_19919);
or U21619 (N_21619,N_16434,N_17279);
nand U21620 (N_21620,N_17820,N_16345);
nand U21621 (N_21621,N_18683,N_19075);
nand U21622 (N_21622,N_15708,N_16427);
nand U21623 (N_21623,N_15774,N_19278);
and U21624 (N_21624,N_18502,N_18716);
and U21625 (N_21625,N_17712,N_19524);
and U21626 (N_21626,N_19465,N_15205);
nor U21627 (N_21627,N_19892,N_19023);
or U21628 (N_21628,N_15297,N_19567);
nand U21629 (N_21629,N_18810,N_16539);
nand U21630 (N_21630,N_19784,N_16866);
nor U21631 (N_21631,N_16446,N_15085);
nand U21632 (N_21632,N_18705,N_16400);
or U21633 (N_21633,N_19459,N_17478);
or U21634 (N_21634,N_17350,N_18201);
and U21635 (N_21635,N_19641,N_18436);
nand U21636 (N_21636,N_19074,N_18505);
nor U21637 (N_21637,N_15131,N_15331);
nand U21638 (N_21638,N_17072,N_17919);
xnor U21639 (N_21639,N_18266,N_16435);
nor U21640 (N_21640,N_19569,N_19350);
and U21641 (N_21641,N_15187,N_18552);
nand U21642 (N_21642,N_16587,N_16650);
nand U21643 (N_21643,N_16070,N_19549);
nor U21644 (N_21644,N_19629,N_17203);
and U21645 (N_21645,N_19209,N_15287);
xnor U21646 (N_21646,N_16426,N_16672);
nor U21647 (N_21647,N_15859,N_16260);
or U21648 (N_21648,N_18631,N_15852);
or U21649 (N_21649,N_19489,N_17155);
xor U21650 (N_21650,N_19576,N_15483);
and U21651 (N_21651,N_16521,N_19969);
nand U21652 (N_21652,N_18739,N_15937);
or U21653 (N_21653,N_17467,N_15662);
and U21654 (N_21654,N_17201,N_16197);
nand U21655 (N_21655,N_15814,N_17838);
or U21656 (N_21656,N_17685,N_17905);
nand U21657 (N_21657,N_15745,N_19201);
nand U21658 (N_21658,N_16954,N_17399);
and U21659 (N_21659,N_17016,N_19223);
nand U21660 (N_21660,N_18165,N_19407);
and U21661 (N_21661,N_15126,N_17009);
and U21662 (N_21662,N_17523,N_15670);
and U21663 (N_21663,N_16896,N_16433);
nand U21664 (N_21664,N_16734,N_17935);
nand U21665 (N_21665,N_18240,N_19870);
xnor U21666 (N_21666,N_18384,N_15482);
nand U21667 (N_21667,N_19531,N_17091);
nand U21668 (N_21668,N_16603,N_18571);
nor U21669 (N_21669,N_19929,N_19450);
xor U21670 (N_21670,N_18824,N_16219);
or U21671 (N_21671,N_15678,N_16042);
or U21672 (N_21672,N_19119,N_15308);
xnor U21673 (N_21673,N_18408,N_18945);
nor U21674 (N_21674,N_17824,N_15418);
nor U21675 (N_21675,N_18527,N_18888);
xnor U21676 (N_21676,N_16295,N_19901);
nor U21677 (N_21677,N_19760,N_19230);
nor U21678 (N_21678,N_17305,N_17045);
nand U21679 (N_21679,N_19420,N_18501);
or U21680 (N_21680,N_19903,N_19141);
and U21681 (N_21681,N_19004,N_15511);
xor U21682 (N_21682,N_19989,N_15261);
nor U21683 (N_21683,N_15054,N_17146);
nor U21684 (N_21684,N_19463,N_15776);
nor U21685 (N_21685,N_18223,N_19395);
nand U21686 (N_21686,N_17059,N_18999);
nor U21687 (N_21687,N_18265,N_19912);
nand U21688 (N_21688,N_16002,N_16785);
and U21689 (N_21689,N_19498,N_15393);
or U21690 (N_21690,N_18652,N_15425);
or U21691 (N_21691,N_15917,N_15460);
nand U21692 (N_21692,N_18017,N_15866);
nor U21693 (N_21693,N_18194,N_15294);
nand U21694 (N_21694,N_16237,N_16083);
nor U21695 (N_21695,N_15353,N_15945);
xor U21696 (N_21696,N_15339,N_18446);
nand U21697 (N_21697,N_16369,N_19242);
nor U21698 (N_21698,N_15019,N_19495);
nand U21699 (N_21699,N_16888,N_16569);
and U21700 (N_21700,N_17128,N_18222);
nor U21701 (N_21701,N_19490,N_16793);
nor U21702 (N_21702,N_16805,N_17209);
nor U21703 (N_21703,N_15665,N_19202);
nor U21704 (N_21704,N_15673,N_16353);
and U21705 (N_21705,N_17160,N_19582);
nor U21706 (N_21706,N_17921,N_19228);
or U21707 (N_21707,N_17691,N_15052);
nand U21708 (N_21708,N_16273,N_17813);
nor U21709 (N_21709,N_18022,N_17916);
nand U21710 (N_21710,N_16323,N_17026);
nand U21711 (N_21711,N_16903,N_18569);
or U21712 (N_21712,N_19573,N_17552);
nand U21713 (N_21713,N_16659,N_16346);
xnor U21714 (N_21714,N_17535,N_18292);
nor U21715 (N_21715,N_17448,N_17779);
nand U21716 (N_21716,N_18764,N_15396);
or U21717 (N_21717,N_19620,N_17429);
or U21718 (N_21718,N_15965,N_15727);
nor U21719 (N_21719,N_18495,N_16149);
nor U21720 (N_21720,N_18951,N_15012);
or U21721 (N_21721,N_15950,N_16863);
and U21722 (N_21722,N_17217,N_18817);
nor U21723 (N_21723,N_16192,N_15196);
nor U21724 (N_21724,N_17086,N_15454);
and U21725 (N_21725,N_17043,N_17300);
nor U21726 (N_21726,N_19806,N_19114);
xor U21727 (N_21727,N_17243,N_18256);
nand U21728 (N_21728,N_16383,N_19511);
nor U21729 (N_21729,N_19093,N_17874);
or U21730 (N_21730,N_17724,N_18700);
nand U21731 (N_21731,N_19591,N_15508);
nand U21732 (N_21732,N_18390,N_15612);
nand U21733 (N_21733,N_16483,N_16612);
nand U21734 (N_21734,N_16959,N_16822);
or U21735 (N_21735,N_19311,N_16332);
xnor U21736 (N_21736,N_19030,N_16309);
xor U21737 (N_21737,N_15669,N_17444);
or U21738 (N_21738,N_19774,N_17600);
and U21739 (N_21739,N_15616,N_17384);
nor U21740 (N_21740,N_18207,N_19337);
nor U21741 (N_21741,N_16238,N_15272);
or U21742 (N_21742,N_16259,N_15420);
nand U21743 (N_21743,N_18537,N_18628);
nor U21744 (N_21744,N_15162,N_16913);
or U21745 (N_21745,N_17376,N_19948);
nor U21746 (N_21746,N_17649,N_17426);
nor U21747 (N_21747,N_18002,N_17284);
nand U21748 (N_21748,N_15901,N_15028);
and U21749 (N_21749,N_16165,N_18727);
or U21750 (N_21750,N_18143,N_16623);
nor U21751 (N_21751,N_19738,N_15474);
nor U21752 (N_21752,N_15369,N_18591);
or U21753 (N_21753,N_15470,N_16756);
nor U21754 (N_21754,N_19196,N_19851);
nand U21755 (N_21755,N_16757,N_15687);
nand U21756 (N_21756,N_15222,N_18965);
or U21757 (N_21757,N_19197,N_17085);
nand U21758 (N_21758,N_17819,N_16644);
nand U21759 (N_21759,N_15087,N_18568);
nand U21760 (N_21760,N_16206,N_17002);
and U21761 (N_21761,N_18629,N_18672);
xnor U21762 (N_21762,N_18036,N_15943);
nor U21763 (N_21763,N_19953,N_17549);
nor U21764 (N_21764,N_18145,N_18353);
and U21765 (N_21765,N_17789,N_16608);
nor U21766 (N_21766,N_15766,N_15824);
nand U21767 (N_21767,N_17216,N_17285);
or U21768 (N_21768,N_18864,N_16892);
and U21769 (N_21769,N_16986,N_15557);
and U21770 (N_21770,N_18800,N_18014);
or U21771 (N_21771,N_16036,N_18886);
nor U21772 (N_21772,N_19659,N_16723);
xnor U21773 (N_21773,N_19247,N_19865);
and U21774 (N_21774,N_16551,N_16049);
nand U21775 (N_21775,N_19516,N_15177);
nor U21776 (N_21776,N_15898,N_19509);
nand U21777 (N_21777,N_17204,N_15034);
nor U21778 (N_21778,N_19264,N_16533);
and U21779 (N_21779,N_18422,N_15002);
nor U21780 (N_21780,N_17449,N_17330);
nand U21781 (N_21781,N_17406,N_16193);
nand U21782 (N_21782,N_19060,N_16726);
nor U21783 (N_21783,N_17358,N_18301);
nor U21784 (N_21784,N_19670,N_17191);
and U21785 (N_21785,N_16795,N_19388);
or U21786 (N_21786,N_17337,N_17342);
or U21787 (N_21787,N_18160,N_19150);
and U21788 (N_21788,N_17555,N_15079);
nand U21789 (N_21789,N_17760,N_17982);
or U21790 (N_21790,N_15156,N_15176);
xnor U21791 (N_21791,N_19376,N_15088);
xor U21792 (N_21792,N_19165,N_18375);
or U21793 (N_21793,N_17179,N_18643);
nand U21794 (N_21794,N_17386,N_16452);
nand U21795 (N_21795,N_18836,N_16486);
nand U21796 (N_21796,N_16142,N_19726);
nor U21797 (N_21797,N_15293,N_16045);
nand U21798 (N_21798,N_16005,N_18570);
nand U21799 (N_21799,N_19424,N_15462);
and U21800 (N_21800,N_18403,N_17018);
or U21801 (N_21801,N_17163,N_18087);
and U21802 (N_21802,N_19663,N_15831);
or U21803 (N_21803,N_18625,N_15755);
xor U21804 (N_21804,N_15231,N_16842);
nor U21805 (N_21805,N_19718,N_15962);
or U21806 (N_21806,N_18083,N_19523);
nand U21807 (N_21807,N_16950,N_18856);
or U21808 (N_21808,N_17309,N_16635);
or U21809 (N_21809,N_15108,N_17145);
and U21810 (N_21810,N_18608,N_17812);
and U21811 (N_21811,N_17036,N_19331);
nand U21812 (N_21812,N_19991,N_16456);
and U21813 (N_21813,N_17447,N_15736);
nand U21814 (N_21814,N_18181,N_15865);
and U21815 (N_21815,N_16764,N_17835);
or U21816 (N_21816,N_16717,N_16624);
or U21817 (N_21817,N_18746,N_19574);
or U21818 (N_21818,N_15927,N_17207);
nand U21819 (N_21819,N_16664,N_19823);
or U21820 (N_21820,N_17293,N_15657);
or U21821 (N_21821,N_17035,N_16213);
or U21822 (N_21822,N_17166,N_17120);
xor U21823 (N_21823,N_18776,N_16420);
nand U21824 (N_21824,N_15057,N_17801);
nand U21825 (N_21825,N_18584,N_17428);
nand U21826 (N_21826,N_15341,N_19819);
or U21827 (N_21827,N_17395,N_19876);
nand U21828 (N_21828,N_15601,N_15402);
nand U21829 (N_21829,N_19599,N_18865);
nor U21830 (N_21830,N_18755,N_18006);
nor U21831 (N_21831,N_17524,N_16351);
and U21832 (N_21832,N_17957,N_17791);
xnor U21833 (N_21833,N_19526,N_17985);
xnor U21834 (N_21834,N_15484,N_17846);
nand U21835 (N_21835,N_16766,N_18336);
or U21836 (N_21836,N_15816,N_16147);
xor U21837 (N_21837,N_17367,N_17056);
nor U21838 (N_21838,N_18334,N_15555);
or U21839 (N_21839,N_18340,N_18018);
or U21840 (N_21840,N_18622,N_17031);
nand U21841 (N_21841,N_15548,N_15014);
nor U21842 (N_21842,N_15032,N_16637);
and U21843 (N_21843,N_18474,N_19192);
or U21844 (N_21844,N_18494,N_16422);
or U21845 (N_21845,N_15158,N_16865);
and U21846 (N_21846,N_16781,N_18126);
and U21847 (N_21847,N_17375,N_17832);
and U21848 (N_21848,N_15837,N_15478);
xnor U21849 (N_21849,N_17023,N_15112);
and U21850 (N_21850,N_16419,N_15255);
or U21851 (N_21851,N_19754,N_15378);
nand U21852 (N_21852,N_16800,N_18450);
or U21853 (N_21853,N_16542,N_16847);
and U21854 (N_21854,N_19853,N_18899);
nor U21855 (N_21855,N_17933,N_16286);
nand U21856 (N_21856,N_16697,N_15783);
and U21857 (N_21857,N_15036,N_16710);
nand U21858 (N_21858,N_18358,N_19720);
or U21859 (N_21859,N_15174,N_16840);
and U21860 (N_21860,N_16804,N_16208);
nor U21861 (N_21861,N_15128,N_18801);
nand U21862 (N_21862,N_18600,N_16543);
nand U21863 (N_21863,N_15571,N_15432);
nor U21864 (N_21864,N_15440,N_17992);
and U21865 (N_21865,N_17470,N_17245);
and U21866 (N_21866,N_17410,N_17019);
or U21867 (N_21867,N_16413,N_19873);
or U21868 (N_21868,N_18076,N_15746);
or U21869 (N_21869,N_18150,N_17445);
and U21870 (N_21870,N_17177,N_15377);
nor U21871 (N_21871,N_15904,N_17438);
or U21872 (N_21872,N_19200,N_15718);
nor U21873 (N_21873,N_17088,N_15345);
nor U21874 (N_21874,N_19721,N_15610);
or U21875 (N_21875,N_18820,N_16886);
and U21876 (N_21876,N_19089,N_19478);
nand U21877 (N_21877,N_16683,N_18099);
nor U21878 (N_21878,N_15361,N_15066);
nor U21879 (N_21879,N_16321,N_19204);
nor U21880 (N_21880,N_19645,N_16152);
nor U21881 (N_21881,N_19785,N_15628);
nand U21882 (N_21882,N_17563,N_19500);
xnor U21883 (N_21883,N_17953,N_15823);
nor U21884 (N_21884,N_18812,N_19073);
xor U21885 (N_21885,N_16138,N_16673);
nor U21886 (N_21886,N_18543,N_19078);
and U21887 (N_21887,N_16464,N_16989);
nor U21888 (N_21888,N_18073,N_16161);
nor U21889 (N_21889,N_17267,N_15426);
nand U21890 (N_21890,N_18164,N_18448);
or U21891 (N_21891,N_17579,N_16350);
nor U21892 (N_21892,N_16718,N_19631);
nand U21893 (N_21893,N_15588,N_17198);
nor U21894 (N_21894,N_19982,N_18644);
or U21895 (N_21895,N_19472,N_16873);
or U21896 (N_21896,N_16915,N_18949);
nand U21897 (N_21897,N_15639,N_16463);
and U21898 (N_21898,N_15999,N_15617);
and U21899 (N_21899,N_18872,N_16600);
nor U21900 (N_21900,N_15658,N_16373);
nor U21901 (N_21901,N_16139,N_15166);
xnor U21902 (N_21902,N_19263,N_18786);
or U21903 (N_21903,N_15782,N_19922);
or U21904 (N_21904,N_16229,N_15729);
and U21905 (N_21905,N_18473,N_17532);
or U21906 (N_21906,N_18620,N_19217);
and U21907 (N_21907,N_15835,N_15747);
or U21908 (N_21908,N_15130,N_16506);
nand U21909 (N_21909,N_19221,N_18349);
or U21910 (N_21910,N_17596,N_19550);
xor U21911 (N_21911,N_15496,N_18112);
or U21912 (N_21912,N_17078,N_15191);
or U21913 (N_21913,N_17946,N_17083);
xnor U21914 (N_21914,N_18841,N_18706);
or U21915 (N_21915,N_19215,N_19627);
nand U21916 (N_21916,N_15929,N_16810);
nand U21917 (N_21917,N_16414,N_18862);
or U21918 (N_21918,N_18092,N_15568);
and U21919 (N_21919,N_15911,N_18063);
nand U21920 (N_21920,N_15912,N_19045);
nor U21921 (N_21921,N_15247,N_18378);
or U21922 (N_21922,N_17109,N_15758);
or U21923 (N_21923,N_15200,N_17842);
or U21924 (N_21924,N_17224,N_15017);
nand U21925 (N_21925,N_15812,N_17740);
xnor U21926 (N_21926,N_17336,N_18284);
nand U21927 (N_21927,N_17744,N_18892);
nor U21928 (N_21928,N_19545,N_15761);
or U21929 (N_21929,N_18995,N_16296);
or U21930 (N_21930,N_18689,N_19130);
or U21931 (N_21931,N_16905,N_16450);
nor U21932 (N_21932,N_17854,N_18406);
xnor U21933 (N_21933,N_17630,N_16568);
nand U21934 (N_21934,N_16548,N_19320);
nor U21935 (N_21935,N_19241,N_17533);
nand U21936 (N_21936,N_16920,N_18413);
nor U21937 (N_21937,N_16665,N_18352);
xnor U21938 (N_21938,N_19497,N_17037);
nor U21939 (N_21939,N_17173,N_18943);
nand U21940 (N_21940,N_16312,N_19983);
nand U21941 (N_21941,N_17955,N_17347);
and U21942 (N_21942,N_18582,N_15442);
or U21943 (N_21943,N_17765,N_18926);
and U21944 (N_21944,N_19920,N_18464);
nor U21945 (N_21945,N_18323,N_17783);
xnor U21946 (N_21946,N_15232,N_18922);
nand U21947 (N_21947,N_15792,N_19921);
or U21948 (N_21948,N_19667,N_19836);
nor U21949 (N_21949,N_19544,N_18575);
xnor U21950 (N_21950,N_16694,N_17242);
nor U21951 (N_21951,N_16210,N_19832);
and U21952 (N_21952,N_17005,N_16384);
or U21953 (N_21953,N_18319,N_16811);
and U21954 (N_21954,N_19214,N_16702);
or U21955 (N_21955,N_18105,N_15220);
nor U21956 (N_21956,N_19696,N_19220);
nand U21957 (N_21957,N_19037,N_19802);
nand U21958 (N_21958,N_16990,N_18743);
nor U21959 (N_21959,N_18674,N_16459);
nor U21960 (N_21960,N_15063,N_18558);
nor U21961 (N_21961,N_18254,N_17932);
xnor U21962 (N_21962,N_16728,N_19039);
nand U21963 (N_21963,N_15160,N_18211);
xnor U21964 (N_21964,N_19713,N_18549);
and U21965 (N_21965,N_15161,N_16853);
nor U21966 (N_21966,N_15499,N_16306);
nor U21967 (N_21967,N_16701,N_15455);
or U21968 (N_21968,N_17288,N_17794);
or U21969 (N_21969,N_15030,N_19692);
xor U21970 (N_21970,N_19283,N_16240);
xnor U21971 (N_21971,N_16609,N_16515);
and U21972 (N_21972,N_16669,N_16358);
and U21973 (N_21973,N_17936,N_15663);
and U21974 (N_21974,N_19056,N_17667);
xnor U21975 (N_21975,N_18594,N_17968);
nand U21976 (N_21976,N_17514,N_18379);
and U21977 (N_21977,N_17274,N_15215);
nand U21978 (N_21978,N_19896,N_19208);
nand U21979 (N_21979,N_16112,N_17491);
and U21980 (N_21980,N_18247,N_17713);
nand U21981 (N_21981,N_19303,N_18360);
nor U21982 (N_21982,N_16335,N_16516);
and U21983 (N_21983,N_15581,N_19971);
and U21984 (N_21984,N_15806,N_15693);
and U21985 (N_21985,N_17907,N_18059);
and U21986 (N_21986,N_16320,N_15249);
nand U21987 (N_21987,N_17773,N_16290);
nand U21988 (N_21988,N_15676,N_15633);
xnor U21989 (N_21989,N_18497,N_18250);
or U21990 (N_21990,N_19542,N_17081);
and U21991 (N_21991,N_18986,N_15569);
or U21992 (N_21992,N_16987,N_16141);
xnor U21993 (N_21993,N_15884,N_15961);
nor U21994 (N_21994,N_16348,N_15552);
nor U21995 (N_21995,N_15120,N_15563);
nand U21996 (N_21996,N_16660,N_17118);
nor U21997 (N_21997,N_15419,N_16761);
and U21998 (N_21998,N_17465,N_15146);
nor U21999 (N_21999,N_15010,N_15078);
nand U22000 (N_22000,N_18137,N_16183);
nand U22001 (N_22001,N_17150,N_16877);
and U22002 (N_22002,N_18415,N_17599);
or U22003 (N_22003,N_17354,N_17951);
or U22004 (N_22004,N_17032,N_15493);
nor U22005 (N_22005,N_16247,N_19640);
nand U22006 (N_22006,N_19224,N_16699);
and U22007 (N_22007,N_17186,N_16578);
and U22008 (N_22008,N_16546,N_19566);
nand U22009 (N_22009,N_17882,N_15064);
nand U22010 (N_22010,N_16808,N_17252);
nor U22011 (N_22011,N_15524,N_18082);
nand U22012 (N_22012,N_16517,N_19012);
xnor U22013 (N_22013,N_18236,N_16378);
and U22014 (N_22014,N_18889,N_16166);
nor U22015 (N_22015,N_18722,N_17656);
nand U22016 (N_22016,N_15951,N_19758);
and U22017 (N_22017,N_18317,N_15277);
or U22018 (N_22018,N_19002,N_18216);
or U22019 (N_22019,N_15631,N_15720);
and U22020 (N_22020,N_15069,N_19757);
nand U22021 (N_22021,N_19797,N_18368);
nor U22022 (N_22022,N_19062,N_15214);
or U22023 (N_22023,N_18487,N_15672);
nor U22024 (N_22024,N_17222,N_17053);
nand U22025 (N_22025,N_17521,N_17340);
nor U22026 (N_22026,N_16562,N_17282);
or U22027 (N_22027,N_15089,N_17721);
nand U22028 (N_22028,N_15467,N_19830);
or U22029 (N_22029,N_19583,N_17244);
nand U22030 (N_22030,N_18791,N_16798);
or U22031 (N_22031,N_15930,N_18267);
and U22032 (N_22032,N_15324,N_16576);
xor U22033 (N_22033,N_16638,N_16220);
or U22034 (N_22034,N_18096,N_19589);
or U22035 (N_22035,N_16750,N_17697);
nand U22036 (N_22036,N_16991,N_16682);
nor U22037 (N_22037,N_19985,N_18033);
and U22038 (N_22038,N_19158,N_17952);
nor U22039 (N_22039,N_19339,N_16164);
nand U22040 (N_22040,N_17833,N_15855);
nand U22041 (N_22041,N_15398,N_16979);
and U22042 (N_22042,N_18159,N_19706);
and U22043 (N_22043,N_15100,N_19938);
xnor U22044 (N_22044,N_16482,N_16500);
xnor U22045 (N_22045,N_17949,N_19962);
or U22046 (N_22046,N_17578,N_17678);
and U22047 (N_22047,N_17909,N_15756);
nand U22048 (N_22048,N_17313,N_17904);
or U22049 (N_22049,N_17694,N_15025);
or U22050 (N_22050,N_19733,N_17332);
and U22051 (N_22051,N_18056,N_19381);
nand U22052 (N_22052,N_18064,N_18598);
or U22053 (N_22053,N_18481,N_15502);
nand U22054 (N_22054,N_18262,N_19305);
nand U22055 (N_22055,N_16029,N_19429);
nand U22056 (N_22056,N_17137,N_16366);
nor U22057 (N_22057,N_17082,N_18361);
nand U22058 (N_22058,N_19115,N_16927);
and U22059 (N_22059,N_17930,N_17840);
xnor U22060 (N_22060,N_19258,N_18782);
or U22061 (N_22061,N_19775,N_15233);
nor U22062 (N_22062,N_16592,N_18028);
nor U22063 (N_22063,N_19309,N_17726);
nor U22064 (N_22064,N_18884,N_16971);
nor U22065 (N_22065,N_19194,N_16557);
nor U22066 (N_22066,N_16675,N_17635);
nor U22067 (N_22067,N_19147,N_19357);
and U22068 (N_22068,N_15072,N_19064);
or U22069 (N_22069,N_16347,N_16949);
nand U22070 (N_22070,N_17196,N_16653);
nor U22071 (N_22071,N_19968,N_19077);
nand U22072 (N_22072,N_16071,N_16221);
nor U22073 (N_22073,N_19136,N_15801);
nor U22074 (N_22074,N_15828,N_16231);
and U22075 (N_22075,N_18807,N_17021);
nor U22076 (N_22076,N_18293,N_19662);
and U22077 (N_22077,N_19685,N_15363);
and U22078 (N_22078,N_17024,N_19646);
or U22079 (N_22079,N_15412,N_19833);
nor U22080 (N_22080,N_17418,N_19173);
and U22081 (N_22081,N_18148,N_19274);
nor U22082 (N_22082,N_18149,N_15545);
nand U22083 (N_22083,N_15889,N_19096);
nand U22084 (N_22084,N_15125,N_15439);
and U22085 (N_22085,N_18667,N_17195);
nand U22086 (N_22086,N_19981,N_19729);
nand U22087 (N_22087,N_18777,N_19323);
xor U22088 (N_22088,N_15320,N_17623);
and U22089 (N_22089,N_16884,N_17880);
or U22090 (N_22090,N_16899,N_15787);
nand U22091 (N_22091,N_17893,N_16398);
or U22092 (N_22092,N_18069,N_17976);
nand U22093 (N_22093,N_19353,N_19448);
or U22094 (N_22094,N_19460,N_17359);
nor U22095 (N_22095,N_16468,N_16815);
or U22096 (N_22096,N_19986,N_17469);
nand U22097 (N_22097,N_18550,N_19171);
nand U22098 (N_22098,N_15757,N_18577);
and U22099 (N_22099,N_18341,N_19094);
nand U22100 (N_22100,N_16019,N_19193);
nand U22101 (N_22101,N_18231,N_15291);
and U22102 (N_22102,N_17861,N_15137);
or U22103 (N_22103,N_17800,N_16868);
xnor U22104 (N_22104,N_18459,N_15875);
nor U22105 (N_22105,N_17262,N_15095);
or U22106 (N_22106,N_16128,N_18034);
xor U22107 (N_22107,N_17328,N_15668);
nor U22108 (N_22108,N_15253,N_18011);
nand U22109 (N_22109,N_19555,N_16088);
nor U22110 (N_22110,N_17343,N_19533);
xor U22111 (N_22111,N_19963,N_17815);
and U22112 (N_22112,N_15538,N_19665);
nand U22113 (N_22113,N_17687,N_16266);
and U22114 (N_22114,N_16380,N_18767);
nand U22115 (N_22115,N_18027,N_17892);
nand U22116 (N_22116,N_15007,N_16487);
and U22117 (N_22117,N_16704,N_15000);
or U22118 (N_22118,N_16778,N_15295);
nor U22119 (N_22119,N_18268,N_18186);
nor U22120 (N_22120,N_18661,N_17334);
nor U22121 (N_22121,N_19051,N_15053);
or U22122 (N_22122,N_15075,N_15317);
and U22123 (N_22123,N_16421,N_15860);
or U22124 (N_22124,N_15642,N_17001);
or U22125 (N_22125,N_16668,N_17115);
and U22126 (N_22126,N_19406,N_18551);
or U22127 (N_22127,N_16155,N_15150);
nor U22128 (N_22128,N_19492,N_15283);
nand U22129 (N_22129,N_15491,N_15350);
or U22130 (N_22130,N_18121,N_15518);
nand U22131 (N_22131,N_19708,N_17881);
nor U22132 (N_22132,N_19354,N_19189);
nand U22133 (N_22133,N_18715,N_15394);
or U22134 (N_22134,N_19924,N_16536);
and U22135 (N_22135,N_18610,N_16354);
or U22136 (N_22136,N_18605,N_17637);
nand U22137 (N_22137,N_15872,N_16200);
nand U22138 (N_22138,N_18432,N_15071);
or U22139 (N_22139,N_18187,N_15654);
nand U22140 (N_22140,N_18840,N_17383);
xnor U22141 (N_22141,N_19290,N_15771);
or U22142 (N_22142,N_15611,N_15182);
and U22143 (N_22143,N_19710,N_17251);
nand U22144 (N_22144,N_18766,N_16839);
nor U22145 (N_22145,N_15888,N_16819);
nor U22146 (N_22146,N_18026,N_17499);
nand U22147 (N_22147,N_16646,N_18903);
or U22148 (N_22148,N_19906,N_17233);
nor U22149 (N_22149,N_15084,N_17462);
nand U22150 (N_22150,N_15695,N_16730);
nand U22151 (N_22151,N_15381,N_16105);
and U22152 (N_22152,N_19595,N_19072);
nor U22153 (N_22153,N_17466,N_15819);
nor U22154 (N_22154,N_17266,N_18151);
nand U22155 (N_22155,N_17158,N_15743);
and U22156 (N_22156,N_19762,N_17826);
xor U22157 (N_22157,N_15717,N_19124);
or U22158 (N_22158,N_15306,N_19952);
nor U22159 (N_22159,N_18060,N_16256);
or U22160 (N_22160,N_17870,N_17593);
nand U22161 (N_22161,N_18259,N_17719);
or U22162 (N_22162,N_19366,N_16203);
xor U22163 (N_22163,N_17855,N_19137);
and U22164 (N_22164,N_15791,N_15224);
or U22165 (N_22165,N_17432,N_18788);
xnor U22166 (N_22166,N_19577,N_15751);
nand U22167 (N_22167,N_18154,N_15645);
nor U22168 (N_22168,N_17541,N_16554);
nor U22169 (N_22169,N_18260,N_19525);
xor U22170 (N_22170,N_15685,N_19581);
xor U22171 (N_22171,N_17868,N_16878);
nor U22172 (N_22172,N_18431,N_19302);
or U22173 (N_22173,N_15805,N_17660);
and U22174 (N_22174,N_18846,N_19596);
and U22175 (N_22175,N_15005,N_18983);
nand U22176 (N_22176,N_15890,N_18433);
and U22177 (N_22177,N_18557,N_18929);
or U22178 (N_22178,N_19844,N_19805);
or U22179 (N_22179,N_19308,N_16162);
or U22180 (N_22180,N_19902,N_15157);
nand U22181 (N_22181,N_18796,N_18708);
nand U22182 (N_22182,N_17864,N_18455);
nor U22183 (N_22183,N_17333,N_15599);
and U22184 (N_22184,N_15029,N_18003);
or U22185 (N_22185,N_16679,N_19187);
xor U22186 (N_22186,N_17190,N_19121);
nand U22187 (N_22187,N_17510,N_16719);
or U22188 (N_22188,N_18016,N_18563);
or U22189 (N_22189,N_16034,N_19992);
nand U22190 (N_22190,N_18041,N_18719);
and U22191 (N_22191,N_18346,N_19386);
or U22192 (N_22192,N_16921,N_18342);
nand U22193 (N_22193,N_16117,N_16995);
nor U22194 (N_22194,N_18685,N_17226);
and U22195 (N_22195,N_17090,N_18763);
or U22196 (N_22196,N_16248,N_19730);
or U22197 (N_22197,N_16059,N_17220);
nand U22198 (N_22198,N_19212,N_17063);
nor U22199 (N_22199,N_15817,N_19910);
xnor U22200 (N_22200,N_18098,N_17489);
or U22201 (N_22201,N_18816,N_18219);
nor U22202 (N_22202,N_16696,N_15597);
xor U22203 (N_22203,N_18939,N_16641);
nor U22204 (N_22204,N_18466,N_19539);
and U22205 (N_22205,N_18067,N_17906);
and U22206 (N_22206,N_17729,N_18179);
nor U22207 (N_22207,N_18373,N_15504);
or U22208 (N_22208,N_17390,N_19723);
nor U22209 (N_22209,N_18616,N_16265);
nand U22210 (N_22210,N_19613,N_17990);
nand U22211 (N_22211,N_16825,N_16262);
and U22212 (N_22212,N_18925,N_19559);
nor U22213 (N_22213,N_16061,N_17594);
and U22214 (N_22214,N_16089,N_18344);
nor U22215 (N_22215,N_17437,N_17924);
nand U22216 (N_22216,N_18214,N_18825);
or U22217 (N_22217,N_18399,N_15802);
or U22218 (N_22218,N_18423,N_15313);
nor U22219 (N_22219,N_17094,N_19091);
and U22220 (N_22220,N_17584,N_18300);
and U22221 (N_22221,N_16773,N_17248);
and U22222 (N_22222,N_16314,N_19689);
or U22223 (N_22223,N_17382,N_17970);
xor U22224 (N_22224,N_15406,N_16444);
xnor U22225 (N_22225,N_15274,N_18217);
nor U22226 (N_22226,N_17034,N_16944);
or U22227 (N_22227,N_18439,N_18425);
nor U22228 (N_22228,N_16559,N_15309);
nand U22229 (N_22229,N_17914,N_15038);
and U22230 (N_22230,N_17927,N_16883);
nand U22231 (N_22231,N_15061,N_17735);
and U22232 (N_22232,N_17790,N_17239);
and U22233 (N_22233,N_19178,N_15887);
and U22234 (N_22234,N_19530,N_15996);
nor U22235 (N_22235,N_19166,N_18588);
nor U22236 (N_22236,N_19438,N_18887);
or U22237 (N_22237,N_16831,N_15209);
nand U22238 (N_22238,N_18230,N_15411);
or U22239 (N_22239,N_19132,N_15206);
nand U22240 (N_22240,N_15550,N_15649);
or U22241 (N_22241,N_16032,N_19881);
nor U22242 (N_22242,N_19099,N_19503);
nor U22243 (N_22243,N_18470,N_18363);
nor U22244 (N_22244,N_17585,N_15958);
nor U22245 (N_22245,N_15878,N_17277);
nand U22246 (N_22246,N_19917,N_19705);
xor U22247 (N_22247,N_16689,N_16188);
nand U22248 (N_22248,N_16513,N_19804);
and U22249 (N_22249,N_19557,N_17008);
or U22250 (N_22250,N_19601,N_15796);
xor U22251 (N_22251,N_15712,N_15533);
or U22252 (N_22252,N_18488,N_19913);
or U22253 (N_22253,N_15680,N_15620);
and U22254 (N_22254,N_16484,N_16226);
or U22255 (N_22255,N_17028,N_15023);
nor U22256 (N_22256,N_18127,N_17827);
and U22257 (N_22257,N_18238,N_15009);
nand U22258 (N_22258,N_16510,N_17604);
or U22259 (N_22259,N_18212,N_17392);
or U22260 (N_22260,N_16118,N_15903);
and U22261 (N_22261,N_18177,N_15964);
nor U22262 (N_22262,N_15646,N_17841);
nor U22263 (N_22263,N_19810,N_15786);
and U22264 (N_22264,N_15376,N_17887);
nor U22265 (N_22265,N_17442,N_16412);
nand U22266 (N_22266,N_16357,N_17998);
and U22267 (N_22267,N_17822,N_18224);
nand U22268 (N_22268,N_16253,N_15803);
nand U22269 (N_22269,N_17944,N_17672);
nand U22270 (N_22270,N_18993,N_19292);
nor U22271 (N_22271,N_18596,N_18065);
and U22272 (N_22272,N_17603,N_15248);
nand U22273 (N_22273,N_17758,N_16662);
nor U22274 (N_22274,N_15551,N_15981);
nand U22275 (N_22275,N_17891,N_17915);
nor U22276 (N_22276,N_15430,N_17335);
nand U22277 (N_22277,N_18282,N_18114);
or U22278 (N_22278,N_16401,N_19061);
nand U22279 (N_22279,N_17054,N_15207);
and U22280 (N_22280,N_18998,N_16695);
or U22281 (N_22281,N_15106,N_15624);
nor U22282 (N_22282,N_16129,N_19413);
and U22283 (N_22283,N_17894,N_16820);
xnor U22284 (N_22284,N_16985,N_19790);
nand U22285 (N_22285,N_17548,N_19964);
nor U22286 (N_22286,N_18460,N_17405);
nand U22287 (N_22287,N_18037,N_16970);
nand U22288 (N_22288,N_15111,N_16573);
xnor U22289 (N_22289,N_16143,N_19658);
nand U22290 (N_22290,N_16969,N_17814);
or U22291 (N_22291,N_19416,N_17737);
and U22292 (N_22292,N_18419,N_17869);
or U22293 (N_22293,N_19427,N_19877);
and U22294 (N_22294,N_15145,N_16479);
or U22295 (N_22295,N_16363,N_16821);
nor U22296 (N_22296,N_19364,N_18768);
xor U22297 (N_22297,N_17079,N_15618);
and U22298 (N_22298,N_18205,N_17530);
nand U22299 (N_22299,N_17456,N_15098);
and U22300 (N_22300,N_16093,N_17948);
or U22301 (N_22301,N_16214,N_16956);
nor U22302 (N_22302,N_15164,N_18400);
or U22303 (N_22303,N_16387,N_18035);
and U22304 (N_22304,N_17730,N_17314);
and U22305 (N_22305,N_17960,N_19840);
nor U22306 (N_22306,N_16334,N_19005);
nand U22307 (N_22307,N_16402,N_19958);
and U22308 (N_22308,N_17261,N_15594);
and U22309 (N_22309,N_17495,N_16591);
nor U22310 (N_22310,N_17488,N_15711);
or U22311 (N_22311,N_16333,N_18960);
nand U22312 (N_22312,N_15485,N_17728);
nor U22313 (N_22313,N_16677,N_19085);
xor U22314 (N_22314,N_15940,N_15739);
nor U22315 (N_22315,N_19693,N_17468);
or U22316 (N_22316,N_17071,N_18997);
and U22317 (N_22317,N_18515,N_19657);
and U22318 (N_22318,N_19995,N_17939);
nor U22319 (N_22319,N_19341,N_19878);
nand U22320 (N_22320,N_18133,N_16532);
or U22321 (N_22321,N_18572,N_15741);
nor U22322 (N_22322,N_18178,N_15715);
nor U22323 (N_22323,N_19765,N_17188);
nor U22324 (N_22324,N_18278,N_19360);
nor U22325 (N_22325,N_19796,N_16527);
nor U22326 (N_22326,N_18209,N_18321);
xor U22327 (N_22327,N_19777,N_19622);
nand U22328 (N_22328,N_18144,N_19286);
nand U22329 (N_22329,N_17474,N_16893);
xor U22330 (N_22330,N_15788,N_17945);
nand U22331 (N_22331,N_16167,N_18401);
nand U22332 (N_22332,N_19205,N_17182);
and U22333 (N_22333,N_18469,N_19180);
and U22334 (N_22334,N_19588,N_16787);
and U22335 (N_22335,N_16254,N_15590);
or U22336 (N_22336,N_17276,N_19252);
nand U22337 (N_22337,N_19621,N_16371);
nor U22338 (N_22338,N_18624,N_17853);
nand U22339 (N_22339,N_17119,N_16817);
xnor U22340 (N_22340,N_16242,N_17734);
or U22341 (N_22341,N_17303,N_15438);
nor U22342 (N_22342,N_19905,N_18462);
nor U22343 (N_22343,N_18516,N_18338);
and U22344 (N_22344,N_19828,N_17046);
nor U22345 (N_22345,N_15302,N_19315);
and U22346 (N_22346,N_19512,N_15351);
or U22347 (N_22347,N_18520,N_16388);
nor U22348 (N_22348,N_15517,N_17979);
nand U22349 (N_22349,N_16741,N_18024);
nand U22350 (N_22350,N_18933,N_18656);
or U22351 (N_22351,N_18784,N_15906);
or U22352 (N_22352,N_16941,N_17041);
or U22353 (N_22353,N_15316,N_16876);
and U22354 (N_22354,N_16391,N_16700);
or U22355 (N_22355,N_16655,N_15573);
and U22356 (N_22356,N_17055,N_16448);
or U22357 (N_22357,N_17051,N_19845);
nand U22358 (N_22358,N_16933,N_17272);
or U22359 (N_22359,N_16330,N_18008);
nor U22360 (N_22360,N_19014,N_15861);
nand U22361 (N_22361,N_17676,N_18524);
and U22362 (N_22362,N_19373,N_16550);
and U22363 (N_22363,N_18329,N_16681);
or U22364 (N_22364,N_15151,N_17828);
or U22365 (N_22365,N_17663,N_15129);
or U22366 (N_22366,N_15186,N_19846);
or U22367 (N_22367,N_17025,N_19295);
nor U22368 (N_22368,N_18809,N_16931);
or U22369 (N_22369,N_15268,N_19907);
and U22370 (N_22370,N_16794,N_18314);
nand U22371 (N_22371,N_19560,N_18891);
and U22372 (N_22372,N_19553,N_17601);
nand U22373 (N_22373,N_19249,N_15021);
nand U22374 (N_22374,N_18161,N_17845);
or U22375 (N_22375,N_17654,N_18618);
and U22376 (N_22376,N_19529,N_17211);
or U22377 (N_22377,N_18666,N_17162);
nor U22378 (N_22378,N_17294,N_15045);
or U22379 (N_22379,N_15346,N_17692);
or U22380 (N_22380,N_17507,N_16946);
nand U22381 (N_22381,N_17296,N_19711);
and U22382 (N_22382,N_16846,N_16759);
xor U22383 (N_22383,N_16255,N_15540);
nor U22384 (N_22384,N_17065,N_15874);
xnor U22385 (N_22385,N_15558,N_17885);
nand U22386 (N_22386,N_17923,N_17144);
nand U22387 (N_22387,N_15469,N_19722);
or U22388 (N_22388,N_18613,N_17231);
nor U22389 (N_22389,N_18276,N_18463);
and U22390 (N_22390,N_18805,N_15319);
nand U22391 (N_22391,N_19348,N_19458);
xnor U22392 (N_22392,N_18528,N_16339);
and U22393 (N_22393,N_15475,N_18245);
xnor U22394 (N_22394,N_19453,N_17000);
and U22395 (N_22395,N_16887,N_18174);
or U22396 (N_22396,N_17598,N_17795);
xor U22397 (N_22397,N_15315,N_15863);
nand U22398 (N_22398,N_15349,N_17401);
and U22399 (N_22399,N_15976,N_19961);
nor U22400 (N_22400,N_18252,N_17908);
nor U22401 (N_22401,N_18157,N_18711);
or U22402 (N_22402,N_15510,N_15201);
nand U22403 (N_22403,N_19277,N_17070);
nor U22404 (N_22404,N_17547,N_16851);
nand U22405 (N_22405,N_16593,N_15799);
and U22406 (N_22406,N_16488,N_18163);
nor U22407 (N_22407,N_15724,N_15694);
or U22408 (N_22408,N_15006,N_18304);
xnor U22409 (N_22409,N_15035,N_19947);
or U22410 (N_22410,N_19298,N_16150);
and U22411 (N_22411,N_18944,N_18213);
and U22412 (N_22412,N_16471,N_18438);
nand U22413 (N_22413,N_15560,N_15702);
nor U22414 (N_22414,N_15238,N_19623);
or U22415 (N_22415,N_16807,N_18441);
or U22416 (N_22416,N_18532,N_17610);
or U22417 (N_22417,N_19698,N_17125);
nor U22418 (N_22418,N_17500,N_16039);
nand U22419 (N_22419,N_18020,N_16425);
nor U22420 (N_22420,N_18395,N_17784);
nor U22421 (N_22421,N_15332,N_19245);
and U22422 (N_22422,N_19281,N_19946);
nor U22423 (N_22423,N_19626,N_18512);
nor U22424 (N_22424,N_19918,N_18015);
xor U22425 (N_22425,N_18540,N_19229);
or U22426 (N_22426,N_16497,N_17651);
xnor U22427 (N_22427,N_16394,N_19127);
nor U22428 (N_22428,N_18530,N_17396);
and U22429 (N_22429,N_18818,N_19632);
and U22430 (N_22430,N_16454,N_17238);
or U22431 (N_22431,N_17295,N_15947);
and U22432 (N_22432,N_16191,N_18911);
and U22433 (N_22433,N_18765,N_18556);
nor U22434 (N_22434,N_15173,N_18576);
and U22435 (N_22435,N_16676,N_16978);
and U22436 (N_22436,N_18980,N_15881);
nor U22437 (N_22437,N_18381,N_15105);
and U22438 (N_22438,N_17926,N_18427);
nor U22439 (N_22439,N_19935,N_17013);
and U22440 (N_22440,N_18590,N_15304);
nand U22441 (N_22441,N_19614,N_15575);
nor U22442 (N_22442,N_15219,N_18458);
nor U22443 (N_22443,N_15603,N_18921);
and U22444 (N_22444,N_16556,N_18091);
nand U22445 (N_22445,N_19617,N_19493);
nand U22446 (N_22446,N_17197,N_16194);
nand U22447 (N_22447,N_16553,N_17321);
or U22448 (N_22448,N_17922,N_19554);
and U22449 (N_22449,N_16731,N_17066);
or U22450 (N_22450,N_19182,N_19869);
and U22451 (N_22451,N_17877,N_16035);
nand U22452 (N_22452,N_15554,N_19578);
or U22453 (N_22453,N_19619,N_19502);
nor U22454 (N_22454,N_19125,N_16407);
nor U22455 (N_22455,N_18156,N_18710);
and U22456 (N_22456,N_18623,N_18696);
or U22457 (N_22457,N_19006,N_17559);
or U22458 (N_22458,N_18518,N_19203);
and U22459 (N_22459,N_18206,N_19941);
nand U22460 (N_22460,N_16754,N_19630);
nand U22461 (N_22461,N_18009,N_16534);
and U22462 (N_22462,N_19411,N_19327);
nand U22463 (N_22463,N_17490,N_17360);
or U22464 (N_22464,N_19269,N_18348);
nor U22465 (N_22465,N_17829,N_16075);
or U22466 (N_22466,N_18389,N_19829);
and U22467 (N_22467,N_19414,N_16018);
nor U22468 (N_22468,N_19974,N_16028);
or U22469 (N_22469,N_19999,N_19856);
nor U22470 (N_22470,N_19324,N_16300);
xnor U22471 (N_22471,N_19972,N_18234);
or U22472 (N_22472,N_19703,N_16298);
or U22473 (N_22473,N_17187,N_16507);
and U22474 (N_22474,N_18482,N_19435);
nand U22475 (N_22475,N_17659,N_19449);
nand U22476 (N_22476,N_16186,N_15172);
nand U22477 (N_22477,N_19688,N_16870);
or U22478 (N_22478,N_18792,N_17497);
nand U22479 (N_22479,N_18724,N_16535);
nand U22480 (N_22480,N_17895,N_18835);
and U22481 (N_22481,N_16449,N_16250);
xor U22482 (N_22482,N_19814,N_17543);
nor U22483 (N_22483,N_17741,N_19813);
and U22484 (N_22484,N_15322,N_15506);
or U22485 (N_22485,N_19359,N_18061);
or U22486 (N_22486,N_17286,N_18215);
or U22487 (N_22487,N_19410,N_16642);
nand U22488 (N_22488,N_17391,N_19385);
or U22489 (N_22489,N_16125,N_17129);
nor U22490 (N_22490,N_18787,N_18869);
nand U22491 (N_22491,N_19279,N_19633);
nor U22492 (N_22492,N_19389,N_17808);
nand U22493 (N_22493,N_19160,N_16514);
xnor U22494 (N_22494,N_17934,N_18115);
nor U22495 (N_22495,N_15392,N_18337);
or U22496 (N_22496,N_15110,N_15413);
nand U22497 (N_22497,N_18684,N_19041);
or U22498 (N_22498,N_17950,N_17010);
and U22499 (N_22499,N_17178,N_16085);
and U22500 (N_22500,N_17683,N_18872);
nand U22501 (N_22501,N_17900,N_17896);
nor U22502 (N_22502,N_19939,N_15856);
nand U22503 (N_22503,N_17424,N_15554);
nor U22504 (N_22504,N_19584,N_16507);
or U22505 (N_22505,N_18675,N_15080);
nand U22506 (N_22506,N_18516,N_18875);
nor U22507 (N_22507,N_15226,N_17191);
xnor U22508 (N_22508,N_17623,N_18592);
and U22509 (N_22509,N_19761,N_16444);
or U22510 (N_22510,N_15121,N_15534);
or U22511 (N_22511,N_19921,N_16660);
xnor U22512 (N_22512,N_15340,N_18135);
and U22513 (N_22513,N_19908,N_15926);
and U22514 (N_22514,N_15151,N_17545);
nand U22515 (N_22515,N_17910,N_17137);
and U22516 (N_22516,N_17537,N_18260);
xnor U22517 (N_22517,N_15992,N_15098);
nor U22518 (N_22518,N_19665,N_18102);
nor U22519 (N_22519,N_17650,N_15199);
xnor U22520 (N_22520,N_19132,N_19804);
or U22521 (N_22521,N_18369,N_19315);
nor U22522 (N_22522,N_17022,N_15651);
and U22523 (N_22523,N_17281,N_19127);
nor U22524 (N_22524,N_17146,N_15824);
nor U22525 (N_22525,N_16782,N_18982);
or U22526 (N_22526,N_17261,N_15872);
nand U22527 (N_22527,N_16278,N_19887);
and U22528 (N_22528,N_16380,N_16327);
or U22529 (N_22529,N_16241,N_18837);
nand U22530 (N_22530,N_15841,N_19460);
or U22531 (N_22531,N_19985,N_15450);
and U22532 (N_22532,N_16830,N_17663);
nand U22533 (N_22533,N_15718,N_19397);
or U22534 (N_22534,N_16532,N_16849);
nor U22535 (N_22535,N_15935,N_19856);
or U22536 (N_22536,N_17155,N_19397);
nand U22537 (N_22537,N_19365,N_16069);
nor U22538 (N_22538,N_18548,N_18362);
and U22539 (N_22539,N_16920,N_19940);
nand U22540 (N_22540,N_19435,N_17226);
and U22541 (N_22541,N_15324,N_19050);
nor U22542 (N_22542,N_18163,N_15861);
and U22543 (N_22543,N_15786,N_15612);
and U22544 (N_22544,N_18489,N_16090);
or U22545 (N_22545,N_17156,N_15578);
or U22546 (N_22546,N_18484,N_18525);
or U22547 (N_22547,N_19738,N_19665);
or U22548 (N_22548,N_16407,N_16840);
nor U22549 (N_22549,N_18157,N_19255);
and U22550 (N_22550,N_15554,N_16152);
nand U22551 (N_22551,N_18541,N_19185);
nor U22552 (N_22552,N_18469,N_16023);
and U22553 (N_22553,N_18145,N_15529);
or U22554 (N_22554,N_17083,N_15980);
nand U22555 (N_22555,N_19275,N_19782);
nor U22556 (N_22556,N_19176,N_16539);
nor U22557 (N_22557,N_16523,N_15260);
and U22558 (N_22558,N_19849,N_18761);
nand U22559 (N_22559,N_18703,N_17896);
nand U22560 (N_22560,N_18370,N_15479);
nand U22561 (N_22561,N_18034,N_16400);
or U22562 (N_22562,N_15079,N_19358);
and U22563 (N_22563,N_15513,N_19447);
nor U22564 (N_22564,N_19039,N_19911);
nand U22565 (N_22565,N_15737,N_16818);
and U22566 (N_22566,N_15416,N_18718);
and U22567 (N_22567,N_18393,N_15155);
or U22568 (N_22568,N_18499,N_15944);
and U22569 (N_22569,N_16484,N_16137);
nand U22570 (N_22570,N_17878,N_16727);
nand U22571 (N_22571,N_16095,N_19104);
nor U22572 (N_22572,N_19592,N_15124);
and U22573 (N_22573,N_16912,N_15347);
or U22574 (N_22574,N_16661,N_17863);
nand U22575 (N_22575,N_15698,N_18308);
nand U22576 (N_22576,N_15923,N_19354);
nor U22577 (N_22577,N_16950,N_18258);
xnor U22578 (N_22578,N_17926,N_15748);
and U22579 (N_22579,N_18760,N_16281);
nor U22580 (N_22580,N_19282,N_19692);
nor U22581 (N_22581,N_19355,N_17281);
or U22582 (N_22582,N_16321,N_15633);
or U22583 (N_22583,N_18799,N_17172);
or U22584 (N_22584,N_17058,N_18215);
and U22585 (N_22585,N_15827,N_16676);
nand U22586 (N_22586,N_17308,N_15334);
nor U22587 (N_22587,N_17271,N_17822);
or U22588 (N_22588,N_16259,N_18384);
and U22589 (N_22589,N_18214,N_18846);
nor U22590 (N_22590,N_18569,N_15942);
nand U22591 (N_22591,N_19823,N_17858);
nor U22592 (N_22592,N_15487,N_18967);
and U22593 (N_22593,N_15902,N_17290);
nor U22594 (N_22594,N_19159,N_18659);
and U22595 (N_22595,N_19887,N_19322);
nor U22596 (N_22596,N_15043,N_15164);
nand U22597 (N_22597,N_16760,N_17716);
or U22598 (N_22598,N_19657,N_18257);
nand U22599 (N_22599,N_18257,N_16454);
xnor U22600 (N_22600,N_19476,N_15940);
and U22601 (N_22601,N_18161,N_16264);
xor U22602 (N_22602,N_16052,N_16352);
nand U22603 (N_22603,N_16777,N_15967);
nor U22604 (N_22604,N_18617,N_17301);
and U22605 (N_22605,N_15543,N_17763);
or U22606 (N_22606,N_19784,N_16006);
and U22607 (N_22607,N_19455,N_19545);
nor U22608 (N_22608,N_19037,N_16954);
nand U22609 (N_22609,N_17887,N_19664);
nand U22610 (N_22610,N_18730,N_18218);
nand U22611 (N_22611,N_16378,N_17694);
nand U22612 (N_22612,N_17616,N_15239);
nor U22613 (N_22613,N_19218,N_15787);
xnor U22614 (N_22614,N_18214,N_17675);
nand U22615 (N_22615,N_17099,N_16815);
nand U22616 (N_22616,N_17903,N_17534);
or U22617 (N_22617,N_19480,N_16531);
nor U22618 (N_22618,N_19737,N_19198);
nor U22619 (N_22619,N_17711,N_19643);
and U22620 (N_22620,N_17155,N_19920);
nor U22621 (N_22621,N_19451,N_15427);
nand U22622 (N_22622,N_16085,N_18521);
nand U22623 (N_22623,N_19068,N_19781);
or U22624 (N_22624,N_16595,N_17389);
and U22625 (N_22625,N_19753,N_18989);
nand U22626 (N_22626,N_18516,N_16785);
nand U22627 (N_22627,N_19545,N_18628);
or U22628 (N_22628,N_18040,N_15285);
or U22629 (N_22629,N_19687,N_17614);
or U22630 (N_22630,N_15073,N_15691);
or U22631 (N_22631,N_19878,N_19591);
or U22632 (N_22632,N_15895,N_17602);
or U22633 (N_22633,N_17204,N_18012);
and U22634 (N_22634,N_19674,N_19207);
and U22635 (N_22635,N_16844,N_17622);
nor U22636 (N_22636,N_17353,N_16346);
or U22637 (N_22637,N_15139,N_16027);
or U22638 (N_22638,N_18285,N_18418);
and U22639 (N_22639,N_18820,N_15947);
and U22640 (N_22640,N_17934,N_18991);
nand U22641 (N_22641,N_17616,N_18626);
nand U22642 (N_22642,N_18478,N_19040);
and U22643 (N_22643,N_17729,N_16828);
nand U22644 (N_22644,N_17996,N_17042);
nand U22645 (N_22645,N_19815,N_16025);
and U22646 (N_22646,N_17770,N_18266);
nand U22647 (N_22647,N_15175,N_19610);
nand U22648 (N_22648,N_16641,N_15915);
nand U22649 (N_22649,N_17887,N_15937);
nand U22650 (N_22650,N_19896,N_16868);
and U22651 (N_22651,N_16623,N_15697);
or U22652 (N_22652,N_18708,N_17786);
nor U22653 (N_22653,N_19807,N_17333);
xnor U22654 (N_22654,N_17236,N_19155);
and U22655 (N_22655,N_18340,N_15301);
nor U22656 (N_22656,N_18282,N_16663);
and U22657 (N_22657,N_19179,N_18900);
nor U22658 (N_22658,N_19009,N_15756);
and U22659 (N_22659,N_17425,N_18356);
and U22660 (N_22660,N_19405,N_16549);
nand U22661 (N_22661,N_15976,N_15213);
nor U22662 (N_22662,N_15925,N_15086);
xnor U22663 (N_22663,N_15103,N_18809);
and U22664 (N_22664,N_19148,N_16378);
and U22665 (N_22665,N_15529,N_15451);
or U22666 (N_22666,N_16049,N_17179);
nand U22667 (N_22667,N_18737,N_15605);
nand U22668 (N_22668,N_17622,N_17836);
and U22669 (N_22669,N_19058,N_16211);
or U22670 (N_22670,N_16374,N_16063);
nand U22671 (N_22671,N_16353,N_15316);
and U22672 (N_22672,N_17611,N_17381);
and U22673 (N_22673,N_18159,N_17821);
and U22674 (N_22674,N_18863,N_18803);
xor U22675 (N_22675,N_15692,N_18638);
xnor U22676 (N_22676,N_15959,N_19843);
nor U22677 (N_22677,N_16069,N_15219);
and U22678 (N_22678,N_17236,N_18295);
and U22679 (N_22679,N_17539,N_18892);
nand U22680 (N_22680,N_18145,N_16621);
and U22681 (N_22681,N_17648,N_15670);
nand U22682 (N_22682,N_16071,N_18536);
nor U22683 (N_22683,N_19891,N_16757);
nand U22684 (N_22684,N_18266,N_18093);
nand U22685 (N_22685,N_16308,N_19773);
nor U22686 (N_22686,N_17955,N_15892);
or U22687 (N_22687,N_19196,N_17763);
or U22688 (N_22688,N_15243,N_16502);
or U22689 (N_22689,N_17032,N_18612);
nand U22690 (N_22690,N_17396,N_15376);
nand U22691 (N_22691,N_19559,N_18044);
nor U22692 (N_22692,N_17292,N_15373);
and U22693 (N_22693,N_17806,N_18099);
xor U22694 (N_22694,N_17720,N_17558);
xnor U22695 (N_22695,N_18140,N_16405);
nor U22696 (N_22696,N_17949,N_17861);
and U22697 (N_22697,N_19155,N_19592);
nand U22698 (N_22698,N_16907,N_15695);
and U22699 (N_22699,N_16026,N_18706);
nor U22700 (N_22700,N_17253,N_15420);
or U22701 (N_22701,N_16267,N_19793);
xnor U22702 (N_22702,N_16582,N_19371);
nor U22703 (N_22703,N_16057,N_19265);
and U22704 (N_22704,N_15882,N_16945);
nor U22705 (N_22705,N_15163,N_19379);
and U22706 (N_22706,N_17792,N_18813);
xor U22707 (N_22707,N_16267,N_16271);
nor U22708 (N_22708,N_18721,N_18411);
nor U22709 (N_22709,N_19131,N_17559);
xor U22710 (N_22710,N_18685,N_18956);
and U22711 (N_22711,N_17739,N_16780);
nor U22712 (N_22712,N_18405,N_15496);
nor U22713 (N_22713,N_16123,N_19940);
nor U22714 (N_22714,N_15891,N_17952);
or U22715 (N_22715,N_17339,N_18477);
xnor U22716 (N_22716,N_17027,N_15043);
and U22717 (N_22717,N_18663,N_19706);
nand U22718 (N_22718,N_15633,N_18203);
nand U22719 (N_22719,N_19566,N_18176);
nor U22720 (N_22720,N_19783,N_15110);
nand U22721 (N_22721,N_18962,N_17544);
nand U22722 (N_22722,N_17257,N_19486);
or U22723 (N_22723,N_16309,N_17952);
or U22724 (N_22724,N_19026,N_18817);
nor U22725 (N_22725,N_16710,N_15604);
nand U22726 (N_22726,N_17235,N_19611);
and U22727 (N_22727,N_18137,N_18241);
xnor U22728 (N_22728,N_15792,N_16958);
nand U22729 (N_22729,N_15508,N_15686);
nand U22730 (N_22730,N_17744,N_16141);
xor U22731 (N_22731,N_16888,N_18071);
nor U22732 (N_22732,N_16418,N_17072);
xor U22733 (N_22733,N_19285,N_17654);
or U22734 (N_22734,N_17793,N_19669);
or U22735 (N_22735,N_15377,N_15304);
and U22736 (N_22736,N_17987,N_18063);
nand U22737 (N_22737,N_16430,N_15719);
nor U22738 (N_22738,N_18078,N_19100);
nor U22739 (N_22739,N_15547,N_16656);
and U22740 (N_22740,N_17766,N_18674);
nand U22741 (N_22741,N_19002,N_17435);
xor U22742 (N_22742,N_18349,N_19162);
or U22743 (N_22743,N_16596,N_19921);
nand U22744 (N_22744,N_16633,N_19627);
xor U22745 (N_22745,N_19115,N_17232);
and U22746 (N_22746,N_15022,N_16102);
nor U22747 (N_22747,N_15971,N_19786);
or U22748 (N_22748,N_15851,N_19089);
nor U22749 (N_22749,N_18657,N_17413);
and U22750 (N_22750,N_16833,N_19988);
nor U22751 (N_22751,N_19392,N_19501);
xor U22752 (N_22752,N_19435,N_18044);
nor U22753 (N_22753,N_17450,N_15280);
or U22754 (N_22754,N_17543,N_18299);
or U22755 (N_22755,N_15490,N_16986);
nand U22756 (N_22756,N_17444,N_16607);
and U22757 (N_22757,N_16069,N_19507);
xor U22758 (N_22758,N_18093,N_15228);
nor U22759 (N_22759,N_19727,N_15171);
or U22760 (N_22760,N_19258,N_17497);
xor U22761 (N_22761,N_19092,N_18962);
nor U22762 (N_22762,N_17331,N_16638);
and U22763 (N_22763,N_16455,N_19996);
nand U22764 (N_22764,N_18123,N_17872);
nor U22765 (N_22765,N_18565,N_19594);
nor U22766 (N_22766,N_17224,N_17183);
or U22767 (N_22767,N_19211,N_18187);
nor U22768 (N_22768,N_19133,N_17876);
and U22769 (N_22769,N_17584,N_19246);
nand U22770 (N_22770,N_19241,N_16690);
nand U22771 (N_22771,N_18669,N_16951);
and U22772 (N_22772,N_17135,N_16712);
and U22773 (N_22773,N_17973,N_19215);
and U22774 (N_22774,N_15674,N_16397);
xnor U22775 (N_22775,N_15434,N_16848);
nor U22776 (N_22776,N_17371,N_17741);
or U22777 (N_22777,N_18562,N_18512);
nand U22778 (N_22778,N_19975,N_15466);
nor U22779 (N_22779,N_18839,N_19155);
nand U22780 (N_22780,N_16196,N_16977);
xor U22781 (N_22781,N_17059,N_18919);
nand U22782 (N_22782,N_16330,N_18839);
nor U22783 (N_22783,N_17906,N_15607);
and U22784 (N_22784,N_16043,N_19392);
or U22785 (N_22785,N_16696,N_18689);
or U22786 (N_22786,N_19949,N_16901);
nand U22787 (N_22787,N_18181,N_19388);
nand U22788 (N_22788,N_18109,N_19073);
xor U22789 (N_22789,N_18892,N_16840);
xnor U22790 (N_22790,N_17692,N_16488);
or U22791 (N_22791,N_19164,N_18232);
and U22792 (N_22792,N_17004,N_19743);
and U22793 (N_22793,N_15402,N_18582);
nand U22794 (N_22794,N_19281,N_15587);
or U22795 (N_22795,N_16839,N_17255);
xnor U22796 (N_22796,N_17560,N_16587);
or U22797 (N_22797,N_16253,N_18174);
or U22798 (N_22798,N_15108,N_15625);
nor U22799 (N_22799,N_15182,N_15167);
nand U22800 (N_22800,N_16726,N_16812);
xnor U22801 (N_22801,N_18603,N_18095);
nand U22802 (N_22802,N_19479,N_17422);
or U22803 (N_22803,N_18907,N_16359);
or U22804 (N_22804,N_19248,N_15010);
nor U22805 (N_22805,N_18488,N_15978);
nor U22806 (N_22806,N_15962,N_19918);
nor U22807 (N_22807,N_18211,N_18208);
or U22808 (N_22808,N_15477,N_19380);
nand U22809 (N_22809,N_16084,N_16043);
nor U22810 (N_22810,N_17506,N_17674);
and U22811 (N_22811,N_18768,N_18742);
xor U22812 (N_22812,N_16669,N_15742);
and U22813 (N_22813,N_18409,N_16750);
xor U22814 (N_22814,N_17223,N_19304);
and U22815 (N_22815,N_15133,N_15634);
nor U22816 (N_22816,N_16501,N_17216);
nand U22817 (N_22817,N_16844,N_16156);
or U22818 (N_22818,N_17700,N_19951);
or U22819 (N_22819,N_17282,N_15760);
xnor U22820 (N_22820,N_15004,N_15387);
xor U22821 (N_22821,N_18425,N_16787);
or U22822 (N_22822,N_15230,N_18994);
or U22823 (N_22823,N_17408,N_17253);
nand U22824 (N_22824,N_17572,N_15778);
and U22825 (N_22825,N_15252,N_19278);
and U22826 (N_22826,N_17777,N_16698);
nor U22827 (N_22827,N_17997,N_19932);
nor U22828 (N_22828,N_16597,N_17153);
nor U22829 (N_22829,N_16235,N_17431);
and U22830 (N_22830,N_19919,N_15125);
nand U22831 (N_22831,N_17735,N_19159);
nor U22832 (N_22832,N_15175,N_19566);
nand U22833 (N_22833,N_18150,N_18960);
nand U22834 (N_22834,N_18926,N_19562);
or U22835 (N_22835,N_15020,N_18790);
nand U22836 (N_22836,N_17843,N_15771);
or U22837 (N_22837,N_15507,N_17943);
nand U22838 (N_22838,N_17212,N_18708);
and U22839 (N_22839,N_18594,N_19899);
nor U22840 (N_22840,N_16205,N_17412);
nand U22841 (N_22841,N_18931,N_19735);
nand U22842 (N_22842,N_19723,N_18804);
nand U22843 (N_22843,N_15717,N_19811);
nand U22844 (N_22844,N_17055,N_16773);
and U22845 (N_22845,N_19968,N_16917);
nand U22846 (N_22846,N_18406,N_15688);
and U22847 (N_22847,N_17732,N_16859);
and U22848 (N_22848,N_19837,N_16846);
xor U22849 (N_22849,N_16010,N_16261);
and U22850 (N_22850,N_19838,N_18261);
and U22851 (N_22851,N_18620,N_19102);
xor U22852 (N_22852,N_18468,N_17075);
nand U22853 (N_22853,N_16546,N_17516);
and U22854 (N_22854,N_16701,N_17515);
xor U22855 (N_22855,N_17382,N_19363);
nor U22856 (N_22856,N_18611,N_16294);
nand U22857 (N_22857,N_16199,N_17834);
nor U22858 (N_22858,N_17928,N_19144);
and U22859 (N_22859,N_18983,N_17510);
xnor U22860 (N_22860,N_19215,N_19586);
nor U22861 (N_22861,N_17425,N_19387);
nor U22862 (N_22862,N_19048,N_18735);
or U22863 (N_22863,N_15566,N_17690);
or U22864 (N_22864,N_17823,N_19165);
and U22865 (N_22865,N_15804,N_16567);
nand U22866 (N_22866,N_15727,N_19416);
nand U22867 (N_22867,N_15884,N_18868);
nand U22868 (N_22868,N_18806,N_19933);
and U22869 (N_22869,N_15377,N_18321);
nor U22870 (N_22870,N_17545,N_16271);
and U22871 (N_22871,N_19049,N_17634);
and U22872 (N_22872,N_18061,N_17214);
xnor U22873 (N_22873,N_18764,N_18570);
xnor U22874 (N_22874,N_16384,N_18762);
or U22875 (N_22875,N_18382,N_17280);
nand U22876 (N_22876,N_15269,N_16444);
or U22877 (N_22877,N_19681,N_17937);
xnor U22878 (N_22878,N_19553,N_19469);
and U22879 (N_22879,N_15169,N_15095);
and U22880 (N_22880,N_16422,N_16993);
or U22881 (N_22881,N_15395,N_15086);
xnor U22882 (N_22882,N_19167,N_16567);
and U22883 (N_22883,N_18428,N_17186);
or U22884 (N_22884,N_19040,N_18404);
nor U22885 (N_22885,N_17517,N_18429);
or U22886 (N_22886,N_16763,N_15217);
xnor U22887 (N_22887,N_18505,N_17501);
nand U22888 (N_22888,N_18322,N_19016);
nor U22889 (N_22889,N_17517,N_17996);
xor U22890 (N_22890,N_19374,N_18489);
nand U22891 (N_22891,N_16868,N_19790);
or U22892 (N_22892,N_17683,N_16443);
or U22893 (N_22893,N_19242,N_17399);
nor U22894 (N_22894,N_15805,N_17221);
and U22895 (N_22895,N_18895,N_17520);
nand U22896 (N_22896,N_15905,N_18857);
nand U22897 (N_22897,N_19596,N_16656);
nor U22898 (N_22898,N_16486,N_19641);
nand U22899 (N_22899,N_19316,N_15239);
or U22900 (N_22900,N_16857,N_17381);
and U22901 (N_22901,N_19581,N_18420);
nand U22902 (N_22902,N_17614,N_18178);
xor U22903 (N_22903,N_17552,N_16832);
or U22904 (N_22904,N_17033,N_15752);
xnor U22905 (N_22905,N_18139,N_18290);
or U22906 (N_22906,N_16739,N_17266);
nand U22907 (N_22907,N_19323,N_18829);
nor U22908 (N_22908,N_15652,N_15436);
nand U22909 (N_22909,N_19340,N_19576);
or U22910 (N_22910,N_16879,N_19775);
or U22911 (N_22911,N_19367,N_16525);
xnor U22912 (N_22912,N_15857,N_15031);
or U22913 (N_22913,N_16591,N_19330);
xnor U22914 (N_22914,N_19127,N_19521);
xnor U22915 (N_22915,N_18570,N_19128);
or U22916 (N_22916,N_19313,N_18389);
nor U22917 (N_22917,N_17587,N_19543);
and U22918 (N_22918,N_16497,N_18557);
or U22919 (N_22919,N_18530,N_16675);
or U22920 (N_22920,N_19666,N_16009);
nor U22921 (N_22921,N_16992,N_16632);
xnor U22922 (N_22922,N_15507,N_19989);
nand U22923 (N_22923,N_18950,N_16883);
nand U22924 (N_22924,N_16385,N_18735);
or U22925 (N_22925,N_15532,N_16075);
nand U22926 (N_22926,N_19871,N_15782);
nand U22927 (N_22927,N_16000,N_16337);
and U22928 (N_22928,N_16816,N_19155);
and U22929 (N_22929,N_17738,N_16771);
and U22930 (N_22930,N_17103,N_18214);
nor U22931 (N_22931,N_17459,N_19800);
xor U22932 (N_22932,N_16472,N_15685);
nand U22933 (N_22933,N_19963,N_18954);
or U22934 (N_22934,N_16112,N_19231);
xnor U22935 (N_22935,N_19652,N_15525);
nand U22936 (N_22936,N_18482,N_17223);
or U22937 (N_22937,N_19010,N_15086);
and U22938 (N_22938,N_15733,N_15596);
or U22939 (N_22939,N_16760,N_15653);
nand U22940 (N_22940,N_15654,N_18265);
and U22941 (N_22941,N_15426,N_19157);
nand U22942 (N_22942,N_16781,N_18610);
nand U22943 (N_22943,N_15351,N_19402);
and U22944 (N_22944,N_18467,N_15338);
nor U22945 (N_22945,N_15047,N_16131);
or U22946 (N_22946,N_19608,N_18324);
and U22947 (N_22947,N_18527,N_15214);
xnor U22948 (N_22948,N_17005,N_19759);
or U22949 (N_22949,N_16989,N_19037);
nor U22950 (N_22950,N_18902,N_17019);
and U22951 (N_22951,N_16811,N_15957);
nand U22952 (N_22952,N_16771,N_17761);
nand U22953 (N_22953,N_18814,N_16721);
nor U22954 (N_22954,N_16930,N_17269);
xor U22955 (N_22955,N_17030,N_18224);
and U22956 (N_22956,N_18987,N_19438);
or U22957 (N_22957,N_17721,N_16857);
or U22958 (N_22958,N_17237,N_18697);
nor U22959 (N_22959,N_16418,N_16140);
nor U22960 (N_22960,N_18232,N_17346);
and U22961 (N_22961,N_17855,N_18096);
and U22962 (N_22962,N_17296,N_15072);
nand U22963 (N_22963,N_19560,N_17244);
or U22964 (N_22964,N_18563,N_18906);
xor U22965 (N_22965,N_19370,N_17349);
and U22966 (N_22966,N_18340,N_15723);
nand U22967 (N_22967,N_18626,N_17443);
or U22968 (N_22968,N_19133,N_18575);
nand U22969 (N_22969,N_16226,N_18697);
nand U22970 (N_22970,N_17825,N_19239);
nand U22971 (N_22971,N_18003,N_18384);
or U22972 (N_22972,N_17593,N_18611);
nand U22973 (N_22973,N_17544,N_18632);
and U22974 (N_22974,N_16169,N_16445);
or U22975 (N_22975,N_17755,N_18333);
nor U22976 (N_22976,N_18443,N_15745);
and U22977 (N_22977,N_19997,N_17092);
or U22978 (N_22978,N_18989,N_16689);
and U22979 (N_22979,N_17180,N_19224);
xor U22980 (N_22980,N_18600,N_15307);
nand U22981 (N_22981,N_17210,N_18870);
nand U22982 (N_22982,N_16128,N_19263);
nor U22983 (N_22983,N_16656,N_17840);
or U22984 (N_22984,N_19596,N_18231);
or U22985 (N_22985,N_16361,N_15012);
nand U22986 (N_22986,N_16104,N_17243);
and U22987 (N_22987,N_16978,N_19309);
nor U22988 (N_22988,N_18583,N_16245);
or U22989 (N_22989,N_17095,N_18124);
nor U22990 (N_22990,N_16182,N_17748);
nor U22991 (N_22991,N_15073,N_15309);
xor U22992 (N_22992,N_15298,N_15560);
nor U22993 (N_22993,N_19957,N_16051);
nand U22994 (N_22994,N_19649,N_19320);
nand U22995 (N_22995,N_19228,N_15852);
nand U22996 (N_22996,N_16963,N_17038);
nor U22997 (N_22997,N_17277,N_18032);
xor U22998 (N_22998,N_15686,N_18681);
nor U22999 (N_22999,N_17276,N_17196);
xnor U23000 (N_23000,N_16597,N_18799);
and U23001 (N_23001,N_18049,N_15075);
xnor U23002 (N_23002,N_18221,N_19016);
or U23003 (N_23003,N_15382,N_16121);
and U23004 (N_23004,N_17984,N_15712);
or U23005 (N_23005,N_16270,N_16610);
nor U23006 (N_23006,N_19620,N_15161);
nor U23007 (N_23007,N_17125,N_15379);
and U23008 (N_23008,N_15828,N_16262);
nand U23009 (N_23009,N_17267,N_19627);
and U23010 (N_23010,N_17671,N_17039);
or U23011 (N_23011,N_15083,N_16300);
nand U23012 (N_23012,N_18621,N_17078);
nor U23013 (N_23013,N_18760,N_18344);
or U23014 (N_23014,N_15574,N_16456);
and U23015 (N_23015,N_15355,N_17380);
or U23016 (N_23016,N_15090,N_18344);
and U23017 (N_23017,N_18818,N_16580);
xnor U23018 (N_23018,N_19577,N_17740);
nor U23019 (N_23019,N_17943,N_19662);
nor U23020 (N_23020,N_16800,N_16006);
nor U23021 (N_23021,N_17024,N_15252);
xnor U23022 (N_23022,N_16041,N_18366);
nor U23023 (N_23023,N_19763,N_16522);
xor U23024 (N_23024,N_16966,N_16509);
xnor U23025 (N_23025,N_15550,N_18780);
nand U23026 (N_23026,N_16490,N_18547);
and U23027 (N_23027,N_15765,N_19584);
and U23028 (N_23028,N_19593,N_17374);
and U23029 (N_23029,N_15062,N_17575);
nor U23030 (N_23030,N_19099,N_16136);
xnor U23031 (N_23031,N_18832,N_16353);
and U23032 (N_23032,N_19121,N_19642);
or U23033 (N_23033,N_19829,N_16113);
nand U23034 (N_23034,N_17680,N_16923);
xor U23035 (N_23035,N_17253,N_16192);
nor U23036 (N_23036,N_17937,N_16996);
nor U23037 (N_23037,N_19319,N_16768);
nor U23038 (N_23038,N_19582,N_18582);
xnor U23039 (N_23039,N_18807,N_18405);
or U23040 (N_23040,N_16429,N_16327);
nor U23041 (N_23041,N_18855,N_15319);
and U23042 (N_23042,N_16849,N_17462);
and U23043 (N_23043,N_16055,N_16679);
nor U23044 (N_23044,N_17462,N_16078);
nand U23045 (N_23045,N_19094,N_16524);
nor U23046 (N_23046,N_17682,N_19131);
and U23047 (N_23047,N_15624,N_19786);
nor U23048 (N_23048,N_17104,N_19812);
nor U23049 (N_23049,N_16074,N_19374);
and U23050 (N_23050,N_18642,N_17362);
nor U23051 (N_23051,N_18800,N_16326);
xnor U23052 (N_23052,N_18314,N_19936);
nand U23053 (N_23053,N_17480,N_17748);
nor U23054 (N_23054,N_18692,N_17667);
nor U23055 (N_23055,N_19945,N_17014);
xor U23056 (N_23056,N_16723,N_17498);
or U23057 (N_23057,N_15422,N_18051);
or U23058 (N_23058,N_15367,N_17725);
nand U23059 (N_23059,N_18775,N_18938);
xor U23060 (N_23060,N_17496,N_15251);
or U23061 (N_23061,N_17666,N_15597);
nand U23062 (N_23062,N_15367,N_19392);
nand U23063 (N_23063,N_19479,N_15135);
nor U23064 (N_23064,N_18541,N_16951);
nand U23065 (N_23065,N_19874,N_17063);
nor U23066 (N_23066,N_17796,N_16268);
nor U23067 (N_23067,N_15767,N_16746);
nor U23068 (N_23068,N_15082,N_16563);
nand U23069 (N_23069,N_17815,N_19995);
or U23070 (N_23070,N_16583,N_17691);
xor U23071 (N_23071,N_18006,N_19466);
or U23072 (N_23072,N_16365,N_16537);
nand U23073 (N_23073,N_18594,N_15492);
xnor U23074 (N_23074,N_19888,N_17055);
nor U23075 (N_23075,N_16940,N_19869);
nand U23076 (N_23076,N_18892,N_15876);
nand U23077 (N_23077,N_17349,N_16232);
and U23078 (N_23078,N_18138,N_16986);
xnor U23079 (N_23079,N_19430,N_17209);
nor U23080 (N_23080,N_15149,N_16007);
nand U23081 (N_23081,N_16878,N_17200);
nor U23082 (N_23082,N_16924,N_17578);
nor U23083 (N_23083,N_15594,N_16997);
nor U23084 (N_23084,N_18668,N_19471);
xnor U23085 (N_23085,N_17958,N_18255);
nand U23086 (N_23086,N_16547,N_19589);
nand U23087 (N_23087,N_18200,N_19929);
and U23088 (N_23088,N_16381,N_19956);
or U23089 (N_23089,N_16779,N_15812);
nor U23090 (N_23090,N_17897,N_19616);
nor U23091 (N_23091,N_17974,N_17584);
and U23092 (N_23092,N_15396,N_19610);
nor U23093 (N_23093,N_19113,N_16768);
nand U23094 (N_23094,N_17262,N_16958);
or U23095 (N_23095,N_18179,N_18467);
and U23096 (N_23096,N_17467,N_17446);
nand U23097 (N_23097,N_19977,N_18802);
nor U23098 (N_23098,N_19516,N_15571);
and U23099 (N_23099,N_15031,N_16575);
and U23100 (N_23100,N_18216,N_19070);
or U23101 (N_23101,N_18470,N_16550);
and U23102 (N_23102,N_16459,N_15008);
xnor U23103 (N_23103,N_18849,N_19237);
xor U23104 (N_23104,N_17023,N_18518);
nor U23105 (N_23105,N_19095,N_17744);
xnor U23106 (N_23106,N_15130,N_18175);
nand U23107 (N_23107,N_19860,N_17928);
nor U23108 (N_23108,N_16329,N_17828);
and U23109 (N_23109,N_18084,N_15075);
nor U23110 (N_23110,N_17143,N_17342);
nand U23111 (N_23111,N_19547,N_18889);
or U23112 (N_23112,N_17595,N_16081);
nand U23113 (N_23113,N_17767,N_18729);
and U23114 (N_23114,N_17652,N_19073);
and U23115 (N_23115,N_15879,N_19457);
nand U23116 (N_23116,N_17368,N_16788);
nor U23117 (N_23117,N_15947,N_16068);
nor U23118 (N_23118,N_15824,N_18637);
and U23119 (N_23119,N_19783,N_18358);
and U23120 (N_23120,N_18144,N_15018);
or U23121 (N_23121,N_18350,N_15028);
or U23122 (N_23122,N_19212,N_18323);
nor U23123 (N_23123,N_15955,N_15599);
nand U23124 (N_23124,N_18429,N_19460);
or U23125 (N_23125,N_19115,N_16018);
nand U23126 (N_23126,N_15830,N_17845);
nor U23127 (N_23127,N_17095,N_16240);
xor U23128 (N_23128,N_16675,N_19708);
nor U23129 (N_23129,N_17342,N_19293);
or U23130 (N_23130,N_16407,N_16672);
and U23131 (N_23131,N_16706,N_16771);
or U23132 (N_23132,N_17429,N_19053);
xnor U23133 (N_23133,N_17612,N_17793);
nor U23134 (N_23134,N_18712,N_16881);
or U23135 (N_23135,N_19246,N_17567);
or U23136 (N_23136,N_18599,N_18870);
nor U23137 (N_23137,N_15403,N_19739);
nand U23138 (N_23138,N_17208,N_18748);
and U23139 (N_23139,N_16536,N_15697);
or U23140 (N_23140,N_16138,N_19220);
or U23141 (N_23141,N_17393,N_19627);
or U23142 (N_23142,N_16181,N_18418);
nand U23143 (N_23143,N_16753,N_15851);
or U23144 (N_23144,N_19450,N_18201);
or U23145 (N_23145,N_16942,N_17889);
nand U23146 (N_23146,N_15411,N_15539);
nor U23147 (N_23147,N_18276,N_16577);
xor U23148 (N_23148,N_18264,N_19939);
or U23149 (N_23149,N_19465,N_17540);
or U23150 (N_23150,N_16907,N_17727);
nor U23151 (N_23151,N_17874,N_19756);
and U23152 (N_23152,N_17993,N_17946);
or U23153 (N_23153,N_19129,N_15194);
nor U23154 (N_23154,N_15254,N_16322);
nand U23155 (N_23155,N_18565,N_17297);
and U23156 (N_23156,N_18104,N_15094);
nor U23157 (N_23157,N_16171,N_15133);
nor U23158 (N_23158,N_17574,N_17069);
nand U23159 (N_23159,N_15384,N_16218);
nor U23160 (N_23160,N_15745,N_19777);
or U23161 (N_23161,N_15816,N_17057);
nor U23162 (N_23162,N_19907,N_15968);
nand U23163 (N_23163,N_19202,N_19857);
xor U23164 (N_23164,N_18052,N_19635);
nor U23165 (N_23165,N_15127,N_15344);
or U23166 (N_23166,N_17114,N_17553);
xnor U23167 (N_23167,N_17231,N_15701);
or U23168 (N_23168,N_17599,N_15311);
nor U23169 (N_23169,N_16141,N_18110);
and U23170 (N_23170,N_19536,N_15116);
xor U23171 (N_23171,N_19425,N_17668);
or U23172 (N_23172,N_19859,N_17055);
nor U23173 (N_23173,N_19687,N_18880);
nand U23174 (N_23174,N_15290,N_18564);
and U23175 (N_23175,N_17502,N_19878);
or U23176 (N_23176,N_18171,N_15602);
nor U23177 (N_23177,N_15395,N_18654);
xnor U23178 (N_23178,N_18284,N_17518);
xnor U23179 (N_23179,N_15321,N_18828);
xnor U23180 (N_23180,N_19826,N_18116);
and U23181 (N_23181,N_19383,N_16167);
nor U23182 (N_23182,N_19392,N_16345);
or U23183 (N_23183,N_15982,N_19445);
nor U23184 (N_23184,N_15046,N_19564);
nand U23185 (N_23185,N_19460,N_17738);
nand U23186 (N_23186,N_18177,N_16810);
or U23187 (N_23187,N_16644,N_17833);
or U23188 (N_23188,N_15939,N_19665);
nor U23189 (N_23189,N_17451,N_16289);
or U23190 (N_23190,N_19151,N_17486);
nor U23191 (N_23191,N_15170,N_18644);
and U23192 (N_23192,N_16196,N_15741);
nand U23193 (N_23193,N_18745,N_19613);
or U23194 (N_23194,N_17247,N_16076);
nor U23195 (N_23195,N_17828,N_15178);
or U23196 (N_23196,N_16502,N_18437);
or U23197 (N_23197,N_19699,N_16099);
nand U23198 (N_23198,N_19226,N_15412);
or U23199 (N_23199,N_19216,N_17812);
nor U23200 (N_23200,N_16563,N_19731);
and U23201 (N_23201,N_15264,N_17994);
and U23202 (N_23202,N_18641,N_15654);
nor U23203 (N_23203,N_17725,N_19410);
and U23204 (N_23204,N_15721,N_16627);
nor U23205 (N_23205,N_18163,N_16927);
and U23206 (N_23206,N_15541,N_19745);
xor U23207 (N_23207,N_19192,N_17445);
nor U23208 (N_23208,N_16616,N_19740);
xnor U23209 (N_23209,N_19266,N_18445);
xor U23210 (N_23210,N_16894,N_16400);
nand U23211 (N_23211,N_15443,N_17767);
xnor U23212 (N_23212,N_16796,N_16072);
or U23213 (N_23213,N_15586,N_15449);
and U23214 (N_23214,N_19292,N_19926);
nand U23215 (N_23215,N_17655,N_16197);
or U23216 (N_23216,N_18097,N_17996);
nor U23217 (N_23217,N_16972,N_19671);
nor U23218 (N_23218,N_18355,N_16811);
nand U23219 (N_23219,N_17142,N_19130);
nor U23220 (N_23220,N_18146,N_18620);
nor U23221 (N_23221,N_15174,N_16625);
or U23222 (N_23222,N_19884,N_17220);
or U23223 (N_23223,N_16287,N_17594);
and U23224 (N_23224,N_16502,N_17749);
nand U23225 (N_23225,N_19144,N_19672);
and U23226 (N_23226,N_15066,N_18869);
or U23227 (N_23227,N_15324,N_15894);
and U23228 (N_23228,N_16320,N_17821);
nor U23229 (N_23229,N_16612,N_19306);
nor U23230 (N_23230,N_15213,N_16531);
and U23231 (N_23231,N_15048,N_16441);
nand U23232 (N_23232,N_16720,N_18172);
nor U23233 (N_23233,N_19981,N_17770);
nor U23234 (N_23234,N_18462,N_19706);
and U23235 (N_23235,N_19559,N_15192);
nor U23236 (N_23236,N_18427,N_18370);
nand U23237 (N_23237,N_15073,N_19597);
or U23238 (N_23238,N_18126,N_18432);
xor U23239 (N_23239,N_18472,N_15732);
nor U23240 (N_23240,N_19771,N_15634);
nand U23241 (N_23241,N_19706,N_18594);
and U23242 (N_23242,N_18831,N_16954);
nor U23243 (N_23243,N_18921,N_19794);
or U23244 (N_23244,N_17785,N_19860);
nor U23245 (N_23245,N_15238,N_15555);
nand U23246 (N_23246,N_15576,N_18126);
nand U23247 (N_23247,N_16212,N_16664);
nor U23248 (N_23248,N_19714,N_15064);
nor U23249 (N_23249,N_15225,N_18247);
nor U23250 (N_23250,N_19865,N_17861);
or U23251 (N_23251,N_16335,N_17995);
and U23252 (N_23252,N_18334,N_17197);
xor U23253 (N_23253,N_15608,N_15341);
or U23254 (N_23254,N_16727,N_15648);
xnor U23255 (N_23255,N_17623,N_16240);
nand U23256 (N_23256,N_19000,N_17183);
nand U23257 (N_23257,N_15872,N_15403);
and U23258 (N_23258,N_15103,N_17495);
nor U23259 (N_23259,N_16673,N_15945);
xnor U23260 (N_23260,N_16628,N_18601);
nand U23261 (N_23261,N_19485,N_17871);
xor U23262 (N_23262,N_15502,N_16647);
nor U23263 (N_23263,N_15330,N_18092);
or U23264 (N_23264,N_19237,N_19187);
and U23265 (N_23265,N_17252,N_18121);
or U23266 (N_23266,N_16997,N_17121);
nand U23267 (N_23267,N_18696,N_15729);
and U23268 (N_23268,N_17617,N_18094);
nand U23269 (N_23269,N_15275,N_19418);
xor U23270 (N_23270,N_15953,N_19636);
xor U23271 (N_23271,N_17815,N_16059);
nor U23272 (N_23272,N_16438,N_16743);
and U23273 (N_23273,N_19172,N_15598);
xor U23274 (N_23274,N_19113,N_16756);
or U23275 (N_23275,N_19346,N_16675);
nand U23276 (N_23276,N_18379,N_18366);
and U23277 (N_23277,N_17918,N_19356);
xor U23278 (N_23278,N_15554,N_15286);
nand U23279 (N_23279,N_17365,N_16576);
nor U23280 (N_23280,N_17182,N_16147);
or U23281 (N_23281,N_18885,N_17922);
or U23282 (N_23282,N_17754,N_18501);
and U23283 (N_23283,N_16208,N_19527);
or U23284 (N_23284,N_17241,N_15689);
nor U23285 (N_23285,N_16550,N_19579);
nor U23286 (N_23286,N_18176,N_19377);
and U23287 (N_23287,N_18900,N_18653);
and U23288 (N_23288,N_18267,N_16905);
nor U23289 (N_23289,N_16965,N_17636);
nand U23290 (N_23290,N_17150,N_15538);
or U23291 (N_23291,N_17189,N_17207);
and U23292 (N_23292,N_19302,N_18974);
nor U23293 (N_23293,N_18746,N_19029);
or U23294 (N_23294,N_19734,N_17078);
xor U23295 (N_23295,N_16342,N_18829);
nor U23296 (N_23296,N_19651,N_19789);
or U23297 (N_23297,N_16118,N_15193);
nand U23298 (N_23298,N_19531,N_18302);
nor U23299 (N_23299,N_19271,N_19069);
or U23300 (N_23300,N_18251,N_16267);
or U23301 (N_23301,N_19634,N_18819);
and U23302 (N_23302,N_18969,N_17861);
nand U23303 (N_23303,N_17627,N_18707);
and U23304 (N_23304,N_17165,N_19476);
nor U23305 (N_23305,N_18742,N_15855);
or U23306 (N_23306,N_18081,N_18255);
or U23307 (N_23307,N_18258,N_18751);
nand U23308 (N_23308,N_15767,N_17510);
nand U23309 (N_23309,N_15189,N_16875);
nor U23310 (N_23310,N_16681,N_19867);
or U23311 (N_23311,N_18518,N_17990);
nor U23312 (N_23312,N_16717,N_15237);
nand U23313 (N_23313,N_16459,N_19835);
and U23314 (N_23314,N_18887,N_18789);
nor U23315 (N_23315,N_16025,N_17881);
and U23316 (N_23316,N_17821,N_19081);
and U23317 (N_23317,N_19680,N_19204);
nand U23318 (N_23318,N_18883,N_19145);
nor U23319 (N_23319,N_15708,N_15358);
nor U23320 (N_23320,N_18241,N_18222);
nand U23321 (N_23321,N_18416,N_19157);
and U23322 (N_23322,N_19167,N_18068);
and U23323 (N_23323,N_17226,N_17327);
nand U23324 (N_23324,N_17618,N_17634);
or U23325 (N_23325,N_19942,N_19509);
nand U23326 (N_23326,N_16452,N_15930);
nor U23327 (N_23327,N_17048,N_16918);
and U23328 (N_23328,N_16686,N_18999);
xor U23329 (N_23329,N_17115,N_16297);
or U23330 (N_23330,N_17534,N_19033);
and U23331 (N_23331,N_16025,N_16715);
or U23332 (N_23332,N_17176,N_15369);
and U23333 (N_23333,N_19277,N_16631);
nand U23334 (N_23334,N_17277,N_18962);
nand U23335 (N_23335,N_16315,N_15329);
xor U23336 (N_23336,N_19032,N_18713);
nand U23337 (N_23337,N_15143,N_15503);
and U23338 (N_23338,N_17179,N_17100);
or U23339 (N_23339,N_19128,N_15313);
nand U23340 (N_23340,N_18315,N_16406);
or U23341 (N_23341,N_17853,N_17274);
and U23342 (N_23342,N_15422,N_16906);
nand U23343 (N_23343,N_15407,N_17555);
nor U23344 (N_23344,N_17563,N_18558);
or U23345 (N_23345,N_15817,N_19710);
nand U23346 (N_23346,N_18877,N_17835);
or U23347 (N_23347,N_17673,N_16466);
nor U23348 (N_23348,N_19751,N_19152);
nor U23349 (N_23349,N_15814,N_15629);
or U23350 (N_23350,N_18510,N_17794);
nor U23351 (N_23351,N_18584,N_15391);
and U23352 (N_23352,N_19805,N_19621);
xnor U23353 (N_23353,N_18265,N_18321);
nor U23354 (N_23354,N_18601,N_17871);
xor U23355 (N_23355,N_18350,N_19132);
or U23356 (N_23356,N_15439,N_19978);
nand U23357 (N_23357,N_17784,N_15801);
xor U23358 (N_23358,N_18390,N_17672);
and U23359 (N_23359,N_19799,N_18722);
and U23360 (N_23360,N_17522,N_17450);
or U23361 (N_23361,N_18113,N_17056);
or U23362 (N_23362,N_17193,N_17810);
or U23363 (N_23363,N_17482,N_18551);
nand U23364 (N_23364,N_15525,N_18968);
and U23365 (N_23365,N_17576,N_19614);
or U23366 (N_23366,N_19282,N_15083);
or U23367 (N_23367,N_18836,N_18691);
and U23368 (N_23368,N_15475,N_18887);
nor U23369 (N_23369,N_17944,N_16473);
nor U23370 (N_23370,N_15766,N_16872);
nand U23371 (N_23371,N_16806,N_16326);
nand U23372 (N_23372,N_17676,N_18819);
or U23373 (N_23373,N_15652,N_17211);
nand U23374 (N_23374,N_15982,N_18236);
nand U23375 (N_23375,N_19846,N_19563);
or U23376 (N_23376,N_17891,N_19775);
nor U23377 (N_23377,N_19494,N_19853);
xnor U23378 (N_23378,N_15982,N_16034);
and U23379 (N_23379,N_16154,N_19013);
xor U23380 (N_23380,N_16701,N_17107);
or U23381 (N_23381,N_18285,N_17833);
or U23382 (N_23382,N_16496,N_15720);
nor U23383 (N_23383,N_16997,N_17542);
nor U23384 (N_23384,N_15594,N_19119);
nor U23385 (N_23385,N_18672,N_18765);
xnor U23386 (N_23386,N_17861,N_16382);
nand U23387 (N_23387,N_17600,N_17698);
or U23388 (N_23388,N_16742,N_17940);
and U23389 (N_23389,N_16901,N_15396);
and U23390 (N_23390,N_15901,N_15309);
or U23391 (N_23391,N_19215,N_19907);
nor U23392 (N_23392,N_19495,N_17186);
or U23393 (N_23393,N_19298,N_17633);
or U23394 (N_23394,N_17737,N_18025);
or U23395 (N_23395,N_19540,N_17894);
nor U23396 (N_23396,N_19998,N_19737);
xor U23397 (N_23397,N_18254,N_15615);
nor U23398 (N_23398,N_19455,N_17776);
or U23399 (N_23399,N_19115,N_16312);
nand U23400 (N_23400,N_17926,N_19017);
and U23401 (N_23401,N_19861,N_19321);
or U23402 (N_23402,N_17694,N_16811);
nor U23403 (N_23403,N_19693,N_16059);
or U23404 (N_23404,N_19444,N_16088);
nand U23405 (N_23405,N_16459,N_17515);
or U23406 (N_23406,N_15576,N_19823);
nor U23407 (N_23407,N_18929,N_16374);
xnor U23408 (N_23408,N_19928,N_19977);
or U23409 (N_23409,N_17313,N_17950);
and U23410 (N_23410,N_15518,N_18401);
nor U23411 (N_23411,N_17415,N_17217);
or U23412 (N_23412,N_17500,N_17335);
nand U23413 (N_23413,N_16451,N_19098);
and U23414 (N_23414,N_16103,N_19939);
xor U23415 (N_23415,N_16909,N_19154);
or U23416 (N_23416,N_19805,N_16384);
nand U23417 (N_23417,N_16449,N_15598);
nand U23418 (N_23418,N_16515,N_18336);
or U23419 (N_23419,N_19878,N_15964);
nand U23420 (N_23420,N_19939,N_19769);
nand U23421 (N_23421,N_18048,N_15087);
or U23422 (N_23422,N_16740,N_18822);
and U23423 (N_23423,N_18356,N_15876);
nor U23424 (N_23424,N_19970,N_18196);
and U23425 (N_23425,N_15154,N_16035);
nand U23426 (N_23426,N_19803,N_17909);
or U23427 (N_23427,N_15590,N_19642);
nand U23428 (N_23428,N_19538,N_16733);
nand U23429 (N_23429,N_15784,N_18908);
and U23430 (N_23430,N_15083,N_19269);
or U23431 (N_23431,N_16513,N_16031);
or U23432 (N_23432,N_17597,N_17991);
and U23433 (N_23433,N_18701,N_16698);
or U23434 (N_23434,N_16201,N_16198);
or U23435 (N_23435,N_19429,N_18333);
nor U23436 (N_23436,N_17831,N_15545);
nor U23437 (N_23437,N_15920,N_18249);
nand U23438 (N_23438,N_18030,N_18700);
nor U23439 (N_23439,N_17537,N_19727);
nand U23440 (N_23440,N_19545,N_16306);
nor U23441 (N_23441,N_15813,N_18342);
and U23442 (N_23442,N_19391,N_15292);
nor U23443 (N_23443,N_17764,N_18621);
nor U23444 (N_23444,N_18456,N_15859);
nand U23445 (N_23445,N_15926,N_17707);
nand U23446 (N_23446,N_16452,N_18081);
nand U23447 (N_23447,N_19845,N_16582);
or U23448 (N_23448,N_19978,N_16305);
and U23449 (N_23449,N_19369,N_19508);
nand U23450 (N_23450,N_17415,N_17739);
nor U23451 (N_23451,N_16660,N_17328);
or U23452 (N_23452,N_18581,N_18959);
nor U23453 (N_23453,N_15826,N_17748);
and U23454 (N_23454,N_18939,N_15431);
or U23455 (N_23455,N_16982,N_19304);
nor U23456 (N_23456,N_16393,N_16943);
or U23457 (N_23457,N_15133,N_18649);
and U23458 (N_23458,N_16937,N_16179);
nand U23459 (N_23459,N_15435,N_19898);
nand U23460 (N_23460,N_19838,N_18390);
or U23461 (N_23461,N_17817,N_18702);
and U23462 (N_23462,N_15696,N_18598);
nand U23463 (N_23463,N_15499,N_18470);
nand U23464 (N_23464,N_19470,N_17830);
or U23465 (N_23465,N_16936,N_17120);
nand U23466 (N_23466,N_15984,N_15224);
or U23467 (N_23467,N_17071,N_19490);
nor U23468 (N_23468,N_15919,N_17787);
nand U23469 (N_23469,N_16452,N_18375);
nor U23470 (N_23470,N_15678,N_19890);
or U23471 (N_23471,N_15501,N_15387);
nand U23472 (N_23472,N_19904,N_19604);
and U23473 (N_23473,N_16686,N_16364);
and U23474 (N_23474,N_18231,N_18711);
xnor U23475 (N_23475,N_17288,N_18597);
and U23476 (N_23476,N_15456,N_18504);
and U23477 (N_23477,N_18198,N_19872);
nand U23478 (N_23478,N_15728,N_15414);
and U23479 (N_23479,N_18222,N_17267);
xnor U23480 (N_23480,N_17932,N_18947);
xor U23481 (N_23481,N_16713,N_15455);
or U23482 (N_23482,N_17282,N_15301);
or U23483 (N_23483,N_18638,N_15625);
nor U23484 (N_23484,N_18353,N_17657);
xor U23485 (N_23485,N_15824,N_18968);
or U23486 (N_23486,N_15569,N_17263);
xor U23487 (N_23487,N_17857,N_15506);
nand U23488 (N_23488,N_19966,N_15245);
or U23489 (N_23489,N_18889,N_15759);
and U23490 (N_23490,N_17379,N_18992);
or U23491 (N_23491,N_18985,N_17068);
nor U23492 (N_23492,N_15411,N_19018);
nor U23493 (N_23493,N_17616,N_16240);
nand U23494 (N_23494,N_18008,N_17003);
xor U23495 (N_23495,N_15501,N_19976);
and U23496 (N_23496,N_18192,N_16364);
and U23497 (N_23497,N_15568,N_18151);
nor U23498 (N_23498,N_17483,N_17011);
nand U23499 (N_23499,N_17571,N_16555);
and U23500 (N_23500,N_16071,N_15091);
or U23501 (N_23501,N_19316,N_15812);
and U23502 (N_23502,N_18224,N_16688);
nand U23503 (N_23503,N_18231,N_15123);
nand U23504 (N_23504,N_19248,N_17455);
and U23505 (N_23505,N_18472,N_19295);
xnor U23506 (N_23506,N_15998,N_17930);
nor U23507 (N_23507,N_16743,N_18145);
nand U23508 (N_23508,N_17915,N_18284);
and U23509 (N_23509,N_15879,N_15254);
or U23510 (N_23510,N_16098,N_18907);
nand U23511 (N_23511,N_16578,N_17759);
nor U23512 (N_23512,N_16983,N_19632);
or U23513 (N_23513,N_17690,N_16888);
nand U23514 (N_23514,N_19829,N_18093);
and U23515 (N_23515,N_16361,N_15557);
or U23516 (N_23516,N_17751,N_15843);
and U23517 (N_23517,N_18050,N_19003);
nand U23518 (N_23518,N_17057,N_16629);
nand U23519 (N_23519,N_15298,N_17994);
and U23520 (N_23520,N_16542,N_18284);
or U23521 (N_23521,N_15762,N_18441);
or U23522 (N_23522,N_19993,N_15961);
nand U23523 (N_23523,N_18366,N_19595);
nand U23524 (N_23524,N_18899,N_16448);
or U23525 (N_23525,N_18912,N_17510);
nand U23526 (N_23526,N_17184,N_17198);
nand U23527 (N_23527,N_16001,N_19163);
nand U23528 (N_23528,N_17354,N_18529);
xnor U23529 (N_23529,N_15279,N_18180);
nor U23530 (N_23530,N_15612,N_18402);
nor U23531 (N_23531,N_18885,N_18752);
xor U23532 (N_23532,N_19001,N_15672);
or U23533 (N_23533,N_17419,N_18767);
and U23534 (N_23534,N_17007,N_16781);
and U23535 (N_23535,N_15264,N_18372);
nand U23536 (N_23536,N_18005,N_17187);
nor U23537 (N_23537,N_18574,N_19226);
or U23538 (N_23538,N_19328,N_15484);
or U23539 (N_23539,N_15193,N_15271);
or U23540 (N_23540,N_18153,N_19659);
xnor U23541 (N_23541,N_16576,N_16561);
or U23542 (N_23542,N_16556,N_17361);
nor U23543 (N_23543,N_19863,N_19557);
and U23544 (N_23544,N_15385,N_16176);
nand U23545 (N_23545,N_16098,N_19253);
nand U23546 (N_23546,N_15786,N_16561);
nand U23547 (N_23547,N_18670,N_16615);
or U23548 (N_23548,N_17567,N_15274);
nand U23549 (N_23549,N_18966,N_18282);
and U23550 (N_23550,N_17829,N_19790);
or U23551 (N_23551,N_19726,N_17244);
xor U23552 (N_23552,N_17351,N_16562);
and U23553 (N_23553,N_15148,N_15851);
and U23554 (N_23554,N_19372,N_18568);
nand U23555 (N_23555,N_17815,N_15734);
and U23556 (N_23556,N_18596,N_19862);
nand U23557 (N_23557,N_17178,N_15688);
nor U23558 (N_23558,N_17486,N_18559);
xor U23559 (N_23559,N_18055,N_18496);
or U23560 (N_23560,N_17336,N_16730);
xnor U23561 (N_23561,N_15529,N_15270);
nand U23562 (N_23562,N_19939,N_19382);
nand U23563 (N_23563,N_15189,N_16493);
nor U23564 (N_23564,N_15428,N_18167);
nor U23565 (N_23565,N_18871,N_17606);
or U23566 (N_23566,N_15726,N_19773);
nor U23567 (N_23567,N_18771,N_15915);
xor U23568 (N_23568,N_17261,N_16780);
nor U23569 (N_23569,N_18823,N_19671);
and U23570 (N_23570,N_19295,N_18122);
nor U23571 (N_23571,N_18362,N_18821);
nor U23572 (N_23572,N_17105,N_18215);
and U23573 (N_23573,N_15326,N_18844);
and U23574 (N_23574,N_15162,N_17864);
and U23575 (N_23575,N_15344,N_17880);
xor U23576 (N_23576,N_18675,N_17803);
or U23577 (N_23577,N_15667,N_15043);
nor U23578 (N_23578,N_18963,N_19420);
nand U23579 (N_23579,N_15813,N_15054);
nor U23580 (N_23580,N_18462,N_17628);
nand U23581 (N_23581,N_18296,N_16829);
nand U23582 (N_23582,N_19875,N_18873);
and U23583 (N_23583,N_17481,N_15578);
and U23584 (N_23584,N_17916,N_16031);
and U23585 (N_23585,N_15646,N_18565);
and U23586 (N_23586,N_19786,N_15507);
nand U23587 (N_23587,N_15114,N_17927);
nand U23588 (N_23588,N_19898,N_16612);
or U23589 (N_23589,N_16256,N_17982);
xor U23590 (N_23590,N_15139,N_17470);
nand U23591 (N_23591,N_15595,N_19007);
nor U23592 (N_23592,N_19785,N_15674);
and U23593 (N_23593,N_18210,N_17133);
and U23594 (N_23594,N_18596,N_17086);
nand U23595 (N_23595,N_15720,N_18741);
nor U23596 (N_23596,N_16849,N_19489);
nand U23597 (N_23597,N_16967,N_16700);
and U23598 (N_23598,N_19724,N_18521);
nor U23599 (N_23599,N_16954,N_18565);
nand U23600 (N_23600,N_18327,N_18260);
nand U23601 (N_23601,N_17403,N_18068);
nor U23602 (N_23602,N_17121,N_16531);
nor U23603 (N_23603,N_15497,N_18377);
and U23604 (N_23604,N_18723,N_17412);
nor U23605 (N_23605,N_16678,N_19785);
and U23606 (N_23606,N_15187,N_19813);
nor U23607 (N_23607,N_17538,N_17665);
or U23608 (N_23608,N_18316,N_17379);
nor U23609 (N_23609,N_19332,N_17774);
nand U23610 (N_23610,N_16095,N_15144);
nor U23611 (N_23611,N_16436,N_18503);
xor U23612 (N_23612,N_16114,N_18871);
and U23613 (N_23613,N_15493,N_18868);
nor U23614 (N_23614,N_17883,N_19159);
or U23615 (N_23615,N_15881,N_16420);
nor U23616 (N_23616,N_17480,N_15447);
or U23617 (N_23617,N_16078,N_18441);
nor U23618 (N_23618,N_19406,N_16713);
and U23619 (N_23619,N_16224,N_19068);
nand U23620 (N_23620,N_16225,N_18768);
nand U23621 (N_23621,N_18298,N_17256);
and U23622 (N_23622,N_17940,N_17084);
or U23623 (N_23623,N_16573,N_18237);
nor U23624 (N_23624,N_15982,N_15979);
nor U23625 (N_23625,N_17357,N_17389);
nor U23626 (N_23626,N_19575,N_17973);
nor U23627 (N_23627,N_15837,N_19717);
and U23628 (N_23628,N_19948,N_16675);
nand U23629 (N_23629,N_19238,N_18703);
nor U23630 (N_23630,N_15141,N_16292);
nor U23631 (N_23631,N_17478,N_16155);
nor U23632 (N_23632,N_18421,N_19005);
and U23633 (N_23633,N_16391,N_19918);
xor U23634 (N_23634,N_18913,N_19934);
or U23635 (N_23635,N_18036,N_19680);
or U23636 (N_23636,N_18231,N_19570);
nor U23637 (N_23637,N_15145,N_19480);
or U23638 (N_23638,N_16735,N_17277);
nor U23639 (N_23639,N_18425,N_17525);
nor U23640 (N_23640,N_17675,N_18778);
nor U23641 (N_23641,N_17115,N_17679);
nor U23642 (N_23642,N_19086,N_18992);
nand U23643 (N_23643,N_17645,N_16196);
and U23644 (N_23644,N_15350,N_15305);
or U23645 (N_23645,N_17131,N_16827);
xnor U23646 (N_23646,N_16910,N_17757);
or U23647 (N_23647,N_17335,N_16595);
nand U23648 (N_23648,N_17054,N_15295);
or U23649 (N_23649,N_15852,N_16084);
or U23650 (N_23650,N_15746,N_16377);
and U23651 (N_23651,N_15183,N_15218);
nand U23652 (N_23652,N_18133,N_16686);
xor U23653 (N_23653,N_15495,N_15183);
nor U23654 (N_23654,N_15636,N_15065);
or U23655 (N_23655,N_19382,N_18346);
or U23656 (N_23656,N_17637,N_15894);
or U23657 (N_23657,N_15505,N_15205);
or U23658 (N_23658,N_18412,N_16577);
nor U23659 (N_23659,N_16927,N_17023);
nor U23660 (N_23660,N_15445,N_15524);
or U23661 (N_23661,N_19535,N_16892);
nor U23662 (N_23662,N_19042,N_19173);
nand U23663 (N_23663,N_19281,N_17903);
and U23664 (N_23664,N_15760,N_15563);
and U23665 (N_23665,N_19798,N_17497);
nand U23666 (N_23666,N_15612,N_15822);
or U23667 (N_23667,N_15435,N_19203);
or U23668 (N_23668,N_19958,N_17260);
xor U23669 (N_23669,N_18365,N_19703);
nor U23670 (N_23670,N_17313,N_16767);
and U23671 (N_23671,N_17859,N_15911);
nand U23672 (N_23672,N_15409,N_17328);
nand U23673 (N_23673,N_16039,N_18036);
and U23674 (N_23674,N_15876,N_19113);
and U23675 (N_23675,N_18129,N_17369);
nand U23676 (N_23676,N_16786,N_16593);
nor U23677 (N_23677,N_17648,N_17377);
or U23678 (N_23678,N_17697,N_18193);
nand U23679 (N_23679,N_16729,N_15678);
nand U23680 (N_23680,N_16109,N_16785);
and U23681 (N_23681,N_19805,N_17803);
or U23682 (N_23682,N_19868,N_19430);
nand U23683 (N_23683,N_17778,N_19229);
nand U23684 (N_23684,N_18858,N_17704);
or U23685 (N_23685,N_19025,N_19503);
nor U23686 (N_23686,N_17217,N_16136);
and U23687 (N_23687,N_15650,N_15512);
nor U23688 (N_23688,N_18316,N_16246);
nand U23689 (N_23689,N_19762,N_19585);
or U23690 (N_23690,N_18477,N_19687);
nor U23691 (N_23691,N_15618,N_18232);
xor U23692 (N_23692,N_15473,N_15575);
or U23693 (N_23693,N_17292,N_15338);
or U23694 (N_23694,N_18310,N_16115);
nor U23695 (N_23695,N_15494,N_17709);
nand U23696 (N_23696,N_19078,N_17508);
nand U23697 (N_23697,N_16562,N_15412);
nand U23698 (N_23698,N_19259,N_17744);
nor U23699 (N_23699,N_17717,N_15167);
xnor U23700 (N_23700,N_15113,N_18712);
or U23701 (N_23701,N_18643,N_15355);
nor U23702 (N_23702,N_16633,N_18862);
xor U23703 (N_23703,N_16541,N_17328);
and U23704 (N_23704,N_16797,N_15194);
nor U23705 (N_23705,N_18597,N_16462);
nor U23706 (N_23706,N_18860,N_19317);
nor U23707 (N_23707,N_19967,N_18563);
or U23708 (N_23708,N_17483,N_15395);
and U23709 (N_23709,N_15392,N_17692);
and U23710 (N_23710,N_19587,N_15436);
xnor U23711 (N_23711,N_19760,N_18518);
and U23712 (N_23712,N_16193,N_19949);
or U23713 (N_23713,N_17701,N_19570);
or U23714 (N_23714,N_16753,N_15329);
and U23715 (N_23715,N_16541,N_18420);
nand U23716 (N_23716,N_17665,N_17283);
and U23717 (N_23717,N_18195,N_15173);
or U23718 (N_23718,N_15647,N_19221);
or U23719 (N_23719,N_15497,N_15421);
xnor U23720 (N_23720,N_17794,N_17773);
or U23721 (N_23721,N_19589,N_15282);
nand U23722 (N_23722,N_18246,N_19688);
nand U23723 (N_23723,N_18647,N_17290);
nand U23724 (N_23724,N_18724,N_16982);
or U23725 (N_23725,N_16179,N_15391);
nor U23726 (N_23726,N_18530,N_15177);
xor U23727 (N_23727,N_19156,N_19409);
or U23728 (N_23728,N_19651,N_15004);
nor U23729 (N_23729,N_15347,N_18237);
nand U23730 (N_23730,N_15971,N_16481);
nor U23731 (N_23731,N_19155,N_18993);
or U23732 (N_23732,N_15727,N_17025);
xnor U23733 (N_23733,N_17750,N_16640);
and U23734 (N_23734,N_15469,N_19006);
nand U23735 (N_23735,N_16569,N_17960);
or U23736 (N_23736,N_15346,N_15198);
and U23737 (N_23737,N_16613,N_19348);
nand U23738 (N_23738,N_16107,N_17790);
nand U23739 (N_23739,N_15564,N_17157);
and U23740 (N_23740,N_16924,N_17534);
nand U23741 (N_23741,N_19935,N_18723);
nand U23742 (N_23742,N_18377,N_18551);
or U23743 (N_23743,N_18558,N_16726);
or U23744 (N_23744,N_19627,N_15547);
nor U23745 (N_23745,N_17696,N_17680);
nor U23746 (N_23746,N_17659,N_17574);
and U23747 (N_23747,N_19985,N_19110);
nor U23748 (N_23748,N_18780,N_15623);
and U23749 (N_23749,N_16552,N_15430);
and U23750 (N_23750,N_17155,N_16711);
nand U23751 (N_23751,N_15133,N_19427);
or U23752 (N_23752,N_17027,N_16809);
nand U23753 (N_23753,N_17676,N_15877);
or U23754 (N_23754,N_17016,N_19202);
nor U23755 (N_23755,N_17433,N_18172);
nand U23756 (N_23756,N_15619,N_17260);
nand U23757 (N_23757,N_17638,N_17537);
and U23758 (N_23758,N_19678,N_19633);
and U23759 (N_23759,N_18862,N_18429);
xor U23760 (N_23760,N_18100,N_16380);
nand U23761 (N_23761,N_15537,N_17637);
nor U23762 (N_23762,N_19236,N_18825);
nor U23763 (N_23763,N_16051,N_15588);
nand U23764 (N_23764,N_16524,N_18806);
nand U23765 (N_23765,N_18720,N_15485);
nor U23766 (N_23766,N_17488,N_19236);
or U23767 (N_23767,N_17369,N_18963);
xor U23768 (N_23768,N_15584,N_19233);
and U23769 (N_23769,N_15418,N_17969);
nand U23770 (N_23770,N_18755,N_16553);
nand U23771 (N_23771,N_15854,N_18470);
or U23772 (N_23772,N_17988,N_16439);
nand U23773 (N_23773,N_15936,N_17441);
nor U23774 (N_23774,N_19835,N_18646);
or U23775 (N_23775,N_18542,N_19976);
or U23776 (N_23776,N_19090,N_18709);
and U23777 (N_23777,N_15981,N_15274);
nor U23778 (N_23778,N_17219,N_15412);
or U23779 (N_23779,N_18544,N_17427);
xnor U23780 (N_23780,N_17074,N_17438);
nor U23781 (N_23781,N_15984,N_17861);
or U23782 (N_23782,N_19724,N_15144);
nor U23783 (N_23783,N_15538,N_18231);
or U23784 (N_23784,N_18578,N_17150);
or U23785 (N_23785,N_18781,N_19393);
nand U23786 (N_23786,N_19640,N_18063);
nor U23787 (N_23787,N_18798,N_17128);
nor U23788 (N_23788,N_16817,N_19962);
nand U23789 (N_23789,N_16547,N_16393);
nand U23790 (N_23790,N_16900,N_15056);
and U23791 (N_23791,N_16886,N_16995);
xnor U23792 (N_23792,N_19000,N_15776);
nor U23793 (N_23793,N_15675,N_15053);
and U23794 (N_23794,N_19210,N_17926);
nor U23795 (N_23795,N_16250,N_19735);
nand U23796 (N_23796,N_18800,N_16842);
and U23797 (N_23797,N_18001,N_19348);
or U23798 (N_23798,N_16047,N_15638);
or U23799 (N_23799,N_17904,N_17090);
or U23800 (N_23800,N_15864,N_16645);
and U23801 (N_23801,N_19415,N_18276);
nor U23802 (N_23802,N_17979,N_17225);
nand U23803 (N_23803,N_19545,N_19320);
nand U23804 (N_23804,N_17770,N_17569);
xor U23805 (N_23805,N_18531,N_17896);
or U23806 (N_23806,N_17260,N_16060);
or U23807 (N_23807,N_18516,N_17371);
nand U23808 (N_23808,N_16781,N_15663);
or U23809 (N_23809,N_17890,N_19781);
or U23810 (N_23810,N_17367,N_15439);
nand U23811 (N_23811,N_17759,N_16649);
nor U23812 (N_23812,N_18842,N_17379);
or U23813 (N_23813,N_17749,N_18417);
nor U23814 (N_23814,N_16114,N_18006);
nand U23815 (N_23815,N_18227,N_17667);
nand U23816 (N_23816,N_15846,N_15786);
or U23817 (N_23817,N_17178,N_18998);
nor U23818 (N_23818,N_18759,N_18486);
and U23819 (N_23819,N_17628,N_18261);
or U23820 (N_23820,N_16037,N_16305);
nand U23821 (N_23821,N_18515,N_15902);
nand U23822 (N_23822,N_16288,N_16406);
and U23823 (N_23823,N_17499,N_17263);
xnor U23824 (N_23824,N_18174,N_16654);
and U23825 (N_23825,N_16642,N_19260);
or U23826 (N_23826,N_17631,N_15064);
nor U23827 (N_23827,N_16681,N_16383);
and U23828 (N_23828,N_18003,N_19488);
or U23829 (N_23829,N_19626,N_19275);
or U23830 (N_23830,N_15411,N_17645);
nand U23831 (N_23831,N_15564,N_15534);
and U23832 (N_23832,N_18676,N_16509);
or U23833 (N_23833,N_19286,N_19563);
xnor U23834 (N_23834,N_19978,N_19316);
xor U23835 (N_23835,N_19592,N_15791);
nand U23836 (N_23836,N_17248,N_19353);
and U23837 (N_23837,N_19792,N_19805);
nand U23838 (N_23838,N_16277,N_17705);
nand U23839 (N_23839,N_19537,N_16096);
or U23840 (N_23840,N_19976,N_16865);
nand U23841 (N_23841,N_17788,N_16194);
or U23842 (N_23842,N_18494,N_15035);
nand U23843 (N_23843,N_18683,N_19382);
and U23844 (N_23844,N_17359,N_16987);
nor U23845 (N_23845,N_17401,N_19965);
xnor U23846 (N_23846,N_17563,N_19664);
and U23847 (N_23847,N_17354,N_19051);
or U23848 (N_23848,N_15686,N_15243);
or U23849 (N_23849,N_17504,N_18289);
nand U23850 (N_23850,N_18459,N_16632);
and U23851 (N_23851,N_16441,N_17880);
or U23852 (N_23852,N_17926,N_18219);
and U23853 (N_23853,N_16636,N_16257);
nand U23854 (N_23854,N_15744,N_18999);
nand U23855 (N_23855,N_15464,N_17229);
nand U23856 (N_23856,N_19106,N_15762);
nor U23857 (N_23857,N_15796,N_18175);
nor U23858 (N_23858,N_18468,N_18411);
and U23859 (N_23859,N_17741,N_17269);
nor U23860 (N_23860,N_16057,N_17444);
nand U23861 (N_23861,N_16404,N_15205);
and U23862 (N_23862,N_18675,N_18038);
nor U23863 (N_23863,N_18097,N_18802);
or U23864 (N_23864,N_17930,N_16613);
and U23865 (N_23865,N_15475,N_18289);
or U23866 (N_23866,N_19427,N_17951);
or U23867 (N_23867,N_17611,N_17345);
and U23868 (N_23868,N_15566,N_19966);
and U23869 (N_23869,N_15610,N_17511);
nand U23870 (N_23870,N_16876,N_15926);
or U23871 (N_23871,N_15103,N_15122);
nor U23872 (N_23872,N_15005,N_17514);
or U23873 (N_23873,N_17116,N_18493);
nor U23874 (N_23874,N_17458,N_19033);
nand U23875 (N_23875,N_17027,N_15825);
nor U23876 (N_23876,N_19598,N_18565);
nor U23877 (N_23877,N_17472,N_15077);
nor U23878 (N_23878,N_19377,N_15382);
and U23879 (N_23879,N_19373,N_19150);
nand U23880 (N_23880,N_16406,N_17150);
or U23881 (N_23881,N_17033,N_16295);
or U23882 (N_23882,N_19875,N_18299);
nor U23883 (N_23883,N_16489,N_15171);
xnor U23884 (N_23884,N_15730,N_18360);
nor U23885 (N_23885,N_15336,N_19973);
and U23886 (N_23886,N_17730,N_19362);
nand U23887 (N_23887,N_17676,N_16527);
or U23888 (N_23888,N_19461,N_18016);
nor U23889 (N_23889,N_18515,N_17476);
or U23890 (N_23890,N_15093,N_15563);
and U23891 (N_23891,N_15299,N_15326);
or U23892 (N_23892,N_15744,N_17806);
and U23893 (N_23893,N_17718,N_16783);
nor U23894 (N_23894,N_19153,N_15896);
or U23895 (N_23895,N_18687,N_15707);
nor U23896 (N_23896,N_16049,N_16093);
nand U23897 (N_23897,N_19331,N_18135);
or U23898 (N_23898,N_19325,N_18483);
nor U23899 (N_23899,N_16572,N_18957);
nand U23900 (N_23900,N_17162,N_15738);
or U23901 (N_23901,N_17293,N_16022);
xor U23902 (N_23902,N_17481,N_19989);
nor U23903 (N_23903,N_19457,N_16193);
and U23904 (N_23904,N_15682,N_19281);
xnor U23905 (N_23905,N_16251,N_16968);
nor U23906 (N_23906,N_18178,N_17691);
nand U23907 (N_23907,N_17628,N_15729);
xor U23908 (N_23908,N_19845,N_17805);
or U23909 (N_23909,N_19119,N_18508);
and U23910 (N_23910,N_19423,N_18196);
or U23911 (N_23911,N_18481,N_15396);
and U23912 (N_23912,N_18154,N_18292);
nand U23913 (N_23913,N_16780,N_16066);
or U23914 (N_23914,N_17905,N_17889);
and U23915 (N_23915,N_16957,N_18059);
nor U23916 (N_23916,N_15330,N_18824);
nor U23917 (N_23917,N_15811,N_17804);
nand U23918 (N_23918,N_18206,N_15881);
or U23919 (N_23919,N_16055,N_15630);
or U23920 (N_23920,N_15324,N_15014);
nor U23921 (N_23921,N_16724,N_16623);
xor U23922 (N_23922,N_17161,N_19802);
nand U23923 (N_23923,N_15018,N_15365);
nand U23924 (N_23924,N_17526,N_17678);
xnor U23925 (N_23925,N_16174,N_18684);
nor U23926 (N_23926,N_16334,N_19882);
and U23927 (N_23927,N_17043,N_19856);
or U23928 (N_23928,N_19489,N_15934);
nand U23929 (N_23929,N_15121,N_16349);
nand U23930 (N_23930,N_18513,N_18518);
nand U23931 (N_23931,N_17052,N_18037);
and U23932 (N_23932,N_16003,N_15962);
nor U23933 (N_23933,N_15672,N_17884);
xnor U23934 (N_23934,N_15058,N_18924);
and U23935 (N_23935,N_19673,N_18951);
or U23936 (N_23936,N_16730,N_19360);
or U23937 (N_23937,N_18408,N_18849);
or U23938 (N_23938,N_16211,N_17964);
and U23939 (N_23939,N_18586,N_16370);
nor U23940 (N_23940,N_17305,N_19627);
or U23941 (N_23941,N_16907,N_19866);
nor U23942 (N_23942,N_19865,N_19521);
or U23943 (N_23943,N_16771,N_15847);
nor U23944 (N_23944,N_15741,N_17951);
nor U23945 (N_23945,N_18110,N_17696);
or U23946 (N_23946,N_16287,N_16295);
or U23947 (N_23947,N_19569,N_15223);
nand U23948 (N_23948,N_15309,N_18544);
or U23949 (N_23949,N_18894,N_19528);
nor U23950 (N_23950,N_18409,N_15298);
and U23951 (N_23951,N_18068,N_15721);
nand U23952 (N_23952,N_17833,N_18754);
nor U23953 (N_23953,N_17343,N_19050);
nand U23954 (N_23954,N_18199,N_16738);
or U23955 (N_23955,N_16387,N_18845);
and U23956 (N_23956,N_19506,N_15424);
nor U23957 (N_23957,N_17031,N_16650);
or U23958 (N_23958,N_19594,N_16079);
nand U23959 (N_23959,N_15830,N_15085);
nand U23960 (N_23960,N_18860,N_17789);
and U23961 (N_23961,N_19819,N_15460);
nand U23962 (N_23962,N_16486,N_15512);
xor U23963 (N_23963,N_16780,N_18934);
nand U23964 (N_23964,N_17700,N_19696);
or U23965 (N_23965,N_19642,N_15253);
and U23966 (N_23966,N_19493,N_19659);
xor U23967 (N_23967,N_15479,N_16749);
or U23968 (N_23968,N_15536,N_16003);
and U23969 (N_23969,N_15546,N_19425);
or U23970 (N_23970,N_19755,N_19459);
nand U23971 (N_23971,N_15858,N_16783);
nor U23972 (N_23972,N_19407,N_18209);
nand U23973 (N_23973,N_15217,N_18194);
or U23974 (N_23974,N_16772,N_17140);
or U23975 (N_23975,N_19622,N_18022);
nor U23976 (N_23976,N_19872,N_17518);
and U23977 (N_23977,N_18107,N_18438);
or U23978 (N_23978,N_16007,N_19429);
nand U23979 (N_23979,N_15468,N_16776);
nand U23980 (N_23980,N_15821,N_19674);
and U23981 (N_23981,N_15258,N_16147);
and U23982 (N_23982,N_16228,N_17803);
and U23983 (N_23983,N_17489,N_18185);
nor U23984 (N_23984,N_15219,N_19268);
nand U23985 (N_23985,N_17278,N_17010);
nor U23986 (N_23986,N_16934,N_18675);
nand U23987 (N_23987,N_16955,N_19843);
or U23988 (N_23988,N_18038,N_19409);
xnor U23989 (N_23989,N_19702,N_18356);
nand U23990 (N_23990,N_17096,N_15149);
or U23991 (N_23991,N_16801,N_16661);
nand U23992 (N_23992,N_16383,N_17406);
or U23993 (N_23993,N_19183,N_17707);
and U23994 (N_23994,N_16026,N_18941);
or U23995 (N_23995,N_17354,N_17410);
and U23996 (N_23996,N_18673,N_15362);
or U23997 (N_23997,N_17849,N_17223);
nand U23998 (N_23998,N_15205,N_19594);
and U23999 (N_23999,N_19432,N_17812);
xor U24000 (N_24000,N_16569,N_19974);
or U24001 (N_24001,N_19908,N_17071);
nand U24002 (N_24002,N_17255,N_16718);
and U24003 (N_24003,N_16672,N_18664);
or U24004 (N_24004,N_16399,N_19095);
or U24005 (N_24005,N_15070,N_19292);
nand U24006 (N_24006,N_16974,N_18948);
and U24007 (N_24007,N_19704,N_19063);
xor U24008 (N_24008,N_19116,N_16436);
and U24009 (N_24009,N_15362,N_16546);
xnor U24010 (N_24010,N_17366,N_17284);
and U24011 (N_24011,N_18193,N_18077);
or U24012 (N_24012,N_17491,N_16196);
or U24013 (N_24013,N_17176,N_16234);
nor U24014 (N_24014,N_15252,N_19045);
nand U24015 (N_24015,N_19697,N_18258);
nand U24016 (N_24016,N_19669,N_15197);
and U24017 (N_24017,N_19037,N_16686);
nor U24018 (N_24018,N_18714,N_18724);
or U24019 (N_24019,N_16040,N_16706);
nand U24020 (N_24020,N_17120,N_16650);
xor U24021 (N_24021,N_17279,N_18969);
or U24022 (N_24022,N_19515,N_19360);
xor U24023 (N_24023,N_16935,N_16439);
and U24024 (N_24024,N_19876,N_18092);
nand U24025 (N_24025,N_18384,N_18278);
nand U24026 (N_24026,N_17353,N_17752);
or U24027 (N_24027,N_17133,N_16842);
nand U24028 (N_24028,N_19264,N_15042);
xnor U24029 (N_24029,N_19084,N_15175);
nor U24030 (N_24030,N_19679,N_17289);
and U24031 (N_24031,N_15607,N_19768);
and U24032 (N_24032,N_18024,N_19324);
xor U24033 (N_24033,N_15025,N_18445);
or U24034 (N_24034,N_19909,N_15817);
xor U24035 (N_24035,N_16936,N_15934);
and U24036 (N_24036,N_16513,N_18659);
or U24037 (N_24037,N_15268,N_18067);
nor U24038 (N_24038,N_17621,N_15372);
nor U24039 (N_24039,N_16230,N_19860);
nand U24040 (N_24040,N_18746,N_15672);
nand U24041 (N_24041,N_18545,N_17811);
and U24042 (N_24042,N_17920,N_15028);
nand U24043 (N_24043,N_19919,N_18924);
and U24044 (N_24044,N_15995,N_18659);
nor U24045 (N_24045,N_16209,N_15387);
nor U24046 (N_24046,N_18006,N_16386);
nor U24047 (N_24047,N_15728,N_19940);
and U24048 (N_24048,N_19843,N_19309);
nor U24049 (N_24049,N_15587,N_17589);
and U24050 (N_24050,N_15350,N_16993);
nor U24051 (N_24051,N_19760,N_15583);
xnor U24052 (N_24052,N_17402,N_15193);
nor U24053 (N_24053,N_18761,N_16770);
nor U24054 (N_24054,N_16048,N_15486);
nand U24055 (N_24055,N_15092,N_18482);
nor U24056 (N_24056,N_19916,N_16529);
or U24057 (N_24057,N_16632,N_16920);
or U24058 (N_24058,N_17647,N_16370);
nand U24059 (N_24059,N_15268,N_18508);
nor U24060 (N_24060,N_15490,N_15008);
nand U24061 (N_24061,N_15699,N_18079);
and U24062 (N_24062,N_15690,N_15609);
nor U24063 (N_24063,N_17423,N_19479);
and U24064 (N_24064,N_18780,N_15718);
and U24065 (N_24065,N_18256,N_15000);
or U24066 (N_24066,N_17883,N_17015);
or U24067 (N_24067,N_18966,N_16718);
nand U24068 (N_24068,N_17341,N_15649);
or U24069 (N_24069,N_15927,N_19541);
or U24070 (N_24070,N_19106,N_15008);
nor U24071 (N_24071,N_16596,N_17504);
and U24072 (N_24072,N_18824,N_18358);
nand U24073 (N_24073,N_18946,N_15848);
nand U24074 (N_24074,N_17135,N_18585);
nand U24075 (N_24075,N_15116,N_16920);
or U24076 (N_24076,N_15949,N_18607);
xnor U24077 (N_24077,N_18240,N_18870);
and U24078 (N_24078,N_19108,N_15568);
nand U24079 (N_24079,N_15277,N_15823);
nor U24080 (N_24080,N_15363,N_18615);
and U24081 (N_24081,N_18068,N_18912);
nand U24082 (N_24082,N_19918,N_18565);
and U24083 (N_24083,N_19722,N_16849);
nor U24084 (N_24084,N_16341,N_17542);
nand U24085 (N_24085,N_17658,N_17117);
and U24086 (N_24086,N_19930,N_18145);
and U24087 (N_24087,N_16911,N_17225);
and U24088 (N_24088,N_17747,N_15802);
nor U24089 (N_24089,N_16763,N_19408);
and U24090 (N_24090,N_19801,N_18859);
or U24091 (N_24091,N_19620,N_19103);
nor U24092 (N_24092,N_17521,N_15903);
nor U24093 (N_24093,N_16973,N_15348);
and U24094 (N_24094,N_17617,N_15051);
and U24095 (N_24095,N_17398,N_15189);
nand U24096 (N_24096,N_16927,N_19882);
nor U24097 (N_24097,N_16518,N_18443);
or U24098 (N_24098,N_15782,N_18963);
nand U24099 (N_24099,N_15253,N_19945);
nand U24100 (N_24100,N_15528,N_17429);
nor U24101 (N_24101,N_15053,N_16702);
or U24102 (N_24102,N_16267,N_18171);
or U24103 (N_24103,N_19570,N_18309);
nand U24104 (N_24104,N_16564,N_19467);
xor U24105 (N_24105,N_19641,N_19990);
and U24106 (N_24106,N_15757,N_18048);
nand U24107 (N_24107,N_16240,N_17834);
nor U24108 (N_24108,N_17689,N_17184);
and U24109 (N_24109,N_17916,N_15928);
or U24110 (N_24110,N_16370,N_16430);
and U24111 (N_24111,N_17074,N_15469);
xnor U24112 (N_24112,N_18525,N_17788);
nor U24113 (N_24113,N_18180,N_18641);
nand U24114 (N_24114,N_18513,N_16461);
nor U24115 (N_24115,N_17985,N_16840);
or U24116 (N_24116,N_17769,N_16462);
and U24117 (N_24117,N_19650,N_16625);
or U24118 (N_24118,N_16272,N_19763);
and U24119 (N_24119,N_15844,N_19277);
and U24120 (N_24120,N_16537,N_17363);
nor U24121 (N_24121,N_18940,N_19730);
or U24122 (N_24122,N_18012,N_19830);
and U24123 (N_24123,N_15818,N_18653);
nor U24124 (N_24124,N_16062,N_16530);
or U24125 (N_24125,N_18626,N_16162);
xor U24126 (N_24126,N_16012,N_16929);
and U24127 (N_24127,N_18646,N_16732);
or U24128 (N_24128,N_18212,N_16922);
and U24129 (N_24129,N_18594,N_18870);
nand U24130 (N_24130,N_15121,N_16890);
nand U24131 (N_24131,N_18897,N_18711);
or U24132 (N_24132,N_19439,N_19790);
and U24133 (N_24133,N_17385,N_19739);
and U24134 (N_24134,N_16708,N_18009);
nand U24135 (N_24135,N_19049,N_19312);
and U24136 (N_24136,N_18180,N_15489);
and U24137 (N_24137,N_19773,N_15840);
nand U24138 (N_24138,N_15485,N_17262);
and U24139 (N_24139,N_19175,N_16290);
nand U24140 (N_24140,N_17283,N_19064);
and U24141 (N_24141,N_18498,N_18162);
or U24142 (N_24142,N_15432,N_19666);
and U24143 (N_24143,N_18532,N_15581);
and U24144 (N_24144,N_17039,N_19938);
and U24145 (N_24145,N_19718,N_19903);
or U24146 (N_24146,N_15026,N_19461);
nand U24147 (N_24147,N_19947,N_17845);
xnor U24148 (N_24148,N_18739,N_15709);
nor U24149 (N_24149,N_18972,N_19704);
nor U24150 (N_24150,N_18808,N_19143);
nor U24151 (N_24151,N_15049,N_18814);
xor U24152 (N_24152,N_17491,N_19182);
xnor U24153 (N_24153,N_19791,N_19484);
or U24154 (N_24154,N_15747,N_16189);
nor U24155 (N_24155,N_16160,N_17856);
xnor U24156 (N_24156,N_19996,N_18801);
xnor U24157 (N_24157,N_18855,N_16856);
nand U24158 (N_24158,N_18226,N_17120);
xor U24159 (N_24159,N_19930,N_16021);
and U24160 (N_24160,N_17623,N_16715);
nand U24161 (N_24161,N_16620,N_17817);
and U24162 (N_24162,N_17875,N_17376);
nor U24163 (N_24163,N_18069,N_17808);
nand U24164 (N_24164,N_15110,N_16919);
or U24165 (N_24165,N_18710,N_16914);
nor U24166 (N_24166,N_18881,N_17036);
or U24167 (N_24167,N_15416,N_18299);
and U24168 (N_24168,N_16651,N_18374);
or U24169 (N_24169,N_17331,N_17638);
nand U24170 (N_24170,N_15534,N_17852);
nor U24171 (N_24171,N_17117,N_18457);
xor U24172 (N_24172,N_19982,N_19053);
nand U24173 (N_24173,N_16495,N_19670);
nor U24174 (N_24174,N_17666,N_17225);
and U24175 (N_24175,N_16408,N_19730);
nand U24176 (N_24176,N_15673,N_17849);
nand U24177 (N_24177,N_17430,N_18783);
or U24178 (N_24178,N_17698,N_18852);
xor U24179 (N_24179,N_16927,N_17704);
nand U24180 (N_24180,N_17878,N_18090);
nand U24181 (N_24181,N_18999,N_17637);
nor U24182 (N_24182,N_15183,N_19306);
and U24183 (N_24183,N_16657,N_18533);
or U24184 (N_24184,N_18514,N_19817);
and U24185 (N_24185,N_17294,N_19968);
and U24186 (N_24186,N_15626,N_18035);
nor U24187 (N_24187,N_16994,N_17522);
nand U24188 (N_24188,N_18114,N_16990);
xnor U24189 (N_24189,N_15662,N_18346);
nor U24190 (N_24190,N_18504,N_19033);
or U24191 (N_24191,N_18320,N_15442);
or U24192 (N_24192,N_15544,N_16746);
or U24193 (N_24193,N_15774,N_17754);
nand U24194 (N_24194,N_18195,N_18376);
and U24195 (N_24195,N_19319,N_17208);
nand U24196 (N_24196,N_15968,N_15169);
or U24197 (N_24197,N_15087,N_15641);
or U24198 (N_24198,N_15631,N_19195);
or U24199 (N_24199,N_18269,N_17144);
nor U24200 (N_24200,N_15480,N_15295);
nand U24201 (N_24201,N_18497,N_19874);
or U24202 (N_24202,N_18148,N_17940);
and U24203 (N_24203,N_19142,N_15392);
nor U24204 (N_24204,N_19046,N_15073);
and U24205 (N_24205,N_17877,N_15011);
and U24206 (N_24206,N_18034,N_15411);
or U24207 (N_24207,N_17911,N_17256);
and U24208 (N_24208,N_15068,N_19842);
nand U24209 (N_24209,N_15086,N_18238);
xnor U24210 (N_24210,N_15786,N_19843);
and U24211 (N_24211,N_18924,N_17185);
or U24212 (N_24212,N_18647,N_16774);
nor U24213 (N_24213,N_17041,N_19575);
nor U24214 (N_24214,N_19093,N_19563);
nor U24215 (N_24215,N_15985,N_17396);
nor U24216 (N_24216,N_15181,N_15583);
and U24217 (N_24217,N_17037,N_18980);
or U24218 (N_24218,N_19886,N_17452);
nand U24219 (N_24219,N_16073,N_19874);
xor U24220 (N_24220,N_18037,N_19149);
and U24221 (N_24221,N_16266,N_18758);
nor U24222 (N_24222,N_17675,N_18326);
and U24223 (N_24223,N_19459,N_17261);
and U24224 (N_24224,N_18424,N_18467);
nand U24225 (N_24225,N_15916,N_19610);
nor U24226 (N_24226,N_15981,N_18874);
or U24227 (N_24227,N_16390,N_17699);
nand U24228 (N_24228,N_18295,N_16678);
xor U24229 (N_24229,N_17649,N_15309);
or U24230 (N_24230,N_16614,N_18880);
and U24231 (N_24231,N_15678,N_18517);
nor U24232 (N_24232,N_17125,N_19680);
or U24233 (N_24233,N_17082,N_17492);
and U24234 (N_24234,N_19703,N_15049);
or U24235 (N_24235,N_18019,N_16941);
and U24236 (N_24236,N_16743,N_18085);
and U24237 (N_24237,N_17376,N_19967);
or U24238 (N_24238,N_19948,N_16877);
and U24239 (N_24239,N_15710,N_16217);
or U24240 (N_24240,N_17348,N_16158);
or U24241 (N_24241,N_16653,N_15579);
nand U24242 (N_24242,N_15731,N_18709);
xnor U24243 (N_24243,N_16405,N_19996);
and U24244 (N_24244,N_15519,N_16045);
nand U24245 (N_24245,N_15583,N_18904);
and U24246 (N_24246,N_17708,N_17681);
and U24247 (N_24247,N_17944,N_15025);
nand U24248 (N_24248,N_18886,N_16512);
and U24249 (N_24249,N_15995,N_15675);
and U24250 (N_24250,N_15477,N_17023);
or U24251 (N_24251,N_16295,N_16263);
xor U24252 (N_24252,N_19456,N_15167);
and U24253 (N_24253,N_15397,N_19467);
and U24254 (N_24254,N_16393,N_17165);
xnor U24255 (N_24255,N_16715,N_16096);
and U24256 (N_24256,N_18995,N_18843);
and U24257 (N_24257,N_17043,N_19549);
or U24258 (N_24258,N_19414,N_15394);
nor U24259 (N_24259,N_17864,N_16400);
or U24260 (N_24260,N_17573,N_18774);
xnor U24261 (N_24261,N_19841,N_19647);
and U24262 (N_24262,N_16687,N_19556);
xor U24263 (N_24263,N_17645,N_18520);
nand U24264 (N_24264,N_17641,N_15045);
nor U24265 (N_24265,N_19762,N_19437);
and U24266 (N_24266,N_15637,N_15718);
nor U24267 (N_24267,N_17577,N_19663);
xnor U24268 (N_24268,N_16484,N_17172);
or U24269 (N_24269,N_19155,N_15533);
nand U24270 (N_24270,N_15022,N_18951);
or U24271 (N_24271,N_16693,N_16109);
nor U24272 (N_24272,N_16969,N_15004);
or U24273 (N_24273,N_17867,N_17968);
and U24274 (N_24274,N_19903,N_15059);
nor U24275 (N_24275,N_18554,N_16216);
or U24276 (N_24276,N_16179,N_17642);
or U24277 (N_24277,N_19958,N_15980);
and U24278 (N_24278,N_19250,N_17828);
or U24279 (N_24279,N_17609,N_17054);
nor U24280 (N_24280,N_15793,N_18140);
nor U24281 (N_24281,N_16381,N_18356);
nand U24282 (N_24282,N_16702,N_18511);
xnor U24283 (N_24283,N_17056,N_16278);
and U24284 (N_24284,N_18090,N_17645);
nand U24285 (N_24285,N_15801,N_15697);
and U24286 (N_24286,N_18189,N_18633);
and U24287 (N_24287,N_18833,N_16518);
nor U24288 (N_24288,N_15911,N_16788);
or U24289 (N_24289,N_16205,N_19900);
xnor U24290 (N_24290,N_19596,N_17798);
or U24291 (N_24291,N_18034,N_17785);
nand U24292 (N_24292,N_18481,N_19166);
nand U24293 (N_24293,N_15388,N_15397);
and U24294 (N_24294,N_17867,N_16852);
nand U24295 (N_24295,N_17056,N_15696);
or U24296 (N_24296,N_19200,N_17931);
nand U24297 (N_24297,N_15303,N_17030);
and U24298 (N_24298,N_17830,N_17602);
nand U24299 (N_24299,N_17285,N_19204);
and U24300 (N_24300,N_17625,N_19567);
and U24301 (N_24301,N_15174,N_15737);
or U24302 (N_24302,N_19600,N_19454);
and U24303 (N_24303,N_18746,N_15654);
and U24304 (N_24304,N_17178,N_15495);
nand U24305 (N_24305,N_18819,N_19492);
nor U24306 (N_24306,N_15345,N_16648);
nand U24307 (N_24307,N_16311,N_18889);
and U24308 (N_24308,N_19033,N_19855);
or U24309 (N_24309,N_16148,N_15241);
nand U24310 (N_24310,N_19578,N_19429);
nand U24311 (N_24311,N_19318,N_17637);
nand U24312 (N_24312,N_16562,N_17699);
nor U24313 (N_24313,N_18879,N_16513);
nand U24314 (N_24314,N_16792,N_18652);
or U24315 (N_24315,N_18920,N_16695);
or U24316 (N_24316,N_16860,N_19972);
or U24317 (N_24317,N_15358,N_15620);
or U24318 (N_24318,N_15363,N_18083);
and U24319 (N_24319,N_15382,N_17435);
or U24320 (N_24320,N_18304,N_16917);
nand U24321 (N_24321,N_15006,N_17849);
or U24322 (N_24322,N_17063,N_16232);
and U24323 (N_24323,N_19530,N_17262);
and U24324 (N_24324,N_19663,N_19044);
nor U24325 (N_24325,N_19609,N_17131);
and U24326 (N_24326,N_16697,N_18711);
nor U24327 (N_24327,N_15944,N_16711);
and U24328 (N_24328,N_18691,N_18804);
nor U24329 (N_24329,N_19155,N_15398);
nor U24330 (N_24330,N_15147,N_18372);
nor U24331 (N_24331,N_19356,N_16951);
and U24332 (N_24332,N_19465,N_17721);
nand U24333 (N_24333,N_19713,N_16497);
and U24334 (N_24334,N_15706,N_15701);
nor U24335 (N_24335,N_18039,N_18572);
or U24336 (N_24336,N_15297,N_15540);
and U24337 (N_24337,N_16759,N_15686);
nor U24338 (N_24338,N_16461,N_19604);
nand U24339 (N_24339,N_16516,N_16519);
and U24340 (N_24340,N_17674,N_17816);
xor U24341 (N_24341,N_17843,N_18574);
xor U24342 (N_24342,N_17634,N_17849);
or U24343 (N_24343,N_18262,N_18965);
and U24344 (N_24344,N_19895,N_19773);
nor U24345 (N_24345,N_15550,N_15029);
and U24346 (N_24346,N_17273,N_19370);
nand U24347 (N_24347,N_15626,N_16123);
xor U24348 (N_24348,N_18602,N_19422);
nand U24349 (N_24349,N_15289,N_18513);
nand U24350 (N_24350,N_19614,N_18202);
or U24351 (N_24351,N_15304,N_15916);
or U24352 (N_24352,N_18635,N_18616);
xor U24353 (N_24353,N_15173,N_17791);
nor U24354 (N_24354,N_19142,N_16928);
or U24355 (N_24355,N_16586,N_17214);
and U24356 (N_24356,N_17182,N_16595);
nor U24357 (N_24357,N_15007,N_16324);
and U24358 (N_24358,N_17236,N_19077);
or U24359 (N_24359,N_18508,N_17980);
or U24360 (N_24360,N_16174,N_15472);
nand U24361 (N_24361,N_15079,N_18402);
and U24362 (N_24362,N_16012,N_16913);
nor U24363 (N_24363,N_15808,N_15360);
or U24364 (N_24364,N_17602,N_18718);
and U24365 (N_24365,N_18707,N_17590);
and U24366 (N_24366,N_15701,N_16831);
nand U24367 (N_24367,N_19967,N_18168);
and U24368 (N_24368,N_15666,N_18682);
and U24369 (N_24369,N_18922,N_18218);
or U24370 (N_24370,N_18949,N_16604);
nand U24371 (N_24371,N_19045,N_19349);
or U24372 (N_24372,N_18827,N_19132);
nor U24373 (N_24373,N_15619,N_17668);
nand U24374 (N_24374,N_16888,N_15107);
nand U24375 (N_24375,N_15475,N_17829);
nand U24376 (N_24376,N_16215,N_15866);
or U24377 (N_24377,N_15080,N_19558);
nand U24378 (N_24378,N_19596,N_19167);
or U24379 (N_24379,N_18957,N_16085);
nor U24380 (N_24380,N_19616,N_15426);
or U24381 (N_24381,N_19813,N_17410);
xnor U24382 (N_24382,N_15895,N_16564);
nor U24383 (N_24383,N_17827,N_18386);
or U24384 (N_24384,N_15235,N_16649);
or U24385 (N_24385,N_19018,N_17325);
and U24386 (N_24386,N_16348,N_19095);
nand U24387 (N_24387,N_16574,N_19808);
nor U24388 (N_24388,N_15110,N_16502);
nand U24389 (N_24389,N_17027,N_15269);
nor U24390 (N_24390,N_18171,N_15503);
xnor U24391 (N_24391,N_19604,N_16480);
nor U24392 (N_24392,N_16243,N_15703);
nand U24393 (N_24393,N_17562,N_19081);
and U24394 (N_24394,N_17072,N_17361);
nor U24395 (N_24395,N_16480,N_15367);
nor U24396 (N_24396,N_19745,N_19877);
nand U24397 (N_24397,N_19862,N_18999);
nand U24398 (N_24398,N_17677,N_19188);
or U24399 (N_24399,N_15628,N_16703);
or U24400 (N_24400,N_18459,N_16220);
and U24401 (N_24401,N_19740,N_16964);
xnor U24402 (N_24402,N_16061,N_19685);
nand U24403 (N_24403,N_17631,N_19206);
nand U24404 (N_24404,N_15973,N_15461);
xnor U24405 (N_24405,N_15309,N_18358);
or U24406 (N_24406,N_17751,N_17637);
nand U24407 (N_24407,N_19744,N_19902);
or U24408 (N_24408,N_19078,N_15114);
or U24409 (N_24409,N_19777,N_17169);
nor U24410 (N_24410,N_15107,N_16051);
or U24411 (N_24411,N_17110,N_17835);
and U24412 (N_24412,N_19980,N_18381);
and U24413 (N_24413,N_17910,N_19879);
or U24414 (N_24414,N_16310,N_17611);
xor U24415 (N_24415,N_15388,N_15389);
or U24416 (N_24416,N_18240,N_19662);
and U24417 (N_24417,N_16179,N_15094);
or U24418 (N_24418,N_19294,N_18256);
or U24419 (N_24419,N_15114,N_17918);
or U24420 (N_24420,N_19402,N_17294);
and U24421 (N_24421,N_18658,N_19321);
nor U24422 (N_24422,N_15561,N_15959);
nand U24423 (N_24423,N_16294,N_17096);
nand U24424 (N_24424,N_15600,N_18269);
or U24425 (N_24425,N_17469,N_17229);
nand U24426 (N_24426,N_19526,N_15758);
or U24427 (N_24427,N_17827,N_17708);
and U24428 (N_24428,N_15942,N_18435);
or U24429 (N_24429,N_19519,N_16745);
and U24430 (N_24430,N_19132,N_19735);
nand U24431 (N_24431,N_15671,N_16506);
and U24432 (N_24432,N_18724,N_15163);
and U24433 (N_24433,N_15124,N_17968);
nor U24434 (N_24434,N_17905,N_15333);
nor U24435 (N_24435,N_18318,N_16213);
xnor U24436 (N_24436,N_18247,N_19342);
nor U24437 (N_24437,N_18768,N_15411);
xnor U24438 (N_24438,N_15845,N_16516);
nor U24439 (N_24439,N_18563,N_16183);
and U24440 (N_24440,N_15376,N_18386);
nor U24441 (N_24441,N_16064,N_16873);
and U24442 (N_24442,N_18123,N_15572);
nand U24443 (N_24443,N_15949,N_15233);
or U24444 (N_24444,N_15913,N_18791);
and U24445 (N_24445,N_19435,N_18024);
nand U24446 (N_24446,N_18326,N_17937);
nand U24447 (N_24447,N_17562,N_16568);
nor U24448 (N_24448,N_15626,N_15333);
nand U24449 (N_24449,N_16934,N_15594);
nand U24450 (N_24450,N_18845,N_15338);
and U24451 (N_24451,N_19091,N_16885);
or U24452 (N_24452,N_17957,N_18502);
xnor U24453 (N_24453,N_18073,N_18501);
or U24454 (N_24454,N_16008,N_17244);
nand U24455 (N_24455,N_18180,N_15370);
nor U24456 (N_24456,N_19575,N_15294);
and U24457 (N_24457,N_17087,N_15539);
or U24458 (N_24458,N_17058,N_17917);
and U24459 (N_24459,N_18756,N_17010);
nand U24460 (N_24460,N_18259,N_19450);
and U24461 (N_24461,N_17197,N_19360);
xnor U24462 (N_24462,N_17617,N_16525);
nand U24463 (N_24463,N_19275,N_16472);
nor U24464 (N_24464,N_17559,N_19649);
nor U24465 (N_24465,N_15535,N_19452);
and U24466 (N_24466,N_19600,N_18050);
nand U24467 (N_24467,N_18180,N_15083);
nand U24468 (N_24468,N_16953,N_18672);
and U24469 (N_24469,N_15929,N_17015);
or U24470 (N_24470,N_15330,N_19513);
xnor U24471 (N_24471,N_16550,N_15292);
and U24472 (N_24472,N_17889,N_17906);
xor U24473 (N_24473,N_18083,N_15863);
or U24474 (N_24474,N_15095,N_19893);
nor U24475 (N_24475,N_15578,N_19677);
and U24476 (N_24476,N_16311,N_15599);
or U24477 (N_24477,N_17902,N_16719);
and U24478 (N_24478,N_15184,N_15213);
nand U24479 (N_24479,N_18125,N_17170);
and U24480 (N_24480,N_17882,N_18620);
xor U24481 (N_24481,N_17810,N_15228);
nor U24482 (N_24482,N_18135,N_16111);
and U24483 (N_24483,N_16623,N_16799);
or U24484 (N_24484,N_16013,N_19659);
or U24485 (N_24485,N_19943,N_19391);
nand U24486 (N_24486,N_16072,N_17675);
nor U24487 (N_24487,N_16076,N_15448);
nand U24488 (N_24488,N_18190,N_15952);
nand U24489 (N_24489,N_17210,N_15181);
nand U24490 (N_24490,N_15919,N_18087);
or U24491 (N_24491,N_15305,N_17515);
nor U24492 (N_24492,N_19562,N_19623);
and U24493 (N_24493,N_17591,N_18567);
and U24494 (N_24494,N_16191,N_19821);
nand U24495 (N_24495,N_16727,N_16966);
and U24496 (N_24496,N_15366,N_18188);
and U24497 (N_24497,N_18531,N_19037);
or U24498 (N_24498,N_19455,N_18102);
nand U24499 (N_24499,N_18449,N_17555);
and U24500 (N_24500,N_19879,N_15596);
or U24501 (N_24501,N_19787,N_19676);
or U24502 (N_24502,N_17284,N_17638);
nand U24503 (N_24503,N_17351,N_17061);
nand U24504 (N_24504,N_15449,N_17295);
nand U24505 (N_24505,N_16768,N_16401);
or U24506 (N_24506,N_15527,N_19457);
xnor U24507 (N_24507,N_18001,N_17528);
and U24508 (N_24508,N_17032,N_17579);
nand U24509 (N_24509,N_19918,N_17256);
nand U24510 (N_24510,N_17595,N_15651);
nand U24511 (N_24511,N_17549,N_15204);
nor U24512 (N_24512,N_17633,N_15544);
xnor U24513 (N_24513,N_15017,N_18886);
or U24514 (N_24514,N_18593,N_18401);
or U24515 (N_24515,N_19076,N_15383);
nand U24516 (N_24516,N_17183,N_15845);
nand U24517 (N_24517,N_18791,N_15285);
nor U24518 (N_24518,N_19954,N_18159);
nor U24519 (N_24519,N_18702,N_19864);
or U24520 (N_24520,N_19415,N_15551);
or U24521 (N_24521,N_16391,N_15026);
xnor U24522 (N_24522,N_17987,N_19203);
xnor U24523 (N_24523,N_19732,N_18820);
nor U24524 (N_24524,N_16644,N_18341);
and U24525 (N_24525,N_17629,N_17439);
and U24526 (N_24526,N_18663,N_16822);
nand U24527 (N_24527,N_16850,N_15162);
and U24528 (N_24528,N_18670,N_15752);
or U24529 (N_24529,N_19168,N_18780);
nand U24530 (N_24530,N_17457,N_18166);
and U24531 (N_24531,N_15231,N_19782);
nor U24532 (N_24532,N_16625,N_19802);
or U24533 (N_24533,N_15718,N_18722);
nand U24534 (N_24534,N_16653,N_19694);
or U24535 (N_24535,N_19871,N_17838);
xnor U24536 (N_24536,N_17314,N_18891);
and U24537 (N_24537,N_18539,N_17807);
nor U24538 (N_24538,N_17592,N_18346);
and U24539 (N_24539,N_18288,N_15905);
or U24540 (N_24540,N_19711,N_18801);
nand U24541 (N_24541,N_15946,N_18489);
xor U24542 (N_24542,N_19496,N_19948);
and U24543 (N_24543,N_16117,N_15735);
nand U24544 (N_24544,N_15506,N_19511);
nand U24545 (N_24545,N_17884,N_19749);
nor U24546 (N_24546,N_17002,N_17854);
or U24547 (N_24547,N_19318,N_15221);
and U24548 (N_24548,N_16882,N_16970);
nand U24549 (N_24549,N_18738,N_18191);
nor U24550 (N_24550,N_18165,N_18564);
or U24551 (N_24551,N_16202,N_16601);
nand U24552 (N_24552,N_15403,N_15305);
nand U24553 (N_24553,N_18525,N_15904);
nand U24554 (N_24554,N_15866,N_16884);
and U24555 (N_24555,N_16589,N_19403);
or U24556 (N_24556,N_17327,N_18040);
and U24557 (N_24557,N_19872,N_16238);
or U24558 (N_24558,N_16450,N_19661);
nand U24559 (N_24559,N_15098,N_19906);
nand U24560 (N_24560,N_19286,N_19387);
or U24561 (N_24561,N_19719,N_18446);
nand U24562 (N_24562,N_18035,N_18298);
xor U24563 (N_24563,N_16557,N_15579);
nor U24564 (N_24564,N_19474,N_18785);
or U24565 (N_24565,N_15254,N_17207);
nor U24566 (N_24566,N_18990,N_15557);
or U24567 (N_24567,N_18298,N_19397);
nor U24568 (N_24568,N_16714,N_15412);
xor U24569 (N_24569,N_19628,N_18174);
xnor U24570 (N_24570,N_16511,N_15646);
nand U24571 (N_24571,N_17724,N_18827);
or U24572 (N_24572,N_16587,N_19984);
nand U24573 (N_24573,N_18100,N_18847);
nand U24574 (N_24574,N_18329,N_18234);
and U24575 (N_24575,N_17574,N_15591);
or U24576 (N_24576,N_19984,N_15144);
and U24577 (N_24577,N_16202,N_19568);
nand U24578 (N_24578,N_16885,N_18188);
nor U24579 (N_24579,N_19744,N_18999);
nand U24580 (N_24580,N_16281,N_19588);
nand U24581 (N_24581,N_16161,N_19193);
nand U24582 (N_24582,N_19719,N_19591);
nor U24583 (N_24583,N_17229,N_15456);
and U24584 (N_24584,N_17051,N_19913);
nand U24585 (N_24585,N_18288,N_15211);
and U24586 (N_24586,N_18353,N_16708);
nor U24587 (N_24587,N_17129,N_19462);
nor U24588 (N_24588,N_16266,N_16052);
nor U24589 (N_24589,N_18067,N_17369);
xnor U24590 (N_24590,N_19789,N_15257);
xnor U24591 (N_24591,N_15168,N_15031);
or U24592 (N_24592,N_18367,N_15393);
xor U24593 (N_24593,N_19289,N_16108);
nand U24594 (N_24594,N_17043,N_18412);
and U24595 (N_24595,N_18998,N_18274);
nor U24596 (N_24596,N_18536,N_18057);
nor U24597 (N_24597,N_18005,N_18300);
nor U24598 (N_24598,N_19170,N_19606);
xnor U24599 (N_24599,N_17714,N_15190);
xor U24600 (N_24600,N_16843,N_15299);
xnor U24601 (N_24601,N_17350,N_18110);
nor U24602 (N_24602,N_16087,N_15423);
or U24603 (N_24603,N_16078,N_16543);
nor U24604 (N_24604,N_19591,N_19748);
xor U24605 (N_24605,N_18613,N_16485);
or U24606 (N_24606,N_19171,N_15560);
or U24607 (N_24607,N_16458,N_17457);
and U24608 (N_24608,N_17615,N_17002);
nor U24609 (N_24609,N_17000,N_18813);
and U24610 (N_24610,N_18071,N_17229);
nor U24611 (N_24611,N_19409,N_18571);
nor U24612 (N_24612,N_19784,N_15324);
or U24613 (N_24613,N_18303,N_15634);
nand U24614 (N_24614,N_19220,N_17943);
and U24615 (N_24615,N_19149,N_15972);
nor U24616 (N_24616,N_16841,N_17493);
nand U24617 (N_24617,N_18707,N_16408);
nand U24618 (N_24618,N_15844,N_15864);
nand U24619 (N_24619,N_19170,N_16421);
xnor U24620 (N_24620,N_19589,N_15871);
nand U24621 (N_24621,N_17973,N_17149);
nor U24622 (N_24622,N_16350,N_18784);
or U24623 (N_24623,N_16342,N_19719);
nor U24624 (N_24624,N_17166,N_15376);
nand U24625 (N_24625,N_16737,N_17747);
nor U24626 (N_24626,N_16985,N_15492);
nor U24627 (N_24627,N_19817,N_18028);
nor U24628 (N_24628,N_15073,N_17892);
nand U24629 (N_24629,N_16032,N_18706);
or U24630 (N_24630,N_18909,N_17416);
or U24631 (N_24631,N_16370,N_19556);
nor U24632 (N_24632,N_16411,N_17825);
xor U24633 (N_24633,N_15973,N_15437);
or U24634 (N_24634,N_19403,N_19176);
or U24635 (N_24635,N_19199,N_15043);
or U24636 (N_24636,N_15659,N_15704);
nor U24637 (N_24637,N_15567,N_19162);
and U24638 (N_24638,N_15460,N_15674);
or U24639 (N_24639,N_15467,N_18721);
nand U24640 (N_24640,N_17943,N_15620);
nand U24641 (N_24641,N_16708,N_15512);
nor U24642 (N_24642,N_19055,N_18942);
and U24643 (N_24643,N_19892,N_17575);
and U24644 (N_24644,N_17650,N_18566);
xnor U24645 (N_24645,N_19605,N_19281);
nor U24646 (N_24646,N_19673,N_15408);
or U24647 (N_24647,N_18502,N_18740);
nand U24648 (N_24648,N_16005,N_15257);
nand U24649 (N_24649,N_18137,N_19320);
or U24650 (N_24650,N_15420,N_17075);
nand U24651 (N_24651,N_18798,N_15518);
nand U24652 (N_24652,N_17922,N_17566);
or U24653 (N_24653,N_16178,N_19666);
nor U24654 (N_24654,N_19600,N_18051);
nor U24655 (N_24655,N_17997,N_16217);
nand U24656 (N_24656,N_16961,N_15289);
and U24657 (N_24657,N_15437,N_19219);
nand U24658 (N_24658,N_15006,N_19483);
nand U24659 (N_24659,N_16329,N_17375);
nor U24660 (N_24660,N_17860,N_17709);
nor U24661 (N_24661,N_16652,N_17542);
or U24662 (N_24662,N_18936,N_19754);
or U24663 (N_24663,N_17653,N_17316);
nor U24664 (N_24664,N_16893,N_18975);
and U24665 (N_24665,N_16909,N_19112);
nor U24666 (N_24666,N_15119,N_18644);
nor U24667 (N_24667,N_17815,N_17265);
xnor U24668 (N_24668,N_18206,N_16483);
or U24669 (N_24669,N_17466,N_15186);
nor U24670 (N_24670,N_18291,N_15374);
nor U24671 (N_24671,N_17636,N_17660);
xnor U24672 (N_24672,N_18446,N_17509);
and U24673 (N_24673,N_19721,N_19386);
nor U24674 (N_24674,N_18684,N_19080);
and U24675 (N_24675,N_18757,N_17800);
xor U24676 (N_24676,N_19917,N_18811);
nor U24677 (N_24677,N_16238,N_15053);
nor U24678 (N_24678,N_16854,N_17593);
or U24679 (N_24679,N_17224,N_15059);
nand U24680 (N_24680,N_18855,N_17538);
and U24681 (N_24681,N_18827,N_16152);
or U24682 (N_24682,N_17664,N_18681);
nor U24683 (N_24683,N_17195,N_19537);
or U24684 (N_24684,N_17597,N_19183);
and U24685 (N_24685,N_18629,N_18618);
xor U24686 (N_24686,N_18375,N_17816);
xor U24687 (N_24687,N_18540,N_16201);
or U24688 (N_24688,N_15287,N_19962);
nor U24689 (N_24689,N_17197,N_16708);
nor U24690 (N_24690,N_16384,N_16007);
or U24691 (N_24691,N_15787,N_17046);
xnor U24692 (N_24692,N_16447,N_19162);
nor U24693 (N_24693,N_16520,N_17108);
xor U24694 (N_24694,N_17030,N_18698);
xor U24695 (N_24695,N_15756,N_19539);
and U24696 (N_24696,N_16701,N_15587);
and U24697 (N_24697,N_19621,N_18871);
and U24698 (N_24698,N_19481,N_19775);
nor U24699 (N_24699,N_15036,N_16646);
or U24700 (N_24700,N_15598,N_16592);
or U24701 (N_24701,N_17198,N_17241);
or U24702 (N_24702,N_18210,N_15961);
or U24703 (N_24703,N_19495,N_18476);
or U24704 (N_24704,N_15642,N_16242);
or U24705 (N_24705,N_16606,N_16396);
or U24706 (N_24706,N_17860,N_17205);
nand U24707 (N_24707,N_18350,N_17721);
nor U24708 (N_24708,N_16646,N_19767);
xnor U24709 (N_24709,N_15667,N_15933);
xor U24710 (N_24710,N_17543,N_15967);
nor U24711 (N_24711,N_16346,N_17581);
nand U24712 (N_24712,N_16238,N_15514);
xnor U24713 (N_24713,N_17118,N_16488);
xnor U24714 (N_24714,N_18908,N_15563);
nand U24715 (N_24715,N_19185,N_16342);
and U24716 (N_24716,N_17770,N_17279);
nor U24717 (N_24717,N_18440,N_15103);
and U24718 (N_24718,N_17201,N_19585);
nand U24719 (N_24719,N_18960,N_16255);
and U24720 (N_24720,N_19964,N_18322);
and U24721 (N_24721,N_16450,N_15982);
nand U24722 (N_24722,N_15750,N_18151);
and U24723 (N_24723,N_17566,N_17975);
nor U24724 (N_24724,N_18610,N_18648);
xnor U24725 (N_24725,N_16481,N_16715);
xnor U24726 (N_24726,N_16192,N_19756);
nand U24727 (N_24727,N_19722,N_19348);
or U24728 (N_24728,N_17413,N_18926);
nor U24729 (N_24729,N_15575,N_16860);
and U24730 (N_24730,N_16694,N_18095);
nand U24731 (N_24731,N_19998,N_17550);
or U24732 (N_24732,N_17411,N_15867);
nand U24733 (N_24733,N_15021,N_17329);
and U24734 (N_24734,N_17232,N_17789);
or U24735 (N_24735,N_18601,N_19370);
and U24736 (N_24736,N_17693,N_19253);
or U24737 (N_24737,N_17124,N_16359);
nand U24738 (N_24738,N_15513,N_15117);
or U24739 (N_24739,N_19343,N_16143);
nor U24740 (N_24740,N_18116,N_18100);
nand U24741 (N_24741,N_17359,N_17573);
and U24742 (N_24742,N_16066,N_16473);
nor U24743 (N_24743,N_18570,N_15275);
or U24744 (N_24744,N_15311,N_19827);
xnor U24745 (N_24745,N_16517,N_17161);
nand U24746 (N_24746,N_15069,N_16730);
and U24747 (N_24747,N_19309,N_15790);
xor U24748 (N_24748,N_17710,N_18811);
xnor U24749 (N_24749,N_16293,N_19444);
nor U24750 (N_24750,N_16928,N_19759);
and U24751 (N_24751,N_19207,N_15399);
nand U24752 (N_24752,N_19858,N_15718);
or U24753 (N_24753,N_16395,N_19978);
nand U24754 (N_24754,N_15476,N_16227);
and U24755 (N_24755,N_18444,N_19724);
xnor U24756 (N_24756,N_16567,N_15210);
xnor U24757 (N_24757,N_16919,N_17423);
nand U24758 (N_24758,N_18161,N_19971);
or U24759 (N_24759,N_15567,N_17411);
or U24760 (N_24760,N_18755,N_19070);
or U24761 (N_24761,N_18173,N_15101);
nor U24762 (N_24762,N_16531,N_18179);
or U24763 (N_24763,N_16136,N_17307);
nand U24764 (N_24764,N_19886,N_17596);
and U24765 (N_24765,N_15642,N_15616);
nor U24766 (N_24766,N_18544,N_19811);
nand U24767 (N_24767,N_16121,N_17956);
nor U24768 (N_24768,N_18319,N_15799);
nor U24769 (N_24769,N_16348,N_19418);
nand U24770 (N_24770,N_15221,N_17298);
xor U24771 (N_24771,N_17431,N_16306);
nand U24772 (N_24772,N_19394,N_19863);
nand U24773 (N_24773,N_17269,N_18660);
or U24774 (N_24774,N_16742,N_17178);
and U24775 (N_24775,N_15592,N_17133);
and U24776 (N_24776,N_16791,N_17855);
and U24777 (N_24777,N_19959,N_19050);
xor U24778 (N_24778,N_16010,N_17979);
or U24779 (N_24779,N_18365,N_18275);
xnor U24780 (N_24780,N_18815,N_18291);
nor U24781 (N_24781,N_18875,N_16822);
and U24782 (N_24782,N_15382,N_15741);
nand U24783 (N_24783,N_17114,N_16436);
nor U24784 (N_24784,N_16560,N_16293);
and U24785 (N_24785,N_17245,N_19932);
or U24786 (N_24786,N_18061,N_15925);
xor U24787 (N_24787,N_19901,N_17635);
nor U24788 (N_24788,N_15710,N_18021);
nand U24789 (N_24789,N_19491,N_18856);
xor U24790 (N_24790,N_18400,N_16387);
or U24791 (N_24791,N_19760,N_15564);
or U24792 (N_24792,N_17565,N_18947);
and U24793 (N_24793,N_18875,N_18401);
nor U24794 (N_24794,N_18165,N_16546);
or U24795 (N_24795,N_18566,N_19246);
nor U24796 (N_24796,N_17173,N_15966);
or U24797 (N_24797,N_19593,N_19904);
and U24798 (N_24798,N_19025,N_18497);
or U24799 (N_24799,N_16926,N_16145);
nand U24800 (N_24800,N_17729,N_16630);
and U24801 (N_24801,N_18780,N_18056);
nor U24802 (N_24802,N_16575,N_16699);
xnor U24803 (N_24803,N_15515,N_17553);
nor U24804 (N_24804,N_18762,N_18302);
and U24805 (N_24805,N_15647,N_18359);
or U24806 (N_24806,N_18564,N_17847);
and U24807 (N_24807,N_16182,N_15675);
xnor U24808 (N_24808,N_17302,N_18695);
or U24809 (N_24809,N_16118,N_15114);
nor U24810 (N_24810,N_19266,N_19234);
or U24811 (N_24811,N_18888,N_18722);
xnor U24812 (N_24812,N_19769,N_16226);
nor U24813 (N_24813,N_17725,N_19676);
xor U24814 (N_24814,N_15180,N_15315);
and U24815 (N_24815,N_16585,N_16444);
and U24816 (N_24816,N_16086,N_17187);
or U24817 (N_24817,N_19846,N_16590);
and U24818 (N_24818,N_17219,N_17705);
and U24819 (N_24819,N_17677,N_15322);
nand U24820 (N_24820,N_16081,N_16513);
xor U24821 (N_24821,N_17119,N_18914);
nor U24822 (N_24822,N_18848,N_15965);
and U24823 (N_24823,N_17526,N_18098);
and U24824 (N_24824,N_16080,N_15713);
xor U24825 (N_24825,N_17264,N_19099);
or U24826 (N_24826,N_19913,N_16318);
nor U24827 (N_24827,N_17617,N_18884);
and U24828 (N_24828,N_17991,N_18557);
or U24829 (N_24829,N_18768,N_18277);
nor U24830 (N_24830,N_16835,N_15588);
or U24831 (N_24831,N_18333,N_17075);
nor U24832 (N_24832,N_19396,N_17348);
xnor U24833 (N_24833,N_16834,N_15292);
or U24834 (N_24834,N_19003,N_17348);
nand U24835 (N_24835,N_19335,N_19505);
nor U24836 (N_24836,N_15197,N_15027);
or U24837 (N_24837,N_16443,N_17327);
and U24838 (N_24838,N_15250,N_18802);
xnor U24839 (N_24839,N_17904,N_17099);
and U24840 (N_24840,N_16822,N_15448);
and U24841 (N_24841,N_18756,N_19188);
and U24842 (N_24842,N_18693,N_17460);
and U24843 (N_24843,N_19465,N_16869);
nor U24844 (N_24844,N_16553,N_18216);
nand U24845 (N_24845,N_18804,N_18395);
or U24846 (N_24846,N_15817,N_17883);
nor U24847 (N_24847,N_15517,N_16315);
nand U24848 (N_24848,N_17666,N_16452);
nor U24849 (N_24849,N_18574,N_17213);
nand U24850 (N_24850,N_19359,N_19625);
or U24851 (N_24851,N_15845,N_19027);
and U24852 (N_24852,N_15829,N_19942);
nand U24853 (N_24853,N_16387,N_16559);
and U24854 (N_24854,N_19361,N_15112);
nor U24855 (N_24855,N_15474,N_18428);
or U24856 (N_24856,N_15387,N_19137);
or U24857 (N_24857,N_16555,N_16128);
nand U24858 (N_24858,N_15039,N_16527);
xnor U24859 (N_24859,N_16207,N_17441);
nor U24860 (N_24860,N_16099,N_15243);
nor U24861 (N_24861,N_18289,N_18709);
nand U24862 (N_24862,N_16007,N_16544);
nor U24863 (N_24863,N_18901,N_17018);
and U24864 (N_24864,N_16983,N_16848);
nor U24865 (N_24865,N_19906,N_17610);
nand U24866 (N_24866,N_17461,N_18258);
or U24867 (N_24867,N_17886,N_15793);
nand U24868 (N_24868,N_16222,N_19746);
nor U24869 (N_24869,N_16037,N_17889);
nand U24870 (N_24870,N_16137,N_16363);
or U24871 (N_24871,N_19472,N_18687);
or U24872 (N_24872,N_19089,N_17574);
or U24873 (N_24873,N_16189,N_18337);
and U24874 (N_24874,N_17875,N_17537);
and U24875 (N_24875,N_19123,N_15388);
xor U24876 (N_24876,N_16127,N_19307);
and U24877 (N_24877,N_18507,N_15289);
xnor U24878 (N_24878,N_17041,N_18513);
or U24879 (N_24879,N_17898,N_15830);
and U24880 (N_24880,N_19445,N_19598);
and U24881 (N_24881,N_19952,N_17209);
xor U24882 (N_24882,N_17330,N_18090);
and U24883 (N_24883,N_16945,N_16572);
and U24884 (N_24884,N_17710,N_16542);
nor U24885 (N_24885,N_18447,N_19341);
xnor U24886 (N_24886,N_15832,N_17662);
nand U24887 (N_24887,N_15429,N_15303);
nor U24888 (N_24888,N_19931,N_17332);
and U24889 (N_24889,N_17463,N_17514);
nand U24890 (N_24890,N_15797,N_19772);
and U24891 (N_24891,N_15258,N_19701);
nand U24892 (N_24892,N_19128,N_15106);
and U24893 (N_24893,N_17434,N_19643);
and U24894 (N_24894,N_15599,N_19474);
nand U24895 (N_24895,N_17453,N_15809);
nor U24896 (N_24896,N_16126,N_15437);
nand U24897 (N_24897,N_17205,N_17118);
nand U24898 (N_24898,N_15495,N_19574);
nand U24899 (N_24899,N_15602,N_15164);
or U24900 (N_24900,N_15087,N_16237);
or U24901 (N_24901,N_18412,N_19580);
and U24902 (N_24902,N_16789,N_15491);
nand U24903 (N_24903,N_15754,N_16688);
and U24904 (N_24904,N_16239,N_17885);
or U24905 (N_24905,N_16401,N_16315);
and U24906 (N_24906,N_19618,N_19636);
or U24907 (N_24907,N_19547,N_17097);
nand U24908 (N_24908,N_15793,N_16520);
xnor U24909 (N_24909,N_16212,N_18711);
nand U24910 (N_24910,N_18070,N_17643);
xnor U24911 (N_24911,N_18105,N_17215);
or U24912 (N_24912,N_16381,N_17335);
nor U24913 (N_24913,N_18404,N_19835);
or U24914 (N_24914,N_18347,N_19249);
or U24915 (N_24915,N_16797,N_18115);
and U24916 (N_24916,N_16673,N_18274);
nor U24917 (N_24917,N_17304,N_17579);
nand U24918 (N_24918,N_15285,N_19409);
or U24919 (N_24919,N_18172,N_19354);
and U24920 (N_24920,N_18042,N_16079);
nand U24921 (N_24921,N_19699,N_18304);
and U24922 (N_24922,N_17693,N_17753);
or U24923 (N_24923,N_18848,N_15424);
nor U24924 (N_24924,N_15313,N_16444);
xnor U24925 (N_24925,N_19260,N_19804);
or U24926 (N_24926,N_18288,N_16585);
and U24927 (N_24927,N_19493,N_19305);
nor U24928 (N_24928,N_19912,N_19580);
nor U24929 (N_24929,N_15199,N_18682);
and U24930 (N_24930,N_17986,N_15624);
nand U24931 (N_24931,N_16098,N_15335);
nand U24932 (N_24932,N_18853,N_19012);
or U24933 (N_24933,N_15140,N_16899);
nor U24934 (N_24934,N_17864,N_16099);
or U24935 (N_24935,N_17670,N_18638);
xnor U24936 (N_24936,N_19771,N_17616);
nor U24937 (N_24937,N_15126,N_18404);
or U24938 (N_24938,N_16648,N_16856);
or U24939 (N_24939,N_16958,N_18500);
nor U24940 (N_24940,N_16587,N_19851);
nand U24941 (N_24941,N_17198,N_19767);
nor U24942 (N_24942,N_16351,N_15203);
nand U24943 (N_24943,N_17554,N_16279);
and U24944 (N_24944,N_18542,N_19032);
or U24945 (N_24945,N_18300,N_16929);
or U24946 (N_24946,N_18590,N_18971);
or U24947 (N_24947,N_19526,N_17306);
nand U24948 (N_24948,N_15043,N_15558);
nor U24949 (N_24949,N_18128,N_16234);
nor U24950 (N_24950,N_18219,N_16848);
and U24951 (N_24951,N_17914,N_16191);
nor U24952 (N_24952,N_19795,N_19887);
and U24953 (N_24953,N_15017,N_19444);
nand U24954 (N_24954,N_16521,N_18998);
nand U24955 (N_24955,N_17807,N_18566);
or U24956 (N_24956,N_16812,N_16923);
or U24957 (N_24957,N_17510,N_19874);
or U24958 (N_24958,N_15211,N_18456);
nand U24959 (N_24959,N_18083,N_17781);
and U24960 (N_24960,N_17276,N_19226);
nand U24961 (N_24961,N_15101,N_18916);
or U24962 (N_24962,N_16588,N_19298);
or U24963 (N_24963,N_18842,N_19441);
nor U24964 (N_24964,N_15936,N_18058);
and U24965 (N_24965,N_15264,N_18641);
xnor U24966 (N_24966,N_18211,N_19465);
and U24967 (N_24967,N_17776,N_19491);
or U24968 (N_24968,N_19039,N_15340);
nand U24969 (N_24969,N_17992,N_15266);
nand U24970 (N_24970,N_17377,N_18493);
and U24971 (N_24971,N_18385,N_19482);
or U24972 (N_24972,N_18961,N_16976);
or U24973 (N_24973,N_16507,N_17523);
and U24974 (N_24974,N_18224,N_15616);
nand U24975 (N_24975,N_16036,N_17412);
nor U24976 (N_24976,N_19882,N_16039);
nor U24977 (N_24977,N_19295,N_16974);
and U24978 (N_24978,N_15851,N_15538);
nor U24979 (N_24979,N_18861,N_17403);
xor U24980 (N_24980,N_19629,N_17323);
or U24981 (N_24981,N_15270,N_19895);
and U24982 (N_24982,N_17108,N_18221);
and U24983 (N_24983,N_16803,N_16285);
nand U24984 (N_24984,N_17721,N_17856);
or U24985 (N_24985,N_19300,N_19536);
and U24986 (N_24986,N_18677,N_15321);
or U24987 (N_24987,N_15529,N_15931);
or U24988 (N_24988,N_18124,N_15842);
xor U24989 (N_24989,N_18843,N_18951);
or U24990 (N_24990,N_17528,N_19202);
nand U24991 (N_24991,N_16740,N_17189);
or U24992 (N_24992,N_18339,N_15265);
nor U24993 (N_24993,N_17438,N_18311);
nand U24994 (N_24994,N_18552,N_15106);
nand U24995 (N_24995,N_15254,N_16476);
nand U24996 (N_24996,N_16798,N_17075);
xor U24997 (N_24997,N_15002,N_16065);
nor U24998 (N_24998,N_15938,N_17318);
and U24999 (N_24999,N_16236,N_17664);
nand U25000 (N_25000,N_20025,N_22325);
or U25001 (N_25001,N_21923,N_22852);
nand U25002 (N_25002,N_21032,N_21138);
nand U25003 (N_25003,N_23373,N_20053);
nand U25004 (N_25004,N_20368,N_23747);
nor U25005 (N_25005,N_24052,N_21519);
nand U25006 (N_25006,N_20580,N_21102);
nand U25007 (N_25007,N_23217,N_24192);
nor U25008 (N_25008,N_21575,N_21941);
and U25009 (N_25009,N_22854,N_23782);
and U25010 (N_25010,N_24157,N_22492);
nor U25011 (N_25011,N_21527,N_21635);
or U25012 (N_25012,N_24206,N_23714);
and U25013 (N_25013,N_20963,N_20761);
and U25014 (N_25014,N_24989,N_21021);
xor U25015 (N_25015,N_23769,N_22539);
nand U25016 (N_25016,N_24167,N_20932);
nor U25017 (N_25017,N_22996,N_21967);
or U25018 (N_25018,N_24194,N_22073);
xnor U25019 (N_25019,N_24208,N_22957);
or U25020 (N_25020,N_20888,N_22262);
and U25021 (N_25021,N_21645,N_21351);
or U25022 (N_25022,N_23377,N_22322);
xor U25023 (N_25023,N_20849,N_21149);
nand U25024 (N_25024,N_24193,N_21412);
nand U25025 (N_25025,N_23923,N_23276);
nor U25026 (N_25026,N_24906,N_21757);
nand U25027 (N_25027,N_20263,N_21819);
or U25028 (N_25028,N_24819,N_23531);
nand U25029 (N_25029,N_24999,N_20667);
xnor U25030 (N_25030,N_20553,N_24951);
nor U25031 (N_25031,N_21835,N_21895);
nor U25032 (N_25032,N_22773,N_20991);
and U25033 (N_25033,N_21993,N_24022);
xor U25034 (N_25034,N_24445,N_22398);
and U25035 (N_25035,N_22764,N_23508);
nand U25036 (N_25036,N_24741,N_24674);
nor U25037 (N_25037,N_21000,N_23817);
nand U25038 (N_25038,N_21413,N_20260);
nand U25039 (N_25039,N_23438,N_23055);
nor U25040 (N_25040,N_22568,N_23402);
or U25041 (N_25041,N_24997,N_22536);
nand U25042 (N_25042,N_24371,N_24720);
and U25043 (N_25043,N_22479,N_21740);
nor U25044 (N_25044,N_22236,N_21337);
nand U25045 (N_25045,N_22446,N_24922);
nand U25046 (N_25046,N_22091,N_21140);
nand U25047 (N_25047,N_22562,N_22085);
xnor U25048 (N_25048,N_20472,N_22849);
and U25049 (N_25049,N_24427,N_22139);
nor U25050 (N_25050,N_22529,N_22108);
nor U25051 (N_25051,N_23052,N_23374);
xor U25052 (N_25052,N_20326,N_20352);
nor U25053 (N_25053,N_20798,N_24304);
and U25054 (N_25054,N_22488,N_23810);
nor U25055 (N_25055,N_23935,N_24385);
or U25056 (N_25056,N_24904,N_20639);
nor U25057 (N_25057,N_21613,N_23223);
or U25058 (N_25058,N_23836,N_21057);
nor U25059 (N_25059,N_22182,N_24354);
nand U25060 (N_25060,N_20382,N_23792);
nand U25061 (N_25061,N_22059,N_21456);
nand U25062 (N_25062,N_22602,N_20807);
xor U25063 (N_25063,N_24518,N_21602);
nor U25064 (N_25064,N_22256,N_24935);
nor U25065 (N_25065,N_23786,N_20790);
or U25066 (N_25066,N_24748,N_22368);
nand U25067 (N_25067,N_22503,N_24242);
or U25068 (N_25068,N_20916,N_20389);
or U25069 (N_25069,N_23283,N_23457);
nand U25070 (N_25070,N_23210,N_20370);
or U25071 (N_25071,N_20254,N_22484);
xnor U25072 (N_25072,N_24154,N_23894);
nand U25073 (N_25073,N_22679,N_23441);
nor U25074 (N_25074,N_24909,N_24308);
nor U25075 (N_25075,N_23173,N_23929);
nor U25076 (N_25076,N_22081,N_20669);
or U25077 (N_25077,N_22978,N_21932);
nor U25078 (N_25078,N_22894,N_20616);
nand U25079 (N_25079,N_21467,N_20152);
nor U25080 (N_25080,N_23167,N_24955);
nor U25081 (N_25081,N_21991,N_20784);
or U25082 (N_25082,N_23633,N_22481);
nor U25083 (N_25083,N_23574,N_20999);
nor U25084 (N_25084,N_20655,N_24293);
or U25085 (N_25085,N_22853,N_24482);
nand U25086 (N_25086,N_21499,N_22991);
or U25087 (N_25087,N_23198,N_24841);
nand U25088 (N_25088,N_23968,N_22842);
nand U25089 (N_25089,N_22131,N_20491);
nand U25090 (N_25090,N_24197,N_21958);
nor U25091 (N_25091,N_24013,N_20678);
xnor U25092 (N_25092,N_24356,N_23043);
or U25093 (N_25093,N_22772,N_21704);
and U25094 (N_25094,N_21099,N_24069);
nor U25095 (N_25095,N_23785,N_24611);
nand U25096 (N_25096,N_22440,N_21262);
nor U25097 (N_25097,N_24333,N_24606);
or U25098 (N_25098,N_21183,N_24563);
nand U25099 (N_25099,N_21350,N_22695);
xnor U25100 (N_25100,N_24639,N_24029);
nor U25101 (N_25101,N_21759,N_21386);
or U25102 (N_25102,N_24164,N_22787);
and U25103 (N_25103,N_20413,N_23370);
or U25104 (N_25104,N_22396,N_24613);
and U25105 (N_25105,N_21511,N_21454);
or U25106 (N_25106,N_23113,N_24127);
xor U25107 (N_25107,N_23356,N_20907);
or U25108 (N_25108,N_20820,N_21994);
nand U25109 (N_25109,N_21079,N_23813);
nor U25110 (N_25110,N_20797,N_22389);
and U25111 (N_25111,N_22856,N_23634);
or U25112 (N_25112,N_24269,N_23330);
nand U25113 (N_25113,N_21399,N_23586);
or U25114 (N_25114,N_23411,N_22395);
nand U25115 (N_25115,N_22950,N_22298);
xor U25116 (N_25116,N_22663,N_22283);
or U25117 (N_25117,N_23134,N_23892);
xor U25118 (N_25118,N_23510,N_20613);
nand U25119 (N_25119,N_22016,N_20008);
nor U25120 (N_25120,N_23641,N_22272);
xnor U25121 (N_25121,N_21807,N_20958);
nand U25122 (N_25122,N_20295,N_22905);
and U25123 (N_25123,N_22190,N_24001);
or U25124 (N_25124,N_21788,N_20680);
and U25125 (N_25125,N_24166,N_24497);
nor U25126 (N_25126,N_21111,N_20994);
xor U25127 (N_25127,N_21273,N_24633);
nor U25128 (N_25128,N_23331,N_24693);
xor U25129 (N_25129,N_23538,N_23607);
nor U25130 (N_25130,N_20138,N_20599);
and U25131 (N_25131,N_23532,N_22666);
and U25132 (N_25132,N_24009,N_22023);
nand U25133 (N_25133,N_20819,N_23970);
or U25134 (N_25134,N_21063,N_22351);
nand U25135 (N_25135,N_24586,N_21563);
and U25136 (N_25136,N_23656,N_24831);
and U25137 (N_25137,N_22227,N_22836);
and U25138 (N_25138,N_22668,N_24018);
or U25139 (N_25139,N_24440,N_24776);
or U25140 (N_25140,N_21416,N_24800);
or U25141 (N_25141,N_24188,N_23521);
or U25142 (N_25142,N_24528,N_20332);
nand U25143 (N_25143,N_21472,N_23159);
and U25144 (N_25144,N_21729,N_20894);
nand U25145 (N_25145,N_23300,N_22526);
and U25146 (N_25146,N_21764,N_24111);
nor U25147 (N_25147,N_23419,N_23175);
or U25148 (N_25148,N_22675,N_21049);
or U25149 (N_25149,N_22341,N_21893);
nand U25150 (N_25150,N_24000,N_23738);
or U25151 (N_25151,N_22265,N_21696);
or U25152 (N_25152,N_23784,N_22051);
nand U25153 (N_25153,N_20383,N_23921);
or U25154 (N_25154,N_21338,N_21841);
or U25155 (N_25155,N_21957,N_23190);
nor U25156 (N_25156,N_24797,N_21629);
nor U25157 (N_25157,N_21571,N_24490);
nand U25158 (N_25158,N_21234,N_23561);
nor U25159 (N_25159,N_24682,N_20538);
nand U25160 (N_25160,N_23773,N_20438);
or U25161 (N_25161,N_23671,N_20752);
nor U25162 (N_25162,N_24458,N_23230);
or U25163 (N_25163,N_22816,N_20369);
and U25164 (N_25164,N_23549,N_20544);
nor U25165 (N_25165,N_24576,N_20592);
and U25166 (N_25166,N_21296,N_22469);
or U25167 (N_25167,N_23044,N_24580);
nor U25168 (N_25168,N_21313,N_22589);
or U25169 (N_25169,N_23736,N_21207);
or U25170 (N_25170,N_23611,N_22399);
xnor U25171 (N_25171,N_20753,N_24179);
or U25172 (N_25172,N_22225,N_20965);
and U25173 (N_25173,N_23599,N_24247);
nor U25174 (N_25174,N_22976,N_22753);
and U25175 (N_25175,N_23407,N_24503);
and U25176 (N_25176,N_20247,N_24931);
nand U25177 (N_25177,N_20080,N_22198);
or U25178 (N_25178,N_23439,N_23511);
and U25179 (N_25179,N_22597,N_22625);
and U25180 (N_25180,N_22353,N_24402);
and U25181 (N_25181,N_22092,N_22439);
nand U25182 (N_25182,N_24950,N_23871);
and U25183 (N_25183,N_20978,N_22366);
nor U25184 (N_25184,N_21647,N_21538);
or U25185 (N_25185,N_21656,N_23896);
nand U25186 (N_25186,N_21294,N_21285);
nand U25187 (N_25187,N_20879,N_21053);
or U25188 (N_25188,N_24737,N_24886);
xnor U25189 (N_25189,N_21084,N_22778);
nor U25190 (N_25190,N_20485,N_24722);
nand U25191 (N_25191,N_20444,N_20933);
nand U25192 (N_25192,N_22473,N_24609);
and U25193 (N_25193,N_24519,N_22904);
or U25194 (N_25194,N_20238,N_23033);
or U25195 (N_25195,N_21278,N_22169);
or U25196 (N_25196,N_20399,N_20955);
or U25197 (N_25197,N_23239,N_22645);
and U25198 (N_25198,N_23496,N_21279);
xnor U25199 (N_25199,N_22590,N_24060);
and U25200 (N_25200,N_23909,N_24716);
or U25201 (N_25201,N_21542,N_21559);
xnor U25202 (N_25202,N_20931,N_23358);
nor U25203 (N_25203,N_21266,N_20898);
or U25204 (N_25204,N_24893,N_20125);
xnor U25205 (N_25205,N_24746,N_22191);
or U25206 (N_25206,N_22549,N_22754);
or U25207 (N_25207,N_21614,N_20590);
or U25208 (N_25208,N_21548,N_20361);
or U25209 (N_25209,N_21693,N_24879);
or U25210 (N_25210,N_21995,N_24843);
and U25211 (N_25211,N_24911,N_20030);
nor U25212 (N_25212,N_21621,N_20749);
or U25213 (N_25213,N_24782,N_20467);
nor U25214 (N_25214,N_22638,N_20433);
or U25215 (N_25215,N_22487,N_23357);
or U25216 (N_25216,N_20257,N_22798);
nor U25217 (N_25217,N_22557,N_21875);
and U25218 (N_25218,N_22113,N_23556);
and U25219 (N_25219,N_22974,N_23152);
xor U25220 (N_25220,N_20064,N_22809);
nand U25221 (N_25221,N_21189,N_22648);
nand U25222 (N_25222,N_21016,N_21155);
nand U25223 (N_25223,N_22047,N_24096);
nor U25224 (N_25224,N_22690,N_20111);
or U25225 (N_25225,N_23690,N_24975);
nand U25226 (N_25226,N_20220,N_20595);
and U25227 (N_25227,N_24521,N_23874);
nand U25228 (N_25228,N_22274,N_21179);
or U25229 (N_25229,N_21275,N_21437);
nor U25230 (N_25230,N_21739,N_20930);
and U25231 (N_25231,N_21312,N_20055);
or U25232 (N_25232,N_23169,N_20642);
nand U25233 (N_25233,N_20007,N_22254);
nand U25234 (N_25234,N_24282,N_24983);
nor U25235 (N_25235,N_21796,N_24813);
and U25236 (N_25236,N_22491,N_21134);
nand U25237 (N_25237,N_21362,N_23533);
nand U25238 (N_25238,N_20240,N_23610);
or U25239 (N_25239,N_21789,N_24806);
nor U25240 (N_25240,N_24448,N_21928);
and U25241 (N_25241,N_21238,N_23852);
or U25242 (N_25242,N_23121,N_21342);
and U25243 (N_25243,N_20414,N_21260);
and U25244 (N_25244,N_24311,N_22197);
nor U25245 (N_25245,N_22636,N_24041);
or U25246 (N_25246,N_21485,N_24361);
nor U25247 (N_25247,N_24801,N_20989);
and U25248 (N_25248,N_22723,N_23686);
or U25249 (N_25249,N_22239,N_22917);
or U25250 (N_25250,N_22915,N_22518);
xor U25251 (N_25251,N_23850,N_24271);
nor U25252 (N_25252,N_21818,N_24697);
nor U25253 (N_25253,N_21202,N_22958);
nand U25254 (N_25254,N_20935,N_24837);
nand U25255 (N_25255,N_24021,N_24736);
or U25256 (N_25256,N_24147,N_22001);
nor U25257 (N_25257,N_21390,N_21763);
nor U25258 (N_25258,N_20788,N_21945);
or U25259 (N_25259,N_21082,N_21340);
or U25260 (N_25260,N_20577,N_23528);
nor U25261 (N_25261,N_22610,N_21826);
nor U25262 (N_25262,N_24554,N_24275);
xnor U25263 (N_25263,N_23910,N_24571);
nand U25264 (N_25264,N_22339,N_22014);
nor U25265 (N_25265,N_22717,N_20388);
xnor U25266 (N_25266,N_24349,N_23762);
nor U25267 (N_25267,N_20113,N_24579);
xnor U25268 (N_25268,N_23158,N_23041);
nand U25269 (N_25269,N_24747,N_20156);
or U25270 (N_25270,N_24120,N_20706);
or U25271 (N_25271,N_22998,N_21723);
nor U25272 (N_25272,N_23189,N_21785);
or U25273 (N_25273,N_24701,N_22329);
or U25274 (N_25274,N_20479,N_22735);
nor U25275 (N_25275,N_22519,N_22940);
and U25276 (N_25276,N_24173,N_24391);
nand U25277 (N_25277,N_24520,N_21980);
or U25278 (N_25278,N_20327,N_20391);
or U25279 (N_25279,N_21930,N_24919);
or U25280 (N_25280,N_20116,N_24536);
nor U25281 (N_25281,N_23887,N_22156);
nor U25282 (N_25282,N_21748,N_23424);
nor U25283 (N_25283,N_22660,N_20237);
and U25284 (N_25284,N_20604,N_20543);
and U25285 (N_25285,N_22622,N_21911);
or U25286 (N_25286,N_22486,N_20922);
nand U25287 (N_25287,N_23423,N_20003);
or U25288 (N_25288,N_22459,N_22613);
or U25289 (N_25289,N_21860,N_23063);
or U25290 (N_25290,N_23501,N_23347);
nor U25291 (N_25291,N_22201,N_20620);
xor U25292 (N_25292,N_21095,N_20631);
nor U25293 (N_25293,N_21062,N_22192);
and U25294 (N_25294,N_22616,N_23753);
and U25295 (N_25295,N_22846,N_21944);
and U25296 (N_25296,N_24065,N_23334);
nor U25297 (N_25297,N_21510,N_21500);
or U25298 (N_25298,N_23366,N_22303);
nor U25299 (N_25299,N_21816,N_24646);
or U25300 (N_25300,N_24733,N_22270);
and U25301 (N_25301,N_24724,N_24794);
nor U25302 (N_25302,N_23464,N_22759);
xor U25303 (N_25303,N_20145,N_24936);
nor U25304 (N_25304,N_23428,N_22466);
and U25305 (N_25305,N_23758,N_22183);
and U25306 (N_25306,N_24265,N_24869);
nand U25307 (N_25307,N_21662,N_23202);
xnor U25308 (N_25308,N_24121,N_23990);
nand U25309 (N_25309,N_23706,N_21355);
nand U25310 (N_25310,N_23224,N_20668);
and U25311 (N_25311,N_23141,N_24507);
nor U25312 (N_25312,N_23642,N_20606);
or U25313 (N_25313,N_24867,N_22388);
and U25314 (N_25314,N_23840,N_23997);
and U25315 (N_25315,N_22026,N_22896);
or U25316 (N_25316,N_24086,N_23195);
xor U25317 (N_25317,N_22825,N_24848);
or U25318 (N_25318,N_22495,N_23488);
and U25319 (N_25319,N_20464,N_22107);
and U25320 (N_25320,N_21825,N_21800);
or U25321 (N_25321,N_21889,N_24700);
nand U25322 (N_25322,N_21961,N_20243);
nand U25323 (N_25323,N_22715,N_22464);
or U25324 (N_25324,N_24155,N_23079);
and U25325 (N_25325,N_23073,N_20823);
xnor U25326 (N_25326,N_20057,N_20634);
nor U25327 (N_25327,N_24900,N_20925);
nand U25328 (N_25328,N_24932,N_24822);
nor U25329 (N_25329,N_22767,N_20151);
or U25330 (N_25330,N_21298,N_21498);
or U25331 (N_25331,N_22651,N_22501);
nand U25332 (N_25332,N_21512,N_22137);
nor U25333 (N_25333,N_22004,N_21714);
and U25334 (N_25334,N_22662,N_23920);
or U25335 (N_25335,N_23998,N_21453);
nor U25336 (N_25336,N_23629,N_24364);
nor U25337 (N_25337,N_23550,N_24760);
nor U25338 (N_25338,N_20360,N_21756);
and U25339 (N_25339,N_22944,N_22707);
xnor U25340 (N_25340,N_21025,N_21537);
nor U25341 (N_25341,N_21839,N_23307);
nor U25342 (N_25342,N_22171,N_20862);
nand U25343 (N_25343,N_21599,N_21212);
or U25344 (N_25344,N_21429,N_21979);
and U25345 (N_25345,N_23380,N_22349);
nand U25346 (N_25346,N_24866,N_24882);
or U25347 (N_25347,N_20283,N_23726);
nor U25348 (N_25348,N_22794,N_20939);
xnor U25349 (N_25349,N_24677,N_22166);
or U25350 (N_25350,N_20617,N_23981);
xnor U25351 (N_25351,N_20512,N_21159);
nor U25352 (N_25352,N_21460,N_24028);
nor U25353 (N_25353,N_23906,N_21828);
nor U25354 (N_25354,N_22637,N_22929);
nand U25355 (N_25355,N_23994,N_23135);
or U25356 (N_25356,N_23529,N_20058);
or U25357 (N_25357,N_21555,N_23797);
or U25358 (N_25358,N_20602,N_22714);
and U25359 (N_25359,N_20246,N_23666);
or U25360 (N_25360,N_20762,N_21786);
nor U25361 (N_25361,N_21859,N_22581);
nand U25362 (N_25362,N_22618,N_23947);
and U25363 (N_25363,N_23685,N_23091);
or U25364 (N_25364,N_20800,N_22154);
xnor U25365 (N_25365,N_22806,N_22851);
or U25366 (N_25366,N_22470,N_20105);
nor U25367 (N_25367,N_23491,N_24469);
and U25368 (N_25368,N_21925,N_20094);
nand U25369 (N_25369,N_22064,N_24793);
or U25370 (N_25370,N_20262,N_21607);
and U25371 (N_25371,N_22890,N_20518);
or U25372 (N_25372,N_20206,N_21047);
and U25373 (N_25373,N_22583,N_22078);
xor U25374 (N_25374,N_22134,N_21968);
nand U25375 (N_25375,N_24549,N_22942);
xnor U25376 (N_25376,N_21104,N_24014);
and U25377 (N_25377,N_21824,N_20778);
nor U25378 (N_25378,N_21906,N_21644);
nand U25379 (N_25379,N_23891,N_21592);
nor U25380 (N_25380,N_20398,N_21473);
nor U25381 (N_25381,N_24446,N_24126);
or U25382 (N_25382,N_20685,N_23716);
nand U25383 (N_25383,N_23737,N_24807);
nor U25384 (N_25384,N_23127,N_22316);
nand U25385 (N_25385,N_22784,N_20333);
or U25386 (N_25386,N_21648,N_21557);
and U25387 (N_25387,N_22728,N_21710);
nand U25388 (N_25388,N_22511,N_23150);
and U25389 (N_25389,N_21843,N_22505);
nor U25390 (N_25390,N_22009,N_20196);
and U25391 (N_25391,N_22121,N_24138);
nand U25392 (N_25392,N_23243,N_23804);
xnor U25393 (N_25393,N_23142,N_22685);
nand U25394 (N_25394,N_20217,N_24943);
or U25395 (N_25395,N_22884,N_20272);
and U25396 (N_25396,N_24073,N_21680);
and U25397 (N_25397,N_20830,N_24338);
nor U25398 (N_25398,N_21131,N_20816);
nor U25399 (N_25399,N_24033,N_20841);
nor U25400 (N_25400,N_23086,N_23339);
nand U25401 (N_25401,N_23614,N_24510);
xor U25402 (N_25402,N_20846,N_22133);
nand U25403 (N_25403,N_24080,N_22011);
nand U25404 (N_25404,N_21291,N_21531);
nor U25405 (N_25405,N_23883,N_24144);
nor U25406 (N_25406,N_24555,N_21496);
or U25407 (N_25407,N_23609,N_22444);
nor U25408 (N_25408,N_21108,N_21410);
or U25409 (N_25409,N_21425,N_20420);
and U25410 (N_25410,N_24079,N_22665);
nand U25411 (N_25411,N_24487,N_21147);
xnor U25412 (N_25412,N_22909,N_20603);
or U25413 (N_25413,N_21314,N_23960);
or U25414 (N_25414,N_20489,N_20640);
and U25415 (N_25415,N_23912,N_22782);
and U25416 (N_25416,N_21735,N_22994);
or U25417 (N_25417,N_20627,N_22098);
and U25418 (N_25418,N_21344,N_23245);
and U25419 (N_25419,N_21589,N_20615);
nor U25420 (N_25420,N_23881,N_24093);
or U25421 (N_25421,N_24332,N_23467);
nand U25422 (N_25422,N_20068,N_21431);
nand U25423 (N_25423,N_23697,N_22623);
nand U25424 (N_25424,N_21105,N_24237);
or U25425 (N_25425,N_20498,N_21752);
nor U25426 (N_25426,N_23333,N_20929);
or U25427 (N_25427,N_23986,N_20101);
nand U25428 (N_25428,N_20244,N_20322);
nand U25429 (N_25429,N_21657,N_23319);
or U25430 (N_25430,N_24235,N_20918);
nand U25431 (N_25431,N_24454,N_22771);
nor U25432 (N_25432,N_22386,N_22312);
or U25433 (N_25433,N_21609,N_24233);
nand U25434 (N_25434,N_24310,N_24163);
and U25435 (N_25435,N_24840,N_24309);
nor U25436 (N_25436,N_20902,N_20833);
nor U25437 (N_25437,N_22509,N_21119);
nor U25438 (N_25438,N_23070,N_22431);
nor U25439 (N_25439,N_20037,N_21409);
nand U25440 (N_25440,N_21722,N_21332);
nor U25441 (N_25441,N_23013,N_24849);
nor U25442 (N_25442,N_22937,N_23101);
nand U25443 (N_25443,N_20059,N_22416);
or U25444 (N_25444,N_24673,N_22530);
and U25445 (N_25445,N_22973,N_23776);
or U25446 (N_25446,N_20131,N_23473);
or U25447 (N_25447,N_21896,N_22641);
nor U25448 (N_25448,N_20724,N_20173);
nor U25449 (N_25449,N_24320,N_20868);
nor U25450 (N_25450,N_22591,N_21664);
or U25451 (N_25451,N_20740,N_22152);
nor U25452 (N_25452,N_24400,N_20195);
and U25453 (N_25453,N_22814,N_20813);
or U25454 (N_25454,N_20066,N_21365);
and U25455 (N_25455,N_20396,N_24108);
or U25456 (N_25456,N_24815,N_23145);
nand U25457 (N_25457,N_20284,N_21805);
or U25458 (N_25458,N_21681,N_20044);
or U25459 (N_25459,N_22263,N_22879);
or U25460 (N_25460,N_23188,N_24923);
or U25461 (N_25461,N_20767,N_24035);
nor U25462 (N_25462,N_20968,N_24566);
nor U25463 (N_25463,N_21576,N_21290);
and U25464 (N_25464,N_21914,N_22523);
xor U25465 (N_25465,N_20488,N_21433);
nor U25466 (N_25466,N_23645,N_23932);
xnor U25467 (N_25467,N_24421,N_20161);
nor U25468 (N_25468,N_22652,N_22063);
or U25469 (N_25469,N_23100,N_22378);
and U25470 (N_25470,N_22172,N_21489);
and U25471 (N_25471,N_23416,N_23936);
or U25472 (N_25472,N_21089,N_20702);
and U25473 (N_25473,N_21056,N_22676);
and U25474 (N_25474,N_22199,N_22456);
and U25475 (N_25475,N_22595,N_23133);
nand U25476 (N_25476,N_23206,N_23745);
nand U25477 (N_25477,N_23824,N_23009);
nand U25478 (N_25478,N_20884,N_24191);
or U25479 (N_25479,N_23130,N_24859);
or U25480 (N_25480,N_24072,N_23272);
nor U25481 (N_25481,N_22148,N_22955);
nor U25482 (N_25482,N_23543,N_22374);
nor U25483 (N_25483,N_23901,N_24861);
nor U25484 (N_25484,N_20435,N_24562);
nand U25485 (N_25485,N_20476,N_20385);
nand U25486 (N_25486,N_24687,N_22164);
nor U25487 (N_25487,N_23658,N_22045);
nor U25488 (N_25488,N_20160,N_24873);
or U25489 (N_25489,N_23360,N_22403);
xor U25490 (N_25490,N_20927,N_20738);
and U25491 (N_25491,N_24903,N_23708);
nor U25492 (N_25492,N_22354,N_21129);
nand U25493 (N_25493,N_24714,N_23525);
xnor U25494 (N_25494,N_20141,N_20802);
nor U25495 (N_25495,N_22919,N_23085);
nand U25496 (N_25496,N_20890,N_22848);
nor U25497 (N_25497,N_21534,N_23075);
nor U25498 (N_25498,N_21211,N_21252);
xor U25499 (N_25499,N_21164,N_20387);
nor U25500 (N_25500,N_21865,N_20757);
and U25501 (N_25501,N_22100,N_21639);
or U25502 (N_25502,N_22251,N_20024);
and U25503 (N_25503,N_23131,N_24303);
nand U25504 (N_25504,N_24378,N_24297);
nand U25505 (N_25505,N_21588,N_24444);
or U25506 (N_25506,N_24336,N_22158);
and U25507 (N_25507,N_23707,N_21243);
or U25508 (N_25508,N_24447,N_21215);
and U25509 (N_25509,N_20231,N_24223);
nor U25510 (N_25510,N_24964,N_22364);
nand U25511 (N_25511,N_23895,N_24413);
or U25512 (N_25512,N_22290,N_24025);
nor U25513 (N_25513,N_22101,N_24838);
nor U25514 (N_25514,N_24212,N_24513);
or U25515 (N_25515,N_20940,N_22828);
and U25516 (N_25516,N_23249,N_21643);
nand U25517 (N_25517,N_23165,N_22604);
or U25518 (N_25518,N_22576,N_24852);
and U25519 (N_25519,N_21231,N_23717);
xnor U25520 (N_25520,N_24387,N_23186);
nand U25521 (N_25521,N_23568,N_24277);
xor U25522 (N_25522,N_21281,N_23280);
nand U25523 (N_25523,N_21514,N_23325);
and U25524 (N_25524,N_20551,N_21902);
nand U25525 (N_25525,N_23934,N_24501);
and U25526 (N_25526,N_23290,N_20375);
nor U25527 (N_25527,N_23696,N_23916);
nand U25528 (N_25528,N_21985,N_24643);
or U25529 (N_25529,N_22337,N_22282);
nor U25530 (N_25530,N_23308,N_20204);
nor U25531 (N_25531,N_23800,N_24056);
and U25532 (N_25532,N_24169,N_23514);
nand U25533 (N_25533,N_21854,N_21136);
or U25534 (N_25534,N_21176,N_22605);
or U25535 (N_25535,N_22483,N_22921);
nor U25536 (N_25536,N_21076,N_21130);
nand U25537 (N_25537,N_21781,N_23177);
or U25538 (N_25538,N_22619,N_23911);
or U25539 (N_25539,N_21815,N_20944);
nor U25540 (N_25540,N_20677,N_21910);
and U25541 (N_25541,N_21276,N_21758);
nand U25542 (N_25542,N_22963,N_21146);
xor U25543 (N_25543,N_23818,N_23823);
nor U25544 (N_25544,N_22678,N_23576);
and U25545 (N_25545,N_21526,N_20719);
xnor U25546 (N_25546,N_21028,N_24266);
nor U25547 (N_25547,N_20273,N_24071);
or U25548 (N_25548,N_23674,N_23343);
nand U25549 (N_25549,N_21829,N_20202);
or U25550 (N_25550,N_23375,N_23160);
nor U25551 (N_25551,N_22918,N_23821);
nor U25552 (N_25552,N_21521,N_20662);
xnor U25553 (N_25553,N_23459,N_21087);
nor U25554 (N_25554,N_21624,N_23434);
nand U25555 (N_25555,N_22196,N_23781);
or U25556 (N_25556,N_22343,N_20222);
nand U25557 (N_25557,N_20765,N_20814);
nor U25558 (N_25558,N_22360,N_21570);
or U25559 (N_25559,N_22713,N_24128);
nand U25560 (N_25560,N_23578,N_21002);
or U25561 (N_25561,N_21356,N_24545);
and U25562 (N_25562,N_23326,N_22693);
nand U25563 (N_25563,N_22281,N_23724);
nor U25564 (N_25564,N_23337,N_24486);
nor U25565 (N_25565,N_24526,N_21442);
nand U25566 (N_25566,N_23191,N_24755);
or U25567 (N_25567,N_24229,N_23861);
nor U25568 (N_25568,N_20528,N_23420);
or U25569 (N_25569,N_21560,N_21697);
or U25570 (N_25570,N_21840,N_20928);
nor U25571 (N_25571,N_23081,N_21667);
xor U25572 (N_25572,N_22476,N_24019);
or U25573 (N_25573,N_20271,N_20536);
nor U25574 (N_25574,N_24102,N_23455);
nand U25575 (N_25575,N_24381,N_21078);
and U25576 (N_25576,N_20162,N_23025);
nor U25577 (N_25577,N_20972,N_24871);
and U25578 (N_25578,N_23028,N_23317);
or U25579 (N_25579,N_22401,N_20612);
and U25580 (N_25580,N_22186,N_22383);
and U25581 (N_25581,N_24088,N_23648);
nor U25582 (N_25582,N_20205,N_23787);
and U25583 (N_25583,N_24498,N_20436);
nand U25584 (N_25584,N_23677,N_20451);
xor U25585 (N_25585,N_22614,N_20892);
xnor U25586 (N_25586,N_22769,N_21832);
or U25587 (N_25587,N_22818,N_22095);
nor U25588 (N_25588,N_22032,N_22141);
nor U25589 (N_25589,N_24731,N_24628);
nor U25590 (N_25590,N_22050,N_22385);
or U25591 (N_25591,N_24564,N_23124);
nand U25592 (N_25592,N_21121,N_20946);
or U25593 (N_25593,N_23474,N_23262);
nand U25594 (N_25594,N_21253,N_20411);
nand U25595 (N_25595,N_22468,N_21209);
and U25596 (N_25596,N_21270,N_23060);
nor U25597 (N_25597,N_21267,N_24842);
nand U25598 (N_25598,N_20676,N_22792);
nor U25599 (N_25599,N_21451,N_22061);
or U25600 (N_25600,N_22430,N_23996);
and U25601 (N_25601,N_20673,N_22302);
nand U25602 (N_25602,N_22797,N_22136);
nor U25603 (N_25603,N_23155,N_21309);
nor U25604 (N_25604,N_22324,N_22427);
nand U25605 (N_25605,N_23396,N_23903);
and U25606 (N_25606,N_20869,N_23289);
and U25607 (N_25607,N_23269,N_22903);
nor U25608 (N_25608,N_22730,N_23842);
nand U25609 (N_25609,N_21573,N_24239);
nand U25610 (N_25610,N_23793,N_20310);
and U25611 (N_25611,N_24256,N_24844);
nor U25612 (N_25612,N_24270,N_22391);
nor U25613 (N_25613,N_23640,N_23316);
or U25614 (N_25614,N_24551,N_23522);
nor U25615 (N_25615,N_21048,N_23809);
nand U25616 (N_25616,N_22512,N_20526);
and U25617 (N_25617,N_24612,N_22621);
nor U25618 (N_25618,N_21019,N_21586);
nor U25619 (N_25619,N_24185,N_21006);
or U25620 (N_25620,N_20109,N_21751);
and U25621 (N_25621,N_20475,N_23875);
nand U25622 (N_25622,N_21227,N_22987);
or U25623 (N_25623,N_23575,N_24135);
nor U25624 (N_25624,N_24790,N_20517);
xor U25625 (N_25625,N_21037,N_21734);
xor U25626 (N_25626,N_24341,N_20176);
nor U25627 (N_25627,N_23702,N_21700);
nand U25628 (N_25628,N_24434,N_21794);
nor U25629 (N_25629,N_22860,N_22422);
and U25630 (N_25630,N_23241,N_20809);
and U25631 (N_25631,N_24343,N_21778);
nor U25632 (N_25632,N_23097,N_20947);
and U25633 (N_25633,N_24665,N_24532);
nor U25634 (N_25634,N_20624,N_23036);
nand U25635 (N_25635,N_21686,N_20727);
nand U25636 (N_25636,N_20893,N_20504);
and U25637 (N_25637,N_22507,N_23417);
nand U25638 (N_25638,N_22489,N_21584);
nand U25639 (N_25639,N_20660,N_24927);
or U25640 (N_25640,N_20985,N_23246);
or U25641 (N_25641,N_23178,N_20400);
xor U25642 (N_25642,N_24032,N_22804);
and U25643 (N_25643,N_22543,N_20643);
and U25644 (N_25644,N_20713,N_23140);
nor U25645 (N_25645,N_24634,N_20026);
or U25646 (N_25646,N_20874,N_24313);
and U25647 (N_25647,N_23489,N_20714);
or U25648 (N_25648,N_21730,N_24038);
nand U25649 (N_25649,N_20618,N_23218);
nor U25650 (N_25650,N_21046,N_21919);
nand U25651 (N_25651,N_23777,N_23363);
nor U25652 (N_25652,N_20229,N_20394);
and U25653 (N_25653,N_20966,N_22318);
nand U25654 (N_25654,N_21846,N_21026);
and U25655 (N_25655,N_21424,N_22938);
and U25656 (N_25656,N_21989,N_23476);
nor U25657 (N_25657,N_24635,N_21192);
or U25658 (N_25658,N_20088,N_22229);
nor U25659 (N_25659,N_22872,N_20521);
nor U25660 (N_25660,N_20633,N_20339);
and U25661 (N_25661,N_24511,N_20574);
and U25662 (N_25662,N_22048,N_20781);
nor U25663 (N_25663,N_23566,N_23978);
and U25664 (N_25664,N_22986,N_20278);
nor U25665 (N_25665,N_22887,N_20537);
nor U25666 (N_25666,N_23477,N_24345);
and U25667 (N_25667,N_21445,N_22686);
nand U25668 (N_25668,N_21827,N_20571);
or U25669 (N_25669,N_21115,N_21983);
nand U25670 (N_25670,N_24896,N_20286);
and U25671 (N_25671,N_20956,N_20952);
and U25672 (N_25672,N_20657,N_23019);
and U25673 (N_25673,N_23770,N_21219);
or U25674 (N_25674,N_21972,N_24679);
nor U25675 (N_25675,N_21083,N_22130);
or U25676 (N_25676,N_22140,N_21640);
nor U25677 (N_25677,N_24203,N_24970);
and U25678 (N_25678,N_22346,N_20137);
or U25679 (N_25679,N_24727,N_22542);
nor U25680 (N_25680,N_21633,N_22964);
nor U25681 (N_25681,N_21707,N_21845);
and U25682 (N_25682,N_22862,N_20224);
or U25683 (N_25683,N_21539,N_21926);
nor U25684 (N_25684,N_22708,N_20213);
or U25685 (N_25685,N_24671,N_20440);
nor U25686 (N_25686,N_23985,N_22706);
nand U25687 (N_25687,N_23435,N_20167);
nand U25688 (N_25688,N_23830,N_21984);
and U25689 (N_25689,N_24407,N_24538);
and U25690 (N_25690,N_21254,N_22408);
nor U25691 (N_25691,N_21011,N_21590);
and U25692 (N_25692,N_22761,N_22603);
and U25693 (N_25693,N_24678,N_23594);
and U25694 (N_25694,N_20381,N_20630);
nand U25695 (N_25695,N_24876,N_21372);
nor U25696 (N_25696,N_23016,N_24565);
xor U25697 (N_25697,N_23010,N_22429);
or U25698 (N_25698,N_24567,N_22554);
nor U25699 (N_25699,N_22727,N_20144);
nand U25700 (N_25700,N_21605,N_20710);
or U25701 (N_25701,N_24370,N_21116);
nor U25702 (N_25702,N_23197,N_21746);
and U25703 (N_25703,N_21598,N_22382);
nor U25704 (N_25704,N_21731,N_22242);
nor U25705 (N_25705,N_20725,N_21072);
or U25706 (N_25706,N_22544,N_24437);
nor U25707 (N_25707,N_23524,N_21886);
xnor U25708 (N_25708,N_24392,N_23761);
and U25709 (N_25709,N_24373,N_22423);
or U25710 (N_25710,N_20021,N_22683);
nor U25711 (N_25711,N_23612,N_24124);
nand U25712 (N_25712,N_24912,N_22830);
or U25713 (N_25713,N_24734,N_21947);
or U25714 (N_25714,N_20157,N_20031);
and U25715 (N_25715,N_21646,N_24845);
or U25716 (N_25716,N_20812,N_21250);
and U25717 (N_25717,N_20306,N_21933);
or U25718 (N_25718,N_22493,N_23042);
nor U25719 (N_25719,N_22810,N_21091);
nor U25720 (N_25720,N_22864,N_22114);
nor U25721 (N_25721,N_20611,N_22005);
and U25722 (N_25722,N_23597,N_22897);
and U25723 (N_25723,N_23967,N_24337);
nor U25724 (N_25724,N_20503,N_24732);
nand U25725 (N_25725,N_20015,N_24418);
and U25726 (N_25726,N_20920,N_21034);
nand U25727 (N_25727,N_23164,N_20839);
nand U25728 (N_25728,N_22218,N_22052);
or U25729 (N_25729,N_23312,N_23463);
nor U25730 (N_25730,N_23233,N_23064);
nor U25731 (N_25731,N_22700,N_21152);
and U25732 (N_25732,N_24207,N_21411);
and U25733 (N_25733,N_22060,N_22044);
and U25734 (N_25734,N_22128,N_23478);
nor U25735 (N_25735,N_21029,N_20771);
nand U25736 (N_25736,N_24803,N_20199);
nor U25737 (N_25737,N_20165,N_24512);
or U25738 (N_25738,N_20579,N_24854);
or U25739 (N_25739,N_24756,N_23277);
or U25740 (N_25740,N_23076,N_21616);
or U25741 (N_25741,N_21682,N_20908);
or U25742 (N_25742,N_20881,N_24307);
nand U25743 (N_25743,N_21727,N_24982);
nor U25744 (N_25744,N_23207,N_23583);
and U25745 (N_25745,N_22125,N_22226);
and U25746 (N_25746,N_22522,N_21122);
nor U25747 (N_25747,N_20748,N_20795);
nor U25748 (N_25748,N_21619,N_23059);
and U25749 (N_25749,N_20232,N_23311);
nor U25750 (N_25750,N_22895,N_20614);
xor U25751 (N_25751,N_20746,N_24597);
nor U25752 (N_25752,N_21393,N_24048);
and U25753 (N_25753,N_24067,N_22228);
nor U25754 (N_25754,N_20358,N_20638);
or U25755 (N_25755,N_20014,N_21903);
nor U25756 (N_25756,N_24502,N_20683);
or U25757 (N_25757,N_21345,N_23625);
or U25758 (N_25758,N_22596,N_21650);
nor U25759 (N_25759,N_20148,N_20523);
or U25760 (N_25760,N_20741,N_21150);
nor U25761 (N_25761,N_20001,N_22321);
nand U25762 (N_25762,N_21986,N_21566);
xor U25763 (N_25763,N_20519,N_24034);
nand U25764 (N_25764,N_20699,N_23021);
nand U25765 (N_25765,N_22205,N_22300);
and U25766 (N_25766,N_20117,N_21475);
and U25767 (N_25767,N_23123,N_22980);
nor U25768 (N_25768,N_21615,N_24616);
or U25769 (N_25769,N_23957,N_21597);
or U25770 (N_25770,N_20835,N_24419);
or U25771 (N_25771,N_22537,N_21814);
or U25772 (N_25772,N_21915,N_20269);
or U25773 (N_25773,N_20529,N_22999);
nor U25774 (N_25774,N_24832,N_21673);
nor U25775 (N_25775,N_23045,N_21811);
and U25776 (N_25776,N_24280,N_24531);
and U25777 (N_25777,N_21359,N_21092);
or U25778 (N_25778,N_22572,N_22087);
nor U25779 (N_25779,N_21162,N_23296);
nor U25780 (N_25780,N_21959,N_24666);
nor U25781 (N_25781,N_21223,N_23351);
xnor U25782 (N_25782,N_23530,N_23421);
nor U25783 (N_25783,N_20428,N_20878);
nand U25784 (N_25784,N_24003,N_22674);
and U25785 (N_25785,N_24578,N_21750);
and U25786 (N_25786,N_20909,N_22257);
or U25787 (N_25787,N_21286,N_22635);
or U25788 (N_25788,N_23361,N_22264);
nor U25789 (N_25789,N_24953,N_22891);
nand U25790 (N_25790,N_20975,N_23115);
nand U25791 (N_25791,N_22545,N_21258);
or U25792 (N_25792,N_20720,N_20743);
nand U25793 (N_25793,N_20324,N_20190);
nand U25794 (N_25794,N_24657,N_24824);
or U25795 (N_25795,N_24995,N_21151);
nor U25796 (N_25796,N_24134,N_20248);
xnor U25797 (N_25797,N_21564,N_21330);
and U25798 (N_25798,N_24181,N_23676);
and U25799 (N_25799,N_20122,N_21610);
or U25800 (N_25800,N_20338,N_22402);
nor U25801 (N_25801,N_21572,N_24986);
nand U25802 (N_25802,N_21248,N_24775);
xnor U25803 (N_25803,N_22912,N_21660);
nor U25804 (N_25804,N_24170,N_20242);
nand U25805 (N_25805,N_20335,N_22328);
nand U25806 (N_25806,N_24058,N_22173);
nor U25807 (N_25807,N_23801,N_22765);
nor U25808 (N_25808,N_20664,N_24706);
or U25809 (N_25809,N_24187,N_21898);
and U25810 (N_25810,N_22617,N_24552);
nand U25811 (N_25811,N_22881,N_24651);
and U25812 (N_25812,N_24753,N_23214);
nor U25813 (N_25813,N_22993,N_21166);
xor U25814 (N_25814,N_20062,N_20653);
and U25815 (N_25815,N_24295,N_22371);
nand U25816 (N_25816,N_24479,N_23185);
xnor U25817 (N_25817,N_22012,N_24417);
or U25818 (N_25818,N_24759,N_20754);
and U25819 (N_25819,N_23376,N_23030);
and U25820 (N_25820,N_24853,N_24718);
nor U25821 (N_25821,N_24189,N_23866);
and U25822 (N_25822,N_21465,N_22241);
or U25823 (N_25823,N_21349,N_24694);
nor U25824 (N_25824,N_21637,N_21524);
or U25825 (N_25825,N_21569,N_21545);
or U25826 (N_25826,N_21198,N_24360);
nand U25827 (N_25827,N_20033,N_22117);
and U25828 (N_25828,N_20046,N_23342);
nand U25829 (N_25829,N_23650,N_20777);
or U25830 (N_25830,N_20096,N_23267);
nor U25831 (N_25831,N_22453,N_24202);
nor U25832 (N_25832,N_23759,N_22736);
or U25833 (N_25833,N_22553,N_22965);
and U25834 (N_25834,N_24262,N_24377);
or U25835 (N_25835,N_20216,N_22342);
nor U25836 (N_25836,N_22550,N_23288);
and U25837 (N_25837,N_24944,N_23050);
nor U25838 (N_25838,N_22409,N_22646);
xnor U25839 (N_25839,N_23595,N_21861);
nand U25840 (N_25840,N_22160,N_21305);
and U25841 (N_25841,N_20290,N_20483);
xnor U25842 (N_25842,N_20961,N_21361);
nor U25843 (N_25843,N_21113,N_20723);
or U25844 (N_25844,N_20482,N_22096);
nand U25845 (N_25845,N_24104,N_23973);
or U25846 (N_25846,N_23746,N_24946);
nor U25847 (N_25847,N_24357,N_22962);
nand U25848 (N_25848,N_22945,N_21156);
and U25849 (N_25849,N_24383,N_24113);
or U25850 (N_25850,N_22943,N_20129);
nor U25851 (N_25851,N_20166,N_24816);
and U25852 (N_25852,N_23553,N_21767);
nor U25853 (N_25853,N_21998,N_21617);
and U25854 (N_25854,N_20127,N_21315);
xnor U25855 (N_25855,N_22320,N_21188);
and U25856 (N_25856,N_23495,N_23453);
nand U25857 (N_25857,N_23944,N_21543);
nand U25858 (N_25858,N_20139,N_24592);
or U25859 (N_25859,N_20870,N_22204);
or U25860 (N_25860,N_21677,N_21831);
xor U25861 (N_25861,N_23889,N_21110);
or U25862 (N_25862,N_24328,N_23893);
nand U25863 (N_25863,N_21237,N_20093);
nand U25864 (N_25864,N_24055,N_21161);
or U25865 (N_25865,N_24175,N_23252);
and U25866 (N_25866,N_21018,N_21582);
nor U25867 (N_25867,N_23591,N_22586);
xnor U25868 (N_25868,N_22189,N_21204);
and U25869 (N_25869,N_22404,N_23832);
xnor U25870 (N_25870,N_20457,N_22234);
or U25871 (N_25871,N_24990,N_21435);
nand U25872 (N_25872,N_23132,N_21240);
or U25873 (N_25873,N_21065,N_22116);
nand U25874 (N_25874,N_20136,N_20739);
nand U25875 (N_25875,N_20251,N_24312);
or U25876 (N_25876,N_20281,N_22672);
or U25877 (N_25877,N_22989,N_23067);
or U25878 (N_25878,N_24097,N_22559);
or U25879 (N_25879,N_20585,N_23722);
nand U25880 (N_25880,N_24940,N_20711);
nor U25881 (N_25881,N_21868,N_20570);
or U25882 (N_25882,N_22961,N_22067);
and U25883 (N_25883,N_21094,N_20960);
and U25884 (N_25884,N_20034,N_21611);
nand U25885 (N_25885,N_20346,N_21101);
nand U25886 (N_25886,N_22471,N_22763);
and U25887 (N_25887,N_20460,N_21905);
nor U25888 (N_25888,N_20227,N_21222);
and U25889 (N_25889,N_20962,N_21387);
nand U25890 (N_25890,N_23108,N_20513);
xor U25891 (N_25891,N_24279,N_21301);
and U25892 (N_25892,N_21909,N_20252);
nand U25893 (N_25893,N_22266,N_21098);
xnor U25894 (N_25894,N_22821,N_22452);
or U25895 (N_25895,N_23783,N_23670);
nor U25896 (N_25896,N_22969,N_21158);
nor U25897 (N_25897,N_23427,N_23877);
and U25898 (N_25898,N_20071,N_22411);
nand U25899 (N_25899,N_22901,N_24621);
or U25900 (N_25900,N_21368,N_21711);
and U25901 (N_25901,N_20721,N_21741);
and U25902 (N_25902,N_23034,N_21769);
or U25903 (N_25903,N_23456,N_21225);
nor U25904 (N_25904,N_21988,N_22547);
nor U25905 (N_25905,N_24376,N_20871);
or U25906 (N_25906,N_21354,N_23739);
xnor U25907 (N_25907,N_21749,N_22340);
nand U25908 (N_25908,N_22033,N_24728);
or U25909 (N_25909,N_23372,N_20681);
or U25910 (N_25910,N_24393,N_22040);
nor U25911 (N_25911,N_24217,N_23682);
and U25912 (N_25912,N_20686,N_20006);
nand U25913 (N_25913,N_21671,N_21373);
or U25914 (N_25914,N_23117,N_21812);
nand U25915 (N_25915,N_23475,N_22527);
and U25916 (N_25916,N_23038,N_20431);
and U25917 (N_25917,N_22010,N_22405);
nor U25918 (N_25918,N_23654,N_22058);
and U25919 (N_25919,N_21706,N_22090);
nor U25920 (N_25920,N_21884,N_24617);
and U25921 (N_25921,N_24384,N_24934);
and U25922 (N_25922,N_23798,N_22217);
or U25923 (N_25923,N_24779,N_22151);
nand U25924 (N_25924,N_21720,N_21488);
xnor U25925 (N_25925,N_24214,N_21771);
nor U25926 (N_25926,N_21728,N_21701);
nand U25927 (N_25927,N_20466,N_24130);
or U25928 (N_25928,N_23993,N_20534);
and U25929 (N_25929,N_21307,N_22827);
and U25930 (N_25930,N_20575,N_22650);
nand U25931 (N_25931,N_24092,N_22516);
or U25932 (N_25932,N_22296,N_21665);
nor U25933 (N_25933,N_21999,N_24799);
and U25934 (N_25934,N_21604,N_20957);
nand U25935 (N_25935,N_21666,N_21385);
nor U25936 (N_25936,N_24451,N_22657);
nand U25937 (N_25937,N_23661,N_20022);
and U25938 (N_25938,N_21074,N_21073);
nor U25939 (N_25939,N_23933,N_20390);
or U25940 (N_25940,N_24228,N_21481);
or U25941 (N_25941,N_21546,N_21163);
nor U25942 (N_25942,N_21316,N_24152);
nor U25943 (N_25943,N_22647,N_20511);
nor U25944 (N_25944,N_21689,N_21263);
nand U25945 (N_25945,N_24401,N_24818);
and U25946 (N_25946,N_20774,N_24227);
or U25947 (N_25947,N_22482,N_21943);
nor U25948 (N_25948,N_23292,N_20313);
and U25949 (N_25949,N_20500,N_20533);
or U25950 (N_25950,N_24367,N_20042);
nand U25951 (N_25951,N_20155,N_20850);
nor U25952 (N_25952,N_24763,N_23196);
xor U25953 (N_25953,N_22038,N_24389);
nor U25954 (N_25954,N_23637,N_24785);
nor U25955 (N_25955,N_23392,N_24524);
nor U25956 (N_25956,N_21495,N_21549);
and U25957 (N_25957,N_22042,N_24645);
and U25958 (N_25958,N_23888,N_21492);
and U25959 (N_25959,N_24620,N_22770);
nand U25960 (N_25960,N_20462,N_22267);
and U25961 (N_25961,N_20214,N_21230);
xor U25962 (N_25962,N_21333,N_23318);
or U25963 (N_25963,N_21096,N_24978);
nor U25964 (N_25964,N_23849,N_20410);
or U25965 (N_25965,N_21304,N_24456);
and U25966 (N_25966,N_21770,N_24176);
xnor U25967 (N_25967,N_20374,N_20547);
nor U25968 (N_25968,N_21551,N_24914);
nor U25969 (N_25969,N_20731,N_23963);
or U25970 (N_25970,N_22742,N_20110);
nor U25971 (N_25971,N_20610,N_24083);
xor U25972 (N_25972,N_24348,N_23945);
and U25973 (N_25973,N_23096,N_20114);
or U25974 (N_25974,N_24575,N_20019);
xnor U25975 (N_25975,N_20808,N_22802);
or U25976 (N_25976,N_21497,N_23608);
nor U25977 (N_25977,N_21556,N_23914);
and U25978 (N_25978,N_22375,N_20477);
or U25979 (N_25979,N_20048,N_22206);
and U25980 (N_25980,N_20622,N_20722);
or U25981 (N_25981,N_23772,N_24825);
or U25982 (N_25982,N_22608,N_23516);
or U25983 (N_25983,N_22178,N_20292);
or U25984 (N_25984,N_21142,N_23503);
nand U25985 (N_25985,N_21503,N_23494);
nor U25986 (N_25986,N_23848,N_23338);
and U25987 (N_25987,N_23105,N_23766);
xor U25988 (N_25988,N_22995,N_22142);
and U25989 (N_25989,N_23281,N_24987);
and U25990 (N_25990,N_24325,N_21462);
nand U25991 (N_25991,N_24290,N_23483);
nor U25992 (N_25992,N_21493,N_24961);
or U25993 (N_25993,N_24875,N_21203);
nand U25994 (N_25994,N_20527,N_23964);
nor U25995 (N_25995,N_24902,N_22631);
and U25996 (N_25996,N_24846,N_20915);
and U25997 (N_25997,N_22057,N_23791);
nand U25998 (N_25998,N_21953,N_20650);
nand U25999 (N_25999,N_24076,N_22642);
or U26000 (N_26000,N_20424,N_23322);
nor U26001 (N_26001,N_22531,N_22384);
and U26002 (N_26002,N_23635,N_24828);
and U26003 (N_26003,N_23949,N_21516);
or U26004 (N_26004,N_24662,N_21817);
nand U26005 (N_26005,N_23639,N_23418);
and U26006 (N_26006,N_21154,N_21685);
nor U26007 (N_26007,N_23106,N_20654);
or U26008 (N_26008,N_22741,N_21620);
or U26009 (N_26009,N_23795,N_22709);
xnor U26010 (N_26010,N_23643,N_21753);
nand U26011 (N_26011,N_24316,N_22348);
nand U26012 (N_26012,N_23399,N_23604);
and U26013 (N_26013,N_21420,N_22161);
xor U26014 (N_26014,N_20560,N_24963);
or U26015 (N_26015,N_23248,N_23228);
nor U26016 (N_26016,N_20469,N_23487);
or U26017 (N_26017,N_21804,N_23433);
and U26018 (N_26018,N_22892,N_22286);
xnor U26019 (N_26019,N_20032,N_23348);
xor U26020 (N_26020,N_24594,N_23941);
or U26021 (N_26021,N_22065,N_20070);
nor U26022 (N_26022,N_21801,N_21334);
nand U26023 (N_26023,N_20478,N_20067);
or U26024 (N_26024,N_24330,N_23865);
and U26025 (N_26025,N_24398,N_21055);
nand U26026 (N_26026,N_20009,N_23003);
nor U26027 (N_26027,N_24477,N_20619);
and U26028 (N_26028,N_22876,N_20443);
or U26029 (N_26029,N_24878,N_21867);
or U26030 (N_26030,N_21692,N_20556);
or U26031 (N_26031,N_24045,N_21809);
nand U26032 (N_26032,N_20432,N_24817);
and U26033 (N_26033,N_23931,N_24051);
nor U26034 (N_26034,N_22216,N_20705);
nor U26035 (N_26035,N_21965,N_22758);
and U26036 (N_26036,N_22317,N_22746);
or U26037 (N_26037,N_23565,N_22315);
nand U26038 (N_26038,N_21335,N_23229);
or U26039 (N_26039,N_20707,N_24278);
or U26040 (N_26040,N_23460,N_21128);
nor U26041 (N_26041,N_22866,N_20426);
or U26042 (N_26042,N_22731,N_20772);
or U26043 (N_26043,N_20301,N_24745);
nand U26044 (N_26044,N_22563,N_22705);
nand U26045 (N_26045,N_23468,N_20321);
and U26046 (N_26046,N_24382,N_21249);
and U26047 (N_26047,N_23313,N_22118);
or U26048 (N_26048,N_24752,N_21799);
and U26049 (N_26049,N_22664,N_23481);
xnor U26050 (N_26050,N_21300,N_22959);
or U26051 (N_26051,N_21182,N_24059);
or U26052 (N_26052,N_21118,N_22436);
and U26053 (N_26053,N_23227,N_24109);
or U26054 (N_26054,N_22692,N_24895);
nor U26055 (N_26055,N_20056,N_23623);
or U26056 (N_26056,N_24394,N_22097);
or U26057 (N_26057,N_24100,N_24359);
nor U26058 (N_26058,N_23977,N_20132);
and U26059 (N_26059,N_24899,N_22432);
nor U26060 (N_26060,N_22570,N_24872);
nand U26061 (N_26061,N_23008,N_21612);
or U26062 (N_26062,N_24105,N_23802);
or U26063 (N_26063,N_22803,N_22299);
nor U26064 (N_26064,N_23698,N_22021);
nand U26065 (N_26065,N_24068,N_23120);
nand U26066 (N_26066,N_21446,N_22982);
nand U26067 (N_26067,N_21567,N_23493);
nand U26068 (N_26068,N_24339,N_20776);
nand U26069 (N_26069,N_24210,N_22748);
nor U26070 (N_26070,N_20572,N_23192);
or U26071 (N_26071,N_21913,N_22927);
nand U26072 (N_26072,N_22379,N_23119);
nor U26073 (N_26073,N_20178,N_24916);
xnor U26074 (N_26074,N_24284,N_23899);
or U26075 (N_26075,N_22628,N_23020);
or U26076 (N_26076,N_20437,N_22801);
xor U26077 (N_26077,N_20363,N_21126);
nor U26078 (N_26078,N_22697,N_21195);
nand U26079 (N_26079,N_21793,N_20971);
and U26080 (N_26080,N_24323,N_22212);
and U26081 (N_26081,N_20689,N_22458);
nor U26082 (N_26082,N_24971,N_24994);
and U26083 (N_26083,N_24541,N_22465);
nand U26084 (N_26084,N_23253,N_24587);
or U26085 (N_26085,N_20810,N_23856);
nor U26086 (N_26086,N_23731,N_21329);
or U26087 (N_26087,N_21897,N_21687);
xnor U26088 (N_26088,N_21480,N_21745);
or U26089 (N_26089,N_22079,N_23846);
nand U26090 (N_26090,N_22819,N_22126);
and U26091 (N_26091,N_23919,N_24464);
or U26092 (N_26092,N_23035,N_22841);
or U26093 (N_26093,N_20323,N_24695);
xor U26094 (N_26094,N_21754,N_24680);
nand U26095 (N_26095,N_23718,N_22832);
xnor U26096 (N_26096,N_23069,N_24517);
nor U26097 (N_26097,N_23336,N_22155);
xor U26098 (N_26098,N_20984,N_21661);
xor U26099 (N_26099,N_20605,N_22911);
and U26100 (N_26100,N_21440,N_21071);
xnor U26101 (N_26101,N_20499,N_23902);
nor U26102 (N_26102,N_20863,N_24286);
nor U26103 (N_26103,N_23653,N_21822);
nor U26104 (N_26104,N_21027,N_21743);
nor U26105 (N_26105,N_20409,N_23469);
xnor U26106 (N_26106,N_24379,N_20942);
nand U26107 (N_26107,N_20865,N_23567);
and U26108 (N_26108,N_22567,N_22120);
and U26109 (N_26109,N_23148,N_23924);
or U26110 (N_26110,N_23991,N_21321);
nand U26111 (N_26111,N_24441,N_21201);
and U26112 (N_26112,N_21167,N_22475);
or U26113 (N_26113,N_24699,N_24276);
or U26114 (N_26114,N_22179,N_21024);
or U26115 (N_26115,N_22478,N_20851);
nor U26116 (N_26116,N_21638,N_23617);
xor U26117 (N_26117,N_20974,N_24363);
nor U26118 (N_26118,N_23305,N_20107);
nor U26119 (N_26119,N_24833,N_23266);
and U26120 (N_26120,N_23437,N_20938);
and U26121 (N_26121,N_22018,N_21288);
nor U26122 (N_26122,N_22224,N_23027);
xnor U26123 (N_26123,N_24211,N_23179);
and U26124 (N_26124,N_23454,N_20423);
or U26125 (N_26125,N_22308,N_24637);
and U26126 (N_26126,N_20787,N_23855);
and U26127 (N_26127,N_22633,N_23461);
or U26128 (N_26128,N_23593,N_20687);
or U26129 (N_26129,N_23328,N_24186);
and U26130 (N_26130,N_20164,N_23812);
or U26131 (N_26131,N_21790,N_22561);
nor U26132 (N_26132,N_23447,N_23007);
nand U26133 (N_26133,N_21033,N_23882);
nor U26134 (N_26134,N_24858,N_20982);
and U26135 (N_26135,N_23484,N_21381);
or U26136 (N_26136,N_24273,N_20828);
and U26137 (N_26137,N_20914,N_21458);
and U26138 (N_26138,N_23168,N_22387);
and U26139 (N_26139,N_22966,N_22249);
nor U26140 (N_26140,N_23854,N_21357);
and U26141 (N_26141,N_21618,N_24664);
nand U26142 (N_26142,N_24905,N_22732);
or U26143 (N_26143,N_24888,N_23984);
nand U26144 (N_26144,N_24119,N_24540);
and U26145 (N_26145,N_23353,N_20296);
xor U26146 (N_26146,N_24095,N_21528);
or U26147 (N_26147,N_23087,N_21415);
and U26148 (N_26148,N_22835,N_20880);
and U26149 (N_26149,N_20943,N_20708);
xor U26150 (N_26150,N_24353,N_22796);
nand U26151 (N_26151,N_22259,N_24346);
xnor U26152 (N_26152,N_22334,N_24751);
or U26153 (N_26153,N_24342,N_21246);
nor U26154 (N_26154,N_23128,N_22829);
and U26155 (N_26155,N_24159,N_20532);
nand U26156 (N_26156,N_24030,N_23626);
xnor U26157 (N_26157,N_21297,N_22857);
nor U26158 (N_26158,N_24959,N_22506);
nor U26159 (N_26159,N_24002,N_21502);
and U26160 (N_26160,N_23703,N_21761);
or U26161 (N_26161,N_22840,N_22357);
nand U26162 (N_26162,N_22355,N_20005);
nor U26163 (N_26163,N_20103,N_22831);
and U26164 (N_26164,N_21581,N_20495);
and U26165 (N_26165,N_20783,N_21626);
nor U26166 (N_26166,N_22954,N_22599);
nand U26167 (N_26167,N_23400,N_21107);
xnor U26168 (N_26168,N_22049,N_21883);
nor U26169 (N_26169,N_21669,N_22533);
nor U26170 (N_26170,N_24046,N_21594);
and U26171 (N_26171,N_22956,N_21948);
nor U26172 (N_26172,N_22451,N_22277);
xnor U26173 (N_26173,N_20715,N_22417);
nor U26174 (N_26174,N_23365,N_22297);
xor U26175 (N_26175,N_20854,N_21066);
and U26176 (N_26176,N_21772,N_24500);
and U26177 (N_26177,N_20146,N_20734);
xor U26178 (N_26178,N_23618,N_22760);
nand U26179 (N_26179,N_24459,N_21766);
and U26180 (N_26180,N_23867,N_24743);
and U26181 (N_26181,N_20377,N_22104);
nand U26182 (N_26182,N_21716,N_20490);
nand U26183 (N_26183,N_24952,N_21169);
xor U26184 (N_26184,N_23440,N_24640);
nor U26185 (N_26185,N_24463,N_20997);
nor U26186 (N_26186,N_23004,N_22874);
and U26187 (N_26187,N_23247,N_24979);
and U26188 (N_26188,N_20671,N_24040);
nand U26189 (N_26189,N_24047,N_20233);
and U26190 (N_26190,N_24918,N_21782);
nor U26191 (N_26191,N_20791,N_24798);
or U26192 (N_26192,N_21360,N_23216);
or U26193 (N_26193,N_22017,N_24856);
or U26194 (N_26194,N_23898,N_20395);
nand U26195 (N_26195,N_20895,N_23431);
nor U26196 (N_26196,N_22510,N_21125);
or U26197 (N_26197,N_23432,N_23605);
or U26198 (N_26198,N_20421,N_20473);
nand U26199 (N_26199,N_21887,N_21908);
nand U26200 (N_26200,N_24980,N_21324);
nand U26201 (N_26201,N_24036,N_24366);
nor U26202 (N_26202,N_24654,N_20609);
nand U26203 (N_26203,N_20515,N_21042);
and U26204 (N_26204,N_21939,N_22029);
and U26205 (N_26205,N_24847,N_20349);
and U26206 (N_26206,N_24957,N_20226);
nor U26207 (N_26207,N_24809,N_22755);
and U26208 (N_26208,N_24958,N_22781);
or U26209 (N_26209,N_24397,N_20729);
or U26210 (N_26210,N_20732,N_21468);
and U26211 (N_26211,N_21148,N_24652);
or U26212 (N_26212,N_24470,N_23215);
or U26213 (N_26213,N_22200,N_20951);
nand U26214 (N_26214,N_20193,N_22319);
and U26215 (N_26215,N_22220,N_24087);
or U26216 (N_26216,N_23757,N_22084);
nor U26217 (N_26217,N_24475,N_22670);
and U26218 (N_26218,N_22843,N_23579);
nand U26219 (N_26219,N_20357,N_23388);
nand U26220 (N_26220,N_23750,N_24443);
nand U26221 (N_26221,N_21040,N_23068);
or U26222 (N_26222,N_20769,N_23341);
and U26223 (N_26223,N_21005,N_23876);
nor U26224 (N_26224,N_21663,N_23570);
nand U26225 (N_26225,N_23144,N_24588);
nor U26226 (N_26226,N_20118,N_22813);
nor U26227 (N_26227,N_21054,N_22238);
and U26228 (N_26228,N_21450,N_22046);
and U26229 (N_26229,N_22558,N_22280);
and U26230 (N_26230,N_23627,N_21007);
and U26231 (N_26231,N_21683,N_24291);
nor U26232 (N_26232,N_22112,N_21242);
nand U26233 (N_26233,N_20192,N_21971);
nor U26234 (N_26234,N_20259,N_23592);
and U26235 (N_26235,N_20069,N_21578);
nor U26236 (N_26236,N_21208,N_23466);
nor U26237 (N_26237,N_23980,N_23615);
nand U26238 (N_26238,N_24007,N_21041);
nor U26239 (N_26239,N_23922,N_22177);
nand U26240 (N_26240,N_23845,N_22392);
and U26241 (N_26241,N_23564,N_21477);
and U26242 (N_26242,N_22143,N_21139);
and U26243 (N_26243,N_21406,N_21226);
nand U26244 (N_26244,N_20128,N_22861);
nor U26245 (N_26245,N_21271,N_24992);
xor U26246 (N_26246,N_23816,N_22992);
nand U26247 (N_26247,N_24857,N_20941);
nor U26248 (N_26248,N_22268,N_24929);
or U26249 (N_26249,N_24153,N_20020);
xnor U26250 (N_26250,N_22144,N_21695);
nor U26251 (N_26251,N_20728,N_22902);
nor U26252 (N_26252,N_22582,N_20154);
nor U26253 (N_26253,N_20912,N_24259);
nand U26254 (N_26254,N_24991,N_22600);
nand U26255 (N_26255,N_23084,N_21144);
nor U26256 (N_26256,N_20508,N_23345);
and U26257 (N_26257,N_20325,N_22435);
and U26258 (N_26258,N_21529,N_20853);
or U26259 (N_26259,N_23425,N_21127);
nand U26260 (N_26260,N_22122,N_23689);
and U26261 (N_26261,N_24887,N_20297);
and U26262 (N_26262,N_23552,N_20379);
nand U26263 (N_26263,N_24572,N_24234);
and U26264 (N_26264,N_24006,N_23498);
nor U26265 (N_26265,N_21871,N_21328);
and U26266 (N_26266,N_24860,N_20453);
or U26267 (N_26267,N_21744,N_21052);
xor U26268 (N_26268,N_20235,N_21513);
nand U26269 (N_26269,N_24462,N_22750);
nand U26270 (N_26270,N_23884,N_20282);
or U26271 (N_26271,N_22219,N_20552);
or U26272 (N_26272,N_24195,N_20672);
or U26273 (N_26273,N_20236,N_22908);
or U26274 (N_26274,N_20502,N_22653);
or U26275 (N_26275,N_23029,N_24942);
nor U26276 (N_26276,N_24416,N_22555);
or U26277 (N_26277,N_20241,N_20416);
or U26278 (N_26278,N_24589,N_24107);
nor U26279 (N_26279,N_22951,N_22015);
or U26280 (N_26280,N_23841,N_24823);
xor U26281 (N_26281,N_23768,N_22644);
nor U26282 (N_26282,N_21535,N_20041);
nand U26283 (N_26283,N_24925,N_21133);
and U26284 (N_26284,N_24604,N_21432);
nand U26285 (N_26285,N_24061,N_22907);
and U26286 (N_26286,N_21216,N_22185);
or U26287 (N_26287,N_21768,N_22757);
and U26288 (N_26288,N_24084,N_22833);
and U26289 (N_26289,N_23555,N_24115);
or U26290 (N_26290,N_22868,N_24094);
nand U26291 (N_26291,N_22968,N_20446);
nor U26292 (N_26292,N_24260,N_21257);
or U26293 (N_26293,N_23537,N_20149);
nand U26294 (N_26294,N_20848,N_21103);
nor U26295 (N_26295,N_21627,N_20270);
xor U26296 (N_26296,N_24090,N_20555);
nand U26297 (N_26297,N_20345,N_21937);
and U26298 (N_26298,N_21837,N_20530);
nand U26299 (N_26299,N_21982,N_21185);
nand U26300 (N_26300,N_23171,N_20397);
nor U26301 (N_26301,N_22785,N_21277);
nor U26302 (N_26302,N_22237,N_20393);
nor U26303 (N_26303,N_21274,N_21881);
nand U26304 (N_26304,N_20792,N_20328);
and U26305 (N_26305,N_21213,N_20520);
and U26306 (N_26306,N_20035,N_21508);
and U26307 (N_26307,N_20569,N_20448);
nand U26308 (N_26308,N_22372,N_20153);
nand U26309 (N_26309,N_24542,N_23774);
nand U26310 (N_26310,N_20100,N_24027);
nand U26311 (N_26311,N_22231,N_21114);
nand U26312 (N_26312,N_23926,N_20261);
nor U26313 (N_26313,N_22377,N_20384);
and U26314 (N_26314,N_22437,N_20539);
nor U26315 (N_26315,N_24791,N_23327);
and U26316 (N_26316,N_21568,N_22145);
nand U26317 (N_26317,N_23445,N_20300);
nand U26318 (N_26318,N_23904,N_22824);
or U26319 (N_26319,N_24915,N_21444);
or U26320 (N_26320,N_22463,N_22811);
xnor U26321 (N_26321,N_23628,N_24850);
and U26322 (N_26322,N_24255,N_21940);
and U26323 (N_26323,N_23749,N_22571);
nand U26324 (N_26324,N_22551,N_21059);
or U26325 (N_26325,N_20568,N_21515);
nor U26326 (N_26326,N_21981,N_22213);
nand U26327 (N_26327,N_21774,N_21375);
or U26328 (N_26328,N_20760,N_22209);
nor U26329 (N_26329,N_22467,N_23847);
nor U26330 (N_26330,N_20986,N_20866);
or U26331 (N_26331,N_23129,N_23324);
nand U26332 (N_26332,N_22394,N_24781);
nand U26333 (N_26333,N_21873,N_22923);
xor U26334 (N_26334,N_24600,N_22933);
xor U26335 (N_26335,N_23390,N_21684);
nand U26336 (N_26336,N_21792,N_23350);
or U26337 (N_26337,N_20903,N_21848);
or U26338 (N_26338,N_22233,N_22885);
nor U26339 (N_26339,N_24764,N_24499);
xnor U26340 (N_26340,N_24851,N_22701);
nor U26341 (N_26341,N_20987,N_21190);
nand U26342 (N_26342,N_22858,N_20450);
nor U26343 (N_26343,N_20656,N_22462);
or U26344 (N_26344,N_22573,N_21823);
or U26345 (N_26345,N_23741,N_22579);
or U26346 (N_26346,N_24118,N_20228);
xor U26347 (N_26347,N_23151,N_21181);
nor U26348 (N_26348,N_20364,N_20959);
xor U26349 (N_26349,N_24305,N_24515);
or U26350 (N_26350,N_20501,N_24415);
or U26351 (N_26351,N_22899,N_23713);
and U26352 (N_26352,N_23942,N_22400);
nand U26353 (N_26353,N_24386,N_21552);
or U26354 (N_26354,N_24920,N_20221);
or U26355 (N_26355,N_23208,N_24151);
or U26356 (N_26356,N_22110,N_20223);
or U26357 (N_26357,N_24136,N_22362);
and U26358 (N_26358,N_24064,N_22407);
nand U26359 (N_26359,N_20336,N_21719);
nor U26360 (N_26360,N_20822,N_24200);
and U26361 (N_26361,N_21117,N_21064);
xnor U26362 (N_26362,N_23200,N_24659);
nor U26363 (N_26363,N_23285,N_22276);
nand U26364 (N_26364,N_24358,N_24789);
or U26365 (N_26365,N_20861,N_21106);
and U26366 (N_26366,N_20356,N_22494);
xnor U26367 (N_26367,N_22977,N_21927);
or U26368 (N_26368,N_20806,N_23005);
nand U26369 (N_26369,N_23975,N_20084);
xor U26370 (N_26370,N_22624,N_23201);
nor U26371 (N_26371,N_20264,N_24599);
or U26372 (N_26372,N_24156,N_24618);
nor U26373 (N_26373,N_23183,N_22834);
xor U26374 (N_26374,N_24543,N_23675);
and U26375 (N_26375,N_21039,N_20587);
or U26376 (N_26376,N_24496,N_23221);
or U26377 (N_26377,N_23622,N_20425);
nand U26378 (N_26378,N_21880,N_22250);
or U26379 (N_26379,N_23665,N_21378);
nand U26380 (N_26380,N_20303,N_20287);
nor U26381 (N_26381,N_21469,N_24703);
or U26382 (N_26382,N_20980,N_21086);
nor U26383 (N_26383,N_24603,N_20474);
nor U26384 (N_26384,N_24414,N_21264);
or U26385 (N_26385,N_21813,N_20378);
and U26386 (N_26386,N_24717,N_23293);
and U26387 (N_26387,N_21235,N_23265);
nand U26388 (N_26388,N_21755,N_20775);
or U26389 (N_26389,N_22335,N_24283);
or U26390 (N_26390,N_21173,N_23723);
nand U26391 (N_26391,N_24669,N_24726);
nand U26392 (N_26392,N_22454,N_23174);
nand U26393 (N_26393,N_22127,N_20858);
nand U26394 (N_26394,N_20090,N_22606);
nand U26395 (N_26395,N_24787,N_23472);
nor U26396 (N_26396,N_22008,N_24103);
and U26397 (N_26397,N_20953,N_21747);
nor U26398 (N_26398,N_24913,N_21705);
and U26399 (N_26399,N_24322,N_21901);
xor U26400 (N_26400,N_23089,N_21929);
and U26401 (N_26401,N_24930,N_24735);
nor U26402 (N_26402,N_20635,N_21476);
nand U26403 (N_26403,N_21856,N_24557);
nor U26404 (N_26404,N_20119,N_20847);
and U26405 (N_26405,N_20359,N_22578);
nand U26406 (N_26406,N_22984,N_20075);
or U26407 (N_26407,N_23048,N_24921);
or U26408 (N_26408,N_22071,N_20412);
or U26409 (N_26409,N_22952,N_20441);
and U26410 (N_26410,N_23094,N_21877);
and U26411 (N_26411,N_22948,N_21160);
and U26412 (N_26412,N_24165,N_24667);
nor U26413 (N_26413,N_24623,N_20456);
or U26414 (N_26414,N_23231,N_23541);
or U26415 (N_26415,N_20578,N_22947);
xnor U26416 (N_26416,N_23582,N_20266);
and U26417 (N_26417,N_23864,N_24765);
nand U26418 (N_26418,N_23209,N_21960);
nand U26419 (N_26419,N_23581,N_22062);
nor U26420 (N_26420,N_21014,N_23820);
nand U26421 (N_26421,N_22598,N_23657);
xor U26422 (N_26422,N_23636,N_23735);
nand U26423 (N_26423,N_21765,N_22088);
nor U26424 (N_26424,N_20926,N_24758);
and U26425 (N_26425,N_21311,N_23088);
nor U26426 (N_26426,N_23448,N_20836);
and U26427 (N_26427,N_23118,N_24638);
nor U26428 (N_26428,N_23789,N_23938);
nand U26429 (N_26429,N_24268,N_24802);
and U26430 (N_26430,N_21220,N_22725);
nand U26431 (N_26431,N_23001,N_22779);
nand U26432 (N_26432,N_22105,N_21798);
nor U26433 (N_26433,N_20316,N_23815);
and U26434 (N_26434,N_23699,N_22030);
and U26435 (N_26435,N_23211,N_21966);
nor U26436 (N_26436,N_22309,N_22609);
nor U26437 (N_26437,N_24054,N_23387);
and U26438 (N_26438,N_23668,N_24670);
nand U26439 (N_26439,N_21392,N_23839);
and U26440 (N_26440,N_20365,N_20189);
xor U26441 (N_26441,N_22546,N_20700);
and U26442 (N_26442,N_20265,N_22313);
nor U26443 (N_26443,N_21196,N_23297);
or U26444 (N_26444,N_23974,N_20827);
xnor U26445 (N_26445,N_21400,N_22412);
nand U26446 (N_26446,N_24581,N_20900);
or U26447 (N_26447,N_22699,N_22370);
nand U26448 (N_26448,N_21530,N_21876);
nand U26449 (N_26449,N_21806,N_20449);
nor U26450 (N_26450,N_20663,N_23354);
or U26451 (N_26451,N_24945,N_20079);
nor U26452 (N_26452,N_21866,N_23807);
and U26453 (N_26453,N_23667,N_23077);
and U26454 (N_26454,N_23310,N_24712);
nor U26455 (N_26455,N_23644,N_20480);
and U26456 (N_26456,N_24184,N_21067);
or U26457 (N_26457,N_21001,N_21272);
nor U26458 (N_26458,N_22291,N_21193);
or U26459 (N_26459,N_22777,N_21141);
xor U26460 (N_26460,N_22269,N_21466);
nand U26461 (N_26461,N_23509,N_21899);
or U26462 (N_26462,N_22025,N_21797);
nor U26463 (N_26463,N_21587,N_22075);
nand U26464 (N_26464,N_24583,N_22428);
or U26465 (N_26465,N_22710,N_23126);
and U26466 (N_26466,N_22922,N_20405);
and U26467 (N_26467,N_23632,N_23779);
xnor U26468 (N_26468,N_22790,N_20924);
nand U26469 (N_26469,N_22253,N_24749);
nand U26470 (N_26470,N_22865,N_21791);
nor U26471 (N_26471,N_22888,N_22304);
and U26472 (N_26472,N_20589,N_22953);
nor U26473 (N_26473,N_20950,N_20115);
or U26474 (N_26474,N_22028,N_21174);
nor U26475 (N_26475,N_23631,N_23184);
and U26476 (N_26476,N_20210,N_23204);
xnor U26477 (N_26477,N_24472,N_20981);
nand U26478 (N_26478,N_21407,N_20320);
nor U26479 (N_26479,N_24777,N_20979);
or U26480 (N_26480,N_21651,N_23588);
xnor U26481 (N_26481,N_22839,N_23928);
nor U26482 (N_26482,N_24484,N_20279);
nand U26483 (N_26483,N_23953,N_23518);
nor U26484 (N_26484,N_23112,N_24171);
nor U26485 (N_26485,N_20921,N_22485);
nand U26486 (N_26486,N_23678,N_20524);
xnor U26487 (N_26487,N_24257,N_24449);
and U26488 (N_26488,N_24744,N_20454);
nor U26489 (N_26489,N_22285,N_20112);
xor U26490 (N_26490,N_22260,N_23527);
or U26491 (N_26491,N_21289,N_22696);
and U26492 (N_26492,N_24101,N_24015);
and U26493 (N_26493,N_23547,N_21339);
nor U26494 (N_26494,N_23827,N_21402);
nor U26495 (N_26495,N_21857,N_21090);
and U26496 (N_26496,N_24523,N_24814);
or U26497 (N_26497,N_22496,N_23822);
or U26498 (N_26498,N_20255,N_21341);
or U26499 (N_26499,N_20988,N_23397);
or U26500 (N_26500,N_21199,N_23279);
or U26501 (N_26501,N_24926,N_20142);
nand U26502 (N_26502,N_22639,N_23176);
and U26503 (N_26503,N_23054,N_22180);
nand U26504 (N_26504,N_21934,N_24321);
and U26505 (N_26505,N_22034,N_22749);
or U26506 (N_26506,N_20996,N_24783);
nand U26507 (N_26507,N_24190,N_23235);
nand U26508 (N_26508,N_21536,N_24898);
or U26509 (N_26509,N_21658,N_24426);
or U26510 (N_26510,N_21322,N_21892);
nor U26511 (N_26511,N_20857,N_23679);
xnor U26512 (N_26512,N_23323,N_22786);
xor U26513 (N_26513,N_24774,N_24424);
or U26514 (N_26514,N_22643,N_24492);
or U26515 (N_26515,N_23024,N_21284);
or U26516 (N_26516,N_23172,N_20976);
xor U26517 (N_26517,N_24826,N_24230);
nand U26518 (N_26518,N_21976,N_21652);
nand U26519 (N_26519,N_22434,N_20309);
nand U26520 (N_26520,N_23669,N_24668);
nand U26521 (N_26521,N_22684,N_21851);
nor U26522 (N_26522,N_21894,N_20082);
or U26523 (N_26523,N_24116,N_23655);
and U26524 (N_26524,N_22474,N_22967);
and U26525 (N_26525,N_23299,N_20768);
xor U26526 (N_26526,N_20207,N_24452);
nor U26527 (N_26527,N_23082,N_24527);
nand U26528 (N_26528,N_21760,N_23999);
and U26529 (N_26529,N_22556,N_22698);
xor U26530 (N_26530,N_24605,N_21779);
nor U26531 (N_26531,N_20353,N_20811);
or U26532 (N_26532,N_24569,N_24168);
nand U26533 (N_26533,N_20855,N_21109);
and U26534 (N_26534,N_20716,N_20554);
or U26535 (N_26535,N_23490,N_20516);
nand U26536 (N_26536,N_24264,N_23426);
or U26537 (N_26537,N_20492,N_21171);
nand U26538 (N_26538,N_22812,N_20901);
xnor U26539 (N_26539,N_23897,N_22630);
and U26540 (N_26540,N_24656,N_20208);
or U26541 (N_26541,N_24884,N_24885);
nand U26542 (N_26542,N_22415,N_21434);
and U26543 (N_26543,N_24890,N_22926);
nor U26544 (N_26544,N_22721,N_20049);
and U26545 (N_26545,N_21987,N_20786);
nor U26546 (N_26546,N_20648,N_22711);
or U26547 (N_26547,N_23263,N_23972);
or U26548 (N_26548,N_22072,N_22419);
or U26549 (N_26549,N_24431,N_20043);
and U26550 (N_26550,N_21426,N_24335);
and U26551 (N_26551,N_24780,N_24302);
and U26552 (N_26552,N_22193,N_22278);
or U26553 (N_26553,N_23170,N_22331);
or U26554 (N_26554,N_20201,N_22418);
nand U26555 (N_26555,N_21912,N_22847);
nand U26556 (N_26556,N_23727,N_23264);
or U26557 (N_26557,N_21417,N_20445);
or U26558 (N_26558,N_22971,N_22941);
nor U26559 (N_26559,N_22168,N_22946);
or U26560 (N_26560,N_22515,N_24839);
and U26561 (N_26561,N_24653,N_21606);
nand U26562 (N_26562,N_24534,N_21044);
nand U26563 (N_26563,N_21352,N_22450);
nand U26564 (N_26564,N_21457,N_21408);
nand U26565 (N_26565,N_21601,N_22380);
and U26566 (N_26566,N_21097,N_22414);
nand U26567 (N_26567,N_24334,N_24063);
nor U26568 (N_26568,N_21081,N_21346);
and U26569 (N_26569,N_24209,N_23125);
or U26570 (N_26570,N_20803,N_23153);
and U26571 (N_26571,N_20249,N_23182);
nand U26572 (N_26572,N_23778,N_22350);
nor U26573 (N_26573,N_20402,N_20852);
nand U26574 (N_26574,N_21653,N_20487);
and U26575 (N_26575,N_22795,N_22039);
or U26576 (N_26576,N_23952,N_20750);
nand U26577 (N_26577,N_22381,N_22560);
nor U26578 (N_26578,N_22584,N_20691);
xnor U26579 (N_26579,N_23146,N_20158);
nand U26580 (N_26580,N_20029,N_20087);
and U26581 (N_26581,N_24070,N_21261);
or U26582 (N_26582,N_21517,N_22517);
nor U26583 (N_26583,N_23040,N_22823);
and U26584 (N_26584,N_24246,N_22680);
or U26585 (N_26585,N_24252,N_22574);
nand U26586 (N_26586,N_21936,N_22443);
nand U26587 (N_26587,N_22774,N_20392);
or U26588 (N_26588,N_24347,N_24369);
xnor U26589 (N_26589,N_22634,N_24988);
and U26590 (N_26590,N_23057,N_24655);
nand U26591 (N_26591,N_21050,N_21554);
or U26592 (N_26592,N_20693,N_21802);
nand U26593 (N_26593,N_22789,N_21389);
and U26594 (N_26594,N_23959,N_20625);
xnor U26595 (N_26595,N_24243,N_20779);
and U26596 (N_26596,N_20340,N_23062);
nand U26597 (N_26597,N_24023,N_22326);
nor U26598 (N_26598,N_20311,N_22066);
nand U26599 (N_26599,N_23693,N_24274);
nor U26600 (N_26600,N_23371,N_21712);
and U26601 (N_26601,N_22240,N_22800);
nor U26602 (N_26602,N_23379,N_23755);
or U26603 (N_26603,N_23805,N_21878);
or U26604 (N_26604,N_21562,N_23515);
nor U26605 (N_26605,N_23219,N_20230);
nand U26606 (N_26606,N_24142,N_24148);
nand U26607 (N_26607,N_22480,N_21318);
or U26608 (N_26608,N_20566,N_24676);
nand U26609 (N_26609,N_22615,N_20875);
and U26610 (N_26610,N_24042,N_22592);
xor U26611 (N_26611,N_22878,N_20665);
and U26612 (N_26612,N_23398,N_20799);
and U26613 (N_26613,N_20628,N_23244);
and U26614 (N_26614,N_23937,N_22314);
xnor U26615 (N_26615,N_21505,N_22089);
nor U26616 (N_26616,N_20291,N_23814);
nor U26617 (N_26617,N_20334,N_23681);
or U26618 (N_26618,N_20095,N_24960);
and U26619 (N_26619,N_23278,N_24106);
nor U26620 (N_26620,N_24375,N_20085);
or U26621 (N_26621,N_24324,N_21858);
nand U26622 (N_26622,N_24263,N_23833);
and U26623 (N_26623,N_24772,N_24855);
nor U26624 (N_26624,N_22235,N_23304);
nor U26625 (N_26625,N_22295,N_20318);
nor U26626 (N_26626,N_24480,N_22985);
or U26627 (N_26627,N_22094,N_24708);
and U26628 (N_26628,N_23869,N_22106);
or U26629 (N_26629,N_23701,N_24504);
and U26630 (N_26630,N_23965,N_21265);
nand U26631 (N_26631,N_20745,N_20859);
xor U26632 (N_26632,N_21353,N_22221);
nand U26633 (N_26633,N_22805,N_23405);
nor U26634 (N_26634,N_23715,N_24117);
nand U26635 (N_26635,N_22013,N_24429);
nor U26636 (N_26636,N_24827,N_24085);
or U26637 (N_26637,N_20047,N_22289);
nor U26638 (N_26638,N_21165,N_24713);
and U26639 (N_26639,N_21631,N_20004);
or U26640 (N_26640,N_21331,N_20074);
or U26641 (N_26641,N_22729,N_20315);
nand U26642 (N_26642,N_22682,N_24684);
nand U26643 (N_26643,N_21888,N_24404);
or U26644 (N_26644,N_20576,N_21585);
and U26645 (N_26645,N_23485,N_23954);
xor U26646 (N_26646,N_20177,N_21217);
nand U26647 (N_26647,N_23989,N_20717);
nand U26648 (N_26648,N_21951,N_20404);
nand U26649 (N_26649,N_20023,N_24607);
or U26650 (N_26650,N_21009,N_20598);
nand U26651 (N_26651,N_24681,N_21008);
nor U26652 (N_26652,N_22007,N_20565);
nor U26653 (N_26653,N_24368,N_24641);
and U26654 (N_26654,N_22541,N_23212);
nand U26655 (N_26655,N_21830,N_22720);
nand U26656 (N_26656,N_24590,N_23256);
nand U26657 (N_26657,N_24891,N_20076);
and U26658 (N_26658,N_22949,N_20186);
and U26659 (N_26659,N_24558,N_24688);
nand U26660 (N_26660,N_20983,N_22780);
nand U26661 (N_26661,N_21596,N_24966);
and U26662 (N_26662,N_24292,N_22601);
nand U26663 (N_26663,N_23502,N_20970);
nor U26664 (N_26664,N_20756,N_22502);
and U26665 (N_26665,N_24467,N_24317);
and U26666 (N_26666,N_23394,N_21842);
nor U26667 (N_26667,N_20121,N_23187);
nor U26668 (N_26668,N_23995,N_23232);
nand U26669 (N_26669,N_24254,N_24004);
and U26670 (N_26670,N_21490,N_22820);
nor U26671 (N_26671,N_24204,N_24901);
nand U26672 (N_26672,N_22593,N_24615);
nor U26673 (N_26673,N_23022,N_24938);
nand U26674 (N_26674,N_23763,N_23662);
or U26675 (N_26675,N_20497,N_22055);
nor U26676 (N_26676,N_22808,N_24889);
nand U26677 (N_26677,N_20621,N_24205);
and U26678 (N_26678,N_21197,N_20052);
nand U26679 (N_26679,N_20258,N_24663);
nand U26680 (N_26680,N_22425,N_24318);
nor U26681 (N_26681,N_23890,N_21058);
or U26682 (N_26682,N_22115,N_24365);
nor U26683 (N_26683,N_24965,N_24411);
nor U26684 (N_26684,N_23946,N_22655);
nand U26685 (N_26685,N_20380,N_22588);
nor U26686 (N_26686,N_24631,N_22783);
nand U26687 (N_26687,N_23506,N_21396);
nor U26688 (N_26688,N_21482,N_23138);
nor U26689 (N_26689,N_20350,N_24771);
nor U26690 (N_26690,N_21487,N_23156);
and U26691 (N_26691,N_21732,N_22068);
or U26692 (N_26692,N_21603,N_21628);
nand U26693 (N_26693,N_22248,N_21852);
or U26694 (N_26694,N_21364,N_22869);
nand U26695 (N_26695,N_24595,N_23930);
nand U26696 (N_26696,N_23831,N_23728);
and U26697 (N_26697,N_22564,N_22077);
xor U26698 (N_26698,N_21672,N_21483);
and U26699 (N_26699,N_22188,N_21484);
nand U26700 (N_26700,N_21659,N_23011);
nor U26701 (N_26701,N_22187,N_20106);
and U26702 (N_26702,N_22691,N_24702);
and U26703 (N_26703,N_23520,N_22500);
or U26704 (N_26704,N_21259,N_23002);
and U26705 (N_26705,N_23226,N_22138);
nor U26706 (N_26706,N_23638,N_22420);
xnor U26707 (N_26707,N_22421,N_21051);
xor U26708 (N_26708,N_21061,N_22979);
or U26709 (N_26709,N_21200,N_22910);
nor U26710 (N_26710,N_24537,N_21269);
nor U26711 (N_26711,N_20342,N_22376);
xnor U26712 (N_26712,N_20531,N_24081);
xnor U26713 (N_26713,N_23157,N_20674);
nand U26714 (N_26714,N_23479,N_24425);
or U26715 (N_26715,N_24020,N_22449);
and U26716 (N_26716,N_21844,N_20696);
nand U26717 (N_26717,N_24625,N_21553);
nor U26718 (N_26718,N_23589,N_20733);
and U26719 (N_26719,N_20843,N_21371);
or U26720 (N_26720,N_21060,N_22149);
nand U26721 (N_26721,N_23775,N_20747);
nor U26722 (N_26722,N_23408,N_23136);
nor U26723 (N_26723,N_20234,N_20245);
nand U26724 (N_26724,N_23444,N_22070);
nand U26725 (N_26725,N_22552,N_22123);
and U26726 (N_26726,N_21872,N_21398);
and U26727 (N_26727,N_23740,N_21292);
and U26728 (N_26728,N_21232,N_20276);
xnor U26729 (N_26729,N_21391,N_20367);
and U26730 (N_26730,N_24812,N_24715);
nor U26731 (N_26731,N_20780,N_24241);
and U26732 (N_26732,N_24993,N_23039);
nand U26733 (N_26733,N_20298,N_20682);
nor U26734 (N_26734,N_24082,N_22538);
xnor U26735 (N_26735,N_23110,N_21879);
and U26736 (N_26736,N_23462,N_24928);
and U26737 (N_26737,N_24692,N_20591);
nor U26738 (N_26738,N_23659,N_21922);
nand U26739 (N_26739,N_23046,N_20679);
and U26740 (N_26740,N_23335,N_23273);
xnor U26741 (N_26741,N_21783,N_23061);
xor U26742 (N_26742,N_24877,N_24868);
and U26743 (N_26743,N_20541,N_20559);
nand U26744 (N_26744,N_21491,N_23367);
nand U26745 (N_26745,N_24535,N_20522);
and U26746 (N_26746,N_21916,N_20992);
nor U26747 (N_26747,N_23948,N_23391);
and U26748 (N_26748,N_20546,N_21239);
xor U26749 (N_26749,N_24548,N_20548);
nor U26750 (N_26750,N_24725,N_23234);
and U26751 (N_26751,N_21023,N_23584);
xor U26752 (N_26752,N_20969,N_20514);
or U26753 (N_26753,N_21369,N_21935);
and U26754 (N_26754,N_20805,N_23534);
or U26755 (N_26755,N_21228,N_20600);
nor U26756 (N_26756,N_20856,N_24698);
or U26757 (N_26757,N_20889,N_23663);
nand U26758 (N_26758,N_22442,N_24705);
or U26759 (N_26759,N_21565,N_21525);
and U26760 (N_26760,N_24272,N_21808);
nand U26761 (N_26761,N_23630,N_22410);
nand U26762 (N_26762,N_23383,N_20937);
or U26763 (N_26763,N_22167,N_20840);
xnor U26764 (N_26764,N_23058,N_23482);
or U26765 (N_26765,N_23090,N_23359);
nor U26766 (N_26766,N_21438,N_22627);
nor U26767 (N_26767,N_21241,N_24630);
nor U26768 (N_26768,N_21035,N_24399);
nor U26769 (N_26769,N_23026,N_22271);
and U26770 (N_26770,N_20038,N_23705);
nand U26771 (N_26771,N_24636,N_21120);
nand U26772 (N_26772,N_20143,N_20209);
and U26773 (N_26773,N_22920,N_21070);
and U26774 (N_26774,N_22461,N_24689);
nor U26775 (N_26775,N_22724,N_22671);
or U26776 (N_26776,N_22056,N_20998);
nor U26777 (N_26777,N_20013,N_22934);
nor U26778 (N_26778,N_23287,N_22255);
nor U26779 (N_26779,N_24784,N_20573);
nor U26780 (N_26780,N_20185,N_23306);
and U26781 (N_26781,N_20439,N_21997);
nand U26782 (N_26782,N_24493,N_24661);
nor U26783 (N_26783,N_23255,N_22983);
or U26784 (N_26784,N_23843,N_24561);
nor U26785 (N_26785,N_23404,N_23143);
xnor U26786 (N_26786,N_23918,N_22762);
nor U26787 (N_26787,N_24226,N_20838);
nand U26788 (N_26788,N_24533,N_21649);
or U26789 (N_26789,N_22211,N_24602);
or U26790 (N_26790,N_24139,N_22080);
or U26791 (N_26791,N_22837,N_20535);
and U26792 (N_26792,N_24149,N_23344);
and U26793 (N_26793,N_24150,N_22223);
nor U26794 (N_26794,N_20083,N_24031);
or U26795 (N_26795,N_22246,N_20401);
and U26796 (N_26796,N_22135,N_21186);
nand U26797 (N_26797,N_21384,N_20891);
nand U26798 (N_26798,N_21642,N_22793);
and U26799 (N_26799,N_24864,N_20212);
xor U26800 (N_26800,N_21862,N_24577);
or U26801 (N_26801,N_21367,N_20447);
nor U26802 (N_26802,N_23799,N_24012);
and U26803 (N_26803,N_23422,N_23673);
nor U26804 (N_26804,N_24350,N_22738);
nand U26805 (N_26805,N_22215,N_22565);
nand U26806 (N_26806,N_23613,N_22447);
nor U26807 (N_26807,N_20054,N_22513);
nor U26808 (N_26808,N_21452,N_23065);
or U26809 (N_26809,N_23857,N_23413);
xor U26810 (N_26810,N_20993,N_20159);
and U26811 (N_26811,N_23563,N_23688);
and U26812 (N_26812,N_23940,N_20695);
or U26813 (N_26813,N_21366,N_24805);
and U26814 (N_26814,N_21327,N_21713);
or U26815 (N_26815,N_24730,N_20804);
nor U26816 (N_26816,N_23315,N_21143);
nor U26817 (N_26817,N_22886,N_22024);
xor U26818 (N_26818,N_21247,N_24658);
and U26819 (N_26819,N_21634,N_20455);
and U26820 (N_26820,N_22292,N_22988);
nand U26821 (N_26821,N_23969,N_23163);
and U26822 (N_26822,N_20759,N_22799);
nand U26823 (N_26823,N_21679,N_22165);
and U26824 (N_26824,N_23018,N_20558);
xnor U26825 (N_26825,N_20641,N_20545);
or U26826 (N_26826,N_21715,N_24141);
nor U26827 (N_26827,N_21863,N_21343);
nand U26828 (N_26828,N_21870,N_23309);
or U26829 (N_26829,N_20594,N_20496);
nand U26830 (N_26830,N_24836,N_20718);
xor U26831 (N_26831,N_20317,N_22153);
or U26832 (N_26832,N_23649,N_21583);
nor U26833 (N_26833,N_23470,N_20371);
nor U26834 (N_26834,N_22791,N_22580);
or U26835 (N_26835,N_23523,N_21921);
nand U26836 (N_26836,N_23560,N_21100);
nor U26837 (N_26837,N_22906,N_22838);
or U26838 (N_26838,N_21780,N_23098);
or U26839 (N_26839,N_23870,N_24550);
and U26840 (N_26840,N_24301,N_20002);
nor U26841 (N_26841,N_20770,N_24709);
and U26842 (N_26842,N_24584,N_24145);
nor U26843 (N_26843,N_24614,N_21421);
nor U26844 (N_26844,N_22037,N_20307);
and U26845 (N_26845,N_21522,N_24248);
nand U26846 (N_26846,N_24985,N_23765);
xor U26847 (N_26847,N_21632,N_20688);
or U26848 (N_26848,N_22036,N_21737);
xnor U26849 (N_26849,N_23395,N_21507);
xor U26850 (N_26850,N_20911,N_22344);
nor U26851 (N_26851,N_20876,N_22521);
xnor U26852 (N_26852,N_21256,N_24632);
and U26853 (N_26853,N_20098,N_24008);
xnor U26854 (N_26854,N_24810,N_20102);
nand U26855 (N_26855,N_24050,N_20355);
and U26856 (N_26856,N_21347,N_21422);
and U26857 (N_26857,N_20277,N_20698);
and U26858 (N_26858,N_20123,N_21904);
or U26859 (N_26859,N_22575,N_24438);
xnor U26860 (N_26860,N_21178,N_22041);
or U26861 (N_26861,N_22293,N_20995);
and U26862 (N_26862,N_22232,N_20250);
or U26863 (N_26863,N_20422,N_22877);
or U26864 (N_26864,N_23240,N_20948);
and U26865 (N_26865,N_20486,N_23458);
or U26866 (N_26866,N_23545,N_24140);
and U26867 (N_26867,N_20415,N_22438);
xnor U26868 (N_26868,N_23771,N_21541);
and U26869 (N_26869,N_24949,N_24298);
and U26870 (N_26870,N_20703,N_24196);
or U26871 (N_26871,N_22850,N_20215);
xor U26872 (N_26872,N_23104,N_20418);
nand U26873 (N_26873,N_24573,N_21080);
nor U26874 (N_26874,N_21430,N_20507);
nand U26875 (N_26875,N_20408,N_22243);
or U26876 (N_26876,N_23251,N_21577);
nand U26877 (N_26877,N_21486,N_23465);
nand U26878 (N_26878,N_21501,N_23355);
and U26879 (N_26879,N_21520,N_20120);
or U26880 (N_26880,N_23573,N_24972);
nand U26881 (N_26881,N_21394,N_23580);
and U26882 (N_26882,N_23683,N_22207);
nor U26883 (N_26883,N_23162,N_23093);
nor U26884 (N_26884,N_21992,N_21494);
or U26885 (N_26885,N_20163,N_20187);
or U26886 (N_26886,N_24685,N_22932);
nor U26887 (N_26887,N_20200,N_22460);
and U26888 (N_26888,N_22722,N_23102);
or U26889 (N_26889,N_23014,N_22093);
or U26890 (N_26890,N_20651,N_23451);
or U26891 (N_26891,N_24396,N_23546);
or U26892 (N_26892,N_22960,N_22202);
nor U26893 (N_26893,N_21395,N_21506);
and U26894 (N_26894,N_20796,N_20794);
nor U26895 (N_26895,N_21418,N_21636);
or U26896 (N_26896,N_21973,N_21836);
and U26897 (N_26897,N_24968,N_24125);
or U26898 (N_26898,N_22656,N_24439);
and U26899 (N_26899,N_20704,N_22413);
nor U26900 (N_26900,N_22703,N_24739);
and U26901 (N_26901,N_23512,N_22752);
xnor U26902 (N_26902,N_22716,N_23340);
or U26903 (N_26903,N_20540,N_23958);
nand U26904 (N_26904,N_23270,N_21382);
nor U26905 (N_26905,N_21942,N_20330);
or U26906 (N_26906,N_21690,N_23542);
and U26907 (N_26907,N_21810,N_23436);
nand U26908 (N_26908,N_23222,N_22744);
and U26909 (N_26909,N_21688,N_23711);
nand U26910 (N_26910,N_21675,N_24213);
nor U26911 (N_26911,N_23275,N_20348);
nor U26912 (N_26912,N_20584,N_24473);
or U26913 (N_26913,N_24380,N_24478);
nand U26914 (N_26914,N_24883,N_21464);
or U26915 (N_26915,N_24750,N_23988);
xnor U26916 (N_26916,N_21479,N_22734);
and U26917 (N_26917,N_24005,N_22305);
and U26918 (N_26918,N_24306,N_21308);
and U26919 (N_26919,N_22043,N_22499);
or U26920 (N_26920,N_21177,N_21471);
or U26921 (N_26921,N_23409,N_22935);
or U26922 (N_26922,N_20659,N_23071);
or U26923 (N_26923,N_23819,N_24428);
and U26924 (N_26924,N_24409,N_23729);
or U26925 (N_26925,N_24420,N_21574);
nand U26926 (N_26926,N_20181,N_24740);
xor U26927 (N_26927,N_24704,N_23271);
nor U26928 (N_26928,N_20372,N_20564);
nor U26929 (N_26929,N_24123,N_21229);
and U26930 (N_26930,N_23694,N_22626);
nor U26931 (N_26931,N_22893,N_23961);
and U26932 (N_26932,N_20294,N_23261);
and U26933 (N_26933,N_23858,N_22498);
nand U26934 (N_26934,N_24403,N_23585);
nor U26935 (N_26935,N_21580,N_20834);
nor U26936 (N_26936,N_21623,N_20175);
nand U26937 (N_26937,N_22352,N_23806);
or U26938 (N_26938,N_22361,N_23983);
nor U26939 (N_26939,N_24218,N_20563);
or U26940 (N_26940,N_22855,N_20376);
xnor U26941 (N_26941,N_23987,N_20147);
nand U26942 (N_26942,N_21702,N_24122);
nand U26943 (N_26943,N_23213,N_23764);
and U26944 (N_26944,N_22245,N_20459);
and U26945 (N_26945,N_24834,N_20063);
nor U26946 (N_26946,N_24894,N_23083);
and U26947 (N_26947,N_21439,N_20821);
or U26948 (N_26948,N_21317,N_24516);
xnor U26949 (N_26949,N_20675,N_24947);
xnor U26950 (N_26950,N_20072,N_20509);
or U26951 (N_26951,N_22916,N_21069);
and U26952 (N_26952,N_23499,N_21172);
nor U26953 (N_26953,N_22939,N_20973);
nor U26954 (N_26954,N_24216,N_23314);
nand U26955 (N_26955,N_23294,N_21533);
and U26956 (N_26956,N_20645,N_23590);
nor U26957 (N_26957,N_20910,N_22667);
and U26958 (N_26958,N_22208,N_24954);
and U26959 (N_26959,N_23734,N_24016);
nand U26960 (N_26960,N_20351,N_22756);
nor U26961 (N_26961,N_20549,N_24077);
nand U26962 (N_26962,N_23939,N_23332);
xnor U26963 (N_26963,N_20588,N_23943);
and U26964 (N_26964,N_23956,N_24585);
or U26965 (N_26965,N_22053,N_23660);
or U26966 (N_26966,N_21088,N_22925);
xnor U26967 (N_26967,N_20078,N_24865);
nand U26968 (N_26968,N_23572,N_20934);
nand U26969 (N_26969,N_24240,N_22054);
nand U26970 (N_26970,N_24112,N_20211);
and U26971 (N_26971,N_20736,N_24114);
or U26972 (N_26972,N_21907,N_23885);
xor U26973 (N_26973,N_22083,N_22294);
and U26974 (N_26974,N_21708,N_22612);
nor U26975 (N_26975,N_24432,N_20586);
nand U26976 (N_26976,N_22640,N_22307);
nor U26977 (N_26977,N_20036,N_21996);
xor U26978 (N_26978,N_22822,N_21738);
nand U26979 (N_26979,N_24956,N_24395);
nand U26980 (N_26980,N_21974,N_20134);
nand U26981 (N_26981,N_23752,N_20896);
nor U26982 (N_26982,N_22393,N_23624);
nand U26983 (N_26983,N_24485,N_21004);
nor U26984 (N_26984,N_20636,N_24410);
xnor U26985 (N_26985,N_23730,N_22147);
nor U26986 (N_26986,N_23544,N_23838);
xor U26987 (N_26987,N_23199,N_24767);
or U26988 (N_26988,N_21470,N_22275);
nor U26989 (N_26989,N_20899,N_24089);
xnor U26990 (N_26990,N_21795,N_22035);
or U26991 (N_26991,N_21168,N_24766);
or U26992 (N_26992,N_21443,N_21137);
and U26993 (N_26993,N_22020,N_21218);
nand U26994 (N_26994,N_22990,N_23412);
xor U26995 (N_26995,N_23619,N_21834);
nand U26996 (N_26996,N_20493,N_23880);
nor U26997 (N_26997,N_21952,N_24489);
and U26998 (N_26998,N_22997,N_24710);
and U26999 (N_26999,N_23193,N_24941);
nor U27000 (N_27000,N_23450,N_21891);
nor U27001 (N_27001,N_20027,N_24539);
or U27002 (N_27002,N_21954,N_20171);
or U27003 (N_27003,N_24062,N_21595);
and U27004 (N_27004,N_24596,N_20018);
nand U27005 (N_27005,N_20582,N_23646);
nor U27006 (N_27006,N_22279,N_23385);
and U27007 (N_27007,N_23742,N_23692);
and U27008 (N_27008,N_21924,N_22900);
or U27009 (N_27009,N_22457,N_21283);
nand U27010 (N_27010,N_24182,N_23554);
nor U27011 (N_27011,N_24253,N_23122);
xor U27012 (N_27012,N_20758,N_24053);
nand U27013 (N_27013,N_21414,N_23603);
and U27014 (N_27014,N_20601,N_20012);
nor U27015 (N_27015,N_22086,N_20430);
and U27016 (N_27016,N_22230,N_20505);
nor U27017 (N_27017,N_22673,N_21310);
and U27018 (N_27018,N_23430,N_22031);
nor U27019 (N_27019,N_23109,N_21625);
nor U27020 (N_27020,N_23254,N_24158);
nand U27021 (N_27021,N_24299,N_23303);
nor U27022 (N_27022,N_23760,N_21077);
nand U27023 (N_27023,N_21031,N_23905);
nand U27024 (N_27024,N_23517,N_23225);
and U27025 (N_27025,N_24917,N_24201);
nand U27026 (N_27026,N_21678,N_23147);
or U27027 (N_27027,N_20886,N_24466);
or U27028 (N_27028,N_23925,N_23720);
or U27029 (N_27029,N_23826,N_22170);
nor U27030 (N_27030,N_22815,N_23951);
nand U27031 (N_27031,N_21145,N_22889);
nor U27032 (N_27032,N_23346,N_21036);
nand U27033 (N_27033,N_20329,N_24829);
or U27034 (N_27034,N_22002,N_22099);
nand U27035 (N_27035,N_23808,N_22681);
nor U27036 (N_27036,N_21293,N_20140);
and U27037 (N_27037,N_22448,N_24221);
nand U27038 (N_27038,N_20194,N_22873);
or U27039 (N_27039,N_20000,N_22082);
nor U27040 (N_27040,N_23449,N_22629);
and U27041 (N_27041,N_20735,N_22027);
nor U27042 (N_27042,N_21676,N_22497);
nand U27043 (N_27043,N_21654,N_21655);
nand U27044 (N_27044,N_23621,N_24907);
nand U27045 (N_27045,N_24285,N_23788);
and U27046 (N_27046,N_21184,N_24405);
and U27047 (N_27047,N_24352,N_23446);
nor U27048 (N_27048,N_21459,N_23557);
and U27049 (N_27049,N_22472,N_22210);
nor U27050 (N_27050,N_23540,N_23710);
and U27051 (N_27051,N_24199,N_20954);
nor U27052 (N_27052,N_20434,N_24133);
and U27053 (N_27053,N_21691,N_20905);
xor U27054 (N_27054,N_24820,N_24219);
nor U27055 (N_27055,N_23194,N_22659);
nor U27056 (N_27056,N_23492,N_21703);
nor U27057 (N_27057,N_23535,N_24778);
xnor U27058 (N_27058,N_23837,N_20304);
nand U27059 (N_27059,N_20362,N_22751);
nand U27060 (N_27060,N_23236,N_23095);
nor U27061 (N_27061,N_23111,N_24514);
nor U27062 (N_27062,N_22863,N_22006);
and U27063 (N_27063,N_23393,N_23526);
xor U27064 (N_27064,N_23979,N_24626);
or U27065 (N_27065,N_24786,N_22718);
nor U27066 (N_27066,N_20608,N_22146);
nor U27067 (N_27067,N_20089,N_22022);
or U27068 (N_27068,N_21523,N_21956);
xor U27069 (N_27069,N_22455,N_24796);
and U27070 (N_27070,N_21600,N_20597);
nor U27071 (N_27071,N_22632,N_23651);
and U27072 (N_27072,N_23562,N_23844);
nor U27073 (N_27073,N_23103,N_24476);
or U27074 (N_27074,N_21849,N_23748);
nand U27075 (N_27075,N_20567,N_22768);
or U27076 (N_27076,N_24881,N_23507);
xnor U27077 (N_27077,N_21970,N_23369);
or U27078 (N_27078,N_23259,N_22373);
nor U27079 (N_27079,N_23950,N_20403);
nor U27080 (N_27080,N_23828,N_21388);
and U27081 (N_27081,N_21132,N_24984);
xnor U27082 (N_27082,N_24874,N_21157);
or U27083 (N_27083,N_20773,N_21736);
nor U27084 (N_27084,N_23329,N_22347);
and U27085 (N_27085,N_24546,N_20525);
and U27086 (N_27086,N_21326,N_24296);
or U27087 (N_27087,N_23559,N_24808);
nand U27088 (N_27088,N_23513,N_24433);
and U27089 (N_27089,N_20818,N_22928);
nand U27090 (N_27090,N_24374,N_23074);
nand U27091 (N_27091,N_20268,N_23571);
xor U27092 (N_27092,N_23321,N_24974);
nand U27093 (N_27093,N_22174,N_20285);
xnor U27094 (N_27094,N_22433,N_24495);
xnor U27095 (N_27095,N_23794,N_21205);
and U27096 (N_27096,N_24245,N_21030);
nor U27097 (N_27097,N_22975,N_20701);
xnor U27098 (N_27098,N_20172,N_24178);
and U27099 (N_27099,N_22261,N_20065);
or U27100 (N_27100,N_20785,N_21853);
nor U27101 (N_27101,N_22306,N_21718);
or U27102 (N_27102,N_23032,N_20312);
or U27103 (N_27103,N_23047,N_20289);
or U27104 (N_27104,N_21020,N_22332);
nand U27105 (N_27105,N_20197,N_20045);
and U27106 (N_27106,N_20452,N_22069);
or U27107 (N_27107,N_24683,N_24049);
nor U27108 (N_27108,N_23853,N_21975);
or U27109 (N_27109,N_23237,N_24225);
nand U27110 (N_27110,N_21775,N_21869);
nand U27111 (N_27111,N_22363,N_20919);
or U27112 (N_27112,N_23099,N_20730);
or U27113 (N_27113,N_20596,N_22184);
or U27114 (N_27114,N_21918,N_21962);
or U27115 (N_27115,N_23725,N_23616);
nor U27116 (N_27116,N_23291,N_21085);
and U27117 (N_27117,N_22658,N_24017);
xor U27118 (N_27118,N_24326,N_21170);
nand U27119 (N_27119,N_22870,N_20061);
and U27120 (N_27120,N_23000,N_24288);
xor U27121 (N_27121,N_22222,N_21978);
or U27122 (N_27122,N_20051,N_21721);
and U27123 (N_27123,N_23414,N_21946);
nand U27124 (N_27124,N_23825,N_22406);
and U27125 (N_27125,N_22766,N_24672);
or U27126 (N_27126,N_23587,N_22132);
nand U27127 (N_27127,N_22273,N_24362);
or U27128 (N_27128,N_21405,N_23927);
and U27129 (N_27129,N_21187,N_23017);
nor U27130 (N_27130,N_20219,N_22688);
or U27131 (N_27131,N_21622,N_23389);
nor U27132 (N_27132,N_23500,N_20637);
nor U27133 (N_27133,N_23410,N_20906);
and U27134 (N_27134,N_23154,N_22338);
or U27135 (N_27135,N_24329,N_20506);
and U27136 (N_27136,N_24099,N_23863);
or U27137 (N_27137,N_24530,N_23548);
nand U27138 (N_27138,N_20218,N_23401);
nor U27139 (N_27139,N_20081,N_23684);
nor U27140 (N_27140,N_23976,N_21379);
nor U27141 (N_27141,N_21532,N_20170);
or U27142 (N_27142,N_20694,N_20666);
and U27143 (N_27143,N_22931,N_23504);
nor U27144 (N_27144,N_21784,N_24622);
and U27145 (N_27145,N_22111,N_20712);
nand U27146 (N_27146,N_21547,N_22726);
or U27147 (N_27147,N_22845,N_21403);
nor U27148 (N_27148,N_22109,N_20168);
or U27149 (N_27149,N_23551,N_23712);
nand U27150 (N_27150,N_24494,N_24762);
xor U27151 (N_27151,N_24525,N_23879);
xor U27152 (N_27152,N_23756,N_24231);
nor U27153 (N_27153,N_22936,N_24412);
xor U27154 (N_27154,N_20883,N_20842);
nor U27155 (N_27155,N_24570,N_22689);
nand U27156 (N_27156,N_21377,N_22367);
nand U27157 (N_27157,N_24962,N_21969);
nor U27158 (N_27158,N_23803,N_24244);
or U27159 (N_27159,N_22258,N_20510);
xnor U27160 (N_27160,N_20923,N_20406);
or U27161 (N_27161,N_24137,N_20872);
or U27162 (N_27162,N_22301,N_20343);
nand U27163 (N_27163,N_23886,N_20964);
or U27164 (N_27164,N_23859,N_21210);
nand U27165 (N_27165,N_23352,N_22669);
or U27166 (N_27166,N_22520,N_20837);
xor U27167 (N_27167,N_20188,N_20550);
or U27168 (N_27168,N_22875,N_20825);
nand U27169 (N_27169,N_21776,N_23384);
and U27170 (N_27170,N_21295,N_22807);
nor U27171 (N_27171,N_21717,N_23917);
xnor U27172 (N_27172,N_20086,N_20468);
xnor U27173 (N_27173,N_22587,N_21777);
or U27174 (N_27174,N_20793,N_21380);
and U27175 (N_27175,N_21123,N_21725);
and U27176 (N_27176,N_24821,N_20458);
nand U27177 (N_27177,N_21579,N_20465);
and U27178 (N_27178,N_20626,N_22737);
or U27179 (N_27179,N_21504,N_21709);
nand U27180 (N_27180,N_22661,N_24769);
and U27181 (N_27181,N_22740,N_21323);
and U27182 (N_27182,N_24788,N_20629);
xor U27183 (N_27183,N_21874,N_24044);
and U27184 (N_27184,N_24372,N_21325);
nand U27185 (N_27185,N_21038,N_24132);
nor U27186 (N_27186,N_23709,N_24948);
or U27187 (N_27187,N_24770,N_24249);
or U27188 (N_27188,N_24024,N_20670);
nor U27189 (N_27189,N_21455,N_21003);
or U27190 (N_27190,N_24340,N_24559);
and U27191 (N_27191,N_23295,N_20267);
nor U27192 (N_27192,N_22594,N_21358);
or U27193 (N_27193,N_22252,N_22534);
or U27194 (N_27194,N_21674,N_24198);
or U27195 (N_27195,N_23298,N_23260);
xor U27196 (N_27196,N_24591,N_20299);
or U27197 (N_27197,N_24011,N_23282);
and U27198 (N_27198,N_20104,N_24344);
nand U27199 (N_27199,N_22336,N_21303);
nand U27200 (N_27200,N_22019,N_21900);
or U27201 (N_27201,N_20225,N_23166);
and U27202 (N_27202,N_20684,N_22288);
xor U27203 (N_27203,N_20427,N_20867);
xnor U27204 (N_27204,N_20860,N_21931);
xor U27205 (N_27205,N_24761,N_21641);
nor U27206 (N_27206,N_24319,N_24465);
nand U27207 (N_27207,N_22981,N_22000);
nor U27208 (N_27208,N_20050,N_20709);
and U27209 (N_27209,N_24172,N_24146);
or U27210 (N_27210,N_21773,N_21068);
or U27211 (N_27211,N_23023,N_22745);
and U27212 (N_27212,N_23721,N_22162);
xor U27213 (N_27213,N_24314,N_23056);
and U27214 (N_27214,N_22844,N_24627);
xor U27215 (N_27215,N_20897,N_20077);
nand U27216 (N_27216,N_20373,N_23652);
nor U27217 (N_27217,N_24795,N_20744);
nand U27218 (N_27218,N_21670,N_24742);
or U27219 (N_27219,N_20179,N_20882);
nand U27220 (N_27220,N_21882,N_24161);
or U27221 (N_27221,N_24574,N_23403);
or U27222 (N_27222,N_22477,N_24686);
nand U27223 (N_27223,N_20887,N_22548);
or U27224 (N_27224,N_24110,N_21694);
and U27225 (N_27225,N_20977,N_21591);
or U27226 (N_27226,N_20256,N_24967);
nor U27227 (N_27227,N_21449,N_20302);
nor U27228 (N_27228,N_24236,N_20040);
nand U27229 (N_27229,N_21015,N_21075);
and U27230 (N_27230,N_20755,N_20652);
or U27231 (N_27231,N_23480,N_23519);
or U27232 (N_27232,N_23971,N_21668);
nand U27233 (N_27233,N_23539,N_20150);
nor U27234 (N_27234,N_22687,N_22397);
nand U27235 (N_27235,N_24057,N_24642);
xor U27236 (N_27236,N_22358,N_21509);
xor U27237 (N_27237,N_20337,N_20097);
nor U27238 (N_27238,N_21963,N_21287);
and U27239 (N_27239,N_22880,N_23114);
nor U27240 (N_27240,N_22159,N_20824);
and U27241 (N_27241,N_21558,N_21427);
and U27242 (N_27242,N_24505,N_23577);
or U27243 (N_27243,N_20135,N_21447);
nand U27244 (N_27244,N_24461,N_21733);
nor U27245 (N_27245,N_21319,N_24529);
or U27246 (N_27246,N_23569,N_20737);
and U27247 (N_27247,N_24455,N_22424);
or U27248 (N_27248,N_24738,N_24598);
or U27249 (N_27249,N_24939,N_22333);
xnor U27250 (N_27250,N_24224,N_21561);
and U27251 (N_27251,N_24707,N_24610);
or U27252 (N_27252,N_23006,N_20751);
nand U27253 (N_27253,N_20644,N_24488);
or U27254 (N_27254,N_22247,N_24039);
or U27255 (N_27255,N_23598,N_23362);
xor U27256 (N_27256,N_23790,N_20016);
nand U27257 (N_27257,N_24568,N_22445);
and U27258 (N_27258,N_21194,N_23301);
and U27259 (N_27259,N_20990,N_23860);
nand U27260 (N_27260,N_20542,N_21955);
and U27261 (N_27261,N_22739,N_21336);
nand U27262 (N_27262,N_20801,N_21608);
and U27263 (N_27263,N_24729,N_22704);
or U27264 (N_27264,N_21206,N_20060);
nor U27265 (N_27265,N_24037,N_21214);
or U27266 (N_27266,N_24835,N_21938);
or U27267 (N_27267,N_22569,N_23596);
nor U27268 (N_27268,N_21833,N_20028);
nor U27269 (N_27269,N_20583,N_21820);
nor U27270 (N_27270,N_21124,N_23284);
nand U27271 (N_27271,N_20463,N_24910);
or U27272 (N_27272,N_20174,N_24422);
nor U27273 (N_27273,N_21383,N_24719);
nor U27274 (N_27274,N_21093,N_24660);
nand U27275 (N_27275,N_24267,N_21419);
or U27276 (N_27276,N_23203,N_20183);
or U27277 (N_27277,N_20632,N_24924);
xor U27278 (N_27278,N_24215,N_21890);
nor U27279 (N_27279,N_22585,N_24327);
nand U27280 (N_27280,N_23378,N_24174);
nand U27281 (N_27281,N_23220,N_20275);
nand U27282 (N_27282,N_22514,N_22103);
and U27283 (N_27283,N_20331,N_21593);
and U27284 (N_27284,N_22129,N_20442);
nor U27285 (N_27285,N_21698,N_22913);
nand U27286 (N_27286,N_23382,N_20417);
and U27287 (N_27287,N_23471,N_20967);
xnor U27288 (N_27288,N_22524,N_22972);
or U27289 (N_27289,N_23780,N_23733);
or U27290 (N_27290,N_23364,N_23687);
nand U27291 (N_27291,N_21175,N_20873);
nand U27292 (N_27292,N_22859,N_21838);
and U27293 (N_27293,N_23873,N_23497);
or U27294 (N_27294,N_22970,N_22076);
or U27295 (N_27295,N_23258,N_20494);
and U27296 (N_27296,N_21245,N_23443);
and U27297 (N_27297,N_20481,N_20011);
nor U27298 (N_27298,N_20764,N_20864);
nor U27299 (N_27299,N_23913,N_23238);
or U27300 (N_27300,N_24091,N_23900);
nand U27301 (N_27301,N_21010,N_23286);
nand U27302 (N_27302,N_24509,N_21742);
nand U27303 (N_27303,N_21363,N_22882);
or U27304 (N_27304,N_20936,N_21630);
or U27305 (N_27305,N_23732,N_20690);
nor U27306 (N_27306,N_21990,N_20766);
or U27307 (N_27307,N_24977,N_24649);
or U27308 (N_27308,N_21950,N_24582);
xnor U27309 (N_27309,N_22930,N_23053);
nand U27310 (N_27310,N_23505,N_23620);
nor U27311 (N_27311,N_22508,N_23862);
or U27312 (N_27312,N_24390,N_24481);
nand U27313 (N_27313,N_23811,N_22345);
and U27314 (N_27314,N_20319,N_22719);
and U27315 (N_27315,N_24556,N_22194);
nor U27316 (N_27316,N_20239,N_21436);
nor U27317 (N_27317,N_20347,N_24232);
or U27318 (N_27318,N_24289,N_24098);
nor U27319 (N_27319,N_21397,N_23680);
nor U27320 (N_27320,N_22914,N_20945);
nand U27321 (N_27321,N_23161,N_21320);
nor U27322 (N_27322,N_23274,N_22620);
nor U27323 (N_27323,N_22163,N_24222);
nand U27324 (N_27324,N_24675,N_21306);
nand U27325 (N_27325,N_22310,N_24351);
nor U27326 (N_27326,N_23704,N_22817);
nor U27327 (N_27327,N_22607,N_22244);
xor U27328 (N_27328,N_24862,N_21540);
nand U27329 (N_27329,N_21401,N_20742);
or U27330 (N_27330,N_22649,N_23664);
nand U27331 (N_27331,N_24331,N_24460);
or U27332 (N_27332,N_23257,N_22284);
nand U27333 (N_27333,N_24468,N_21847);
nand U27334 (N_27334,N_20623,N_20182);
nand U27335 (N_27335,N_24180,N_21017);
or U27336 (N_27336,N_20407,N_22490);
xor U27337 (N_27337,N_24976,N_24026);
or U27338 (N_27338,N_24010,N_23139);
nor U27339 (N_27339,N_20829,N_20288);
and U27340 (N_27340,N_21299,N_23966);
or U27341 (N_27341,N_24435,N_20831);
nor U27342 (N_27342,N_21949,N_24629);
and U27343 (N_27343,N_23691,N_20845);
and U27344 (N_27344,N_23242,N_24043);
or U27345 (N_27345,N_23486,N_21885);
or U27346 (N_27346,N_24624,N_22898);
nor U27347 (N_27347,N_21255,N_20470);
nand U27348 (N_27348,N_23829,N_20647);
or U27349 (N_27349,N_23955,N_21404);
xor U27350 (N_27350,N_21478,N_23137);
or U27351 (N_27351,N_24457,N_21112);
and U27352 (N_27352,N_22214,N_20646);
nor U27353 (N_27353,N_24870,N_24754);
and U27354 (N_27354,N_24294,N_23601);
and U27355 (N_27355,N_21803,N_22871);
nor U27356 (N_27356,N_21022,N_20557);
nand U27357 (N_27357,N_21370,N_21699);
nand U27358 (N_27358,N_22611,N_24711);
and U27359 (N_27359,N_22528,N_23744);
nand U27360 (N_27360,N_22426,N_22327);
nand U27361 (N_27361,N_23302,N_22181);
xnor U27362 (N_27362,N_23907,N_20885);
and U27363 (N_27363,N_24281,N_24691);
nor U27364 (N_27364,N_21977,N_24160);
xor U27365 (N_27365,N_24474,N_23767);
nor U27366 (N_27366,N_20280,N_23205);
xor U27367 (N_27367,N_24300,N_23386);
or U27368 (N_27368,N_24251,N_22003);
nor U27369 (N_27369,N_20692,N_20429);
nor U27370 (N_27370,N_21964,N_22566);
nor U27371 (N_27371,N_21762,N_22677);
and U27372 (N_27372,N_21244,N_21135);
nand U27373 (N_27373,N_20917,N_24220);
nand U27374 (N_27374,N_24830,N_23796);
and U27375 (N_27375,N_23037,N_21268);
or U27376 (N_27376,N_24522,N_24238);
nor U27377 (N_27377,N_23672,N_22369);
xnor U27378 (N_27378,N_23149,N_23107);
nand U27379 (N_27379,N_22356,N_22712);
or U27380 (N_27380,N_21282,N_23743);
nor U27381 (N_27381,N_20484,N_24450);
or U27382 (N_27382,N_23181,N_21474);
or U27383 (N_27383,N_23719,N_23180);
and U27384 (N_27384,N_24937,N_20344);
nand U27385 (N_27385,N_24483,N_21850);
nand U27386 (N_27386,N_20815,N_22532);
nand U27387 (N_27387,N_24162,N_20293);
nand U27388 (N_27388,N_24355,N_21302);
nor U27389 (N_27389,N_24183,N_24601);
nand U27390 (N_27390,N_24131,N_24723);
and U27391 (N_27391,N_24608,N_23442);
nor U27392 (N_27392,N_24998,N_24650);
nor U27393 (N_27393,N_22359,N_24143);
nand U27394 (N_27394,N_22150,N_21920);
or U27395 (N_27395,N_20010,N_23051);
nand U27396 (N_27396,N_22776,N_21043);
xnor U27397 (N_27397,N_20726,N_20419);
nand U27398 (N_27398,N_20184,N_24553);
nand U27399 (N_27399,N_23452,N_22157);
xnor U27400 (N_27400,N_23982,N_21348);
and U27401 (N_27401,N_24442,N_20561);
nand U27402 (N_27402,N_24453,N_20039);
or U27403 (N_27403,N_20949,N_22287);
xor U27404 (N_27404,N_24996,N_22504);
and U27405 (N_27405,N_22577,N_24933);
or U27406 (N_27406,N_21012,N_23695);
xnor U27407 (N_27407,N_23320,N_24547);
nand U27408 (N_27408,N_23080,N_22775);
or U27409 (N_27409,N_23429,N_21428);
nand U27410 (N_27410,N_23868,N_23406);
nand U27411 (N_27411,N_20877,N_22747);
or U27412 (N_27412,N_21821,N_22654);
or U27413 (N_27413,N_24250,N_20092);
nand U27414 (N_27414,N_22124,N_24773);
nor U27415 (N_27415,N_23078,N_23349);
and U27416 (N_27416,N_24973,N_21550);
or U27417 (N_27417,N_21376,N_23116);
and U27418 (N_27418,N_20649,N_23754);
xnor U27419 (N_27419,N_20826,N_24619);
or U27420 (N_27420,N_23962,N_21864);
or U27421 (N_27421,N_24074,N_22867);
nand U27422 (N_27422,N_20471,N_20593);
nand U27423 (N_27423,N_20169,N_24258);
and U27424 (N_27424,N_23600,N_20697);
nand U27425 (N_27425,N_22119,N_21463);
nor U27426 (N_27426,N_24908,N_23012);
xnor U27427 (N_27427,N_20017,N_20904);
and U27428 (N_27428,N_20126,N_21236);
or U27429 (N_27429,N_20253,N_24066);
nand U27430 (N_27430,N_24792,N_24696);
or U27431 (N_27431,N_23915,N_24593);
or U27432 (N_27432,N_24644,N_22330);
nand U27433 (N_27433,N_23415,N_20461);
and U27434 (N_27434,N_20581,N_24423);
and U27435 (N_27435,N_20782,N_24544);
or U27436 (N_27436,N_22311,N_22525);
nand U27437 (N_27437,N_24757,N_20198);
nor U27438 (N_27438,N_23015,N_21448);
nand U27439 (N_27439,N_24315,N_23250);
or U27440 (N_27440,N_20341,N_24506);
and U27441 (N_27441,N_24863,N_20366);
nand U27442 (N_27442,N_23878,N_24436);
xor U27443 (N_27443,N_22540,N_22883);
and U27444 (N_27444,N_21726,N_22102);
xor U27445 (N_27445,N_21180,N_23834);
nand U27446 (N_27446,N_22323,N_22733);
or U27447 (N_27447,N_23049,N_22826);
or U27448 (N_27448,N_20073,N_20133);
nor U27449 (N_27449,N_21045,N_21233);
and U27450 (N_27450,N_23031,N_20274);
xor U27451 (N_27451,N_20191,N_23992);
nand U27452 (N_27452,N_21153,N_20354);
nand U27453 (N_27453,N_21224,N_21221);
xnor U27454 (N_27454,N_20108,N_24690);
or U27455 (N_27455,N_24969,N_24287);
xor U27456 (N_27456,N_24430,N_23602);
nor U27457 (N_27457,N_24471,N_24897);
and U27458 (N_27458,N_23381,N_20124);
nor U27459 (N_27459,N_23700,N_20091);
nor U27460 (N_27460,N_22365,N_20305);
nor U27461 (N_27461,N_21013,N_23647);
nor U27462 (N_27462,N_22203,N_22924);
nand U27463 (N_27463,N_23872,N_21280);
or U27464 (N_27464,N_21518,N_22743);
nor U27465 (N_27465,N_23066,N_23368);
nand U27466 (N_27466,N_21251,N_22195);
nand U27467 (N_27467,N_20203,N_24177);
nand U27468 (N_27468,N_24388,N_22175);
nand U27469 (N_27469,N_20817,N_22390);
nand U27470 (N_27470,N_24491,N_24129);
nand U27471 (N_27471,N_21855,N_21423);
or U27472 (N_27472,N_24261,N_23558);
nor U27473 (N_27473,N_23851,N_24721);
nand U27474 (N_27474,N_24560,N_24406);
and U27475 (N_27475,N_20180,N_22788);
and U27476 (N_27476,N_21191,N_21374);
nor U27477 (N_27477,N_20099,N_23751);
or U27478 (N_27478,N_23268,N_21724);
and U27479 (N_27479,N_24768,N_22441);
xnor U27480 (N_27480,N_22535,N_21787);
or U27481 (N_27481,N_20844,N_21544);
nor U27482 (N_27482,N_23606,N_24508);
nand U27483 (N_27483,N_22694,N_23835);
and U27484 (N_27484,N_20562,N_24648);
nand U27485 (N_27485,N_20658,N_24647);
or U27486 (N_27486,N_20607,N_24078);
nor U27487 (N_27487,N_24880,N_20130);
or U27488 (N_27488,N_24804,N_23536);
xor U27489 (N_27489,N_22074,N_24981);
and U27490 (N_27490,N_21461,N_24892);
nand U27491 (N_27491,N_20308,N_20913);
nor U27492 (N_27492,N_23908,N_20314);
xor U27493 (N_27493,N_20661,N_24075);
or U27494 (N_27494,N_22702,N_20763);
or U27495 (N_27495,N_22176,N_20789);
or U27496 (N_27496,N_23092,N_21917);
and U27497 (N_27497,N_20832,N_24408);
nand U27498 (N_27498,N_20386,N_23072);
and U27499 (N_27499,N_24811,N_21441);
and U27500 (N_27500,N_20573,N_20363);
xor U27501 (N_27501,N_23099,N_21535);
or U27502 (N_27502,N_24119,N_24055);
or U27503 (N_27503,N_21269,N_23689);
nor U27504 (N_27504,N_24145,N_22938);
and U27505 (N_27505,N_24434,N_21695);
nand U27506 (N_27506,N_20345,N_21401);
xor U27507 (N_27507,N_22972,N_22553);
nand U27508 (N_27508,N_21500,N_21059);
or U27509 (N_27509,N_23972,N_23043);
nor U27510 (N_27510,N_20838,N_22312);
and U27511 (N_27511,N_23369,N_24338);
or U27512 (N_27512,N_20525,N_20315);
nand U27513 (N_27513,N_24652,N_22531);
nor U27514 (N_27514,N_22141,N_20912);
or U27515 (N_27515,N_20671,N_24326);
nor U27516 (N_27516,N_20358,N_24920);
nand U27517 (N_27517,N_21941,N_24196);
and U27518 (N_27518,N_24255,N_20969);
and U27519 (N_27519,N_21717,N_20279);
or U27520 (N_27520,N_20627,N_22584);
nor U27521 (N_27521,N_21828,N_21014);
or U27522 (N_27522,N_22271,N_22842);
nor U27523 (N_27523,N_22568,N_24576);
xnor U27524 (N_27524,N_20119,N_21524);
nor U27525 (N_27525,N_22623,N_24314);
xnor U27526 (N_27526,N_20525,N_24121);
or U27527 (N_27527,N_21298,N_24643);
xor U27528 (N_27528,N_22800,N_23164);
or U27529 (N_27529,N_20204,N_23555);
and U27530 (N_27530,N_22810,N_21240);
xnor U27531 (N_27531,N_24339,N_23405);
xor U27532 (N_27532,N_20410,N_21671);
or U27533 (N_27533,N_20094,N_22085);
nor U27534 (N_27534,N_24728,N_24912);
nand U27535 (N_27535,N_23979,N_21038);
and U27536 (N_27536,N_24674,N_21423);
or U27537 (N_27537,N_20546,N_20267);
nor U27538 (N_27538,N_24917,N_23872);
nand U27539 (N_27539,N_21767,N_24050);
xor U27540 (N_27540,N_22495,N_22346);
nand U27541 (N_27541,N_20746,N_24961);
nor U27542 (N_27542,N_24715,N_23516);
nand U27543 (N_27543,N_21417,N_21851);
nor U27544 (N_27544,N_21787,N_22726);
nand U27545 (N_27545,N_20828,N_20927);
and U27546 (N_27546,N_21324,N_24989);
nand U27547 (N_27547,N_23632,N_23688);
nand U27548 (N_27548,N_20117,N_21200);
nor U27549 (N_27549,N_20313,N_22623);
nor U27550 (N_27550,N_24907,N_24305);
nor U27551 (N_27551,N_24558,N_24870);
nor U27552 (N_27552,N_24925,N_23064);
xor U27553 (N_27553,N_21211,N_23734);
nand U27554 (N_27554,N_24630,N_23220);
and U27555 (N_27555,N_21344,N_24834);
and U27556 (N_27556,N_22231,N_21548);
nor U27557 (N_27557,N_20445,N_21399);
nor U27558 (N_27558,N_24195,N_20956);
nor U27559 (N_27559,N_22256,N_23848);
or U27560 (N_27560,N_20197,N_22045);
xnor U27561 (N_27561,N_21818,N_20513);
nor U27562 (N_27562,N_20620,N_23604);
nand U27563 (N_27563,N_23506,N_21584);
and U27564 (N_27564,N_21001,N_22418);
and U27565 (N_27565,N_23736,N_20473);
nor U27566 (N_27566,N_23701,N_20468);
nor U27567 (N_27567,N_23118,N_23525);
nand U27568 (N_27568,N_24486,N_24244);
or U27569 (N_27569,N_22801,N_24401);
nor U27570 (N_27570,N_21554,N_23181);
nor U27571 (N_27571,N_23200,N_23012);
and U27572 (N_27572,N_21207,N_24499);
xnor U27573 (N_27573,N_24552,N_22396);
or U27574 (N_27574,N_24311,N_22359);
or U27575 (N_27575,N_23484,N_20277);
nor U27576 (N_27576,N_20643,N_21626);
nand U27577 (N_27577,N_24012,N_23329);
and U27578 (N_27578,N_22982,N_21092);
or U27579 (N_27579,N_23953,N_20984);
nand U27580 (N_27580,N_24394,N_21587);
nor U27581 (N_27581,N_23622,N_22887);
and U27582 (N_27582,N_20519,N_20474);
or U27583 (N_27583,N_21711,N_23562);
nor U27584 (N_27584,N_20221,N_20835);
nor U27585 (N_27585,N_20941,N_22842);
xnor U27586 (N_27586,N_23457,N_24411);
nor U27587 (N_27587,N_24109,N_21194);
nor U27588 (N_27588,N_23930,N_23562);
nor U27589 (N_27589,N_22521,N_23951);
nor U27590 (N_27590,N_22056,N_22747);
or U27591 (N_27591,N_20652,N_23480);
or U27592 (N_27592,N_23816,N_21357);
and U27593 (N_27593,N_22140,N_24141);
xor U27594 (N_27594,N_22706,N_24434);
nor U27595 (N_27595,N_22200,N_23129);
nand U27596 (N_27596,N_22352,N_20034);
nand U27597 (N_27597,N_24557,N_24806);
or U27598 (N_27598,N_24642,N_24221);
and U27599 (N_27599,N_23021,N_21449);
or U27600 (N_27600,N_23466,N_20022);
or U27601 (N_27601,N_21283,N_20114);
nand U27602 (N_27602,N_20409,N_22207);
xnor U27603 (N_27603,N_22481,N_24149);
or U27604 (N_27604,N_20702,N_22803);
and U27605 (N_27605,N_24211,N_24972);
and U27606 (N_27606,N_21549,N_21544);
or U27607 (N_27607,N_24202,N_20008);
xnor U27608 (N_27608,N_22635,N_20571);
and U27609 (N_27609,N_24825,N_24329);
nor U27610 (N_27610,N_24941,N_24244);
and U27611 (N_27611,N_23633,N_24647);
nand U27612 (N_27612,N_23898,N_20756);
and U27613 (N_27613,N_23616,N_21057);
nor U27614 (N_27614,N_20570,N_20015);
or U27615 (N_27615,N_22444,N_20688);
or U27616 (N_27616,N_24640,N_23997);
nand U27617 (N_27617,N_20946,N_24378);
xor U27618 (N_27618,N_24690,N_24113);
nand U27619 (N_27619,N_20597,N_23912);
or U27620 (N_27620,N_23719,N_21246);
or U27621 (N_27621,N_24559,N_21506);
or U27622 (N_27622,N_20648,N_21228);
nand U27623 (N_27623,N_22322,N_20244);
nor U27624 (N_27624,N_24512,N_22574);
nor U27625 (N_27625,N_22198,N_24710);
or U27626 (N_27626,N_21160,N_22928);
nor U27627 (N_27627,N_23084,N_21159);
xnor U27628 (N_27628,N_24241,N_20420);
xor U27629 (N_27629,N_23073,N_20569);
xnor U27630 (N_27630,N_22095,N_21010);
nor U27631 (N_27631,N_24043,N_21229);
or U27632 (N_27632,N_24691,N_20152);
and U27633 (N_27633,N_24135,N_24513);
nand U27634 (N_27634,N_24101,N_22714);
nor U27635 (N_27635,N_24135,N_22168);
or U27636 (N_27636,N_24049,N_24596);
nand U27637 (N_27637,N_22322,N_21469);
or U27638 (N_27638,N_24648,N_24589);
and U27639 (N_27639,N_21254,N_20510);
and U27640 (N_27640,N_22452,N_23144);
nand U27641 (N_27641,N_24695,N_20914);
and U27642 (N_27642,N_23349,N_21075);
and U27643 (N_27643,N_21029,N_23497);
and U27644 (N_27644,N_23749,N_21437);
nand U27645 (N_27645,N_20538,N_23086);
nand U27646 (N_27646,N_21356,N_21060);
nand U27647 (N_27647,N_20544,N_21160);
or U27648 (N_27648,N_20914,N_23928);
nor U27649 (N_27649,N_22235,N_24132);
or U27650 (N_27650,N_22896,N_21794);
nor U27651 (N_27651,N_20609,N_23755);
xnor U27652 (N_27652,N_20622,N_21598);
nand U27653 (N_27653,N_24989,N_23632);
or U27654 (N_27654,N_20501,N_22178);
nand U27655 (N_27655,N_20435,N_24933);
nor U27656 (N_27656,N_23798,N_24859);
nor U27657 (N_27657,N_22800,N_21763);
or U27658 (N_27658,N_22297,N_24188);
and U27659 (N_27659,N_24463,N_23223);
and U27660 (N_27660,N_20556,N_23443);
or U27661 (N_27661,N_20992,N_20673);
nand U27662 (N_27662,N_22796,N_22574);
and U27663 (N_27663,N_23409,N_23002);
nor U27664 (N_27664,N_24817,N_22788);
nand U27665 (N_27665,N_23436,N_24082);
xnor U27666 (N_27666,N_22563,N_21132);
nand U27667 (N_27667,N_20256,N_22629);
or U27668 (N_27668,N_24551,N_23131);
nor U27669 (N_27669,N_20430,N_21787);
or U27670 (N_27670,N_20926,N_22399);
nand U27671 (N_27671,N_21797,N_22725);
and U27672 (N_27672,N_23838,N_20665);
nor U27673 (N_27673,N_23222,N_24325);
nand U27674 (N_27674,N_21405,N_22291);
xor U27675 (N_27675,N_22671,N_20134);
nor U27676 (N_27676,N_21839,N_24910);
nor U27677 (N_27677,N_20381,N_23979);
and U27678 (N_27678,N_24601,N_22907);
nor U27679 (N_27679,N_21145,N_22062);
xor U27680 (N_27680,N_24836,N_22970);
xnor U27681 (N_27681,N_22144,N_21563);
nand U27682 (N_27682,N_23628,N_21948);
nand U27683 (N_27683,N_22923,N_21180);
xnor U27684 (N_27684,N_22530,N_22154);
nor U27685 (N_27685,N_22527,N_23007);
or U27686 (N_27686,N_22583,N_21892);
nand U27687 (N_27687,N_23888,N_24555);
or U27688 (N_27688,N_24321,N_21324);
nor U27689 (N_27689,N_22087,N_22975);
nand U27690 (N_27690,N_22095,N_21580);
or U27691 (N_27691,N_22673,N_23935);
or U27692 (N_27692,N_21520,N_24036);
nand U27693 (N_27693,N_24746,N_24166);
or U27694 (N_27694,N_20171,N_23465);
and U27695 (N_27695,N_24517,N_20164);
nand U27696 (N_27696,N_20411,N_24227);
nor U27697 (N_27697,N_20178,N_21887);
nand U27698 (N_27698,N_24609,N_24755);
and U27699 (N_27699,N_23480,N_24639);
nand U27700 (N_27700,N_24253,N_21309);
nand U27701 (N_27701,N_22626,N_22628);
nor U27702 (N_27702,N_23129,N_23090);
and U27703 (N_27703,N_22499,N_20619);
xnor U27704 (N_27704,N_24400,N_23099);
nor U27705 (N_27705,N_24081,N_20188);
nor U27706 (N_27706,N_20174,N_20639);
nor U27707 (N_27707,N_24108,N_23863);
nor U27708 (N_27708,N_21491,N_22022);
and U27709 (N_27709,N_21149,N_21432);
or U27710 (N_27710,N_23008,N_21697);
nor U27711 (N_27711,N_21429,N_21087);
nor U27712 (N_27712,N_22472,N_23370);
nor U27713 (N_27713,N_20460,N_22434);
nor U27714 (N_27714,N_23281,N_22870);
nor U27715 (N_27715,N_21085,N_24140);
and U27716 (N_27716,N_20198,N_24557);
and U27717 (N_27717,N_24642,N_20925);
nor U27718 (N_27718,N_20246,N_23944);
nor U27719 (N_27719,N_24025,N_22906);
nor U27720 (N_27720,N_22122,N_21589);
nand U27721 (N_27721,N_22021,N_23606);
nand U27722 (N_27722,N_20620,N_20240);
and U27723 (N_27723,N_20501,N_22718);
or U27724 (N_27724,N_23420,N_23131);
xnor U27725 (N_27725,N_20190,N_21156);
nand U27726 (N_27726,N_22581,N_21450);
nand U27727 (N_27727,N_24505,N_22848);
nor U27728 (N_27728,N_22242,N_22919);
and U27729 (N_27729,N_22072,N_20470);
and U27730 (N_27730,N_21964,N_24533);
and U27731 (N_27731,N_20627,N_21430);
nand U27732 (N_27732,N_23716,N_23723);
nor U27733 (N_27733,N_20406,N_22092);
nand U27734 (N_27734,N_21510,N_22451);
or U27735 (N_27735,N_23595,N_22040);
or U27736 (N_27736,N_20650,N_20472);
and U27737 (N_27737,N_20909,N_23075);
and U27738 (N_27738,N_21908,N_24021);
xnor U27739 (N_27739,N_22311,N_24930);
nand U27740 (N_27740,N_23705,N_23123);
or U27741 (N_27741,N_23944,N_23333);
nor U27742 (N_27742,N_23661,N_24504);
xnor U27743 (N_27743,N_23885,N_24579);
nor U27744 (N_27744,N_20683,N_21018);
nand U27745 (N_27745,N_22579,N_23134);
or U27746 (N_27746,N_23001,N_24021);
xnor U27747 (N_27747,N_20413,N_20631);
and U27748 (N_27748,N_21011,N_20474);
nor U27749 (N_27749,N_24264,N_21498);
nand U27750 (N_27750,N_21679,N_22022);
or U27751 (N_27751,N_20294,N_20662);
nand U27752 (N_27752,N_20696,N_23468);
nand U27753 (N_27753,N_20181,N_23686);
nor U27754 (N_27754,N_23172,N_24860);
or U27755 (N_27755,N_22738,N_21287);
nor U27756 (N_27756,N_20754,N_23643);
or U27757 (N_27757,N_23416,N_23526);
and U27758 (N_27758,N_24001,N_24126);
nand U27759 (N_27759,N_23038,N_21101);
nand U27760 (N_27760,N_20262,N_20633);
nand U27761 (N_27761,N_20258,N_22612);
nand U27762 (N_27762,N_21242,N_24154);
and U27763 (N_27763,N_23060,N_23221);
or U27764 (N_27764,N_20101,N_20980);
xor U27765 (N_27765,N_21778,N_21009);
or U27766 (N_27766,N_22615,N_21867);
or U27767 (N_27767,N_20568,N_24438);
nand U27768 (N_27768,N_20947,N_21378);
and U27769 (N_27769,N_21914,N_23428);
nand U27770 (N_27770,N_24059,N_20238);
nand U27771 (N_27771,N_24993,N_21333);
or U27772 (N_27772,N_22312,N_23696);
xor U27773 (N_27773,N_22262,N_20816);
or U27774 (N_27774,N_24942,N_23696);
and U27775 (N_27775,N_22400,N_23295);
or U27776 (N_27776,N_20355,N_23435);
or U27777 (N_27777,N_23057,N_21133);
or U27778 (N_27778,N_20819,N_20269);
xor U27779 (N_27779,N_23863,N_23758);
or U27780 (N_27780,N_20607,N_24896);
and U27781 (N_27781,N_21284,N_21706);
and U27782 (N_27782,N_22992,N_23211);
or U27783 (N_27783,N_22853,N_24281);
nor U27784 (N_27784,N_20320,N_23752);
or U27785 (N_27785,N_21375,N_24318);
nor U27786 (N_27786,N_22166,N_20662);
nor U27787 (N_27787,N_20892,N_24896);
nor U27788 (N_27788,N_20896,N_21434);
nor U27789 (N_27789,N_23952,N_23408);
xnor U27790 (N_27790,N_21301,N_20990);
or U27791 (N_27791,N_23330,N_21435);
nor U27792 (N_27792,N_22754,N_23317);
nand U27793 (N_27793,N_22998,N_23211);
and U27794 (N_27794,N_22931,N_24526);
nand U27795 (N_27795,N_22550,N_22819);
xor U27796 (N_27796,N_20566,N_21356);
and U27797 (N_27797,N_22722,N_21971);
and U27798 (N_27798,N_21385,N_23833);
nor U27799 (N_27799,N_20832,N_23679);
xnor U27800 (N_27800,N_21142,N_22913);
nor U27801 (N_27801,N_24493,N_20017);
and U27802 (N_27802,N_23083,N_21819);
nand U27803 (N_27803,N_20956,N_23099);
nand U27804 (N_27804,N_24486,N_21045);
or U27805 (N_27805,N_20996,N_21416);
nor U27806 (N_27806,N_24377,N_24804);
and U27807 (N_27807,N_24206,N_23097);
and U27808 (N_27808,N_21172,N_20441);
or U27809 (N_27809,N_20014,N_20762);
nor U27810 (N_27810,N_20829,N_24521);
nor U27811 (N_27811,N_21002,N_22123);
and U27812 (N_27812,N_22943,N_23706);
nand U27813 (N_27813,N_22783,N_20108);
nand U27814 (N_27814,N_20208,N_20164);
or U27815 (N_27815,N_22365,N_23452);
and U27816 (N_27816,N_21741,N_22488);
nand U27817 (N_27817,N_22312,N_20873);
and U27818 (N_27818,N_24290,N_22281);
or U27819 (N_27819,N_22591,N_24666);
or U27820 (N_27820,N_24069,N_23552);
nand U27821 (N_27821,N_23972,N_24491);
xor U27822 (N_27822,N_20921,N_24602);
and U27823 (N_27823,N_24291,N_24234);
or U27824 (N_27824,N_23636,N_20274);
nand U27825 (N_27825,N_24401,N_24992);
nor U27826 (N_27826,N_21824,N_24815);
nand U27827 (N_27827,N_21543,N_24026);
or U27828 (N_27828,N_21413,N_22155);
and U27829 (N_27829,N_23633,N_24408);
nand U27830 (N_27830,N_20227,N_20880);
nor U27831 (N_27831,N_21791,N_23482);
and U27832 (N_27832,N_22040,N_21572);
or U27833 (N_27833,N_22078,N_24879);
and U27834 (N_27834,N_20292,N_21571);
or U27835 (N_27835,N_22459,N_23521);
or U27836 (N_27836,N_20299,N_20806);
or U27837 (N_27837,N_21883,N_20151);
nor U27838 (N_27838,N_24162,N_20921);
nor U27839 (N_27839,N_23556,N_24949);
nand U27840 (N_27840,N_23777,N_23329);
xnor U27841 (N_27841,N_20853,N_23353);
or U27842 (N_27842,N_22502,N_21083);
nand U27843 (N_27843,N_22126,N_20989);
nor U27844 (N_27844,N_22149,N_21853);
or U27845 (N_27845,N_24703,N_20487);
or U27846 (N_27846,N_24638,N_23352);
nand U27847 (N_27847,N_23201,N_24771);
nand U27848 (N_27848,N_24772,N_22489);
nand U27849 (N_27849,N_23802,N_24467);
or U27850 (N_27850,N_21802,N_22793);
and U27851 (N_27851,N_21613,N_20377);
or U27852 (N_27852,N_20711,N_24941);
nor U27853 (N_27853,N_20874,N_24415);
nor U27854 (N_27854,N_20110,N_20060);
nand U27855 (N_27855,N_21836,N_23730);
and U27856 (N_27856,N_22530,N_22367);
nor U27857 (N_27857,N_21726,N_20379);
or U27858 (N_27858,N_23406,N_23023);
nor U27859 (N_27859,N_20894,N_20603);
or U27860 (N_27860,N_23886,N_24995);
or U27861 (N_27861,N_20816,N_21220);
nor U27862 (N_27862,N_24821,N_20400);
and U27863 (N_27863,N_24723,N_24048);
and U27864 (N_27864,N_22875,N_22063);
or U27865 (N_27865,N_20707,N_24382);
nor U27866 (N_27866,N_20767,N_23282);
nor U27867 (N_27867,N_24684,N_24167);
and U27868 (N_27868,N_23226,N_24225);
nand U27869 (N_27869,N_22256,N_20707);
nand U27870 (N_27870,N_20399,N_22515);
nor U27871 (N_27871,N_22656,N_22120);
xnor U27872 (N_27872,N_21223,N_21778);
nor U27873 (N_27873,N_24255,N_24369);
nand U27874 (N_27874,N_23653,N_20663);
or U27875 (N_27875,N_22492,N_20488);
or U27876 (N_27876,N_23377,N_23222);
nand U27877 (N_27877,N_22765,N_20105);
nor U27878 (N_27878,N_24338,N_22971);
nand U27879 (N_27879,N_21986,N_23859);
nor U27880 (N_27880,N_20684,N_22139);
nand U27881 (N_27881,N_21957,N_24617);
nand U27882 (N_27882,N_20831,N_20084);
or U27883 (N_27883,N_21204,N_24742);
or U27884 (N_27884,N_22301,N_23282);
nor U27885 (N_27885,N_24134,N_24480);
nand U27886 (N_27886,N_21602,N_21252);
or U27887 (N_27887,N_20301,N_21402);
nor U27888 (N_27888,N_23160,N_22117);
xor U27889 (N_27889,N_23873,N_24440);
and U27890 (N_27890,N_23019,N_21793);
or U27891 (N_27891,N_24134,N_21197);
xor U27892 (N_27892,N_23212,N_24757);
nand U27893 (N_27893,N_23908,N_22109);
xor U27894 (N_27894,N_23079,N_24163);
or U27895 (N_27895,N_23365,N_23777);
nand U27896 (N_27896,N_24176,N_20868);
and U27897 (N_27897,N_23130,N_24880);
nand U27898 (N_27898,N_24762,N_23659);
nand U27899 (N_27899,N_23188,N_20581);
and U27900 (N_27900,N_21199,N_20492);
nor U27901 (N_27901,N_22861,N_22471);
or U27902 (N_27902,N_21635,N_24245);
nor U27903 (N_27903,N_22418,N_20140);
or U27904 (N_27904,N_24071,N_21651);
nand U27905 (N_27905,N_24439,N_22480);
and U27906 (N_27906,N_21528,N_23398);
nor U27907 (N_27907,N_20133,N_23919);
nand U27908 (N_27908,N_23250,N_21656);
nor U27909 (N_27909,N_23195,N_21079);
nand U27910 (N_27910,N_23335,N_20389);
nor U27911 (N_27911,N_23127,N_23926);
xor U27912 (N_27912,N_21528,N_22858);
nor U27913 (N_27913,N_24510,N_23228);
nand U27914 (N_27914,N_20061,N_22858);
or U27915 (N_27915,N_23765,N_23031);
and U27916 (N_27916,N_21598,N_23958);
nor U27917 (N_27917,N_24647,N_20051);
xor U27918 (N_27918,N_23605,N_24299);
and U27919 (N_27919,N_22117,N_22579);
or U27920 (N_27920,N_22441,N_20228);
and U27921 (N_27921,N_23806,N_20672);
nand U27922 (N_27922,N_22381,N_20094);
nor U27923 (N_27923,N_23231,N_24677);
or U27924 (N_27924,N_23439,N_22699);
nor U27925 (N_27925,N_23052,N_23398);
nand U27926 (N_27926,N_23980,N_20327);
nand U27927 (N_27927,N_23321,N_22606);
and U27928 (N_27928,N_20498,N_20586);
xor U27929 (N_27929,N_24814,N_23136);
and U27930 (N_27930,N_23219,N_20659);
and U27931 (N_27931,N_22479,N_23790);
and U27932 (N_27932,N_20228,N_20745);
xnor U27933 (N_27933,N_23710,N_20093);
xnor U27934 (N_27934,N_22050,N_22267);
nor U27935 (N_27935,N_22380,N_21796);
xnor U27936 (N_27936,N_23620,N_20109);
and U27937 (N_27937,N_22329,N_20518);
nand U27938 (N_27938,N_24416,N_20515);
xnor U27939 (N_27939,N_22339,N_21628);
or U27940 (N_27940,N_24256,N_21393);
and U27941 (N_27941,N_22553,N_24742);
xor U27942 (N_27942,N_21310,N_21357);
or U27943 (N_27943,N_24771,N_24276);
nor U27944 (N_27944,N_24367,N_22384);
or U27945 (N_27945,N_21782,N_20051);
or U27946 (N_27946,N_23698,N_23655);
or U27947 (N_27947,N_23558,N_21914);
xor U27948 (N_27948,N_22045,N_24886);
and U27949 (N_27949,N_24809,N_22785);
nor U27950 (N_27950,N_24756,N_24623);
and U27951 (N_27951,N_20399,N_20484);
or U27952 (N_27952,N_22698,N_22623);
or U27953 (N_27953,N_22448,N_20704);
nand U27954 (N_27954,N_20609,N_22703);
or U27955 (N_27955,N_22038,N_24156);
nand U27956 (N_27956,N_20525,N_20153);
and U27957 (N_27957,N_20132,N_21745);
or U27958 (N_27958,N_23290,N_22258);
xnor U27959 (N_27959,N_23099,N_20193);
or U27960 (N_27960,N_21719,N_21073);
nand U27961 (N_27961,N_24895,N_21683);
or U27962 (N_27962,N_21277,N_22895);
xor U27963 (N_27963,N_22009,N_22521);
xnor U27964 (N_27964,N_20279,N_24718);
or U27965 (N_27965,N_24959,N_21631);
nor U27966 (N_27966,N_22991,N_24947);
nor U27967 (N_27967,N_22033,N_23368);
or U27968 (N_27968,N_21026,N_22245);
nor U27969 (N_27969,N_24923,N_21123);
nor U27970 (N_27970,N_24692,N_21152);
nor U27971 (N_27971,N_21964,N_22387);
and U27972 (N_27972,N_23512,N_20670);
nor U27973 (N_27973,N_21939,N_22062);
nor U27974 (N_27974,N_20137,N_23373);
or U27975 (N_27975,N_21003,N_20444);
nand U27976 (N_27976,N_22497,N_23191);
and U27977 (N_27977,N_21024,N_22228);
and U27978 (N_27978,N_24955,N_21906);
and U27979 (N_27979,N_23155,N_20031);
nand U27980 (N_27980,N_20428,N_22947);
nor U27981 (N_27981,N_23181,N_24539);
nand U27982 (N_27982,N_20853,N_24958);
xor U27983 (N_27983,N_23810,N_22653);
or U27984 (N_27984,N_22473,N_24284);
and U27985 (N_27985,N_21205,N_24843);
nand U27986 (N_27986,N_22544,N_21771);
and U27987 (N_27987,N_22970,N_21804);
nand U27988 (N_27988,N_24269,N_23499);
or U27989 (N_27989,N_24588,N_22633);
and U27990 (N_27990,N_22703,N_24394);
nand U27991 (N_27991,N_24905,N_20086);
or U27992 (N_27992,N_22685,N_23048);
nor U27993 (N_27993,N_22511,N_22139);
nor U27994 (N_27994,N_20343,N_23222);
xor U27995 (N_27995,N_22903,N_20085);
nor U27996 (N_27996,N_23732,N_20090);
or U27997 (N_27997,N_21416,N_21435);
nor U27998 (N_27998,N_22602,N_23311);
or U27999 (N_27999,N_24022,N_22915);
nand U28000 (N_28000,N_21196,N_23648);
nor U28001 (N_28001,N_20200,N_22351);
or U28002 (N_28002,N_24704,N_21785);
nor U28003 (N_28003,N_22240,N_23865);
nand U28004 (N_28004,N_22148,N_20818);
nor U28005 (N_28005,N_22003,N_22794);
nand U28006 (N_28006,N_21604,N_20440);
or U28007 (N_28007,N_21359,N_22451);
or U28008 (N_28008,N_24482,N_22393);
and U28009 (N_28009,N_24860,N_21065);
nand U28010 (N_28010,N_24026,N_21495);
and U28011 (N_28011,N_24855,N_21942);
and U28012 (N_28012,N_21039,N_23693);
nor U28013 (N_28013,N_24614,N_24022);
nand U28014 (N_28014,N_20502,N_21922);
and U28015 (N_28015,N_20428,N_23478);
xor U28016 (N_28016,N_21072,N_22954);
or U28017 (N_28017,N_23718,N_20904);
or U28018 (N_28018,N_23044,N_23102);
xnor U28019 (N_28019,N_24147,N_23441);
nor U28020 (N_28020,N_20387,N_22165);
or U28021 (N_28021,N_22868,N_23219);
nand U28022 (N_28022,N_22837,N_23797);
or U28023 (N_28023,N_22810,N_24512);
xor U28024 (N_28024,N_24514,N_24079);
and U28025 (N_28025,N_20954,N_24624);
and U28026 (N_28026,N_20766,N_23393);
or U28027 (N_28027,N_21659,N_22458);
nand U28028 (N_28028,N_20949,N_21248);
or U28029 (N_28029,N_22958,N_20308);
or U28030 (N_28030,N_24016,N_20403);
and U28031 (N_28031,N_22376,N_20690);
nor U28032 (N_28032,N_21597,N_20445);
or U28033 (N_28033,N_20356,N_22922);
and U28034 (N_28034,N_24657,N_21144);
and U28035 (N_28035,N_24841,N_20194);
nor U28036 (N_28036,N_24202,N_21886);
or U28037 (N_28037,N_20698,N_20719);
or U28038 (N_28038,N_20454,N_23295);
and U28039 (N_28039,N_21031,N_23023);
and U28040 (N_28040,N_20236,N_22603);
nand U28041 (N_28041,N_24519,N_21136);
nor U28042 (N_28042,N_21493,N_21782);
or U28043 (N_28043,N_22829,N_23767);
and U28044 (N_28044,N_22462,N_20772);
nand U28045 (N_28045,N_23929,N_24104);
or U28046 (N_28046,N_23785,N_22461);
or U28047 (N_28047,N_23766,N_22664);
nand U28048 (N_28048,N_24583,N_23344);
nor U28049 (N_28049,N_24200,N_21963);
or U28050 (N_28050,N_21950,N_20400);
nand U28051 (N_28051,N_22142,N_23084);
nand U28052 (N_28052,N_24969,N_24688);
nand U28053 (N_28053,N_22580,N_23078);
or U28054 (N_28054,N_20714,N_23421);
xor U28055 (N_28055,N_24953,N_22723);
or U28056 (N_28056,N_21132,N_20264);
nor U28057 (N_28057,N_23994,N_22990);
and U28058 (N_28058,N_20640,N_20096);
nor U28059 (N_28059,N_21634,N_21293);
nor U28060 (N_28060,N_22926,N_24754);
nand U28061 (N_28061,N_22448,N_23870);
nand U28062 (N_28062,N_21597,N_24993);
nor U28063 (N_28063,N_21709,N_22294);
or U28064 (N_28064,N_24130,N_23765);
nand U28065 (N_28065,N_21721,N_24825);
nand U28066 (N_28066,N_21524,N_20459);
nor U28067 (N_28067,N_23430,N_22249);
nand U28068 (N_28068,N_24657,N_23569);
nand U28069 (N_28069,N_20696,N_24660);
nor U28070 (N_28070,N_23258,N_20197);
or U28071 (N_28071,N_20965,N_21471);
and U28072 (N_28072,N_23229,N_22498);
nor U28073 (N_28073,N_24841,N_24190);
or U28074 (N_28074,N_22181,N_20370);
nor U28075 (N_28075,N_23250,N_21439);
or U28076 (N_28076,N_20699,N_21574);
and U28077 (N_28077,N_24165,N_24363);
nand U28078 (N_28078,N_21295,N_20919);
nor U28079 (N_28079,N_21298,N_20209);
nor U28080 (N_28080,N_24155,N_23448);
nor U28081 (N_28081,N_20833,N_22409);
nor U28082 (N_28082,N_21027,N_21952);
xnor U28083 (N_28083,N_23606,N_20062);
and U28084 (N_28084,N_23420,N_23116);
nor U28085 (N_28085,N_23722,N_24397);
nor U28086 (N_28086,N_21149,N_24336);
nor U28087 (N_28087,N_20721,N_23872);
xor U28088 (N_28088,N_23099,N_21368);
nand U28089 (N_28089,N_23778,N_20802);
nand U28090 (N_28090,N_21343,N_24372);
nand U28091 (N_28091,N_21334,N_21538);
nand U28092 (N_28092,N_24921,N_22940);
or U28093 (N_28093,N_23282,N_21391);
or U28094 (N_28094,N_20145,N_22619);
or U28095 (N_28095,N_24605,N_21135);
and U28096 (N_28096,N_22007,N_24026);
or U28097 (N_28097,N_21562,N_20124);
nor U28098 (N_28098,N_24929,N_24772);
nand U28099 (N_28099,N_22961,N_21822);
nor U28100 (N_28100,N_22153,N_23993);
or U28101 (N_28101,N_21869,N_24301);
nor U28102 (N_28102,N_24304,N_23464);
or U28103 (N_28103,N_24738,N_24501);
nand U28104 (N_28104,N_22733,N_24081);
or U28105 (N_28105,N_24687,N_21158);
or U28106 (N_28106,N_22608,N_24432);
or U28107 (N_28107,N_24368,N_23096);
nor U28108 (N_28108,N_21884,N_21441);
nor U28109 (N_28109,N_21133,N_20461);
nor U28110 (N_28110,N_21908,N_22951);
nor U28111 (N_28111,N_24969,N_22920);
and U28112 (N_28112,N_24368,N_23201);
nor U28113 (N_28113,N_22241,N_24211);
and U28114 (N_28114,N_22897,N_20825);
nor U28115 (N_28115,N_24146,N_22537);
and U28116 (N_28116,N_20472,N_22743);
nor U28117 (N_28117,N_20817,N_22704);
nand U28118 (N_28118,N_20351,N_21477);
and U28119 (N_28119,N_21978,N_24238);
nor U28120 (N_28120,N_20970,N_22262);
xor U28121 (N_28121,N_22985,N_20394);
nand U28122 (N_28122,N_20502,N_22261);
nand U28123 (N_28123,N_22308,N_22050);
and U28124 (N_28124,N_20688,N_24054);
xor U28125 (N_28125,N_24341,N_23616);
and U28126 (N_28126,N_22002,N_22961);
nand U28127 (N_28127,N_20896,N_24455);
or U28128 (N_28128,N_23990,N_24305);
or U28129 (N_28129,N_24986,N_23952);
xnor U28130 (N_28130,N_22725,N_22812);
nor U28131 (N_28131,N_20132,N_20040);
and U28132 (N_28132,N_24828,N_23926);
and U28133 (N_28133,N_24470,N_22925);
xnor U28134 (N_28134,N_21297,N_20279);
or U28135 (N_28135,N_23116,N_20415);
or U28136 (N_28136,N_21498,N_23717);
nor U28137 (N_28137,N_24021,N_22035);
or U28138 (N_28138,N_20044,N_22376);
nor U28139 (N_28139,N_21741,N_24301);
and U28140 (N_28140,N_21748,N_20642);
nand U28141 (N_28141,N_21245,N_22719);
nand U28142 (N_28142,N_20420,N_21261);
xor U28143 (N_28143,N_23775,N_22024);
nor U28144 (N_28144,N_24911,N_24721);
nand U28145 (N_28145,N_23729,N_20635);
nor U28146 (N_28146,N_24327,N_21056);
or U28147 (N_28147,N_20247,N_23397);
and U28148 (N_28148,N_21567,N_21406);
nor U28149 (N_28149,N_20445,N_20054);
and U28150 (N_28150,N_20783,N_22574);
or U28151 (N_28151,N_22891,N_20858);
nand U28152 (N_28152,N_22333,N_24293);
nand U28153 (N_28153,N_22656,N_24468);
and U28154 (N_28154,N_24334,N_20411);
nor U28155 (N_28155,N_22461,N_24932);
nand U28156 (N_28156,N_20951,N_22108);
nor U28157 (N_28157,N_21227,N_24640);
nand U28158 (N_28158,N_23628,N_23209);
or U28159 (N_28159,N_21610,N_24839);
nand U28160 (N_28160,N_23382,N_22565);
nand U28161 (N_28161,N_21387,N_22609);
and U28162 (N_28162,N_20655,N_20662);
and U28163 (N_28163,N_20313,N_21880);
and U28164 (N_28164,N_20010,N_23699);
or U28165 (N_28165,N_24456,N_24243);
nand U28166 (N_28166,N_22972,N_24032);
and U28167 (N_28167,N_21057,N_24872);
and U28168 (N_28168,N_24008,N_23705);
and U28169 (N_28169,N_21967,N_23263);
nand U28170 (N_28170,N_20888,N_24318);
or U28171 (N_28171,N_23474,N_23683);
xnor U28172 (N_28172,N_22750,N_21547);
nand U28173 (N_28173,N_23651,N_20860);
nor U28174 (N_28174,N_23611,N_21588);
nand U28175 (N_28175,N_22962,N_24770);
nor U28176 (N_28176,N_24916,N_21268);
nand U28177 (N_28177,N_24748,N_22665);
nor U28178 (N_28178,N_21155,N_20909);
or U28179 (N_28179,N_24548,N_20299);
nand U28180 (N_28180,N_20870,N_24700);
nand U28181 (N_28181,N_23587,N_20110);
nor U28182 (N_28182,N_23282,N_22842);
or U28183 (N_28183,N_23336,N_21389);
nor U28184 (N_28184,N_21489,N_22391);
nor U28185 (N_28185,N_21976,N_21250);
or U28186 (N_28186,N_21818,N_23700);
or U28187 (N_28187,N_20657,N_23595);
xor U28188 (N_28188,N_24933,N_24318);
nand U28189 (N_28189,N_23528,N_22341);
nor U28190 (N_28190,N_21723,N_21894);
nand U28191 (N_28191,N_24682,N_23612);
and U28192 (N_28192,N_24087,N_23426);
or U28193 (N_28193,N_23740,N_20308);
and U28194 (N_28194,N_24836,N_24793);
and U28195 (N_28195,N_20684,N_21825);
and U28196 (N_28196,N_20422,N_20906);
or U28197 (N_28197,N_22598,N_20257);
or U28198 (N_28198,N_21619,N_21301);
and U28199 (N_28199,N_21430,N_22645);
nand U28200 (N_28200,N_22785,N_23461);
nand U28201 (N_28201,N_21421,N_21191);
nand U28202 (N_28202,N_22796,N_24976);
and U28203 (N_28203,N_24228,N_24344);
and U28204 (N_28204,N_21382,N_22136);
or U28205 (N_28205,N_24014,N_23062);
or U28206 (N_28206,N_23786,N_22202);
xor U28207 (N_28207,N_24058,N_23123);
nand U28208 (N_28208,N_22303,N_23781);
nor U28209 (N_28209,N_24429,N_20897);
nand U28210 (N_28210,N_24240,N_20274);
and U28211 (N_28211,N_21217,N_24094);
xnor U28212 (N_28212,N_22461,N_24969);
and U28213 (N_28213,N_23707,N_20591);
and U28214 (N_28214,N_20490,N_20835);
and U28215 (N_28215,N_22765,N_20582);
or U28216 (N_28216,N_23084,N_24097);
and U28217 (N_28217,N_23254,N_22454);
nand U28218 (N_28218,N_20916,N_23538);
nand U28219 (N_28219,N_22109,N_23039);
or U28220 (N_28220,N_22403,N_22350);
nand U28221 (N_28221,N_23484,N_22580);
or U28222 (N_28222,N_22455,N_22273);
or U28223 (N_28223,N_20030,N_23923);
nand U28224 (N_28224,N_24242,N_21138);
or U28225 (N_28225,N_24132,N_24278);
nor U28226 (N_28226,N_22620,N_24495);
or U28227 (N_28227,N_24924,N_21349);
or U28228 (N_28228,N_23611,N_20247);
nand U28229 (N_28229,N_24757,N_22426);
nor U28230 (N_28230,N_22879,N_23836);
nor U28231 (N_28231,N_22200,N_22953);
nand U28232 (N_28232,N_24196,N_23543);
and U28233 (N_28233,N_22445,N_24255);
xnor U28234 (N_28234,N_23167,N_20077);
xnor U28235 (N_28235,N_21375,N_24501);
nor U28236 (N_28236,N_20799,N_24530);
or U28237 (N_28237,N_22884,N_22127);
xor U28238 (N_28238,N_22443,N_23011);
xor U28239 (N_28239,N_20744,N_24129);
nand U28240 (N_28240,N_22266,N_22660);
nor U28241 (N_28241,N_22986,N_22580);
nor U28242 (N_28242,N_22730,N_20220);
or U28243 (N_28243,N_22699,N_20296);
nor U28244 (N_28244,N_22139,N_21933);
or U28245 (N_28245,N_20161,N_24039);
or U28246 (N_28246,N_24645,N_20557);
xnor U28247 (N_28247,N_20200,N_21345);
nor U28248 (N_28248,N_23962,N_20689);
and U28249 (N_28249,N_24925,N_23456);
nor U28250 (N_28250,N_22569,N_20837);
and U28251 (N_28251,N_22391,N_21692);
nor U28252 (N_28252,N_24204,N_21718);
or U28253 (N_28253,N_23233,N_24794);
nor U28254 (N_28254,N_23187,N_22525);
and U28255 (N_28255,N_24769,N_23787);
xnor U28256 (N_28256,N_21336,N_24751);
or U28257 (N_28257,N_21747,N_22306);
nand U28258 (N_28258,N_21849,N_20976);
xnor U28259 (N_28259,N_22046,N_23141);
nor U28260 (N_28260,N_23516,N_21933);
xor U28261 (N_28261,N_24296,N_21429);
nor U28262 (N_28262,N_23570,N_23194);
nor U28263 (N_28263,N_20777,N_24542);
nor U28264 (N_28264,N_20304,N_22991);
nor U28265 (N_28265,N_24496,N_20002);
or U28266 (N_28266,N_23570,N_22464);
xnor U28267 (N_28267,N_22699,N_20919);
nor U28268 (N_28268,N_22203,N_24878);
and U28269 (N_28269,N_21524,N_24748);
nand U28270 (N_28270,N_23989,N_21412);
nand U28271 (N_28271,N_21195,N_24273);
nor U28272 (N_28272,N_20669,N_21338);
and U28273 (N_28273,N_21142,N_21941);
and U28274 (N_28274,N_22885,N_20382);
nor U28275 (N_28275,N_24650,N_23288);
nor U28276 (N_28276,N_20159,N_22523);
xnor U28277 (N_28277,N_21854,N_22221);
nor U28278 (N_28278,N_20817,N_20118);
nor U28279 (N_28279,N_23542,N_21611);
nor U28280 (N_28280,N_22771,N_23435);
and U28281 (N_28281,N_21409,N_23684);
nor U28282 (N_28282,N_24571,N_20448);
and U28283 (N_28283,N_23676,N_23694);
nand U28284 (N_28284,N_23282,N_21327);
nand U28285 (N_28285,N_23982,N_20095);
nand U28286 (N_28286,N_24036,N_22376);
and U28287 (N_28287,N_21316,N_22165);
xnor U28288 (N_28288,N_23182,N_24515);
nand U28289 (N_28289,N_22737,N_20179);
xor U28290 (N_28290,N_20730,N_20240);
or U28291 (N_28291,N_22847,N_22684);
or U28292 (N_28292,N_20802,N_23987);
nor U28293 (N_28293,N_21293,N_23171);
xor U28294 (N_28294,N_22311,N_24099);
nand U28295 (N_28295,N_23247,N_23827);
nand U28296 (N_28296,N_24419,N_20515);
xor U28297 (N_28297,N_24750,N_24345);
and U28298 (N_28298,N_22465,N_23801);
and U28299 (N_28299,N_21384,N_20922);
and U28300 (N_28300,N_22906,N_23236);
nand U28301 (N_28301,N_22877,N_24345);
or U28302 (N_28302,N_24777,N_24442);
and U28303 (N_28303,N_20152,N_24815);
or U28304 (N_28304,N_22117,N_24084);
nand U28305 (N_28305,N_23347,N_23519);
nand U28306 (N_28306,N_22877,N_22729);
xor U28307 (N_28307,N_21520,N_24369);
and U28308 (N_28308,N_22259,N_22744);
or U28309 (N_28309,N_23576,N_24899);
and U28310 (N_28310,N_21754,N_21970);
or U28311 (N_28311,N_21109,N_21187);
and U28312 (N_28312,N_24779,N_22266);
nor U28313 (N_28313,N_22244,N_21802);
or U28314 (N_28314,N_20483,N_23351);
xnor U28315 (N_28315,N_23042,N_24015);
nor U28316 (N_28316,N_22271,N_22753);
nor U28317 (N_28317,N_24319,N_22288);
nor U28318 (N_28318,N_24621,N_20200);
or U28319 (N_28319,N_21623,N_24860);
nand U28320 (N_28320,N_23881,N_20934);
or U28321 (N_28321,N_22297,N_23796);
and U28322 (N_28322,N_22934,N_22294);
nor U28323 (N_28323,N_21495,N_21293);
and U28324 (N_28324,N_21745,N_20340);
nor U28325 (N_28325,N_22564,N_22488);
nand U28326 (N_28326,N_21888,N_21008);
nand U28327 (N_28327,N_22205,N_24538);
nor U28328 (N_28328,N_20948,N_20087);
or U28329 (N_28329,N_24352,N_24301);
nor U28330 (N_28330,N_21008,N_23692);
nand U28331 (N_28331,N_21799,N_20553);
nand U28332 (N_28332,N_22413,N_21226);
and U28333 (N_28333,N_20289,N_23359);
nand U28334 (N_28334,N_24151,N_24315);
nand U28335 (N_28335,N_20469,N_21734);
nor U28336 (N_28336,N_22627,N_20719);
nor U28337 (N_28337,N_20108,N_23139);
and U28338 (N_28338,N_24468,N_22473);
nor U28339 (N_28339,N_24675,N_24799);
and U28340 (N_28340,N_24108,N_21237);
and U28341 (N_28341,N_20557,N_24762);
nand U28342 (N_28342,N_23957,N_21889);
or U28343 (N_28343,N_21639,N_21308);
and U28344 (N_28344,N_23381,N_24281);
or U28345 (N_28345,N_20527,N_23031);
nand U28346 (N_28346,N_23142,N_20293);
nor U28347 (N_28347,N_24911,N_24852);
or U28348 (N_28348,N_23101,N_23590);
and U28349 (N_28349,N_22852,N_23240);
or U28350 (N_28350,N_20522,N_22781);
or U28351 (N_28351,N_20570,N_21326);
or U28352 (N_28352,N_24702,N_21456);
xnor U28353 (N_28353,N_24142,N_24855);
or U28354 (N_28354,N_21621,N_22439);
or U28355 (N_28355,N_23923,N_22419);
and U28356 (N_28356,N_24323,N_24042);
nand U28357 (N_28357,N_22611,N_24353);
nand U28358 (N_28358,N_22022,N_24660);
or U28359 (N_28359,N_21541,N_24541);
nor U28360 (N_28360,N_24987,N_21407);
or U28361 (N_28361,N_22454,N_22769);
nand U28362 (N_28362,N_20337,N_24322);
nand U28363 (N_28363,N_22459,N_23647);
or U28364 (N_28364,N_22661,N_23386);
and U28365 (N_28365,N_24921,N_24177);
and U28366 (N_28366,N_20464,N_20610);
and U28367 (N_28367,N_22333,N_21952);
nand U28368 (N_28368,N_22322,N_23953);
and U28369 (N_28369,N_23269,N_21553);
nor U28370 (N_28370,N_20493,N_20464);
nand U28371 (N_28371,N_20245,N_20106);
and U28372 (N_28372,N_22379,N_23481);
and U28373 (N_28373,N_24198,N_24825);
nand U28374 (N_28374,N_20652,N_23397);
nand U28375 (N_28375,N_24401,N_21392);
nand U28376 (N_28376,N_24778,N_23821);
and U28377 (N_28377,N_21433,N_21239);
and U28378 (N_28378,N_24358,N_21502);
nor U28379 (N_28379,N_23305,N_22442);
and U28380 (N_28380,N_24004,N_24709);
nor U28381 (N_28381,N_21760,N_23486);
nand U28382 (N_28382,N_20787,N_20789);
nand U28383 (N_28383,N_20388,N_23506);
and U28384 (N_28384,N_21307,N_24745);
or U28385 (N_28385,N_21078,N_21501);
nand U28386 (N_28386,N_24628,N_20680);
xnor U28387 (N_28387,N_21352,N_24235);
and U28388 (N_28388,N_20293,N_23564);
nor U28389 (N_28389,N_24453,N_23881);
and U28390 (N_28390,N_24537,N_22491);
nand U28391 (N_28391,N_20562,N_22679);
or U28392 (N_28392,N_24002,N_23648);
xor U28393 (N_28393,N_23402,N_20285);
nor U28394 (N_28394,N_21375,N_24830);
or U28395 (N_28395,N_24617,N_20730);
or U28396 (N_28396,N_23212,N_21816);
and U28397 (N_28397,N_20311,N_22932);
or U28398 (N_28398,N_22662,N_23061);
nor U28399 (N_28399,N_22320,N_24856);
nand U28400 (N_28400,N_23635,N_22477);
nand U28401 (N_28401,N_24656,N_20563);
xnor U28402 (N_28402,N_23008,N_22193);
xor U28403 (N_28403,N_23377,N_23759);
or U28404 (N_28404,N_23912,N_24883);
xor U28405 (N_28405,N_21300,N_24003);
or U28406 (N_28406,N_21030,N_20992);
nand U28407 (N_28407,N_24863,N_22553);
nand U28408 (N_28408,N_21130,N_20061);
or U28409 (N_28409,N_23928,N_23832);
and U28410 (N_28410,N_24367,N_23207);
nand U28411 (N_28411,N_24271,N_24626);
nand U28412 (N_28412,N_21837,N_20262);
or U28413 (N_28413,N_22785,N_24723);
nand U28414 (N_28414,N_23907,N_23342);
nor U28415 (N_28415,N_22183,N_22280);
nor U28416 (N_28416,N_23182,N_24298);
and U28417 (N_28417,N_21117,N_23746);
and U28418 (N_28418,N_21734,N_23763);
nor U28419 (N_28419,N_22820,N_22510);
nor U28420 (N_28420,N_22356,N_22493);
nand U28421 (N_28421,N_20563,N_21218);
or U28422 (N_28422,N_21433,N_21010);
or U28423 (N_28423,N_24725,N_21112);
or U28424 (N_28424,N_20865,N_21089);
and U28425 (N_28425,N_20612,N_20793);
nor U28426 (N_28426,N_23754,N_23082);
nand U28427 (N_28427,N_23376,N_24721);
xnor U28428 (N_28428,N_22557,N_20873);
nand U28429 (N_28429,N_24772,N_23513);
and U28430 (N_28430,N_23567,N_24596);
or U28431 (N_28431,N_20226,N_20076);
nand U28432 (N_28432,N_24916,N_22000);
nor U28433 (N_28433,N_22552,N_24939);
nor U28434 (N_28434,N_24926,N_22540);
xor U28435 (N_28435,N_20904,N_22892);
and U28436 (N_28436,N_20751,N_22406);
or U28437 (N_28437,N_24679,N_22976);
nor U28438 (N_28438,N_20845,N_22303);
and U28439 (N_28439,N_24480,N_21918);
nand U28440 (N_28440,N_23169,N_21453);
xor U28441 (N_28441,N_20616,N_23110);
nand U28442 (N_28442,N_22728,N_22992);
nor U28443 (N_28443,N_22612,N_23318);
and U28444 (N_28444,N_23932,N_22202);
or U28445 (N_28445,N_20944,N_24132);
nand U28446 (N_28446,N_20346,N_22400);
nand U28447 (N_28447,N_20510,N_21423);
nor U28448 (N_28448,N_21361,N_23596);
or U28449 (N_28449,N_21565,N_24410);
or U28450 (N_28450,N_22949,N_20374);
nor U28451 (N_28451,N_23731,N_22997);
or U28452 (N_28452,N_23080,N_24511);
nor U28453 (N_28453,N_24828,N_23716);
and U28454 (N_28454,N_20073,N_23396);
nor U28455 (N_28455,N_23516,N_20003);
nor U28456 (N_28456,N_20947,N_21298);
nand U28457 (N_28457,N_23566,N_24370);
nor U28458 (N_28458,N_21478,N_24634);
nor U28459 (N_28459,N_20365,N_22563);
xor U28460 (N_28460,N_24091,N_21559);
or U28461 (N_28461,N_21637,N_22731);
nor U28462 (N_28462,N_20474,N_21179);
nor U28463 (N_28463,N_24501,N_21175);
and U28464 (N_28464,N_21157,N_23373);
or U28465 (N_28465,N_21393,N_23961);
or U28466 (N_28466,N_23930,N_20900);
nor U28467 (N_28467,N_20556,N_20085);
or U28468 (N_28468,N_24660,N_20015);
nor U28469 (N_28469,N_20444,N_24641);
or U28470 (N_28470,N_22463,N_24076);
or U28471 (N_28471,N_24011,N_21482);
nor U28472 (N_28472,N_22011,N_21126);
nand U28473 (N_28473,N_23278,N_24723);
and U28474 (N_28474,N_21591,N_24610);
nand U28475 (N_28475,N_21097,N_23412);
and U28476 (N_28476,N_21219,N_22568);
nand U28477 (N_28477,N_23126,N_24319);
nand U28478 (N_28478,N_21445,N_22939);
nor U28479 (N_28479,N_24235,N_23395);
nor U28480 (N_28480,N_21960,N_22470);
nand U28481 (N_28481,N_22522,N_20815);
xnor U28482 (N_28482,N_22633,N_23844);
nand U28483 (N_28483,N_21990,N_24562);
nor U28484 (N_28484,N_21270,N_22709);
or U28485 (N_28485,N_22096,N_23921);
or U28486 (N_28486,N_24529,N_24965);
nor U28487 (N_28487,N_22488,N_20670);
nor U28488 (N_28488,N_20863,N_22701);
nor U28489 (N_28489,N_20480,N_24058);
nor U28490 (N_28490,N_24760,N_21408);
xor U28491 (N_28491,N_24992,N_24037);
nand U28492 (N_28492,N_21164,N_20087);
and U28493 (N_28493,N_24944,N_24235);
xnor U28494 (N_28494,N_21452,N_22811);
nand U28495 (N_28495,N_21255,N_23461);
nand U28496 (N_28496,N_20370,N_24116);
nor U28497 (N_28497,N_24364,N_23401);
or U28498 (N_28498,N_21777,N_21370);
nand U28499 (N_28499,N_23010,N_24769);
or U28500 (N_28500,N_22276,N_24106);
or U28501 (N_28501,N_22443,N_20017);
nand U28502 (N_28502,N_21467,N_24600);
nor U28503 (N_28503,N_22920,N_20445);
or U28504 (N_28504,N_24538,N_23067);
xor U28505 (N_28505,N_24808,N_24759);
or U28506 (N_28506,N_23703,N_23436);
nand U28507 (N_28507,N_22808,N_20610);
nor U28508 (N_28508,N_22378,N_23175);
nand U28509 (N_28509,N_23760,N_23111);
nor U28510 (N_28510,N_23933,N_21707);
nand U28511 (N_28511,N_23510,N_24174);
and U28512 (N_28512,N_24471,N_20127);
xnor U28513 (N_28513,N_21646,N_23405);
nand U28514 (N_28514,N_23451,N_21048);
nor U28515 (N_28515,N_20304,N_23713);
nand U28516 (N_28516,N_23686,N_23359);
and U28517 (N_28517,N_21379,N_23193);
and U28518 (N_28518,N_22716,N_22693);
nand U28519 (N_28519,N_24953,N_23479);
nor U28520 (N_28520,N_21941,N_21024);
nor U28521 (N_28521,N_22255,N_20451);
nand U28522 (N_28522,N_20969,N_20190);
xnor U28523 (N_28523,N_21703,N_24986);
or U28524 (N_28524,N_23309,N_23879);
or U28525 (N_28525,N_23442,N_23417);
or U28526 (N_28526,N_23241,N_20856);
nor U28527 (N_28527,N_22836,N_21316);
nand U28528 (N_28528,N_22653,N_21077);
nand U28529 (N_28529,N_23029,N_24664);
or U28530 (N_28530,N_22589,N_22178);
nor U28531 (N_28531,N_20511,N_21261);
nand U28532 (N_28532,N_20739,N_21538);
and U28533 (N_28533,N_23661,N_20565);
and U28534 (N_28534,N_22598,N_24434);
xor U28535 (N_28535,N_24905,N_24452);
or U28536 (N_28536,N_20064,N_23584);
nand U28537 (N_28537,N_23540,N_21911);
and U28538 (N_28538,N_24947,N_23904);
xnor U28539 (N_28539,N_21829,N_20190);
nand U28540 (N_28540,N_21440,N_22440);
nor U28541 (N_28541,N_24337,N_22571);
nand U28542 (N_28542,N_20672,N_20468);
and U28543 (N_28543,N_22377,N_20120);
or U28544 (N_28544,N_20518,N_21630);
or U28545 (N_28545,N_20483,N_20196);
and U28546 (N_28546,N_24705,N_22207);
or U28547 (N_28547,N_21136,N_23806);
or U28548 (N_28548,N_21916,N_24485);
xor U28549 (N_28549,N_23954,N_22455);
and U28550 (N_28550,N_21678,N_24176);
nand U28551 (N_28551,N_21179,N_22672);
or U28552 (N_28552,N_20734,N_24281);
or U28553 (N_28553,N_24534,N_20366);
or U28554 (N_28554,N_22284,N_22191);
and U28555 (N_28555,N_24708,N_24385);
or U28556 (N_28556,N_20971,N_20836);
nand U28557 (N_28557,N_24425,N_21881);
nor U28558 (N_28558,N_23636,N_23179);
and U28559 (N_28559,N_20722,N_23888);
or U28560 (N_28560,N_21871,N_22293);
nand U28561 (N_28561,N_21585,N_21775);
and U28562 (N_28562,N_20354,N_23167);
nand U28563 (N_28563,N_24385,N_23973);
or U28564 (N_28564,N_22994,N_21558);
and U28565 (N_28565,N_22553,N_21654);
or U28566 (N_28566,N_24228,N_21778);
and U28567 (N_28567,N_24363,N_23792);
nor U28568 (N_28568,N_21880,N_22364);
nor U28569 (N_28569,N_20237,N_24385);
or U28570 (N_28570,N_22779,N_20100);
nor U28571 (N_28571,N_24235,N_24845);
nor U28572 (N_28572,N_24852,N_22041);
xor U28573 (N_28573,N_22664,N_24400);
and U28574 (N_28574,N_20036,N_23390);
or U28575 (N_28575,N_22071,N_23318);
or U28576 (N_28576,N_20994,N_20231);
or U28577 (N_28577,N_20019,N_22932);
nand U28578 (N_28578,N_22255,N_21029);
and U28579 (N_28579,N_23347,N_23475);
nor U28580 (N_28580,N_20603,N_23497);
nand U28581 (N_28581,N_23417,N_24712);
and U28582 (N_28582,N_22069,N_22587);
and U28583 (N_28583,N_21918,N_24364);
xnor U28584 (N_28584,N_20594,N_24958);
nor U28585 (N_28585,N_23649,N_24418);
nand U28586 (N_28586,N_21081,N_24455);
nand U28587 (N_28587,N_23102,N_20048);
nand U28588 (N_28588,N_22107,N_21473);
or U28589 (N_28589,N_21844,N_20238);
nand U28590 (N_28590,N_24405,N_24953);
or U28591 (N_28591,N_22860,N_22571);
nand U28592 (N_28592,N_24201,N_24572);
nor U28593 (N_28593,N_22916,N_24093);
nor U28594 (N_28594,N_23772,N_22027);
nor U28595 (N_28595,N_24299,N_20093);
or U28596 (N_28596,N_24185,N_24223);
nand U28597 (N_28597,N_21338,N_22190);
and U28598 (N_28598,N_21945,N_20506);
xor U28599 (N_28599,N_21282,N_23471);
and U28600 (N_28600,N_21079,N_21009);
nor U28601 (N_28601,N_22708,N_22757);
and U28602 (N_28602,N_23078,N_24957);
or U28603 (N_28603,N_22790,N_20226);
nor U28604 (N_28604,N_22377,N_20127);
and U28605 (N_28605,N_20488,N_21767);
or U28606 (N_28606,N_24111,N_20580);
nand U28607 (N_28607,N_24715,N_21511);
and U28608 (N_28608,N_20667,N_22284);
nor U28609 (N_28609,N_24787,N_20645);
xor U28610 (N_28610,N_22722,N_24542);
or U28611 (N_28611,N_20711,N_23149);
or U28612 (N_28612,N_20055,N_20027);
and U28613 (N_28613,N_22011,N_22893);
xnor U28614 (N_28614,N_22487,N_24498);
nor U28615 (N_28615,N_20605,N_24234);
and U28616 (N_28616,N_23185,N_21182);
nand U28617 (N_28617,N_21155,N_20455);
or U28618 (N_28618,N_20842,N_23466);
nand U28619 (N_28619,N_21844,N_20388);
and U28620 (N_28620,N_24680,N_23731);
or U28621 (N_28621,N_21600,N_23706);
or U28622 (N_28622,N_22433,N_20333);
or U28623 (N_28623,N_22396,N_23521);
xnor U28624 (N_28624,N_20701,N_22906);
nor U28625 (N_28625,N_20598,N_23597);
and U28626 (N_28626,N_24283,N_24598);
or U28627 (N_28627,N_20594,N_21765);
or U28628 (N_28628,N_20468,N_22815);
or U28629 (N_28629,N_24783,N_22063);
and U28630 (N_28630,N_21770,N_23549);
and U28631 (N_28631,N_21365,N_24124);
or U28632 (N_28632,N_22794,N_20661);
and U28633 (N_28633,N_22911,N_23720);
nor U28634 (N_28634,N_22430,N_22543);
and U28635 (N_28635,N_22038,N_24725);
nor U28636 (N_28636,N_22214,N_24122);
and U28637 (N_28637,N_22092,N_21748);
nand U28638 (N_28638,N_20632,N_22379);
or U28639 (N_28639,N_21533,N_21036);
nand U28640 (N_28640,N_24032,N_22275);
nand U28641 (N_28641,N_24848,N_24471);
and U28642 (N_28642,N_20458,N_21596);
nor U28643 (N_28643,N_20170,N_23915);
xor U28644 (N_28644,N_23637,N_22504);
or U28645 (N_28645,N_21190,N_20541);
and U28646 (N_28646,N_21927,N_22697);
nand U28647 (N_28647,N_23100,N_22334);
or U28648 (N_28648,N_20389,N_24159);
nor U28649 (N_28649,N_22283,N_22963);
nor U28650 (N_28650,N_24779,N_22186);
xnor U28651 (N_28651,N_20034,N_24917);
or U28652 (N_28652,N_21383,N_21772);
nor U28653 (N_28653,N_24617,N_24075);
nand U28654 (N_28654,N_22380,N_20795);
nand U28655 (N_28655,N_21651,N_22816);
xor U28656 (N_28656,N_23081,N_24485);
and U28657 (N_28657,N_20708,N_20125);
xor U28658 (N_28658,N_22194,N_23756);
and U28659 (N_28659,N_20332,N_21953);
nand U28660 (N_28660,N_22834,N_20626);
or U28661 (N_28661,N_21713,N_20187);
or U28662 (N_28662,N_21250,N_23267);
nand U28663 (N_28663,N_21265,N_20920);
nand U28664 (N_28664,N_23630,N_23576);
nor U28665 (N_28665,N_21098,N_24851);
or U28666 (N_28666,N_20918,N_24888);
nand U28667 (N_28667,N_21106,N_22403);
and U28668 (N_28668,N_23025,N_24860);
nand U28669 (N_28669,N_20725,N_23974);
nor U28670 (N_28670,N_21475,N_23077);
or U28671 (N_28671,N_22307,N_20474);
and U28672 (N_28672,N_24171,N_23419);
xor U28673 (N_28673,N_21812,N_24561);
nor U28674 (N_28674,N_20858,N_20654);
nor U28675 (N_28675,N_24500,N_21752);
xnor U28676 (N_28676,N_23885,N_23679);
nor U28677 (N_28677,N_23179,N_23651);
nor U28678 (N_28678,N_20074,N_22772);
nor U28679 (N_28679,N_22884,N_20987);
nor U28680 (N_28680,N_24848,N_21894);
nor U28681 (N_28681,N_23046,N_21287);
or U28682 (N_28682,N_21274,N_24590);
or U28683 (N_28683,N_23012,N_20249);
nand U28684 (N_28684,N_21555,N_20841);
nand U28685 (N_28685,N_23195,N_23144);
nand U28686 (N_28686,N_24576,N_24977);
nor U28687 (N_28687,N_24165,N_21193);
nor U28688 (N_28688,N_23784,N_23125);
nor U28689 (N_28689,N_22782,N_24921);
nand U28690 (N_28690,N_22829,N_22782);
nor U28691 (N_28691,N_22941,N_24060);
xor U28692 (N_28692,N_20909,N_22674);
or U28693 (N_28693,N_21086,N_24011);
nor U28694 (N_28694,N_21992,N_22559);
or U28695 (N_28695,N_20397,N_22799);
nand U28696 (N_28696,N_23688,N_22635);
nand U28697 (N_28697,N_24569,N_24382);
nand U28698 (N_28698,N_23598,N_21387);
nand U28699 (N_28699,N_21087,N_24498);
and U28700 (N_28700,N_22311,N_24958);
or U28701 (N_28701,N_21754,N_20511);
or U28702 (N_28702,N_23136,N_24963);
nand U28703 (N_28703,N_23649,N_20718);
or U28704 (N_28704,N_24828,N_24238);
nand U28705 (N_28705,N_24298,N_23809);
or U28706 (N_28706,N_22454,N_24887);
nor U28707 (N_28707,N_20142,N_23393);
nand U28708 (N_28708,N_20279,N_23786);
or U28709 (N_28709,N_24996,N_21598);
nor U28710 (N_28710,N_23834,N_22170);
nor U28711 (N_28711,N_23189,N_23126);
and U28712 (N_28712,N_20832,N_21223);
nand U28713 (N_28713,N_22640,N_20863);
or U28714 (N_28714,N_24603,N_21289);
nor U28715 (N_28715,N_20567,N_23942);
nor U28716 (N_28716,N_20157,N_20668);
nand U28717 (N_28717,N_21680,N_21099);
or U28718 (N_28718,N_23793,N_22712);
nand U28719 (N_28719,N_20722,N_22608);
nand U28720 (N_28720,N_21987,N_22147);
nor U28721 (N_28721,N_22442,N_21419);
xnor U28722 (N_28722,N_23537,N_20402);
nand U28723 (N_28723,N_24593,N_24528);
nor U28724 (N_28724,N_22150,N_24357);
or U28725 (N_28725,N_20242,N_23392);
nor U28726 (N_28726,N_20135,N_24015);
and U28727 (N_28727,N_20726,N_24319);
or U28728 (N_28728,N_20569,N_20455);
or U28729 (N_28729,N_24269,N_22269);
and U28730 (N_28730,N_23273,N_20593);
nor U28731 (N_28731,N_24737,N_23150);
xor U28732 (N_28732,N_20397,N_20938);
nand U28733 (N_28733,N_24741,N_24940);
nand U28734 (N_28734,N_21631,N_23930);
or U28735 (N_28735,N_23632,N_24871);
or U28736 (N_28736,N_20971,N_24626);
or U28737 (N_28737,N_23059,N_22953);
or U28738 (N_28738,N_23018,N_24550);
and U28739 (N_28739,N_24066,N_21659);
or U28740 (N_28740,N_24876,N_20937);
and U28741 (N_28741,N_21090,N_21818);
nand U28742 (N_28742,N_21606,N_20855);
or U28743 (N_28743,N_20189,N_23619);
nand U28744 (N_28744,N_24889,N_21665);
nor U28745 (N_28745,N_24537,N_20840);
nand U28746 (N_28746,N_22502,N_24137);
or U28747 (N_28747,N_23392,N_20809);
and U28748 (N_28748,N_24225,N_21197);
nand U28749 (N_28749,N_21084,N_24706);
and U28750 (N_28750,N_23617,N_24116);
and U28751 (N_28751,N_23462,N_22572);
nor U28752 (N_28752,N_22987,N_22070);
xnor U28753 (N_28753,N_24948,N_23749);
or U28754 (N_28754,N_23069,N_24584);
or U28755 (N_28755,N_24689,N_20444);
and U28756 (N_28756,N_21010,N_23377);
or U28757 (N_28757,N_20846,N_20883);
and U28758 (N_28758,N_20805,N_20771);
or U28759 (N_28759,N_24473,N_23370);
nor U28760 (N_28760,N_21993,N_24827);
nor U28761 (N_28761,N_22762,N_21424);
or U28762 (N_28762,N_21693,N_20322);
and U28763 (N_28763,N_23372,N_24108);
and U28764 (N_28764,N_21270,N_24198);
or U28765 (N_28765,N_23049,N_22732);
xor U28766 (N_28766,N_20005,N_21614);
and U28767 (N_28767,N_20313,N_20886);
nand U28768 (N_28768,N_20771,N_24775);
nand U28769 (N_28769,N_23144,N_21243);
nand U28770 (N_28770,N_24565,N_23839);
or U28771 (N_28771,N_24294,N_24127);
nor U28772 (N_28772,N_21332,N_23457);
nand U28773 (N_28773,N_23149,N_21483);
nand U28774 (N_28774,N_23171,N_24713);
nand U28775 (N_28775,N_21240,N_20857);
xnor U28776 (N_28776,N_23459,N_23083);
nand U28777 (N_28777,N_21569,N_23664);
or U28778 (N_28778,N_21626,N_23006);
nor U28779 (N_28779,N_24167,N_22226);
and U28780 (N_28780,N_21698,N_22318);
nand U28781 (N_28781,N_23344,N_20186);
nor U28782 (N_28782,N_20859,N_22708);
nand U28783 (N_28783,N_20110,N_21832);
xnor U28784 (N_28784,N_23302,N_20072);
nand U28785 (N_28785,N_23429,N_22297);
nand U28786 (N_28786,N_23660,N_23188);
nor U28787 (N_28787,N_23176,N_23377);
xor U28788 (N_28788,N_22975,N_23251);
nand U28789 (N_28789,N_21383,N_21897);
or U28790 (N_28790,N_22572,N_22787);
xnor U28791 (N_28791,N_21242,N_20453);
nand U28792 (N_28792,N_23340,N_21609);
and U28793 (N_28793,N_22486,N_21652);
or U28794 (N_28794,N_20430,N_20468);
nor U28795 (N_28795,N_21755,N_22322);
nor U28796 (N_28796,N_23141,N_24462);
nand U28797 (N_28797,N_20021,N_21384);
or U28798 (N_28798,N_22493,N_23271);
nor U28799 (N_28799,N_24992,N_20249);
nand U28800 (N_28800,N_21249,N_24830);
nand U28801 (N_28801,N_21742,N_24464);
or U28802 (N_28802,N_21493,N_24948);
xnor U28803 (N_28803,N_20739,N_20911);
nor U28804 (N_28804,N_22487,N_23496);
nand U28805 (N_28805,N_22493,N_24505);
nand U28806 (N_28806,N_24168,N_24669);
or U28807 (N_28807,N_21336,N_22158);
xnor U28808 (N_28808,N_21644,N_21056);
nor U28809 (N_28809,N_20596,N_20057);
nor U28810 (N_28810,N_22893,N_22083);
nand U28811 (N_28811,N_24241,N_23783);
and U28812 (N_28812,N_23637,N_21077);
nand U28813 (N_28813,N_22817,N_23082);
nor U28814 (N_28814,N_23282,N_24386);
nor U28815 (N_28815,N_21262,N_21638);
nand U28816 (N_28816,N_20079,N_21816);
or U28817 (N_28817,N_21356,N_20937);
nor U28818 (N_28818,N_24843,N_21026);
nor U28819 (N_28819,N_20371,N_21980);
or U28820 (N_28820,N_24393,N_22994);
nor U28821 (N_28821,N_24439,N_23488);
nor U28822 (N_28822,N_23282,N_23357);
nand U28823 (N_28823,N_22714,N_20333);
nand U28824 (N_28824,N_24233,N_21274);
nand U28825 (N_28825,N_24280,N_21205);
nand U28826 (N_28826,N_20834,N_23615);
nor U28827 (N_28827,N_20326,N_20920);
nor U28828 (N_28828,N_20235,N_23585);
and U28829 (N_28829,N_20059,N_21753);
nand U28830 (N_28830,N_20232,N_24935);
nand U28831 (N_28831,N_20361,N_22923);
and U28832 (N_28832,N_21271,N_21851);
or U28833 (N_28833,N_24945,N_23878);
and U28834 (N_28834,N_20514,N_24485);
nor U28835 (N_28835,N_23335,N_21421);
or U28836 (N_28836,N_20468,N_24470);
or U28837 (N_28837,N_24149,N_23485);
and U28838 (N_28838,N_21826,N_23893);
nand U28839 (N_28839,N_24456,N_21843);
and U28840 (N_28840,N_23539,N_24826);
and U28841 (N_28841,N_23930,N_20259);
or U28842 (N_28842,N_24084,N_23087);
and U28843 (N_28843,N_20314,N_21929);
and U28844 (N_28844,N_20183,N_22701);
or U28845 (N_28845,N_20858,N_22042);
or U28846 (N_28846,N_20280,N_23609);
nand U28847 (N_28847,N_23426,N_20895);
nand U28848 (N_28848,N_21238,N_21206);
nand U28849 (N_28849,N_23605,N_23541);
nand U28850 (N_28850,N_22835,N_20440);
nor U28851 (N_28851,N_23485,N_21824);
or U28852 (N_28852,N_24917,N_23613);
xor U28853 (N_28853,N_21512,N_22591);
or U28854 (N_28854,N_22809,N_24378);
nand U28855 (N_28855,N_23927,N_23428);
nor U28856 (N_28856,N_20931,N_22454);
nor U28857 (N_28857,N_20046,N_22449);
or U28858 (N_28858,N_22647,N_24022);
nand U28859 (N_28859,N_21785,N_20221);
or U28860 (N_28860,N_21840,N_21656);
and U28861 (N_28861,N_23481,N_22397);
or U28862 (N_28862,N_20630,N_23505);
nand U28863 (N_28863,N_21797,N_21179);
nand U28864 (N_28864,N_23946,N_23903);
xor U28865 (N_28865,N_22616,N_22648);
or U28866 (N_28866,N_23480,N_21617);
nor U28867 (N_28867,N_21820,N_22456);
and U28868 (N_28868,N_20826,N_20774);
nor U28869 (N_28869,N_21338,N_22891);
and U28870 (N_28870,N_22922,N_24847);
nand U28871 (N_28871,N_22942,N_21444);
or U28872 (N_28872,N_21418,N_24276);
nor U28873 (N_28873,N_23813,N_23684);
nor U28874 (N_28874,N_21901,N_20107);
and U28875 (N_28875,N_24750,N_21216);
nand U28876 (N_28876,N_24218,N_20314);
nor U28877 (N_28877,N_22848,N_23631);
nand U28878 (N_28878,N_20087,N_23742);
nor U28879 (N_28879,N_24004,N_22683);
or U28880 (N_28880,N_20465,N_21444);
or U28881 (N_28881,N_20463,N_22674);
and U28882 (N_28882,N_21226,N_20690);
nand U28883 (N_28883,N_21709,N_24039);
xnor U28884 (N_28884,N_24113,N_23735);
and U28885 (N_28885,N_23459,N_22095);
or U28886 (N_28886,N_23488,N_23186);
nand U28887 (N_28887,N_22765,N_23056);
or U28888 (N_28888,N_21297,N_20163);
nand U28889 (N_28889,N_20864,N_24924);
and U28890 (N_28890,N_24304,N_22701);
nor U28891 (N_28891,N_24812,N_20839);
nand U28892 (N_28892,N_24416,N_22847);
nor U28893 (N_28893,N_22653,N_22672);
nand U28894 (N_28894,N_20286,N_23871);
and U28895 (N_28895,N_23506,N_21548);
nand U28896 (N_28896,N_23815,N_24210);
and U28897 (N_28897,N_23756,N_22188);
nor U28898 (N_28898,N_20258,N_24930);
xor U28899 (N_28899,N_21098,N_23819);
or U28900 (N_28900,N_23334,N_22909);
or U28901 (N_28901,N_21664,N_21218);
nand U28902 (N_28902,N_23607,N_23845);
nand U28903 (N_28903,N_24096,N_23175);
nor U28904 (N_28904,N_23275,N_21748);
nor U28905 (N_28905,N_20435,N_20387);
nor U28906 (N_28906,N_20417,N_22357);
nor U28907 (N_28907,N_21139,N_20440);
and U28908 (N_28908,N_21017,N_21455);
or U28909 (N_28909,N_20341,N_23424);
nand U28910 (N_28910,N_24998,N_23570);
nor U28911 (N_28911,N_20484,N_20987);
nor U28912 (N_28912,N_23037,N_22243);
and U28913 (N_28913,N_21888,N_21781);
nor U28914 (N_28914,N_24741,N_22193);
xnor U28915 (N_28915,N_21848,N_22872);
and U28916 (N_28916,N_22112,N_20861);
or U28917 (N_28917,N_20598,N_24834);
and U28918 (N_28918,N_23564,N_22578);
or U28919 (N_28919,N_20177,N_20578);
nand U28920 (N_28920,N_24607,N_20757);
nor U28921 (N_28921,N_23859,N_21125);
or U28922 (N_28922,N_24295,N_23397);
nand U28923 (N_28923,N_22410,N_21469);
xnor U28924 (N_28924,N_22753,N_24056);
nand U28925 (N_28925,N_23606,N_24641);
or U28926 (N_28926,N_24261,N_22596);
nand U28927 (N_28927,N_21002,N_23224);
nor U28928 (N_28928,N_20666,N_24055);
and U28929 (N_28929,N_22009,N_23339);
nor U28930 (N_28930,N_24173,N_22425);
or U28931 (N_28931,N_24849,N_24156);
nor U28932 (N_28932,N_20772,N_20037);
and U28933 (N_28933,N_20434,N_23036);
nor U28934 (N_28934,N_21704,N_21902);
or U28935 (N_28935,N_21859,N_22669);
nand U28936 (N_28936,N_24299,N_24408);
nor U28937 (N_28937,N_23519,N_23911);
nand U28938 (N_28938,N_22113,N_20990);
nand U28939 (N_28939,N_24010,N_24097);
nand U28940 (N_28940,N_20759,N_20705);
nor U28941 (N_28941,N_23334,N_24590);
nor U28942 (N_28942,N_22174,N_24177);
or U28943 (N_28943,N_21492,N_20505);
or U28944 (N_28944,N_24385,N_22995);
nand U28945 (N_28945,N_23890,N_20848);
nor U28946 (N_28946,N_24583,N_22855);
nor U28947 (N_28947,N_20539,N_20200);
nand U28948 (N_28948,N_21837,N_23801);
and U28949 (N_28949,N_22192,N_20837);
or U28950 (N_28950,N_23277,N_24989);
nand U28951 (N_28951,N_23250,N_20220);
nand U28952 (N_28952,N_20185,N_21983);
and U28953 (N_28953,N_22806,N_20515);
nor U28954 (N_28954,N_20864,N_22796);
nor U28955 (N_28955,N_23842,N_23880);
nand U28956 (N_28956,N_22782,N_21728);
nor U28957 (N_28957,N_22637,N_23225);
nand U28958 (N_28958,N_22135,N_22353);
and U28959 (N_28959,N_21982,N_21139);
and U28960 (N_28960,N_24546,N_21721);
nand U28961 (N_28961,N_20805,N_22029);
nor U28962 (N_28962,N_20892,N_23383);
or U28963 (N_28963,N_22057,N_22832);
nor U28964 (N_28964,N_21017,N_20263);
or U28965 (N_28965,N_23243,N_23424);
xor U28966 (N_28966,N_22638,N_23057);
nand U28967 (N_28967,N_21082,N_23710);
and U28968 (N_28968,N_20729,N_20901);
nor U28969 (N_28969,N_24260,N_20568);
nor U28970 (N_28970,N_22254,N_22973);
nand U28971 (N_28971,N_24077,N_23389);
and U28972 (N_28972,N_21346,N_21870);
or U28973 (N_28973,N_22421,N_24487);
nor U28974 (N_28974,N_20878,N_20231);
xnor U28975 (N_28975,N_20269,N_21689);
nor U28976 (N_28976,N_23482,N_22379);
nand U28977 (N_28977,N_21520,N_22350);
or U28978 (N_28978,N_23744,N_24771);
nor U28979 (N_28979,N_23395,N_22150);
and U28980 (N_28980,N_22750,N_20201);
or U28981 (N_28981,N_22890,N_24678);
nor U28982 (N_28982,N_20504,N_23684);
nand U28983 (N_28983,N_20731,N_21471);
nor U28984 (N_28984,N_23980,N_21208);
nor U28985 (N_28985,N_24964,N_20160);
nor U28986 (N_28986,N_24627,N_21389);
nor U28987 (N_28987,N_24250,N_21624);
nand U28988 (N_28988,N_20479,N_20874);
or U28989 (N_28989,N_24763,N_23907);
nand U28990 (N_28990,N_20588,N_23773);
nand U28991 (N_28991,N_23698,N_20250);
nor U28992 (N_28992,N_24346,N_23463);
or U28993 (N_28993,N_24461,N_20617);
nand U28994 (N_28994,N_23987,N_21448);
and U28995 (N_28995,N_23211,N_23856);
and U28996 (N_28996,N_22832,N_21823);
xnor U28997 (N_28997,N_22589,N_20473);
and U28998 (N_28998,N_24677,N_23125);
nand U28999 (N_28999,N_22113,N_20566);
nor U29000 (N_29000,N_24615,N_24650);
or U29001 (N_29001,N_22991,N_20037);
and U29002 (N_29002,N_24658,N_23609);
nor U29003 (N_29003,N_23997,N_21587);
nand U29004 (N_29004,N_20376,N_23146);
xnor U29005 (N_29005,N_22339,N_20463);
or U29006 (N_29006,N_22636,N_21492);
or U29007 (N_29007,N_24722,N_23602);
xor U29008 (N_29008,N_23088,N_22659);
and U29009 (N_29009,N_23929,N_22300);
nand U29010 (N_29010,N_23116,N_24035);
and U29011 (N_29011,N_24572,N_23201);
or U29012 (N_29012,N_23665,N_22484);
nand U29013 (N_29013,N_24959,N_22330);
nand U29014 (N_29014,N_22529,N_22724);
nor U29015 (N_29015,N_20597,N_23370);
nand U29016 (N_29016,N_20206,N_24433);
xor U29017 (N_29017,N_21391,N_24685);
nand U29018 (N_29018,N_23294,N_22173);
nor U29019 (N_29019,N_21611,N_20331);
xor U29020 (N_29020,N_21906,N_24353);
or U29021 (N_29021,N_22072,N_23268);
nor U29022 (N_29022,N_21682,N_23757);
or U29023 (N_29023,N_21236,N_24194);
or U29024 (N_29024,N_20244,N_23783);
or U29025 (N_29025,N_21049,N_20519);
nor U29026 (N_29026,N_24347,N_24299);
nand U29027 (N_29027,N_20144,N_20294);
nand U29028 (N_29028,N_24968,N_22056);
and U29029 (N_29029,N_20396,N_24043);
or U29030 (N_29030,N_22293,N_20049);
and U29031 (N_29031,N_23235,N_21315);
or U29032 (N_29032,N_24275,N_24991);
nor U29033 (N_29033,N_24411,N_24904);
or U29034 (N_29034,N_24975,N_20131);
nor U29035 (N_29035,N_24595,N_20008);
or U29036 (N_29036,N_23780,N_20494);
nor U29037 (N_29037,N_24088,N_24623);
nor U29038 (N_29038,N_24383,N_23041);
and U29039 (N_29039,N_24283,N_22088);
nor U29040 (N_29040,N_21038,N_24784);
nand U29041 (N_29041,N_21699,N_22264);
nand U29042 (N_29042,N_22021,N_24250);
and U29043 (N_29043,N_22022,N_21672);
and U29044 (N_29044,N_23494,N_22277);
and U29045 (N_29045,N_22939,N_22784);
nor U29046 (N_29046,N_21130,N_24199);
nand U29047 (N_29047,N_21337,N_21211);
nor U29048 (N_29048,N_24522,N_23198);
and U29049 (N_29049,N_21191,N_21838);
nand U29050 (N_29050,N_22615,N_23797);
nand U29051 (N_29051,N_20823,N_23054);
nand U29052 (N_29052,N_23262,N_22816);
or U29053 (N_29053,N_23818,N_20314);
and U29054 (N_29054,N_20944,N_24347);
and U29055 (N_29055,N_24330,N_24583);
nand U29056 (N_29056,N_23411,N_21372);
nand U29057 (N_29057,N_21483,N_21301);
or U29058 (N_29058,N_23904,N_21260);
and U29059 (N_29059,N_24445,N_21339);
nand U29060 (N_29060,N_24095,N_24083);
and U29061 (N_29061,N_20943,N_23204);
and U29062 (N_29062,N_20640,N_23105);
and U29063 (N_29063,N_21015,N_23861);
nand U29064 (N_29064,N_23948,N_22570);
or U29065 (N_29065,N_21822,N_22287);
and U29066 (N_29066,N_20133,N_24858);
nor U29067 (N_29067,N_22216,N_20168);
and U29068 (N_29068,N_21502,N_23036);
or U29069 (N_29069,N_23671,N_20481);
and U29070 (N_29070,N_21942,N_20141);
or U29071 (N_29071,N_21428,N_22250);
and U29072 (N_29072,N_20935,N_21466);
and U29073 (N_29073,N_22868,N_24892);
and U29074 (N_29074,N_23219,N_21974);
and U29075 (N_29075,N_24399,N_24544);
nor U29076 (N_29076,N_23122,N_21605);
or U29077 (N_29077,N_20927,N_21111);
and U29078 (N_29078,N_23969,N_22542);
and U29079 (N_29079,N_21049,N_21874);
nand U29080 (N_29080,N_22339,N_23512);
or U29081 (N_29081,N_21718,N_21009);
nand U29082 (N_29082,N_20579,N_22284);
nand U29083 (N_29083,N_24892,N_21512);
nand U29084 (N_29084,N_22356,N_22020);
nor U29085 (N_29085,N_24797,N_24884);
nor U29086 (N_29086,N_23215,N_22387);
or U29087 (N_29087,N_24639,N_20141);
nand U29088 (N_29088,N_24987,N_20166);
and U29089 (N_29089,N_24184,N_23739);
or U29090 (N_29090,N_22470,N_24638);
xor U29091 (N_29091,N_24328,N_20737);
xnor U29092 (N_29092,N_20268,N_21564);
nand U29093 (N_29093,N_21374,N_23100);
xor U29094 (N_29094,N_20524,N_20742);
and U29095 (N_29095,N_23089,N_24602);
nand U29096 (N_29096,N_24673,N_22248);
nor U29097 (N_29097,N_20220,N_20346);
nand U29098 (N_29098,N_22609,N_22753);
nor U29099 (N_29099,N_23032,N_21772);
nor U29100 (N_29100,N_24721,N_20479);
nor U29101 (N_29101,N_21227,N_20261);
or U29102 (N_29102,N_21524,N_22358);
or U29103 (N_29103,N_21324,N_23651);
or U29104 (N_29104,N_24932,N_20098);
xor U29105 (N_29105,N_24904,N_20285);
xor U29106 (N_29106,N_20215,N_22282);
or U29107 (N_29107,N_20437,N_23474);
or U29108 (N_29108,N_24940,N_23479);
and U29109 (N_29109,N_20743,N_23093);
nor U29110 (N_29110,N_23619,N_20172);
xnor U29111 (N_29111,N_22827,N_20450);
nand U29112 (N_29112,N_22427,N_22859);
nand U29113 (N_29113,N_21316,N_20821);
or U29114 (N_29114,N_22206,N_23392);
or U29115 (N_29115,N_22131,N_22312);
or U29116 (N_29116,N_21464,N_20862);
nor U29117 (N_29117,N_23903,N_21072);
or U29118 (N_29118,N_20389,N_21890);
nand U29119 (N_29119,N_21965,N_24721);
xor U29120 (N_29120,N_21837,N_24456);
and U29121 (N_29121,N_23908,N_20358);
or U29122 (N_29122,N_21672,N_23389);
nor U29123 (N_29123,N_20337,N_24465);
nor U29124 (N_29124,N_22811,N_23998);
nand U29125 (N_29125,N_24253,N_22677);
nand U29126 (N_29126,N_21748,N_24611);
nor U29127 (N_29127,N_24014,N_22455);
nor U29128 (N_29128,N_23969,N_24576);
or U29129 (N_29129,N_24051,N_20695);
nand U29130 (N_29130,N_21591,N_21103);
nor U29131 (N_29131,N_23859,N_21586);
nor U29132 (N_29132,N_23909,N_24946);
or U29133 (N_29133,N_21518,N_22736);
nand U29134 (N_29134,N_23954,N_21867);
nand U29135 (N_29135,N_24039,N_21166);
and U29136 (N_29136,N_20294,N_23586);
and U29137 (N_29137,N_20886,N_23849);
nor U29138 (N_29138,N_22150,N_23815);
xor U29139 (N_29139,N_22449,N_23725);
nand U29140 (N_29140,N_24768,N_22988);
nand U29141 (N_29141,N_23783,N_22803);
nand U29142 (N_29142,N_21301,N_23902);
xor U29143 (N_29143,N_21010,N_21203);
nor U29144 (N_29144,N_24808,N_20195);
or U29145 (N_29145,N_22260,N_23310);
nand U29146 (N_29146,N_22708,N_24779);
and U29147 (N_29147,N_21468,N_23459);
and U29148 (N_29148,N_23461,N_24963);
nand U29149 (N_29149,N_23860,N_21629);
or U29150 (N_29150,N_22528,N_21742);
and U29151 (N_29151,N_24729,N_23606);
nor U29152 (N_29152,N_21571,N_24084);
nor U29153 (N_29153,N_21516,N_24404);
and U29154 (N_29154,N_20852,N_21766);
or U29155 (N_29155,N_22052,N_24151);
and U29156 (N_29156,N_24961,N_22529);
and U29157 (N_29157,N_20549,N_21144);
or U29158 (N_29158,N_21874,N_22263);
xnor U29159 (N_29159,N_20824,N_23074);
and U29160 (N_29160,N_21136,N_24340);
or U29161 (N_29161,N_20794,N_24863);
and U29162 (N_29162,N_21057,N_23560);
and U29163 (N_29163,N_24723,N_21646);
and U29164 (N_29164,N_22973,N_22555);
and U29165 (N_29165,N_20026,N_24770);
and U29166 (N_29166,N_22525,N_21749);
nor U29167 (N_29167,N_20049,N_24317);
or U29168 (N_29168,N_21596,N_22880);
or U29169 (N_29169,N_20069,N_20256);
and U29170 (N_29170,N_20142,N_22059);
and U29171 (N_29171,N_22615,N_21387);
nand U29172 (N_29172,N_20750,N_24921);
nand U29173 (N_29173,N_20245,N_23951);
xnor U29174 (N_29174,N_24141,N_23192);
nand U29175 (N_29175,N_21895,N_20698);
nor U29176 (N_29176,N_20030,N_21641);
xnor U29177 (N_29177,N_23520,N_22033);
nor U29178 (N_29178,N_21411,N_24829);
nand U29179 (N_29179,N_20980,N_20945);
nand U29180 (N_29180,N_24477,N_21426);
nand U29181 (N_29181,N_21638,N_24764);
and U29182 (N_29182,N_23367,N_22857);
or U29183 (N_29183,N_23847,N_23796);
or U29184 (N_29184,N_23133,N_24511);
nand U29185 (N_29185,N_24461,N_20760);
nor U29186 (N_29186,N_21867,N_22013);
and U29187 (N_29187,N_22625,N_20576);
or U29188 (N_29188,N_22051,N_23670);
xnor U29189 (N_29189,N_24044,N_21751);
nand U29190 (N_29190,N_23985,N_22195);
or U29191 (N_29191,N_24079,N_20883);
or U29192 (N_29192,N_20705,N_22197);
nand U29193 (N_29193,N_20900,N_23172);
and U29194 (N_29194,N_20684,N_22262);
or U29195 (N_29195,N_24756,N_21022);
nor U29196 (N_29196,N_20969,N_24540);
or U29197 (N_29197,N_21451,N_21726);
and U29198 (N_29198,N_21707,N_22441);
nand U29199 (N_29199,N_22730,N_23452);
nor U29200 (N_29200,N_20758,N_20986);
or U29201 (N_29201,N_22351,N_23457);
and U29202 (N_29202,N_21812,N_23510);
and U29203 (N_29203,N_23418,N_23900);
and U29204 (N_29204,N_20487,N_20062);
nor U29205 (N_29205,N_22527,N_24024);
or U29206 (N_29206,N_22708,N_23854);
nor U29207 (N_29207,N_23403,N_21425);
xnor U29208 (N_29208,N_24671,N_21288);
nor U29209 (N_29209,N_22750,N_23050);
nand U29210 (N_29210,N_23975,N_22377);
nor U29211 (N_29211,N_23153,N_23715);
nand U29212 (N_29212,N_24768,N_22420);
or U29213 (N_29213,N_24303,N_21187);
and U29214 (N_29214,N_24373,N_20618);
or U29215 (N_29215,N_24085,N_21196);
xor U29216 (N_29216,N_22107,N_21278);
nand U29217 (N_29217,N_24795,N_21268);
xnor U29218 (N_29218,N_20882,N_20392);
or U29219 (N_29219,N_21625,N_23474);
nand U29220 (N_29220,N_20770,N_23555);
nand U29221 (N_29221,N_22030,N_22698);
nand U29222 (N_29222,N_24543,N_21504);
nand U29223 (N_29223,N_20137,N_22054);
or U29224 (N_29224,N_23793,N_24883);
and U29225 (N_29225,N_20157,N_21239);
nor U29226 (N_29226,N_22493,N_21938);
xnor U29227 (N_29227,N_22213,N_24429);
nand U29228 (N_29228,N_22402,N_22147);
and U29229 (N_29229,N_23601,N_22230);
nor U29230 (N_29230,N_21413,N_23699);
nand U29231 (N_29231,N_23727,N_23106);
nor U29232 (N_29232,N_24927,N_24326);
and U29233 (N_29233,N_23824,N_24818);
nand U29234 (N_29234,N_23377,N_21186);
nor U29235 (N_29235,N_23343,N_24244);
nor U29236 (N_29236,N_24744,N_23876);
nand U29237 (N_29237,N_20813,N_20586);
xor U29238 (N_29238,N_23579,N_22419);
and U29239 (N_29239,N_24619,N_22000);
nor U29240 (N_29240,N_20870,N_24153);
nor U29241 (N_29241,N_22423,N_20175);
nor U29242 (N_29242,N_21269,N_20106);
nand U29243 (N_29243,N_23464,N_24527);
nor U29244 (N_29244,N_24828,N_20676);
xor U29245 (N_29245,N_22614,N_20629);
or U29246 (N_29246,N_23555,N_24006);
nand U29247 (N_29247,N_23376,N_22420);
nand U29248 (N_29248,N_23631,N_20945);
and U29249 (N_29249,N_21702,N_20239);
xnor U29250 (N_29250,N_24877,N_22793);
and U29251 (N_29251,N_21531,N_23221);
or U29252 (N_29252,N_24456,N_21045);
or U29253 (N_29253,N_23871,N_23308);
or U29254 (N_29254,N_23588,N_21420);
xnor U29255 (N_29255,N_21435,N_21340);
nand U29256 (N_29256,N_22632,N_22924);
and U29257 (N_29257,N_20397,N_24873);
or U29258 (N_29258,N_24107,N_22303);
or U29259 (N_29259,N_23761,N_21008);
nor U29260 (N_29260,N_20158,N_22628);
and U29261 (N_29261,N_24440,N_23452);
nand U29262 (N_29262,N_22072,N_23866);
nor U29263 (N_29263,N_21945,N_21470);
xnor U29264 (N_29264,N_20499,N_20949);
and U29265 (N_29265,N_23448,N_20998);
and U29266 (N_29266,N_22655,N_22299);
nor U29267 (N_29267,N_24305,N_22034);
and U29268 (N_29268,N_23080,N_23348);
or U29269 (N_29269,N_23065,N_20738);
or U29270 (N_29270,N_20217,N_22924);
nor U29271 (N_29271,N_21790,N_22941);
nand U29272 (N_29272,N_21752,N_21288);
nand U29273 (N_29273,N_21597,N_24681);
and U29274 (N_29274,N_21622,N_24491);
nand U29275 (N_29275,N_20697,N_21312);
nor U29276 (N_29276,N_21151,N_23094);
nand U29277 (N_29277,N_23899,N_20594);
nand U29278 (N_29278,N_24893,N_21885);
nor U29279 (N_29279,N_22166,N_21243);
nor U29280 (N_29280,N_24048,N_24817);
and U29281 (N_29281,N_21821,N_21134);
xnor U29282 (N_29282,N_21837,N_20267);
nor U29283 (N_29283,N_23915,N_21151);
nor U29284 (N_29284,N_22659,N_23466);
nand U29285 (N_29285,N_21792,N_23625);
or U29286 (N_29286,N_20728,N_22613);
or U29287 (N_29287,N_21900,N_20256);
and U29288 (N_29288,N_24767,N_22331);
or U29289 (N_29289,N_23941,N_22695);
or U29290 (N_29290,N_24486,N_20647);
nor U29291 (N_29291,N_23189,N_20795);
nand U29292 (N_29292,N_24235,N_24593);
and U29293 (N_29293,N_24381,N_21800);
nor U29294 (N_29294,N_20015,N_22152);
or U29295 (N_29295,N_22192,N_23517);
nand U29296 (N_29296,N_21787,N_24338);
or U29297 (N_29297,N_24147,N_21338);
nand U29298 (N_29298,N_22090,N_23864);
nand U29299 (N_29299,N_23499,N_20983);
nor U29300 (N_29300,N_22697,N_21536);
nand U29301 (N_29301,N_21962,N_23449);
nand U29302 (N_29302,N_21212,N_23560);
nand U29303 (N_29303,N_23464,N_23487);
nand U29304 (N_29304,N_20852,N_23429);
or U29305 (N_29305,N_20550,N_21242);
nand U29306 (N_29306,N_24683,N_20333);
nand U29307 (N_29307,N_20741,N_23304);
nand U29308 (N_29308,N_21419,N_23411);
nor U29309 (N_29309,N_24108,N_22958);
nand U29310 (N_29310,N_22902,N_23573);
nand U29311 (N_29311,N_22219,N_21536);
nand U29312 (N_29312,N_21146,N_23833);
nor U29313 (N_29313,N_21222,N_22241);
nand U29314 (N_29314,N_21657,N_23682);
and U29315 (N_29315,N_24820,N_24860);
nand U29316 (N_29316,N_24075,N_23240);
nor U29317 (N_29317,N_24956,N_21909);
nand U29318 (N_29318,N_22245,N_24186);
nor U29319 (N_29319,N_20851,N_21733);
nor U29320 (N_29320,N_20244,N_23155);
xor U29321 (N_29321,N_23321,N_24657);
and U29322 (N_29322,N_23224,N_22580);
nand U29323 (N_29323,N_21727,N_20225);
nor U29324 (N_29324,N_22584,N_22500);
nand U29325 (N_29325,N_22617,N_20638);
nor U29326 (N_29326,N_23611,N_20017);
nand U29327 (N_29327,N_21109,N_20568);
xor U29328 (N_29328,N_21406,N_21706);
xor U29329 (N_29329,N_24318,N_23043);
xnor U29330 (N_29330,N_20743,N_21105);
and U29331 (N_29331,N_24221,N_21112);
nor U29332 (N_29332,N_23802,N_24029);
nor U29333 (N_29333,N_24016,N_24951);
nand U29334 (N_29334,N_22569,N_22549);
and U29335 (N_29335,N_23047,N_21654);
nand U29336 (N_29336,N_20362,N_23020);
or U29337 (N_29337,N_22823,N_22890);
nor U29338 (N_29338,N_20668,N_20482);
nand U29339 (N_29339,N_24599,N_24273);
nor U29340 (N_29340,N_23364,N_23481);
or U29341 (N_29341,N_23744,N_24195);
or U29342 (N_29342,N_23969,N_22258);
or U29343 (N_29343,N_21130,N_24808);
nand U29344 (N_29344,N_22820,N_22853);
nor U29345 (N_29345,N_20047,N_22912);
nand U29346 (N_29346,N_23092,N_20403);
or U29347 (N_29347,N_23935,N_23258);
or U29348 (N_29348,N_24861,N_20296);
xor U29349 (N_29349,N_21770,N_22196);
nor U29350 (N_29350,N_22063,N_23576);
nor U29351 (N_29351,N_24371,N_22313);
or U29352 (N_29352,N_23561,N_22934);
nor U29353 (N_29353,N_20087,N_22798);
nand U29354 (N_29354,N_22086,N_24742);
nor U29355 (N_29355,N_23767,N_22639);
and U29356 (N_29356,N_23780,N_24746);
or U29357 (N_29357,N_24855,N_24212);
nand U29358 (N_29358,N_24392,N_24626);
nand U29359 (N_29359,N_22847,N_22599);
nand U29360 (N_29360,N_22146,N_22510);
or U29361 (N_29361,N_23302,N_22486);
or U29362 (N_29362,N_22214,N_22965);
nand U29363 (N_29363,N_20680,N_24893);
nor U29364 (N_29364,N_22800,N_20399);
nor U29365 (N_29365,N_24762,N_22663);
and U29366 (N_29366,N_23695,N_20555);
and U29367 (N_29367,N_20069,N_20784);
xnor U29368 (N_29368,N_23684,N_23268);
xor U29369 (N_29369,N_21422,N_24468);
xnor U29370 (N_29370,N_22570,N_22923);
or U29371 (N_29371,N_20057,N_21480);
xnor U29372 (N_29372,N_22383,N_21885);
nor U29373 (N_29373,N_21829,N_22637);
nand U29374 (N_29374,N_21533,N_23109);
and U29375 (N_29375,N_23361,N_24067);
and U29376 (N_29376,N_22674,N_22455);
or U29377 (N_29377,N_21404,N_22385);
or U29378 (N_29378,N_22409,N_23598);
or U29379 (N_29379,N_24815,N_24196);
nand U29380 (N_29380,N_24243,N_23188);
or U29381 (N_29381,N_24683,N_24151);
xor U29382 (N_29382,N_22285,N_22522);
and U29383 (N_29383,N_23786,N_24018);
and U29384 (N_29384,N_21123,N_22565);
and U29385 (N_29385,N_22930,N_24922);
xnor U29386 (N_29386,N_23731,N_23309);
nor U29387 (N_29387,N_23067,N_21690);
nor U29388 (N_29388,N_21470,N_24897);
xor U29389 (N_29389,N_24974,N_24539);
or U29390 (N_29390,N_20627,N_20377);
and U29391 (N_29391,N_24016,N_20922);
and U29392 (N_29392,N_20256,N_24099);
or U29393 (N_29393,N_20201,N_21032);
or U29394 (N_29394,N_23541,N_24723);
xnor U29395 (N_29395,N_23398,N_21634);
nor U29396 (N_29396,N_20673,N_24088);
or U29397 (N_29397,N_20591,N_23108);
or U29398 (N_29398,N_23227,N_21055);
nand U29399 (N_29399,N_21383,N_22646);
nor U29400 (N_29400,N_22140,N_23236);
or U29401 (N_29401,N_22396,N_24146);
or U29402 (N_29402,N_20167,N_23229);
nand U29403 (N_29403,N_21399,N_21503);
or U29404 (N_29404,N_24335,N_21895);
nor U29405 (N_29405,N_22238,N_24839);
nand U29406 (N_29406,N_20609,N_24673);
nor U29407 (N_29407,N_24706,N_20683);
nor U29408 (N_29408,N_22564,N_23419);
nand U29409 (N_29409,N_21679,N_24327);
nand U29410 (N_29410,N_24443,N_24133);
nor U29411 (N_29411,N_22624,N_20165);
and U29412 (N_29412,N_21259,N_21436);
and U29413 (N_29413,N_20682,N_22121);
and U29414 (N_29414,N_23043,N_24750);
and U29415 (N_29415,N_24011,N_24353);
xor U29416 (N_29416,N_22554,N_22237);
nand U29417 (N_29417,N_23916,N_22311);
or U29418 (N_29418,N_24102,N_21619);
nand U29419 (N_29419,N_24052,N_20851);
xor U29420 (N_29420,N_20942,N_22913);
nand U29421 (N_29421,N_20084,N_23155);
and U29422 (N_29422,N_21542,N_21034);
nor U29423 (N_29423,N_24653,N_21199);
or U29424 (N_29424,N_24398,N_22775);
nor U29425 (N_29425,N_22308,N_24430);
nand U29426 (N_29426,N_21381,N_20887);
nand U29427 (N_29427,N_24696,N_20586);
xnor U29428 (N_29428,N_24710,N_22330);
and U29429 (N_29429,N_22064,N_23360);
nand U29430 (N_29430,N_22185,N_20666);
and U29431 (N_29431,N_23888,N_23875);
or U29432 (N_29432,N_21323,N_21924);
nor U29433 (N_29433,N_23960,N_24602);
nor U29434 (N_29434,N_20112,N_20016);
nand U29435 (N_29435,N_20673,N_21603);
or U29436 (N_29436,N_20578,N_20118);
xor U29437 (N_29437,N_22063,N_20549);
and U29438 (N_29438,N_23391,N_23232);
and U29439 (N_29439,N_21339,N_23819);
nor U29440 (N_29440,N_23348,N_22483);
or U29441 (N_29441,N_22050,N_22805);
nand U29442 (N_29442,N_22148,N_24628);
nand U29443 (N_29443,N_21880,N_23232);
nor U29444 (N_29444,N_24451,N_22557);
or U29445 (N_29445,N_21255,N_24912);
nor U29446 (N_29446,N_23932,N_24118);
or U29447 (N_29447,N_24252,N_24298);
xor U29448 (N_29448,N_22073,N_24397);
and U29449 (N_29449,N_21669,N_20315);
or U29450 (N_29450,N_23111,N_20801);
or U29451 (N_29451,N_21614,N_22724);
or U29452 (N_29452,N_21600,N_21678);
nand U29453 (N_29453,N_21525,N_22032);
nor U29454 (N_29454,N_22018,N_22671);
or U29455 (N_29455,N_22474,N_20588);
nand U29456 (N_29456,N_21346,N_20832);
nor U29457 (N_29457,N_23922,N_24239);
xnor U29458 (N_29458,N_24665,N_21086);
xnor U29459 (N_29459,N_20879,N_21290);
nand U29460 (N_29460,N_21393,N_20875);
nor U29461 (N_29461,N_22902,N_23529);
and U29462 (N_29462,N_22900,N_24276);
or U29463 (N_29463,N_22162,N_24444);
and U29464 (N_29464,N_22180,N_21932);
nor U29465 (N_29465,N_21188,N_21072);
nor U29466 (N_29466,N_22678,N_21851);
nor U29467 (N_29467,N_23599,N_20901);
nand U29468 (N_29468,N_23237,N_23769);
or U29469 (N_29469,N_22607,N_21882);
or U29470 (N_29470,N_20376,N_22463);
nor U29471 (N_29471,N_22982,N_24306);
nand U29472 (N_29472,N_20801,N_21034);
nor U29473 (N_29473,N_22855,N_22468);
or U29474 (N_29474,N_20002,N_22119);
nand U29475 (N_29475,N_21928,N_22576);
or U29476 (N_29476,N_22456,N_23246);
nand U29477 (N_29477,N_23409,N_22109);
or U29478 (N_29478,N_22996,N_23588);
nand U29479 (N_29479,N_21581,N_23454);
nand U29480 (N_29480,N_24981,N_20304);
or U29481 (N_29481,N_21110,N_22175);
nand U29482 (N_29482,N_21870,N_23159);
nand U29483 (N_29483,N_21936,N_24977);
nand U29484 (N_29484,N_23214,N_20692);
xor U29485 (N_29485,N_20232,N_23387);
nor U29486 (N_29486,N_22872,N_24616);
or U29487 (N_29487,N_23648,N_21199);
and U29488 (N_29488,N_20069,N_22700);
and U29489 (N_29489,N_24565,N_23069);
or U29490 (N_29490,N_23166,N_23738);
nand U29491 (N_29491,N_21309,N_21365);
nand U29492 (N_29492,N_23019,N_23619);
and U29493 (N_29493,N_23615,N_23675);
or U29494 (N_29494,N_23293,N_22423);
nand U29495 (N_29495,N_22781,N_23098);
nor U29496 (N_29496,N_22173,N_23915);
or U29497 (N_29497,N_23953,N_23128);
or U29498 (N_29498,N_24232,N_23067);
and U29499 (N_29499,N_20072,N_24316);
and U29500 (N_29500,N_21462,N_23813);
nand U29501 (N_29501,N_22358,N_23893);
nor U29502 (N_29502,N_24076,N_22182);
nor U29503 (N_29503,N_22185,N_23766);
nand U29504 (N_29504,N_21434,N_20354);
nand U29505 (N_29505,N_23374,N_20287);
or U29506 (N_29506,N_24255,N_20918);
nor U29507 (N_29507,N_23106,N_21823);
or U29508 (N_29508,N_20669,N_20149);
and U29509 (N_29509,N_22173,N_23664);
and U29510 (N_29510,N_21021,N_23199);
or U29511 (N_29511,N_23210,N_21807);
and U29512 (N_29512,N_24383,N_21825);
xor U29513 (N_29513,N_22980,N_24972);
and U29514 (N_29514,N_22116,N_23389);
nand U29515 (N_29515,N_20027,N_22299);
nor U29516 (N_29516,N_22880,N_23723);
xnor U29517 (N_29517,N_21752,N_23341);
and U29518 (N_29518,N_22171,N_20972);
and U29519 (N_29519,N_22339,N_23086);
or U29520 (N_29520,N_24813,N_20041);
nand U29521 (N_29521,N_23497,N_24845);
or U29522 (N_29522,N_22657,N_22913);
and U29523 (N_29523,N_21231,N_21456);
or U29524 (N_29524,N_23100,N_21081);
nor U29525 (N_29525,N_24629,N_23107);
xnor U29526 (N_29526,N_21789,N_24037);
xnor U29527 (N_29527,N_22936,N_21347);
nor U29528 (N_29528,N_20219,N_24803);
and U29529 (N_29529,N_22018,N_20591);
nand U29530 (N_29530,N_24411,N_23233);
nand U29531 (N_29531,N_21864,N_20652);
or U29532 (N_29532,N_22109,N_24747);
nor U29533 (N_29533,N_21149,N_20230);
or U29534 (N_29534,N_21832,N_21985);
or U29535 (N_29535,N_24578,N_20284);
and U29536 (N_29536,N_23780,N_20925);
or U29537 (N_29537,N_22375,N_24174);
nor U29538 (N_29538,N_21861,N_23374);
and U29539 (N_29539,N_20221,N_24497);
nand U29540 (N_29540,N_24606,N_24532);
nor U29541 (N_29541,N_21685,N_22024);
nand U29542 (N_29542,N_21571,N_22352);
nor U29543 (N_29543,N_22055,N_22970);
and U29544 (N_29544,N_23935,N_22114);
nand U29545 (N_29545,N_21685,N_20926);
nor U29546 (N_29546,N_22882,N_23450);
or U29547 (N_29547,N_21097,N_22678);
or U29548 (N_29548,N_20660,N_20863);
nor U29549 (N_29549,N_20106,N_24381);
or U29550 (N_29550,N_22275,N_24438);
nand U29551 (N_29551,N_23424,N_23004);
and U29552 (N_29552,N_24307,N_21654);
nor U29553 (N_29553,N_20291,N_20668);
or U29554 (N_29554,N_20786,N_20911);
and U29555 (N_29555,N_22121,N_22941);
nand U29556 (N_29556,N_23187,N_20681);
nor U29557 (N_29557,N_23084,N_24146);
and U29558 (N_29558,N_21868,N_22880);
nand U29559 (N_29559,N_23159,N_21610);
nor U29560 (N_29560,N_20538,N_21628);
xnor U29561 (N_29561,N_24209,N_20429);
nor U29562 (N_29562,N_21997,N_23103);
and U29563 (N_29563,N_23803,N_22738);
or U29564 (N_29564,N_24210,N_21922);
nor U29565 (N_29565,N_24112,N_22492);
or U29566 (N_29566,N_20929,N_22760);
and U29567 (N_29567,N_24432,N_24927);
nor U29568 (N_29568,N_24422,N_23773);
nand U29569 (N_29569,N_21061,N_23372);
nand U29570 (N_29570,N_20034,N_22558);
and U29571 (N_29571,N_23916,N_22593);
nor U29572 (N_29572,N_23489,N_23243);
nor U29573 (N_29573,N_22893,N_24604);
nand U29574 (N_29574,N_20575,N_23017);
nor U29575 (N_29575,N_23697,N_23601);
and U29576 (N_29576,N_22332,N_24774);
and U29577 (N_29577,N_24439,N_21300);
nor U29578 (N_29578,N_23558,N_22187);
nand U29579 (N_29579,N_24675,N_24413);
nor U29580 (N_29580,N_23909,N_22686);
and U29581 (N_29581,N_23306,N_20063);
nand U29582 (N_29582,N_21225,N_21327);
and U29583 (N_29583,N_20480,N_23567);
or U29584 (N_29584,N_24983,N_21064);
nand U29585 (N_29585,N_24655,N_21441);
or U29586 (N_29586,N_22868,N_21418);
or U29587 (N_29587,N_21357,N_21633);
nor U29588 (N_29588,N_20510,N_23803);
xnor U29589 (N_29589,N_21934,N_20733);
xor U29590 (N_29590,N_23073,N_20869);
or U29591 (N_29591,N_23065,N_22516);
or U29592 (N_29592,N_20184,N_23101);
xnor U29593 (N_29593,N_24079,N_22161);
or U29594 (N_29594,N_21959,N_23815);
and U29595 (N_29595,N_22525,N_22709);
nor U29596 (N_29596,N_22856,N_21335);
nor U29597 (N_29597,N_23960,N_20010);
nor U29598 (N_29598,N_23281,N_22554);
nand U29599 (N_29599,N_24157,N_22181);
nor U29600 (N_29600,N_24806,N_21948);
or U29601 (N_29601,N_22245,N_21792);
nand U29602 (N_29602,N_21362,N_21058);
nand U29603 (N_29603,N_23063,N_21363);
nand U29604 (N_29604,N_23299,N_24699);
nor U29605 (N_29605,N_22889,N_24138);
or U29606 (N_29606,N_23465,N_21120);
nor U29607 (N_29607,N_21170,N_21463);
nand U29608 (N_29608,N_20387,N_23433);
nor U29609 (N_29609,N_23345,N_23443);
xor U29610 (N_29610,N_24814,N_24941);
xnor U29611 (N_29611,N_22645,N_20535);
nand U29612 (N_29612,N_20470,N_24744);
xor U29613 (N_29613,N_23319,N_21991);
or U29614 (N_29614,N_21823,N_23695);
and U29615 (N_29615,N_23133,N_21134);
nor U29616 (N_29616,N_20958,N_20316);
nand U29617 (N_29617,N_22394,N_24963);
nor U29618 (N_29618,N_23337,N_21367);
and U29619 (N_29619,N_20147,N_23132);
and U29620 (N_29620,N_20832,N_23737);
nor U29621 (N_29621,N_20831,N_24190);
or U29622 (N_29622,N_24828,N_22692);
and U29623 (N_29623,N_24437,N_22725);
xnor U29624 (N_29624,N_24676,N_21876);
xnor U29625 (N_29625,N_21845,N_22606);
nand U29626 (N_29626,N_20375,N_22333);
and U29627 (N_29627,N_20777,N_24726);
nor U29628 (N_29628,N_23077,N_22648);
or U29629 (N_29629,N_24576,N_24382);
and U29630 (N_29630,N_21190,N_20563);
and U29631 (N_29631,N_20025,N_23775);
and U29632 (N_29632,N_24231,N_20169);
or U29633 (N_29633,N_21691,N_23377);
xnor U29634 (N_29634,N_23861,N_22528);
nor U29635 (N_29635,N_23392,N_20199);
or U29636 (N_29636,N_23714,N_22583);
nand U29637 (N_29637,N_22743,N_22225);
nor U29638 (N_29638,N_23394,N_22767);
and U29639 (N_29639,N_24106,N_20926);
and U29640 (N_29640,N_23395,N_20946);
nand U29641 (N_29641,N_23118,N_24269);
nor U29642 (N_29642,N_21834,N_21000);
and U29643 (N_29643,N_24943,N_20588);
and U29644 (N_29644,N_20087,N_24401);
or U29645 (N_29645,N_21007,N_23118);
nand U29646 (N_29646,N_21455,N_21262);
nor U29647 (N_29647,N_21703,N_20269);
nor U29648 (N_29648,N_23474,N_22681);
xor U29649 (N_29649,N_21249,N_22708);
and U29650 (N_29650,N_23997,N_23017);
xor U29651 (N_29651,N_23914,N_22050);
and U29652 (N_29652,N_22182,N_20987);
nand U29653 (N_29653,N_23669,N_24170);
and U29654 (N_29654,N_21142,N_24029);
xor U29655 (N_29655,N_20167,N_20865);
nand U29656 (N_29656,N_22233,N_21874);
xnor U29657 (N_29657,N_22237,N_21683);
and U29658 (N_29658,N_22006,N_21222);
nand U29659 (N_29659,N_20221,N_20934);
nor U29660 (N_29660,N_22728,N_21130);
and U29661 (N_29661,N_22033,N_24902);
nor U29662 (N_29662,N_20101,N_24787);
nand U29663 (N_29663,N_22759,N_20341);
nand U29664 (N_29664,N_23649,N_23840);
and U29665 (N_29665,N_23179,N_24128);
xnor U29666 (N_29666,N_22001,N_22067);
or U29667 (N_29667,N_23091,N_23316);
or U29668 (N_29668,N_24889,N_22560);
or U29669 (N_29669,N_22696,N_21047);
and U29670 (N_29670,N_23586,N_21372);
and U29671 (N_29671,N_21702,N_22268);
and U29672 (N_29672,N_21332,N_24327);
and U29673 (N_29673,N_23572,N_23311);
or U29674 (N_29674,N_20158,N_20479);
and U29675 (N_29675,N_23431,N_24652);
xor U29676 (N_29676,N_20840,N_21190);
nand U29677 (N_29677,N_22934,N_24403);
and U29678 (N_29678,N_23111,N_20983);
and U29679 (N_29679,N_24301,N_20719);
xnor U29680 (N_29680,N_24083,N_23025);
nor U29681 (N_29681,N_24200,N_24248);
nand U29682 (N_29682,N_23216,N_21708);
and U29683 (N_29683,N_21237,N_23698);
nand U29684 (N_29684,N_21843,N_20881);
nand U29685 (N_29685,N_23720,N_21507);
xor U29686 (N_29686,N_23050,N_24546);
nand U29687 (N_29687,N_24960,N_24736);
nand U29688 (N_29688,N_20469,N_22823);
nor U29689 (N_29689,N_20307,N_20364);
and U29690 (N_29690,N_24478,N_21886);
xor U29691 (N_29691,N_20272,N_20251);
nor U29692 (N_29692,N_24547,N_23467);
and U29693 (N_29693,N_24958,N_20947);
nand U29694 (N_29694,N_24595,N_24616);
or U29695 (N_29695,N_22413,N_20228);
nor U29696 (N_29696,N_20529,N_21019);
nand U29697 (N_29697,N_23958,N_20696);
xor U29698 (N_29698,N_22170,N_24467);
and U29699 (N_29699,N_24391,N_24123);
or U29700 (N_29700,N_24378,N_23526);
and U29701 (N_29701,N_23054,N_24119);
nand U29702 (N_29702,N_24353,N_22569);
and U29703 (N_29703,N_24144,N_24155);
or U29704 (N_29704,N_22304,N_21141);
or U29705 (N_29705,N_20467,N_21982);
nand U29706 (N_29706,N_24826,N_21196);
nor U29707 (N_29707,N_22674,N_21913);
or U29708 (N_29708,N_23195,N_23217);
and U29709 (N_29709,N_21948,N_24398);
or U29710 (N_29710,N_23960,N_21426);
or U29711 (N_29711,N_22832,N_24913);
or U29712 (N_29712,N_22043,N_20679);
xor U29713 (N_29713,N_24596,N_23552);
nand U29714 (N_29714,N_21052,N_20559);
nor U29715 (N_29715,N_20004,N_20957);
nand U29716 (N_29716,N_21000,N_21385);
and U29717 (N_29717,N_21582,N_20745);
nor U29718 (N_29718,N_24089,N_22041);
and U29719 (N_29719,N_21960,N_23613);
and U29720 (N_29720,N_22495,N_22205);
nand U29721 (N_29721,N_23928,N_22130);
nor U29722 (N_29722,N_21030,N_21271);
or U29723 (N_29723,N_24180,N_22419);
or U29724 (N_29724,N_23913,N_21153);
or U29725 (N_29725,N_22536,N_20846);
xor U29726 (N_29726,N_24382,N_20004);
and U29727 (N_29727,N_23548,N_20007);
nand U29728 (N_29728,N_20060,N_23988);
nand U29729 (N_29729,N_20948,N_20926);
or U29730 (N_29730,N_24390,N_21995);
or U29731 (N_29731,N_20199,N_20842);
nand U29732 (N_29732,N_24214,N_24953);
or U29733 (N_29733,N_20484,N_24598);
nor U29734 (N_29734,N_20787,N_23458);
or U29735 (N_29735,N_21959,N_24342);
and U29736 (N_29736,N_20836,N_22639);
xnor U29737 (N_29737,N_24349,N_21578);
nand U29738 (N_29738,N_21919,N_20511);
and U29739 (N_29739,N_21790,N_22995);
nand U29740 (N_29740,N_22231,N_20740);
nand U29741 (N_29741,N_24522,N_21223);
xor U29742 (N_29742,N_22476,N_24350);
or U29743 (N_29743,N_21174,N_20450);
nand U29744 (N_29744,N_21101,N_22176);
and U29745 (N_29745,N_24414,N_23384);
nand U29746 (N_29746,N_22666,N_24440);
and U29747 (N_29747,N_24492,N_23106);
xnor U29748 (N_29748,N_21545,N_22533);
nor U29749 (N_29749,N_21209,N_21736);
and U29750 (N_29750,N_24713,N_22816);
nor U29751 (N_29751,N_23375,N_21293);
xnor U29752 (N_29752,N_21075,N_24381);
or U29753 (N_29753,N_20653,N_22712);
nand U29754 (N_29754,N_23292,N_22035);
nand U29755 (N_29755,N_24422,N_23497);
and U29756 (N_29756,N_21228,N_24310);
or U29757 (N_29757,N_21262,N_22575);
nand U29758 (N_29758,N_22190,N_23534);
nor U29759 (N_29759,N_20690,N_20902);
nor U29760 (N_29760,N_23096,N_20869);
xor U29761 (N_29761,N_23601,N_24481);
nor U29762 (N_29762,N_20642,N_22696);
nand U29763 (N_29763,N_21170,N_23413);
or U29764 (N_29764,N_24178,N_21205);
xnor U29765 (N_29765,N_21883,N_24382);
nor U29766 (N_29766,N_23313,N_22006);
nand U29767 (N_29767,N_24950,N_24400);
nor U29768 (N_29768,N_23898,N_21521);
nor U29769 (N_29769,N_20021,N_23614);
xor U29770 (N_29770,N_21527,N_22440);
nand U29771 (N_29771,N_23211,N_21206);
nor U29772 (N_29772,N_20152,N_23787);
xnor U29773 (N_29773,N_20788,N_21838);
nor U29774 (N_29774,N_23308,N_21110);
nand U29775 (N_29775,N_21426,N_24606);
or U29776 (N_29776,N_22990,N_23734);
nor U29777 (N_29777,N_22427,N_23968);
nor U29778 (N_29778,N_23038,N_20278);
or U29779 (N_29779,N_21496,N_20388);
and U29780 (N_29780,N_21027,N_20007);
nor U29781 (N_29781,N_23954,N_20071);
and U29782 (N_29782,N_22815,N_21859);
nor U29783 (N_29783,N_23297,N_20396);
nand U29784 (N_29784,N_23884,N_21077);
nor U29785 (N_29785,N_22143,N_24743);
and U29786 (N_29786,N_24421,N_20677);
nand U29787 (N_29787,N_21172,N_23291);
and U29788 (N_29788,N_22495,N_24349);
nand U29789 (N_29789,N_22158,N_22485);
nand U29790 (N_29790,N_23603,N_21236);
nor U29791 (N_29791,N_21639,N_20013);
nand U29792 (N_29792,N_22073,N_23291);
nand U29793 (N_29793,N_23727,N_21778);
and U29794 (N_29794,N_23285,N_24849);
and U29795 (N_29795,N_20971,N_24047);
nand U29796 (N_29796,N_21234,N_23605);
or U29797 (N_29797,N_22393,N_21685);
and U29798 (N_29798,N_21508,N_22085);
xnor U29799 (N_29799,N_24270,N_23361);
and U29800 (N_29800,N_20150,N_22663);
or U29801 (N_29801,N_22524,N_22159);
nor U29802 (N_29802,N_23479,N_21161);
nor U29803 (N_29803,N_20216,N_22903);
or U29804 (N_29804,N_22433,N_24870);
or U29805 (N_29805,N_22970,N_21881);
nand U29806 (N_29806,N_23942,N_22623);
xnor U29807 (N_29807,N_24734,N_23904);
nand U29808 (N_29808,N_20275,N_24832);
nor U29809 (N_29809,N_21333,N_24908);
nand U29810 (N_29810,N_22770,N_23458);
nand U29811 (N_29811,N_22326,N_21920);
nand U29812 (N_29812,N_23756,N_22086);
nor U29813 (N_29813,N_24946,N_21151);
nand U29814 (N_29814,N_24451,N_21727);
and U29815 (N_29815,N_20347,N_20894);
nor U29816 (N_29816,N_22627,N_22660);
nor U29817 (N_29817,N_24385,N_24981);
and U29818 (N_29818,N_20741,N_22345);
nand U29819 (N_29819,N_22193,N_21566);
and U29820 (N_29820,N_20873,N_22673);
nor U29821 (N_29821,N_21367,N_22840);
or U29822 (N_29822,N_23902,N_23266);
or U29823 (N_29823,N_24585,N_24202);
and U29824 (N_29824,N_22301,N_20518);
and U29825 (N_29825,N_22904,N_22591);
nor U29826 (N_29826,N_21026,N_23760);
nand U29827 (N_29827,N_23341,N_24254);
nand U29828 (N_29828,N_22423,N_22521);
xor U29829 (N_29829,N_23851,N_20630);
and U29830 (N_29830,N_22972,N_20758);
or U29831 (N_29831,N_20776,N_21207);
and U29832 (N_29832,N_23967,N_21820);
or U29833 (N_29833,N_22563,N_22308);
nand U29834 (N_29834,N_20921,N_23964);
and U29835 (N_29835,N_20711,N_20404);
or U29836 (N_29836,N_22837,N_20660);
and U29837 (N_29837,N_20369,N_22036);
nor U29838 (N_29838,N_20110,N_20439);
nand U29839 (N_29839,N_21016,N_22803);
or U29840 (N_29840,N_24363,N_24059);
nand U29841 (N_29841,N_24227,N_22867);
or U29842 (N_29842,N_24484,N_24654);
nand U29843 (N_29843,N_20427,N_21084);
or U29844 (N_29844,N_21538,N_24236);
xor U29845 (N_29845,N_23111,N_23075);
xor U29846 (N_29846,N_22303,N_21542);
nor U29847 (N_29847,N_20589,N_24823);
nand U29848 (N_29848,N_21692,N_22959);
or U29849 (N_29849,N_22615,N_24439);
or U29850 (N_29850,N_24661,N_22253);
nand U29851 (N_29851,N_22340,N_22548);
and U29852 (N_29852,N_22603,N_21218);
or U29853 (N_29853,N_24169,N_23917);
and U29854 (N_29854,N_24989,N_23725);
or U29855 (N_29855,N_20170,N_23671);
or U29856 (N_29856,N_23369,N_23741);
xnor U29857 (N_29857,N_23571,N_22902);
nand U29858 (N_29858,N_22056,N_23203);
nor U29859 (N_29859,N_23512,N_21653);
nand U29860 (N_29860,N_23812,N_21885);
nor U29861 (N_29861,N_20046,N_24722);
nor U29862 (N_29862,N_20096,N_22136);
xor U29863 (N_29863,N_24631,N_20506);
nor U29864 (N_29864,N_20602,N_20825);
or U29865 (N_29865,N_22440,N_24201);
xnor U29866 (N_29866,N_22856,N_21556);
xor U29867 (N_29867,N_20050,N_22204);
or U29868 (N_29868,N_20692,N_24676);
nand U29869 (N_29869,N_23684,N_24738);
or U29870 (N_29870,N_20150,N_22023);
nand U29871 (N_29871,N_22905,N_23746);
nand U29872 (N_29872,N_24440,N_24038);
nor U29873 (N_29873,N_20876,N_22064);
and U29874 (N_29874,N_23179,N_22815);
or U29875 (N_29875,N_20390,N_21939);
xor U29876 (N_29876,N_22259,N_23265);
xor U29877 (N_29877,N_24402,N_22848);
nand U29878 (N_29878,N_20809,N_20565);
or U29879 (N_29879,N_22393,N_23063);
nand U29880 (N_29880,N_22263,N_24038);
or U29881 (N_29881,N_22576,N_24522);
nand U29882 (N_29882,N_23093,N_21489);
and U29883 (N_29883,N_22470,N_24380);
xor U29884 (N_29884,N_24431,N_22007);
nor U29885 (N_29885,N_20937,N_20084);
nor U29886 (N_29886,N_20972,N_22325);
nor U29887 (N_29887,N_20862,N_23516);
xnor U29888 (N_29888,N_24938,N_21234);
nor U29889 (N_29889,N_24364,N_23861);
nand U29890 (N_29890,N_22735,N_22997);
or U29891 (N_29891,N_21496,N_20320);
nand U29892 (N_29892,N_22056,N_22862);
and U29893 (N_29893,N_22477,N_20936);
or U29894 (N_29894,N_20693,N_24933);
nand U29895 (N_29895,N_22287,N_22286);
xnor U29896 (N_29896,N_23411,N_21530);
nand U29897 (N_29897,N_21929,N_21786);
or U29898 (N_29898,N_23110,N_22834);
or U29899 (N_29899,N_20050,N_21355);
nor U29900 (N_29900,N_23265,N_21898);
and U29901 (N_29901,N_21364,N_21399);
nand U29902 (N_29902,N_22737,N_20682);
nand U29903 (N_29903,N_23354,N_23275);
xor U29904 (N_29904,N_23437,N_23321);
and U29905 (N_29905,N_21103,N_20703);
xnor U29906 (N_29906,N_23178,N_24454);
nand U29907 (N_29907,N_21359,N_22074);
xor U29908 (N_29908,N_24902,N_22647);
nand U29909 (N_29909,N_22076,N_20303);
or U29910 (N_29910,N_24963,N_22183);
or U29911 (N_29911,N_24715,N_21664);
nor U29912 (N_29912,N_24458,N_20243);
or U29913 (N_29913,N_20919,N_22687);
or U29914 (N_29914,N_24657,N_22460);
or U29915 (N_29915,N_21562,N_23936);
nor U29916 (N_29916,N_23640,N_22093);
and U29917 (N_29917,N_24402,N_23195);
and U29918 (N_29918,N_21899,N_24617);
and U29919 (N_29919,N_22162,N_22274);
nand U29920 (N_29920,N_21379,N_24961);
or U29921 (N_29921,N_21230,N_21374);
and U29922 (N_29922,N_24609,N_20390);
nor U29923 (N_29923,N_20754,N_21232);
nand U29924 (N_29924,N_22980,N_23122);
nand U29925 (N_29925,N_21360,N_21627);
or U29926 (N_29926,N_22368,N_20140);
or U29927 (N_29927,N_21181,N_22564);
and U29928 (N_29928,N_20520,N_22678);
xnor U29929 (N_29929,N_20716,N_22213);
xnor U29930 (N_29930,N_22893,N_23184);
and U29931 (N_29931,N_24212,N_20977);
and U29932 (N_29932,N_24044,N_24826);
nor U29933 (N_29933,N_23086,N_23357);
or U29934 (N_29934,N_23072,N_21506);
or U29935 (N_29935,N_23904,N_23685);
and U29936 (N_29936,N_20032,N_21121);
or U29937 (N_29937,N_20490,N_20090);
and U29938 (N_29938,N_20072,N_21158);
xor U29939 (N_29939,N_22328,N_24479);
or U29940 (N_29940,N_24581,N_20392);
and U29941 (N_29941,N_24849,N_24304);
and U29942 (N_29942,N_22419,N_20754);
or U29943 (N_29943,N_21672,N_21837);
or U29944 (N_29944,N_21409,N_24768);
or U29945 (N_29945,N_23213,N_23001);
or U29946 (N_29946,N_22396,N_20655);
xor U29947 (N_29947,N_22751,N_24204);
nand U29948 (N_29948,N_21437,N_22527);
xor U29949 (N_29949,N_24825,N_20839);
nor U29950 (N_29950,N_22461,N_20272);
nor U29951 (N_29951,N_22872,N_23029);
and U29952 (N_29952,N_20423,N_20519);
xnor U29953 (N_29953,N_20951,N_21209);
nand U29954 (N_29954,N_23827,N_21141);
xor U29955 (N_29955,N_23796,N_21858);
or U29956 (N_29956,N_24869,N_20163);
and U29957 (N_29957,N_20217,N_23604);
and U29958 (N_29958,N_22560,N_20758);
nor U29959 (N_29959,N_20035,N_20741);
nor U29960 (N_29960,N_20005,N_23238);
and U29961 (N_29961,N_21164,N_21235);
and U29962 (N_29962,N_24654,N_22445);
xnor U29963 (N_29963,N_22953,N_23021);
or U29964 (N_29964,N_24868,N_23168);
and U29965 (N_29965,N_22990,N_24043);
or U29966 (N_29966,N_20712,N_20714);
or U29967 (N_29967,N_23606,N_22702);
or U29968 (N_29968,N_21839,N_20967);
or U29969 (N_29969,N_23462,N_23240);
nor U29970 (N_29970,N_23626,N_24728);
nand U29971 (N_29971,N_24020,N_22259);
and U29972 (N_29972,N_24896,N_23333);
nor U29973 (N_29973,N_22255,N_20078);
nand U29974 (N_29974,N_21497,N_24681);
nor U29975 (N_29975,N_21306,N_21181);
nor U29976 (N_29976,N_21201,N_20509);
and U29977 (N_29977,N_23593,N_24440);
nor U29978 (N_29978,N_20206,N_23747);
or U29979 (N_29979,N_23599,N_21755);
or U29980 (N_29980,N_20556,N_24796);
and U29981 (N_29981,N_23095,N_21783);
xnor U29982 (N_29982,N_23325,N_23238);
nand U29983 (N_29983,N_23543,N_21033);
nand U29984 (N_29984,N_22073,N_24264);
nand U29985 (N_29985,N_22941,N_24466);
or U29986 (N_29986,N_24096,N_21862);
nand U29987 (N_29987,N_24660,N_24915);
and U29988 (N_29988,N_24462,N_23154);
or U29989 (N_29989,N_24619,N_22294);
xnor U29990 (N_29990,N_23651,N_24692);
or U29991 (N_29991,N_24670,N_24654);
nand U29992 (N_29992,N_24211,N_21709);
or U29993 (N_29993,N_22505,N_24875);
nor U29994 (N_29994,N_21516,N_22675);
or U29995 (N_29995,N_21166,N_22225);
and U29996 (N_29996,N_21294,N_20293);
nor U29997 (N_29997,N_22040,N_20376);
nor U29998 (N_29998,N_24183,N_22131);
or U29999 (N_29999,N_21644,N_20262);
nor UO_0 (O_0,N_27577,N_29152);
or UO_1 (O_1,N_25140,N_29427);
or UO_2 (O_2,N_25498,N_28790);
nand UO_3 (O_3,N_26307,N_29860);
or UO_4 (O_4,N_28822,N_28947);
or UO_5 (O_5,N_28967,N_28220);
nand UO_6 (O_6,N_29561,N_26740);
and UO_7 (O_7,N_27456,N_25733);
and UO_8 (O_8,N_28875,N_26277);
and UO_9 (O_9,N_27295,N_25470);
nor UO_10 (O_10,N_25037,N_26578);
nor UO_11 (O_11,N_29522,N_27882);
or UO_12 (O_12,N_26021,N_25615);
or UO_13 (O_13,N_25387,N_25755);
nand UO_14 (O_14,N_29090,N_29096);
xor UO_15 (O_15,N_27662,N_29308);
nor UO_16 (O_16,N_28903,N_27602);
and UO_17 (O_17,N_28463,N_26311);
nand UO_18 (O_18,N_28593,N_25801);
and UO_19 (O_19,N_28548,N_28631);
or UO_20 (O_20,N_26859,N_28510);
xnor UO_21 (O_21,N_26582,N_29932);
and UO_22 (O_22,N_28478,N_26677);
xnor UO_23 (O_23,N_26264,N_25393);
nor UO_24 (O_24,N_27192,N_28295);
and UO_25 (O_25,N_29099,N_25036);
and UO_26 (O_26,N_27770,N_27055);
nand UO_27 (O_27,N_26174,N_25463);
nor UO_28 (O_28,N_27816,N_29844);
xnor UO_29 (O_29,N_25886,N_27496);
xor UO_30 (O_30,N_28171,N_25850);
and UO_31 (O_31,N_29148,N_25233);
nand UO_32 (O_32,N_27961,N_25218);
nor UO_33 (O_33,N_25374,N_27125);
nor UO_34 (O_34,N_26825,N_27629);
and UO_35 (O_35,N_27255,N_28092);
or UO_36 (O_36,N_29451,N_27252);
nor UO_37 (O_37,N_29618,N_28433);
and UO_38 (O_38,N_28994,N_26798);
xnor UO_39 (O_39,N_28412,N_29394);
nor UO_40 (O_40,N_26478,N_29219);
or UO_41 (O_41,N_26010,N_29486);
and UO_42 (O_42,N_26160,N_28824);
nor UO_43 (O_43,N_26569,N_26351);
nor UO_44 (O_44,N_27635,N_25605);
and UO_45 (O_45,N_25416,N_26992);
or UO_46 (O_46,N_27665,N_27915);
or UO_47 (O_47,N_26732,N_26465);
xnor UO_48 (O_48,N_29717,N_29011);
or UO_49 (O_49,N_26220,N_29075);
or UO_50 (O_50,N_27265,N_28852);
or UO_51 (O_51,N_26399,N_29491);
nand UO_52 (O_52,N_29432,N_28577);
nor UO_53 (O_53,N_25096,N_25468);
and UO_54 (O_54,N_29140,N_29098);
or UO_55 (O_55,N_25684,N_27573);
xnor UO_56 (O_56,N_26909,N_26947);
nand UO_57 (O_57,N_28665,N_26247);
or UO_58 (O_58,N_29224,N_27321);
and UO_59 (O_59,N_28883,N_25234);
and UO_60 (O_60,N_28739,N_25133);
or UO_61 (O_61,N_27960,N_28746);
or UO_62 (O_62,N_29318,N_25555);
and UO_63 (O_63,N_29156,N_29094);
nor UO_64 (O_64,N_29577,N_27824);
and UO_65 (O_65,N_25952,N_25297);
xor UO_66 (O_66,N_26916,N_26919);
nor UO_67 (O_67,N_28411,N_29867);
xor UO_68 (O_68,N_27913,N_25413);
and UO_69 (O_69,N_27521,N_27760);
or UO_70 (O_70,N_27468,N_26376);
xnor UO_71 (O_71,N_28218,N_25095);
xor UO_72 (O_72,N_25355,N_28833);
nor UO_73 (O_73,N_28009,N_25381);
nor UO_74 (O_74,N_29169,N_26537);
xnor UO_75 (O_75,N_29952,N_28260);
nor UO_76 (O_76,N_27334,N_25197);
xnor UO_77 (O_77,N_26790,N_26000);
nor UO_78 (O_78,N_26441,N_25711);
or UO_79 (O_79,N_29263,N_26603);
or UO_80 (O_80,N_28719,N_26756);
nor UO_81 (O_81,N_27845,N_27394);
nand UO_82 (O_82,N_29728,N_27452);
and UO_83 (O_83,N_28675,N_25103);
nand UO_84 (O_84,N_28781,N_29509);
nand UO_85 (O_85,N_27438,N_25843);
nand UO_86 (O_86,N_27962,N_28986);
xor UO_87 (O_87,N_25967,N_29780);
and UO_88 (O_88,N_27091,N_26258);
xor UO_89 (O_89,N_27068,N_28470);
and UO_90 (O_90,N_29572,N_28603);
nand UO_91 (O_91,N_28678,N_27707);
and UO_92 (O_92,N_29549,N_26608);
or UO_93 (O_93,N_26402,N_25501);
or UO_94 (O_94,N_28374,N_29609);
and UO_95 (O_95,N_27355,N_28204);
nand UO_96 (O_96,N_25090,N_25497);
nand UO_97 (O_97,N_25761,N_26443);
and UO_98 (O_98,N_29584,N_28841);
nor UO_99 (O_99,N_28382,N_29573);
xnor UO_100 (O_100,N_27583,N_28048);
nor UO_101 (O_101,N_29824,N_27776);
or UO_102 (O_102,N_26629,N_28810);
nor UO_103 (O_103,N_29276,N_27850);
or UO_104 (O_104,N_25922,N_27793);
xor UO_105 (O_105,N_26965,N_26291);
nand UO_106 (O_106,N_28045,N_27465);
and UO_107 (O_107,N_28467,N_26554);
or UO_108 (O_108,N_27600,N_29137);
or UO_109 (O_109,N_25180,N_29842);
and UO_110 (O_110,N_25784,N_26684);
nor UO_111 (O_111,N_28894,N_26730);
and UO_112 (O_112,N_25964,N_27945);
xor UO_113 (O_113,N_29757,N_26286);
nand UO_114 (O_114,N_27397,N_29665);
or UO_115 (O_115,N_26967,N_25324);
and UO_116 (O_116,N_27152,N_25421);
xor UO_117 (O_117,N_26060,N_27656);
nor UO_118 (O_118,N_27758,N_26869);
or UO_119 (O_119,N_26079,N_25541);
nand UO_120 (O_120,N_27360,N_28848);
nor UO_121 (O_121,N_29288,N_29259);
and UO_122 (O_122,N_26648,N_29056);
nand UO_123 (O_123,N_28307,N_29859);
or UO_124 (O_124,N_25496,N_28932);
and UO_125 (O_125,N_27721,N_27242);
or UO_126 (O_126,N_28721,N_29848);
and UO_127 (O_127,N_27145,N_25802);
nand UO_128 (O_128,N_26389,N_29045);
and UO_129 (O_129,N_27174,N_28962);
and UO_130 (O_130,N_29307,N_28673);
and UO_131 (O_131,N_25548,N_28256);
and UO_132 (O_132,N_29419,N_28611);
nor UO_133 (O_133,N_25602,N_28963);
xor UO_134 (O_134,N_26321,N_26707);
xor UO_135 (O_135,N_29913,N_26202);
nor UO_136 (O_136,N_25766,N_25962);
or UO_137 (O_137,N_28562,N_28031);
nand UO_138 (O_138,N_26081,N_25792);
and UO_139 (O_139,N_25848,N_26904);
nor UO_140 (O_140,N_29500,N_29654);
nor UO_141 (O_141,N_25499,N_27118);
and UO_142 (O_142,N_27273,N_25607);
or UO_143 (O_143,N_27504,N_26394);
and UO_144 (O_144,N_26696,N_28844);
nor UO_145 (O_145,N_29479,N_29878);
nor UO_146 (O_146,N_26150,N_27270);
or UO_147 (O_147,N_28038,N_25327);
nand UO_148 (O_148,N_26946,N_28647);
nand UO_149 (O_149,N_27918,N_27023);
nor UO_150 (O_150,N_29193,N_27005);
nor UO_151 (O_151,N_27875,N_26990);
nand UO_152 (O_152,N_27740,N_29548);
xnor UO_153 (O_153,N_25271,N_27117);
nor UO_154 (O_154,N_26057,N_29110);
or UO_155 (O_155,N_26974,N_25671);
and UO_156 (O_156,N_29969,N_25776);
nand UO_157 (O_157,N_25670,N_25478);
nor UO_158 (O_158,N_28710,N_28688);
nor UO_159 (O_159,N_29511,N_27839);
or UO_160 (O_160,N_25214,N_26780);
nor UO_161 (O_161,N_26642,N_27378);
nor UO_162 (O_162,N_26646,N_29035);
nor UO_163 (O_163,N_26833,N_25181);
and UO_164 (O_164,N_29590,N_29959);
nand UO_165 (O_165,N_26425,N_28332);
or UO_166 (O_166,N_29070,N_27140);
nand UO_167 (O_167,N_25681,N_29192);
and UO_168 (O_168,N_28612,N_27347);
and UO_169 (O_169,N_27634,N_27115);
nor UO_170 (O_170,N_27214,N_25721);
nand UO_171 (O_171,N_25786,N_25390);
or UO_172 (O_172,N_27136,N_25150);
nor UO_173 (O_173,N_25448,N_28081);
xor UO_174 (O_174,N_26935,N_26930);
nor UO_175 (O_175,N_27474,N_28971);
nor UO_176 (O_176,N_25731,N_27407);
nor UO_177 (O_177,N_27018,N_28169);
and UO_178 (O_178,N_27354,N_25065);
nand UO_179 (O_179,N_26293,N_26420);
and UO_180 (O_180,N_28733,N_27829);
nand UO_181 (O_181,N_29089,N_26120);
and UO_182 (O_182,N_26616,N_27861);
nand UO_183 (O_183,N_25379,N_27402);
and UO_184 (O_184,N_29723,N_28838);
and UO_185 (O_185,N_28314,N_29117);
nand UO_186 (O_186,N_28403,N_26250);
nor UO_187 (O_187,N_29686,N_26979);
and UO_188 (O_188,N_26352,N_29138);
xnor UO_189 (O_189,N_28907,N_27232);
and UO_190 (O_190,N_25395,N_27783);
or UO_191 (O_191,N_27040,N_29950);
nor UO_192 (O_192,N_29888,N_29813);
nor UO_193 (O_193,N_25488,N_28042);
xor UO_194 (O_194,N_29413,N_27135);
and UO_195 (O_195,N_27028,N_28112);
nand UO_196 (O_196,N_25397,N_27715);
and UO_197 (O_197,N_25408,N_28343);
or UO_198 (O_198,N_28780,N_28447);
or UO_199 (O_199,N_26136,N_26226);
xnor UO_200 (O_200,N_27033,N_26530);
nor UO_201 (O_201,N_28622,N_27931);
and UO_202 (O_202,N_27823,N_29247);
and UO_203 (O_203,N_25252,N_28444);
nand UO_204 (O_204,N_25335,N_26404);
nor UO_205 (O_205,N_27919,N_29870);
nor UO_206 (O_206,N_29828,N_25998);
nand UO_207 (O_207,N_28247,N_27653);
nand UO_208 (O_208,N_26454,N_28359);
nor UO_209 (O_209,N_25457,N_25779);
or UO_210 (O_210,N_26503,N_29114);
nor UO_211 (O_211,N_26559,N_27350);
and UO_212 (O_212,N_25080,N_27299);
nor UO_213 (O_213,N_28634,N_29274);
nor UO_214 (O_214,N_26176,N_27080);
nor UO_215 (O_215,N_28293,N_28684);
nor UO_216 (O_216,N_28047,N_27925);
nor UO_217 (O_217,N_25108,N_29528);
or UO_218 (O_218,N_29547,N_25929);
or UO_219 (O_219,N_29311,N_26933);
nand UO_220 (O_220,N_26487,N_26787);
nor UO_221 (O_221,N_25578,N_25226);
and UO_222 (O_222,N_26847,N_25807);
and UO_223 (O_223,N_29295,N_26157);
nor UO_224 (O_224,N_27904,N_25727);
and UO_225 (O_225,N_29050,N_29532);
nand UO_226 (O_226,N_27595,N_29814);
nand UO_227 (O_227,N_27283,N_28582);
nor UO_228 (O_228,N_26469,N_25956);
nand UO_229 (O_229,N_27717,N_26498);
xnor UO_230 (O_230,N_27754,N_27672);
nand UO_231 (O_231,N_29406,N_27512);
and UO_232 (O_232,N_29630,N_28428);
xnor UO_233 (O_233,N_29146,N_25078);
xnor UO_234 (O_234,N_27943,N_29688);
or UO_235 (O_235,N_27902,N_27327);
and UO_236 (O_236,N_29321,N_25049);
and UO_237 (O_237,N_27290,N_25020);
nand UO_238 (O_238,N_26364,N_28130);
or UO_239 (O_239,N_26126,N_28876);
or UO_240 (O_240,N_28913,N_28807);
and UO_241 (O_241,N_25575,N_28750);
and UO_242 (O_242,N_29091,N_25034);
nand UO_243 (O_243,N_28787,N_25383);
nor UO_244 (O_244,N_27011,N_27563);
nor UO_245 (O_245,N_28165,N_27072);
and UO_246 (O_246,N_26521,N_28159);
xor UO_247 (O_247,N_26335,N_26369);
nand UO_248 (O_248,N_26551,N_25314);
or UO_249 (O_249,N_25299,N_29253);
nor UO_250 (O_250,N_29123,N_26205);
nor UO_251 (O_251,N_28223,N_25586);
and UO_252 (O_252,N_29296,N_29816);
or UO_253 (O_253,N_29104,N_26628);
nand UO_254 (O_254,N_28866,N_26011);
and UO_255 (O_255,N_26076,N_28415);
nor UO_256 (O_256,N_25606,N_28214);
xnor UO_257 (O_257,N_25378,N_29013);
and UO_258 (O_258,N_27741,N_25860);
or UO_259 (O_259,N_27618,N_27690);
xor UO_260 (O_260,N_29450,N_25870);
or UO_261 (O_261,N_26806,N_28728);
or UO_262 (O_262,N_26535,N_26432);
and UO_263 (O_263,N_26957,N_25147);
xor UO_264 (O_264,N_27719,N_25447);
or UO_265 (O_265,N_26816,N_27864);
nor UO_266 (O_266,N_28453,N_28830);
or UO_267 (O_267,N_26127,N_28754);
nor UO_268 (O_268,N_28532,N_27082);
nor UO_269 (O_269,N_27049,N_29923);
nor UO_270 (O_270,N_25024,N_26312);
xnor UO_271 (O_271,N_29739,N_26107);
nand UO_272 (O_272,N_29368,N_27257);
or UO_273 (O_273,N_29917,N_27188);
or UO_274 (O_274,N_25859,N_25895);
or UO_275 (O_275,N_28834,N_29157);
nand UO_276 (O_276,N_26953,N_26148);
nand UO_277 (O_277,N_29447,N_29069);
and UO_278 (O_278,N_29107,N_26319);
nand UO_279 (O_279,N_27597,N_28414);
nand UO_280 (O_280,N_27832,N_29709);
or UO_281 (O_281,N_27070,N_25570);
nor UO_282 (O_282,N_29407,N_29657);
and UO_283 (O_283,N_27694,N_27485);
or UO_284 (O_284,N_26959,N_27289);
or UO_285 (O_285,N_25898,N_25655);
and UO_286 (O_286,N_29810,N_28878);
nor UO_287 (O_287,N_26731,N_26095);
nor UO_288 (O_288,N_27891,N_28858);
nand UO_289 (O_289,N_27297,N_25106);
and UO_290 (O_290,N_25510,N_25946);
xnor UO_291 (O_291,N_29902,N_28525);
xnor UO_292 (O_292,N_29443,N_25628);
nand UO_293 (O_293,N_28677,N_26769);
nor UO_294 (O_294,N_28817,N_27970);
or UO_295 (O_295,N_25783,N_26759);
nand UO_296 (O_296,N_29189,N_27047);
xor UO_297 (O_297,N_29212,N_27235);
or UO_298 (O_298,N_27073,N_29005);
or UO_299 (O_299,N_28095,N_26981);
and UO_300 (O_300,N_27734,N_25120);
nor UO_301 (O_301,N_29294,N_25056);
nand UO_302 (O_302,N_29513,N_26357);
nand UO_303 (O_303,N_26625,N_26221);
xor UO_304 (O_304,N_25275,N_25660);
nand UO_305 (O_305,N_27604,N_27599);
xor UO_306 (O_306,N_27886,N_27948);
nor UO_307 (O_307,N_28759,N_25333);
or UO_308 (O_308,N_26378,N_28556);
nor UO_309 (O_309,N_29760,N_29641);
nor UO_310 (O_310,N_25620,N_26103);
nor UO_311 (O_311,N_29150,N_26179);
xor UO_312 (O_312,N_27746,N_27625);
or UO_313 (O_313,N_28504,N_29749);
nor UO_314 (O_314,N_25196,N_29310);
and UO_315 (O_315,N_27302,N_26660);
or UO_316 (O_316,N_25622,N_27054);
or UO_317 (O_317,N_28311,N_25845);
nand UO_318 (O_318,N_27965,N_27292);
or UO_319 (O_319,N_26733,N_28396);
nand UO_320 (O_320,N_25194,N_29664);
and UO_321 (O_321,N_25089,N_25518);
nor UO_322 (O_322,N_27930,N_27837);
nor UO_323 (O_323,N_28869,N_28155);
nor UO_324 (O_324,N_28319,N_29428);
or UO_325 (O_325,N_26259,N_25608);
or UO_326 (O_326,N_27554,N_27658);
nor UO_327 (O_327,N_26068,N_26750);
nor UO_328 (O_328,N_25186,N_27916);
and UO_329 (O_329,N_28884,N_28208);
or UO_330 (O_330,N_28197,N_26856);
and UO_331 (O_331,N_26842,N_26962);
nor UO_332 (O_332,N_27165,N_28101);
or UO_333 (O_333,N_29200,N_27834);
nand UO_334 (O_334,N_28079,N_29036);
and UO_335 (O_335,N_29984,N_25893);
nor UO_336 (O_336,N_26994,N_29744);
xor UO_337 (O_337,N_25283,N_27567);
or UO_338 (O_338,N_28249,N_29747);
xor UO_339 (O_339,N_26114,N_25869);
and UO_340 (O_340,N_25014,N_25785);
nand UO_341 (O_341,N_26390,N_27728);
nor UO_342 (O_342,N_25673,N_28476);
and UO_343 (O_343,N_26477,N_28541);
nand UO_344 (O_344,N_28458,N_25572);
nand UO_345 (O_345,N_25365,N_29093);
xor UO_346 (O_346,N_29163,N_26279);
and UO_347 (O_347,N_26742,N_28867);
nand UO_348 (O_348,N_29553,N_28707);
or UO_349 (O_349,N_29994,N_25115);
or UO_350 (O_350,N_27836,N_29442);
and UO_351 (O_351,N_29585,N_25529);
xnor UO_352 (O_352,N_27045,N_26523);
nor UO_353 (O_353,N_28025,N_25905);
and UO_354 (O_354,N_29784,N_25124);
xor UO_355 (O_355,N_25760,N_26145);
nor UO_356 (O_356,N_29403,N_27820);
or UO_357 (O_357,N_26146,N_28644);
and UO_358 (O_358,N_25101,N_26896);
and UO_359 (O_359,N_29468,N_27151);
nor UO_360 (O_360,N_29121,N_25941);
nand UO_361 (O_361,N_25460,N_25352);
or UO_362 (O_362,N_27977,N_25212);
nand UO_363 (O_363,N_25914,N_29229);
or UO_364 (O_364,N_29769,N_28923);
and UO_365 (O_365,N_29740,N_25771);
and UO_366 (O_366,N_27419,N_28316);
nor UO_367 (O_367,N_27408,N_27213);
xor UO_368 (O_368,N_29835,N_26186);
or UO_369 (O_369,N_29282,N_26789);
or UO_370 (O_370,N_28351,N_25098);
and UO_371 (O_371,N_25694,N_29668);
nor UO_372 (O_372,N_26803,N_27443);
nor UO_373 (O_373,N_25705,N_26617);
nor UO_374 (O_374,N_27128,N_27412);
nand UO_375 (O_375,N_25517,N_28119);
and UO_376 (O_376,N_26003,N_28544);
nand UO_377 (O_377,N_25306,N_28599);
xor UO_378 (O_378,N_26257,N_27827);
nand UO_379 (O_379,N_27053,N_26452);
and UO_380 (O_380,N_26864,N_29417);
xnor UO_381 (O_381,N_27342,N_25944);
nand UO_382 (O_382,N_26051,N_29425);
nor UO_383 (O_383,N_29476,N_25153);
nand UO_384 (O_384,N_25060,N_27052);
nor UO_385 (O_385,N_28229,N_25267);
xor UO_386 (O_386,N_26895,N_29153);
and UO_387 (O_387,N_28845,N_25256);
nand UO_388 (O_388,N_25303,N_29650);
nor UO_389 (O_389,N_28920,N_27897);
and UO_390 (O_390,N_28252,N_26032);
and UO_391 (O_391,N_29087,N_28902);
nand UO_392 (O_392,N_29440,N_26718);
nand UO_393 (O_393,N_28439,N_26137);
nand UO_394 (O_394,N_27475,N_27466);
nor UO_395 (O_395,N_25752,N_26231);
nand UO_396 (O_396,N_26239,N_27365);
nand UO_397 (O_397,N_25063,N_25823);
or UO_398 (O_398,N_28406,N_26570);
or UO_399 (O_399,N_28765,N_28660);
and UO_400 (O_400,N_25667,N_28085);
nand UO_401 (O_401,N_25000,N_25729);
nand UO_402 (O_402,N_27581,N_26343);
nand UO_403 (O_403,N_27341,N_26500);
nor UO_404 (O_404,N_26456,N_27139);
and UO_405 (O_405,N_28680,N_28764);
nor UO_406 (O_406,N_26671,N_25289);
xor UO_407 (O_407,N_29675,N_28956);
and UO_408 (O_408,N_26006,N_25701);
xor UO_409 (O_409,N_29405,N_25617);
or UO_410 (O_410,N_26344,N_28564);
or UO_411 (O_411,N_25099,N_28114);
nand UO_412 (O_412,N_28370,N_25152);
xnor UO_413 (O_413,N_29347,N_26828);
nor UO_414 (O_414,N_26837,N_26647);
nand UO_415 (O_415,N_25966,N_26689);
and UO_416 (O_416,N_28699,N_27863);
or UO_417 (O_417,N_29329,N_29213);
or UO_418 (O_418,N_25739,N_25524);
nand UO_419 (O_419,N_25744,N_25041);
or UO_420 (O_420,N_25320,N_27374);
and UO_421 (O_421,N_25634,N_29017);
nand UO_422 (O_422,N_27453,N_25698);
nand UO_423 (O_423,N_27523,N_27017);
nand UO_424 (O_424,N_28589,N_26034);
and UO_425 (O_425,N_29948,N_27967);
or UO_426 (O_426,N_29601,N_26639);
and UO_427 (O_427,N_29845,N_29402);
xor UO_428 (O_428,N_29614,N_27933);
xnor UO_429 (O_429,N_28703,N_27805);
nor UO_430 (O_430,N_29024,N_26327);
nand UO_431 (O_431,N_29762,N_26835);
nand UO_432 (O_432,N_27250,N_26119);
and UO_433 (O_433,N_29016,N_26388);
or UO_434 (O_434,N_28288,N_29682);
nand UO_435 (O_435,N_27349,N_26409);
and UO_436 (O_436,N_25238,N_29088);
nor UO_437 (O_437,N_27106,N_29569);
nand UO_438 (O_438,N_29946,N_27790);
xor UO_439 (O_439,N_26907,N_29438);
nor UO_440 (O_440,N_28327,N_27821);
and UO_441 (O_441,N_26875,N_26485);
nor UO_442 (O_442,N_25205,N_26256);
and UO_443 (O_443,N_27020,N_27607);
xor UO_444 (O_444,N_25775,N_29076);
nor UO_445 (O_445,N_27540,N_29985);
nand UO_446 (O_446,N_29864,N_28373);
nand UO_447 (O_447,N_25668,N_28346);
nor UO_448 (O_448,N_27574,N_26565);
or UO_449 (O_449,N_27294,N_25897);
nand UO_450 (O_450,N_28182,N_28957);
nor UO_451 (O_451,N_27089,N_29542);
nand UO_452 (O_452,N_28215,N_28793);
nor UO_453 (O_453,N_25122,N_29115);
nor UO_454 (O_454,N_28206,N_26330);
nand UO_455 (O_455,N_29851,N_25616);
nor UO_456 (O_456,N_26096,N_25010);
or UO_457 (O_457,N_28129,N_27142);
nor UO_458 (O_458,N_27878,N_29400);
xnor UO_459 (O_459,N_26260,N_28741);
or UO_460 (O_460,N_25830,N_26296);
or UO_461 (O_461,N_28409,N_29342);
nor UO_462 (O_462,N_27676,N_27366);
and UO_463 (O_463,N_29904,N_28140);
and UO_464 (O_464,N_29627,N_26724);
nor UO_465 (O_465,N_26960,N_27825);
nor UO_466 (O_466,N_29628,N_28979);
nand UO_467 (O_467,N_25533,N_26852);
nor UO_468 (O_468,N_28168,N_28184);
or UO_469 (O_469,N_28672,N_26001);
nand UO_470 (O_470,N_28146,N_28050);
and UO_471 (O_471,N_29891,N_27701);
nand UO_472 (O_472,N_26717,N_29343);
xor UO_473 (O_473,N_25975,N_25596);
or UO_474 (O_474,N_26575,N_26923);
nand UO_475 (O_475,N_28485,N_28887);
xnor UO_476 (O_476,N_28714,N_27752);
nor UO_477 (O_477,N_27792,N_27876);
and UO_478 (O_478,N_27367,N_28928);
and UO_479 (O_479,N_26222,N_29431);
and UO_480 (O_480,N_27048,N_29309);
nor UO_481 (O_481,N_25647,N_26849);
nand UO_482 (O_482,N_27030,N_26194);
or UO_483 (O_483,N_25139,N_26690);
nand UO_484 (O_484,N_29279,N_29201);
xnor UO_485 (O_485,N_29655,N_27695);
nand UO_486 (O_486,N_25407,N_25135);
or UO_487 (O_487,N_29021,N_28304);
nor UO_488 (O_488,N_28070,N_25232);
nand UO_489 (O_489,N_27808,N_25431);
nor UO_490 (O_490,N_25988,N_27134);
or UO_491 (O_491,N_28642,N_25357);
nand UO_492 (O_492,N_29836,N_28657);
nor UO_493 (O_493,N_28438,N_28041);
nor UO_494 (O_494,N_25219,N_26016);
and UO_495 (O_495,N_28667,N_26218);
or UO_496 (O_496,N_28970,N_26592);
or UO_497 (O_497,N_25302,N_28181);
and UO_498 (O_498,N_25822,N_25505);
nor UO_499 (O_499,N_25949,N_27680);
nand UO_500 (O_500,N_25040,N_29260);
nand UO_501 (O_501,N_29202,N_28605);
nor UO_502 (O_502,N_26538,N_28579);
nand UO_503 (O_503,N_27708,N_27692);
nand UO_504 (O_504,N_25899,N_25423);
nand UO_505 (O_505,N_27233,N_26743);
and UO_506 (O_506,N_27667,N_28639);
nand UO_507 (O_507,N_25305,N_25285);
or UO_508 (O_508,N_26140,N_29940);
nor UO_509 (O_509,N_25486,N_29471);
and UO_510 (O_510,N_29911,N_26952);
xor UO_511 (O_511,N_29947,N_29589);
nor UO_512 (O_512,N_28726,N_25706);
and UO_513 (O_513,N_26391,N_25174);
and UO_514 (O_514,N_28850,N_27398);
nor UO_515 (O_515,N_26713,N_27497);
or UO_516 (O_516,N_26880,N_29919);
nor UO_517 (O_517,N_26457,N_29458);
and UO_518 (O_518,N_26020,N_29194);
nor UO_519 (O_519,N_28259,N_27437);
and UO_520 (O_520,N_25747,N_26384);
nand UO_521 (O_521,N_29748,N_26812);
or UO_522 (O_522,N_27186,N_28488);
nor UO_523 (O_523,N_25494,N_26802);
and UO_524 (O_524,N_28910,N_29061);
nand UO_525 (O_525,N_29699,N_25676);
or UO_526 (O_526,N_28212,N_28098);
nand UO_527 (O_527,N_27535,N_29131);
and UO_528 (O_528,N_26059,N_25313);
nor UO_529 (O_529,N_27949,N_26162);
nor UO_530 (O_530,N_29633,N_29214);
xor UO_531 (O_531,N_26490,N_26426);
or UO_532 (O_532,N_26185,N_28618);
nand UO_533 (O_533,N_27450,N_26099);
and UO_534 (O_534,N_29292,N_29422);
or UO_535 (O_535,N_29944,N_26522);
and UO_536 (O_536,N_28334,N_27051);
nor UO_537 (O_537,N_27146,N_28075);
and UO_538 (O_538,N_26453,N_28349);
nand UO_539 (O_539,N_28555,N_26014);
xnor UO_540 (O_540,N_29285,N_26810);
nor UO_541 (O_541,N_26492,N_25254);
nand UO_542 (O_542,N_29990,N_28508);
nand UO_543 (O_543,N_26720,N_27517);
nand UO_544 (O_544,N_28904,N_28918);
xor UO_545 (O_545,N_25483,N_27110);
nand UO_546 (O_546,N_28076,N_25459);
nand UO_547 (O_547,N_26729,N_28551);
nor UO_548 (O_548,N_26187,N_26314);
and UO_549 (O_549,N_28682,N_26203);
and UO_550 (O_550,N_27212,N_27555);
nand UO_551 (O_551,N_27220,N_25853);
nand UO_552 (O_552,N_25871,N_26383);
nand UO_553 (O_553,N_25902,N_29783);
or UO_554 (O_554,N_29795,N_25609);
or UO_555 (O_555,N_29336,N_26488);
xnor UO_556 (O_556,N_28794,N_27938);
and UO_557 (O_557,N_28625,N_26872);
or UO_558 (O_558,N_29711,N_27377);
nand UO_559 (O_559,N_26037,N_26154);
nand UO_560 (O_560,N_26637,N_27800);
or UO_561 (O_561,N_29979,N_29291);
nor UO_562 (O_562,N_27149,N_25591);
nand UO_563 (O_563,N_28698,N_29457);
or UO_564 (O_564,N_26062,N_29485);
nor UO_565 (O_565,N_27236,N_26741);
or UO_566 (O_566,N_25295,N_27100);
nand UO_567 (O_567,N_29452,N_29191);
or UO_568 (O_568,N_29286,N_26511);
nand UO_569 (O_569,N_27464,N_29171);
and UO_570 (O_570,N_25341,N_26340);
nor UO_571 (O_571,N_29872,N_28299);
or UO_572 (O_572,N_25334,N_29698);
or UO_573 (O_573,N_29401,N_29350);
and UO_574 (O_574,N_26797,N_27368);
nand UO_575 (O_575,N_28694,N_27390);
or UO_576 (O_576,N_26212,N_25130);
or UO_577 (O_577,N_29225,N_26448);
or UO_578 (O_578,N_28454,N_26436);
nor UO_579 (O_579,N_26621,N_26117);
or UO_580 (O_580,N_29517,N_26366);
xnor UO_581 (O_581,N_27009,N_29498);
and UO_582 (O_582,N_29726,N_25707);
nor UO_583 (O_583,N_26489,N_27209);
xor UO_584 (O_584,N_29503,N_27078);
or UO_585 (O_585,N_29703,N_28473);
or UO_586 (O_586,N_27705,N_28813);
and UO_587 (O_587,N_26737,N_25151);
xor UO_588 (O_588,N_27206,N_27994);
or UO_589 (O_589,N_28376,N_25279);
and UO_590 (O_590,N_26542,N_26586);
or UO_591 (O_591,N_29380,N_26029);
xnor UO_592 (O_592,N_27105,N_25424);
or UO_593 (O_593,N_29588,N_28093);
and UO_594 (O_594,N_27847,N_29954);
or UO_595 (O_595,N_29666,N_29580);
or UO_596 (O_596,N_25026,N_27530);
nand UO_597 (O_597,N_27616,N_29807);
and UO_598 (O_598,N_25084,N_28935);
and UO_599 (O_599,N_27160,N_25748);
and UO_600 (O_600,N_27278,N_26313);
nor UO_601 (O_601,N_26190,N_26768);
xnor UO_602 (O_602,N_27346,N_29606);
nand UO_603 (O_603,N_29649,N_26640);
nand UO_604 (O_604,N_28683,N_25366);
or UO_605 (O_605,N_28799,N_26105);
and UO_606 (O_606,N_28980,N_28421);
or UO_607 (O_607,N_25086,N_29843);
or UO_608 (O_608,N_28198,N_25528);
nor UO_609 (O_609,N_25412,N_26371);
and UO_610 (O_610,N_29858,N_25852);
nand UO_611 (O_611,N_25636,N_29731);
and UO_612 (O_612,N_28117,N_28364);
or UO_613 (O_613,N_26914,N_27014);
xor UO_614 (O_614,N_28153,N_28823);
nand UO_615 (O_615,N_25434,N_26866);
nand UO_616 (O_616,N_28174,N_28232);
or UO_617 (O_617,N_28811,N_27296);
xor UO_618 (O_618,N_27534,N_29474);
nor UO_619 (O_619,N_26606,N_27060);
xor UO_620 (O_620,N_25117,N_27323);
xor UO_621 (O_621,N_28898,N_26948);
nand UO_622 (O_622,N_26987,N_26289);
and UO_623 (O_623,N_27436,N_26813);
and UO_624 (O_624,N_27689,N_29124);
and UO_625 (O_625,N_29887,N_25426);
nor UO_626 (O_626,N_28791,N_29916);
nor UO_627 (O_627,N_26098,N_27987);
or UO_628 (O_628,N_25027,N_26066);
and UO_629 (O_629,N_28496,N_27711);
nor UO_630 (O_630,N_26173,N_27371);
and UO_631 (O_631,N_27771,N_25980);
nand UO_632 (O_632,N_27972,N_29111);
nand UO_633 (O_633,N_28292,N_29690);
nand UO_634 (O_634,N_27156,N_27230);
nor UO_635 (O_635,N_25974,N_26623);
and UO_636 (O_636,N_29448,N_25985);
xor UO_637 (O_637,N_26885,N_25677);
nand UO_638 (O_638,N_28567,N_29672);
xnor UO_639 (O_639,N_25043,N_27881);
xor UO_640 (O_640,N_26329,N_27778);
or UO_641 (O_641,N_28100,N_27831);
nor UO_642 (O_642,N_26080,N_26093);
and UO_643 (O_643,N_28188,N_26408);
xor UO_644 (O_644,N_28437,N_26238);
and UO_645 (O_645,N_27853,N_28951);
nand UO_646 (O_646,N_25440,N_25051);
or UO_647 (O_647,N_29238,N_28952);
or UO_648 (O_648,N_26549,N_26821);
and UO_649 (O_649,N_28027,N_28104);
nor UO_650 (O_650,N_28797,N_27589);
nand UO_651 (O_651,N_29085,N_27835);
nor UO_652 (O_652,N_27435,N_25737);
nand UO_653 (O_653,N_29529,N_28772);
nor UO_654 (O_654,N_27247,N_26493);
nand UO_655 (O_655,N_27263,N_27934);
or UO_656 (O_656,N_27985,N_25888);
and UO_657 (O_657,N_28568,N_29395);
or UO_658 (O_658,N_27944,N_29871);
nand UO_659 (O_659,N_25556,N_27958);
or UO_660 (O_660,N_28966,N_25322);
nor UO_661 (O_661,N_28116,N_28254);
nor UO_662 (O_662,N_26359,N_27059);
nor UO_663 (O_663,N_26604,N_28404);
nor UO_664 (O_664,N_27502,N_25759);
or UO_665 (O_665,N_26232,N_25513);
and UO_666 (O_666,N_29015,N_27384);
nand UO_667 (O_667,N_26699,N_25259);
or UO_668 (O_668,N_27941,N_27312);
or UO_669 (O_669,N_25224,N_29866);
nand UO_670 (O_670,N_25664,N_25877);
nand UO_671 (O_671,N_25225,N_27542);
xor UO_672 (O_672,N_29176,N_27173);
or UO_673 (O_673,N_29415,N_26346);
nand UO_674 (O_674,N_27651,N_25384);
or UO_675 (O_675,N_26999,N_26225);
or UO_676 (O_676,N_25623,N_26451);
nor UO_677 (O_677,N_25948,N_27343);
or UO_678 (O_678,N_29550,N_28827);
nor UO_679 (O_679,N_27027,N_29190);
nor UO_680 (O_680,N_25207,N_27927);
nor UO_681 (O_681,N_28999,N_25545);
nand UO_682 (O_682,N_29449,N_26084);
or UO_683 (O_683,N_29359,N_28840);
or UO_684 (O_684,N_26834,N_28880);
nor UO_685 (O_685,N_26901,N_28602);
nand UO_686 (O_686,N_26631,N_29998);
and UO_687 (O_687,N_27426,N_25203);
xnor UO_688 (O_688,N_27062,N_26770);
nand UO_689 (O_689,N_29268,N_27578);
xor UO_690 (O_690,N_26261,N_27733);
nand UO_691 (O_691,N_26871,N_26412);
nor UO_692 (O_692,N_29249,N_28925);
or UO_693 (O_693,N_28016,N_25745);
or UO_694 (O_694,N_26650,N_29470);
nor UO_695 (O_695,N_26072,N_27391);
and UO_696 (O_696,N_26236,N_26761);
xor UO_697 (O_697,N_25451,N_26860);
or UO_698 (O_698,N_25428,N_28124);
and UO_699 (O_699,N_26168,N_26118);
nand UO_700 (O_700,N_26941,N_27457);
nand UO_701 (O_701,N_25316,N_28598);
and UO_702 (O_702,N_27291,N_28713);
nor UO_703 (O_703,N_26970,N_29554);
and UO_704 (O_704,N_25185,N_29314);
nor UO_705 (O_705,N_25751,N_27594);
nor UO_706 (O_706,N_29079,N_25960);
nor UO_707 (O_707,N_28617,N_29181);
nor UO_708 (O_708,N_29512,N_28594);
nor UO_709 (O_709,N_27133,N_27887);
nor UO_710 (O_710,N_27763,N_27267);
or UO_711 (O_711,N_28135,N_29411);
nor UO_712 (O_712,N_29390,N_29064);
nand UO_713 (O_713,N_25872,N_26323);
nand UO_714 (O_714,N_25167,N_25507);
nand UO_715 (O_715,N_27491,N_27936);
nand UO_716 (O_716,N_28109,N_28652);
and UO_717 (O_717,N_26367,N_28068);
and UO_718 (O_718,N_26468,N_28915);
nor UO_719 (O_719,N_26749,N_29313);
nand UO_720 (O_720,N_29430,N_29333);
nand UO_721 (O_721,N_29803,N_27980);
or UO_722 (O_722,N_27169,N_25953);
nand UO_723 (O_723,N_27460,N_25458);
xnor UO_724 (O_724,N_28122,N_25336);
and UO_725 (O_725,N_29177,N_28289);
and UO_726 (O_726,N_26685,N_29849);
or UO_727 (O_727,N_26064,N_29332);
nor UO_728 (O_728,N_26867,N_26071);
nor UO_729 (O_729,N_25906,N_26892);
nor UO_730 (O_730,N_27196,N_26779);
xor UO_731 (O_731,N_28063,N_26106);
or UO_732 (O_732,N_27753,N_28484);
or UO_733 (O_733,N_26287,N_27553);
or UO_734 (O_734,N_25163,N_28697);
nor UO_735 (O_735,N_28847,N_29173);
nand UO_736 (O_736,N_27802,N_27458);
nand UO_737 (O_737,N_28614,N_25491);
nor UO_738 (O_738,N_27481,N_27182);
nand UO_739 (O_739,N_28842,N_25579);
nand UO_740 (O_740,N_29785,N_26755);
and UO_741 (O_741,N_28442,N_27781);
or UO_742 (O_742,N_25894,N_29109);
or UO_743 (O_743,N_26823,N_28219);
or UO_744 (O_744,N_26552,N_29620);
and UO_745 (O_745,N_27171,N_29393);
nor UO_746 (O_746,N_25938,N_29634);
or UO_747 (O_747,N_29582,N_27687);
nor UO_748 (O_748,N_27353,N_26562);
and UO_749 (O_749,N_26199,N_26206);
or UO_750 (O_750,N_27726,N_27159);
nand UO_751 (O_751,N_28549,N_29520);
and UO_752 (O_752,N_25882,N_25045);
nand UO_753 (O_753,N_25066,N_26877);
and UO_754 (O_754,N_25450,N_25323);
nor UO_755 (O_755,N_26379,N_27854);
and UO_756 (O_756,N_25223,N_27614);
and UO_757 (O_757,N_28399,N_25144);
or UO_758 (O_758,N_26227,N_25569);
nor UO_759 (O_759,N_25590,N_27087);
xnor UO_760 (O_760,N_27415,N_29961);
or UO_761 (O_761,N_26984,N_26046);
and UO_762 (O_762,N_27190,N_29120);
or UO_763 (O_763,N_26921,N_26809);
nand UO_764 (O_764,N_26476,N_26995);
xnor UO_765 (O_765,N_27488,N_27075);
or UO_766 (O_766,N_26262,N_26085);
nor UO_767 (O_767,N_25127,N_28988);
nor UO_768 (O_768,N_28938,N_25614);
or UO_769 (O_769,N_25091,N_25400);
nor UO_770 (O_770,N_28294,N_28731);
nand UO_771 (O_771,N_27505,N_28596);
xor UO_772 (O_772,N_25261,N_29564);
nand UO_773 (O_773,N_28738,N_27476);
and UO_774 (O_774,N_29376,N_26484);
nor UO_775 (O_775,N_28446,N_26470);
nor UO_776 (O_776,N_25963,N_25138);
nand UO_777 (O_777,N_27743,N_29768);
nor UO_778 (O_778,N_29679,N_27389);
nor UO_779 (O_779,N_28275,N_28195);
nand UO_780 (O_780,N_25444,N_25580);
nand UO_781 (O_781,N_29647,N_25654);
and UO_782 (O_782,N_25128,N_28342);
xnor UO_783 (O_783,N_25255,N_28032);
nand UO_784 (O_784,N_25959,N_26794);
and UO_785 (O_785,N_28662,N_25925);
and UO_786 (O_786,N_26615,N_28565);
xor UO_787 (O_787,N_29315,N_26557);
xnor UO_788 (O_788,N_25142,N_28906);
nand UO_789 (O_789,N_28245,N_25884);
nor UO_790 (O_790,N_29281,N_28331);
nand UO_791 (O_791,N_28060,N_26245);
nand UO_792 (O_792,N_27215,N_25149);
xnor UO_793 (O_793,N_28640,N_27564);
and UO_794 (O_794,N_29708,N_26912);
or UO_795 (O_795,N_29059,N_29621);
or UO_796 (O_796,N_27102,N_26002);
and UO_797 (O_797,N_27245,N_28690);
nor UO_798 (O_798,N_25639,N_28018);
nor UO_799 (O_799,N_29971,N_25164);
nor UO_800 (O_800,N_29481,N_27280);
and UO_801 (O_801,N_29416,N_26027);
nor UO_802 (O_802,N_25746,N_29974);
or UO_803 (O_803,N_29043,N_27946);
or UO_804 (O_804,N_26031,N_25044);
nand UO_805 (O_805,N_27858,N_28849);
nand UO_806 (O_806,N_26697,N_25035);
xnor UO_807 (O_807,N_28000,N_28136);
and UO_808 (O_808,N_28006,N_28471);
nor UO_809 (O_809,N_26925,N_29898);
xor UO_810 (O_810,N_29965,N_28937);
nand UO_811 (O_811,N_25565,N_27037);
nor UO_812 (O_812,N_26170,N_26585);
nor UO_813 (O_813,N_29754,N_28115);
and UO_814 (O_814,N_26751,N_28199);
nor UO_815 (O_815,N_25274,N_28505);
or UO_816 (O_816,N_29487,N_28248);
and UO_817 (O_817,N_29041,N_28262);
or UO_818 (O_818,N_29755,N_25251);
nor UO_819 (O_819,N_27541,N_28241);
nor UO_820 (O_820,N_29775,N_26028);
nor UO_821 (O_821,N_28864,N_26956);
nand UO_822 (O_822,N_27720,N_27483);
nor UO_823 (O_823,N_26792,N_29988);
xnor UO_824 (O_824,N_25435,N_27427);
and UO_825 (O_825,N_27649,N_27330);
or UO_826 (O_826,N_25758,N_28983);
nor UO_827 (O_827,N_25770,N_27274);
nor UO_828 (O_828,N_25201,N_25772);
or UO_829 (O_829,N_26294,N_27851);
nor UO_830 (O_830,N_27112,N_25774);
or UO_831 (O_831,N_28228,N_28871);
and UO_832 (O_832,N_26128,N_27373);
and UO_833 (O_833,N_26431,N_29833);
nor UO_834 (O_834,N_26868,N_28992);
and UO_835 (O_835,N_25803,N_27648);
nor UO_836 (O_836,N_28086,N_28227);
nand UO_837 (O_837,N_25939,N_26161);
xor UO_838 (O_838,N_26301,N_29808);
nor UO_839 (O_839,N_26043,N_28046);
nand UO_840 (O_840,N_29031,N_27755);
xnor UO_841 (O_841,N_25819,N_25053);
and UO_842 (O_842,N_25360,N_26241);
nand UO_843 (O_843,N_25277,N_29037);
nand UO_844 (O_844,N_27871,N_28853);
nand UO_845 (O_845,N_28011,N_28147);
nor UO_846 (O_846,N_25840,N_26614);
or UO_847 (O_847,N_28173,N_26113);
nor UO_848 (O_848,N_29782,N_29837);
and UO_849 (O_849,N_28522,N_26495);
nor UO_850 (O_850,N_25855,N_27090);
nand UO_851 (O_851,N_28643,N_26381);
and UO_852 (O_852,N_25874,N_26350);
and UO_853 (O_853,N_28279,N_28695);
or UO_854 (O_854,N_26077,N_29499);
or UO_855 (O_855,N_25926,N_26672);
xor UO_856 (O_856,N_25984,N_28084);
xor UO_857 (O_857,N_26499,N_27951);
xnor UO_858 (O_858,N_28535,N_28655);
and UO_859 (O_859,N_28627,N_29248);
and UO_860 (O_860,N_26791,N_29032);
nor UO_861 (O_861,N_25055,N_25791);
nand UO_862 (O_862,N_26045,N_26215);
and UO_863 (O_863,N_25532,N_25347);
or UO_864 (O_864,N_27906,N_27846);
or UO_865 (O_865,N_29933,N_29681);
or UO_866 (O_866,N_29182,N_29685);
or UO_867 (O_867,N_28519,N_26711);
nand UO_868 (O_868,N_28225,N_27525);
nand UO_869 (O_869,N_28651,N_25371);
xor UO_870 (O_870,N_28233,N_29773);
nor UO_871 (O_871,N_26473,N_26198);
or UO_872 (O_872,N_27234,N_26475);
and UO_873 (O_873,N_25057,N_26430);
and UO_874 (O_874,N_29264,N_28489);
and UO_875 (O_875,N_28851,N_26055);
xor UO_876 (O_876,N_28924,N_25824);
and UO_877 (O_877,N_28604,N_28110);
nor UO_878 (O_878,N_27786,N_25813);
or UO_879 (O_879,N_28105,N_28088);
or UO_880 (O_880,N_27202,N_26278);
xor UO_881 (O_881,N_27298,N_25439);
and UO_882 (O_882,N_28091,N_27010);
and UO_883 (O_883,N_26539,N_27867);
nand UO_884 (O_884,N_26772,N_26655);
nor UO_885 (O_885,N_29560,N_29973);
xnor UO_886 (O_886,N_27421,N_25931);
nor UO_887 (O_887,N_29526,N_27266);
and UO_888 (O_888,N_27153,N_29196);
nand UO_889 (O_889,N_27959,N_26534);
and UO_890 (O_890,N_28818,N_26836);
and UO_891 (O_891,N_26725,N_28255);
or UO_892 (O_892,N_25016,N_27199);
and UO_893 (O_893,N_29882,N_29790);
nor UO_894 (O_894,N_29603,N_26434);
xnor UO_895 (O_895,N_25420,N_27372);
or UO_896 (O_896,N_29195,N_26067);
or UO_897 (O_897,N_26691,N_28151);
and UO_898 (O_898,N_29022,N_25452);
nand UO_899 (O_899,N_26748,N_27262);
nor UO_900 (O_900,N_27731,N_28286);
nor UO_901 (O_901,N_26405,N_26998);
and UO_902 (O_902,N_27038,N_26110);
nand UO_903 (O_903,N_29184,N_27484);
nor UO_904 (O_904,N_25641,N_27543);
and UO_905 (O_905,N_29970,N_27872);
or UO_906 (O_906,N_29218,N_26180);
and UO_907 (O_907,N_27315,N_28908);
nand UO_908 (O_908,N_26017,N_27329);
nand UO_909 (O_909,N_28524,N_28363);
xnor UO_910 (O_910,N_29518,N_27901);
nand UO_911 (O_911,N_26633,N_28196);
nand UO_912 (O_912,N_27138,N_25411);
nor UO_913 (O_913,N_26634,N_29465);
and UO_914 (O_914,N_27392,N_26428);
xor UO_915 (O_915,N_26270,N_28277);
and UO_916 (O_916,N_26191,N_28337);
xnor UO_917 (O_917,N_26310,N_29543);
nor UO_918 (O_918,N_25618,N_27332);
or UO_919 (O_919,N_26048,N_26982);
or UO_920 (O_920,N_28236,N_27668);
nand UO_921 (O_921,N_26265,N_25943);
nor UO_922 (O_922,N_25753,N_29492);
nor UO_923 (O_923,N_26547,N_26502);
nor UO_924 (O_924,N_29262,N_26295);
nor UO_925 (O_925,N_25017,N_27991);
and UO_926 (O_926,N_25441,N_28771);
and UO_927 (O_927,N_27406,N_26131);
or UO_928 (O_928,N_29976,N_26680);
nand UO_929 (O_929,N_27413,N_25626);
nand UO_930 (O_930,N_28580,N_29719);
nand UO_931 (O_931,N_27132,N_27922);
nor UO_932 (O_932,N_26726,N_28284);
nand UO_933 (O_933,N_26739,N_25188);
nand UO_934 (O_934,N_27666,N_25266);
or UO_935 (O_935,N_29025,N_25342);
or UO_936 (O_936,N_25114,N_25268);
nand UO_937 (O_937,N_26165,N_27094);
nand UO_938 (O_938,N_26858,N_25750);
and UO_939 (O_939,N_26899,N_27031);
or UO_940 (O_940,N_25364,N_28487);
or UO_941 (O_941,N_28203,N_28040);
nor UO_942 (O_942,N_27300,N_26387);
or UO_943 (O_943,N_28982,N_28661);
xor UO_944 (O_944,N_26590,N_25723);
or UO_945 (O_945,N_27981,N_25003);
and UO_946 (O_946,N_25951,N_28322);
nor UO_947 (O_947,N_27240,N_27923);
or UO_948 (O_948,N_25604,N_28691);
and UO_949 (O_949,N_25244,N_29906);
nand UO_950 (O_950,N_27098,N_28757);
and UO_951 (O_951,N_27947,N_28015);
nand UO_952 (O_952,N_28779,N_28789);
or UO_953 (O_953,N_28257,N_28786);
and UO_954 (O_954,N_28595,N_25240);
xnor UO_955 (O_955,N_27688,N_27531);
nand UO_956 (O_956,N_28435,N_27639);
nor UO_957 (O_957,N_27462,N_28514);
nand UO_958 (O_958,N_27370,N_29331);
nor UO_959 (O_959,N_27852,N_27900);
and UO_960 (O_960,N_29801,N_27841);
or UO_961 (O_961,N_28192,N_27914);
and UO_962 (O_962,N_27633,N_27439);
nor UO_963 (O_963,N_25691,N_26063);
nand UO_964 (O_964,N_28265,N_27963);
nor UO_965 (O_965,N_29636,N_28766);
and UO_966 (O_966,N_29945,N_25597);
and UO_967 (O_967,N_29381,N_26075);
nor UO_968 (O_968,N_25583,N_27729);
or UO_969 (O_969,N_25179,N_25028);
nor UO_970 (O_970,N_26855,N_26087);
nor UO_971 (O_971,N_26519,N_28681);
and UO_972 (O_972,N_26526,N_28036);
nor UO_973 (O_973,N_29936,N_26795);
nand UO_974 (O_974,N_25104,N_25137);
nand UO_975 (O_975,N_29832,N_25291);
and UO_976 (O_976,N_28216,N_27571);
nor UO_977 (O_977,N_26807,N_27609);
xnor UO_978 (O_978,N_25317,N_29216);
xnor UO_979 (O_979,N_25726,N_25594);
and UO_980 (O_980,N_29889,N_27470);
and UO_981 (O_981,N_27697,N_29165);
or UO_982 (O_982,N_29467,N_26566);
xnor UO_983 (O_983,N_29704,N_29581);
or UO_984 (O_984,N_27431,N_25950);
nand UO_985 (O_985,N_29527,N_29340);
nor UO_986 (O_986,N_26958,N_25574);
nor UO_987 (O_987,N_28656,N_25730);
nor UO_988 (O_988,N_28502,N_27326);
nand UO_989 (O_989,N_25480,N_25183);
or UO_990 (O_990,N_28901,N_27092);
nand UO_991 (O_991,N_29058,N_25543);
nand UO_992 (O_992,N_28222,N_25154);
nor UO_993 (O_993,N_27702,N_25560);
and UO_994 (O_994,N_26975,N_27654);
or UO_995 (O_995,N_28860,N_25319);
nor UO_996 (O_996,N_28309,N_27756);
and UO_997 (O_997,N_25881,N_29997);
nand UO_998 (O_998,N_29397,N_25585);
and UO_999 (O_999,N_29920,N_29250);
nor UO_1000 (O_1000,N_26471,N_26516);
nor UO_1001 (O_1001,N_25191,N_28111);
xnor UO_1002 (O_1002,N_26268,N_29545);
xor UO_1003 (O_1003,N_26328,N_28133);
or UO_1004 (O_1004,N_28609,N_27910);
xnor UO_1005 (O_1005,N_25361,N_28801);
and UO_1006 (O_1006,N_28244,N_26304);
nand UO_1007 (O_1007,N_29256,N_28014);
xnor UO_1008 (O_1008,N_27647,N_28193);
nor UO_1009 (O_1009,N_27650,N_27107);
nand UO_1010 (O_1010,N_27978,N_27495);
nor UO_1011 (O_1011,N_28053,N_25001);
and UO_1012 (O_1012,N_28408,N_29706);
nor UO_1013 (O_1013,N_27924,N_25258);
nand UO_1014 (O_1014,N_28034,N_26444);
or UO_1015 (O_1015,N_26224,N_25198);
nand UO_1016 (O_1016,N_29399,N_26058);
and UO_1017 (O_1017,N_28491,N_29890);
or UO_1018 (O_1018,N_25192,N_29305);
nor UO_1019 (O_1019,N_28870,N_27903);
xor UO_1020 (O_1020,N_25100,N_26116);
or UO_1021 (O_1021,N_25213,N_29925);
or UO_1022 (O_1022,N_29996,N_25158);
and UO_1023 (O_1023,N_28497,N_28686);
or UO_1024 (O_1024,N_29352,N_28668);
nand UO_1025 (O_1025,N_28557,N_28624);
xnor UO_1026 (O_1026,N_28338,N_28940);
nand UO_1027 (O_1027,N_27550,N_25260);
and UO_1028 (O_1028,N_28872,N_26800);
nor UO_1029 (O_1029,N_29078,N_28090);
xor UO_1030 (O_1030,N_29510,N_25292);
or UO_1031 (O_1031,N_26318,N_25999);
xor UO_1032 (O_1032,N_27071,N_28231);
or UO_1033 (O_1033,N_26676,N_27905);
and UO_1034 (O_1034,N_25175,N_28916);
xor UO_1035 (O_1035,N_26662,N_29591);
or UO_1036 (O_1036,N_29139,N_26266);
xnor UO_1037 (O_1037,N_28049,N_28523);
and UO_1038 (O_1038,N_28654,N_29915);
xnor UO_1039 (O_1039,N_28553,N_27177);
nor UO_1040 (O_1040,N_29434,N_28058);
nor UO_1041 (O_1041,N_29825,N_29765);
and UO_1042 (O_1042,N_25767,N_29557);
nor UO_1043 (O_1043,N_28418,N_27081);
nor UO_1044 (O_1044,N_28976,N_27275);
and UO_1045 (O_1045,N_26407,N_29678);
and UO_1046 (O_1046,N_29280,N_27433);
nand UO_1047 (O_1047,N_25937,N_28325);
nand UO_1048 (O_1048,N_28584,N_29705);
nand UO_1049 (O_1049,N_28630,N_26561);
nand UO_1050 (O_1050,N_27767,N_25278);
or UO_1051 (O_1051,N_26712,N_27063);
xnor UO_1052 (O_1052,N_25389,N_26588);
nand UO_1053 (O_1053,N_26977,N_27345);
nor UO_1054 (O_1054,N_26532,N_26666);
nand UO_1055 (O_1055,N_25429,N_25851);
or UO_1056 (O_1056,N_29514,N_29896);
and UO_1057 (O_1057,N_29804,N_25523);
nor UO_1058 (O_1058,N_25515,N_29562);
or UO_1059 (O_1059,N_27762,N_29290);
xnor UO_1060 (O_1060,N_26709,N_28499);
nand UO_1061 (O_1061,N_28372,N_28620);
xor UO_1062 (O_1062,N_25644,N_25582);
and UO_1063 (O_1063,N_27164,N_28137);
or UO_1064 (O_1064,N_29551,N_29538);
nand UO_1065 (O_1065,N_26845,N_28356);
nand UO_1066 (O_1066,N_29635,N_29531);
nor UO_1067 (O_1067,N_27777,N_29424);
or UO_1068 (O_1068,N_28717,N_27706);
or UO_1069 (O_1069,N_25742,N_28466);
xnor UO_1070 (O_1070,N_28221,N_25052);
or UO_1071 (O_1071,N_29612,N_26543);
nand UO_1072 (O_1072,N_27545,N_29594);
nor UO_1073 (O_1073,N_27780,N_25187);
and UO_1074 (O_1074,N_27547,N_25887);
nor UO_1075 (O_1075,N_25356,N_25112);
or UO_1076 (O_1076,N_25508,N_27784);
or UO_1077 (O_1077,N_26403,N_29930);
nand UO_1078 (O_1078,N_25248,N_25989);
nor UO_1079 (O_1079,N_26413,N_29226);
and UO_1080 (O_1080,N_26442,N_25042);
or UO_1081 (O_1081,N_28460,N_29439);
and UO_1082 (O_1082,N_25465,N_29033);
nand UO_1083 (O_1083,N_26682,N_27516);
or UO_1084 (O_1084,N_25666,N_26727);
nor UO_1085 (O_1085,N_28450,N_28578);
nand UO_1086 (O_1086,N_26092,N_25372);
nand UO_1087 (O_1087,N_26508,N_26917);
nor UO_1088 (O_1088,N_26598,N_25889);
or UO_1089 (O_1089,N_28390,N_26881);
nor UO_1090 (O_1090,N_26047,N_26385);
or UO_1091 (O_1091,N_29145,N_27116);
and UO_1092 (O_1092,N_26155,N_27477);
nor UO_1093 (O_1093,N_29587,N_29644);
or UO_1094 (O_1094,N_26934,N_29245);
or UO_1095 (O_1095,N_28718,N_26922);
nand UO_1096 (O_1096,N_28243,N_29992);
xnor UO_1097 (O_1097,N_27324,N_26777);
nand UO_1098 (O_1098,N_27803,N_27161);
and UO_1099 (O_1099,N_28905,N_27013);
nor UO_1100 (O_1100,N_26694,N_29475);
nor UO_1101 (O_1101,N_28302,N_27885);
xnor UO_1102 (O_1102,N_29068,N_29312);
or UO_1103 (O_1103,N_25362,N_25241);
or UO_1104 (O_1104,N_27935,N_28103);
or UO_1105 (O_1105,N_25455,N_26244);
nor UO_1106 (O_1106,N_27219,N_29289);
nor UO_1107 (O_1107,N_25156,N_25697);
nor UO_1108 (O_1108,N_29831,N_27993);
nor UO_1109 (O_1109,N_29730,N_25558);
or UO_1110 (O_1110,N_28650,N_27417);
or UO_1111 (O_1111,N_27403,N_27200);
and UO_1112 (O_1112,N_28895,N_29370);
nor UO_1113 (O_1113,N_29597,N_26796);
nand UO_1114 (O_1114,N_25764,N_28814);
or UO_1115 (O_1115,N_29143,N_26658);
nand UO_1116 (O_1116,N_25011,N_29651);
xnor UO_1117 (O_1117,N_25502,N_27952);
or UO_1118 (O_1118,N_28017,N_25083);
nor UO_1119 (O_1119,N_25102,N_25354);
nand UO_1120 (O_1120,N_28071,N_25832);
nand UO_1121 (O_1121,N_28226,N_27764);
nor UO_1122 (O_1122,N_27682,N_27920);
nand UO_1123 (O_1123,N_26555,N_28725);
nor UO_1124 (O_1124,N_25640,N_26983);
and UO_1125 (O_1125,N_29787,N_26018);
nor UO_1126 (O_1126,N_28368,N_27029);
or UO_1127 (O_1127,N_29983,N_29727);
nand UO_1128 (O_1128,N_29382,N_28708);
or UO_1129 (O_1129,N_29166,N_28563);
and UO_1130 (O_1130,N_27414,N_27207);
nor UO_1131 (O_1131,N_25778,N_29968);
or UO_1132 (O_1132,N_29982,N_28958);
nor UO_1133 (O_1133,N_25769,N_29611);
nand UO_1134 (O_1134,N_25427,N_27067);
and UO_1135 (O_1135,N_28440,N_28819);
xor UO_1136 (O_1136,N_28326,N_29222);
nor UO_1137 (O_1137,N_26681,N_29694);
and UO_1138 (O_1138,N_29712,N_25713);
nand UO_1139 (O_1139,N_26862,N_29558);
nand UO_1140 (O_1140,N_26246,N_27019);
xnor UO_1141 (O_1141,N_29763,N_25665);
or UO_1142 (O_1142,N_28974,N_25456);
or UO_1143 (O_1143,N_25111,N_29640);
nand UO_1144 (O_1144,N_26466,N_27895);
or UO_1145 (O_1145,N_29809,N_25210);
or UO_1146 (O_1146,N_25368,N_28978);
or UO_1147 (O_1147,N_26657,N_27264);
nor UO_1148 (O_1148,N_26297,N_27718);
nor UO_1149 (O_1149,N_26918,N_27569);
and UO_1150 (O_1150,N_27992,N_26091);
nand UO_1151 (O_1151,N_28270,N_27724);
nor UO_1152 (O_1152,N_28785,N_26435);
xor UO_1153 (O_1153,N_27660,N_27501);
or UO_1154 (O_1154,N_28998,N_25294);
nor UO_1155 (O_1155,N_26024,N_29365);
or UO_1156 (O_1156,N_25612,N_25835);
nand UO_1157 (O_1157,N_28960,N_26572);
nand UO_1158 (O_1158,N_28832,N_25800);
nand UO_1159 (O_1159,N_27890,N_25978);
and UO_1160 (O_1160,N_27429,N_29918);
or UO_1161 (O_1161,N_28792,N_28461);
nor UO_1162 (O_1162,N_25863,N_26783);
xor UO_1163 (O_1163,N_26558,N_27856);
nand UO_1164 (O_1164,N_28089,N_27801);
nor UO_1165 (O_1165,N_27251,N_27806);
nand UO_1166 (O_1166,N_29283,N_29604);
nor UO_1167 (O_1167,N_26040,N_28836);
nand UO_1168 (O_1168,N_26525,N_29715);
and UO_1169 (O_1169,N_27195,N_29535);
or UO_1170 (O_1170,N_28498,N_27176);
nor UO_1171 (O_1171,N_28099,N_25059);
xor UO_1172 (O_1172,N_25388,N_28948);
and UO_1173 (O_1173,N_26363,N_25940);
and UO_1174 (O_1174,N_25903,N_28802);
nand UO_1175 (O_1175,N_25825,N_26839);
nand UO_1176 (O_1176,N_27276,N_26368);
nor UO_1177 (O_1177,N_25461,N_25328);
or UO_1178 (O_1178,N_29480,N_29793);
and UO_1179 (O_1179,N_26449,N_26844);
nor UO_1180 (O_1180,N_29839,N_29879);
nor UO_1181 (O_1181,N_28863,N_27894);
nand UO_1182 (O_1182,N_28706,N_29466);
nand UO_1183 (O_1183,N_29802,N_29330);
nor UO_1184 (O_1184,N_28828,N_25307);
or UO_1185 (O_1185,N_27788,N_25539);
nand UO_1186 (O_1186,N_27507,N_29537);
nand UO_1187 (O_1187,N_27303,N_25688);
and UO_1188 (O_1188,N_29388,N_29570);
nor UO_1189 (O_1189,N_26494,N_28865);
and UO_1190 (O_1190,N_25658,N_28881);
and UO_1191 (O_1191,N_27243,N_25296);
and UO_1192 (O_1192,N_28669,N_28981);
nor UO_1193 (O_1193,N_29638,N_26820);
nor UO_1194 (O_1194,N_29071,N_25703);
and UO_1195 (O_1195,N_29725,N_28755);
or UO_1196 (O_1196,N_29901,N_25568);
nand UO_1197 (O_1197,N_26746,N_27865);
nand UO_1198 (O_1198,N_29855,N_26233);
xnor UO_1199 (O_1199,N_28500,N_29269);
xnor UO_1200 (O_1200,N_25909,N_26316);
nor UO_1201 (O_1201,N_25125,N_29893);
nand UO_1202 (O_1202,N_25177,N_26281);
or UO_1203 (O_1203,N_26025,N_25695);
or UO_1204 (O_1204,N_29766,N_28398);
xor UO_1205 (O_1205,N_26207,N_27810);
nand UO_1206 (O_1206,N_27998,N_25675);
nor UO_1207 (O_1207,N_26805,N_26023);
and UO_1208 (O_1208,N_26300,N_25237);
nand UO_1209 (O_1209,N_27129,N_25217);
and UO_1210 (O_1210,N_28560,N_25249);
and UO_1211 (O_1211,N_28897,N_27351);
nor UO_1212 (O_1212,N_28995,N_25449);
and UO_1213 (O_1213,N_28335,N_25971);
xnor UO_1214 (O_1214,N_28194,N_28142);
and UO_1215 (O_1215,N_28583,N_25687);
nand UO_1216 (O_1216,N_28144,N_26424);
and UO_1217 (O_1217,N_27544,N_29496);
or UO_1218 (O_1218,N_28953,N_26533);
nand UO_1219 (O_1219,N_27570,N_27789);
nand UO_1220 (O_1220,N_29160,N_25704);
nor UO_1221 (O_1221,N_29600,N_29062);
xnor UO_1222 (O_1222,N_28720,N_28266);
and UO_1223 (O_1223,N_28526,N_27691);
xnor UO_1224 (O_1224,N_25464,N_29266);
or UO_1225 (O_1225,N_27703,N_29105);
nor UO_1226 (O_1226,N_29167,N_25077);
and UO_1227 (O_1227,N_25146,N_29135);
nand UO_1228 (O_1228,N_26455,N_28517);
nor UO_1229 (O_1229,N_29029,N_28635);
nor UO_1230 (O_1230,N_28931,N_29408);
or UO_1231 (O_1231,N_28874,N_29546);
nand UO_1232 (O_1232,N_28477,N_27511);
nand UO_1233 (O_1233,N_26004,N_26945);
or UO_1234 (O_1234,N_29223,N_29020);
nand UO_1235 (O_1235,N_28391,N_26653);
or UO_1236 (O_1236,N_27722,N_27386);
nand UO_1237 (O_1237,N_28175,N_25857);
or UO_1238 (O_1238,N_28354,N_26591);
or UO_1239 (O_1239,N_27175,N_25134);
or UO_1240 (O_1240,N_29598,N_28106);
nand UO_1241 (O_1241,N_29175,N_29669);
nor UO_1242 (O_1242,N_28701,N_29101);
nor UO_1243 (O_1243,N_25074,N_25910);
and UO_1244 (O_1244,N_27126,N_29892);
xor UO_1245 (O_1245,N_25506,N_29366);
xnor UO_1246 (O_1246,N_29147,N_26651);
or UO_1247 (O_1247,N_27757,N_26336);
and UO_1248 (O_1248,N_27400,N_27623);
nor UO_1249 (O_1249,N_28282,N_28899);
or UO_1250 (O_1250,N_27328,N_25009);
and UO_1251 (O_1251,N_25085,N_28339);
nand UO_1252 (O_1252,N_29593,N_26531);
and UO_1253 (O_1253,N_26217,N_29771);
nand UO_1254 (O_1254,N_25638,N_28132);
and UO_1255 (O_1255,N_26971,N_25404);
or UO_1256 (O_1256,N_28945,N_28687);
or UO_1257 (O_1257,N_28749,N_29258);
nand UO_1258 (O_1258,N_29991,N_25808);
or UO_1259 (O_1259,N_29894,N_28997);
or UO_1260 (O_1260,N_27562,N_28816);
xor UO_1261 (O_1261,N_25563,N_26213);
nand UO_1262 (O_1262,N_29774,N_26201);
or UO_1263 (O_1263,N_26624,N_29862);
nand UO_1264 (O_1264,N_27593,N_27950);
or UO_1265 (O_1265,N_26125,N_29039);
and UO_1266 (O_1266,N_26891,N_28054);
nand UO_1267 (O_1267,N_28469,N_26669);
or UO_1268 (O_1268,N_28663,N_27224);
xor UO_1269 (O_1269,N_29957,N_29776);
nor UO_1270 (O_1270,N_26406,N_25247);
nand UO_1271 (O_1271,N_29743,N_27430);
and UO_1272 (O_1272,N_29798,N_27480);
and UO_1273 (O_1273,N_28912,N_26169);
nor UO_1274 (O_1274,N_25547,N_26234);
nor UO_1275 (O_1275,N_27144,N_25521);
or UO_1276 (O_1276,N_26661,N_25525);
or UO_1277 (O_1277,N_29046,N_27241);
nand UO_1278 (O_1278,N_29158,N_28003);
nor UO_1279 (O_1279,N_27024,N_26283);
nand UO_1280 (O_1280,N_26415,N_28441);
and UO_1281 (O_1281,N_28712,N_29142);
or UO_1282 (O_1282,N_29197,N_27249);
nand UO_1283 (O_1283,N_29134,N_25867);
and UO_1284 (O_1284,N_26305,N_29713);
nor UO_1285 (O_1285,N_26786,N_29003);
or UO_1286 (O_1286,N_29541,N_28886);
nor UO_1287 (O_1287,N_26664,N_26108);
nand UO_1288 (O_1288,N_26143,N_28369);
or UO_1289 (O_1289,N_25215,N_27041);
nor UO_1290 (O_1290,N_28676,N_28890);
nor UO_1291 (O_1291,N_25454,N_28729);
nand UO_1292 (O_1292,N_26627,N_25375);
nand UO_1293 (O_1293,N_28420,N_25839);
and UO_1294 (O_1294,N_29183,N_29579);
or UO_1295 (O_1295,N_25589,N_28587);
and UO_1296 (O_1296,N_27185,N_25861);
or UO_1297 (O_1297,N_28324,N_29469);
and UO_1298 (O_1298,N_29086,N_29255);
and UO_1299 (O_1299,N_29113,N_25868);
and UO_1300 (O_1300,N_29144,N_28518);
nor UO_1301 (O_1301,N_27416,N_25942);
and UO_1302 (O_1302,N_28283,N_28475);
nor UO_1303 (O_1303,N_27463,N_25875);
nand UO_1304 (O_1304,N_29065,N_28740);
or UO_1305 (O_1305,N_29868,N_28149);
and UO_1306 (O_1306,N_27503,N_25131);
or UO_1307 (O_1307,N_26189,N_29519);
nor UO_1308 (O_1308,N_27184,N_29966);
nor UO_1309 (O_1309,N_25789,N_26763);
xor UO_1310 (O_1310,N_25797,N_25646);
nor UO_1311 (O_1311,N_29328,N_26972);
nand UO_1312 (O_1312,N_25250,N_28798);
nor UO_1313 (O_1313,N_26315,N_28278);
nand UO_1314 (O_1314,N_25022,N_28554);
nor UO_1315 (O_1315,N_27387,N_28540);
and UO_1316 (O_1316,N_29805,N_27320);
nor UO_1317 (O_1317,N_26649,N_26109);
or UO_1318 (O_1318,N_27358,N_27652);
nor UO_1319 (O_1319,N_26282,N_27193);
and UO_1320 (O_1320,N_26564,N_27500);
or UO_1321 (O_1321,N_26626,N_25717);
xor UO_1322 (O_1322,N_29907,N_25955);
nand UO_1323 (O_1323,N_25738,N_25637);
nand UO_1324 (O_1324,N_25298,N_25414);
nand UO_1325 (O_1325,N_28930,N_29610);
xnor UO_1326 (O_1326,N_28474,N_29221);
and UO_1327 (O_1327,N_26524,N_27926);
or UO_1328 (O_1328,N_29770,N_27975);
nor UO_1329 (O_1329,N_29385,N_27937);
nand UO_1330 (O_1330,N_25601,N_29244);
nor UO_1331 (O_1331,N_28944,N_29217);
nor UO_1332 (O_1332,N_25503,N_27999);
and UO_1333 (O_1333,N_25161,N_28804);
nor UO_1334 (O_1334,N_28955,N_27079);
or UO_1335 (O_1335,N_26427,N_27239);
nand UO_1336 (O_1336,N_27401,N_29857);
and UO_1337 (O_1337,N_25689,N_25805);
and UO_1338 (O_1338,N_26193,N_26988);
or UO_1339 (O_1339,N_27745,N_29980);
or UO_1340 (O_1340,N_25936,N_27785);
or UO_1341 (O_1341,N_28760,N_28285);
xnor UO_1342 (O_1342,N_25918,N_27744);
and UO_1343 (O_1343,N_25220,N_28145);
or UO_1344 (O_1344,N_28972,N_29445);
nor UO_1345 (O_1345,N_25928,N_25067);
nor UO_1346 (O_1346,N_26123,N_26560);
xnor UO_1347 (O_1347,N_28328,N_28770);
or UO_1348 (O_1348,N_26767,N_27641);
or UO_1349 (O_1349,N_29576,N_25994);
and UO_1350 (O_1350,N_27376,N_27096);
and UO_1351 (O_1351,N_27749,N_29955);
xnor UO_1352 (O_1352,N_28432,N_26708);
nand UO_1353 (O_1353,N_28623,N_29575);
or UO_1354 (O_1354,N_29583,N_27424);
nor UO_1355 (O_1355,N_29000,N_26377);
and UO_1356 (O_1356,N_27917,N_26854);
nand UO_1357 (O_1357,N_27866,N_27331);
xor UO_1358 (O_1358,N_27699,N_25157);
nor UO_1359 (O_1359,N_28615,N_28509);
and UO_1360 (O_1360,N_29924,N_25199);
or UO_1361 (O_1361,N_26209,N_25410);
nand UO_1362 (O_1362,N_29938,N_26022);
or UO_1363 (O_1363,N_26913,N_28348);
xor UO_1364 (O_1364,N_26049,N_26290);
or UO_1365 (O_1365,N_28213,N_26978);
nor UO_1366 (O_1366,N_28900,N_28067);
nand UO_1367 (O_1367,N_26438,N_25917);
nor UO_1368 (O_1368,N_28459,N_26440);
xnor UO_1369 (O_1369,N_25419,N_27735);
and UO_1370 (O_1370,N_25710,N_25923);
nor UO_1371 (O_1371,N_28743,N_25908);
and UO_1372 (O_1372,N_26667,N_26090);
nor UO_1373 (O_1373,N_29030,N_26698);
and UO_1374 (O_1374,N_28312,N_25272);
and UO_1375 (O_1375,N_27056,N_26888);
and UO_1376 (O_1376,N_29693,N_27601);
nand UO_1377 (O_1377,N_27869,N_26178);
nor UO_1378 (O_1378,N_25005,N_28207);
nor UO_1379 (O_1379,N_26130,N_29900);
nand UO_1380 (O_1380,N_28164,N_29420);
nor UO_1381 (O_1381,N_26838,N_26237);
nor UO_1382 (O_1382,N_27761,N_29325);
xor UO_1383 (O_1383,N_26038,N_29670);
and UO_1384 (O_1384,N_29530,N_28062);
or UO_1385 (O_1385,N_29745,N_27248);
and UO_1386 (O_1386,N_25409,N_25553);
nand UO_1387 (O_1387,N_26100,N_27685);
nor UO_1388 (O_1388,N_25653,N_27870);
and UO_1389 (O_1389,N_25265,N_28235);
nor UO_1390 (O_1390,N_26861,N_25386);
nor UO_1391 (O_1391,N_29846,N_29662);
xor UO_1392 (O_1392,N_27311,N_28512);
or UO_1393 (O_1393,N_26670,N_26229);
or UO_1394 (O_1394,N_25348,N_28959);
or UO_1395 (O_1395,N_25804,N_26242);
or UO_1396 (O_1396,N_25340,N_28934);
nand UO_1397 (O_1397,N_26683,N_29733);
nor UO_1398 (O_1398,N_28795,N_29881);
and UO_1399 (O_1399,N_26678,N_25806);
nor UO_1400 (O_1400,N_26890,N_29525);
and UO_1401 (O_1401,N_26906,N_26302);
xor UO_1402 (O_1402,N_26870,N_26645);
nor UO_1403 (O_1403,N_25864,N_25178);
nor UO_1404 (O_1404,N_27189,N_27335);
and UO_1405 (O_1405,N_28734,N_26338);
nor UO_1406 (O_1406,N_25293,N_28021);
nor UO_1407 (O_1407,N_25195,N_29130);
nand UO_1408 (O_1408,N_25007,N_25500);
nand UO_1409 (O_1409,N_26620,N_26898);
nor UO_1410 (O_1410,N_25968,N_28585);
xnor UO_1411 (O_1411,N_29023,N_25398);
and UO_1412 (O_1412,N_25595,N_27114);
nor UO_1413 (O_1413,N_25847,N_25610);
nand UO_1414 (O_1414,N_28653,N_26375);
and UO_1415 (O_1415,N_25118,N_29326);
or UO_1416 (O_1416,N_25756,N_25976);
and UO_1417 (O_1417,N_26263,N_29073);
or UO_1418 (O_1418,N_29317,N_27539);
nand UO_1419 (O_1419,N_28462,N_25715);
or UO_1420 (O_1420,N_27208,N_26074);
or UO_1421 (O_1421,N_28298,N_26361);
nand UO_1422 (O_1422,N_28679,N_28056);
and UO_1423 (O_1423,N_25814,N_26159);
nor UO_1424 (O_1424,N_26609,N_26584);
nand UO_1425 (O_1425,N_27748,N_26041);
nor UO_1426 (O_1426,N_28641,N_26061);
nor UO_1427 (O_1427,N_26734,N_26007);
nor UO_1428 (O_1428,N_29794,N_29676);
nand UO_1429 (O_1429,N_27043,N_27579);
or UO_1430 (O_1430,N_27446,N_27759);
xor UO_1431 (O_1431,N_27626,N_29502);
and UO_1432 (O_1432,N_25321,N_28566);
and UO_1433 (O_1433,N_27269,N_29149);
nor UO_1434 (O_1434,N_26636,N_28305);
nor UO_1435 (O_1435,N_27716,N_27619);
nor UO_1436 (O_1436,N_26808,N_29254);
nor UO_1437 (O_1437,N_29789,N_25373);
and UO_1438 (O_1438,N_28896,N_29379);
nor UO_1439 (O_1439,N_26757,N_25088);
nor UO_1440 (O_1440,N_27253,N_26513);
and UO_1441 (O_1441,N_26902,N_27281);
nand UO_1442 (O_1442,N_29823,N_29349);
and UO_1443 (O_1443,N_26182,N_25530);
and UO_1444 (O_1444,N_26692,N_29338);
nand UO_1445 (O_1445,N_25841,N_26332);
nor UO_1446 (O_1446,N_28511,N_25973);
and UO_1447 (O_1447,N_26518,N_29829);
nor UO_1448 (O_1448,N_25725,N_27111);
nor UO_1449 (O_1449,N_25921,N_27646);
nand UO_1450 (O_1450,N_25075,N_25309);
nor UO_1451 (O_1451,N_26094,N_29051);
xnor UO_1452 (O_1452,N_28839,N_29660);
nor UO_1453 (O_1453,N_26745,N_26887);
and UO_1454 (O_1454,N_29233,N_27833);
xnor UO_1455 (O_1455,N_29483,N_28559);
nor UO_1456 (O_1456,N_25669,N_28727);
or UO_1457 (O_1457,N_28638,N_28538);
nand UO_1458 (O_1458,N_27655,N_27216);
nor UO_1459 (O_1459,N_27157,N_29389);
and UO_1460 (O_1460,N_29615,N_25833);
xnor UO_1461 (O_1461,N_25004,N_28426);
or UO_1462 (O_1462,N_29301,N_25657);
nor UO_1463 (O_1463,N_27203,N_28410);
nor UO_1464 (O_1464,N_27119,N_28395);
nor UO_1465 (O_1465,N_26773,N_28671);
nand UO_1466 (O_1466,N_26474,N_28315);
and UO_1467 (O_1467,N_26240,N_26439);
nand UO_1468 (O_1468,N_28217,N_26252);
nor UO_1469 (O_1469,N_26963,N_29351);
or UO_1470 (O_1470,N_26188,N_29746);
xnor UO_1471 (O_1471,N_27809,N_28094);
and UO_1472 (O_1472,N_25013,N_29179);
xor UO_1473 (O_1473,N_26822,N_29346);
nor UO_1474 (O_1474,N_28200,N_27382);
or UO_1475 (O_1475,N_26931,N_25230);
or UO_1476 (O_1476,N_29659,N_29761);
nand UO_1477 (O_1477,N_25561,N_29377);
or UO_1478 (O_1478,N_29297,N_29937);
nor UO_1479 (O_1479,N_29007,N_29964);
or UO_1480 (O_1480,N_29034,N_29128);
nor UO_1481 (O_1481,N_28843,N_27794);
and UO_1482 (O_1482,N_25699,N_25445);
or UO_1483 (O_1483,N_27471,N_27538);
xnor UO_1484 (O_1484,N_26276,N_27714);
nor UO_1485 (O_1485,N_25740,N_26042);
and UO_1486 (O_1486,N_27288,N_27677);
nand UO_1487 (O_1487,N_27804,N_29646);
nand UO_1488 (O_1488,N_28425,N_28889);
and UO_1489 (O_1489,N_27170,N_27113);
nor UO_1490 (O_1490,N_26050,N_26355);
or UO_1491 (O_1491,N_28150,N_25566);
and UO_1492 (O_1492,N_25015,N_26459);
nor UO_1493 (O_1493,N_27396,N_28417);
or UO_1494 (O_1494,N_25924,N_28019);
and UO_1495 (O_1495,N_28597,N_27844);
nand UO_1496 (O_1496,N_29943,N_27282);
nand UO_1497 (O_1497,N_25402,N_27287);
nand UO_1498 (O_1498,N_29241,N_29738);
xnor UO_1499 (O_1499,N_28783,N_25473);
nor UO_1500 (O_1500,N_29228,N_29800);
nand UO_1501 (O_1501,N_25489,N_27380);
nor UO_1502 (O_1502,N_28443,N_25712);
or UO_1503 (O_1503,N_29354,N_28385);
xnor UO_1504 (O_1504,N_25236,N_25661);
nand UO_1505 (O_1505,N_28885,N_27409);
nor UO_1506 (O_1506,N_28808,N_29596);
nor UO_1507 (O_1507,N_28061,N_28143);
or UO_1508 (O_1508,N_25155,N_27670);
nor UO_1509 (O_1509,N_25453,N_28082);
and UO_1510 (O_1510,N_25836,N_25878);
nand UO_1511 (O_1511,N_26673,N_29962);
nor UO_1512 (O_1512,N_26771,N_27526);
nor UO_1513 (O_1513,N_27026,N_26104);
nor UO_1514 (O_1514,N_28340,N_25535);
and UO_1515 (O_1515,N_29242,N_28503);
xnor UO_1516 (O_1516,N_28954,N_27381);
and UO_1517 (O_1517,N_27322,N_28434);
and UO_1518 (O_1518,N_27843,N_28080);
nand UO_1519 (O_1519,N_27605,N_28123);
and UO_1520 (O_1520,N_29187,N_26167);
and UO_1521 (O_1521,N_25741,N_27849);
and UO_1522 (O_1522,N_27576,N_28646);
and UO_1523 (O_1523,N_25682,N_26483);
nor UO_1524 (O_1524,N_26736,N_25345);
xor UO_1525 (O_1525,N_28185,N_29631);
and UO_1526 (O_1526,N_29339,N_25732);
nor UO_1527 (O_1527,N_29209,N_27747);
or UO_1528 (O_1528,N_27513,N_29623);
or UO_1529 (O_1529,N_28702,N_29348);
nand UO_1530 (O_1530,N_28272,N_28445);
nor UO_1531 (O_1531,N_27293,N_28209);
nor UO_1532 (O_1532,N_28732,N_28321);
nand UO_1533 (O_1533,N_29516,N_28685);
nand UO_1534 (O_1534,N_28711,N_27838);
nor UO_1535 (O_1535,N_26728,N_28177);
or UO_1536 (O_1536,N_26005,N_28138);
nand UO_1537 (O_1537,N_29436,N_26546);
nor UO_1538 (O_1538,N_25765,N_27108);
or UO_1539 (O_1539,N_25559,N_25891);
nand UO_1540 (O_1540,N_28837,N_27840);
and UO_1541 (O_1541,N_27198,N_28026);
or UO_1542 (O_1542,N_25550,N_27942);
nor UO_1543 (O_1543,N_26317,N_25394);
nand UO_1544 (O_1544,N_26715,N_28493);
nand UO_1545 (O_1545,N_27879,N_29960);
or UO_1546 (O_1546,N_28715,N_26505);
or UO_1547 (O_1547,N_28761,N_28506);
and UO_1548 (O_1548,N_29559,N_29304);
or UO_1549 (O_1549,N_27314,N_27997);
and UO_1550 (O_1550,N_26618,N_25584);
nand UO_1551 (O_1551,N_27046,N_25990);
and UO_1552 (O_1552,N_26019,N_28087);
and UO_1553 (O_1553,N_26607,N_25892);
xnor UO_1554 (O_1554,N_28472,N_26910);
or UO_1555 (O_1555,N_29607,N_26195);
or UO_1556 (O_1556,N_29724,N_27404);
and UO_1557 (O_1557,N_26587,N_27423);
and UO_1558 (O_1558,N_29574,N_28465);
nand UO_1559 (O_1559,N_28528,N_27973);
and UO_1560 (O_1560,N_26078,N_26865);
and UO_1561 (O_1561,N_26905,N_26347);
nor UO_1562 (O_1562,N_26514,N_25032);
nand UO_1563 (O_1563,N_26411,N_29373);
nand UO_1564 (O_1564,N_28154,N_26365);
nor UO_1565 (O_1565,N_29103,N_26550);
nand UO_1566 (O_1566,N_26395,N_27884);
or UO_1567 (O_1567,N_29482,N_28516);
nor UO_1568 (O_1568,N_26462,N_26817);
or UO_1569 (O_1569,N_29963,N_25204);
and UO_1570 (O_1570,N_25462,N_28531);
nor UO_1571 (O_1571,N_29658,N_29639);
nor UO_1572 (O_1572,N_28570,N_29781);
nand UO_1573 (O_1573,N_26400,N_26652);
or UO_1574 (O_1574,N_29619,N_28601);
nand UO_1575 (O_1575,N_28909,N_27640);
nand UO_1576 (O_1576,N_26362,N_28569);
xor UO_1577 (O_1577,N_28608,N_26386);
nor UO_1578 (O_1578,N_27042,N_26929);
and UO_1579 (O_1579,N_25796,N_29364);
nor UO_1580 (O_1580,N_29459,N_26688);
nand UO_1581 (O_1581,N_29524,N_29186);
and UO_1582 (O_1582,N_27284,N_25932);
nor UO_1583 (O_1583,N_28413,N_29817);
and UO_1584 (O_1584,N_29796,N_28534);
xor UO_1585 (O_1585,N_25385,N_29617);
nor UO_1586 (O_1586,N_28744,N_29885);
nor UO_1587 (O_1587,N_27319,N_26993);
nand UO_1588 (O_1588,N_25162,N_29298);
and UO_1589 (O_1589,N_26251,N_26744);
nand UO_1590 (O_1590,N_26292,N_29616);
or UO_1591 (O_1591,N_26273,N_28347);
or UO_1592 (O_1592,N_28380,N_26701);
and UO_1593 (O_1593,N_26950,N_29999);
and UO_1594 (O_1594,N_27669,N_28035);
or UO_1595 (O_1595,N_29935,N_28427);
nand UO_1596 (O_1596,N_28747,N_26501);
nor UO_1597 (O_1597,N_26932,N_26504);
or UO_1598 (O_1598,N_27774,N_29028);
nand UO_1599 (O_1599,N_26576,N_27995);
nand UO_1600 (O_1600,N_28024,N_28246);
nor UO_1601 (O_1601,N_25492,N_25724);
nand UO_1602 (O_1602,N_27637,N_29671);
or UO_1603 (O_1603,N_26900,N_29127);
nor UO_1604 (O_1604,N_27172,N_25603);
xnor UO_1605 (O_1605,N_26955,N_25399);
nor UO_1606 (O_1606,N_29391,N_27440);
or UO_1607 (O_1607,N_27880,N_25554);
nor UO_1608 (O_1608,N_26752,N_26675);
nor UO_1609 (O_1609,N_28575,N_27486);
and UO_1610 (O_1610,N_26054,N_28360);
and UO_1611 (O_1611,N_28189,N_25330);
or UO_1612 (O_1612,N_28507,N_25674);
nand UO_1613 (O_1613,N_27815,N_29929);
and UO_1614 (O_1614,N_28619,N_27393);
and UO_1615 (O_1615,N_28891,N_25132);
and UO_1616 (O_1616,N_25969,N_27363);
or UO_1617 (O_1617,N_25809,N_25901);
nand UO_1618 (O_1618,N_26111,N_25504);
nor UO_1619 (O_1619,N_27304,N_28402);
nand UO_1620 (O_1620,N_25121,N_29074);
xnor UO_1621 (O_1621,N_28479,N_27000);
or UO_1622 (O_1622,N_27489,N_29082);
or UO_1623 (O_1623,N_27218,N_26857);
and UO_1624 (O_1624,N_27766,N_26491);
and UO_1625 (O_1625,N_27050,N_25184);
and UO_1626 (O_1626,N_26467,N_25846);
xnor UO_1627 (O_1627,N_26392,N_26611);
or UO_1628 (O_1628,N_26039,N_27674);
or UO_1629 (O_1629,N_27336,N_28274);
or UO_1630 (O_1630,N_28859,N_28705);
xor UO_1631 (O_1631,N_27976,N_27907);
and UO_1632 (O_1632,N_27822,N_25540);
nor UO_1633 (O_1633,N_25520,N_25023);
nand UO_1634 (O_1634,N_29363,N_29361);
or UO_1635 (O_1635,N_27221,N_26840);
nor UO_1636 (O_1636,N_29815,N_29141);
or UO_1637 (O_1637,N_27179,N_27222);
xor UO_1638 (O_1638,N_29386,N_25401);
nand UO_1639 (O_1639,N_27364,N_26373);
nor UO_1640 (O_1640,N_25418,N_29613);
nor UO_1641 (O_1641,N_25415,N_29344);
nor UO_1642 (O_1642,N_29396,N_25477);
nor UO_1643 (O_1643,N_29555,N_27383);
nand UO_1644 (O_1644,N_28361,N_25571);
nand UO_1645 (O_1645,N_26949,N_27508);
nor UO_1646 (O_1646,N_26723,N_29497);
nand UO_1647 (O_1647,N_29521,N_26641);
or UO_1648 (O_1648,N_25227,N_25073);
nor UO_1649 (O_1649,N_25062,N_28301);
and UO_1650 (O_1650,N_29811,N_28057);
nand UO_1651 (O_1651,N_27348,N_26811);
nor UO_1652 (O_1652,N_27560,N_25170);
nand UO_1653 (O_1653,N_26721,N_26228);
nand UO_1654 (O_1654,N_28933,N_28964);
nand UO_1655 (O_1655,N_25312,N_27493);
and UO_1656 (O_1656,N_28633,N_29038);
nand UO_1657 (O_1657,N_29454,N_25972);
nor UO_1658 (O_1658,N_26419,N_26613);
xor UO_1659 (O_1659,N_28250,N_27001);
nand UO_1660 (O_1660,N_28313,N_25467);
nor UO_1661 (O_1661,N_26496,N_26517);
nor UO_1662 (O_1662,N_26873,N_28806);
xnor UO_1663 (O_1663,N_29240,N_29235);
or UO_1664 (O_1664,N_26600,N_29975);
and UO_1665 (O_1665,N_25516,N_25141);
and UO_1666 (O_1666,N_26056,N_25257);
xnor UO_1667 (O_1667,N_28367,N_28490);
or UO_1668 (O_1668,N_26274,N_26747);
and UO_1669 (O_1669,N_25200,N_28456);
and UO_1670 (O_1670,N_26414,N_25437);
or UO_1671 (O_1671,N_27939,N_26345);
xnor UO_1672 (O_1672,N_26599,N_25714);
and UO_1673 (O_1673,N_26124,N_25343);
or UO_1674 (O_1674,N_27036,N_26961);
nand UO_1675 (O_1675,N_26507,N_27103);
nor UO_1676 (O_1676,N_26879,N_26339);
nor UO_1677 (O_1677,N_26147,N_27008);
and UO_1678 (O_1678,N_27811,N_26778);
nand UO_1679 (O_1679,N_25562,N_28287);
nand UO_1680 (O_1680,N_25700,N_29168);
nor UO_1681 (O_1681,N_25911,N_25495);
nand UO_1682 (O_1682,N_27590,N_28825);
and UO_1683 (O_1683,N_25820,N_27420);
and UO_1684 (O_1684,N_26115,N_27893);
nand UO_1685 (O_1685,N_29095,N_25534);
or UO_1686 (O_1686,N_26181,N_28350);
and UO_1687 (O_1687,N_26216,N_25913);
and UO_1688 (O_1688,N_29505,N_27568);
and UO_1689 (O_1689,N_29899,N_25919);
nor UO_1690 (O_1690,N_27163,N_28752);
and UO_1691 (O_1691,N_28748,N_25728);
xnor UO_1692 (O_1692,N_26360,N_26009);
nand UO_1693 (O_1693,N_25613,N_28629);
nor UO_1694 (O_1694,N_29014,N_25811);
nor UO_1695 (O_1695,N_26197,N_25329);
or UO_1696 (O_1696,N_28375,N_26776);
or UO_1697 (O_1697,N_29602,N_28574);
and UO_1698 (O_1698,N_26208,N_29567);
or UO_1699 (O_1699,N_27868,N_27955);
and UO_1700 (O_1700,N_27097,N_28029);
and UO_1701 (O_1701,N_25981,N_27002);
nor UO_1702 (O_1702,N_26908,N_25581);
nor UO_1703 (O_1703,N_27807,N_26015);
xor UO_1704 (O_1704,N_25325,N_25380);
or UO_1705 (O_1705,N_25136,N_29042);
or UO_1706 (O_1706,N_26331,N_25652);
or UO_1707 (O_1707,N_26674,N_29568);
nor UO_1708 (O_1708,N_28416,N_27644);
nand UO_1709 (O_1709,N_26714,N_28261);
and UO_1710 (O_1710,N_27585,N_26303);
nand UO_1711 (O_1711,N_27799,N_27385);
or UO_1712 (O_1712,N_27455,N_25113);
nand UO_1713 (O_1713,N_28929,N_25648);
nor UO_1714 (O_1714,N_29626,N_29838);
xnor UO_1715 (O_1715,N_27338,N_25685);
and UO_1716 (O_1716,N_27451,N_29515);
nand UO_1717 (O_1717,N_28985,N_29410);
or UO_1718 (O_1718,N_26184,N_25720);
and UO_1719 (O_1719,N_26102,N_29523);
xor UO_1720 (O_1720,N_29874,N_25880);
and UO_1721 (O_1721,N_25781,N_28336);
nand UO_1722 (O_1722,N_28125,N_29941);
or UO_1723 (O_1723,N_29164,N_26686);
or UO_1724 (O_1724,N_26422,N_27034);
nand UO_1725 (O_1725,N_26129,N_25904);
xor UO_1726 (O_1726,N_25446,N_26788);
nor UO_1727 (O_1727,N_25573,N_29455);
and UO_1728 (O_1728,N_25527,N_26472);
nor UO_1729 (O_1729,N_25391,N_25490);
nor UO_1730 (O_1730,N_27620,N_29714);
and UO_1731 (O_1731,N_28632,N_26421);
nand UO_1732 (O_1732,N_29939,N_28303);
nor UO_1733 (O_1733,N_27979,N_28588);
nor UO_1734 (O_1734,N_26243,N_27883);
nor UO_1735 (O_1735,N_25844,N_25842);
and UO_1736 (O_1736,N_29084,N_26151);
nand UO_1737 (O_1737,N_29360,N_28778);
nor UO_1738 (O_1738,N_28501,N_28571);
and UO_1739 (O_1739,N_25281,N_28010);
nor UO_1740 (O_1740,N_27313,N_27454);
nor UO_1741 (O_1741,N_29210,N_27954);
nor UO_1742 (O_1742,N_25382,N_25148);
nor UO_1743 (O_1743,N_26070,N_28543);
nor UO_1744 (O_1744,N_27411,N_29877);
nor UO_1745 (O_1745,N_26026,N_26200);
and UO_1746 (O_1746,N_29155,N_29684);
and UO_1747 (O_1747,N_26774,N_27127);
and UO_1748 (O_1748,N_25683,N_29533);
or UO_1749 (O_1749,N_26156,N_25631);
xnor UO_1750 (O_1750,N_27183,N_29055);
or UO_1751 (O_1751,N_29374,N_26571);
or UO_1752 (O_1752,N_27369,N_25883);
nor UO_1753 (O_1753,N_25790,N_25678);
xnor UO_1754 (O_1754,N_25993,N_28946);
and UO_1755 (O_1755,N_27842,N_29821);
nor UO_1756 (O_1756,N_25107,N_27307);
xnor UO_1757 (O_1757,N_29799,N_26463);
nor UO_1758 (O_1758,N_26445,N_29437);
and UO_1759 (O_1759,N_25087,N_25567);
and UO_1760 (O_1760,N_26253,N_28127);
and UO_1761 (O_1761,N_25795,N_29605);
or UO_1762 (O_1762,N_26705,N_28191);
or UO_1763 (O_1763,N_27632,N_27004);
xnor UO_1764 (O_1764,N_26545,N_29414);
nor UO_1765 (O_1765,N_25143,N_29205);
nor UO_1766 (O_1766,N_25353,N_26738);
or UO_1767 (O_1767,N_26353,N_29494);
nor UO_1768 (O_1768,N_27227,N_28689);
nor UO_1769 (O_1769,N_28542,N_28436);
nor UO_1770 (O_1770,N_28358,N_27057);
or UO_1771 (O_1771,N_28126,N_29850);
nor UO_1772 (O_1772,N_27180,N_29369);
and UO_1773 (O_1773,N_25443,N_25367);
nand UO_1774 (O_1774,N_28758,N_25564);
or UO_1775 (O_1775,N_27552,N_26760);
and UO_1776 (O_1776,N_26481,N_25145);
and UO_1777 (O_1777,N_28846,N_27557);
nand UO_1778 (O_1778,N_28357,N_29720);
nor UO_1779 (O_1779,N_29106,N_27877);
nor UO_1780 (O_1780,N_28108,N_29674);
nor UO_1781 (O_1781,N_29972,N_28039);
or UO_1782 (O_1782,N_29384,N_27223);
xnor UO_1783 (O_1783,N_29211,N_26153);
or UO_1784 (O_1784,N_26938,N_25472);
nor UO_1785 (O_1785,N_25827,N_26968);
or UO_1786 (O_1786,N_28296,N_29934);
nand UO_1787 (O_1787,N_29697,N_25482);
xnor UO_1788 (O_1788,N_26410,N_26515);
nor UO_1789 (O_1789,N_28547,N_29759);
nor UO_1790 (O_1790,N_27983,N_25512);
nand UO_1791 (O_1791,N_26814,N_27120);
nor UO_1792 (O_1792,N_27285,N_25977);
xor UO_1793 (O_1793,N_28769,N_28716);
and UO_1794 (O_1794,N_29162,N_26936);
or UO_1795 (O_1795,N_28782,N_26433);
nand UO_1796 (O_1796,N_25815,N_26382);
or UO_1797 (O_1797,N_25777,N_29989);
nor UO_1798 (O_1798,N_25442,N_27150);
and UO_1799 (O_1799,N_25094,N_27434);
nand UO_1800 (O_1800,N_25743,N_27606);
nand UO_1801 (O_1801,N_25068,N_25406);
nand UO_1802 (O_1802,N_27709,N_27996);
or UO_1803 (O_1803,N_27524,N_29270);
xnor UO_1804 (O_1804,N_29863,N_27615);
nor UO_1805 (O_1805,N_25600,N_26214);
nand UO_1806 (O_1806,N_27317,N_27684);
and UO_1807 (O_1807,N_29701,N_29446);
or UO_1808 (O_1808,N_28996,N_27889);
nand UO_1809 (O_1809,N_27817,N_28007);
or UO_1810 (O_1810,N_26577,N_26164);
nor UO_1811 (O_1811,N_27124,N_25126);
nand UO_1812 (O_1812,N_29852,N_29057);
or UO_1813 (O_1813,N_28648,N_27310);
nor UO_1814 (O_1814,N_27624,N_28128);
xor UO_1815 (O_1815,N_29677,N_25702);
or UO_1816 (O_1816,N_26527,N_27678);
nor UO_1817 (O_1817,N_26033,N_27518);
nand UO_1818 (O_1818,N_26644,N_25165);
or UO_1819 (O_1819,N_29643,N_29398);
nor UO_1820 (O_1820,N_25958,N_25338);
or UO_1821 (O_1821,N_29118,N_29702);
nor UO_1822 (O_1822,N_25557,N_29278);
or UO_1823 (O_1823,N_26766,N_29002);
nand UO_1824 (O_1824,N_28264,N_26574);
and UO_1825 (O_1825,N_25359,N_27921);
and UO_1826 (O_1826,N_29691,N_25780);
xor UO_1827 (O_1827,N_25768,N_26703);
nor UO_1828 (O_1828,N_28163,N_26911);
nor UO_1829 (O_1829,N_25837,N_25110);
nor UO_1830 (O_1830,N_27591,N_29019);
or UO_1831 (O_1831,N_28429,N_25991);
nor UO_1832 (O_1832,N_25109,N_28139);
nor UO_1833 (O_1833,N_29981,N_26580);
or UO_1834 (O_1834,N_28037,N_27225);
nor UO_1835 (O_1835,N_29220,N_27957);
or UO_1836 (O_1836,N_28942,N_29357);
and UO_1837 (O_1837,N_29462,N_27565);
nand UO_1838 (O_1838,N_28378,N_27514);
nor UO_1839 (O_1839,N_27953,N_29372);
nor UO_1840 (O_1840,N_28919,N_28939);
or UO_1841 (O_1841,N_27147,N_29102);
or UO_1842 (O_1842,N_29261,N_25337);
nand UO_1843 (O_1843,N_25377,N_26927);
xor UO_1844 (O_1844,N_27742,N_27316);
or UO_1845 (O_1845,N_26460,N_28494);
nor UO_1846 (O_1846,N_26097,N_25549);
nand UO_1847 (O_1847,N_28666,N_26876);
nor UO_1848 (O_1848,N_26372,N_29922);
nor UO_1849 (O_1849,N_26529,N_28102);
and UO_1850 (O_1850,N_27244,N_28187);
xnor UO_1851 (O_1851,N_25222,N_25834);
nor UO_1852 (O_1852,N_29335,N_27642);
nand UO_1853 (O_1853,N_29006,N_29506);
nor UO_1854 (O_1854,N_25856,N_27432);
or UO_1855 (O_1855,N_28205,N_27536);
xnor UO_1856 (O_1856,N_26548,N_27395);
nand UO_1857 (O_1857,N_27448,N_27099);
or UO_1858 (O_1858,N_26012,N_27461);
or UO_1859 (O_1859,N_26654,N_29490);
nor UO_1860 (O_1860,N_25430,N_28064);
and UO_1861 (O_1861,N_26138,N_28723);
and UO_1862 (O_1862,N_25828,N_28268);
nor UO_1863 (O_1863,N_28857,N_26464);
nand UO_1864 (O_1864,N_26782,N_29489);
or UO_1865 (O_1865,N_26894,N_28926);
xor UO_1866 (O_1866,N_29927,N_27773);
xor UO_1867 (O_1867,N_26284,N_27074);
and UO_1868 (O_1868,N_28805,N_27194);
nand UO_1869 (O_1869,N_27444,N_26393);
nand UO_1870 (O_1870,N_25716,N_26735);
or UO_1871 (O_1871,N_27226,N_29049);
nor UO_1872 (O_1872,N_29100,N_27988);
nand UO_1873 (O_1873,N_25479,N_27077);
nor UO_1874 (O_1874,N_25854,N_28422);
and UO_1875 (O_1875,N_25907,N_25076);
nor UO_1876 (O_1876,N_29230,N_29753);
and UO_1877 (O_1877,N_27025,N_28271);
nand UO_1878 (O_1878,N_26939,N_28166);
nor UO_1879 (O_1879,N_28800,N_26141);
or UO_1880 (O_1880,N_28591,N_25286);
nor UO_1881 (O_1881,N_25474,N_27122);
nand UO_1882 (O_1882,N_25436,N_27093);
and UO_1883 (O_1883,N_26693,N_28297);
nor UO_1884 (O_1884,N_26230,N_28809);
nand UO_1885 (O_1885,N_29392,N_27527);
or UO_1886 (O_1886,N_27812,N_27874);
nor UO_1887 (O_1887,N_27622,N_26920);
nor UO_1888 (O_1888,N_29154,N_29876);
nor UO_1889 (O_1889,N_28561,N_26679);
and UO_1890 (O_1890,N_26086,N_28157);
and UO_1891 (O_1891,N_29429,N_29949);
nor UO_1892 (O_1892,N_27737,N_26973);
nand UO_1893 (O_1893,N_25979,N_27698);
nor UO_1894 (O_1894,N_28074,N_28821);
nor UO_1895 (O_1895,N_27713,N_25598);
nand UO_1896 (O_1896,N_29092,N_28273);
and UO_1897 (O_1897,N_26827,N_27083);
nor UO_1898 (O_1898,N_25526,N_26158);
xnor UO_1899 (O_1899,N_26991,N_26396);
nand UO_1900 (O_1900,N_29729,N_29571);
nor UO_1901 (O_1901,N_25983,N_25216);
nand UO_1902 (O_1902,N_25123,N_29819);
nand UO_1903 (O_1903,N_28152,N_27339);
nor UO_1904 (O_1904,N_29883,N_26013);
nor UO_1905 (O_1905,N_28419,N_28393);
nand UO_1906 (O_1906,N_28674,N_27238);
or UO_1907 (O_1907,N_27551,N_26506);
nand UO_1908 (O_1908,N_26255,N_27819);
nand UO_1909 (O_1909,N_29271,N_28664);
nor UO_1910 (O_1910,N_25159,N_27830);
or UO_1911 (O_1911,N_25493,N_29303);
nand UO_1912 (O_1912,N_26843,N_28394);
and UO_1913 (O_1913,N_27305,N_28306);
nand UO_1914 (O_1914,N_28763,N_26804);
xnor UO_1915 (O_1915,N_26630,N_28043);
or UO_1916 (O_1916,N_27986,N_28788);
nor UO_1917 (O_1917,N_26171,N_28670);
or UO_1918 (O_1918,N_27596,N_26704);
xnor UO_1919 (O_1919,N_28572,N_29756);
nand UO_1920 (O_1920,N_25718,N_28943);
nand UO_1921 (O_1921,N_29501,N_28280);
or UO_1922 (O_1922,N_29067,N_28879);
and UO_1923 (O_1923,N_25097,N_25290);
nand UO_1924 (O_1924,N_27405,N_27928);
and UO_1925 (O_1925,N_27478,N_28530);
nand UO_1926 (O_1926,N_28397,N_28230);
xor UO_1927 (O_1927,N_25890,N_25576);
or UO_1928 (O_1928,N_25947,N_25432);
nand UO_1929 (O_1929,N_28486,N_25029);
or UO_1930 (O_1930,N_28148,N_25119);
nand UO_1931 (O_1931,N_28310,N_25031);
and UO_1932 (O_1932,N_28464,N_25050);
nand UO_1933 (O_1933,N_29460,N_27798);
or UO_1934 (O_1934,N_28796,N_29441);
and UO_1935 (O_1935,N_26665,N_27509);
nor UO_1936 (O_1936,N_27217,N_27256);
xnor UO_1937 (O_1937,N_26144,N_25202);
xnor UO_1938 (O_1938,N_25173,N_25006);
nand UO_1939 (O_1939,N_29009,N_27765);
nor UO_1940 (O_1940,N_29751,N_28083);
or UO_1941 (O_1941,N_29172,N_27657);
and UO_1942 (O_1942,N_27490,N_25242);
and UO_1943 (O_1943,N_26210,N_26976);
and UO_1944 (O_1944,N_28613,N_29767);
and UO_1945 (O_1945,N_27459,N_27032);
nand UO_1946 (O_1946,N_28300,N_25788);
and UO_1947 (O_1947,N_26163,N_25749);
nand UO_1948 (O_1948,N_28520,N_29048);
nor UO_1949 (O_1949,N_25304,N_28401);
nor UO_1950 (O_1950,N_27039,N_29302);
nor UO_1951 (O_1951,N_27016,N_25469);
nand UO_1952 (O_1952,N_26486,N_27769);
nand UO_1953 (O_1953,N_28330,N_26985);
nor UO_1954 (O_1954,N_26172,N_25070);
nor UO_1955 (O_1955,N_28186,N_28405);
and UO_1956 (O_1956,N_26528,N_27498);
xor UO_1957 (O_1957,N_27559,N_27211);
nand UO_1958 (O_1958,N_25696,N_28777);
nand UO_1959 (O_1959,N_25273,N_28829);
nand UO_1960 (O_1960,N_28495,N_26249);
nor UO_1961 (O_1961,N_27892,N_25048);
nor UO_1962 (O_1962,N_28815,N_26337);
nand UO_1963 (O_1963,N_29908,N_29673);
nand UO_1964 (O_1964,N_28318,N_25593);
or UO_1965 (O_1965,N_29129,N_27158);
or UO_1966 (O_1966,N_26510,N_28118);
and UO_1967 (O_1967,N_27966,N_26632);
or UO_1968 (O_1968,N_29047,N_28581);
or UO_1969 (O_1969,N_26596,N_26480);
or UO_1970 (O_1970,N_28386,N_25656);
nand UO_1971 (O_1971,N_28267,N_28468);
or UO_1972 (O_1972,N_27259,N_27586);
nor UO_1973 (O_1973,N_28586,N_29453);
nor UO_1974 (O_1974,N_28365,N_26719);
and UO_1975 (O_1975,N_27229,N_29320);
xnor UO_1976 (O_1976,N_25485,N_27627);
and UO_1977 (O_1977,N_25403,N_28751);
nand UO_1978 (O_1978,N_26540,N_26758);
or UO_1979 (O_1979,N_26223,N_25522);
and UO_1980 (O_1980,N_25358,N_27086);
and UO_1981 (O_1981,N_29337,N_26082);
and UO_1982 (O_1982,N_29293,N_25332);
xnor UO_1983 (O_1983,N_29066,N_25873);
nor UO_1984 (O_1984,N_26940,N_29265);
or UO_1985 (O_1985,N_27519,N_29507);
or UO_1986 (O_1986,N_28044,N_29508);
nand UO_1987 (O_1987,N_25735,N_25318);
and UO_1988 (O_1988,N_28961,N_28051);
nand UO_1989 (O_1989,N_29854,N_27797);
nor UO_1990 (O_1990,N_25519,N_29116);
nor UO_1991 (O_1991,N_26073,N_26874);
xnor UO_1992 (O_1992,N_28202,N_25787);
xnor UO_1993 (O_1993,N_29178,N_27681);
or UO_1994 (O_1994,N_26088,N_27361);
nand UO_1995 (O_1995,N_26132,N_25663);
nor UO_1996 (O_1996,N_28366,N_28158);
and UO_1997 (O_1997,N_28329,N_28183);
and UO_1998 (O_1998,N_28253,N_29080);
nand UO_1999 (O_1999,N_29742,N_28452);
and UO_2000 (O_2000,N_26509,N_29052);
and UO_2001 (O_2001,N_28990,N_28917);
and UO_2002 (O_2002,N_27254,N_27095);
or UO_2003 (O_2003,N_26219,N_25799);
and UO_2004 (O_2004,N_28407,N_29358);
and UO_2005 (O_2005,N_27228,N_26142);
nand UO_2006 (O_2006,N_25546,N_28291);
and UO_2007 (O_2007,N_26320,N_29977);
and UO_2008 (O_2008,N_27584,N_27301);
nor UO_2009 (O_2009,N_29316,N_27388);
nor UO_2010 (O_2010,N_26267,N_29161);
or UO_2011 (O_2011,N_27268,N_29077);
nor UO_2012 (O_2012,N_29119,N_25129);
or UO_2013 (O_2013,N_27379,N_25957);
or UO_2014 (O_2014,N_25476,N_27964);
nor UO_2015 (O_2015,N_27712,N_26989);
xnor UO_2016 (O_2016,N_25417,N_28882);
nor UO_2017 (O_2017,N_27210,N_29423);
nor UO_2018 (O_2018,N_27873,N_27779);
or UO_2019 (O_2019,N_29151,N_25054);
xnor UO_2020 (O_2020,N_25709,N_28753);
nand UO_2021 (O_2021,N_26926,N_27855);
nand UO_2022 (O_2022,N_28012,N_28709);
nand UO_2023 (O_2023,N_29287,N_26275);
or UO_2024 (O_2024,N_27003,N_25284);
and UO_2025 (O_2025,N_27246,N_26710);
and UO_2026 (O_2026,N_25810,N_27191);
nor UO_2027 (O_2027,N_26196,N_26706);
or UO_2028 (O_2028,N_29383,N_25821);
or UO_2029 (O_2029,N_25280,N_27061);
and UO_2030 (O_2030,N_27528,N_25945);
or UO_2031 (O_2031,N_29246,N_25995);
xor UO_2032 (O_2032,N_26271,N_29792);
or UO_2033 (O_2033,N_26461,N_29895);
or UO_2034 (O_2034,N_26753,N_27154);
and UO_2035 (O_2035,N_25033,N_26573);
xor UO_2036 (O_2036,N_27546,N_27645);
nor UO_2037 (O_2037,N_27592,N_26482);
nor UO_2038 (O_2038,N_26583,N_26824);
nand UO_2039 (O_2039,N_25934,N_25514);
or UO_2040 (O_2040,N_28078,N_28649);
and UO_2041 (O_2041,N_25754,N_29478);
nand UO_2042 (O_2042,N_25927,N_25997);
xnor UO_2043 (O_2043,N_26306,N_26044);
nor UO_2044 (O_2044,N_28190,N_28539);
nand UO_2045 (O_2045,N_29081,N_25422);
and UO_2046 (O_2046,N_26799,N_28156);
xor UO_2047 (O_2047,N_29656,N_26622);
nor UO_2048 (O_2048,N_27352,N_25627);
and UO_2049 (O_2049,N_26446,N_25264);
and UO_2050 (O_2050,N_28251,N_26447);
or UO_2051 (O_2051,N_25632,N_26595);
or UO_2052 (O_2052,N_28107,N_29375);
or UO_2053 (O_2053,N_27725,N_26101);
nand UO_2054 (O_2054,N_25642,N_27956);
nand UO_2055 (O_2055,N_28451,N_28033);
nor UO_2056 (O_2056,N_26166,N_28013);
nor UO_2057 (O_2057,N_29926,N_26601);
xnor UO_2058 (O_2058,N_28355,N_25552);
nand UO_2059 (O_2059,N_29788,N_29861);
or UO_2060 (O_2060,N_29786,N_28371);
and UO_2061 (O_2061,N_29355,N_27069);
or UO_2062 (O_2062,N_29539,N_28353);
or UO_2063 (O_2063,N_26841,N_26479);
nor UO_2064 (O_2064,N_26687,N_29903);
and UO_2065 (O_2065,N_27362,N_29716);
and UO_2066 (O_2066,N_27356,N_29812);
nand UO_2067 (O_2067,N_27472,N_28991);
and UO_2068 (O_2068,N_26924,N_26597);
nor UO_2069 (O_2069,N_28210,N_27308);
or UO_2070 (O_2070,N_27608,N_27131);
or UO_2071 (O_2071,N_27340,N_27007);
and UO_2072 (O_2072,N_26954,N_29083);
xor UO_2073 (O_2073,N_28550,N_28737);
or UO_2074 (O_2074,N_29236,N_29472);
nor UO_2075 (O_2075,N_26579,N_28121);
xnor UO_2076 (O_2076,N_25862,N_27558);
xnor UO_2077 (O_2077,N_26889,N_26370);
and UO_2078 (O_2078,N_27909,N_25351);
nor UO_2079 (O_2079,N_27162,N_27612);
nor UO_2080 (O_2080,N_25992,N_29504);
or UO_2081 (O_2081,N_28768,N_28423);
or UO_2082 (O_2082,N_26397,N_25471);
nor UO_2083 (O_2083,N_27109,N_29345);
and UO_2084 (O_2084,N_26285,N_25624);
nand UO_2085 (O_2085,N_28430,N_27104);
or UO_2086 (O_2086,N_26754,N_29534);
nor UO_2087 (O_2087,N_25762,N_25190);
or UO_2088 (O_2088,N_28977,N_27279);
nor UO_2089 (O_2089,N_26762,N_26423);
nor UO_2090 (O_2090,N_29791,N_26589);
xor UO_2091 (O_2091,N_28065,N_28826);
nand UO_2092 (O_2092,N_29418,N_28529);
nor UO_2093 (O_2093,N_25954,N_27659);
or UO_2094 (O_2094,N_29806,N_27166);
nor UO_2095 (O_2095,N_29736,N_29910);
nor UO_2096 (O_2096,N_26437,N_29433);
and UO_2097 (O_2097,N_29695,N_27603);
and UO_2098 (O_2098,N_29473,N_26380);
nand UO_2099 (O_2099,N_25896,N_25722);
xnor UO_2100 (O_2100,N_27492,N_27510);
and UO_2101 (O_2101,N_25986,N_28936);
or UO_2102 (O_2102,N_27357,N_27723);
nand UO_2103 (O_2103,N_29942,N_25105);
or UO_2104 (O_2104,N_25630,N_25858);
and UO_2105 (O_2105,N_28161,N_27473);
nand UO_2106 (O_2106,N_26069,N_27736);
nor UO_2107 (O_2107,N_27663,N_26793);
nand UO_2108 (O_2108,N_29435,N_29689);
nand UO_2109 (O_2109,N_28922,N_26450);
nand UO_2110 (O_2110,N_29444,N_28536);
nor UO_2111 (O_2111,N_29897,N_29595);
nand UO_2112 (O_2112,N_29956,N_26418);
nand UO_2113 (O_2113,N_25544,N_28658);
and UO_2114 (O_2114,N_29300,N_27686);
and UO_2115 (O_2115,N_26568,N_28558);
nand UO_2116 (O_2116,N_26663,N_28028);
xor UO_2117 (O_2117,N_25643,N_27813);
nor UO_2118 (O_2118,N_26183,N_27515);
nand UO_2119 (O_2119,N_26036,N_27168);
and UO_2120 (O_2120,N_29772,N_29404);
and UO_2121 (O_2121,N_25069,N_26944);
nand UO_2122 (O_2122,N_25339,N_28552);
or UO_2123 (O_2123,N_25619,N_25690);
or UO_2124 (O_2124,N_26354,N_25879);
and UO_2125 (O_2125,N_29012,N_25350);
nand UO_2126 (O_2126,N_25719,N_25326);
nand UO_2127 (O_2127,N_25169,N_26309);
and UO_2128 (O_2128,N_26429,N_28628);
nor UO_2129 (O_2129,N_25475,N_25209);
xor UO_2130 (O_2130,N_28362,N_25229);
nor UO_2131 (O_2131,N_28784,N_26356);
xnor UO_2132 (O_2132,N_26884,N_25263);
nand UO_2133 (O_2133,N_25331,N_25282);
nand UO_2134 (O_2134,N_26083,N_27598);
nand UO_2135 (O_2135,N_26556,N_28616);
or UO_2136 (O_2136,N_28387,N_28344);
nor UO_2137 (O_2137,N_27137,N_28281);
nand UO_2138 (O_2138,N_29208,N_29010);
nand UO_2139 (O_2139,N_28645,N_26826);
xnor UO_2140 (O_2140,N_27506,N_25577);
xnor UO_2141 (O_2141,N_25116,N_25038);
or UO_2142 (O_2142,N_29060,N_28180);
nand UO_2143 (O_2143,N_25734,N_27782);
nand UO_2144 (O_2144,N_25081,N_27990);
or UO_2145 (O_2145,N_28001,N_27494);
and UO_2146 (O_2146,N_28160,N_28131);
or UO_2147 (O_2147,N_28276,N_27610);
nand UO_2148 (O_2148,N_28162,N_27272);
and UO_2149 (O_2149,N_26702,N_29188);
or UO_2150 (O_2150,N_27359,N_25798);
or UO_2151 (O_2151,N_27425,N_25008);
and UO_2152 (O_2152,N_29735,N_27768);
nand UO_2153 (O_2153,N_29199,N_25072);
nor UO_2154 (O_2154,N_27848,N_29170);
nand UO_2155 (O_2155,N_27101,N_27187);
nor UO_2156 (O_2156,N_28167,N_29371);
xnor UO_2157 (O_2157,N_29132,N_25551);
nor UO_2158 (O_2158,N_29323,N_29112);
and UO_2159 (O_2159,N_27065,N_28172);
or UO_2160 (O_2160,N_26581,N_25866);
or UO_2161 (O_2161,N_29198,N_29645);
nand UO_2162 (O_2162,N_27260,N_27021);
and UO_2163 (O_2163,N_27899,N_27814);
or UO_2164 (O_2164,N_26997,N_29488);
and UO_2165 (O_2165,N_25930,N_28941);
nand UO_2166 (O_2166,N_28736,N_29737);
and UO_2167 (O_2167,N_26668,N_25369);
and UO_2168 (O_2168,N_29126,N_28606);
nand UO_2169 (O_2169,N_27012,N_29847);
and UO_2170 (O_2170,N_29203,N_29875);
xnor UO_2171 (O_2171,N_28449,N_27696);
nand UO_2172 (O_2172,N_29097,N_27441);
nand UO_2173 (O_2173,N_26594,N_25211);
and UO_2174 (O_2174,N_29921,N_29053);
xor UO_2175 (O_2175,N_28855,N_27022);
nor UO_2176 (O_2176,N_27862,N_25487);
or UO_2177 (O_2177,N_26829,N_29319);
and UO_2178 (O_2178,N_27727,N_28269);
nand UO_2179 (O_2179,N_29700,N_29027);
or UO_2180 (O_2180,N_26850,N_29928);
nor UO_2181 (O_2181,N_26299,N_26398);
or UO_2182 (O_2182,N_28969,N_29680);
and UO_2183 (O_2183,N_29841,N_28776);
or UO_2184 (O_2184,N_27984,N_25649);
or UO_2185 (O_2185,N_27580,N_25189);
or UO_2186 (O_2186,N_27529,N_26605);
or UO_2187 (O_2187,N_29978,N_25633);
nand UO_2188 (O_2188,N_29777,N_25538);
nand UO_2189 (O_2189,N_29667,N_26831);
nand UO_2190 (O_2190,N_28400,N_26520);
nor UO_2191 (O_2191,N_27664,N_28927);
nor UO_2192 (O_2192,N_29696,N_25782);
nand UO_2193 (O_2193,N_29040,N_27006);
and UO_2194 (O_2194,N_29886,N_29231);
nor UO_2195 (O_2195,N_27532,N_27261);
and UO_2196 (O_2196,N_25243,N_25058);
or UO_2197 (O_2197,N_25511,N_29026);
or UO_2198 (O_2198,N_29797,N_26053);
nand UO_2199 (O_2199,N_25865,N_29625);
nand UO_2200 (O_2200,N_29818,N_27969);
or UO_2201 (O_2201,N_29273,N_26416);
nor UO_2202 (O_2202,N_28431,N_28621);
nand UO_2203 (O_2203,N_28290,N_29299);
xor UO_2204 (O_2204,N_29624,N_26512);
and UO_2205 (O_2205,N_28383,N_27148);
or UO_2206 (O_2206,N_27929,N_28113);
xor UO_2207 (O_2207,N_29206,N_29608);
nand UO_2208 (O_2208,N_28742,N_26553);
and UO_2209 (O_2209,N_25160,N_26716);
nand UO_2210 (O_2210,N_27375,N_28756);
nor UO_2211 (O_2211,N_26832,N_28610);
nand UO_2212 (O_2212,N_29239,N_28333);
and UO_2213 (O_2213,N_29827,N_25030);
and UO_2214 (O_2214,N_25621,N_28527);
or UO_2215 (O_2215,N_27058,N_28341);
nand UO_2216 (O_2216,N_26980,N_28693);
or UO_2217 (O_2217,N_29324,N_25793);
nor UO_2218 (O_2218,N_26112,N_26269);
or UO_2219 (O_2219,N_28730,N_27277);
nor UO_2220 (O_2220,N_27795,N_25079);
nor UO_2221 (O_2221,N_25245,N_27638);
or UO_2222 (O_2222,N_26969,N_29873);
nor UO_2223 (O_2223,N_25826,N_29993);
and UO_2224 (O_2224,N_28234,N_25531);
nand UO_2225 (O_2225,N_28178,N_25433);
or UO_2226 (O_2226,N_28237,N_27896);
nor UO_2227 (O_2227,N_25363,N_27467);
and UO_2228 (O_2228,N_28424,N_29456);
nor UO_2229 (O_2229,N_29856,N_25438);
nor UO_2230 (O_2230,N_28696,N_25344);
and UO_2231 (O_2231,N_29484,N_25405);
nor UO_2232 (O_2232,N_25288,N_28854);
nand UO_2233 (O_2233,N_27582,N_28573);
nand UO_2234 (O_2234,N_27487,N_27566);
nand UO_2235 (O_2235,N_28492,N_27818);
or UO_2236 (O_2236,N_29820,N_28735);
nand UO_2237 (O_2237,N_29018,N_27750);
nor UO_2238 (O_2238,N_26943,N_26342);
nand UO_2239 (O_2239,N_27044,N_28097);
nor UO_2240 (O_2240,N_26942,N_25629);
and UO_2241 (O_2241,N_28950,N_29063);
or UO_2242 (O_2242,N_25900,N_25599);
and UO_2243 (O_2243,N_29652,N_25346);
nor UO_2244 (O_2244,N_28636,N_26322);
xnor UO_2245 (O_2245,N_27422,N_25542);
or UO_2246 (O_2246,N_25672,N_28911);
xnor UO_2247 (O_2247,N_26030,N_25686);
nor UO_2248 (O_2248,N_28480,N_27333);
and UO_2249 (O_2249,N_27940,N_29718);
nand UO_2250 (O_2250,N_27205,N_28384);
nor UO_2251 (O_2251,N_25276,N_29556);
xor UO_2252 (O_2252,N_28345,N_25171);
nand UO_2253 (O_2253,N_25965,N_28533);
or UO_2254 (O_2254,N_29834,N_29008);
xor UO_2255 (O_2255,N_25231,N_28030);
nand UO_2256 (O_2256,N_28179,N_28745);
nor UO_2257 (O_2257,N_26272,N_29136);
and UO_2258 (O_2258,N_27318,N_27258);
nor UO_2259 (O_2259,N_29880,N_26089);
or UO_2260 (O_2260,N_26897,N_29207);
and UO_2261 (O_2261,N_26308,N_28072);
nand UO_2262 (O_2262,N_29914,N_25466);
and UO_2263 (O_2263,N_28975,N_29001);
and UO_2264 (O_2264,N_28775,N_27911);
nor UO_2265 (O_2265,N_29463,N_27912);
nor UO_2266 (O_2266,N_27772,N_27449);
nor UO_2267 (O_2267,N_27588,N_27445);
or UO_2268 (O_2268,N_27076,N_25206);
nand UO_2269 (O_2269,N_25916,N_29327);
nand UO_2270 (O_2270,N_26765,N_25176);
xor UO_2271 (O_2271,N_28176,N_25982);
or UO_2272 (O_2272,N_28455,N_26204);
nor UO_2273 (O_2273,N_27974,N_25920);
nor UO_2274 (O_2274,N_28521,N_28914);
nor UO_2275 (O_2275,N_26937,N_29461);
or UO_2276 (O_2276,N_29232,N_28812);
or UO_2277 (O_2277,N_28774,N_26008);
and UO_2278 (O_2278,N_29227,N_28877);
xnor UO_2279 (O_2279,N_27630,N_27482);
nor UO_2280 (O_2280,N_25659,N_27575);
and UO_2281 (O_2281,N_25239,N_25611);
and UO_2282 (O_2282,N_25970,N_25509);
xor UO_2283 (O_2283,N_25047,N_28004);
nor UO_2284 (O_2284,N_27167,N_25736);
nand UO_2285 (O_2285,N_26951,N_25915);
nor UO_2286 (O_2286,N_27306,N_27613);
and UO_2287 (O_2287,N_28626,N_29958);
nand UO_2288 (O_2288,N_27155,N_27088);
nor UO_2289 (O_2289,N_27898,N_28389);
and UO_2290 (O_2290,N_26035,N_29237);
nor UO_2291 (O_2291,N_28546,N_25002);
and UO_2292 (O_2292,N_27631,N_25484);
or UO_2293 (O_2293,N_29661,N_27628);
nand UO_2294 (O_2294,N_29629,N_29830);
and UO_2295 (O_2295,N_29722,N_26349);
nand UO_2296 (O_2296,N_28537,N_28892);
xnor UO_2297 (O_2297,N_29125,N_29378);
or UO_2298 (O_2298,N_28482,N_25818);
nor UO_2299 (O_2299,N_26458,N_29353);
nor UO_2300 (O_2300,N_29734,N_27587);
nand UO_2301 (O_2301,N_28201,N_26401);
xor UO_2302 (O_2302,N_29234,N_27549);
and UO_2303 (O_2303,N_28600,N_28481);
or UO_2304 (O_2304,N_26280,N_29251);
and UO_2305 (O_2305,N_28949,N_27732);
nor UO_2306 (O_2306,N_25392,N_28576);
nand UO_2307 (O_2307,N_28989,N_28352);
nor UO_2308 (O_2308,N_27982,N_25961);
or UO_2309 (O_2309,N_25287,N_25838);
nor UO_2310 (O_2310,N_28258,N_27888);
and UO_2311 (O_2311,N_27410,N_26052);
or UO_2312 (O_2312,N_28868,N_29367);
and UO_2313 (O_2313,N_29865,N_26358);
xnor UO_2314 (O_2314,N_25481,N_25831);
nand UO_2315 (O_2315,N_26541,N_28993);
nand UO_2316 (O_2316,N_26886,N_29637);
nand UO_2317 (O_2317,N_26374,N_26122);
nand UO_2318 (O_2318,N_27775,N_28308);
or UO_2319 (O_2319,N_29277,N_28965);
and UO_2320 (O_2320,N_29931,N_27197);
nor UO_2321 (O_2321,N_27399,N_26497);
nand UO_2322 (O_2322,N_27085,N_25269);
xor UO_2323 (O_2323,N_26638,N_28008);
or UO_2324 (O_2324,N_26964,N_27989);
or UO_2325 (O_2325,N_25996,N_28700);
nor UO_2326 (O_2326,N_27617,N_26235);
and UO_2327 (O_2327,N_28893,N_26915);
or UO_2328 (O_2328,N_27469,N_25301);
nand UO_2329 (O_2329,N_28238,N_28968);
and UO_2330 (O_2330,N_29710,N_28263);
and UO_2331 (O_2331,N_29267,N_26851);
and UO_2332 (O_2332,N_26536,N_27084);
xor UO_2333 (O_2333,N_28861,N_29322);
nor UO_2334 (O_2334,N_27548,N_28722);
nor UO_2335 (O_2335,N_25166,N_27520);
or UO_2336 (O_2336,N_27201,N_29552);
nor UO_2337 (O_2337,N_29732,N_26848);
nor UO_2338 (O_2338,N_29752,N_26775);
nand UO_2339 (O_2339,N_28513,N_27675);
xor UO_2340 (O_2340,N_28515,N_25270);
and UO_2341 (O_2341,N_26878,N_27796);
and UO_2342 (O_2342,N_27204,N_25935);
or UO_2343 (O_2343,N_26801,N_29174);
or UO_2344 (O_2344,N_26781,N_28240);
or UO_2345 (O_2345,N_27181,N_26134);
nor UO_2346 (O_2346,N_29306,N_28607);
nor UO_2347 (O_2347,N_25829,N_29779);
xor UO_2348 (O_2348,N_26593,N_29951);
nand UO_2349 (O_2349,N_29544,N_27860);
nand UO_2350 (O_2350,N_25692,N_26139);
nand UO_2351 (O_2351,N_28069,N_27968);
or UO_2352 (O_2352,N_25885,N_27309);
nor UO_2353 (O_2353,N_26149,N_29648);
or UO_2354 (O_2354,N_29741,N_25071);
nor UO_2355 (O_2355,N_25235,N_28377);
and UO_2356 (O_2356,N_26192,N_29853);
and UO_2357 (O_2357,N_26248,N_26325);
nor UO_2358 (O_2358,N_26135,N_27683);
nor UO_2359 (O_2359,N_27428,N_27572);
nand UO_2360 (O_2360,N_28134,N_25093);
nor UO_2361 (O_2361,N_25651,N_27857);
and UO_2362 (O_2362,N_27479,N_26544);
or UO_2363 (O_2363,N_26722,N_28002);
and UO_2364 (O_2364,N_29540,N_29341);
xnor UO_2365 (O_2365,N_28984,N_28055);
nand UO_2366 (O_2366,N_26903,N_27121);
and UO_2367 (O_2367,N_25537,N_25311);
and UO_2368 (O_2368,N_29122,N_28381);
nor UO_2369 (O_2369,N_25039,N_27673);
nand UO_2370 (O_2370,N_25816,N_28831);
nor UO_2371 (O_2371,N_27679,N_28022);
nor UO_2372 (O_2372,N_25300,N_26177);
nor UO_2373 (O_2373,N_26065,N_28767);
xnor UO_2374 (O_2374,N_27704,N_27971);
and UO_2375 (O_2375,N_29778,N_29133);
nand UO_2376 (O_2376,N_27123,N_27908);
and UO_2377 (O_2377,N_26288,N_29108);
or UO_2378 (O_2378,N_27751,N_25425);
or UO_2379 (O_2379,N_26333,N_28052);
nand UO_2380 (O_2380,N_28005,N_29334);
xor UO_2381 (O_2381,N_27231,N_28724);
and UO_2382 (O_2382,N_27337,N_27671);
xor UO_2383 (O_2383,N_25262,N_27828);
nor UO_2384 (O_2384,N_29159,N_28659);
nor UO_2385 (O_2385,N_27015,N_29750);
and UO_2386 (O_2386,N_29721,N_25061);
nor UO_2387 (O_2387,N_28704,N_28242);
nand UO_2388 (O_2388,N_27537,N_29565);
nand UO_2389 (O_2389,N_29004,N_29356);
or UO_2390 (O_2390,N_29421,N_29869);
and UO_2391 (O_2391,N_29707,N_29884);
or UO_2392 (O_2392,N_27271,N_27787);
and UO_2393 (O_2393,N_28448,N_28211);
and UO_2394 (O_2394,N_27826,N_29826);
and UO_2395 (O_2395,N_28059,N_26334);
or UO_2396 (O_2396,N_28392,N_26853);
or UO_2397 (O_2397,N_25168,N_29622);
or UO_2398 (O_2398,N_29072,N_25012);
xor UO_2399 (O_2399,N_29953,N_25817);
or UO_2400 (O_2400,N_28141,N_25876);
nor UO_2401 (O_2401,N_25645,N_25376);
and UO_2402 (O_2402,N_26635,N_25193);
or UO_2403 (O_2403,N_29204,N_27442);
nor UO_2404 (O_2404,N_27447,N_28592);
or UO_2405 (O_2405,N_28856,N_28692);
or UO_2406 (O_2406,N_29272,N_26893);
nor UO_2407 (O_2407,N_29477,N_28457);
and UO_2408 (O_2408,N_29986,N_27143);
and UO_2409 (O_2409,N_28096,N_27178);
and UO_2410 (O_2410,N_26815,N_28637);
xnor UO_2411 (O_2411,N_28073,N_26659);
nor UO_2412 (O_2412,N_29758,N_27739);
or UO_2413 (O_2413,N_27141,N_25536);
or UO_2414 (O_2414,N_25763,N_29362);
or UO_2415 (O_2415,N_28224,N_29840);
or UO_2416 (O_2416,N_26152,N_25592);
nor UO_2417 (O_2417,N_29215,N_27730);
nand UO_2418 (O_2418,N_27066,N_27738);
nor UO_2419 (O_2419,N_26211,N_29180);
or UO_2420 (O_2420,N_26986,N_25019);
and UO_2421 (O_2421,N_27636,N_26341);
nor UO_2422 (O_2422,N_28077,N_29987);
and UO_2423 (O_2423,N_29493,N_26298);
nor UO_2424 (O_2424,N_29566,N_29044);
and UO_2425 (O_2425,N_25812,N_26764);
nand UO_2426 (O_2426,N_25208,N_27561);
and UO_2427 (O_2427,N_29909,N_26996);
and UO_2428 (O_2428,N_26254,N_29054);
nor UO_2429 (O_2429,N_29599,N_26656);
nor UO_2430 (O_2430,N_28835,N_29536);
or UO_2431 (O_2431,N_29495,N_29409);
and UO_2432 (O_2432,N_25182,N_28762);
nand UO_2433 (O_2433,N_25933,N_27522);
nor UO_2434 (O_2434,N_29764,N_29683);
and UO_2435 (O_2435,N_28323,N_25092);
or UO_2436 (O_2436,N_26882,N_25849);
xor UO_2437 (O_2437,N_27611,N_26928);
nor UO_2438 (O_2438,N_25315,N_28888);
nor UO_2439 (O_2439,N_28973,N_29642);
and UO_2440 (O_2440,N_29912,N_27499);
or UO_2441 (O_2441,N_27859,N_26326);
xor UO_2442 (O_2442,N_29663,N_28773);
nand UO_2443 (O_2443,N_26612,N_28862);
or UO_2444 (O_2444,N_25349,N_28379);
nor UO_2445 (O_2445,N_26602,N_29243);
and UO_2446 (O_2446,N_26563,N_25228);
and UO_2447 (O_2447,N_29967,N_25662);
nor UO_2448 (O_2448,N_28066,N_25221);
or UO_2449 (O_2449,N_27791,N_27064);
and UO_2450 (O_2450,N_27325,N_25018);
nand UO_2451 (O_2451,N_28545,N_27710);
or UO_2452 (O_2452,N_25794,N_25396);
nor UO_2453 (O_2453,N_25253,N_25987);
nand UO_2454 (O_2454,N_26619,N_28483);
nor UO_2455 (O_2455,N_25693,N_29275);
or UO_2456 (O_2456,N_29284,N_25679);
nand UO_2457 (O_2457,N_26785,N_26348);
nor UO_2458 (O_2458,N_27035,N_25587);
nor UO_2459 (O_2459,N_29257,N_25172);
and UO_2460 (O_2460,N_27621,N_25370);
and UO_2461 (O_2461,N_27418,N_26966);
and UO_2462 (O_2462,N_29822,N_26819);
or UO_2463 (O_2463,N_29905,N_25064);
nand UO_2464 (O_2464,N_27932,N_29586);
and UO_2465 (O_2465,N_28170,N_25912);
and UO_2466 (O_2466,N_26175,N_29578);
or UO_2467 (O_2467,N_27344,N_26846);
or UO_2468 (O_2468,N_28317,N_29185);
and UO_2469 (O_2469,N_26784,N_29252);
and UO_2470 (O_2470,N_26121,N_29387);
xnor UO_2471 (O_2471,N_28388,N_26883);
or UO_2472 (O_2472,N_29563,N_28023);
nor UO_2473 (O_2473,N_25046,N_29592);
and UO_2474 (O_2474,N_29632,N_29653);
or UO_2475 (O_2475,N_25588,N_26863);
nand UO_2476 (O_2476,N_25308,N_28873);
or UO_2477 (O_2477,N_28803,N_29426);
and UO_2478 (O_2478,N_29687,N_25680);
nor UO_2479 (O_2479,N_25310,N_27533);
xnor UO_2480 (O_2480,N_28320,N_26830);
and UO_2481 (O_2481,N_26133,N_26610);
nand UO_2482 (O_2482,N_25082,N_25650);
or UO_2483 (O_2483,N_26643,N_26818);
nand UO_2484 (O_2484,N_29412,N_28120);
or UO_2485 (O_2485,N_26567,N_29995);
xor UO_2486 (O_2486,N_25708,N_27286);
or UO_2487 (O_2487,N_25021,N_27130);
nand UO_2488 (O_2488,N_25025,N_27556);
xnor UO_2489 (O_2489,N_28239,N_27643);
nor UO_2490 (O_2490,N_28020,N_26700);
nand UO_2491 (O_2491,N_28921,N_27661);
nor UO_2492 (O_2492,N_25625,N_29692);
nor UO_2493 (O_2493,N_25246,N_25773);
nor UO_2494 (O_2494,N_28590,N_27700);
or UO_2495 (O_2495,N_26695,N_25635);
and UO_2496 (O_2496,N_28820,N_27237);
nor UO_2497 (O_2497,N_26324,N_29464);
nor UO_2498 (O_2498,N_28987,N_26417);
nand UO_2499 (O_2499,N_27693,N_25757);
nor UO_2500 (O_2500,N_26024,N_25598);
nand UO_2501 (O_2501,N_25199,N_27079);
xnor UO_2502 (O_2502,N_28808,N_26517);
nand UO_2503 (O_2503,N_25879,N_27419);
nor UO_2504 (O_2504,N_28567,N_25860);
nor UO_2505 (O_2505,N_29856,N_28287);
or UO_2506 (O_2506,N_25794,N_27956);
nor UO_2507 (O_2507,N_29647,N_25878);
or UO_2508 (O_2508,N_25552,N_26674);
or UO_2509 (O_2509,N_26063,N_27805);
nor UO_2510 (O_2510,N_26363,N_26388);
or UO_2511 (O_2511,N_29330,N_28898);
and UO_2512 (O_2512,N_27257,N_26569);
nand UO_2513 (O_2513,N_29144,N_27757);
or UO_2514 (O_2514,N_27796,N_29228);
xnor UO_2515 (O_2515,N_26084,N_28926);
and UO_2516 (O_2516,N_28540,N_29234);
nor UO_2517 (O_2517,N_25924,N_29642);
nand UO_2518 (O_2518,N_26893,N_28593);
or UO_2519 (O_2519,N_28217,N_26920);
and UO_2520 (O_2520,N_28706,N_29777);
xor UO_2521 (O_2521,N_25482,N_27500);
or UO_2522 (O_2522,N_29593,N_28183);
nand UO_2523 (O_2523,N_28382,N_29308);
or UO_2524 (O_2524,N_26110,N_25341);
or UO_2525 (O_2525,N_26666,N_26165);
nor UO_2526 (O_2526,N_27145,N_29894);
and UO_2527 (O_2527,N_26299,N_29317);
or UO_2528 (O_2528,N_25807,N_25500);
nand UO_2529 (O_2529,N_26370,N_28448);
nand UO_2530 (O_2530,N_25485,N_28788);
nor UO_2531 (O_2531,N_27772,N_26059);
nand UO_2532 (O_2532,N_25762,N_28369);
or UO_2533 (O_2533,N_27678,N_27878);
and UO_2534 (O_2534,N_26489,N_28406);
nor UO_2535 (O_2535,N_29559,N_25238);
nand UO_2536 (O_2536,N_27786,N_25001);
nand UO_2537 (O_2537,N_25235,N_27407);
xnor UO_2538 (O_2538,N_28926,N_28813);
and UO_2539 (O_2539,N_27046,N_29227);
nand UO_2540 (O_2540,N_29972,N_25783);
nor UO_2541 (O_2541,N_27626,N_28678);
or UO_2542 (O_2542,N_27510,N_27309);
nand UO_2543 (O_2543,N_25704,N_25549);
and UO_2544 (O_2544,N_28018,N_29450);
nor UO_2545 (O_2545,N_27885,N_26286);
nor UO_2546 (O_2546,N_26107,N_25576);
or UO_2547 (O_2547,N_29588,N_25971);
xor UO_2548 (O_2548,N_29033,N_28586);
nand UO_2549 (O_2549,N_27812,N_27679);
nand UO_2550 (O_2550,N_29132,N_28069);
nor UO_2551 (O_2551,N_28068,N_28346);
nor UO_2552 (O_2552,N_26770,N_25091);
or UO_2553 (O_2553,N_27949,N_25999);
or UO_2554 (O_2554,N_27220,N_26757);
nor UO_2555 (O_2555,N_29048,N_26323);
nand UO_2556 (O_2556,N_26342,N_28887);
nor UO_2557 (O_2557,N_28898,N_25823);
or UO_2558 (O_2558,N_29278,N_28146);
and UO_2559 (O_2559,N_29037,N_28854);
nand UO_2560 (O_2560,N_29934,N_25325);
nand UO_2561 (O_2561,N_27215,N_26436);
and UO_2562 (O_2562,N_27310,N_25519);
or UO_2563 (O_2563,N_26151,N_26083);
nand UO_2564 (O_2564,N_29162,N_29239);
nor UO_2565 (O_2565,N_29938,N_28829);
nor UO_2566 (O_2566,N_26990,N_27824);
xnor UO_2567 (O_2567,N_26880,N_28300);
or UO_2568 (O_2568,N_28531,N_27954);
or UO_2569 (O_2569,N_29299,N_25905);
and UO_2570 (O_2570,N_28123,N_27512);
and UO_2571 (O_2571,N_27133,N_28878);
nor UO_2572 (O_2572,N_26320,N_27156);
xnor UO_2573 (O_2573,N_29994,N_29959);
or UO_2574 (O_2574,N_29494,N_29270);
xor UO_2575 (O_2575,N_27093,N_25820);
and UO_2576 (O_2576,N_27477,N_29045);
nand UO_2577 (O_2577,N_26496,N_28039);
xnor UO_2578 (O_2578,N_28764,N_27381);
and UO_2579 (O_2579,N_27978,N_28101);
nand UO_2580 (O_2580,N_26302,N_29342);
or UO_2581 (O_2581,N_25356,N_28973);
nand UO_2582 (O_2582,N_26486,N_25865);
and UO_2583 (O_2583,N_29713,N_28258);
and UO_2584 (O_2584,N_25241,N_27487);
nand UO_2585 (O_2585,N_26816,N_27955);
or UO_2586 (O_2586,N_29307,N_28608);
nor UO_2587 (O_2587,N_27607,N_25175);
and UO_2588 (O_2588,N_26734,N_29971);
and UO_2589 (O_2589,N_27358,N_28523);
or UO_2590 (O_2590,N_25377,N_27321);
or UO_2591 (O_2591,N_25197,N_28070);
nor UO_2592 (O_2592,N_28247,N_26767);
nand UO_2593 (O_2593,N_29971,N_25562);
and UO_2594 (O_2594,N_27866,N_29483);
and UO_2595 (O_2595,N_25736,N_28525);
nand UO_2596 (O_2596,N_25005,N_26013);
nor UO_2597 (O_2597,N_29410,N_26018);
xor UO_2598 (O_2598,N_27260,N_26716);
nor UO_2599 (O_2599,N_26695,N_25451);
xor UO_2600 (O_2600,N_28290,N_27028);
nand UO_2601 (O_2601,N_28586,N_27243);
nand UO_2602 (O_2602,N_25636,N_26015);
nand UO_2603 (O_2603,N_28808,N_28262);
or UO_2604 (O_2604,N_28737,N_26752);
and UO_2605 (O_2605,N_26904,N_28257);
or UO_2606 (O_2606,N_28964,N_25059);
and UO_2607 (O_2607,N_29594,N_27025);
and UO_2608 (O_2608,N_27565,N_29862);
or UO_2609 (O_2609,N_25695,N_26884);
nor UO_2610 (O_2610,N_29448,N_25754);
or UO_2611 (O_2611,N_27786,N_29553);
and UO_2612 (O_2612,N_28885,N_26865);
nand UO_2613 (O_2613,N_28916,N_25734);
or UO_2614 (O_2614,N_28618,N_29929);
nor UO_2615 (O_2615,N_28365,N_26800);
nor UO_2616 (O_2616,N_27414,N_29448);
and UO_2617 (O_2617,N_28291,N_29144);
and UO_2618 (O_2618,N_25927,N_29229);
and UO_2619 (O_2619,N_25128,N_28027);
nor UO_2620 (O_2620,N_28861,N_25572);
and UO_2621 (O_2621,N_29537,N_29607);
nor UO_2622 (O_2622,N_25708,N_29725);
nor UO_2623 (O_2623,N_28272,N_29384);
nor UO_2624 (O_2624,N_29783,N_26854);
and UO_2625 (O_2625,N_29282,N_25160);
and UO_2626 (O_2626,N_26946,N_27390);
and UO_2627 (O_2627,N_25684,N_28985);
nand UO_2628 (O_2628,N_27915,N_29055);
nand UO_2629 (O_2629,N_25575,N_29801);
or UO_2630 (O_2630,N_26995,N_29289);
or UO_2631 (O_2631,N_26290,N_27904);
or UO_2632 (O_2632,N_29282,N_26703);
or UO_2633 (O_2633,N_25942,N_25871);
or UO_2634 (O_2634,N_28957,N_27029);
and UO_2635 (O_2635,N_27194,N_26958);
nor UO_2636 (O_2636,N_28531,N_27070);
xor UO_2637 (O_2637,N_26123,N_27465);
or UO_2638 (O_2638,N_25797,N_28286);
nand UO_2639 (O_2639,N_28813,N_28904);
nand UO_2640 (O_2640,N_25910,N_29850);
nand UO_2641 (O_2641,N_29947,N_25336);
nor UO_2642 (O_2642,N_26274,N_26082);
nand UO_2643 (O_2643,N_27703,N_26164);
xor UO_2644 (O_2644,N_28628,N_29897);
nand UO_2645 (O_2645,N_27801,N_25326);
nand UO_2646 (O_2646,N_25659,N_29044);
nor UO_2647 (O_2647,N_27801,N_28103);
nand UO_2648 (O_2648,N_29771,N_25726);
and UO_2649 (O_2649,N_26885,N_29303);
and UO_2650 (O_2650,N_28365,N_27608);
or UO_2651 (O_2651,N_25530,N_26649);
nor UO_2652 (O_2652,N_27273,N_28864);
or UO_2653 (O_2653,N_28711,N_25978);
or UO_2654 (O_2654,N_25414,N_26691);
and UO_2655 (O_2655,N_28906,N_26937);
nand UO_2656 (O_2656,N_28210,N_27081);
or UO_2657 (O_2657,N_25796,N_28012);
nand UO_2658 (O_2658,N_27832,N_29946);
or UO_2659 (O_2659,N_25273,N_29946);
nor UO_2660 (O_2660,N_29202,N_28677);
and UO_2661 (O_2661,N_25265,N_26305);
xor UO_2662 (O_2662,N_26858,N_26124);
and UO_2663 (O_2663,N_29866,N_28010);
or UO_2664 (O_2664,N_27019,N_27150);
nor UO_2665 (O_2665,N_28980,N_26217);
or UO_2666 (O_2666,N_25215,N_29398);
and UO_2667 (O_2667,N_28794,N_26037);
nand UO_2668 (O_2668,N_27737,N_26749);
xnor UO_2669 (O_2669,N_26460,N_28891);
nand UO_2670 (O_2670,N_28649,N_28032);
or UO_2671 (O_2671,N_29970,N_27580);
nand UO_2672 (O_2672,N_29850,N_27466);
nand UO_2673 (O_2673,N_26031,N_29944);
and UO_2674 (O_2674,N_28645,N_27941);
nor UO_2675 (O_2675,N_29934,N_28417);
nor UO_2676 (O_2676,N_26165,N_26983);
nor UO_2677 (O_2677,N_28890,N_27135);
nand UO_2678 (O_2678,N_27687,N_28003);
nor UO_2679 (O_2679,N_25180,N_25803);
or UO_2680 (O_2680,N_25027,N_28568);
xor UO_2681 (O_2681,N_28720,N_26133);
and UO_2682 (O_2682,N_29374,N_27946);
xnor UO_2683 (O_2683,N_28157,N_27229);
and UO_2684 (O_2684,N_29735,N_25993);
xor UO_2685 (O_2685,N_28964,N_25695);
nand UO_2686 (O_2686,N_28095,N_25600);
or UO_2687 (O_2687,N_27529,N_26335);
nand UO_2688 (O_2688,N_25175,N_25105);
and UO_2689 (O_2689,N_25781,N_25763);
and UO_2690 (O_2690,N_26789,N_28950);
nand UO_2691 (O_2691,N_28011,N_29436);
and UO_2692 (O_2692,N_25355,N_26151);
and UO_2693 (O_2693,N_26402,N_28707);
nor UO_2694 (O_2694,N_29489,N_25870);
nand UO_2695 (O_2695,N_29147,N_26780);
or UO_2696 (O_2696,N_25606,N_29147);
or UO_2697 (O_2697,N_26945,N_26177);
or UO_2698 (O_2698,N_26051,N_28770);
xnor UO_2699 (O_2699,N_26787,N_28996);
and UO_2700 (O_2700,N_29074,N_29156);
nor UO_2701 (O_2701,N_25210,N_28491);
nor UO_2702 (O_2702,N_29835,N_27986);
xor UO_2703 (O_2703,N_29586,N_26735);
nor UO_2704 (O_2704,N_26354,N_25150);
or UO_2705 (O_2705,N_28424,N_28321);
or UO_2706 (O_2706,N_27665,N_25149);
nor UO_2707 (O_2707,N_25091,N_29271);
or UO_2708 (O_2708,N_25275,N_28106);
nor UO_2709 (O_2709,N_27582,N_27792);
nor UO_2710 (O_2710,N_25021,N_26125);
nand UO_2711 (O_2711,N_28855,N_27322);
nand UO_2712 (O_2712,N_25236,N_25994);
xnor UO_2713 (O_2713,N_29771,N_26123);
or UO_2714 (O_2714,N_29636,N_26329);
and UO_2715 (O_2715,N_26915,N_25745);
and UO_2716 (O_2716,N_26772,N_28416);
nand UO_2717 (O_2717,N_27797,N_29501);
nor UO_2718 (O_2718,N_25813,N_29751);
nand UO_2719 (O_2719,N_27734,N_25741);
xor UO_2720 (O_2720,N_29174,N_29331);
xor UO_2721 (O_2721,N_26815,N_29330);
and UO_2722 (O_2722,N_28426,N_27045);
xnor UO_2723 (O_2723,N_26528,N_29344);
nand UO_2724 (O_2724,N_25184,N_25044);
or UO_2725 (O_2725,N_28940,N_27507);
nor UO_2726 (O_2726,N_27135,N_27634);
nand UO_2727 (O_2727,N_28791,N_29476);
xnor UO_2728 (O_2728,N_26782,N_28245);
and UO_2729 (O_2729,N_28162,N_25584);
and UO_2730 (O_2730,N_28166,N_25448);
nand UO_2731 (O_2731,N_28689,N_25973);
nand UO_2732 (O_2732,N_27758,N_27193);
nand UO_2733 (O_2733,N_25634,N_28115);
nand UO_2734 (O_2734,N_28764,N_25704);
nor UO_2735 (O_2735,N_26248,N_26663);
nand UO_2736 (O_2736,N_26005,N_26625);
nand UO_2737 (O_2737,N_27754,N_26538);
and UO_2738 (O_2738,N_26807,N_26315);
nor UO_2739 (O_2739,N_29073,N_25184);
or UO_2740 (O_2740,N_27114,N_28180);
nand UO_2741 (O_2741,N_27507,N_27325);
nand UO_2742 (O_2742,N_25194,N_27310);
or UO_2743 (O_2743,N_28729,N_26624);
and UO_2744 (O_2744,N_27982,N_25153);
nand UO_2745 (O_2745,N_26399,N_25601);
and UO_2746 (O_2746,N_29440,N_25645);
or UO_2747 (O_2747,N_27526,N_25006);
nand UO_2748 (O_2748,N_29270,N_28498);
xor UO_2749 (O_2749,N_27371,N_29831);
nor UO_2750 (O_2750,N_27218,N_29782);
nor UO_2751 (O_2751,N_26877,N_25009);
xor UO_2752 (O_2752,N_28917,N_26037);
nand UO_2753 (O_2753,N_26988,N_28022);
nand UO_2754 (O_2754,N_29024,N_25963);
or UO_2755 (O_2755,N_25854,N_29513);
nor UO_2756 (O_2756,N_27599,N_28165);
nor UO_2757 (O_2757,N_25402,N_29212);
or UO_2758 (O_2758,N_26245,N_26970);
nand UO_2759 (O_2759,N_26385,N_25457);
and UO_2760 (O_2760,N_29992,N_29430);
nor UO_2761 (O_2761,N_27060,N_26662);
and UO_2762 (O_2762,N_26330,N_29844);
xor UO_2763 (O_2763,N_26725,N_28116);
or UO_2764 (O_2764,N_27827,N_27942);
or UO_2765 (O_2765,N_28319,N_25915);
or UO_2766 (O_2766,N_26814,N_29897);
xnor UO_2767 (O_2767,N_28487,N_27712);
or UO_2768 (O_2768,N_28217,N_28832);
or UO_2769 (O_2769,N_28305,N_29479);
nand UO_2770 (O_2770,N_28671,N_27878);
xor UO_2771 (O_2771,N_25756,N_28369);
and UO_2772 (O_2772,N_26399,N_26976);
or UO_2773 (O_2773,N_28219,N_25752);
nor UO_2774 (O_2774,N_27083,N_27322);
or UO_2775 (O_2775,N_29485,N_28194);
nand UO_2776 (O_2776,N_27290,N_29179);
xnor UO_2777 (O_2777,N_27411,N_29742);
nand UO_2778 (O_2778,N_25934,N_27087);
and UO_2779 (O_2779,N_27202,N_26362);
nand UO_2780 (O_2780,N_28991,N_25309);
nand UO_2781 (O_2781,N_25597,N_27666);
nand UO_2782 (O_2782,N_27291,N_28322);
or UO_2783 (O_2783,N_28346,N_28624);
or UO_2784 (O_2784,N_26431,N_27687);
nand UO_2785 (O_2785,N_26740,N_25875);
nor UO_2786 (O_2786,N_26877,N_29243);
nand UO_2787 (O_2787,N_28315,N_29898);
nand UO_2788 (O_2788,N_25821,N_26377);
and UO_2789 (O_2789,N_29463,N_25371);
and UO_2790 (O_2790,N_28323,N_25001);
or UO_2791 (O_2791,N_27978,N_27814);
nand UO_2792 (O_2792,N_29009,N_27025);
and UO_2793 (O_2793,N_27853,N_29723);
nand UO_2794 (O_2794,N_26091,N_25319);
or UO_2795 (O_2795,N_27465,N_27668);
nor UO_2796 (O_2796,N_28264,N_25613);
nand UO_2797 (O_2797,N_27790,N_26249);
and UO_2798 (O_2798,N_25224,N_25267);
and UO_2799 (O_2799,N_29299,N_26489);
or UO_2800 (O_2800,N_28366,N_27819);
xnor UO_2801 (O_2801,N_25645,N_28870);
and UO_2802 (O_2802,N_28211,N_25504);
nor UO_2803 (O_2803,N_26003,N_27637);
nand UO_2804 (O_2804,N_29343,N_27511);
or UO_2805 (O_2805,N_25374,N_28362);
nand UO_2806 (O_2806,N_29398,N_26281);
or UO_2807 (O_2807,N_28391,N_28223);
and UO_2808 (O_2808,N_29157,N_25749);
nand UO_2809 (O_2809,N_25961,N_29530);
nor UO_2810 (O_2810,N_26831,N_29826);
nor UO_2811 (O_2811,N_27691,N_25991);
xnor UO_2812 (O_2812,N_27332,N_28444);
nor UO_2813 (O_2813,N_28908,N_28972);
nor UO_2814 (O_2814,N_29230,N_27642);
nor UO_2815 (O_2815,N_29257,N_29827);
and UO_2816 (O_2816,N_25262,N_26617);
and UO_2817 (O_2817,N_26300,N_27379);
and UO_2818 (O_2818,N_27218,N_28025);
nor UO_2819 (O_2819,N_28746,N_26608);
and UO_2820 (O_2820,N_28494,N_27226);
or UO_2821 (O_2821,N_27479,N_26242);
or UO_2822 (O_2822,N_25451,N_26063);
xor UO_2823 (O_2823,N_29719,N_25066);
nor UO_2824 (O_2824,N_27751,N_25991);
nor UO_2825 (O_2825,N_26077,N_26574);
nand UO_2826 (O_2826,N_28383,N_27530);
or UO_2827 (O_2827,N_26307,N_26092);
nand UO_2828 (O_2828,N_28658,N_29966);
nor UO_2829 (O_2829,N_25700,N_26279);
nor UO_2830 (O_2830,N_25283,N_28638);
or UO_2831 (O_2831,N_26168,N_28029);
nor UO_2832 (O_2832,N_27563,N_26324);
nand UO_2833 (O_2833,N_26693,N_28166);
nor UO_2834 (O_2834,N_25979,N_29462);
nor UO_2835 (O_2835,N_25386,N_28580);
nand UO_2836 (O_2836,N_25858,N_25160);
nor UO_2837 (O_2837,N_28317,N_27870);
nand UO_2838 (O_2838,N_27511,N_29165);
and UO_2839 (O_2839,N_26410,N_26615);
nand UO_2840 (O_2840,N_28925,N_28431);
nand UO_2841 (O_2841,N_29395,N_29379);
nor UO_2842 (O_2842,N_25027,N_26321);
xor UO_2843 (O_2843,N_25564,N_29793);
or UO_2844 (O_2844,N_28925,N_27257);
and UO_2845 (O_2845,N_28360,N_27394);
nor UO_2846 (O_2846,N_29396,N_25576);
and UO_2847 (O_2847,N_29033,N_25215);
or UO_2848 (O_2848,N_29050,N_26123);
nand UO_2849 (O_2849,N_27291,N_28805);
and UO_2850 (O_2850,N_28035,N_26161);
nor UO_2851 (O_2851,N_27319,N_27709);
xor UO_2852 (O_2852,N_28924,N_25183);
nand UO_2853 (O_2853,N_27720,N_26728);
or UO_2854 (O_2854,N_27595,N_26441);
nand UO_2855 (O_2855,N_29934,N_28663);
or UO_2856 (O_2856,N_27919,N_27013);
and UO_2857 (O_2857,N_27388,N_26625);
nor UO_2858 (O_2858,N_29959,N_26911);
nor UO_2859 (O_2859,N_28471,N_29125);
xnor UO_2860 (O_2860,N_27760,N_26577);
nand UO_2861 (O_2861,N_26015,N_28404);
nor UO_2862 (O_2862,N_27861,N_29890);
nand UO_2863 (O_2863,N_25645,N_29735);
and UO_2864 (O_2864,N_28484,N_27763);
and UO_2865 (O_2865,N_25208,N_25717);
and UO_2866 (O_2866,N_27365,N_27398);
nor UO_2867 (O_2867,N_28149,N_26544);
or UO_2868 (O_2868,N_29251,N_29026);
or UO_2869 (O_2869,N_26475,N_28663);
nand UO_2870 (O_2870,N_29526,N_28593);
and UO_2871 (O_2871,N_27035,N_25398);
or UO_2872 (O_2872,N_25667,N_25291);
nor UO_2873 (O_2873,N_28705,N_29562);
nor UO_2874 (O_2874,N_28266,N_29340);
nand UO_2875 (O_2875,N_25725,N_26272);
nor UO_2876 (O_2876,N_28461,N_28941);
nand UO_2877 (O_2877,N_26387,N_29841);
xor UO_2878 (O_2878,N_26420,N_29594);
nand UO_2879 (O_2879,N_29379,N_29848);
or UO_2880 (O_2880,N_27820,N_28487);
nand UO_2881 (O_2881,N_26130,N_25428);
nand UO_2882 (O_2882,N_26728,N_25862);
and UO_2883 (O_2883,N_25936,N_28244);
nand UO_2884 (O_2884,N_27131,N_27712);
and UO_2885 (O_2885,N_27817,N_26248);
nor UO_2886 (O_2886,N_27369,N_26407);
and UO_2887 (O_2887,N_27979,N_27350);
or UO_2888 (O_2888,N_26183,N_28182);
nand UO_2889 (O_2889,N_28176,N_26457);
nand UO_2890 (O_2890,N_29300,N_27101);
nor UO_2891 (O_2891,N_25307,N_29240);
nor UO_2892 (O_2892,N_29201,N_28605);
or UO_2893 (O_2893,N_26319,N_26694);
and UO_2894 (O_2894,N_29188,N_28431);
nor UO_2895 (O_2895,N_29234,N_26361);
nor UO_2896 (O_2896,N_29869,N_28225);
or UO_2897 (O_2897,N_25010,N_25345);
or UO_2898 (O_2898,N_26800,N_25123);
and UO_2899 (O_2899,N_29990,N_27245);
and UO_2900 (O_2900,N_26347,N_26633);
or UO_2901 (O_2901,N_28808,N_25964);
or UO_2902 (O_2902,N_27581,N_29818);
nand UO_2903 (O_2903,N_28144,N_29499);
and UO_2904 (O_2904,N_26358,N_27114);
or UO_2905 (O_2905,N_25106,N_28059);
and UO_2906 (O_2906,N_28476,N_28757);
nand UO_2907 (O_2907,N_25550,N_26552);
and UO_2908 (O_2908,N_25748,N_27124);
or UO_2909 (O_2909,N_25001,N_26113);
nor UO_2910 (O_2910,N_26373,N_29162);
nor UO_2911 (O_2911,N_26944,N_29958);
or UO_2912 (O_2912,N_26032,N_27371);
xor UO_2913 (O_2913,N_26217,N_27543);
nor UO_2914 (O_2914,N_26058,N_25130);
and UO_2915 (O_2915,N_27700,N_28684);
nand UO_2916 (O_2916,N_25451,N_28726);
nor UO_2917 (O_2917,N_28081,N_28758);
and UO_2918 (O_2918,N_26024,N_26999);
and UO_2919 (O_2919,N_29286,N_29556);
or UO_2920 (O_2920,N_25871,N_26616);
xnor UO_2921 (O_2921,N_28583,N_26021);
xnor UO_2922 (O_2922,N_27676,N_25138);
nand UO_2923 (O_2923,N_29570,N_29659);
nor UO_2924 (O_2924,N_25906,N_25588);
nor UO_2925 (O_2925,N_28270,N_26656);
nand UO_2926 (O_2926,N_25489,N_25032);
xor UO_2927 (O_2927,N_27285,N_25365);
or UO_2928 (O_2928,N_28985,N_27706);
and UO_2929 (O_2929,N_29199,N_25561);
xor UO_2930 (O_2930,N_25234,N_29098);
xnor UO_2931 (O_2931,N_29574,N_29805);
or UO_2932 (O_2932,N_25900,N_27480);
nor UO_2933 (O_2933,N_29156,N_27679);
nor UO_2934 (O_2934,N_27103,N_26698);
or UO_2935 (O_2935,N_28369,N_29003);
nand UO_2936 (O_2936,N_25610,N_29482);
nand UO_2937 (O_2937,N_26035,N_25256);
or UO_2938 (O_2938,N_25648,N_27454);
and UO_2939 (O_2939,N_28848,N_27978);
nor UO_2940 (O_2940,N_28445,N_29767);
nor UO_2941 (O_2941,N_28187,N_28388);
or UO_2942 (O_2942,N_25951,N_28691);
and UO_2943 (O_2943,N_25691,N_29095);
xnor UO_2944 (O_2944,N_29088,N_29487);
xnor UO_2945 (O_2945,N_27192,N_28689);
and UO_2946 (O_2946,N_25277,N_26115);
nand UO_2947 (O_2947,N_25312,N_29280);
or UO_2948 (O_2948,N_26840,N_27960);
xor UO_2949 (O_2949,N_27966,N_27921);
nor UO_2950 (O_2950,N_26138,N_28838);
and UO_2951 (O_2951,N_26371,N_26425);
and UO_2952 (O_2952,N_26431,N_25457);
or UO_2953 (O_2953,N_28367,N_26127);
nor UO_2954 (O_2954,N_29961,N_26456);
nor UO_2955 (O_2955,N_26652,N_27952);
and UO_2956 (O_2956,N_28925,N_26728);
nand UO_2957 (O_2957,N_28179,N_29699);
and UO_2958 (O_2958,N_25101,N_27252);
xor UO_2959 (O_2959,N_26124,N_29114);
or UO_2960 (O_2960,N_25609,N_29652);
and UO_2961 (O_2961,N_25675,N_26463);
nand UO_2962 (O_2962,N_27191,N_29919);
xor UO_2963 (O_2963,N_29412,N_27300);
or UO_2964 (O_2964,N_25730,N_28708);
nor UO_2965 (O_2965,N_25147,N_27929);
or UO_2966 (O_2966,N_27065,N_26477);
or UO_2967 (O_2967,N_26701,N_27977);
nand UO_2968 (O_2968,N_29875,N_26325);
and UO_2969 (O_2969,N_29131,N_27802);
or UO_2970 (O_2970,N_26244,N_27235);
xor UO_2971 (O_2971,N_25196,N_29864);
and UO_2972 (O_2972,N_25959,N_29018);
or UO_2973 (O_2973,N_25654,N_27777);
or UO_2974 (O_2974,N_27651,N_25580);
xnor UO_2975 (O_2975,N_29000,N_29206);
nor UO_2976 (O_2976,N_29665,N_25709);
and UO_2977 (O_2977,N_28806,N_25027);
xor UO_2978 (O_2978,N_25527,N_27652);
and UO_2979 (O_2979,N_29502,N_26740);
or UO_2980 (O_2980,N_28685,N_29703);
nor UO_2981 (O_2981,N_29264,N_26158);
and UO_2982 (O_2982,N_26258,N_28748);
or UO_2983 (O_2983,N_25311,N_26198);
nor UO_2984 (O_2984,N_26835,N_25653);
nor UO_2985 (O_2985,N_25559,N_26177);
nand UO_2986 (O_2986,N_25390,N_27690);
nand UO_2987 (O_2987,N_25302,N_29102);
and UO_2988 (O_2988,N_28839,N_26852);
or UO_2989 (O_2989,N_29614,N_27294);
xor UO_2990 (O_2990,N_28172,N_29127);
and UO_2991 (O_2991,N_25276,N_29376);
and UO_2992 (O_2992,N_29247,N_27119);
or UO_2993 (O_2993,N_25650,N_29903);
and UO_2994 (O_2994,N_25679,N_25756);
nand UO_2995 (O_2995,N_28908,N_27059);
nor UO_2996 (O_2996,N_27386,N_28399);
and UO_2997 (O_2997,N_26641,N_26603);
nor UO_2998 (O_2998,N_28457,N_26936);
xor UO_2999 (O_2999,N_28847,N_28929);
and UO_3000 (O_3000,N_26958,N_25167);
nor UO_3001 (O_3001,N_27788,N_25917);
and UO_3002 (O_3002,N_27172,N_25916);
or UO_3003 (O_3003,N_29718,N_29828);
nand UO_3004 (O_3004,N_27688,N_25408);
nand UO_3005 (O_3005,N_26453,N_25403);
nand UO_3006 (O_3006,N_29219,N_25507);
and UO_3007 (O_3007,N_25691,N_26010);
nand UO_3008 (O_3008,N_29494,N_28118);
or UO_3009 (O_3009,N_29628,N_28849);
xnor UO_3010 (O_3010,N_29730,N_25029);
and UO_3011 (O_3011,N_27750,N_27630);
xnor UO_3012 (O_3012,N_29880,N_26971);
xnor UO_3013 (O_3013,N_29560,N_29593);
nand UO_3014 (O_3014,N_27302,N_28760);
nand UO_3015 (O_3015,N_27538,N_29477);
or UO_3016 (O_3016,N_27236,N_27301);
nand UO_3017 (O_3017,N_26579,N_26581);
nand UO_3018 (O_3018,N_29856,N_27783);
and UO_3019 (O_3019,N_27768,N_25645);
nand UO_3020 (O_3020,N_29810,N_29173);
or UO_3021 (O_3021,N_25534,N_28172);
nand UO_3022 (O_3022,N_26063,N_29976);
and UO_3023 (O_3023,N_29640,N_25791);
and UO_3024 (O_3024,N_26917,N_26368);
and UO_3025 (O_3025,N_29827,N_25225);
nor UO_3026 (O_3026,N_26903,N_27459);
nand UO_3027 (O_3027,N_28597,N_27702);
nand UO_3028 (O_3028,N_25886,N_28299);
nor UO_3029 (O_3029,N_29245,N_26487);
nand UO_3030 (O_3030,N_28363,N_27386);
or UO_3031 (O_3031,N_28247,N_25263);
nor UO_3032 (O_3032,N_27837,N_27171);
nand UO_3033 (O_3033,N_26373,N_27124);
or UO_3034 (O_3034,N_29045,N_28510);
or UO_3035 (O_3035,N_29056,N_28416);
xnor UO_3036 (O_3036,N_26809,N_25287);
or UO_3037 (O_3037,N_27265,N_27175);
nor UO_3038 (O_3038,N_25726,N_26949);
nand UO_3039 (O_3039,N_29800,N_29596);
nor UO_3040 (O_3040,N_26620,N_27996);
nor UO_3041 (O_3041,N_27034,N_29118);
and UO_3042 (O_3042,N_26978,N_29546);
or UO_3043 (O_3043,N_29172,N_29025);
nand UO_3044 (O_3044,N_27784,N_27490);
nand UO_3045 (O_3045,N_25212,N_29069);
xor UO_3046 (O_3046,N_27395,N_29969);
nor UO_3047 (O_3047,N_27723,N_26676);
nand UO_3048 (O_3048,N_25362,N_29870);
and UO_3049 (O_3049,N_28722,N_25693);
and UO_3050 (O_3050,N_26206,N_27966);
nand UO_3051 (O_3051,N_28414,N_27632);
nand UO_3052 (O_3052,N_27445,N_27601);
and UO_3053 (O_3053,N_26467,N_28610);
nand UO_3054 (O_3054,N_27364,N_25873);
and UO_3055 (O_3055,N_29102,N_25198);
and UO_3056 (O_3056,N_29793,N_27746);
xnor UO_3057 (O_3057,N_28291,N_27043);
xnor UO_3058 (O_3058,N_26619,N_25007);
nand UO_3059 (O_3059,N_29607,N_26800);
nor UO_3060 (O_3060,N_26185,N_28083);
or UO_3061 (O_3061,N_26880,N_29646);
nor UO_3062 (O_3062,N_28983,N_29373);
and UO_3063 (O_3063,N_26736,N_26300);
nand UO_3064 (O_3064,N_25500,N_28990);
and UO_3065 (O_3065,N_26663,N_27553);
nor UO_3066 (O_3066,N_26284,N_28654);
nor UO_3067 (O_3067,N_25293,N_28986);
nor UO_3068 (O_3068,N_26948,N_28228);
and UO_3069 (O_3069,N_25035,N_29781);
or UO_3070 (O_3070,N_26117,N_29593);
and UO_3071 (O_3071,N_29689,N_25937);
xnor UO_3072 (O_3072,N_29105,N_29580);
and UO_3073 (O_3073,N_29459,N_29928);
or UO_3074 (O_3074,N_26516,N_29343);
nand UO_3075 (O_3075,N_26878,N_28384);
or UO_3076 (O_3076,N_25584,N_28344);
and UO_3077 (O_3077,N_26855,N_26609);
nor UO_3078 (O_3078,N_28070,N_27750);
or UO_3079 (O_3079,N_29929,N_28688);
nor UO_3080 (O_3080,N_28000,N_29531);
nand UO_3081 (O_3081,N_26299,N_29327);
and UO_3082 (O_3082,N_25345,N_28911);
nor UO_3083 (O_3083,N_26200,N_28637);
or UO_3084 (O_3084,N_25250,N_27557);
or UO_3085 (O_3085,N_27322,N_27607);
nor UO_3086 (O_3086,N_29567,N_29062);
xor UO_3087 (O_3087,N_28999,N_25071);
or UO_3088 (O_3088,N_28426,N_25272);
or UO_3089 (O_3089,N_25905,N_27073);
and UO_3090 (O_3090,N_25764,N_27789);
xor UO_3091 (O_3091,N_26235,N_27451);
xnor UO_3092 (O_3092,N_25358,N_25243);
or UO_3093 (O_3093,N_27057,N_25897);
nor UO_3094 (O_3094,N_25297,N_26197);
xor UO_3095 (O_3095,N_29299,N_27625);
nor UO_3096 (O_3096,N_25389,N_25591);
nand UO_3097 (O_3097,N_28342,N_28468);
nand UO_3098 (O_3098,N_25579,N_25790);
nand UO_3099 (O_3099,N_29303,N_27396);
and UO_3100 (O_3100,N_26354,N_27222);
or UO_3101 (O_3101,N_25514,N_29118);
nand UO_3102 (O_3102,N_26678,N_25458);
nor UO_3103 (O_3103,N_27761,N_28785);
or UO_3104 (O_3104,N_29752,N_28924);
and UO_3105 (O_3105,N_29023,N_26327);
and UO_3106 (O_3106,N_27189,N_26489);
nor UO_3107 (O_3107,N_26204,N_25552);
or UO_3108 (O_3108,N_25343,N_27630);
nor UO_3109 (O_3109,N_25857,N_28469);
nor UO_3110 (O_3110,N_28588,N_27238);
and UO_3111 (O_3111,N_29017,N_25982);
nor UO_3112 (O_3112,N_25730,N_27700);
or UO_3113 (O_3113,N_27477,N_25581);
or UO_3114 (O_3114,N_28715,N_28582);
nand UO_3115 (O_3115,N_26583,N_28772);
and UO_3116 (O_3116,N_27073,N_25714);
and UO_3117 (O_3117,N_27147,N_25856);
or UO_3118 (O_3118,N_28839,N_28910);
nand UO_3119 (O_3119,N_28299,N_27366);
xnor UO_3120 (O_3120,N_27808,N_27310);
or UO_3121 (O_3121,N_26378,N_27572);
nand UO_3122 (O_3122,N_26717,N_28917);
nor UO_3123 (O_3123,N_27014,N_28696);
nor UO_3124 (O_3124,N_29791,N_29134);
and UO_3125 (O_3125,N_26620,N_27445);
nor UO_3126 (O_3126,N_25926,N_25595);
and UO_3127 (O_3127,N_27399,N_27205);
or UO_3128 (O_3128,N_27216,N_27495);
nand UO_3129 (O_3129,N_28592,N_26283);
or UO_3130 (O_3130,N_29673,N_28964);
nor UO_3131 (O_3131,N_25908,N_25105);
nor UO_3132 (O_3132,N_27408,N_27489);
or UO_3133 (O_3133,N_29823,N_26257);
and UO_3134 (O_3134,N_25672,N_27594);
and UO_3135 (O_3135,N_28920,N_25957);
or UO_3136 (O_3136,N_26074,N_26812);
nand UO_3137 (O_3137,N_27994,N_27589);
nand UO_3138 (O_3138,N_29258,N_29025);
or UO_3139 (O_3139,N_26819,N_27157);
and UO_3140 (O_3140,N_27198,N_26153);
nor UO_3141 (O_3141,N_25684,N_26971);
nand UO_3142 (O_3142,N_27836,N_29168);
nand UO_3143 (O_3143,N_25321,N_27554);
and UO_3144 (O_3144,N_27161,N_28663);
or UO_3145 (O_3145,N_28680,N_25121);
nand UO_3146 (O_3146,N_26300,N_27518);
xnor UO_3147 (O_3147,N_25500,N_27043);
nand UO_3148 (O_3148,N_25658,N_29527);
or UO_3149 (O_3149,N_27000,N_25201);
or UO_3150 (O_3150,N_25573,N_29445);
nor UO_3151 (O_3151,N_25917,N_26966);
or UO_3152 (O_3152,N_27268,N_27422);
or UO_3153 (O_3153,N_28970,N_29885);
xnor UO_3154 (O_3154,N_26513,N_27225);
nor UO_3155 (O_3155,N_28284,N_27805);
xnor UO_3156 (O_3156,N_26667,N_28451);
xnor UO_3157 (O_3157,N_27922,N_27206);
nor UO_3158 (O_3158,N_28010,N_29013);
or UO_3159 (O_3159,N_25251,N_29966);
nand UO_3160 (O_3160,N_26870,N_25492);
nor UO_3161 (O_3161,N_27267,N_28099);
and UO_3162 (O_3162,N_28437,N_26628);
nor UO_3163 (O_3163,N_26767,N_29410);
and UO_3164 (O_3164,N_25686,N_25793);
or UO_3165 (O_3165,N_26970,N_28801);
nor UO_3166 (O_3166,N_26288,N_25015);
nand UO_3167 (O_3167,N_26313,N_27295);
nand UO_3168 (O_3168,N_26911,N_29607);
and UO_3169 (O_3169,N_28475,N_25517);
nand UO_3170 (O_3170,N_26238,N_28493);
and UO_3171 (O_3171,N_26397,N_26152);
xnor UO_3172 (O_3172,N_26235,N_28858);
and UO_3173 (O_3173,N_28199,N_25136);
or UO_3174 (O_3174,N_25648,N_27702);
nand UO_3175 (O_3175,N_28799,N_28098);
nand UO_3176 (O_3176,N_29232,N_29576);
or UO_3177 (O_3177,N_29698,N_29979);
nor UO_3178 (O_3178,N_27924,N_25675);
and UO_3179 (O_3179,N_27972,N_29515);
or UO_3180 (O_3180,N_25661,N_25489);
and UO_3181 (O_3181,N_29787,N_25924);
and UO_3182 (O_3182,N_28938,N_28829);
nor UO_3183 (O_3183,N_28887,N_29334);
nor UO_3184 (O_3184,N_25075,N_27586);
xnor UO_3185 (O_3185,N_28490,N_28603);
nor UO_3186 (O_3186,N_25513,N_29107);
and UO_3187 (O_3187,N_28043,N_29909);
nand UO_3188 (O_3188,N_28849,N_27993);
nand UO_3189 (O_3189,N_25817,N_26647);
and UO_3190 (O_3190,N_26287,N_27535);
nor UO_3191 (O_3191,N_26181,N_29976);
nand UO_3192 (O_3192,N_27412,N_29891);
or UO_3193 (O_3193,N_29946,N_29113);
and UO_3194 (O_3194,N_27741,N_28875);
or UO_3195 (O_3195,N_26900,N_25153);
nor UO_3196 (O_3196,N_27274,N_28589);
or UO_3197 (O_3197,N_26536,N_27166);
nor UO_3198 (O_3198,N_25608,N_29458);
nor UO_3199 (O_3199,N_27467,N_25898);
nor UO_3200 (O_3200,N_26942,N_25073);
nand UO_3201 (O_3201,N_29374,N_26747);
nor UO_3202 (O_3202,N_29233,N_29897);
or UO_3203 (O_3203,N_28647,N_29220);
or UO_3204 (O_3204,N_26306,N_29232);
and UO_3205 (O_3205,N_27613,N_26676);
nand UO_3206 (O_3206,N_25680,N_25429);
nor UO_3207 (O_3207,N_29842,N_28263);
nor UO_3208 (O_3208,N_28162,N_28543);
or UO_3209 (O_3209,N_29838,N_26681);
nor UO_3210 (O_3210,N_29538,N_28473);
nor UO_3211 (O_3211,N_26018,N_28667);
nand UO_3212 (O_3212,N_26452,N_26559);
nand UO_3213 (O_3213,N_25438,N_29504);
or UO_3214 (O_3214,N_29806,N_26516);
nor UO_3215 (O_3215,N_29471,N_26590);
or UO_3216 (O_3216,N_26512,N_25117);
or UO_3217 (O_3217,N_25739,N_29114);
xnor UO_3218 (O_3218,N_26380,N_27100);
nand UO_3219 (O_3219,N_29619,N_25160);
nand UO_3220 (O_3220,N_27976,N_29976);
nand UO_3221 (O_3221,N_29317,N_29243);
nor UO_3222 (O_3222,N_29681,N_25570);
and UO_3223 (O_3223,N_26879,N_25992);
or UO_3224 (O_3224,N_26737,N_28312);
or UO_3225 (O_3225,N_26470,N_29338);
nor UO_3226 (O_3226,N_26313,N_26825);
nand UO_3227 (O_3227,N_25979,N_28704);
nor UO_3228 (O_3228,N_28601,N_25587);
nand UO_3229 (O_3229,N_27320,N_28339);
nand UO_3230 (O_3230,N_25538,N_26670);
nor UO_3231 (O_3231,N_29736,N_28777);
or UO_3232 (O_3232,N_26262,N_26119);
nand UO_3233 (O_3233,N_27217,N_27894);
nor UO_3234 (O_3234,N_27171,N_27824);
nand UO_3235 (O_3235,N_25132,N_26014);
and UO_3236 (O_3236,N_26046,N_27998);
nand UO_3237 (O_3237,N_25948,N_28800);
nand UO_3238 (O_3238,N_28706,N_28272);
or UO_3239 (O_3239,N_27104,N_25726);
nand UO_3240 (O_3240,N_25305,N_29785);
nand UO_3241 (O_3241,N_28149,N_29393);
and UO_3242 (O_3242,N_27419,N_25016);
or UO_3243 (O_3243,N_25497,N_25716);
or UO_3244 (O_3244,N_29747,N_26763);
or UO_3245 (O_3245,N_26793,N_25033);
and UO_3246 (O_3246,N_28215,N_26513);
xnor UO_3247 (O_3247,N_27044,N_25259);
and UO_3248 (O_3248,N_29083,N_29713);
xnor UO_3249 (O_3249,N_25524,N_26208);
nor UO_3250 (O_3250,N_27017,N_25007);
nor UO_3251 (O_3251,N_28611,N_28014);
or UO_3252 (O_3252,N_26684,N_25703);
nand UO_3253 (O_3253,N_25923,N_29620);
and UO_3254 (O_3254,N_26546,N_29831);
nand UO_3255 (O_3255,N_25576,N_26416);
and UO_3256 (O_3256,N_28295,N_26973);
and UO_3257 (O_3257,N_27918,N_29774);
nand UO_3258 (O_3258,N_27828,N_29499);
or UO_3259 (O_3259,N_28092,N_29738);
or UO_3260 (O_3260,N_25620,N_29281);
and UO_3261 (O_3261,N_25093,N_28392);
and UO_3262 (O_3262,N_28682,N_25496);
nor UO_3263 (O_3263,N_26119,N_25307);
nand UO_3264 (O_3264,N_28635,N_27097);
xnor UO_3265 (O_3265,N_29257,N_29760);
and UO_3266 (O_3266,N_29257,N_28679);
nor UO_3267 (O_3267,N_28761,N_29552);
nor UO_3268 (O_3268,N_26477,N_29448);
and UO_3269 (O_3269,N_27978,N_26449);
or UO_3270 (O_3270,N_25502,N_28804);
nand UO_3271 (O_3271,N_29815,N_28878);
and UO_3272 (O_3272,N_27922,N_27639);
and UO_3273 (O_3273,N_26315,N_25639);
or UO_3274 (O_3274,N_28798,N_25927);
nand UO_3275 (O_3275,N_26348,N_28098);
and UO_3276 (O_3276,N_25693,N_26342);
or UO_3277 (O_3277,N_28666,N_27531);
nand UO_3278 (O_3278,N_26168,N_28162);
or UO_3279 (O_3279,N_28666,N_26313);
nand UO_3280 (O_3280,N_25782,N_26541);
nand UO_3281 (O_3281,N_29840,N_25342);
or UO_3282 (O_3282,N_26876,N_26056);
and UO_3283 (O_3283,N_29368,N_25972);
nor UO_3284 (O_3284,N_28931,N_26760);
nand UO_3285 (O_3285,N_25637,N_29774);
nand UO_3286 (O_3286,N_26301,N_26098);
nor UO_3287 (O_3287,N_25143,N_28039);
nand UO_3288 (O_3288,N_26023,N_26087);
or UO_3289 (O_3289,N_28950,N_26296);
nand UO_3290 (O_3290,N_27885,N_26955);
nand UO_3291 (O_3291,N_28174,N_29670);
nand UO_3292 (O_3292,N_28736,N_29603);
and UO_3293 (O_3293,N_29427,N_29032);
and UO_3294 (O_3294,N_26781,N_25878);
nand UO_3295 (O_3295,N_29786,N_26344);
and UO_3296 (O_3296,N_27686,N_29411);
or UO_3297 (O_3297,N_25776,N_28210);
and UO_3298 (O_3298,N_27298,N_29629);
nor UO_3299 (O_3299,N_29142,N_25520);
or UO_3300 (O_3300,N_28357,N_26841);
or UO_3301 (O_3301,N_25350,N_26970);
nor UO_3302 (O_3302,N_26550,N_27973);
and UO_3303 (O_3303,N_26624,N_29031);
and UO_3304 (O_3304,N_25038,N_26601);
nor UO_3305 (O_3305,N_25091,N_26928);
nor UO_3306 (O_3306,N_26579,N_28908);
or UO_3307 (O_3307,N_28557,N_25559);
nor UO_3308 (O_3308,N_28760,N_26573);
and UO_3309 (O_3309,N_25011,N_25606);
nand UO_3310 (O_3310,N_25493,N_27697);
nand UO_3311 (O_3311,N_25766,N_28225);
nor UO_3312 (O_3312,N_26880,N_29960);
nor UO_3313 (O_3313,N_29692,N_27514);
or UO_3314 (O_3314,N_28741,N_28839);
nor UO_3315 (O_3315,N_27073,N_27892);
xor UO_3316 (O_3316,N_27961,N_28943);
and UO_3317 (O_3317,N_25151,N_28582);
or UO_3318 (O_3318,N_27256,N_26495);
and UO_3319 (O_3319,N_25577,N_27973);
and UO_3320 (O_3320,N_28477,N_27224);
or UO_3321 (O_3321,N_27766,N_29991);
and UO_3322 (O_3322,N_27626,N_27432);
or UO_3323 (O_3323,N_27783,N_27341);
xor UO_3324 (O_3324,N_27403,N_25455);
nand UO_3325 (O_3325,N_29503,N_26712);
nand UO_3326 (O_3326,N_25053,N_28585);
or UO_3327 (O_3327,N_29857,N_28739);
nor UO_3328 (O_3328,N_25802,N_25075);
and UO_3329 (O_3329,N_29035,N_25055);
or UO_3330 (O_3330,N_26484,N_26809);
nor UO_3331 (O_3331,N_25525,N_28483);
nor UO_3332 (O_3332,N_28061,N_25368);
nand UO_3333 (O_3333,N_29665,N_28388);
nor UO_3334 (O_3334,N_27744,N_25262);
xnor UO_3335 (O_3335,N_25996,N_28143);
or UO_3336 (O_3336,N_28270,N_26904);
nor UO_3337 (O_3337,N_27972,N_25973);
and UO_3338 (O_3338,N_28965,N_29925);
nor UO_3339 (O_3339,N_25305,N_29816);
xor UO_3340 (O_3340,N_27356,N_27408);
or UO_3341 (O_3341,N_26874,N_25650);
xor UO_3342 (O_3342,N_25672,N_29904);
and UO_3343 (O_3343,N_29826,N_29439);
or UO_3344 (O_3344,N_26285,N_29048);
nand UO_3345 (O_3345,N_27356,N_27864);
nand UO_3346 (O_3346,N_29701,N_28577);
or UO_3347 (O_3347,N_28484,N_26236);
xnor UO_3348 (O_3348,N_27619,N_25446);
or UO_3349 (O_3349,N_28147,N_28723);
nand UO_3350 (O_3350,N_28102,N_27007);
nand UO_3351 (O_3351,N_25767,N_26571);
or UO_3352 (O_3352,N_28735,N_28759);
xnor UO_3353 (O_3353,N_29372,N_27845);
and UO_3354 (O_3354,N_26911,N_28765);
and UO_3355 (O_3355,N_27138,N_25866);
and UO_3356 (O_3356,N_28322,N_26169);
and UO_3357 (O_3357,N_27403,N_28380);
nor UO_3358 (O_3358,N_28857,N_28878);
and UO_3359 (O_3359,N_27636,N_28608);
or UO_3360 (O_3360,N_25613,N_29840);
or UO_3361 (O_3361,N_28191,N_25262);
nor UO_3362 (O_3362,N_29721,N_27401);
nor UO_3363 (O_3363,N_26073,N_26596);
nor UO_3364 (O_3364,N_27946,N_26175);
nor UO_3365 (O_3365,N_28974,N_26068);
or UO_3366 (O_3366,N_27277,N_29356);
and UO_3367 (O_3367,N_26845,N_27506);
xnor UO_3368 (O_3368,N_29608,N_29497);
and UO_3369 (O_3369,N_28593,N_25798);
nand UO_3370 (O_3370,N_28998,N_27339);
nor UO_3371 (O_3371,N_25026,N_26382);
and UO_3372 (O_3372,N_26607,N_25336);
or UO_3373 (O_3373,N_27839,N_25932);
nor UO_3374 (O_3374,N_28329,N_26311);
or UO_3375 (O_3375,N_28285,N_25375);
nor UO_3376 (O_3376,N_25956,N_26433);
and UO_3377 (O_3377,N_25601,N_28158);
and UO_3378 (O_3378,N_29160,N_27510);
nand UO_3379 (O_3379,N_27245,N_25383);
xnor UO_3380 (O_3380,N_28797,N_27715);
nor UO_3381 (O_3381,N_26053,N_28557);
nand UO_3382 (O_3382,N_28197,N_25181);
nand UO_3383 (O_3383,N_28456,N_28732);
nor UO_3384 (O_3384,N_25495,N_25740);
nor UO_3385 (O_3385,N_29375,N_26178);
nand UO_3386 (O_3386,N_27014,N_25410);
nand UO_3387 (O_3387,N_28149,N_28256);
nand UO_3388 (O_3388,N_28433,N_25146);
nor UO_3389 (O_3389,N_26905,N_28388);
and UO_3390 (O_3390,N_28076,N_29762);
or UO_3391 (O_3391,N_29797,N_27592);
and UO_3392 (O_3392,N_28211,N_27544);
nand UO_3393 (O_3393,N_26820,N_25078);
or UO_3394 (O_3394,N_25772,N_28960);
or UO_3395 (O_3395,N_28625,N_29736);
nor UO_3396 (O_3396,N_29127,N_27564);
or UO_3397 (O_3397,N_27624,N_28854);
nand UO_3398 (O_3398,N_25426,N_25703);
nand UO_3399 (O_3399,N_28539,N_26517);
or UO_3400 (O_3400,N_25588,N_26163);
or UO_3401 (O_3401,N_29598,N_25462);
nand UO_3402 (O_3402,N_28489,N_29704);
or UO_3403 (O_3403,N_25400,N_26030);
nor UO_3404 (O_3404,N_27464,N_26199);
nor UO_3405 (O_3405,N_25588,N_29286);
nor UO_3406 (O_3406,N_27120,N_25143);
xnor UO_3407 (O_3407,N_28124,N_28489);
nand UO_3408 (O_3408,N_27800,N_27109);
xnor UO_3409 (O_3409,N_27448,N_25373);
or UO_3410 (O_3410,N_27840,N_29539);
or UO_3411 (O_3411,N_25878,N_27628);
nor UO_3412 (O_3412,N_28686,N_28138);
nand UO_3413 (O_3413,N_26731,N_25961);
or UO_3414 (O_3414,N_25212,N_25498);
nand UO_3415 (O_3415,N_28956,N_28859);
or UO_3416 (O_3416,N_29901,N_26043);
nand UO_3417 (O_3417,N_26688,N_25408);
nor UO_3418 (O_3418,N_27443,N_26536);
and UO_3419 (O_3419,N_28719,N_27880);
nor UO_3420 (O_3420,N_25199,N_27073);
nand UO_3421 (O_3421,N_29731,N_28803);
nor UO_3422 (O_3422,N_28355,N_27151);
or UO_3423 (O_3423,N_29915,N_28889);
and UO_3424 (O_3424,N_29851,N_29052);
nand UO_3425 (O_3425,N_27946,N_28049);
nand UO_3426 (O_3426,N_29886,N_29737);
nand UO_3427 (O_3427,N_25146,N_28661);
nor UO_3428 (O_3428,N_25285,N_25902);
and UO_3429 (O_3429,N_29553,N_25093);
nand UO_3430 (O_3430,N_28314,N_28701);
nor UO_3431 (O_3431,N_25840,N_28964);
or UO_3432 (O_3432,N_27253,N_28060);
nor UO_3433 (O_3433,N_26474,N_29217);
nor UO_3434 (O_3434,N_27296,N_25144);
or UO_3435 (O_3435,N_26309,N_28739);
nand UO_3436 (O_3436,N_27616,N_29258);
and UO_3437 (O_3437,N_28391,N_26499);
nor UO_3438 (O_3438,N_25643,N_28010);
and UO_3439 (O_3439,N_27256,N_29101);
xnor UO_3440 (O_3440,N_28208,N_27892);
nor UO_3441 (O_3441,N_27601,N_29234);
or UO_3442 (O_3442,N_29582,N_29186);
or UO_3443 (O_3443,N_29266,N_25912);
or UO_3444 (O_3444,N_25541,N_28483);
nand UO_3445 (O_3445,N_27554,N_26479);
nand UO_3446 (O_3446,N_25550,N_29747);
or UO_3447 (O_3447,N_25862,N_27617);
or UO_3448 (O_3448,N_27153,N_28445);
and UO_3449 (O_3449,N_27345,N_26348);
xnor UO_3450 (O_3450,N_26928,N_25379);
nand UO_3451 (O_3451,N_28831,N_25752);
or UO_3452 (O_3452,N_27016,N_25373);
xnor UO_3453 (O_3453,N_27940,N_28764);
and UO_3454 (O_3454,N_28656,N_28326);
and UO_3455 (O_3455,N_27350,N_28760);
nand UO_3456 (O_3456,N_25544,N_26230);
and UO_3457 (O_3457,N_27409,N_26908);
and UO_3458 (O_3458,N_29937,N_27548);
nand UO_3459 (O_3459,N_26012,N_29542);
nor UO_3460 (O_3460,N_27541,N_26576);
and UO_3461 (O_3461,N_28438,N_27301);
or UO_3462 (O_3462,N_27842,N_25009);
nor UO_3463 (O_3463,N_26490,N_28458);
nand UO_3464 (O_3464,N_27122,N_28703);
nor UO_3465 (O_3465,N_25182,N_25295);
and UO_3466 (O_3466,N_28937,N_26109);
nor UO_3467 (O_3467,N_29292,N_26421);
xor UO_3468 (O_3468,N_28856,N_28408);
nor UO_3469 (O_3469,N_26313,N_28917);
xor UO_3470 (O_3470,N_27736,N_25671);
nand UO_3471 (O_3471,N_28243,N_29359);
nand UO_3472 (O_3472,N_26557,N_27379);
nor UO_3473 (O_3473,N_29579,N_29330);
nand UO_3474 (O_3474,N_28428,N_27079);
and UO_3475 (O_3475,N_25750,N_27468);
and UO_3476 (O_3476,N_29770,N_26667);
or UO_3477 (O_3477,N_27363,N_29743);
or UO_3478 (O_3478,N_26288,N_25336);
nand UO_3479 (O_3479,N_26418,N_25595);
nor UO_3480 (O_3480,N_29099,N_25661);
and UO_3481 (O_3481,N_27259,N_28790);
nor UO_3482 (O_3482,N_25751,N_26278);
nand UO_3483 (O_3483,N_25050,N_27318);
nand UO_3484 (O_3484,N_26902,N_29657);
or UO_3485 (O_3485,N_25197,N_27466);
nor UO_3486 (O_3486,N_25120,N_27341);
or UO_3487 (O_3487,N_29048,N_28990);
nor UO_3488 (O_3488,N_25517,N_28156);
or UO_3489 (O_3489,N_28305,N_27095);
xor UO_3490 (O_3490,N_26447,N_25917);
nor UO_3491 (O_3491,N_26306,N_28748);
nand UO_3492 (O_3492,N_26826,N_27145);
nand UO_3493 (O_3493,N_28431,N_25950);
and UO_3494 (O_3494,N_28711,N_29043);
nor UO_3495 (O_3495,N_29230,N_25268);
nand UO_3496 (O_3496,N_27378,N_26180);
and UO_3497 (O_3497,N_27526,N_28287);
or UO_3498 (O_3498,N_28625,N_29783);
nand UO_3499 (O_3499,N_27473,N_26134);
endmodule