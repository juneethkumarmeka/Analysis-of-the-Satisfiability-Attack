module basic_500_3000_500_60_levels_1xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_220,In_296);
or U1 (N_1,In_84,In_155);
nand U2 (N_2,In_40,In_79);
and U3 (N_3,In_159,In_483);
and U4 (N_4,In_30,In_490);
nor U5 (N_5,In_131,In_294);
nor U6 (N_6,In_283,In_422);
or U7 (N_7,In_140,In_107);
nand U8 (N_8,In_487,In_417);
or U9 (N_9,In_6,In_161);
nand U10 (N_10,In_254,In_173);
or U11 (N_11,In_177,In_32);
nor U12 (N_12,In_243,In_102);
nor U13 (N_13,In_34,In_89);
nor U14 (N_14,In_150,In_116);
and U15 (N_15,In_394,In_104);
or U16 (N_16,In_337,In_201);
nand U17 (N_17,In_316,In_47);
or U18 (N_18,In_1,In_50);
nor U19 (N_19,In_176,In_48);
xnor U20 (N_20,In_474,In_469);
nor U21 (N_21,In_299,In_330);
or U22 (N_22,In_389,In_54);
and U23 (N_23,In_142,In_251);
or U24 (N_24,In_206,In_308);
nand U25 (N_25,In_278,In_479);
or U26 (N_26,In_314,In_385);
and U27 (N_27,In_402,In_74);
and U28 (N_28,In_309,In_171);
nor U29 (N_29,In_441,In_378);
or U30 (N_30,In_231,In_492);
or U31 (N_31,In_181,In_364);
or U32 (N_32,In_349,In_59);
nor U33 (N_33,In_398,In_331);
or U34 (N_34,In_415,In_27);
nand U35 (N_35,In_383,In_467);
nand U36 (N_36,In_478,In_499);
and U37 (N_37,In_183,In_332);
or U38 (N_38,In_222,In_37);
nor U39 (N_39,In_443,In_285);
nand U40 (N_40,In_120,In_138);
or U41 (N_41,In_65,In_369);
and U42 (N_42,In_93,In_397);
or U43 (N_43,In_117,In_62);
and U44 (N_44,In_444,In_382);
nor U45 (N_45,In_261,In_72);
nor U46 (N_46,In_184,In_212);
nor U47 (N_47,In_286,In_384);
nand U48 (N_48,In_160,In_310);
nor U49 (N_49,In_108,In_192);
and U50 (N_50,In_236,In_36);
or U51 (N_51,In_143,In_46);
or U52 (N_52,In_28,In_247);
nor U53 (N_53,In_260,N_4);
nor U54 (N_54,N_17,In_223);
nand U55 (N_55,In_453,In_434);
nor U56 (N_56,In_421,N_25);
xor U57 (N_57,In_328,In_282);
or U58 (N_58,In_262,In_169);
nor U59 (N_59,In_185,In_439);
nand U60 (N_60,In_127,In_489);
or U61 (N_61,In_227,In_420);
or U62 (N_62,In_114,In_357);
nand U63 (N_63,In_480,In_472);
and U64 (N_64,In_21,In_484);
or U65 (N_65,In_372,In_174);
or U66 (N_66,In_438,In_179);
nand U67 (N_67,In_488,In_284);
nor U68 (N_68,In_313,In_76);
nor U69 (N_69,In_321,In_404);
and U70 (N_70,In_263,In_18);
nand U71 (N_71,In_462,In_256);
nand U72 (N_72,In_187,In_375);
and U73 (N_73,In_23,In_408);
or U74 (N_74,N_30,In_66);
nor U75 (N_75,In_178,In_358);
nand U76 (N_76,In_43,In_210);
nor U77 (N_77,In_344,In_392);
or U78 (N_78,In_9,In_53);
or U79 (N_79,In_39,In_141);
nand U80 (N_80,In_495,In_426);
and U81 (N_81,In_377,In_188);
or U82 (N_82,In_475,In_339);
nor U83 (N_83,In_476,In_7);
nand U84 (N_84,In_352,N_26);
nor U85 (N_85,In_134,In_55);
and U86 (N_86,In_246,N_22);
or U87 (N_87,N_29,In_370);
and U88 (N_88,In_235,In_380);
nor U89 (N_89,In_342,In_355);
or U90 (N_90,In_335,In_306);
nand U91 (N_91,N_46,In_348);
and U92 (N_92,In_58,N_7);
nand U93 (N_93,In_482,In_418);
or U94 (N_94,In_497,In_461);
nor U95 (N_95,In_362,N_27);
or U96 (N_96,In_265,In_468);
nand U97 (N_97,In_80,In_437);
nand U98 (N_98,In_24,In_29);
and U99 (N_99,In_295,In_287);
or U100 (N_100,In_267,N_84);
or U101 (N_101,In_428,In_317);
or U102 (N_102,N_57,N_44);
and U103 (N_103,In_113,In_412);
or U104 (N_104,In_148,In_202);
and U105 (N_105,In_414,N_68);
and U106 (N_106,In_244,N_9);
nor U107 (N_107,In_99,In_360);
or U108 (N_108,In_237,In_407);
and U109 (N_109,In_224,In_153);
nor U110 (N_110,In_145,In_226);
and U111 (N_111,In_471,In_464);
and U112 (N_112,In_106,In_205);
nor U113 (N_113,In_424,N_62);
nor U114 (N_114,In_359,In_351);
nor U115 (N_115,In_406,In_374);
nand U116 (N_116,N_89,In_423);
nand U117 (N_117,In_110,In_111);
and U118 (N_118,In_279,N_71);
or U119 (N_119,In_14,In_356);
and U120 (N_120,In_366,In_92);
nor U121 (N_121,In_290,N_80);
and U122 (N_122,In_242,N_90);
and U123 (N_123,In_60,In_221);
or U124 (N_124,In_388,In_139);
and U125 (N_125,In_368,In_228);
nor U126 (N_126,N_19,In_132);
and U127 (N_127,In_268,In_491);
nand U128 (N_128,In_272,In_191);
nor U129 (N_129,N_51,N_12);
nand U130 (N_130,N_92,In_363);
nand U131 (N_131,N_72,In_238);
nand U132 (N_132,In_22,In_189);
or U133 (N_133,In_97,In_83);
or U134 (N_134,In_301,In_214);
nor U135 (N_135,In_123,In_391);
or U136 (N_136,N_95,In_137);
or U137 (N_137,In_121,In_162);
or U138 (N_138,In_165,In_10);
nand U139 (N_139,In_91,In_190);
nand U140 (N_140,N_59,In_96);
nand U141 (N_141,In_15,In_115);
or U142 (N_142,In_195,In_101);
or U143 (N_143,In_460,N_53);
and U144 (N_144,In_387,N_55);
nand U145 (N_145,In_73,In_56);
nor U146 (N_146,N_15,In_302);
nand U147 (N_147,In_152,In_86);
and U148 (N_148,In_209,N_63);
or U149 (N_149,In_456,N_21);
or U150 (N_150,In_354,In_82);
xor U151 (N_151,In_20,In_304);
and U152 (N_152,N_135,N_77);
or U153 (N_153,In_281,N_3);
and U154 (N_154,N_50,In_225);
and U155 (N_155,In_49,In_31);
and U156 (N_156,In_493,N_112);
or U157 (N_157,In_35,In_449);
nor U158 (N_158,In_186,N_121);
and U159 (N_159,N_1,In_182);
and U160 (N_160,In_130,In_442);
nand U161 (N_161,In_118,N_54);
and U162 (N_162,In_38,In_57);
nand U163 (N_163,N_28,In_95);
and U164 (N_164,N_100,In_250);
nor U165 (N_165,N_134,N_39);
nor U166 (N_166,In_459,N_113);
and U167 (N_167,In_324,In_429);
and U168 (N_168,In_4,N_137);
and U169 (N_169,In_416,N_41);
and U170 (N_170,In_230,In_269);
nand U171 (N_171,In_336,In_255);
or U172 (N_172,In_297,In_11);
nand U173 (N_173,In_87,In_41);
nor U174 (N_174,N_45,In_470);
nand U175 (N_175,N_66,In_240);
or U176 (N_176,In_446,In_19);
nand U177 (N_177,In_291,In_311);
and U178 (N_178,N_60,N_70);
or U179 (N_179,In_419,In_129);
or U180 (N_180,In_447,In_325);
and U181 (N_181,In_253,In_207);
nand U182 (N_182,N_32,N_18);
nor U183 (N_183,In_376,In_180);
xor U184 (N_184,N_82,In_67);
and U185 (N_185,N_52,N_142);
and U186 (N_186,In_373,In_203);
nor U187 (N_187,In_463,In_63);
nor U188 (N_188,N_96,In_413);
or U189 (N_189,N_109,In_498);
nor U190 (N_190,In_194,In_77);
and U191 (N_191,N_97,In_379);
and U192 (N_192,In_300,In_109);
nor U193 (N_193,N_117,N_145);
and U194 (N_194,N_40,N_5);
or U195 (N_195,N_35,In_307);
and U196 (N_196,In_327,In_338);
nor U197 (N_197,In_440,In_425);
nor U198 (N_198,In_346,N_138);
nand U199 (N_199,N_148,N_49);
and U200 (N_200,In_208,In_473);
or U201 (N_201,In_289,In_322);
or U202 (N_202,N_47,In_258);
or U203 (N_203,N_43,N_179);
or U204 (N_204,In_13,N_93);
nor U205 (N_205,In_409,In_275);
nor U206 (N_206,N_76,N_157);
and U207 (N_207,N_159,In_450);
nand U208 (N_208,In_445,N_103);
nor U209 (N_209,In_229,In_26);
and U210 (N_210,In_257,In_241);
or U211 (N_211,In_303,In_167);
nor U212 (N_212,In_193,In_198);
or U213 (N_213,N_10,N_173);
nand U214 (N_214,In_494,In_44);
and U215 (N_215,In_395,N_120);
or U216 (N_216,N_20,N_192);
or U217 (N_217,In_340,N_164);
and U218 (N_218,N_183,N_175);
nor U219 (N_219,N_64,N_86);
or U220 (N_220,In_431,N_67);
nor U221 (N_221,In_103,N_11);
nor U222 (N_222,In_158,In_12);
and U223 (N_223,In_320,In_496);
nand U224 (N_224,In_273,N_136);
nand U225 (N_225,In_100,N_184);
or U226 (N_226,In_51,N_107);
and U227 (N_227,N_8,In_200);
and U228 (N_228,N_31,N_153);
nand U229 (N_229,N_58,In_276);
nand U230 (N_230,N_130,N_126);
nand U231 (N_231,N_176,N_79);
or U232 (N_232,In_170,N_81);
and U233 (N_233,In_410,N_199);
nand U234 (N_234,In_146,In_458);
or U235 (N_235,In_298,N_110);
or U236 (N_236,N_139,N_185);
and U237 (N_237,In_457,N_133);
nor U238 (N_238,In_333,In_319);
and U239 (N_239,In_305,In_293);
or U240 (N_240,In_168,N_85);
nor U241 (N_241,In_135,In_280);
nand U242 (N_242,In_288,In_78);
and U243 (N_243,N_172,In_329);
nand U244 (N_244,In_292,In_216);
nand U245 (N_245,N_13,N_123);
nor U246 (N_246,N_144,In_393);
and U247 (N_247,N_0,N_162);
nand U248 (N_248,N_118,In_52);
or U249 (N_249,In_64,In_334);
nand U250 (N_250,In_433,In_264);
nor U251 (N_251,N_167,In_454);
or U252 (N_252,In_400,In_81);
or U253 (N_253,In_144,N_37);
nor U254 (N_254,N_108,In_390);
and U255 (N_255,In_312,N_216);
nand U256 (N_256,In_218,N_111);
or U257 (N_257,N_132,N_191);
and U258 (N_258,N_200,N_240);
and U259 (N_259,N_61,In_126);
or U260 (N_260,In_259,N_116);
and U261 (N_261,In_133,N_187);
and U262 (N_262,N_170,In_315);
and U263 (N_263,N_160,N_236);
and U264 (N_264,N_226,N_83);
nand U265 (N_265,In_401,N_165);
and U266 (N_266,N_24,N_87);
and U267 (N_267,N_244,N_168);
or U268 (N_268,N_78,In_465);
xnor U269 (N_269,In_481,N_131);
and U270 (N_270,N_114,N_242);
nand U271 (N_271,N_104,In_248);
and U272 (N_272,N_155,N_65);
nand U273 (N_273,N_16,In_75);
nand U274 (N_274,N_188,In_68);
or U275 (N_275,In_452,In_213);
nand U276 (N_276,In_239,N_33);
nand U277 (N_277,In_3,N_231);
or U278 (N_278,In_69,N_237);
nor U279 (N_279,N_189,In_172);
nor U280 (N_280,N_224,In_85);
nor U281 (N_281,N_182,N_180);
xnor U282 (N_282,In_5,In_151);
nand U283 (N_283,N_23,In_71);
nor U284 (N_284,In_234,N_127);
nand U285 (N_285,N_218,In_245);
or U286 (N_286,N_171,In_361);
or U287 (N_287,N_221,In_367);
nor U288 (N_288,In_381,N_143);
nand U289 (N_289,N_248,In_318);
or U290 (N_290,In_403,In_455);
nor U291 (N_291,N_213,N_239);
nor U292 (N_292,In_345,In_0);
or U293 (N_293,In_411,N_234);
nand U294 (N_294,In_270,N_38);
nor U295 (N_295,N_158,In_163);
nor U296 (N_296,In_154,N_219);
nand U297 (N_297,N_220,In_427);
nor U298 (N_298,In_266,In_119);
and U299 (N_299,In_252,N_233);
and U300 (N_300,N_251,In_8);
or U301 (N_301,N_295,N_195);
nand U302 (N_302,N_193,N_285);
or U303 (N_303,In_341,N_250);
nor U304 (N_304,N_150,N_296);
nor U305 (N_305,N_73,N_260);
nand U306 (N_306,N_247,N_297);
and U307 (N_307,N_181,N_299);
nor U308 (N_308,N_101,In_451);
and U309 (N_309,In_196,In_164);
or U310 (N_310,In_347,N_196);
nand U311 (N_311,N_152,N_206);
or U312 (N_312,In_98,In_25);
nor U313 (N_313,N_230,In_486);
nand U314 (N_314,N_258,In_233);
or U315 (N_315,In_136,N_56);
or U316 (N_316,N_278,N_156);
and U317 (N_317,N_245,N_276);
nand U318 (N_318,In_219,N_94);
or U319 (N_319,In_277,N_215);
xor U320 (N_320,N_122,N_163);
nor U321 (N_321,N_253,N_287);
and U322 (N_322,In_42,N_91);
nand U323 (N_323,In_70,N_105);
nand U324 (N_324,N_280,In_112);
and U325 (N_325,N_256,In_166);
nand U326 (N_326,In_353,N_190);
or U327 (N_327,In_430,N_261);
nor U328 (N_328,In_88,In_156);
or U329 (N_329,N_166,N_254);
and U330 (N_330,In_396,N_263);
and U331 (N_331,N_279,N_228);
nor U332 (N_332,In_105,N_194);
and U333 (N_333,N_255,N_262);
nor U334 (N_334,In_211,N_217);
and U335 (N_335,N_284,N_169);
and U336 (N_336,N_214,N_293);
nor U337 (N_337,N_222,N_34);
nor U338 (N_338,N_235,N_161);
nand U339 (N_339,N_2,N_269);
nor U340 (N_340,In_147,In_17);
nor U341 (N_341,N_203,In_232);
nor U342 (N_342,N_128,In_435);
nor U343 (N_343,In_350,N_268);
nand U344 (N_344,N_294,N_281);
and U345 (N_345,N_88,In_45);
nor U346 (N_346,N_177,N_288);
nor U347 (N_347,In_405,N_102);
nand U348 (N_348,N_98,N_291);
nand U349 (N_349,In_371,N_225);
nand U350 (N_350,N_42,N_198);
or U351 (N_351,N_303,N_349);
or U352 (N_352,N_69,N_316);
or U353 (N_353,N_323,In_343);
nand U354 (N_354,N_335,N_266);
and U355 (N_355,N_210,N_312);
nand U356 (N_356,In_90,N_310);
or U357 (N_357,N_274,In_323);
and U358 (N_358,N_207,In_466);
or U359 (N_359,N_331,In_436);
nand U360 (N_360,N_209,N_267);
and U361 (N_361,N_227,In_61);
nor U362 (N_362,N_348,N_325);
and U363 (N_363,N_252,In_33);
nand U364 (N_364,N_106,N_336);
nor U365 (N_365,In_274,N_298);
and U366 (N_366,N_241,In_122);
or U367 (N_367,N_275,N_124);
or U368 (N_368,N_283,N_319);
nor U369 (N_369,N_322,N_115);
or U370 (N_370,In_249,In_215);
and U371 (N_371,N_339,N_334);
nand U372 (N_372,N_201,N_205);
xnor U373 (N_373,N_243,N_304);
or U374 (N_374,N_344,N_6);
and U375 (N_375,N_272,N_202);
and U376 (N_376,N_265,N_277);
and U377 (N_377,N_119,N_308);
or U378 (N_378,N_178,N_282);
nand U379 (N_379,N_74,In_432);
nor U380 (N_380,N_212,In_477);
and U381 (N_381,N_223,N_273);
or U382 (N_382,N_309,N_328);
nor U383 (N_383,N_197,N_264);
or U384 (N_384,N_147,N_307);
and U385 (N_385,N_246,N_338);
nor U386 (N_386,N_301,N_330);
and U387 (N_387,In_16,N_337);
and U388 (N_388,N_300,N_75);
or U389 (N_389,N_332,N_125);
nor U390 (N_390,In_197,N_259);
or U391 (N_391,N_151,N_329);
or U392 (N_392,N_232,In_128);
and U393 (N_393,N_343,In_157);
nor U394 (N_394,N_333,N_306);
nand U395 (N_395,N_174,In_125);
nor U396 (N_396,In_199,N_129);
and U397 (N_397,N_238,N_48);
and U398 (N_398,N_140,N_154);
nand U399 (N_399,N_270,N_346);
nor U400 (N_400,N_383,N_353);
and U401 (N_401,N_378,In_448);
nor U402 (N_402,N_341,N_385);
or U403 (N_403,N_386,N_361);
nor U404 (N_404,N_374,N_204);
nand U405 (N_405,N_320,N_359);
and U406 (N_406,In_386,N_373);
nor U407 (N_407,N_396,N_324);
nor U408 (N_408,N_345,N_141);
nor U409 (N_409,N_292,N_350);
and U410 (N_410,In_175,N_390);
and U411 (N_411,N_372,In_365);
or U412 (N_412,N_211,In_204);
nor U413 (N_413,N_352,In_399);
nand U414 (N_414,N_365,N_355);
nor U415 (N_415,N_286,In_124);
and U416 (N_416,N_229,In_94);
nand U417 (N_417,N_397,N_302);
and U418 (N_418,N_357,N_249);
and U419 (N_419,N_340,N_399);
and U420 (N_420,N_388,In_326);
nor U421 (N_421,N_375,N_389);
nor U422 (N_422,N_354,N_395);
nand U423 (N_423,N_370,N_364);
or U424 (N_424,N_356,N_358);
or U425 (N_425,N_318,N_366);
nand U426 (N_426,N_149,N_381);
nor U427 (N_427,N_311,N_347);
nand U428 (N_428,N_376,N_382);
or U429 (N_429,N_146,N_384);
nor U430 (N_430,N_342,N_257);
and U431 (N_431,In_271,N_186);
nor U432 (N_432,N_391,N_327);
xor U433 (N_433,N_14,N_377);
xnor U434 (N_434,N_380,N_362);
or U435 (N_435,N_367,N_369);
or U436 (N_436,N_314,N_271);
or U437 (N_437,N_36,N_326);
or U438 (N_438,N_290,N_313);
and U439 (N_439,In_2,N_371);
or U440 (N_440,N_379,N_315);
nor U441 (N_441,N_387,N_392);
nor U442 (N_442,N_99,N_360);
xor U443 (N_443,N_305,N_398);
and U444 (N_444,N_394,N_351);
and U445 (N_445,N_363,N_393);
nor U446 (N_446,N_368,In_217);
nor U447 (N_447,In_485,N_321);
or U448 (N_448,N_208,N_289);
nor U449 (N_449,In_149,N_317);
nor U450 (N_450,N_445,N_429);
nand U451 (N_451,N_413,N_406);
nand U452 (N_452,N_407,N_440);
or U453 (N_453,N_412,N_402);
and U454 (N_454,N_443,N_419);
or U455 (N_455,N_435,N_421);
nor U456 (N_456,N_438,N_437);
nand U457 (N_457,N_446,N_439);
or U458 (N_458,N_425,N_444);
and U459 (N_459,N_418,N_420);
nor U460 (N_460,N_422,N_423);
nand U461 (N_461,N_424,N_426);
nand U462 (N_462,N_434,N_448);
and U463 (N_463,N_401,N_431);
nand U464 (N_464,N_404,N_441);
or U465 (N_465,N_400,N_447);
and U466 (N_466,N_436,N_409);
or U467 (N_467,N_405,N_427);
nand U468 (N_468,N_433,N_428);
nor U469 (N_469,N_449,N_403);
nor U470 (N_470,N_414,N_416);
nand U471 (N_471,N_430,N_415);
nand U472 (N_472,N_411,N_417);
and U473 (N_473,N_408,N_442);
nor U474 (N_474,N_432,N_410);
and U475 (N_475,N_419,N_418);
xnor U476 (N_476,N_408,N_424);
xnor U477 (N_477,N_433,N_415);
or U478 (N_478,N_426,N_433);
and U479 (N_479,N_425,N_449);
and U480 (N_480,N_419,N_424);
nor U481 (N_481,N_447,N_415);
nand U482 (N_482,N_410,N_447);
nor U483 (N_483,N_443,N_402);
nand U484 (N_484,N_436,N_423);
or U485 (N_485,N_437,N_427);
nand U486 (N_486,N_427,N_425);
xnor U487 (N_487,N_421,N_401);
nand U488 (N_488,N_448,N_424);
and U489 (N_489,N_448,N_436);
or U490 (N_490,N_443,N_445);
and U491 (N_491,N_438,N_406);
or U492 (N_492,N_408,N_429);
nand U493 (N_493,N_444,N_422);
nor U494 (N_494,N_433,N_414);
and U495 (N_495,N_428,N_431);
nand U496 (N_496,N_403,N_409);
nand U497 (N_497,N_441,N_419);
nor U498 (N_498,N_402,N_430);
nor U499 (N_499,N_432,N_400);
nand U500 (N_500,N_458,N_482);
nor U501 (N_501,N_495,N_461);
and U502 (N_502,N_492,N_471);
and U503 (N_503,N_494,N_497);
nor U504 (N_504,N_491,N_490);
nand U505 (N_505,N_498,N_465);
nand U506 (N_506,N_456,N_484);
and U507 (N_507,N_470,N_463);
and U508 (N_508,N_487,N_493);
or U509 (N_509,N_477,N_462);
and U510 (N_510,N_483,N_457);
nand U511 (N_511,N_452,N_464);
or U512 (N_512,N_455,N_466);
and U513 (N_513,N_473,N_489);
or U514 (N_514,N_476,N_486);
and U515 (N_515,N_451,N_496);
or U516 (N_516,N_454,N_469);
nor U517 (N_517,N_499,N_475);
or U518 (N_518,N_488,N_481);
and U519 (N_519,N_485,N_480);
and U520 (N_520,N_478,N_459);
nor U521 (N_521,N_474,N_479);
and U522 (N_522,N_453,N_468);
nand U523 (N_523,N_460,N_467);
and U524 (N_524,N_450,N_472);
nor U525 (N_525,N_470,N_456);
or U526 (N_526,N_485,N_463);
or U527 (N_527,N_489,N_495);
nor U528 (N_528,N_466,N_497);
or U529 (N_529,N_461,N_471);
nor U530 (N_530,N_498,N_488);
nand U531 (N_531,N_468,N_488);
and U532 (N_532,N_485,N_495);
or U533 (N_533,N_454,N_471);
nor U534 (N_534,N_487,N_479);
nor U535 (N_535,N_479,N_498);
or U536 (N_536,N_454,N_457);
nand U537 (N_537,N_493,N_450);
nor U538 (N_538,N_495,N_459);
nor U539 (N_539,N_477,N_467);
or U540 (N_540,N_487,N_460);
nor U541 (N_541,N_481,N_454);
or U542 (N_542,N_498,N_499);
or U543 (N_543,N_466,N_464);
and U544 (N_544,N_481,N_453);
nor U545 (N_545,N_457,N_455);
nor U546 (N_546,N_490,N_463);
and U547 (N_547,N_450,N_487);
nand U548 (N_548,N_469,N_484);
nand U549 (N_549,N_463,N_455);
nand U550 (N_550,N_514,N_507);
nor U551 (N_551,N_515,N_531);
or U552 (N_552,N_543,N_505);
nor U553 (N_553,N_506,N_541);
nand U554 (N_554,N_509,N_548);
nand U555 (N_555,N_502,N_547);
xnor U556 (N_556,N_532,N_539);
and U557 (N_557,N_546,N_519);
nand U558 (N_558,N_527,N_533);
and U559 (N_559,N_534,N_530);
nor U560 (N_560,N_508,N_549);
or U561 (N_561,N_523,N_537);
nand U562 (N_562,N_544,N_517);
nand U563 (N_563,N_520,N_536);
and U564 (N_564,N_540,N_538);
and U565 (N_565,N_522,N_516);
nand U566 (N_566,N_525,N_545);
nand U567 (N_567,N_513,N_528);
xor U568 (N_568,N_511,N_535);
and U569 (N_569,N_529,N_512);
nand U570 (N_570,N_524,N_542);
nor U571 (N_571,N_526,N_503);
nor U572 (N_572,N_501,N_500);
nand U573 (N_573,N_521,N_510);
nand U574 (N_574,N_518,N_504);
or U575 (N_575,N_535,N_522);
nor U576 (N_576,N_533,N_530);
nand U577 (N_577,N_513,N_502);
nor U578 (N_578,N_511,N_520);
or U579 (N_579,N_538,N_539);
xor U580 (N_580,N_516,N_538);
or U581 (N_581,N_532,N_506);
or U582 (N_582,N_512,N_545);
nand U583 (N_583,N_500,N_545);
or U584 (N_584,N_541,N_520);
nand U585 (N_585,N_508,N_504);
nor U586 (N_586,N_506,N_540);
nand U587 (N_587,N_545,N_524);
or U588 (N_588,N_527,N_548);
nand U589 (N_589,N_540,N_524);
and U590 (N_590,N_522,N_521);
or U591 (N_591,N_517,N_518);
or U592 (N_592,N_521,N_535);
nand U593 (N_593,N_506,N_512);
or U594 (N_594,N_537,N_535);
and U595 (N_595,N_502,N_521);
nand U596 (N_596,N_526,N_544);
or U597 (N_597,N_505,N_507);
xnor U598 (N_598,N_511,N_528);
and U599 (N_599,N_533,N_524);
or U600 (N_600,N_596,N_586);
nor U601 (N_601,N_595,N_564);
nand U602 (N_602,N_592,N_552);
nor U603 (N_603,N_587,N_562);
and U604 (N_604,N_570,N_551);
nand U605 (N_605,N_572,N_584);
nor U606 (N_606,N_556,N_594);
and U607 (N_607,N_588,N_571);
nand U608 (N_608,N_590,N_576);
or U609 (N_609,N_598,N_557);
or U610 (N_610,N_559,N_591);
nand U611 (N_611,N_573,N_599);
nand U612 (N_612,N_555,N_593);
nor U613 (N_613,N_583,N_597);
or U614 (N_614,N_563,N_581);
nand U615 (N_615,N_568,N_569);
xor U616 (N_616,N_558,N_580);
or U617 (N_617,N_553,N_554);
nand U618 (N_618,N_582,N_575);
nand U619 (N_619,N_550,N_574);
nand U620 (N_620,N_567,N_561);
and U621 (N_621,N_577,N_565);
nand U622 (N_622,N_578,N_560);
or U623 (N_623,N_579,N_566);
and U624 (N_624,N_589,N_585);
nand U625 (N_625,N_587,N_591);
nand U626 (N_626,N_582,N_588);
or U627 (N_627,N_555,N_563);
and U628 (N_628,N_582,N_583);
nand U629 (N_629,N_559,N_553);
or U630 (N_630,N_562,N_570);
nor U631 (N_631,N_575,N_591);
nor U632 (N_632,N_594,N_598);
nor U633 (N_633,N_556,N_557);
or U634 (N_634,N_559,N_575);
nand U635 (N_635,N_564,N_570);
or U636 (N_636,N_551,N_561);
or U637 (N_637,N_585,N_594);
nor U638 (N_638,N_563,N_578);
nand U639 (N_639,N_551,N_584);
nor U640 (N_640,N_572,N_561);
nand U641 (N_641,N_573,N_584);
nor U642 (N_642,N_584,N_565);
and U643 (N_643,N_584,N_563);
and U644 (N_644,N_554,N_598);
nor U645 (N_645,N_550,N_566);
nor U646 (N_646,N_590,N_595);
nand U647 (N_647,N_592,N_589);
nor U648 (N_648,N_599,N_568);
nand U649 (N_649,N_578,N_585);
and U650 (N_650,N_621,N_640);
and U651 (N_651,N_631,N_607);
nor U652 (N_652,N_644,N_614);
nand U653 (N_653,N_649,N_629);
nand U654 (N_654,N_613,N_600);
or U655 (N_655,N_622,N_642);
or U656 (N_656,N_602,N_610);
nand U657 (N_657,N_615,N_630);
or U658 (N_658,N_628,N_646);
nand U659 (N_659,N_623,N_601);
and U660 (N_660,N_647,N_626);
nand U661 (N_661,N_632,N_627);
nor U662 (N_662,N_635,N_604);
or U663 (N_663,N_648,N_643);
nand U664 (N_664,N_616,N_609);
nand U665 (N_665,N_608,N_611);
nand U666 (N_666,N_636,N_612);
nand U667 (N_667,N_638,N_625);
or U668 (N_668,N_603,N_641);
nand U669 (N_669,N_645,N_639);
nand U670 (N_670,N_606,N_620);
and U671 (N_671,N_619,N_624);
nand U672 (N_672,N_617,N_618);
and U673 (N_673,N_634,N_605);
nor U674 (N_674,N_637,N_633);
or U675 (N_675,N_632,N_640);
nor U676 (N_676,N_609,N_608);
or U677 (N_677,N_601,N_645);
and U678 (N_678,N_609,N_601);
or U679 (N_679,N_605,N_646);
and U680 (N_680,N_602,N_634);
and U681 (N_681,N_644,N_641);
nor U682 (N_682,N_635,N_613);
nand U683 (N_683,N_613,N_647);
and U684 (N_684,N_641,N_616);
nand U685 (N_685,N_608,N_620);
nand U686 (N_686,N_626,N_644);
or U687 (N_687,N_641,N_643);
and U688 (N_688,N_616,N_631);
nand U689 (N_689,N_612,N_643);
or U690 (N_690,N_633,N_610);
and U691 (N_691,N_625,N_637);
and U692 (N_692,N_602,N_615);
nand U693 (N_693,N_624,N_640);
and U694 (N_694,N_648,N_614);
nand U695 (N_695,N_639,N_621);
or U696 (N_696,N_624,N_621);
or U697 (N_697,N_624,N_631);
nor U698 (N_698,N_628,N_609);
nand U699 (N_699,N_620,N_639);
xnor U700 (N_700,N_662,N_669);
nand U701 (N_701,N_695,N_670);
nand U702 (N_702,N_698,N_667);
or U703 (N_703,N_658,N_664);
or U704 (N_704,N_681,N_659);
nand U705 (N_705,N_651,N_689);
and U706 (N_706,N_676,N_697);
nand U707 (N_707,N_673,N_672);
nand U708 (N_708,N_680,N_686);
nor U709 (N_709,N_654,N_668);
nor U710 (N_710,N_685,N_661);
and U711 (N_711,N_652,N_688);
nand U712 (N_712,N_684,N_675);
or U713 (N_713,N_682,N_683);
and U714 (N_714,N_678,N_671);
or U715 (N_715,N_665,N_694);
nand U716 (N_716,N_655,N_666);
or U717 (N_717,N_692,N_653);
or U718 (N_718,N_690,N_691);
nand U719 (N_719,N_674,N_663);
and U720 (N_720,N_677,N_699);
or U721 (N_721,N_679,N_687);
nand U722 (N_722,N_650,N_657);
nand U723 (N_723,N_656,N_696);
and U724 (N_724,N_693,N_660);
or U725 (N_725,N_660,N_658);
nor U726 (N_726,N_672,N_682);
or U727 (N_727,N_698,N_668);
and U728 (N_728,N_677,N_651);
and U729 (N_729,N_652,N_690);
and U730 (N_730,N_690,N_663);
nor U731 (N_731,N_672,N_675);
nand U732 (N_732,N_695,N_692);
or U733 (N_733,N_659,N_670);
nand U734 (N_734,N_651,N_668);
nand U735 (N_735,N_658,N_681);
or U736 (N_736,N_685,N_657);
or U737 (N_737,N_691,N_667);
nand U738 (N_738,N_665,N_676);
nor U739 (N_739,N_651,N_656);
or U740 (N_740,N_657,N_688);
and U741 (N_741,N_692,N_684);
or U742 (N_742,N_691,N_662);
or U743 (N_743,N_653,N_689);
nor U744 (N_744,N_680,N_695);
and U745 (N_745,N_662,N_656);
nor U746 (N_746,N_696,N_655);
and U747 (N_747,N_694,N_659);
and U748 (N_748,N_697,N_667);
and U749 (N_749,N_678,N_673);
nand U750 (N_750,N_728,N_716);
nand U751 (N_751,N_732,N_735);
and U752 (N_752,N_721,N_705);
or U753 (N_753,N_713,N_714);
or U754 (N_754,N_701,N_727);
nor U755 (N_755,N_718,N_711);
or U756 (N_756,N_702,N_734);
or U757 (N_757,N_715,N_744);
and U758 (N_758,N_740,N_719);
and U759 (N_759,N_738,N_736);
xor U760 (N_760,N_725,N_709);
and U761 (N_761,N_706,N_746);
nor U762 (N_762,N_708,N_737);
nor U763 (N_763,N_748,N_733);
and U764 (N_764,N_745,N_730);
nand U765 (N_765,N_720,N_729);
nor U766 (N_766,N_743,N_710);
and U767 (N_767,N_739,N_742);
or U768 (N_768,N_749,N_741);
and U769 (N_769,N_723,N_700);
or U770 (N_770,N_722,N_707);
and U771 (N_771,N_747,N_703);
or U772 (N_772,N_726,N_712);
nand U773 (N_773,N_724,N_704);
nor U774 (N_774,N_717,N_731);
nor U775 (N_775,N_733,N_717);
or U776 (N_776,N_736,N_706);
and U777 (N_777,N_741,N_701);
nand U778 (N_778,N_700,N_735);
and U779 (N_779,N_737,N_704);
nor U780 (N_780,N_708,N_727);
nor U781 (N_781,N_711,N_710);
xnor U782 (N_782,N_717,N_724);
nor U783 (N_783,N_743,N_733);
nor U784 (N_784,N_738,N_737);
nand U785 (N_785,N_727,N_721);
and U786 (N_786,N_712,N_715);
nand U787 (N_787,N_733,N_706);
nand U788 (N_788,N_738,N_735);
and U789 (N_789,N_720,N_727);
or U790 (N_790,N_725,N_739);
or U791 (N_791,N_734,N_704);
nor U792 (N_792,N_711,N_744);
or U793 (N_793,N_748,N_720);
nand U794 (N_794,N_707,N_738);
nor U795 (N_795,N_739,N_714);
or U796 (N_796,N_731,N_714);
nand U797 (N_797,N_716,N_730);
or U798 (N_798,N_731,N_707);
nand U799 (N_799,N_708,N_702);
or U800 (N_800,N_783,N_788);
nand U801 (N_801,N_779,N_776);
nand U802 (N_802,N_754,N_773);
nand U803 (N_803,N_762,N_787);
nor U804 (N_804,N_785,N_768);
nor U805 (N_805,N_791,N_756);
or U806 (N_806,N_753,N_750);
nor U807 (N_807,N_782,N_755);
or U808 (N_808,N_777,N_763);
nor U809 (N_809,N_784,N_795);
nand U810 (N_810,N_781,N_771);
or U811 (N_811,N_793,N_772);
nor U812 (N_812,N_770,N_775);
xor U813 (N_813,N_799,N_797);
and U814 (N_814,N_798,N_774);
nor U815 (N_815,N_761,N_792);
nand U816 (N_816,N_794,N_764);
or U817 (N_817,N_752,N_766);
nor U818 (N_818,N_751,N_769);
or U819 (N_819,N_789,N_758);
nand U820 (N_820,N_790,N_796);
nand U821 (N_821,N_780,N_757);
or U822 (N_822,N_765,N_760);
and U823 (N_823,N_759,N_767);
nor U824 (N_824,N_778,N_786);
nand U825 (N_825,N_768,N_753);
nand U826 (N_826,N_768,N_793);
and U827 (N_827,N_794,N_782);
nand U828 (N_828,N_796,N_763);
or U829 (N_829,N_788,N_758);
nand U830 (N_830,N_752,N_753);
or U831 (N_831,N_770,N_767);
nor U832 (N_832,N_755,N_791);
or U833 (N_833,N_790,N_781);
nand U834 (N_834,N_759,N_754);
and U835 (N_835,N_781,N_769);
nand U836 (N_836,N_782,N_787);
and U837 (N_837,N_789,N_750);
and U838 (N_838,N_750,N_790);
nand U839 (N_839,N_756,N_784);
or U840 (N_840,N_783,N_787);
nor U841 (N_841,N_791,N_793);
or U842 (N_842,N_752,N_763);
and U843 (N_843,N_795,N_773);
nor U844 (N_844,N_792,N_779);
nor U845 (N_845,N_778,N_755);
and U846 (N_846,N_782,N_788);
nand U847 (N_847,N_760,N_784);
and U848 (N_848,N_781,N_780);
xor U849 (N_849,N_750,N_768);
and U850 (N_850,N_805,N_814);
nor U851 (N_851,N_829,N_847);
nor U852 (N_852,N_816,N_817);
nand U853 (N_853,N_842,N_819);
nand U854 (N_854,N_820,N_809);
and U855 (N_855,N_807,N_846);
and U856 (N_856,N_838,N_833);
xnor U857 (N_857,N_841,N_812);
or U858 (N_858,N_826,N_811);
and U859 (N_859,N_825,N_818);
or U860 (N_860,N_803,N_835);
and U861 (N_861,N_827,N_848);
nand U862 (N_862,N_804,N_810);
or U863 (N_863,N_849,N_830);
or U864 (N_864,N_836,N_834);
and U865 (N_865,N_801,N_843);
nand U866 (N_866,N_815,N_821);
and U867 (N_867,N_840,N_845);
or U868 (N_868,N_832,N_822);
or U869 (N_869,N_824,N_844);
nor U870 (N_870,N_831,N_823);
xor U871 (N_871,N_806,N_837);
nand U872 (N_872,N_802,N_828);
nand U873 (N_873,N_813,N_839);
or U874 (N_874,N_808,N_800);
or U875 (N_875,N_843,N_803);
nand U876 (N_876,N_826,N_830);
nand U877 (N_877,N_805,N_806);
and U878 (N_878,N_838,N_823);
and U879 (N_879,N_825,N_804);
or U880 (N_880,N_839,N_804);
nand U881 (N_881,N_836,N_826);
nor U882 (N_882,N_812,N_807);
nor U883 (N_883,N_823,N_835);
nor U884 (N_884,N_831,N_845);
and U885 (N_885,N_834,N_822);
and U886 (N_886,N_834,N_848);
or U887 (N_887,N_824,N_848);
nor U888 (N_888,N_847,N_819);
nand U889 (N_889,N_833,N_817);
nor U890 (N_890,N_827,N_823);
and U891 (N_891,N_826,N_812);
or U892 (N_892,N_815,N_827);
nor U893 (N_893,N_849,N_821);
and U894 (N_894,N_843,N_826);
nor U895 (N_895,N_816,N_835);
and U896 (N_896,N_818,N_848);
and U897 (N_897,N_846,N_823);
and U898 (N_898,N_814,N_840);
or U899 (N_899,N_846,N_802);
nor U900 (N_900,N_899,N_871);
and U901 (N_901,N_856,N_897);
nor U902 (N_902,N_854,N_864);
and U903 (N_903,N_877,N_891);
or U904 (N_904,N_862,N_890);
nand U905 (N_905,N_855,N_867);
or U906 (N_906,N_888,N_883);
or U907 (N_907,N_868,N_857);
nor U908 (N_908,N_879,N_869);
nor U909 (N_909,N_851,N_892);
or U910 (N_910,N_893,N_852);
and U911 (N_911,N_889,N_860);
nand U912 (N_912,N_873,N_896);
or U913 (N_913,N_884,N_895);
nand U914 (N_914,N_898,N_876);
or U915 (N_915,N_885,N_858);
or U916 (N_916,N_882,N_894);
or U917 (N_917,N_880,N_853);
and U918 (N_918,N_886,N_887);
or U919 (N_919,N_870,N_859);
or U920 (N_920,N_861,N_850);
or U921 (N_921,N_863,N_865);
nor U922 (N_922,N_878,N_881);
nor U923 (N_923,N_866,N_874);
nor U924 (N_924,N_872,N_875);
or U925 (N_925,N_893,N_869);
and U926 (N_926,N_852,N_872);
and U927 (N_927,N_881,N_898);
or U928 (N_928,N_881,N_861);
nor U929 (N_929,N_858,N_886);
nand U930 (N_930,N_867,N_882);
xnor U931 (N_931,N_873,N_855);
nor U932 (N_932,N_850,N_895);
and U933 (N_933,N_856,N_851);
nor U934 (N_934,N_892,N_855);
nor U935 (N_935,N_869,N_892);
nor U936 (N_936,N_898,N_861);
nand U937 (N_937,N_871,N_882);
nor U938 (N_938,N_892,N_895);
nand U939 (N_939,N_869,N_858);
nor U940 (N_940,N_897,N_878);
and U941 (N_941,N_860,N_858);
nor U942 (N_942,N_870,N_875);
nor U943 (N_943,N_873,N_875);
and U944 (N_944,N_888,N_893);
or U945 (N_945,N_874,N_898);
or U946 (N_946,N_858,N_882);
and U947 (N_947,N_855,N_869);
nand U948 (N_948,N_879,N_896);
or U949 (N_949,N_862,N_891);
nand U950 (N_950,N_930,N_932);
or U951 (N_951,N_942,N_919);
nand U952 (N_952,N_900,N_927);
nand U953 (N_953,N_910,N_941);
nand U954 (N_954,N_911,N_913);
or U955 (N_955,N_905,N_938);
nor U956 (N_956,N_922,N_929);
or U957 (N_957,N_907,N_947);
nor U958 (N_958,N_944,N_908);
nand U959 (N_959,N_914,N_901);
and U960 (N_960,N_936,N_917);
nor U961 (N_961,N_935,N_923);
and U962 (N_962,N_924,N_920);
nand U963 (N_963,N_939,N_931);
or U964 (N_964,N_946,N_906);
or U965 (N_965,N_934,N_933);
nand U966 (N_966,N_928,N_925);
and U967 (N_967,N_902,N_916);
nand U968 (N_968,N_918,N_904);
nor U969 (N_969,N_921,N_912);
or U970 (N_970,N_903,N_948);
nand U971 (N_971,N_909,N_943);
and U972 (N_972,N_945,N_926);
or U973 (N_973,N_949,N_940);
and U974 (N_974,N_937,N_915);
or U975 (N_975,N_902,N_943);
or U976 (N_976,N_920,N_923);
nor U977 (N_977,N_907,N_908);
and U978 (N_978,N_913,N_902);
nor U979 (N_979,N_941,N_920);
and U980 (N_980,N_911,N_947);
or U981 (N_981,N_903,N_924);
nand U982 (N_982,N_905,N_917);
nor U983 (N_983,N_916,N_918);
and U984 (N_984,N_940,N_910);
or U985 (N_985,N_938,N_940);
nor U986 (N_986,N_931,N_940);
and U987 (N_987,N_911,N_907);
nand U988 (N_988,N_935,N_922);
or U989 (N_989,N_934,N_931);
and U990 (N_990,N_924,N_917);
nand U991 (N_991,N_912,N_906);
nor U992 (N_992,N_919,N_912);
or U993 (N_993,N_925,N_920);
nand U994 (N_994,N_904,N_942);
nand U995 (N_995,N_904,N_902);
nor U996 (N_996,N_930,N_928);
and U997 (N_997,N_940,N_933);
or U998 (N_998,N_916,N_936);
or U999 (N_999,N_946,N_917);
nand U1000 (N_1000,N_955,N_953);
nand U1001 (N_1001,N_980,N_979);
or U1002 (N_1002,N_951,N_990);
and U1003 (N_1003,N_988,N_996);
nand U1004 (N_1004,N_971,N_956);
nor U1005 (N_1005,N_958,N_991);
nor U1006 (N_1006,N_982,N_998);
and U1007 (N_1007,N_952,N_963);
nand U1008 (N_1008,N_954,N_999);
xnor U1009 (N_1009,N_964,N_992);
or U1010 (N_1010,N_961,N_966);
and U1011 (N_1011,N_959,N_977);
nand U1012 (N_1012,N_950,N_967);
nand U1013 (N_1013,N_972,N_995);
nor U1014 (N_1014,N_993,N_987);
and U1015 (N_1015,N_970,N_997);
and U1016 (N_1016,N_994,N_978);
nand U1017 (N_1017,N_957,N_968);
and U1018 (N_1018,N_976,N_969);
or U1019 (N_1019,N_974,N_965);
nor U1020 (N_1020,N_989,N_983);
nand U1021 (N_1021,N_960,N_962);
and U1022 (N_1022,N_986,N_975);
nor U1023 (N_1023,N_981,N_973);
nor U1024 (N_1024,N_984,N_985);
or U1025 (N_1025,N_979,N_989);
nor U1026 (N_1026,N_968,N_987);
or U1027 (N_1027,N_955,N_997);
nand U1028 (N_1028,N_951,N_992);
or U1029 (N_1029,N_980,N_988);
or U1030 (N_1030,N_989,N_965);
nor U1031 (N_1031,N_991,N_962);
or U1032 (N_1032,N_971,N_968);
nand U1033 (N_1033,N_950,N_980);
or U1034 (N_1034,N_952,N_950);
nor U1035 (N_1035,N_987,N_955);
nor U1036 (N_1036,N_976,N_993);
or U1037 (N_1037,N_982,N_967);
and U1038 (N_1038,N_950,N_987);
nor U1039 (N_1039,N_980,N_956);
and U1040 (N_1040,N_960,N_988);
nor U1041 (N_1041,N_984,N_975);
nand U1042 (N_1042,N_956,N_996);
nand U1043 (N_1043,N_998,N_973);
or U1044 (N_1044,N_974,N_952);
or U1045 (N_1045,N_975,N_974);
nand U1046 (N_1046,N_980,N_987);
nor U1047 (N_1047,N_957,N_996);
nor U1048 (N_1048,N_970,N_995);
nand U1049 (N_1049,N_991,N_998);
or U1050 (N_1050,N_1021,N_1028);
or U1051 (N_1051,N_1003,N_1015);
and U1052 (N_1052,N_1018,N_1013);
and U1053 (N_1053,N_1036,N_1041);
nand U1054 (N_1054,N_1016,N_1047);
nand U1055 (N_1055,N_1002,N_1019);
and U1056 (N_1056,N_1039,N_1045);
nor U1057 (N_1057,N_1008,N_1007);
or U1058 (N_1058,N_1011,N_1001);
nand U1059 (N_1059,N_1033,N_1046);
and U1060 (N_1060,N_1030,N_1026);
and U1061 (N_1061,N_1020,N_1049);
nor U1062 (N_1062,N_1014,N_1006);
nor U1063 (N_1063,N_1040,N_1037);
nor U1064 (N_1064,N_1042,N_1012);
xnor U1065 (N_1065,N_1043,N_1044);
nor U1066 (N_1066,N_1029,N_1031);
nand U1067 (N_1067,N_1017,N_1023);
and U1068 (N_1068,N_1048,N_1025);
nand U1069 (N_1069,N_1038,N_1034);
nor U1070 (N_1070,N_1027,N_1035);
and U1071 (N_1071,N_1024,N_1004);
nand U1072 (N_1072,N_1000,N_1032);
and U1073 (N_1073,N_1005,N_1009);
nand U1074 (N_1074,N_1022,N_1010);
and U1075 (N_1075,N_1031,N_1015);
nor U1076 (N_1076,N_1040,N_1047);
and U1077 (N_1077,N_1014,N_1041);
and U1078 (N_1078,N_1035,N_1018);
and U1079 (N_1079,N_1048,N_1011);
nand U1080 (N_1080,N_1029,N_1040);
nor U1081 (N_1081,N_1000,N_1005);
nor U1082 (N_1082,N_1042,N_1014);
nand U1083 (N_1083,N_1040,N_1048);
nor U1084 (N_1084,N_1047,N_1049);
nor U1085 (N_1085,N_1040,N_1018);
or U1086 (N_1086,N_1025,N_1017);
nor U1087 (N_1087,N_1038,N_1046);
nand U1088 (N_1088,N_1011,N_1009);
nor U1089 (N_1089,N_1042,N_1043);
nand U1090 (N_1090,N_1005,N_1030);
and U1091 (N_1091,N_1036,N_1034);
and U1092 (N_1092,N_1041,N_1016);
and U1093 (N_1093,N_1000,N_1022);
nor U1094 (N_1094,N_1033,N_1037);
and U1095 (N_1095,N_1023,N_1025);
and U1096 (N_1096,N_1010,N_1028);
or U1097 (N_1097,N_1038,N_1037);
nor U1098 (N_1098,N_1032,N_1008);
nor U1099 (N_1099,N_1005,N_1045);
nand U1100 (N_1100,N_1096,N_1099);
nand U1101 (N_1101,N_1081,N_1091);
xnor U1102 (N_1102,N_1087,N_1064);
nand U1103 (N_1103,N_1080,N_1085);
or U1104 (N_1104,N_1053,N_1054);
and U1105 (N_1105,N_1065,N_1084);
nand U1106 (N_1106,N_1052,N_1070);
xnor U1107 (N_1107,N_1078,N_1092);
nor U1108 (N_1108,N_1089,N_1094);
nand U1109 (N_1109,N_1067,N_1079);
and U1110 (N_1110,N_1075,N_1069);
or U1111 (N_1111,N_1088,N_1073);
or U1112 (N_1112,N_1076,N_1058);
and U1113 (N_1113,N_1055,N_1066);
or U1114 (N_1114,N_1095,N_1093);
nand U1115 (N_1115,N_1062,N_1060);
and U1116 (N_1116,N_1083,N_1074);
nor U1117 (N_1117,N_1086,N_1059);
nand U1118 (N_1118,N_1057,N_1090);
and U1119 (N_1119,N_1077,N_1051);
or U1120 (N_1120,N_1050,N_1063);
or U1121 (N_1121,N_1071,N_1098);
and U1122 (N_1122,N_1056,N_1082);
nand U1123 (N_1123,N_1061,N_1068);
nand U1124 (N_1124,N_1097,N_1072);
and U1125 (N_1125,N_1096,N_1057);
nor U1126 (N_1126,N_1090,N_1077);
or U1127 (N_1127,N_1056,N_1070);
and U1128 (N_1128,N_1081,N_1095);
and U1129 (N_1129,N_1091,N_1071);
nand U1130 (N_1130,N_1086,N_1061);
or U1131 (N_1131,N_1098,N_1099);
nand U1132 (N_1132,N_1065,N_1095);
or U1133 (N_1133,N_1079,N_1065);
nor U1134 (N_1134,N_1061,N_1062);
nor U1135 (N_1135,N_1051,N_1091);
and U1136 (N_1136,N_1079,N_1050);
or U1137 (N_1137,N_1081,N_1092);
and U1138 (N_1138,N_1069,N_1082);
or U1139 (N_1139,N_1099,N_1089);
nor U1140 (N_1140,N_1054,N_1095);
nand U1141 (N_1141,N_1053,N_1077);
and U1142 (N_1142,N_1078,N_1087);
nor U1143 (N_1143,N_1082,N_1067);
and U1144 (N_1144,N_1050,N_1073);
and U1145 (N_1145,N_1064,N_1051);
nand U1146 (N_1146,N_1066,N_1084);
and U1147 (N_1147,N_1077,N_1075);
and U1148 (N_1148,N_1078,N_1055);
nand U1149 (N_1149,N_1054,N_1073);
nand U1150 (N_1150,N_1143,N_1116);
or U1151 (N_1151,N_1147,N_1114);
nand U1152 (N_1152,N_1122,N_1136);
nand U1153 (N_1153,N_1111,N_1118);
nand U1154 (N_1154,N_1108,N_1126);
nor U1155 (N_1155,N_1115,N_1101);
and U1156 (N_1156,N_1113,N_1148);
and U1157 (N_1157,N_1100,N_1145);
nand U1158 (N_1158,N_1134,N_1129);
or U1159 (N_1159,N_1119,N_1142);
nor U1160 (N_1160,N_1149,N_1135);
nand U1161 (N_1161,N_1125,N_1112);
or U1162 (N_1162,N_1104,N_1120);
and U1163 (N_1163,N_1146,N_1105);
nand U1164 (N_1164,N_1132,N_1106);
nand U1165 (N_1165,N_1140,N_1139);
and U1166 (N_1166,N_1124,N_1127);
nand U1167 (N_1167,N_1109,N_1137);
nor U1168 (N_1168,N_1128,N_1141);
or U1169 (N_1169,N_1121,N_1138);
nand U1170 (N_1170,N_1130,N_1107);
or U1171 (N_1171,N_1102,N_1133);
nor U1172 (N_1172,N_1110,N_1117);
or U1173 (N_1173,N_1103,N_1131);
xnor U1174 (N_1174,N_1144,N_1123);
and U1175 (N_1175,N_1142,N_1129);
and U1176 (N_1176,N_1139,N_1143);
or U1177 (N_1177,N_1135,N_1136);
nand U1178 (N_1178,N_1103,N_1144);
or U1179 (N_1179,N_1114,N_1145);
nor U1180 (N_1180,N_1116,N_1114);
nand U1181 (N_1181,N_1116,N_1103);
nor U1182 (N_1182,N_1111,N_1142);
nand U1183 (N_1183,N_1135,N_1101);
or U1184 (N_1184,N_1142,N_1130);
nor U1185 (N_1185,N_1126,N_1129);
nor U1186 (N_1186,N_1143,N_1103);
or U1187 (N_1187,N_1136,N_1112);
nand U1188 (N_1188,N_1133,N_1132);
nor U1189 (N_1189,N_1133,N_1129);
and U1190 (N_1190,N_1138,N_1137);
and U1191 (N_1191,N_1118,N_1141);
or U1192 (N_1192,N_1126,N_1107);
or U1193 (N_1193,N_1131,N_1105);
nand U1194 (N_1194,N_1104,N_1149);
xnor U1195 (N_1195,N_1132,N_1136);
nor U1196 (N_1196,N_1120,N_1135);
and U1197 (N_1197,N_1109,N_1100);
nand U1198 (N_1198,N_1146,N_1118);
nand U1199 (N_1199,N_1136,N_1123);
nand U1200 (N_1200,N_1156,N_1180);
nand U1201 (N_1201,N_1195,N_1177);
nand U1202 (N_1202,N_1157,N_1179);
nand U1203 (N_1203,N_1191,N_1184);
nor U1204 (N_1204,N_1190,N_1199);
and U1205 (N_1205,N_1154,N_1152);
nor U1206 (N_1206,N_1168,N_1165);
or U1207 (N_1207,N_1166,N_1155);
or U1208 (N_1208,N_1153,N_1178);
nand U1209 (N_1209,N_1197,N_1198);
nand U1210 (N_1210,N_1183,N_1169);
or U1211 (N_1211,N_1187,N_1170);
nand U1212 (N_1212,N_1189,N_1193);
and U1213 (N_1213,N_1151,N_1164);
and U1214 (N_1214,N_1161,N_1162);
nor U1215 (N_1215,N_1176,N_1150);
or U1216 (N_1216,N_1185,N_1192);
and U1217 (N_1217,N_1196,N_1167);
nor U1218 (N_1218,N_1182,N_1175);
xnor U1219 (N_1219,N_1159,N_1194);
nor U1220 (N_1220,N_1158,N_1172);
nand U1221 (N_1221,N_1160,N_1173);
or U1222 (N_1222,N_1171,N_1174);
and U1223 (N_1223,N_1186,N_1163);
and U1224 (N_1224,N_1181,N_1188);
nor U1225 (N_1225,N_1165,N_1169);
nand U1226 (N_1226,N_1155,N_1192);
or U1227 (N_1227,N_1171,N_1172);
nor U1228 (N_1228,N_1178,N_1198);
and U1229 (N_1229,N_1166,N_1192);
nor U1230 (N_1230,N_1169,N_1155);
nor U1231 (N_1231,N_1198,N_1182);
nor U1232 (N_1232,N_1171,N_1164);
or U1233 (N_1233,N_1159,N_1175);
or U1234 (N_1234,N_1169,N_1177);
nor U1235 (N_1235,N_1194,N_1186);
nor U1236 (N_1236,N_1162,N_1178);
nand U1237 (N_1237,N_1171,N_1177);
nand U1238 (N_1238,N_1164,N_1192);
nor U1239 (N_1239,N_1156,N_1185);
nand U1240 (N_1240,N_1163,N_1173);
nand U1241 (N_1241,N_1187,N_1180);
and U1242 (N_1242,N_1183,N_1186);
nand U1243 (N_1243,N_1174,N_1164);
nor U1244 (N_1244,N_1151,N_1153);
nand U1245 (N_1245,N_1196,N_1160);
nor U1246 (N_1246,N_1153,N_1158);
or U1247 (N_1247,N_1162,N_1184);
nand U1248 (N_1248,N_1183,N_1162);
nor U1249 (N_1249,N_1166,N_1164);
nand U1250 (N_1250,N_1209,N_1205);
nor U1251 (N_1251,N_1211,N_1218);
or U1252 (N_1252,N_1239,N_1241);
or U1253 (N_1253,N_1201,N_1234);
and U1254 (N_1254,N_1206,N_1232);
and U1255 (N_1255,N_1217,N_1236);
and U1256 (N_1256,N_1212,N_1220);
nand U1257 (N_1257,N_1214,N_1227);
nor U1258 (N_1258,N_1229,N_1233);
or U1259 (N_1259,N_1210,N_1208);
and U1260 (N_1260,N_1225,N_1235);
and U1261 (N_1261,N_1203,N_1228);
and U1262 (N_1262,N_1240,N_1230);
nand U1263 (N_1263,N_1243,N_1248);
or U1264 (N_1264,N_1216,N_1246);
nand U1265 (N_1265,N_1249,N_1231);
nor U1266 (N_1266,N_1245,N_1244);
or U1267 (N_1267,N_1223,N_1226);
and U1268 (N_1268,N_1202,N_1207);
nand U1269 (N_1269,N_1200,N_1224);
and U1270 (N_1270,N_1213,N_1222);
nand U1271 (N_1271,N_1238,N_1204);
nand U1272 (N_1272,N_1219,N_1247);
nand U1273 (N_1273,N_1215,N_1237);
and U1274 (N_1274,N_1221,N_1242);
nor U1275 (N_1275,N_1218,N_1224);
nand U1276 (N_1276,N_1238,N_1230);
nand U1277 (N_1277,N_1236,N_1223);
nand U1278 (N_1278,N_1207,N_1209);
nor U1279 (N_1279,N_1243,N_1221);
nand U1280 (N_1280,N_1246,N_1209);
or U1281 (N_1281,N_1232,N_1243);
or U1282 (N_1282,N_1221,N_1225);
or U1283 (N_1283,N_1205,N_1239);
nand U1284 (N_1284,N_1248,N_1206);
nor U1285 (N_1285,N_1211,N_1220);
or U1286 (N_1286,N_1215,N_1228);
and U1287 (N_1287,N_1208,N_1242);
nor U1288 (N_1288,N_1233,N_1240);
nor U1289 (N_1289,N_1221,N_1244);
or U1290 (N_1290,N_1226,N_1248);
nor U1291 (N_1291,N_1245,N_1202);
or U1292 (N_1292,N_1207,N_1237);
or U1293 (N_1293,N_1248,N_1207);
and U1294 (N_1294,N_1237,N_1214);
nand U1295 (N_1295,N_1223,N_1235);
nand U1296 (N_1296,N_1234,N_1247);
or U1297 (N_1297,N_1241,N_1243);
nand U1298 (N_1298,N_1233,N_1249);
or U1299 (N_1299,N_1247,N_1224);
and U1300 (N_1300,N_1291,N_1253);
and U1301 (N_1301,N_1259,N_1265);
or U1302 (N_1302,N_1277,N_1284);
and U1303 (N_1303,N_1299,N_1255);
and U1304 (N_1304,N_1257,N_1258);
nor U1305 (N_1305,N_1278,N_1289);
nand U1306 (N_1306,N_1288,N_1287);
nand U1307 (N_1307,N_1285,N_1294);
or U1308 (N_1308,N_1262,N_1266);
nor U1309 (N_1309,N_1279,N_1270);
nor U1310 (N_1310,N_1256,N_1275);
nand U1311 (N_1311,N_1251,N_1298);
nand U1312 (N_1312,N_1264,N_1271);
nand U1313 (N_1313,N_1281,N_1273);
nor U1314 (N_1314,N_1272,N_1268);
nor U1315 (N_1315,N_1295,N_1267);
and U1316 (N_1316,N_1269,N_1297);
or U1317 (N_1317,N_1283,N_1250);
or U1318 (N_1318,N_1260,N_1274);
nand U1319 (N_1319,N_1261,N_1290);
nor U1320 (N_1320,N_1293,N_1280);
nand U1321 (N_1321,N_1282,N_1254);
nand U1322 (N_1322,N_1263,N_1296);
nand U1323 (N_1323,N_1286,N_1252);
or U1324 (N_1324,N_1292,N_1276);
or U1325 (N_1325,N_1265,N_1252);
nor U1326 (N_1326,N_1293,N_1256);
or U1327 (N_1327,N_1251,N_1282);
nand U1328 (N_1328,N_1295,N_1258);
xor U1329 (N_1329,N_1251,N_1289);
nor U1330 (N_1330,N_1296,N_1269);
nor U1331 (N_1331,N_1262,N_1276);
and U1332 (N_1332,N_1279,N_1288);
nor U1333 (N_1333,N_1266,N_1298);
and U1334 (N_1334,N_1252,N_1275);
nand U1335 (N_1335,N_1282,N_1267);
or U1336 (N_1336,N_1273,N_1277);
xnor U1337 (N_1337,N_1259,N_1287);
or U1338 (N_1338,N_1287,N_1281);
or U1339 (N_1339,N_1289,N_1254);
or U1340 (N_1340,N_1268,N_1285);
nand U1341 (N_1341,N_1296,N_1259);
nand U1342 (N_1342,N_1295,N_1259);
nand U1343 (N_1343,N_1297,N_1289);
nand U1344 (N_1344,N_1284,N_1280);
nor U1345 (N_1345,N_1290,N_1289);
or U1346 (N_1346,N_1288,N_1257);
or U1347 (N_1347,N_1287,N_1297);
or U1348 (N_1348,N_1260,N_1279);
or U1349 (N_1349,N_1266,N_1286);
nand U1350 (N_1350,N_1325,N_1328);
and U1351 (N_1351,N_1314,N_1341);
and U1352 (N_1352,N_1304,N_1313);
or U1353 (N_1353,N_1343,N_1323);
or U1354 (N_1354,N_1307,N_1301);
and U1355 (N_1355,N_1306,N_1327);
nor U1356 (N_1356,N_1331,N_1334);
or U1357 (N_1357,N_1319,N_1336);
and U1358 (N_1358,N_1348,N_1311);
xor U1359 (N_1359,N_1320,N_1302);
nor U1360 (N_1360,N_1322,N_1317);
nand U1361 (N_1361,N_1316,N_1329);
and U1362 (N_1362,N_1324,N_1309);
or U1363 (N_1363,N_1300,N_1305);
nand U1364 (N_1364,N_1308,N_1315);
nand U1365 (N_1365,N_1342,N_1346);
nor U1366 (N_1366,N_1318,N_1349);
nand U1367 (N_1367,N_1345,N_1321);
or U1368 (N_1368,N_1344,N_1303);
and U1369 (N_1369,N_1310,N_1337);
nor U1370 (N_1370,N_1335,N_1339);
and U1371 (N_1371,N_1326,N_1340);
nand U1372 (N_1372,N_1338,N_1330);
and U1373 (N_1373,N_1312,N_1333);
nand U1374 (N_1374,N_1347,N_1332);
nand U1375 (N_1375,N_1331,N_1314);
nand U1376 (N_1376,N_1312,N_1306);
and U1377 (N_1377,N_1337,N_1349);
and U1378 (N_1378,N_1327,N_1334);
and U1379 (N_1379,N_1328,N_1347);
or U1380 (N_1380,N_1336,N_1333);
nor U1381 (N_1381,N_1333,N_1343);
and U1382 (N_1382,N_1323,N_1342);
nor U1383 (N_1383,N_1310,N_1342);
nor U1384 (N_1384,N_1344,N_1302);
nor U1385 (N_1385,N_1333,N_1302);
nor U1386 (N_1386,N_1345,N_1302);
nand U1387 (N_1387,N_1314,N_1348);
nand U1388 (N_1388,N_1344,N_1333);
nor U1389 (N_1389,N_1341,N_1305);
or U1390 (N_1390,N_1302,N_1337);
or U1391 (N_1391,N_1324,N_1312);
or U1392 (N_1392,N_1311,N_1306);
or U1393 (N_1393,N_1307,N_1309);
or U1394 (N_1394,N_1320,N_1319);
or U1395 (N_1395,N_1331,N_1313);
nor U1396 (N_1396,N_1337,N_1331);
nand U1397 (N_1397,N_1304,N_1327);
and U1398 (N_1398,N_1310,N_1336);
nor U1399 (N_1399,N_1343,N_1315);
nor U1400 (N_1400,N_1370,N_1361);
nor U1401 (N_1401,N_1375,N_1355);
xnor U1402 (N_1402,N_1368,N_1394);
nor U1403 (N_1403,N_1393,N_1350);
and U1404 (N_1404,N_1383,N_1359);
and U1405 (N_1405,N_1386,N_1395);
nor U1406 (N_1406,N_1354,N_1373);
nor U1407 (N_1407,N_1358,N_1392);
nor U1408 (N_1408,N_1387,N_1382);
or U1409 (N_1409,N_1388,N_1363);
or U1410 (N_1410,N_1374,N_1353);
and U1411 (N_1411,N_1377,N_1384);
nor U1412 (N_1412,N_1365,N_1364);
or U1413 (N_1413,N_1369,N_1399);
xnor U1414 (N_1414,N_1376,N_1390);
nor U1415 (N_1415,N_1371,N_1351);
or U1416 (N_1416,N_1381,N_1397);
or U1417 (N_1417,N_1367,N_1379);
nor U1418 (N_1418,N_1360,N_1389);
or U1419 (N_1419,N_1391,N_1380);
nor U1420 (N_1420,N_1378,N_1385);
nor U1421 (N_1421,N_1352,N_1366);
and U1422 (N_1422,N_1356,N_1362);
or U1423 (N_1423,N_1398,N_1357);
nand U1424 (N_1424,N_1396,N_1372);
nor U1425 (N_1425,N_1376,N_1384);
nand U1426 (N_1426,N_1357,N_1355);
or U1427 (N_1427,N_1352,N_1390);
xor U1428 (N_1428,N_1388,N_1382);
and U1429 (N_1429,N_1351,N_1367);
nand U1430 (N_1430,N_1369,N_1370);
nand U1431 (N_1431,N_1360,N_1351);
or U1432 (N_1432,N_1384,N_1365);
and U1433 (N_1433,N_1370,N_1384);
nor U1434 (N_1434,N_1362,N_1377);
and U1435 (N_1435,N_1365,N_1371);
nor U1436 (N_1436,N_1374,N_1390);
or U1437 (N_1437,N_1350,N_1365);
nand U1438 (N_1438,N_1387,N_1353);
and U1439 (N_1439,N_1386,N_1376);
and U1440 (N_1440,N_1379,N_1369);
or U1441 (N_1441,N_1368,N_1382);
nor U1442 (N_1442,N_1362,N_1391);
and U1443 (N_1443,N_1358,N_1354);
nor U1444 (N_1444,N_1378,N_1367);
and U1445 (N_1445,N_1376,N_1399);
or U1446 (N_1446,N_1386,N_1351);
nand U1447 (N_1447,N_1352,N_1376);
nor U1448 (N_1448,N_1381,N_1375);
nor U1449 (N_1449,N_1358,N_1352);
and U1450 (N_1450,N_1419,N_1402);
nor U1451 (N_1451,N_1431,N_1415);
and U1452 (N_1452,N_1433,N_1432);
nand U1453 (N_1453,N_1413,N_1447);
or U1454 (N_1454,N_1425,N_1409);
and U1455 (N_1455,N_1446,N_1435);
or U1456 (N_1456,N_1441,N_1444);
nor U1457 (N_1457,N_1445,N_1434);
and U1458 (N_1458,N_1407,N_1418);
and U1459 (N_1459,N_1404,N_1417);
or U1460 (N_1460,N_1428,N_1439);
and U1461 (N_1461,N_1401,N_1411);
or U1462 (N_1462,N_1436,N_1424);
nand U1463 (N_1463,N_1422,N_1442);
nor U1464 (N_1464,N_1406,N_1438);
or U1465 (N_1465,N_1405,N_1423);
nor U1466 (N_1466,N_1408,N_1427);
nor U1467 (N_1467,N_1400,N_1443);
or U1468 (N_1468,N_1420,N_1437);
nor U1469 (N_1469,N_1426,N_1410);
nand U1470 (N_1470,N_1448,N_1430);
nand U1471 (N_1471,N_1449,N_1412);
or U1472 (N_1472,N_1429,N_1403);
or U1473 (N_1473,N_1416,N_1421);
and U1474 (N_1474,N_1440,N_1414);
nand U1475 (N_1475,N_1420,N_1400);
or U1476 (N_1476,N_1428,N_1431);
or U1477 (N_1477,N_1424,N_1440);
nor U1478 (N_1478,N_1412,N_1420);
or U1479 (N_1479,N_1416,N_1444);
nor U1480 (N_1480,N_1435,N_1433);
nor U1481 (N_1481,N_1415,N_1410);
nor U1482 (N_1482,N_1434,N_1422);
and U1483 (N_1483,N_1410,N_1418);
and U1484 (N_1484,N_1416,N_1449);
nand U1485 (N_1485,N_1429,N_1414);
and U1486 (N_1486,N_1440,N_1446);
and U1487 (N_1487,N_1400,N_1403);
and U1488 (N_1488,N_1445,N_1437);
or U1489 (N_1489,N_1411,N_1431);
or U1490 (N_1490,N_1423,N_1415);
or U1491 (N_1491,N_1406,N_1433);
and U1492 (N_1492,N_1413,N_1416);
and U1493 (N_1493,N_1420,N_1426);
nor U1494 (N_1494,N_1428,N_1418);
nand U1495 (N_1495,N_1429,N_1416);
or U1496 (N_1496,N_1411,N_1437);
or U1497 (N_1497,N_1408,N_1424);
and U1498 (N_1498,N_1422,N_1420);
nand U1499 (N_1499,N_1410,N_1434);
nand U1500 (N_1500,N_1496,N_1470);
nor U1501 (N_1501,N_1454,N_1466);
nor U1502 (N_1502,N_1468,N_1462);
or U1503 (N_1503,N_1488,N_1493);
or U1504 (N_1504,N_1472,N_1453);
or U1505 (N_1505,N_1499,N_1451);
nor U1506 (N_1506,N_1452,N_1461);
nand U1507 (N_1507,N_1475,N_1465);
or U1508 (N_1508,N_1497,N_1474);
nor U1509 (N_1509,N_1491,N_1477);
nor U1510 (N_1510,N_1467,N_1478);
and U1511 (N_1511,N_1458,N_1476);
nand U1512 (N_1512,N_1490,N_1489);
and U1513 (N_1513,N_1464,N_1455);
nor U1514 (N_1514,N_1494,N_1498);
nand U1515 (N_1515,N_1485,N_1484);
nand U1516 (N_1516,N_1473,N_1471);
and U1517 (N_1517,N_1487,N_1495);
nand U1518 (N_1518,N_1463,N_1480);
and U1519 (N_1519,N_1492,N_1457);
nor U1520 (N_1520,N_1450,N_1479);
nor U1521 (N_1521,N_1456,N_1469);
or U1522 (N_1522,N_1483,N_1486);
or U1523 (N_1523,N_1482,N_1459);
and U1524 (N_1524,N_1481,N_1460);
and U1525 (N_1525,N_1496,N_1483);
nand U1526 (N_1526,N_1483,N_1498);
nor U1527 (N_1527,N_1480,N_1482);
xor U1528 (N_1528,N_1484,N_1488);
nand U1529 (N_1529,N_1499,N_1474);
nand U1530 (N_1530,N_1465,N_1457);
nor U1531 (N_1531,N_1485,N_1466);
nand U1532 (N_1532,N_1459,N_1457);
nor U1533 (N_1533,N_1468,N_1450);
and U1534 (N_1534,N_1467,N_1484);
nand U1535 (N_1535,N_1496,N_1472);
or U1536 (N_1536,N_1486,N_1453);
and U1537 (N_1537,N_1465,N_1472);
or U1538 (N_1538,N_1479,N_1470);
and U1539 (N_1539,N_1486,N_1496);
and U1540 (N_1540,N_1482,N_1496);
nor U1541 (N_1541,N_1460,N_1464);
and U1542 (N_1542,N_1469,N_1492);
nor U1543 (N_1543,N_1476,N_1492);
nand U1544 (N_1544,N_1451,N_1477);
nor U1545 (N_1545,N_1489,N_1488);
and U1546 (N_1546,N_1451,N_1459);
or U1547 (N_1547,N_1491,N_1463);
and U1548 (N_1548,N_1486,N_1457);
nor U1549 (N_1549,N_1498,N_1477);
nand U1550 (N_1550,N_1540,N_1500);
nor U1551 (N_1551,N_1546,N_1521);
nand U1552 (N_1552,N_1538,N_1516);
and U1553 (N_1553,N_1515,N_1531);
xor U1554 (N_1554,N_1514,N_1522);
or U1555 (N_1555,N_1523,N_1512);
and U1556 (N_1556,N_1505,N_1506);
nand U1557 (N_1557,N_1511,N_1501);
and U1558 (N_1558,N_1507,N_1536);
nor U1559 (N_1559,N_1535,N_1542);
and U1560 (N_1560,N_1527,N_1541);
or U1561 (N_1561,N_1509,N_1502);
nor U1562 (N_1562,N_1528,N_1530);
nor U1563 (N_1563,N_1548,N_1526);
or U1564 (N_1564,N_1508,N_1525);
nor U1565 (N_1565,N_1510,N_1533);
nor U1566 (N_1566,N_1539,N_1503);
nand U1567 (N_1567,N_1534,N_1544);
nand U1568 (N_1568,N_1504,N_1543);
nor U1569 (N_1569,N_1537,N_1524);
nand U1570 (N_1570,N_1520,N_1549);
nand U1571 (N_1571,N_1518,N_1545);
and U1572 (N_1572,N_1529,N_1547);
and U1573 (N_1573,N_1513,N_1532);
and U1574 (N_1574,N_1517,N_1519);
nand U1575 (N_1575,N_1529,N_1531);
nor U1576 (N_1576,N_1514,N_1532);
and U1577 (N_1577,N_1527,N_1503);
nor U1578 (N_1578,N_1504,N_1535);
nor U1579 (N_1579,N_1524,N_1506);
or U1580 (N_1580,N_1526,N_1524);
or U1581 (N_1581,N_1516,N_1539);
nor U1582 (N_1582,N_1500,N_1541);
or U1583 (N_1583,N_1547,N_1540);
nand U1584 (N_1584,N_1524,N_1504);
or U1585 (N_1585,N_1542,N_1547);
and U1586 (N_1586,N_1537,N_1517);
or U1587 (N_1587,N_1540,N_1516);
or U1588 (N_1588,N_1537,N_1501);
nand U1589 (N_1589,N_1525,N_1515);
nor U1590 (N_1590,N_1541,N_1528);
or U1591 (N_1591,N_1523,N_1514);
or U1592 (N_1592,N_1507,N_1509);
or U1593 (N_1593,N_1516,N_1506);
nor U1594 (N_1594,N_1544,N_1526);
nor U1595 (N_1595,N_1528,N_1514);
and U1596 (N_1596,N_1544,N_1525);
nor U1597 (N_1597,N_1546,N_1503);
and U1598 (N_1598,N_1542,N_1543);
nor U1599 (N_1599,N_1545,N_1503);
nand U1600 (N_1600,N_1561,N_1586);
and U1601 (N_1601,N_1592,N_1575);
and U1602 (N_1602,N_1584,N_1591);
and U1603 (N_1603,N_1588,N_1576);
or U1604 (N_1604,N_1577,N_1559);
and U1605 (N_1605,N_1569,N_1556);
and U1606 (N_1606,N_1555,N_1552);
or U1607 (N_1607,N_1578,N_1595);
xor U1608 (N_1608,N_1554,N_1572);
or U1609 (N_1609,N_1581,N_1551);
and U1610 (N_1610,N_1599,N_1594);
nor U1611 (N_1611,N_1596,N_1579);
nand U1612 (N_1612,N_1582,N_1564);
and U1613 (N_1613,N_1585,N_1589);
or U1614 (N_1614,N_1558,N_1562);
or U1615 (N_1615,N_1571,N_1557);
nor U1616 (N_1616,N_1593,N_1550);
nand U1617 (N_1617,N_1567,N_1583);
nand U1618 (N_1618,N_1590,N_1565);
nand U1619 (N_1619,N_1566,N_1553);
nand U1620 (N_1620,N_1574,N_1587);
nor U1621 (N_1621,N_1568,N_1598);
nor U1622 (N_1622,N_1563,N_1573);
nor U1623 (N_1623,N_1560,N_1597);
and U1624 (N_1624,N_1580,N_1570);
nor U1625 (N_1625,N_1592,N_1552);
nor U1626 (N_1626,N_1551,N_1557);
and U1627 (N_1627,N_1568,N_1577);
and U1628 (N_1628,N_1565,N_1569);
nor U1629 (N_1629,N_1588,N_1557);
and U1630 (N_1630,N_1595,N_1557);
nand U1631 (N_1631,N_1589,N_1571);
and U1632 (N_1632,N_1558,N_1563);
nor U1633 (N_1633,N_1587,N_1551);
nor U1634 (N_1634,N_1592,N_1559);
nor U1635 (N_1635,N_1593,N_1552);
or U1636 (N_1636,N_1582,N_1580);
nor U1637 (N_1637,N_1564,N_1580);
nor U1638 (N_1638,N_1581,N_1555);
and U1639 (N_1639,N_1562,N_1556);
nor U1640 (N_1640,N_1575,N_1599);
nor U1641 (N_1641,N_1567,N_1575);
nand U1642 (N_1642,N_1559,N_1596);
nor U1643 (N_1643,N_1575,N_1576);
nor U1644 (N_1644,N_1591,N_1564);
nand U1645 (N_1645,N_1574,N_1577);
and U1646 (N_1646,N_1576,N_1577);
nor U1647 (N_1647,N_1596,N_1599);
and U1648 (N_1648,N_1565,N_1572);
or U1649 (N_1649,N_1588,N_1562);
or U1650 (N_1650,N_1646,N_1618);
nand U1651 (N_1651,N_1615,N_1617);
nand U1652 (N_1652,N_1609,N_1604);
or U1653 (N_1653,N_1629,N_1602);
nand U1654 (N_1654,N_1613,N_1640);
nand U1655 (N_1655,N_1633,N_1643);
or U1656 (N_1656,N_1606,N_1611);
nor U1657 (N_1657,N_1645,N_1614);
nor U1658 (N_1658,N_1647,N_1619);
or U1659 (N_1659,N_1636,N_1601);
nand U1660 (N_1660,N_1649,N_1621);
and U1661 (N_1661,N_1634,N_1637);
and U1662 (N_1662,N_1635,N_1641);
nand U1663 (N_1663,N_1605,N_1608);
and U1664 (N_1664,N_1642,N_1638);
and U1665 (N_1665,N_1628,N_1620);
or U1666 (N_1666,N_1612,N_1622);
nor U1667 (N_1667,N_1627,N_1648);
and U1668 (N_1668,N_1625,N_1623);
and U1669 (N_1669,N_1603,N_1631);
or U1670 (N_1670,N_1624,N_1610);
and U1671 (N_1671,N_1616,N_1630);
nand U1672 (N_1672,N_1644,N_1632);
and U1673 (N_1673,N_1626,N_1639);
nor U1674 (N_1674,N_1600,N_1607);
and U1675 (N_1675,N_1602,N_1617);
nor U1676 (N_1676,N_1609,N_1600);
nand U1677 (N_1677,N_1630,N_1636);
nand U1678 (N_1678,N_1627,N_1613);
or U1679 (N_1679,N_1612,N_1641);
or U1680 (N_1680,N_1612,N_1600);
or U1681 (N_1681,N_1614,N_1609);
and U1682 (N_1682,N_1622,N_1642);
nand U1683 (N_1683,N_1624,N_1625);
or U1684 (N_1684,N_1613,N_1633);
nor U1685 (N_1685,N_1629,N_1634);
nand U1686 (N_1686,N_1603,N_1615);
or U1687 (N_1687,N_1601,N_1643);
or U1688 (N_1688,N_1615,N_1632);
and U1689 (N_1689,N_1633,N_1647);
and U1690 (N_1690,N_1624,N_1601);
and U1691 (N_1691,N_1606,N_1625);
and U1692 (N_1692,N_1601,N_1646);
and U1693 (N_1693,N_1636,N_1625);
or U1694 (N_1694,N_1620,N_1633);
or U1695 (N_1695,N_1612,N_1603);
and U1696 (N_1696,N_1648,N_1649);
nand U1697 (N_1697,N_1632,N_1639);
or U1698 (N_1698,N_1645,N_1627);
or U1699 (N_1699,N_1634,N_1645);
and U1700 (N_1700,N_1662,N_1689);
nand U1701 (N_1701,N_1660,N_1668);
nand U1702 (N_1702,N_1659,N_1658);
nand U1703 (N_1703,N_1674,N_1691);
and U1704 (N_1704,N_1687,N_1690);
nor U1705 (N_1705,N_1698,N_1676);
or U1706 (N_1706,N_1697,N_1664);
nand U1707 (N_1707,N_1686,N_1652);
nor U1708 (N_1708,N_1669,N_1667);
xor U1709 (N_1709,N_1693,N_1656);
or U1710 (N_1710,N_1680,N_1694);
or U1711 (N_1711,N_1681,N_1657);
and U1712 (N_1712,N_1695,N_1688);
nand U1713 (N_1713,N_1671,N_1692);
nand U1714 (N_1714,N_1673,N_1666);
nor U1715 (N_1715,N_1684,N_1696);
nand U1716 (N_1716,N_1670,N_1655);
and U1717 (N_1717,N_1654,N_1699);
or U1718 (N_1718,N_1672,N_1661);
nor U1719 (N_1719,N_1683,N_1653);
nor U1720 (N_1720,N_1677,N_1663);
nor U1721 (N_1721,N_1678,N_1650);
nor U1722 (N_1722,N_1685,N_1665);
or U1723 (N_1723,N_1682,N_1675);
and U1724 (N_1724,N_1651,N_1679);
and U1725 (N_1725,N_1654,N_1688);
nor U1726 (N_1726,N_1655,N_1694);
and U1727 (N_1727,N_1678,N_1664);
nor U1728 (N_1728,N_1655,N_1683);
nor U1729 (N_1729,N_1684,N_1669);
and U1730 (N_1730,N_1691,N_1669);
nand U1731 (N_1731,N_1678,N_1686);
nor U1732 (N_1732,N_1657,N_1668);
nand U1733 (N_1733,N_1660,N_1691);
or U1734 (N_1734,N_1657,N_1661);
or U1735 (N_1735,N_1663,N_1689);
nand U1736 (N_1736,N_1670,N_1678);
or U1737 (N_1737,N_1685,N_1695);
nor U1738 (N_1738,N_1650,N_1690);
nor U1739 (N_1739,N_1658,N_1672);
and U1740 (N_1740,N_1650,N_1694);
or U1741 (N_1741,N_1660,N_1655);
and U1742 (N_1742,N_1675,N_1689);
nor U1743 (N_1743,N_1687,N_1657);
and U1744 (N_1744,N_1683,N_1662);
or U1745 (N_1745,N_1668,N_1652);
or U1746 (N_1746,N_1656,N_1663);
and U1747 (N_1747,N_1654,N_1675);
nand U1748 (N_1748,N_1653,N_1680);
or U1749 (N_1749,N_1695,N_1697);
nor U1750 (N_1750,N_1741,N_1723);
nor U1751 (N_1751,N_1711,N_1701);
nand U1752 (N_1752,N_1714,N_1736);
or U1753 (N_1753,N_1720,N_1702);
and U1754 (N_1754,N_1735,N_1724);
nor U1755 (N_1755,N_1749,N_1705);
xnor U1756 (N_1756,N_1729,N_1706);
nor U1757 (N_1757,N_1746,N_1708);
nand U1758 (N_1758,N_1732,N_1745);
nor U1759 (N_1759,N_1731,N_1709);
and U1760 (N_1760,N_1722,N_1747);
nand U1761 (N_1761,N_1734,N_1715);
and U1762 (N_1762,N_1744,N_1728);
or U1763 (N_1763,N_1742,N_1725);
and U1764 (N_1764,N_1710,N_1703);
nor U1765 (N_1765,N_1721,N_1739);
nor U1766 (N_1766,N_1726,N_1730);
or U1767 (N_1767,N_1700,N_1707);
nor U1768 (N_1768,N_1719,N_1748);
nand U1769 (N_1769,N_1743,N_1713);
nand U1770 (N_1770,N_1733,N_1738);
nand U1771 (N_1771,N_1718,N_1737);
or U1772 (N_1772,N_1712,N_1740);
nor U1773 (N_1773,N_1727,N_1717);
nand U1774 (N_1774,N_1716,N_1704);
nand U1775 (N_1775,N_1713,N_1721);
nor U1776 (N_1776,N_1702,N_1704);
nand U1777 (N_1777,N_1719,N_1730);
nor U1778 (N_1778,N_1743,N_1721);
nor U1779 (N_1779,N_1742,N_1739);
nor U1780 (N_1780,N_1713,N_1709);
and U1781 (N_1781,N_1743,N_1712);
and U1782 (N_1782,N_1704,N_1701);
or U1783 (N_1783,N_1740,N_1728);
or U1784 (N_1784,N_1717,N_1720);
nand U1785 (N_1785,N_1727,N_1719);
and U1786 (N_1786,N_1705,N_1742);
nand U1787 (N_1787,N_1745,N_1739);
or U1788 (N_1788,N_1734,N_1738);
and U1789 (N_1789,N_1710,N_1729);
nand U1790 (N_1790,N_1701,N_1734);
or U1791 (N_1791,N_1720,N_1736);
nor U1792 (N_1792,N_1704,N_1710);
or U1793 (N_1793,N_1720,N_1745);
nor U1794 (N_1794,N_1742,N_1744);
and U1795 (N_1795,N_1742,N_1734);
and U1796 (N_1796,N_1718,N_1711);
nand U1797 (N_1797,N_1707,N_1740);
nor U1798 (N_1798,N_1731,N_1724);
nor U1799 (N_1799,N_1746,N_1720);
or U1800 (N_1800,N_1796,N_1785);
nor U1801 (N_1801,N_1755,N_1764);
nand U1802 (N_1802,N_1793,N_1790);
and U1803 (N_1803,N_1762,N_1768);
and U1804 (N_1804,N_1799,N_1792);
or U1805 (N_1805,N_1772,N_1794);
and U1806 (N_1806,N_1767,N_1795);
or U1807 (N_1807,N_1775,N_1781);
nand U1808 (N_1808,N_1766,N_1752);
nor U1809 (N_1809,N_1787,N_1776);
or U1810 (N_1810,N_1779,N_1782);
or U1811 (N_1811,N_1773,N_1786);
and U1812 (N_1812,N_1754,N_1798);
or U1813 (N_1813,N_1751,N_1789);
nor U1814 (N_1814,N_1777,N_1770);
or U1815 (N_1815,N_1763,N_1784);
and U1816 (N_1816,N_1778,N_1780);
nand U1817 (N_1817,N_1760,N_1774);
or U1818 (N_1818,N_1750,N_1788);
nand U1819 (N_1819,N_1783,N_1759);
nor U1820 (N_1820,N_1756,N_1771);
nand U1821 (N_1821,N_1761,N_1765);
nor U1822 (N_1822,N_1753,N_1757);
or U1823 (N_1823,N_1758,N_1797);
and U1824 (N_1824,N_1769,N_1791);
nand U1825 (N_1825,N_1784,N_1757);
and U1826 (N_1826,N_1766,N_1781);
nand U1827 (N_1827,N_1786,N_1790);
or U1828 (N_1828,N_1769,N_1796);
and U1829 (N_1829,N_1781,N_1776);
nand U1830 (N_1830,N_1771,N_1784);
nand U1831 (N_1831,N_1771,N_1799);
and U1832 (N_1832,N_1757,N_1799);
nand U1833 (N_1833,N_1794,N_1773);
nor U1834 (N_1834,N_1764,N_1777);
or U1835 (N_1835,N_1754,N_1761);
nand U1836 (N_1836,N_1755,N_1789);
or U1837 (N_1837,N_1770,N_1797);
nor U1838 (N_1838,N_1752,N_1765);
or U1839 (N_1839,N_1785,N_1795);
or U1840 (N_1840,N_1760,N_1763);
nand U1841 (N_1841,N_1757,N_1781);
nand U1842 (N_1842,N_1772,N_1759);
and U1843 (N_1843,N_1792,N_1776);
or U1844 (N_1844,N_1785,N_1752);
and U1845 (N_1845,N_1768,N_1793);
nand U1846 (N_1846,N_1787,N_1768);
nand U1847 (N_1847,N_1761,N_1770);
and U1848 (N_1848,N_1774,N_1783);
nand U1849 (N_1849,N_1771,N_1755);
nor U1850 (N_1850,N_1847,N_1829);
and U1851 (N_1851,N_1832,N_1809);
or U1852 (N_1852,N_1822,N_1820);
or U1853 (N_1853,N_1827,N_1810);
or U1854 (N_1854,N_1817,N_1800);
nor U1855 (N_1855,N_1803,N_1831);
and U1856 (N_1856,N_1841,N_1845);
or U1857 (N_1857,N_1848,N_1844);
and U1858 (N_1858,N_1821,N_1812);
nor U1859 (N_1859,N_1843,N_1839);
nor U1860 (N_1860,N_1811,N_1816);
or U1861 (N_1861,N_1813,N_1823);
nor U1862 (N_1862,N_1801,N_1828);
and U1863 (N_1863,N_1840,N_1825);
nor U1864 (N_1864,N_1802,N_1838);
and U1865 (N_1865,N_1815,N_1833);
nand U1866 (N_1866,N_1849,N_1846);
nand U1867 (N_1867,N_1835,N_1804);
nand U1868 (N_1868,N_1808,N_1814);
nand U1869 (N_1869,N_1837,N_1836);
nor U1870 (N_1870,N_1824,N_1805);
and U1871 (N_1871,N_1830,N_1826);
nor U1872 (N_1872,N_1806,N_1807);
and U1873 (N_1873,N_1819,N_1818);
and U1874 (N_1874,N_1842,N_1834);
nand U1875 (N_1875,N_1835,N_1828);
or U1876 (N_1876,N_1819,N_1803);
and U1877 (N_1877,N_1825,N_1806);
nand U1878 (N_1878,N_1824,N_1809);
nand U1879 (N_1879,N_1818,N_1836);
or U1880 (N_1880,N_1841,N_1800);
or U1881 (N_1881,N_1831,N_1842);
and U1882 (N_1882,N_1819,N_1826);
and U1883 (N_1883,N_1816,N_1847);
or U1884 (N_1884,N_1811,N_1820);
and U1885 (N_1885,N_1800,N_1809);
nor U1886 (N_1886,N_1849,N_1800);
or U1887 (N_1887,N_1821,N_1824);
nor U1888 (N_1888,N_1827,N_1820);
or U1889 (N_1889,N_1836,N_1839);
or U1890 (N_1890,N_1805,N_1810);
and U1891 (N_1891,N_1846,N_1848);
or U1892 (N_1892,N_1811,N_1801);
nor U1893 (N_1893,N_1823,N_1843);
or U1894 (N_1894,N_1829,N_1834);
nand U1895 (N_1895,N_1836,N_1827);
or U1896 (N_1896,N_1824,N_1844);
nand U1897 (N_1897,N_1818,N_1808);
nor U1898 (N_1898,N_1834,N_1825);
or U1899 (N_1899,N_1812,N_1832);
or U1900 (N_1900,N_1871,N_1862);
nand U1901 (N_1901,N_1869,N_1855);
nand U1902 (N_1902,N_1877,N_1878);
or U1903 (N_1903,N_1865,N_1879);
or U1904 (N_1904,N_1866,N_1858);
and U1905 (N_1905,N_1874,N_1895);
and U1906 (N_1906,N_1897,N_1875);
and U1907 (N_1907,N_1853,N_1850);
and U1908 (N_1908,N_1857,N_1896);
and U1909 (N_1909,N_1888,N_1894);
nand U1910 (N_1910,N_1868,N_1887);
and U1911 (N_1911,N_1885,N_1883);
nand U1912 (N_1912,N_1893,N_1860);
xor U1913 (N_1913,N_1891,N_1870);
or U1914 (N_1914,N_1859,N_1890);
nand U1915 (N_1915,N_1881,N_1864);
or U1916 (N_1916,N_1861,N_1876);
nand U1917 (N_1917,N_1886,N_1852);
and U1918 (N_1918,N_1867,N_1898);
nand U1919 (N_1919,N_1889,N_1899);
and U1920 (N_1920,N_1856,N_1851);
nor U1921 (N_1921,N_1863,N_1880);
or U1922 (N_1922,N_1873,N_1882);
nor U1923 (N_1923,N_1872,N_1854);
and U1924 (N_1924,N_1884,N_1892);
and U1925 (N_1925,N_1891,N_1856);
and U1926 (N_1926,N_1857,N_1897);
nand U1927 (N_1927,N_1863,N_1869);
or U1928 (N_1928,N_1883,N_1869);
nand U1929 (N_1929,N_1855,N_1892);
nand U1930 (N_1930,N_1892,N_1886);
or U1931 (N_1931,N_1877,N_1886);
and U1932 (N_1932,N_1892,N_1873);
or U1933 (N_1933,N_1867,N_1859);
and U1934 (N_1934,N_1853,N_1887);
and U1935 (N_1935,N_1874,N_1885);
nor U1936 (N_1936,N_1884,N_1876);
nand U1937 (N_1937,N_1854,N_1884);
nand U1938 (N_1938,N_1895,N_1862);
or U1939 (N_1939,N_1887,N_1884);
nor U1940 (N_1940,N_1856,N_1878);
nand U1941 (N_1941,N_1881,N_1863);
or U1942 (N_1942,N_1871,N_1856);
or U1943 (N_1943,N_1877,N_1884);
nor U1944 (N_1944,N_1893,N_1880);
nor U1945 (N_1945,N_1879,N_1876);
nand U1946 (N_1946,N_1898,N_1850);
nor U1947 (N_1947,N_1854,N_1858);
nand U1948 (N_1948,N_1888,N_1853);
nor U1949 (N_1949,N_1884,N_1861);
nor U1950 (N_1950,N_1936,N_1914);
or U1951 (N_1951,N_1938,N_1912);
and U1952 (N_1952,N_1949,N_1920);
nor U1953 (N_1953,N_1925,N_1931);
or U1954 (N_1954,N_1928,N_1948);
nor U1955 (N_1955,N_1941,N_1918);
and U1956 (N_1956,N_1911,N_1903);
and U1957 (N_1957,N_1900,N_1915);
or U1958 (N_1958,N_1930,N_1919);
nand U1959 (N_1959,N_1932,N_1909);
and U1960 (N_1960,N_1945,N_1924);
or U1961 (N_1961,N_1933,N_1944);
nor U1962 (N_1962,N_1917,N_1929);
and U1963 (N_1963,N_1916,N_1901);
or U1964 (N_1964,N_1904,N_1926);
nor U1965 (N_1965,N_1943,N_1910);
or U1966 (N_1966,N_1922,N_1947);
and U1967 (N_1967,N_1934,N_1940);
and U1968 (N_1968,N_1927,N_1937);
nor U1969 (N_1969,N_1902,N_1942);
and U1970 (N_1970,N_1913,N_1923);
and U1971 (N_1971,N_1939,N_1946);
or U1972 (N_1972,N_1905,N_1908);
nand U1973 (N_1973,N_1921,N_1906);
nor U1974 (N_1974,N_1935,N_1907);
nor U1975 (N_1975,N_1916,N_1938);
or U1976 (N_1976,N_1932,N_1936);
nand U1977 (N_1977,N_1916,N_1931);
and U1978 (N_1978,N_1901,N_1907);
nand U1979 (N_1979,N_1948,N_1941);
nand U1980 (N_1980,N_1913,N_1929);
nor U1981 (N_1981,N_1947,N_1933);
nor U1982 (N_1982,N_1941,N_1902);
or U1983 (N_1983,N_1937,N_1906);
or U1984 (N_1984,N_1936,N_1901);
nor U1985 (N_1985,N_1927,N_1947);
and U1986 (N_1986,N_1900,N_1949);
or U1987 (N_1987,N_1927,N_1903);
and U1988 (N_1988,N_1905,N_1936);
nand U1989 (N_1989,N_1901,N_1948);
or U1990 (N_1990,N_1934,N_1946);
nor U1991 (N_1991,N_1919,N_1933);
or U1992 (N_1992,N_1926,N_1916);
nand U1993 (N_1993,N_1914,N_1928);
or U1994 (N_1994,N_1921,N_1943);
nand U1995 (N_1995,N_1917,N_1915);
or U1996 (N_1996,N_1910,N_1917);
nand U1997 (N_1997,N_1904,N_1901);
nor U1998 (N_1998,N_1930,N_1936);
or U1999 (N_1999,N_1941,N_1922);
nand U2000 (N_2000,N_1991,N_1974);
and U2001 (N_2001,N_1997,N_1964);
nor U2002 (N_2002,N_1973,N_1957);
or U2003 (N_2003,N_1953,N_1963);
or U2004 (N_2004,N_1977,N_1969);
and U2005 (N_2005,N_1992,N_1960);
and U2006 (N_2006,N_1987,N_1959);
and U2007 (N_2007,N_1968,N_1980);
nand U2008 (N_2008,N_1999,N_1983);
nor U2009 (N_2009,N_1961,N_1971);
nor U2010 (N_2010,N_1998,N_1958);
or U2011 (N_2011,N_1950,N_1989);
nand U2012 (N_2012,N_1984,N_1995);
or U2013 (N_2013,N_1996,N_1979);
or U2014 (N_2014,N_1972,N_1981);
nand U2015 (N_2015,N_1985,N_1976);
or U2016 (N_2016,N_1988,N_1982);
nand U2017 (N_2017,N_1955,N_1978);
or U2018 (N_2018,N_1954,N_1994);
nor U2019 (N_2019,N_1967,N_1962);
and U2020 (N_2020,N_1966,N_1952);
nand U2021 (N_2021,N_1990,N_1986);
nand U2022 (N_2022,N_1951,N_1975);
nor U2023 (N_2023,N_1965,N_1993);
nor U2024 (N_2024,N_1970,N_1956);
nor U2025 (N_2025,N_1969,N_1967);
and U2026 (N_2026,N_1982,N_1963);
xnor U2027 (N_2027,N_1977,N_1958);
nor U2028 (N_2028,N_1978,N_1992);
nor U2029 (N_2029,N_1975,N_1978);
or U2030 (N_2030,N_1974,N_1977);
and U2031 (N_2031,N_1973,N_1959);
nor U2032 (N_2032,N_1956,N_1986);
and U2033 (N_2033,N_1977,N_1972);
and U2034 (N_2034,N_1972,N_1961);
nor U2035 (N_2035,N_1968,N_1972);
xnor U2036 (N_2036,N_1981,N_1996);
and U2037 (N_2037,N_1996,N_1986);
nor U2038 (N_2038,N_1972,N_1955);
or U2039 (N_2039,N_1982,N_1999);
and U2040 (N_2040,N_1972,N_1986);
nor U2041 (N_2041,N_1972,N_1954);
or U2042 (N_2042,N_1987,N_1998);
and U2043 (N_2043,N_1988,N_1995);
and U2044 (N_2044,N_1989,N_1986);
or U2045 (N_2045,N_1966,N_1967);
and U2046 (N_2046,N_1986,N_1993);
nand U2047 (N_2047,N_1993,N_1967);
nor U2048 (N_2048,N_1971,N_1978);
or U2049 (N_2049,N_1999,N_1952);
or U2050 (N_2050,N_2035,N_2022);
and U2051 (N_2051,N_2037,N_2023);
and U2052 (N_2052,N_2039,N_2009);
nor U2053 (N_2053,N_2015,N_2049);
or U2054 (N_2054,N_2041,N_2027);
nand U2055 (N_2055,N_2024,N_2020);
and U2056 (N_2056,N_2014,N_2042);
nor U2057 (N_2057,N_2002,N_2006);
or U2058 (N_2058,N_2026,N_2032);
nand U2059 (N_2059,N_2028,N_2047);
and U2060 (N_2060,N_2016,N_2013);
and U2061 (N_2061,N_2040,N_2003);
and U2062 (N_2062,N_2044,N_2025);
nand U2063 (N_2063,N_2005,N_2019);
and U2064 (N_2064,N_2031,N_2017);
or U2065 (N_2065,N_2034,N_2048);
and U2066 (N_2066,N_2018,N_2046);
and U2067 (N_2067,N_2029,N_2033);
and U2068 (N_2068,N_2010,N_2008);
nand U2069 (N_2069,N_2000,N_2038);
nand U2070 (N_2070,N_2043,N_2030);
or U2071 (N_2071,N_2012,N_2045);
nor U2072 (N_2072,N_2001,N_2007);
nand U2073 (N_2073,N_2036,N_2004);
nor U2074 (N_2074,N_2021,N_2011);
and U2075 (N_2075,N_2032,N_2012);
or U2076 (N_2076,N_2031,N_2025);
or U2077 (N_2077,N_2041,N_2006);
or U2078 (N_2078,N_2026,N_2033);
or U2079 (N_2079,N_2044,N_2011);
or U2080 (N_2080,N_2002,N_2047);
nand U2081 (N_2081,N_2014,N_2026);
and U2082 (N_2082,N_2037,N_2012);
nand U2083 (N_2083,N_2029,N_2039);
or U2084 (N_2084,N_2013,N_2004);
nor U2085 (N_2085,N_2035,N_2037);
nor U2086 (N_2086,N_2021,N_2042);
nand U2087 (N_2087,N_2030,N_2013);
and U2088 (N_2088,N_2008,N_2034);
nand U2089 (N_2089,N_2037,N_2030);
nand U2090 (N_2090,N_2032,N_2037);
nor U2091 (N_2091,N_2045,N_2032);
or U2092 (N_2092,N_2001,N_2018);
nand U2093 (N_2093,N_2020,N_2000);
nor U2094 (N_2094,N_2000,N_2019);
nor U2095 (N_2095,N_2048,N_2039);
or U2096 (N_2096,N_2023,N_2004);
and U2097 (N_2097,N_2030,N_2048);
nand U2098 (N_2098,N_2003,N_2047);
nand U2099 (N_2099,N_2039,N_2013);
and U2100 (N_2100,N_2092,N_2091);
or U2101 (N_2101,N_2070,N_2079);
nand U2102 (N_2102,N_2090,N_2069);
nand U2103 (N_2103,N_2054,N_2061);
nor U2104 (N_2104,N_2080,N_2073);
xor U2105 (N_2105,N_2066,N_2062);
nand U2106 (N_2106,N_2085,N_2088);
nor U2107 (N_2107,N_2059,N_2081);
and U2108 (N_2108,N_2057,N_2077);
and U2109 (N_2109,N_2056,N_2074);
nor U2110 (N_2110,N_2095,N_2055);
nor U2111 (N_2111,N_2087,N_2097);
or U2112 (N_2112,N_2093,N_2051);
and U2113 (N_2113,N_2064,N_2065);
nor U2114 (N_2114,N_2071,N_2098);
nand U2115 (N_2115,N_2084,N_2075);
or U2116 (N_2116,N_2089,N_2058);
and U2117 (N_2117,N_2082,N_2072);
and U2118 (N_2118,N_2094,N_2068);
and U2119 (N_2119,N_2052,N_2060);
nand U2120 (N_2120,N_2096,N_2078);
or U2121 (N_2121,N_2067,N_2063);
or U2122 (N_2122,N_2053,N_2050);
or U2123 (N_2123,N_2086,N_2083);
and U2124 (N_2124,N_2076,N_2099);
nor U2125 (N_2125,N_2081,N_2057);
or U2126 (N_2126,N_2096,N_2051);
or U2127 (N_2127,N_2084,N_2080);
xor U2128 (N_2128,N_2074,N_2077);
nand U2129 (N_2129,N_2092,N_2050);
nand U2130 (N_2130,N_2069,N_2050);
or U2131 (N_2131,N_2099,N_2093);
xor U2132 (N_2132,N_2076,N_2070);
nand U2133 (N_2133,N_2077,N_2079);
and U2134 (N_2134,N_2061,N_2073);
nor U2135 (N_2135,N_2092,N_2079);
or U2136 (N_2136,N_2075,N_2092);
nor U2137 (N_2137,N_2082,N_2057);
or U2138 (N_2138,N_2085,N_2053);
nor U2139 (N_2139,N_2065,N_2052);
or U2140 (N_2140,N_2063,N_2050);
nor U2141 (N_2141,N_2080,N_2088);
nand U2142 (N_2142,N_2087,N_2098);
nand U2143 (N_2143,N_2058,N_2091);
or U2144 (N_2144,N_2052,N_2090);
nor U2145 (N_2145,N_2088,N_2084);
and U2146 (N_2146,N_2071,N_2089);
and U2147 (N_2147,N_2082,N_2081);
and U2148 (N_2148,N_2084,N_2058);
nor U2149 (N_2149,N_2074,N_2050);
nor U2150 (N_2150,N_2104,N_2111);
and U2151 (N_2151,N_2110,N_2132);
nor U2152 (N_2152,N_2144,N_2102);
nand U2153 (N_2153,N_2108,N_2101);
or U2154 (N_2154,N_2113,N_2121);
nor U2155 (N_2155,N_2105,N_2129);
nand U2156 (N_2156,N_2147,N_2120);
and U2157 (N_2157,N_2134,N_2139);
or U2158 (N_2158,N_2103,N_2124);
and U2159 (N_2159,N_2112,N_2148);
and U2160 (N_2160,N_2116,N_2142);
and U2161 (N_2161,N_2109,N_2135);
nor U2162 (N_2162,N_2133,N_2100);
or U2163 (N_2163,N_2141,N_2118);
nor U2164 (N_2164,N_2123,N_2131);
nor U2165 (N_2165,N_2122,N_2128);
nand U2166 (N_2166,N_2149,N_2107);
nor U2167 (N_2167,N_2126,N_2145);
and U2168 (N_2168,N_2140,N_2106);
or U2169 (N_2169,N_2125,N_2127);
or U2170 (N_2170,N_2137,N_2146);
nand U2171 (N_2171,N_2115,N_2136);
or U2172 (N_2172,N_2117,N_2138);
nand U2173 (N_2173,N_2119,N_2143);
or U2174 (N_2174,N_2114,N_2130);
and U2175 (N_2175,N_2115,N_2137);
or U2176 (N_2176,N_2123,N_2111);
nor U2177 (N_2177,N_2112,N_2137);
nor U2178 (N_2178,N_2139,N_2140);
and U2179 (N_2179,N_2134,N_2111);
nand U2180 (N_2180,N_2116,N_2147);
nand U2181 (N_2181,N_2132,N_2125);
nand U2182 (N_2182,N_2103,N_2119);
or U2183 (N_2183,N_2118,N_2147);
nand U2184 (N_2184,N_2141,N_2148);
and U2185 (N_2185,N_2123,N_2119);
nand U2186 (N_2186,N_2146,N_2130);
nor U2187 (N_2187,N_2129,N_2125);
nor U2188 (N_2188,N_2124,N_2125);
nand U2189 (N_2189,N_2129,N_2147);
nor U2190 (N_2190,N_2108,N_2132);
nor U2191 (N_2191,N_2126,N_2128);
nor U2192 (N_2192,N_2141,N_2143);
nor U2193 (N_2193,N_2121,N_2148);
and U2194 (N_2194,N_2117,N_2105);
nor U2195 (N_2195,N_2148,N_2136);
nand U2196 (N_2196,N_2140,N_2137);
and U2197 (N_2197,N_2135,N_2136);
nand U2198 (N_2198,N_2138,N_2113);
or U2199 (N_2199,N_2140,N_2126);
nand U2200 (N_2200,N_2185,N_2154);
and U2201 (N_2201,N_2167,N_2189);
and U2202 (N_2202,N_2188,N_2182);
or U2203 (N_2203,N_2159,N_2170);
or U2204 (N_2204,N_2151,N_2193);
and U2205 (N_2205,N_2180,N_2169);
nor U2206 (N_2206,N_2161,N_2164);
nor U2207 (N_2207,N_2166,N_2195);
and U2208 (N_2208,N_2168,N_2150);
or U2209 (N_2209,N_2152,N_2165);
or U2210 (N_2210,N_2181,N_2186);
nand U2211 (N_2211,N_2156,N_2173);
or U2212 (N_2212,N_2175,N_2177);
or U2213 (N_2213,N_2174,N_2197);
or U2214 (N_2214,N_2194,N_2176);
or U2215 (N_2215,N_2155,N_2163);
nor U2216 (N_2216,N_2171,N_2183);
nor U2217 (N_2217,N_2196,N_2157);
nand U2218 (N_2218,N_2179,N_2153);
or U2219 (N_2219,N_2158,N_2187);
nand U2220 (N_2220,N_2190,N_2192);
or U2221 (N_2221,N_2191,N_2184);
and U2222 (N_2222,N_2160,N_2199);
or U2223 (N_2223,N_2172,N_2198);
nor U2224 (N_2224,N_2162,N_2178);
and U2225 (N_2225,N_2152,N_2160);
nor U2226 (N_2226,N_2158,N_2193);
nand U2227 (N_2227,N_2177,N_2158);
nor U2228 (N_2228,N_2169,N_2177);
nand U2229 (N_2229,N_2155,N_2196);
and U2230 (N_2230,N_2154,N_2177);
and U2231 (N_2231,N_2150,N_2180);
or U2232 (N_2232,N_2164,N_2195);
nor U2233 (N_2233,N_2162,N_2151);
and U2234 (N_2234,N_2184,N_2179);
nor U2235 (N_2235,N_2161,N_2186);
xor U2236 (N_2236,N_2174,N_2178);
nand U2237 (N_2237,N_2161,N_2178);
nor U2238 (N_2238,N_2174,N_2161);
nor U2239 (N_2239,N_2152,N_2161);
nand U2240 (N_2240,N_2189,N_2191);
or U2241 (N_2241,N_2184,N_2188);
and U2242 (N_2242,N_2164,N_2152);
and U2243 (N_2243,N_2150,N_2172);
nor U2244 (N_2244,N_2163,N_2156);
nand U2245 (N_2245,N_2199,N_2197);
nand U2246 (N_2246,N_2193,N_2177);
nor U2247 (N_2247,N_2186,N_2199);
nand U2248 (N_2248,N_2168,N_2199);
nand U2249 (N_2249,N_2163,N_2183);
or U2250 (N_2250,N_2212,N_2237);
or U2251 (N_2251,N_2226,N_2207);
or U2252 (N_2252,N_2249,N_2239);
nor U2253 (N_2253,N_2220,N_2205);
or U2254 (N_2254,N_2240,N_2242);
nand U2255 (N_2255,N_2201,N_2247);
nand U2256 (N_2256,N_2219,N_2200);
and U2257 (N_2257,N_2215,N_2235);
nand U2258 (N_2258,N_2246,N_2209);
nand U2259 (N_2259,N_2222,N_2229);
nor U2260 (N_2260,N_2204,N_2231);
nand U2261 (N_2261,N_2228,N_2214);
or U2262 (N_2262,N_2227,N_2230);
and U2263 (N_2263,N_2243,N_2248);
and U2264 (N_2264,N_2244,N_2221);
or U2265 (N_2265,N_2213,N_2225);
nand U2266 (N_2266,N_2236,N_2211);
or U2267 (N_2267,N_2238,N_2224);
nor U2268 (N_2268,N_2202,N_2223);
nand U2269 (N_2269,N_2203,N_2216);
nand U2270 (N_2270,N_2210,N_2233);
or U2271 (N_2271,N_2245,N_2232);
nor U2272 (N_2272,N_2241,N_2234);
or U2273 (N_2273,N_2206,N_2208);
or U2274 (N_2274,N_2217,N_2218);
or U2275 (N_2275,N_2200,N_2229);
or U2276 (N_2276,N_2220,N_2236);
or U2277 (N_2277,N_2234,N_2206);
and U2278 (N_2278,N_2225,N_2229);
nand U2279 (N_2279,N_2212,N_2242);
and U2280 (N_2280,N_2226,N_2242);
and U2281 (N_2281,N_2215,N_2211);
nand U2282 (N_2282,N_2202,N_2230);
or U2283 (N_2283,N_2231,N_2227);
or U2284 (N_2284,N_2207,N_2229);
or U2285 (N_2285,N_2224,N_2221);
or U2286 (N_2286,N_2219,N_2234);
nand U2287 (N_2287,N_2238,N_2227);
or U2288 (N_2288,N_2217,N_2220);
nor U2289 (N_2289,N_2204,N_2241);
xor U2290 (N_2290,N_2231,N_2241);
nand U2291 (N_2291,N_2216,N_2218);
and U2292 (N_2292,N_2207,N_2248);
or U2293 (N_2293,N_2232,N_2229);
nand U2294 (N_2294,N_2236,N_2204);
nand U2295 (N_2295,N_2218,N_2200);
and U2296 (N_2296,N_2233,N_2215);
or U2297 (N_2297,N_2249,N_2217);
or U2298 (N_2298,N_2208,N_2249);
or U2299 (N_2299,N_2242,N_2203);
or U2300 (N_2300,N_2283,N_2251);
or U2301 (N_2301,N_2284,N_2268);
or U2302 (N_2302,N_2273,N_2260);
nand U2303 (N_2303,N_2286,N_2266);
and U2304 (N_2304,N_2269,N_2276);
nor U2305 (N_2305,N_2292,N_2264);
nand U2306 (N_2306,N_2285,N_2256);
xnor U2307 (N_2307,N_2282,N_2274);
or U2308 (N_2308,N_2299,N_2261);
nor U2309 (N_2309,N_2288,N_2293);
nand U2310 (N_2310,N_2296,N_2265);
nand U2311 (N_2311,N_2272,N_2267);
xnor U2312 (N_2312,N_2270,N_2252);
or U2313 (N_2313,N_2275,N_2279);
and U2314 (N_2314,N_2253,N_2259);
nand U2315 (N_2315,N_2258,N_2287);
and U2316 (N_2316,N_2262,N_2255);
and U2317 (N_2317,N_2294,N_2291);
and U2318 (N_2318,N_2257,N_2281);
nand U2319 (N_2319,N_2254,N_2289);
nor U2320 (N_2320,N_2263,N_2280);
or U2321 (N_2321,N_2295,N_2277);
or U2322 (N_2322,N_2297,N_2271);
nor U2323 (N_2323,N_2290,N_2250);
and U2324 (N_2324,N_2278,N_2298);
and U2325 (N_2325,N_2274,N_2279);
and U2326 (N_2326,N_2289,N_2293);
nand U2327 (N_2327,N_2270,N_2293);
nor U2328 (N_2328,N_2276,N_2271);
and U2329 (N_2329,N_2264,N_2272);
or U2330 (N_2330,N_2273,N_2292);
xnor U2331 (N_2331,N_2292,N_2260);
nor U2332 (N_2332,N_2292,N_2291);
and U2333 (N_2333,N_2283,N_2298);
or U2334 (N_2334,N_2285,N_2271);
or U2335 (N_2335,N_2277,N_2256);
and U2336 (N_2336,N_2281,N_2258);
or U2337 (N_2337,N_2274,N_2287);
nor U2338 (N_2338,N_2263,N_2283);
xnor U2339 (N_2339,N_2268,N_2298);
nand U2340 (N_2340,N_2265,N_2275);
and U2341 (N_2341,N_2253,N_2297);
xor U2342 (N_2342,N_2284,N_2259);
and U2343 (N_2343,N_2299,N_2276);
nand U2344 (N_2344,N_2258,N_2259);
nor U2345 (N_2345,N_2251,N_2259);
nor U2346 (N_2346,N_2251,N_2265);
nand U2347 (N_2347,N_2295,N_2252);
or U2348 (N_2348,N_2269,N_2298);
xor U2349 (N_2349,N_2264,N_2258);
and U2350 (N_2350,N_2337,N_2303);
and U2351 (N_2351,N_2322,N_2348);
or U2352 (N_2352,N_2327,N_2323);
and U2353 (N_2353,N_2331,N_2326);
nand U2354 (N_2354,N_2316,N_2314);
or U2355 (N_2355,N_2300,N_2344);
or U2356 (N_2356,N_2332,N_2320);
or U2357 (N_2357,N_2333,N_2341);
nand U2358 (N_2358,N_2305,N_2329);
nor U2359 (N_2359,N_2343,N_2310);
nor U2360 (N_2360,N_2313,N_2346);
nor U2361 (N_2361,N_2302,N_2321);
and U2362 (N_2362,N_2324,N_2336);
or U2363 (N_2363,N_2306,N_2318);
nor U2364 (N_2364,N_2340,N_2345);
or U2365 (N_2365,N_2315,N_2301);
xor U2366 (N_2366,N_2330,N_2319);
nand U2367 (N_2367,N_2308,N_2311);
nand U2368 (N_2368,N_2338,N_2317);
and U2369 (N_2369,N_2349,N_2325);
or U2370 (N_2370,N_2307,N_2334);
or U2371 (N_2371,N_2335,N_2304);
or U2372 (N_2372,N_2339,N_2342);
nand U2373 (N_2373,N_2347,N_2312);
nor U2374 (N_2374,N_2328,N_2309);
or U2375 (N_2375,N_2301,N_2316);
xnor U2376 (N_2376,N_2313,N_2304);
and U2377 (N_2377,N_2318,N_2310);
nor U2378 (N_2378,N_2301,N_2346);
or U2379 (N_2379,N_2326,N_2303);
nand U2380 (N_2380,N_2312,N_2329);
and U2381 (N_2381,N_2334,N_2309);
or U2382 (N_2382,N_2309,N_2306);
nand U2383 (N_2383,N_2324,N_2321);
nor U2384 (N_2384,N_2302,N_2344);
nand U2385 (N_2385,N_2342,N_2340);
nor U2386 (N_2386,N_2331,N_2309);
nand U2387 (N_2387,N_2345,N_2308);
nor U2388 (N_2388,N_2309,N_2333);
and U2389 (N_2389,N_2305,N_2302);
nor U2390 (N_2390,N_2329,N_2330);
xor U2391 (N_2391,N_2323,N_2339);
and U2392 (N_2392,N_2341,N_2313);
or U2393 (N_2393,N_2344,N_2308);
and U2394 (N_2394,N_2330,N_2314);
and U2395 (N_2395,N_2338,N_2309);
nor U2396 (N_2396,N_2335,N_2327);
nor U2397 (N_2397,N_2330,N_2303);
nor U2398 (N_2398,N_2317,N_2309);
and U2399 (N_2399,N_2339,N_2319);
or U2400 (N_2400,N_2395,N_2358);
and U2401 (N_2401,N_2390,N_2363);
and U2402 (N_2402,N_2380,N_2382);
nand U2403 (N_2403,N_2378,N_2359);
or U2404 (N_2404,N_2351,N_2364);
or U2405 (N_2405,N_2379,N_2396);
nor U2406 (N_2406,N_2370,N_2381);
nor U2407 (N_2407,N_2398,N_2355);
nor U2408 (N_2408,N_2365,N_2383);
and U2409 (N_2409,N_2357,N_2367);
or U2410 (N_2410,N_2391,N_2385);
and U2411 (N_2411,N_2384,N_2389);
nand U2412 (N_2412,N_2368,N_2386);
or U2413 (N_2413,N_2373,N_2350);
xnor U2414 (N_2414,N_2353,N_2366);
nand U2415 (N_2415,N_2393,N_2371);
or U2416 (N_2416,N_2377,N_2375);
and U2417 (N_2417,N_2372,N_2354);
nor U2418 (N_2418,N_2356,N_2360);
nand U2419 (N_2419,N_2362,N_2369);
nand U2420 (N_2420,N_2399,N_2361);
or U2421 (N_2421,N_2352,N_2376);
and U2422 (N_2422,N_2388,N_2387);
nand U2423 (N_2423,N_2392,N_2394);
and U2424 (N_2424,N_2397,N_2374);
and U2425 (N_2425,N_2366,N_2388);
and U2426 (N_2426,N_2368,N_2397);
nand U2427 (N_2427,N_2365,N_2399);
nand U2428 (N_2428,N_2378,N_2397);
nand U2429 (N_2429,N_2371,N_2351);
nand U2430 (N_2430,N_2379,N_2376);
and U2431 (N_2431,N_2393,N_2372);
or U2432 (N_2432,N_2382,N_2381);
nand U2433 (N_2433,N_2355,N_2399);
nor U2434 (N_2434,N_2382,N_2396);
or U2435 (N_2435,N_2364,N_2371);
nand U2436 (N_2436,N_2388,N_2350);
and U2437 (N_2437,N_2396,N_2395);
nand U2438 (N_2438,N_2359,N_2396);
and U2439 (N_2439,N_2366,N_2351);
and U2440 (N_2440,N_2374,N_2351);
nand U2441 (N_2441,N_2354,N_2365);
and U2442 (N_2442,N_2360,N_2358);
nor U2443 (N_2443,N_2351,N_2352);
and U2444 (N_2444,N_2374,N_2393);
nor U2445 (N_2445,N_2374,N_2356);
nand U2446 (N_2446,N_2377,N_2398);
nor U2447 (N_2447,N_2364,N_2358);
nor U2448 (N_2448,N_2359,N_2394);
or U2449 (N_2449,N_2364,N_2375);
nand U2450 (N_2450,N_2447,N_2423);
and U2451 (N_2451,N_2433,N_2435);
nand U2452 (N_2452,N_2425,N_2443);
and U2453 (N_2453,N_2431,N_2424);
nor U2454 (N_2454,N_2413,N_2430);
nor U2455 (N_2455,N_2429,N_2440);
or U2456 (N_2456,N_2410,N_2411);
nand U2457 (N_2457,N_2415,N_2407);
nand U2458 (N_2458,N_2426,N_2439);
and U2459 (N_2459,N_2417,N_2420);
nor U2460 (N_2460,N_2406,N_2422);
nor U2461 (N_2461,N_2409,N_2437);
nand U2462 (N_2462,N_2444,N_2408);
or U2463 (N_2463,N_2412,N_2449);
nand U2464 (N_2464,N_2400,N_2442);
and U2465 (N_2465,N_2414,N_2448);
or U2466 (N_2466,N_2402,N_2416);
nor U2467 (N_2467,N_2404,N_2418);
nand U2468 (N_2468,N_2428,N_2432);
or U2469 (N_2469,N_2419,N_2446);
nor U2470 (N_2470,N_2436,N_2441);
nand U2471 (N_2471,N_2438,N_2427);
nand U2472 (N_2472,N_2421,N_2401);
nand U2473 (N_2473,N_2403,N_2405);
nor U2474 (N_2474,N_2445,N_2434);
nand U2475 (N_2475,N_2425,N_2411);
nor U2476 (N_2476,N_2400,N_2402);
or U2477 (N_2477,N_2429,N_2443);
nor U2478 (N_2478,N_2436,N_2401);
nor U2479 (N_2479,N_2433,N_2425);
nand U2480 (N_2480,N_2404,N_2435);
nand U2481 (N_2481,N_2410,N_2413);
or U2482 (N_2482,N_2407,N_2418);
nor U2483 (N_2483,N_2449,N_2438);
or U2484 (N_2484,N_2410,N_2446);
nand U2485 (N_2485,N_2431,N_2442);
or U2486 (N_2486,N_2441,N_2431);
and U2487 (N_2487,N_2421,N_2438);
nor U2488 (N_2488,N_2409,N_2427);
nor U2489 (N_2489,N_2428,N_2407);
or U2490 (N_2490,N_2403,N_2445);
nand U2491 (N_2491,N_2405,N_2419);
and U2492 (N_2492,N_2438,N_2415);
nand U2493 (N_2493,N_2402,N_2448);
nand U2494 (N_2494,N_2429,N_2446);
xor U2495 (N_2495,N_2432,N_2429);
nand U2496 (N_2496,N_2406,N_2410);
nand U2497 (N_2497,N_2447,N_2415);
nand U2498 (N_2498,N_2435,N_2400);
nand U2499 (N_2499,N_2408,N_2420);
xnor U2500 (N_2500,N_2474,N_2450);
nand U2501 (N_2501,N_2462,N_2480);
nor U2502 (N_2502,N_2496,N_2466);
nor U2503 (N_2503,N_2458,N_2486);
nand U2504 (N_2504,N_2464,N_2492);
and U2505 (N_2505,N_2468,N_2471);
or U2506 (N_2506,N_2454,N_2473);
or U2507 (N_2507,N_2476,N_2452);
or U2508 (N_2508,N_2484,N_2475);
or U2509 (N_2509,N_2465,N_2477);
and U2510 (N_2510,N_2463,N_2497);
and U2511 (N_2511,N_2467,N_2489);
nor U2512 (N_2512,N_2487,N_2478);
and U2513 (N_2513,N_2455,N_2460);
nor U2514 (N_2514,N_2472,N_2483);
nand U2515 (N_2515,N_2461,N_2485);
nor U2516 (N_2516,N_2453,N_2495);
nor U2517 (N_2517,N_2499,N_2494);
nor U2518 (N_2518,N_2470,N_2451);
or U2519 (N_2519,N_2469,N_2491);
nor U2520 (N_2520,N_2459,N_2488);
nand U2521 (N_2521,N_2490,N_2481);
nand U2522 (N_2522,N_2457,N_2456);
or U2523 (N_2523,N_2493,N_2498);
and U2524 (N_2524,N_2479,N_2482);
or U2525 (N_2525,N_2492,N_2457);
nor U2526 (N_2526,N_2499,N_2470);
and U2527 (N_2527,N_2497,N_2450);
or U2528 (N_2528,N_2479,N_2495);
or U2529 (N_2529,N_2457,N_2477);
nand U2530 (N_2530,N_2479,N_2498);
or U2531 (N_2531,N_2459,N_2497);
and U2532 (N_2532,N_2453,N_2480);
or U2533 (N_2533,N_2495,N_2457);
nand U2534 (N_2534,N_2456,N_2484);
nor U2535 (N_2535,N_2478,N_2457);
nor U2536 (N_2536,N_2465,N_2488);
nor U2537 (N_2537,N_2493,N_2488);
nor U2538 (N_2538,N_2467,N_2474);
and U2539 (N_2539,N_2469,N_2460);
nand U2540 (N_2540,N_2466,N_2493);
or U2541 (N_2541,N_2490,N_2482);
nor U2542 (N_2542,N_2464,N_2479);
or U2543 (N_2543,N_2468,N_2475);
and U2544 (N_2544,N_2492,N_2489);
or U2545 (N_2545,N_2470,N_2459);
nor U2546 (N_2546,N_2468,N_2462);
or U2547 (N_2547,N_2470,N_2458);
nand U2548 (N_2548,N_2484,N_2467);
and U2549 (N_2549,N_2469,N_2466);
or U2550 (N_2550,N_2545,N_2531);
nand U2551 (N_2551,N_2532,N_2524);
nand U2552 (N_2552,N_2520,N_2507);
nand U2553 (N_2553,N_2519,N_2528);
and U2554 (N_2554,N_2527,N_2548);
or U2555 (N_2555,N_2546,N_2513);
or U2556 (N_2556,N_2542,N_2530);
nor U2557 (N_2557,N_2504,N_2506);
or U2558 (N_2558,N_2511,N_2529);
and U2559 (N_2559,N_2505,N_2541);
nor U2560 (N_2560,N_2534,N_2547);
or U2561 (N_2561,N_2517,N_2537);
or U2562 (N_2562,N_2514,N_2533);
and U2563 (N_2563,N_2538,N_2512);
nand U2564 (N_2564,N_2549,N_2502);
or U2565 (N_2565,N_2503,N_2525);
nor U2566 (N_2566,N_2500,N_2516);
nand U2567 (N_2567,N_2515,N_2508);
nand U2568 (N_2568,N_2536,N_2510);
nand U2569 (N_2569,N_2535,N_2543);
nor U2570 (N_2570,N_2518,N_2522);
nand U2571 (N_2571,N_2539,N_2501);
or U2572 (N_2572,N_2523,N_2509);
nand U2573 (N_2573,N_2526,N_2540);
nor U2574 (N_2574,N_2544,N_2521);
or U2575 (N_2575,N_2541,N_2542);
and U2576 (N_2576,N_2548,N_2533);
and U2577 (N_2577,N_2529,N_2503);
nand U2578 (N_2578,N_2535,N_2526);
or U2579 (N_2579,N_2512,N_2520);
nand U2580 (N_2580,N_2523,N_2525);
and U2581 (N_2581,N_2536,N_2529);
nor U2582 (N_2582,N_2523,N_2508);
and U2583 (N_2583,N_2532,N_2549);
or U2584 (N_2584,N_2534,N_2525);
or U2585 (N_2585,N_2531,N_2516);
or U2586 (N_2586,N_2545,N_2540);
or U2587 (N_2587,N_2511,N_2516);
nor U2588 (N_2588,N_2506,N_2539);
and U2589 (N_2589,N_2505,N_2518);
and U2590 (N_2590,N_2518,N_2510);
and U2591 (N_2591,N_2518,N_2506);
nor U2592 (N_2592,N_2501,N_2513);
nor U2593 (N_2593,N_2546,N_2514);
nor U2594 (N_2594,N_2544,N_2509);
and U2595 (N_2595,N_2541,N_2539);
or U2596 (N_2596,N_2539,N_2543);
nand U2597 (N_2597,N_2549,N_2538);
nor U2598 (N_2598,N_2501,N_2547);
and U2599 (N_2599,N_2543,N_2515);
nor U2600 (N_2600,N_2592,N_2584);
nor U2601 (N_2601,N_2586,N_2593);
and U2602 (N_2602,N_2567,N_2550);
nand U2603 (N_2603,N_2595,N_2562);
nand U2604 (N_2604,N_2555,N_2553);
or U2605 (N_2605,N_2580,N_2599);
nor U2606 (N_2606,N_2583,N_2574);
or U2607 (N_2607,N_2576,N_2559);
or U2608 (N_2608,N_2585,N_2578);
xnor U2609 (N_2609,N_2551,N_2552);
nor U2610 (N_2610,N_2579,N_2590);
nor U2611 (N_2611,N_2598,N_2558);
and U2612 (N_2612,N_2581,N_2588);
nand U2613 (N_2613,N_2556,N_2570);
nor U2614 (N_2614,N_2557,N_2565);
nor U2615 (N_2615,N_2577,N_2597);
and U2616 (N_2616,N_2572,N_2569);
nand U2617 (N_2617,N_2591,N_2594);
or U2618 (N_2618,N_2560,N_2573);
or U2619 (N_2619,N_2587,N_2596);
or U2620 (N_2620,N_2575,N_2568);
nor U2621 (N_2621,N_2571,N_2561);
nand U2622 (N_2622,N_2554,N_2582);
nor U2623 (N_2623,N_2566,N_2563);
nor U2624 (N_2624,N_2589,N_2564);
and U2625 (N_2625,N_2587,N_2598);
nand U2626 (N_2626,N_2561,N_2599);
or U2627 (N_2627,N_2589,N_2572);
nor U2628 (N_2628,N_2562,N_2579);
and U2629 (N_2629,N_2556,N_2598);
and U2630 (N_2630,N_2550,N_2558);
and U2631 (N_2631,N_2559,N_2580);
and U2632 (N_2632,N_2563,N_2591);
and U2633 (N_2633,N_2576,N_2565);
nor U2634 (N_2634,N_2579,N_2552);
or U2635 (N_2635,N_2555,N_2587);
or U2636 (N_2636,N_2587,N_2586);
nor U2637 (N_2637,N_2571,N_2591);
and U2638 (N_2638,N_2595,N_2588);
and U2639 (N_2639,N_2587,N_2557);
or U2640 (N_2640,N_2585,N_2571);
nand U2641 (N_2641,N_2599,N_2596);
and U2642 (N_2642,N_2552,N_2558);
and U2643 (N_2643,N_2596,N_2583);
or U2644 (N_2644,N_2594,N_2563);
nor U2645 (N_2645,N_2578,N_2586);
or U2646 (N_2646,N_2563,N_2571);
nand U2647 (N_2647,N_2561,N_2556);
or U2648 (N_2648,N_2565,N_2554);
nand U2649 (N_2649,N_2555,N_2575);
nand U2650 (N_2650,N_2612,N_2620);
or U2651 (N_2651,N_2645,N_2601);
nand U2652 (N_2652,N_2606,N_2649);
nand U2653 (N_2653,N_2629,N_2624);
or U2654 (N_2654,N_2635,N_2637);
or U2655 (N_2655,N_2639,N_2614);
and U2656 (N_2656,N_2618,N_2627);
nor U2657 (N_2657,N_2610,N_2647);
or U2658 (N_2658,N_2607,N_2642);
nor U2659 (N_2659,N_2615,N_2640);
nor U2660 (N_2660,N_2638,N_2619);
nor U2661 (N_2661,N_2603,N_2628);
or U2662 (N_2662,N_2636,N_2634);
or U2663 (N_2663,N_2622,N_2641);
nand U2664 (N_2664,N_2623,N_2633);
or U2665 (N_2665,N_2602,N_2608);
and U2666 (N_2666,N_2631,N_2632);
nor U2667 (N_2667,N_2617,N_2643);
or U2668 (N_2668,N_2616,N_2611);
and U2669 (N_2669,N_2625,N_2604);
nand U2670 (N_2670,N_2600,N_2621);
nand U2671 (N_2671,N_2646,N_2626);
nand U2672 (N_2672,N_2644,N_2648);
xor U2673 (N_2673,N_2609,N_2613);
or U2674 (N_2674,N_2630,N_2605);
or U2675 (N_2675,N_2640,N_2643);
nor U2676 (N_2676,N_2610,N_2628);
or U2677 (N_2677,N_2625,N_2621);
or U2678 (N_2678,N_2611,N_2625);
and U2679 (N_2679,N_2639,N_2644);
or U2680 (N_2680,N_2645,N_2642);
nand U2681 (N_2681,N_2628,N_2643);
xnor U2682 (N_2682,N_2643,N_2647);
and U2683 (N_2683,N_2601,N_2646);
and U2684 (N_2684,N_2648,N_2607);
nand U2685 (N_2685,N_2603,N_2634);
nand U2686 (N_2686,N_2623,N_2604);
or U2687 (N_2687,N_2626,N_2613);
and U2688 (N_2688,N_2600,N_2627);
nand U2689 (N_2689,N_2626,N_2604);
or U2690 (N_2690,N_2610,N_2648);
or U2691 (N_2691,N_2627,N_2641);
and U2692 (N_2692,N_2601,N_2622);
and U2693 (N_2693,N_2645,N_2630);
nor U2694 (N_2694,N_2645,N_2638);
nand U2695 (N_2695,N_2608,N_2619);
or U2696 (N_2696,N_2606,N_2636);
and U2697 (N_2697,N_2622,N_2630);
nand U2698 (N_2698,N_2626,N_2618);
nand U2699 (N_2699,N_2649,N_2614);
nor U2700 (N_2700,N_2691,N_2654);
nor U2701 (N_2701,N_2697,N_2659);
or U2702 (N_2702,N_2661,N_2670);
nor U2703 (N_2703,N_2688,N_2667);
nor U2704 (N_2704,N_2678,N_2696);
and U2705 (N_2705,N_2660,N_2655);
and U2706 (N_2706,N_2692,N_2693);
nor U2707 (N_2707,N_2669,N_2676);
or U2708 (N_2708,N_2662,N_2690);
or U2709 (N_2709,N_2677,N_2698);
nand U2710 (N_2710,N_2699,N_2658);
nand U2711 (N_2711,N_2653,N_2664);
nor U2712 (N_2712,N_2681,N_2665);
and U2713 (N_2713,N_2674,N_2680);
nor U2714 (N_2714,N_2695,N_2679);
xnor U2715 (N_2715,N_2684,N_2685);
nor U2716 (N_2716,N_2652,N_2657);
and U2717 (N_2717,N_2650,N_2673);
nand U2718 (N_2718,N_2694,N_2682);
nor U2719 (N_2719,N_2672,N_2668);
and U2720 (N_2720,N_2666,N_2683);
nor U2721 (N_2721,N_2671,N_2689);
nor U2722 (N_2722,N_2675,N_2686);
or U2723 (N_2723,N_2687,N_2656);
and U2724 (N_2724,N_2663,N_2651);
or U2725 (N_2725,N_2659,N_2670);
or U2726 (N_2726,N_2652,N_2678);
nand U2727 (N_2727,N_2678,N_2693);
or U2728 (N_2728,N_2669,N_2666);
nor U2729 (N_2729,N_2699,N_2690);
or U2730 (N_2730,N_2693,N_2661);
and U2731 (N_2731,N_2691,N_2657);
nand U2732 (N_2732,N_2686,N_2654);
nand U2733 (N_2733,N_2666,N_2678);
or U2734 (N_2734,N_2693,N_2679);
and U2735 (N_2735,N_2695,N_2668);
nand U2736 (N_2736,N_2691,N_2687);
nor U2737 (N_2737,N_2698,N_2672);
and U2738 (N_2738,N_2656,N_2681);
and U2739 (N_2739,N_2667,N_2674);
nor U2740 (N_2740,N_2690,N_2681);
and U2741 (N_2741,N_2680,N_2692);
nor U2742 (N_2742,N_2684,N_2653);
nand U2743 (N_2743,N_2689,N_2676);
or U2744 (N_2744,N_2661,N_2690);
and U2745 (N_2745,N_2657,N_2690);
nand U2746 (N_2746,N_2656,N_2688);
nor U2747 (N_2747,N_2655,N_2684);
and U2748 (N_2748,N_2699,N_2688);
nand U2749 (N_2749,N_2667,N_2651);
and U2750 (N_2750,N_2748,N_2730);
nor U2751 (N_2751,N_2735,N_2716);
nor U2752 (N_2752,N_2736,N_2705);
and U2753 (N_2753,N_2745,N_2724);
and U2754 (N_2754,N_2701,N_2728);
nand U2755 (N_2755,N_2737,N_2723);
nand U2756 (N_2756,N_2733,N_2702);
nor U2757 (N_2757,N_2704,N_2746);
nor U2758 (N_2758,N_2742,N_2712);
nor U2759 (N_2759,N_2715,N_2707);
nand U2760 (N_2760,N_2721,N_2725);
nor U2761 (N_2761,N_2710,N_2706);
or U2762 (N_2762,N_2727,N_2738);
xnor U2763 (N_2763,N_2741,N_2722);
and U2764 (N_2764,N_2703,N_2749);
nor U2765 (N_2765,N_2740,N_2714);
and U2766 (N_2766,N_2731,N_2747);
nand U2767 (N_2767,N_2732,N_2739);
nand U2768 (N_2768,N_2743,N_2729);
nand U2769 (N_2769,N_2718,N_2744);
or U2770 (N_2770,N_2717,N_2719);
xnor U2771 (N_2771,N_2708,N_2726);
nor U2772 (N_2772,N_2711,N_2700);
or U2773 (N_2773,N_2709,N_2734);
and U2774 (N_2774,N_2713,N_2720);
and U2775 (N_2775,N_2734,N_2721);
nor U2776 (N_2776,N_2746,N_2703);
nand U2777 (N_2777,N_2734,N_2739);
or U2778 (N_2778,N_2742,N_2731);
and U2779 (N_2779,N_2745,N_2726);
and U2780 (N_2780,N_2747,N_2725);
or U2781 (N_2781,N_2701,N_2719);
or U2782 (N_2782,N_2744,N_2749);
nor U2783 (N_2783,N_2708,N_2710);
and U2784 (N_2784,N_2745,N_2729);
or U2785 (N_2785,N_2718,N_2720);
nand U2786 (N_2786,N_2736,N_2714);
nand U2787 (N_2787,N_2715,N_2720);
nand U2788 (N_2788,N_2725,N_2718);
and U2789 (N_2789,N_2742,N_2715);
and U2790 (N_2790,N_2703,N_2724);
nor U2791 (N_2791,N_2737,N_2717);
and U2792 (N_2792,N_2730,N_2742);
or U2793 (N_2793,N_2733,N_2741);
or U2794 (N_2794,N_2736,N_2723);
nand U2795 (N_2795,N_2746,N_2707);
nand U2796 (N_2796,N_2725,N_2713);
or U2797 (N_2797,N_2726,N_2749);
nor U2798 (N_2798,N_2726,N_2721);
or U2799 (N_2799,N_2743,N_2744);
and U2800 (N_2800,N_2763,N_2783);
and U2801 (N_2801,N_2796,N_2779);
nor U2802 (N_2802,N_2758,N_2773);
nand U2803 (N_2803,N_2775,N_2765);
nand U2804 (N_2804,N_2788,N_2759);
and U2805 (N_2805,N_2787,N_2791);
nor U2806 (N_2806,N_2781,N_2754);
nand U2807 (N_2807,N_2760,N_2785);
nand U2808 (N_2808,N_2772,N_2789);
nor U2809 (N_2809,N_2795,N_2792);
nor U2810 (N_2810,N_2756,N_2793);
nand U2811 (N_2811,N_2768,N_2776);
nand U2812 (N_2812,N_2798,N_2786);
or U2813 (N_2813,N_2799,N_2761);
nor U2814 (N_2814,N_2750,N_2777);
nand U2815 (N_2815,N_2757,N_2752);
or U2816 (N_2816,N_2764,N_2769);
nand U2817 (N_2817,N_2784,N_2767);
and U2818 (N_2818,N_2797,N_2762);
nand U2819 (N_2819,N_2753,N_2794);
nand U2820 (N_2820,N_2751,N_2780);
or U2821 (N_2821,N_2770,N_2771);
nand U2822 (N_2822,N_2782,N_2774);
and U2823 (N_2823,N_2790,N_2778);
nor U2824 (N_2824,N_2755,N_2766);
and U2825 (N_2825,N_2784,N_2794);
nor U2826 (N_2826,N_2781,N_2789);
or U2827 (N_2827,N_2774,N_2752);
nand U2828 (N_2828,N_2777,N_2776);
nor U2829 (N_2829,N_2781,N_2785);
and U2830 (N_2830,N_2774,N_2771);
nand U2831 (N_2831,N_2771,N_2782);
and U2832 (N_2832,N_2771,N_2784);
nor U2833 (N_2833,N_2766,N_2753);
or U2834 (N_2834,N_2766,N_2758);
or U2835 (N_2835,N_2767,N_2750);
and U2836 (N_2836,N_2756,N_2794);
and U2837 (N_2837,N_2795,N_2793);
nor U2838 (N_2838,N_2792,N_2783);
nand U2839 (N_2839,N_2764,N_2790);
nand U2840 (N_2840,N_2790,N_2787);
nor U2841 (N_2841,N_2788,N_2763);
or U2842 (N_2842,N_2788,N_2761);
and U2843 (N_2843,N_2762,N_2775);
nor U2844 (N_2844,N_2794,N_2790);
and U2845 (N_2845,N_2779,N_2766);
and U2846 (N_2846,N_2767,N_2764);
and U2847 (N_2847,N_2798,N_2779);
nor U2848 (N_2848,N_2764,N_2792);
or U2849 (N_2849,N_2797,N_2795);
or U2850 (N_2850,N_2847,N_2836);
and U2851 (N_2851,N_2849,N_2808);
nor U2852 (N_2852,N_2828,N_2824);
nor U2853 (N_2853,N_2821,N_2812);
and U2854 (N_2854,N_2832,N_2846);
nand U2855 (N_2855,N_2815,N_2819);
and U2856 (N_2856,N_2833,N_2802);
nor U2857 (N_2857,N_2843,N_2806);
nor U2858 (N_2858,N_2800,N_2844);
nor U2859 (N_2859,N_2840,N_2801);
or U2860 (N_2860,N_2839,N_2822);
and U2861 (N_2861,N_2825,N_2813);
nor U2862 (N_2862,N_2820,N_2827);
nor U2863 (N_2863,N_2818,N_2835);
and U2864 (N_2864,N_2816,N_2803);
nor U2865 (N_2865,N_2830,N_2807);
nor U2866 (N_2866,N_2838,N_2841);
or U2867 (N_2867,N_2834,N_2809);
nand U2868 (N_2868,N_2837,N_2848);
and U2869 (N_2869,N_2845,N_2811);
or U2870 (N_2870,N_2817,N_2842);
nand U2871 (N_2871,N_2805,N_2826);
nand U2872 (N_2872,N_2814,N_2829);
or U2873 (N_2873,N_2810,N_2804);
or U2874 (N_2874,N_2823,N_2831);
nand U2875 (N_2875,N_2815,N_2846);
or U2876 (N_2876,N_2842,N_2836);
nor U2877 (N_2877,N_2804,N_2833);
nand U2878 (N_2878,N_2843,N_2811);
or U2879 (N_2879,N_2845,N_2829);
nor U2880 (N_2880,N_2834,N_2813);
nor U2881 (N_2881,N_2808,N_2837);
nand U2882 (N_2882,N_2809,N_2807);
or U2883 (N_2883,N_2842,N_2802);
nor U2884 (N_2884,N_2842,N_2830);
xor U2885 (N_2885,N_2806,N_2838);
nor U2886 (N_2886,N_2825,N_2838);
or U2887 (N_2887,N_2823,N_2801);
xnor U2888 (N_2888,N_2814,N_2818);
or U2889 (N_2889,N_2842,N_2848);
nand U2890 (N_2890,N_2805,N_2842);
nand U2891 (N_2891,N_2823,N_2849);
nand U2892 (N_2892,N_2805,N_2848);
and U2893 (N_2893,N_2813,N_2843);
nor U2894 (N_2894,N_2821,N_2841);
nor U2895 (N_2895,N_2820,N_2816);
nand U2896 (N_2896,N_2836,N_2820);
nor U2897 (N_2897,N_2826,N_2821);
nand U2898 (N_2898,N_2838,N_2805);
or U2899 (N_2899,N_2842,N_2808);
or U2900 (N_2900,N_2879,N_2891);
nor U2901 (N_2901,N_2866,N_2852);
or U2902 (N_2902,N_2857,N_2859);
nor U2903 (N_2903,N_2878,N_2882);
nand U2904 (N_2904,N_2870,N_2893);
nand U2905 (N_2905,N_2850,N_2877);
nand U2906 (N_2906,N_2851,N_2854);
nand U2907 (N_2907,N_2863,N_2895);
or U2908 (N_2908,N_2864,N_2890);
nand U2909 (N_2909,N_2886,N_2856);
and U2910 (N_2910,N_2867,N_2899);
nand U2911 (N_2911,N_2894,N_2873);
or U2912 (N_2912,N_2868,N_2887);
nand U2913 (N_2913,N_2855,N_2874);
nand U2914 (N_2914,N_2884,N_2871);
or U2915 (N_2915,N_2889,N_2865);
nor U2916 (N_2916,N_2881,N_2876);
or U2917 (N_2917,N_2875,N_2898);
or U2918 (N_2918,N_2869,N_2883);
or U2919 (N_2919,N_2885,N_2880);
or U2920 (N_2920,N_2862,N_2860);
xnor U2921 (N_2921,N_2888,N_2858);
xor U2922 (N_2922,N_2897,N_2892);
nand U2923 (N_2923,N_2853,N_2896);
nand U2924 (N_2924,N_2872,N_2861);
or U2925 (N_2925,N_2869,N_2876);
nand U2926 (N_2926,N_2862,N_2880);
nand U2927 (N_2927,N_2871,N_2853);
nor U2928 (N_2928,N_2890,N_2884);
nand U2929 (N_2929,N_2853,N_2878);
nand U2930 (N_2930,N_2860,N_2884);
nor U2931 (N_2931,N_2881,N_2891);
nor U2932 (N_2932,N_2887,N_2852);
and U2933 (N_2933,N_2881,N_2879);
or U2934 (N_2934,N_2891,N_2883);
nor U2935 (N_2935,N_2879,N_2896);
nor U2936 (N_2936,N_2878,N_2854);
and U2937 (N_2937,N_2869,N_2881);
or U2938 (N_2938,N_2897,N_2887);
and U2939 (N_2939,N_2859,N_2891);
or U2940 (N_2940,N_2874,N_2858);
nand U2941 (N_2941,N_2899,N_2883);
and U2942 (N_2942,N_2863,N_2896);
or U2943 (N_2943,N_2879,N_2863);
nor U2944 (N_2944,N_2869,N_2886);
nor U2945 (N_2945,N_2877,N_2859);
nand U2946 (N_2946,N_2873,N_2855);
and U2947 (N_2947,N_2864,N_2897);
nor U2948 (N_2948,N_2882,N_2867);
nor U2949 (N_2949,N_2896,N_2859);
nand U2950 (N_2950,N_2938,N_2924);
nor U2951 (N_2951,N_2904,N_2900);
nand U2952 (N_2952,N_2921,N_2901);
or U2953 (N_2953,N_2932,N_2949);
nand U2954 (N_2954,N_2930,N_2948);
xor U2955 (N_2955,N_2905,N_2908);
or U2956 (N_2956,N_2936,N_2942);
and U2957 (N_2957,N_2903,N_2941);
or U2958 (N_2958,N_2920,N_2946);
or U2959 (N_2959,N_2939,N_2935);
or U2960 (N_2960,N_2927,N_2928);
and U2961 (N_2961,N_2914,N_2915);
or U2962 (N_2962,N_2906,N_2945);
and U2963 (N_2963,N_2925,N_2916);
nor U2964 (N_2964,N_2926,N_2922);
nand U2965 (N_2965,N_2923,N_2910);
or U2966 (N_2966,N_2913,N_2931);
nor U2967 (N_2967,N_2934,N_2933);
nand U2968 (N_2968,N_2911,N_2944);
and U2969 (N_2969,N_2907,N_2909);
nand U2970 (N_2970,N_2902,N_2912);
nand U2971 (N_2971,N_2937,N_2918);
and U2972 (N_2972,N_2947,N_2929);
nand U2973 (N_2973,N_2919,N_2943);
nand U2974 (N_2974,N_2940,N_2917);
nor U2975 (N_2975,N_2908,N_2901);
nand U2976 (N_2976,N_2917,N_2914);
nor U2977 (N_2977,N_2948,N_2940);
nand U2978 (N_2978,N_2933,N_2912);
and U2979 (N_2979,N_2920,N_2940);
or U2980 (N_2980,N_2918,N_2948);
nand U2981 (N_2981,N_2916,N_2927);
nand U2982 (N_2982,N_2914,N_2908);
or U2983 (N_2983,N_2925,N_2932);
nand U2984 (N_2984,N_2916,N_2921);
nor U2985 (N_2985,N_2949,N_2948);
nand U2986 (N_2986,N_2930,N_2933);
nor U2987 (N_2987,N_2924,N_2928);
nor U2988 (N_2988,N_2948,N_2905);
nor U2989 (N_2989,N_2903,N_2948);
and U2990 (N_2990,N_2939,N_2946);
or U2991 (N_2991,N_2904,N_2942);
and U2992 (N_2992,N_2907,N_2935);
nor U2993 (N_2993,N_2936,N_2904);
nand U2994 (N_2994,N_2915,N_2935);
or U2995 (N_2995,N_2914,N_2923);
and U2996 (N_2996,N_2946,N_2927);
or U2997 (N_2997,N_2915,N_2945);
and U2998 (N_2998,N_2939,N_2938);
or U2999 (N_2999,N_2947,N_2919);
or UO_0 (O_0,N_2973,N_2952);
or UO_1 (O_1,N_2967,N_2966);
and UO_2 (O_2,N_2991,N_2983);
or UO_3 (O_3,N_2990,N_2962);
nand UO_4 (O_4,N_2988,N_2964);
xor UO_5 (O_5,N_2979,N_2994);
or UO_6 (O_6,N_2970,N_2961);
and UO_7 (O_7,N_2953,N_2963);
or UO_8 (O_8,N_2984,N_2993);
nor UO_9 (O_9,N_2978,N_2969);
nand UO_10 (O_10,N_2960,N_2998);
and UO_11 (O_11,N_2951,N_2974);
or UO_12 (O_12,N_2965,N_2959);
or UO_13 (O_13,N_2996,N_2976);
nor UO_14 (O_14,N_2989,N_2985);
nand UO_15 (O_15,N_2995,N_2954);
nand UO_16 (O_16,N_2972,N_2997);
nor UO_17 (O_17,N_2980,N_2975);
nand UO_18 (O_18,N_2982,N_2992);
or UO_19 (O_19,N_2955,N_2956);
nand UO_20 (O_20,N_2986,N_2971);
nand UO_21 (O_21,N_2968,N_2987);
or UO_22 (O_22,N_2999,N_2950);
nor UO_23 (O_23,N_2957,N_2981);
nor UO_24 (O_24,N_2977,N_2958);
nor UO_25 (O_25,N_2961,N_2996);
nor UO_26 (O_26,N_2979,N_2984);
or UO_27 (O_27,N_2950,N_2951);
and UO_28 (O_28,N_2963,N_2972);
nor UO_29 (O_29,N_2982,N_2978);
nor UO_30 (O_30,N_2953,N_2960);
nor UO_31 (O_31,N_2970,N_2987);
nor UO_32 (O_32,N_2990,N_2971);
nor UO_33 (O_33,N_2998,N_2955);
or UO_34 (O_34,N_2965,N_2973);
or UO_35 (O_35,N_2964,N_2994);
nor UO_36 (O_36,N_2971,N_2961);
nand UO_37 (O_37,N_2983,N_2986);
nor UO_38 (O_38,N_2970,N_2985);
and UO_39 (O_39,N_2966,N_2972);
xnor UO_40 (O_40,N_2979,N_2958);
and UO_41 (O_41,N_2990,N_2975);
or UO_42 (O_42,N_2974,N_2971);
nand UO_43 (O_43,N_2977,N_2992);
or UO_44 (O_44,N_2961,N_2992);
nor UO_45 (O_45,N_2986,N_2968);
nand UO_46 (O_46,N_2968,N_2988);
nor UO_47 (O_47,N_2993,N_2979);
or UO_48 (O_48,N_2992,N_2952);
and UO_49 (O_49,N_2964,N_2963);
or UO_50 (O_50,N_2950,N_2952);
nand UO_51 (O_51,N_2967,N_2983);
nand UO_52 (O_52,N_2964,N_2962);
and UO_53 (O_53,N_2974,N_2969);
or UO_54 (O_54,N_2991,N_2989);
and UO_55 (O_55,N_2963,N_2950);
or UO_56 (O_56,N_2968,N_2959);
or UO_57 (O_57,N_2970,N_2977);
nand UO_58 (O_58,N_2999,N_2962);
nand UO_59 (O_59,N_2991,N_2970);
or UO_60 (O_60,N_2997,N_2960);
nand UO_61 (O_61,N_2986,N_2960);
or UO_62 (O_62,N_2981,N_2959);
nor UO_63 (O_63,N_2976,N_2980);
nor UO_64 (O_64,N_2984,N_2973);
or UO_65 (O_65,N_2975,N_2953);
or UO_66 (O_66,N_2972,N_2993);
nor UO_67 (O_67,N_2983,N_2960);
nand UO_68 (O_68,N_2958,N_2997);
and UO_69 (O_69,N_2989,N_2992);
nor UO_70 (O_70,N_2992,N_2956);
nor UO_71 (O_71,N_2993,N_2978);
nand UO_72 (O_72,N_2992,N_2963);
or UO_73 (O_73,N_2957,N_2990);
nand UO_74 (O_74,N_2969,N_2959);
nand UO_75 (O_75,N_2959,N_2957);
and UO_76 (O_76,N_2996,N_2995);
nor UO_77 (O_77,N_2980,N_2972);
or UO_78 (O_78,N_2964,N_2983);
and UO_79 (O_79,N_2962,N_2978);
and UO_80 (O_80,N_2999,N_2963);
nor UO_81 (O_81,N_2972,N_2987);
nand UO_82 (O_82,N_2990,N_2959);
nand UO_83 (O_83,N_2996,N_2985);
and UO_84 (O_84,N_2998,N_2975);
nor UO_85 (O_85,N_2997,N_2964);
or UO_86 (O_86,N_2965,N_2975);
nand UO_87 (O_87,N_2962,N_2955);
nand UO_88 (O_88,N_2969,N_2989);
nand UO_89 (O_89,N_2981,N_2963);
or UO_90 (O_90,N_2985,N_2953);
or UO_91 (O_91,N_2991,N_2962);
or UO_92 (O_92,N_2979,N_2981);
or UO_93 (O_93,N_2996,N_2983);
or UO_94 (O_94,N_2999,N_2989);
and UO_95 (O_95,N_2950,N_2980);
or UO_96 (O_96,N_2953,N_2951);
and UO_97 (O_97,N_2974,N_2968);
nor UO_98 (O_98,N_2997,N_2989);
or UO_99 (O_99,N_2977,N_2951);
nand UO_100 (O_100,N_2957,N_2975);
nand UO_101 (O_101,N_2973,N_2991);
nand UO_102 (O_102,N_2995,N_2971);
nor UO_103 (O_103,N_2950,N_2960);
or UO_104 (O_104,N_2984,N_2978);
and UO_105 (O_105,N_2968,N_2993);
nor UO_106 (O_106,N_2999,N_2990);
and UO_107 (O_107,N_2996,N_2955);
or UO_108 (O_108,N_2998,N_2971);
or UO_109 (O_109,N_2963,N_2984);
or UO_110 (O_110,N_2974,N_2980);
or UO_111 (O_111,N_2964,N_2966);
or UO_112 (O_112,N_2993,N_2989);
nor UO_113 (O_113,N_2959,N_2955);
or UO_114 (O_114,N_2985,N_2971);
or UO_115 (O_115,N_2962,N_2956);
nand UO_116 (O_116,N_2981,N_2950);
nand UO_117 (O_117,N_2958,N_2993);
nand UO_118 (O_118,N_2991,N_2965);
or UO_119 (O_119,N_2953,N_2952);
and UO_120 (O_120,N_2993,N_2983);
nor UO_121 (O_121,N_2977,N_2974);
and UO_122 (O_122,N_2996,N_2998);
nor UO_123 (O_123,N_2959,N_2996);
and UO_124 (O_124,N_2951,N_2961);
nor UO_125 (O_125,N_2967,N_2992);
nand UO_126 (O_126,N_2988,N_2980);
nor UO_127 (O_127,N_2988,N_2950);
or UO_128 (O_128,N_2979,N_2954);
nor UO_129 (O_129,N_2956,N_2998);
nor UO_130 (O_130,N_2950,N_2965);
nor UO_131 (O_131,N_2987,N_2963);
or UO_132 (O_132,N_2971,N_2950);
and UO_133 (O_133,N_2970,N_2957);
nor UO_134 (O_134,N_2951,N_2956);
or UO_135 (O_135,N_2990,N_2979);
nor UO_136 (O_136,N_2990,N_2963);
and UO_137 (O_137,N_2997,N_2983);
and UO_138 (O_138,N_2993,N_2960);
nand UO_139 (O_139,N_2974,N_2954);
nor UO_140 (O_140,N_2980,N_2963);
or UO_141 (O_141,N_2971,N_2976);
or UO_142 (O_142,N_2983,N_2969);
nand UO_143 (O_143,N_2974,N_2988);
nand UO_144 (O_144,N_2972,N_2971);
and UO_145 (O_145,N_2950,N_2984);
nor UO_146 (O_146,N_2962,N_2994);
or UO_147 (O_147,N_2983,N_2989);
nand UO_148 (O_148,N_2980,N_2966);
and UO_149 (O_149,N_2953,N_2962);
nor UO_150 (O_150,N_2977,N_2962);
or UO_151 (O_151,N_2966,N_2989);
nand UO_152 (O_152,N_2999,N_2968);
and UO_153 (O_153,N_2996,N_2993);
nor UO_154 (O_154,N_2973,N_2976);
nand UO_155 (O_155,N_2994,N_2995);
nor UO_156 (O_156,N_2975,N_2970);
nor UO_157 (O_157,N_2973,N_2960);
or UO_158 (O_158,N_2989,N_2981);
nand UO_159 (O_159,N_2988,N_2977);
nor UO_160 (O_160,N_2975,N_2962);
and UO_161 (O_161,N_2952,N_2985);
nand UO_162 (O_162,N_2973,N_2964);
nor UO_163 (O_163,N_2952,N_2998);
nand UO_164 (O_164,N_2963,N_2966);
nor UO_165 (O_165,N_2977,N_2996);
and UO_166 (O_166,N_2952,N_2996);
nand UO_167 (O_167,N_2993,N_2977);
nor UO_168 (O_168,N_2956,N_2954);
nand UO_169 (O_169,N_2970,N_2978);
and UO_170 (O_170,N_2990,N_2955);
nand UO_171 (O_171,N_2979,N_2972);
and UO_172 (O_172,N_2984,N_2955);
or UO_173 (O_173,N_2954,N_2952);
and UO_174 (O_174,N_2962,N_2984);
or UO_175 (O_175,N_2998,N_2957);
nand UO_176 (O_176,N_2963,N_2974);
or UO_177 (O_177,N_2956,N_2950);
nor UO_178 (O_178,N_2956,N_2984);
nor UO_179 (O_179,N_2982,N_2993);
or UO_180 (O_180,N_2966,N_2952);
or UO_181 (O_181,N_2968,N_2998);
nand UO_182 (O_182,N_2981,N_2971);
nand UO_183 (O_183,N_2999,N_2984);
nand UO_184 (O_184,N_2959,N_2978);
nand UO_185 (O_185,N_2990,N_2966);
or UO_186 (O_186,N_2990,N_2980);
or UO_187 (O_187,N_2951,N_2964);
and UO_188 (O_188,N_2951,N_2957);
nand UO_189 (O_189,N_2993,N_2992);
nand UO_190 (O_190,N_2981,N_2967);
nor UO_191 (O_191,N_2955,N_2997);
or UO_192 (O_192,N_2950,N_2961);
and UO_193 (O_193,N_2964,N_2981);
or UO_194 (O_194,N_2972,N_2957);
and UO_195 (O_195,N_2951,N_2968);
nand UO_196 (O_196,N_2991,N_2972);
and UO_197 (O_197,N_2980,N_2991);
and UO_198 (O_198,N_2983,N_2994);
nand UO_199 (O_199,N_2965,N_2952);
and UO_200 (O_200,N_2990,N_2976);
or UO_201 (O_201,N_2969,N_2950);
nor UO_202 (O_202,N_2983,N_2981);
and UO_203 (O_203,N_2967,N_2956);
or UO_204 (O_204,N_2988,N_2956);
or UO_205 (O_205,N_2965,N_2970);
or UO_206 (O_206,N_2980,N_2983);
nand UO_207 (O_207,N_2971,N_2966);
and UO_208 (O_208,N_2972,N_2956);
nor UO_209 (O_209,N_2954,N_2978);
or UO_210 (O_210,N_2983,N_2957);
nand UO_211 (O_211,N_2980,N_2993);
or UO_212 (O_212,N_2972,N_2953);
or UO_213 (O_213,N_2989,N_2977);
and UO_214 (O_214,N_2990,N_2984);
and UO_215 (O_215,N_2971,N_2984);
and UO_216 (O_216,N_2972,N_2999);
nand UO_217 (O_217,N_2976,N_2967);
and UO_218 (O_218,N_2975,N_2983);
nand UO_219 (O_219,N_2994,N_2963);
and UO_220 (O_220,N_2994,N_2957);
nor UO_221 (O_221,N_2975,N_2992);
nor UO_222 (O_222,N_2981,N_2953);
or UO_223 (O_223,N_2972,N_2982);
or UO_224 (O_224,N_2994,N_2978);
nand UO_225 (O_225,N_2976,N_2975);
nor UO_226 (O_226,N_2960,N_2982);
nor UO_227 (O_227,N_2962,N_2974);
or UO_228 (O_228,N_2968,N_2960);
and UO_229 (O_229,N_2994,N_2974);
and UO_230 (O_230,N_2980,N_2955);
and UO_231 (O_231,N_2968,N_2985);
nand UO_232 (O_232,N_2969,N_2951);
nor UO_233 (O_233,N_2992,N_2991);
nand UO_234 (O_234,N_2951,N_2991);
xnor UO_235 (O_235,N_2998,N_2976);
or UO_236 (O_236,N_2984,N_2996);
or UO_237 (O_237,N_2996,N_2956);
xnor UO_238 (O_238,N_2959,N_2988);
and UO_239 (O_239,N_2952,N_2977);
or UO_240 (O_240,N_2954,N_2971);
nor UO_241 (O_241,N_2965,N_2981);
nor UO_242 (O_242,N_2962,N_2952);
and UO_243 (O_243,N_2966,N_2959);
nor UO_244 (O_244,N_2956,N_2960);
nor UO_245 (O_245,N_2980,N_2985);
nor UO_246 (O_246,N_2971,N_2968);
nor UO_247 (O_247,N_2952,N_2964);
and UO_248 (O_248,N_2995,N_2960);
or UO_249 (O_249,N_2967,N_2978);
or UO_250 (O_250,N_2999,N_2964);
nand UO_251 (O_251,N_2983,N_2985);
and UO_252 (O_252,N_2971,N_2963);
or UO_253 (O_253,N_2995,N_2980);
nand UO_254 (O_254,N_2996,N_2950);
nor UO_255 (O_255,N_2980,N_2994);
and UO_256 (O_256,N_2967,N_2952);
and UO_257 (O_257,N_2978,N_2980);
nor UO_258 (O_258,N_2979,N_2988);
nor UO_259 (O_259,N_2975,N_2973);
nor UO_260 (O_260,N_2980,N_2977);
and UO_261 (O_261,N_2991,N_2977);
nor UO_262 (O_262,N_2990,N_2977);
nand UO_263 (O_263,N_2975,N_2959);
nor UO_264 (O_264,N_2979,N_2955);
nor UO_265 (O_265,N_2981,N_2958);
or UO_266 (O_266,N_2985,N_2974);
and UO_267 (O_267,N_2972,N_2960);
or UO_268 (O_268,N_2994,N_2951);
nor UO_269 (O_269,N_2956,N_2991);
nor UO_270 (O_270,N_2960,N_2951);
nor UO_271 (O_271,N_2977,N_2987);
and UO_272 (O_272,N_2988,N_2997);
nor UO_273 (O_273,N_2977,N_2979);
nand UO_274 (O_274,N_2959,N_2984);
and UO_275 (O_275,N_2961,N_2962);
nand UO_276 (O_276,N_2957,N_2988);
xnor UO_277 (O_277,N_2982,N_2983);
nor UO_278 (O_278,N_2999,N_2960);
nand UO_279 (O_279,N_2959,N_2953);
or UO_280 (O_280,N_2975,N_2977);
and UO_281 (O_281,N_2967,N_2980);
nand UO_282 (O_282,N_2987,N_2959);
and UO_283 (O_283,N_2960,N_2957);
or UO_284 (O_284,N_2985,N_2961);
or UO_285 (O_285,N_2956,N_2976);
and UO_286 (O_286,N_2995,N_2970);
or UO_287 (O_287,N_2963,N_2978);
xor UO_288 (O_288,N_2967,N_2986);
or UO_289 (O_289,N_2965,N_2989);
or UO_290 (O_290,N_2978,N_2985);
or UO_291 (O_291,N_2959,N_2997);
or UO_292 (O_292,N_2986,N_2997);
or UO_293 (O_293,N_2961,N_2967);
nor UO_294 (O_294,N_2963,N_2997);
and UO_295 (O_295,N_2990,N_2986);
and UO_296 (O_296,N_2997,N_2971);
nor UO_297 (O_297,N_2976,N_2953);
or UO_298 (O_298,N_2984,N_2965);
or UO_299 (O_299,N_2967,N_2989);
nor UO_300 (O_300,N_2989,N_2974);
and UO_301 (O_301,N_2984,N_2964);
and UO_302 (O_302,N_2983,N_2973);
nand UO_303 (O_303,N_2997,N_2954);
nand UO_304 (O_304,N_2996,N_2966);
and UO_305 (O_305,N_2986,N_2975);
nor UO_306 (O_306,N_2961,N_2986);
nor UO_307 (O_307,N_2998,N_2951);
nand UO_308 (O_308,N_2986,N_2984);
or UO_309 (O_309,N_2992,N_2987);
xnor UO_310 (O_310,N_2986,N_2987);
and UO_311 (O_311,N_2950,N_2990);
nand UO_312 (O_312,N_2993,N_2970);
and UO_313 (O_313,N_2958,N_2991);
or UO_314 (O_314,N_2961,N_2963);
or UO_315 (O_315,N_2979,N_2968);
nor UO_316 (O_316,N_2954,N_2966);
nand UO_317 (O_317,N_2988,N_2971);
nand UO_318 (O_318,N_2990,N_2989);
and UO_319 (O_319,N_2989,N_2959);
and UO_320 (O_320,N_2977,N_2999);
and UO_321 (O_321,N_2994,N_2952);
and UO_322 (O_322,N_2981,N_2968);
nand UO_323 (O_323,N_2959,N_2958);
nand UO_324 (O_324,N_2986,N_2965);
and UO_325 (O_325,N_2967,N_2995);
or UO_326 (O_326,N_2971,N_2996);
xnor UO_327 (O_327,N_2953,N_2986);
nor UO_328 (O_328,N_2979,N_2998);
nor UO_329 (O_329,N_2976,N_2974);
and UO_330 (O_330,N_2989,N_2982);
and UO_331 (O_331,N_2979,N_2996);
xor UO_332 (O_332,N_2956,N_2964);
nand UO_333 (O_333,N_2969,N_2963);
and UO_334 (O_334,N_2990,N_2981);
nand UO_335 (O_335,N_2962,N_2970);
or UO_336 (O_336,N_2963,N_2967);
and UO_337 (O_337,N_2959,N_2993);
and UO_338 (O_338,N_2992,N_2974);
nand UO_339 (O_339,N_2983,N_2998);
and UO_340 (O_340,N_2965,N_2967);
and UO_341 (O_341,N_2957,N_2987);
and UO_342 (O_342,N_2977,N_2968);
and UO_343 (O_343,N_2991,N_2985);
and UO_344 (O_344,N_2979,N_2995);
and UO_345 (O_345,N_2955,N_2951);
and UO_346 (O_346,N_2969,N_2993);
nand UO_347 (O_347,N_2966,N_2970);
nor UO_348 (O_348,N_2958,N_2983);
nand UO_349 (O_349,N_2978,N_2955);
or UO_350 (O_350,N_2975,N_2966);
and UO_351 (O_351,N_2975,N_2991);
and UO_352 (O_352,N_2957,N_2978);
nand UO_353 (O_353,N_2977,N_2964);
nor UO_354 (O_354,N_2994,N_2990);
nor UO_355 (O_355,N_2956,N_2981);
or UO_356 (O_356,N_2964,N_2971);
or UO_357 (O_357,N_2966,N_2951);
and UO_358 (O_358,N_2979,N_2985);
and UO_359 (O_359,N_2989,N_2980);
nor UO_360 (O_360,N_2983,N_2978);
nand UO_361 (O_361,N_2972,N_2973);
or UO_362 (O_362,N_2980,N_2981);
and UO_363 (O_363,N_2999,N_2991);
and UO_364 (O_364,N_2970,N_2951);
and UO_365 (O_365,N_2985,N_2956);
and UO_366 (O_366,N_2987,N_2974);
nand UO_367 (O_367,N_2976,N_2965);
and UO_368 (O_368,N_2992,N_2994);
nand UO_369 (O_369,N_2951,N_2995);
nor UO_370 (O_370,N_2953,N_2995);
nand UO_371 (O_371,N_2952,N_2960);
nand UO_372 (O_372,N_2974,N_2953);
or UO_373 (O_373,N_2991,N_2978);
or UO_374 (O_374,N_2957,N_2979);
nand UO_375 (O_375,N_2987,N_2999);
and UO_376 (O_376,N_2988,N_2962);
nand UO_377 (O_377,N_2998,N_2977);
nand UO_378 (O_378,N_2978,N_2974);
or UO_379 (O_379,N_2976,N_2999);
and UO_380 (O_380,N_2995,N_2993);
nor UO_381 (O_381,N_2973,N_2955);
nand UO_382 (O_382,N_2957,N_2993);
nor UO_383 (O_383,N_2998,N_2965);
nor UO_384 (O_384,N_2996,N_2988);
or UO_385 (O_385,N_2979,N_2950);
nor UO_386 (O_386,N_2990,N_2965);
nand UO_387 (O_387,N_2968,N_2976);
and UO_388 (O_388,N_2956,N_2978);
nor UO_389 (O_389,N_2980,N_2987);
nor UO_390 (O_390,N_2969,N_2996);
nor UO_391 (O_391,N_2958,N_2987);
nor UO_392 (O_392,N_2967,N_2950);
nand UO_393 (O_393,N_2953,N_2993);
or UO_394 (O_394,N_2970,N_2967);
nor UO_395 (O_395,N_2970,N_2952);
or UO_396 (O_396,N_2986,N_2982);
nor UO_397 (O_397,N_2986,N_2959);
and UO_398 (O_398,N_2950,N_2985);
nand UO_399 (O_399,N_2958,N_2961);
nand UO_400 (O_400,N_2977,N_2983);
or UO_401 (O_401,N_2971,N_2993);
or UO_402 (O_402,N_2994,N_2958);
nand UO_403 (O_403,N_2975,N_2960);
or UO_404 (O_404,N_2999,N_2971);
nand UO_405 (O_405,N_2996,N_2957);
or UO_406 (O_406,N_2960,N_2955);
and UO_407 (O_407,N_2960,N_2963);
or UO_408 (O_408,N_2995,N_2957);
and UO_409 (O_409,N_2987,N_2979);
nand UO_410 (O_410,N_2982,N_2984);
nand UO_411 (O_411,N_2950,N_2959);
nor UO_412 (O_412,N_2982,N_2968);
and UO_413 (O_413,N_2976,N_2977);
or UO_414 (O_414,N_2988,N_2991);
or UO_415 (O_415,N_2960,N_2970);
nor UO_416 (O_416,N_2964,N_2974);
nor UO_417 (O_417,N_2953,N_2958);
nor UO_418 (O_418,N_2961,N_2955);
nand UO_419 (O_419,N_2985,N_2977);
nor UO_420 (O_420,N_2988,N_2966);
nand UO_421 (O_421,N_2987,N_2954);
nand UO_422 (O_422,N_2982,N_2991);
nand UO_423 (O_423,N_2994,N_2975);
xnor UO_424 (O_424,N_2987,N_2971);
and UO_425 (O_425,N_2988,N_2969);
nand UO_426 (O_426,N_2962,N_2972);
or UO_427 (O_427,N_2999,N_2974);
nor UO_428 (O_428,N_2972,N_2955);
or UO_429 (O_429,N_2953,N_2990);
and UO_430 (O_430,N_2962,N_2971);
nand UO_431 (O_431,N_2992,N_2971);
or UO_432 (O_432,N_2971,N_2994);
nor UO_433 (O_433,N_2972,N_2983);
nor UO_434 (O_434,N_2978,N_2989);
and UO_435 (O_435,N_2954,N_2988);
nor UO_436 (O_436,N_2957,N_2997);
and UO_437 (O_437,N_2964,N_2955);
and UO_438 (O_438,N_2974,N_2983);
nor UO_439 (O_439,N_2976,N_2962);
and UO_440 (O_440,N_2972,N_2974);
or UO_441 (O_441,N_2956,N_2995);
nor UO_442 (O_442,N_2954,N_2967);
and UO_443 (O_443,N_2982,N_2979);
and UO_444 (O_444,N_2953,N_2999);
nor UO_445 (O_445,N_2958,N_2982);
nand UO_446 (O_446,N_2977,N_2971);
and UO_447 (O_447,N_2984,N_2980);
or UO_448 (O_448,N_2987,N_2976);
and UO_449 (O_449,N_2961,N_2984);
nor UO_450 (O_450,N_2989,N_2957);
nand UO_451 (O_451,N_2961,N_2993);
or UO_452 (O_452,N_2985,N_2981);
nor UO_453 (O_453,N_2959,N_2985);
nand UO_454 (O_454,N_2996,N_2990);
nand UO_455 (O_455,N_2958,N_2972);
and UO_456 (O_456,N_2988,N_2972);
or UO_457 (O_457,N_2963,N_2965);
nor UO_458 (O_458,N_2976,N_2983);
or UO_459 (O_459,N_2962,N_2996);
nand UO_460 (O_460,N_2956,N_2957);
nor UO_461 (O_461,N_2976,N_2997);
or UO_462 (O_462,N_2987,N_2998);
or UO_463 (O_463,N_2974,N_2982);
and UO_464 (O_464,N_2967,N_2951);
or UO_465 (O_465,N_2954,N_2950);
nor UO_466 (O_466,N_2976,N_2982);
nor UO_467 (O_467,N_2966,N_2998);
and UO_468 (O_468,N_2980,N_2954);
nor UO_469 (O_469,N_2960,N_2990);
nor UO_470 (O_470,N_2973,N_2971);
nand UO_471 (O_471,N_2998,N_2984);
nor UO_472 (O_472,N_2979,N_2970);
and UO_473 (O_473,N_2952,N_2983);
nor UO_474 (O_474,N_2987,N_2956);
nand UO_475 (O_475,N_2986,N_2969);
or UO_476 (O_476,N_2952,N_2989);
or UO_477 (O_477,N_2953,N_2968);
and UO_478 (O_478,N_2973,N_2999);
xnor UO_479 (O_479,N_2977,N_2957);
or UO_480 (O_480,N_2979,N_2960);
nor UO_481 (O_481,N_2960,N_2954);
nand UO_482 (O_482,N_2980,N_2951);
nor UO_483 (O_483,N_2986,N_2998);
nor UO_484 (O_484,N_2968,N_2969);
nand UO_485 (O_485,N_2997,N_2992);
nand UO_486 (O_486,N_2960,N_2964);
and UO_487 (O_487,N_2976,N_2955);
nand UO_488 (O_488,N_2998,N_2964);
or UO_489 (O_489,N_2962,N_2998);
nand UO_490 (O_490,N_2952,N_2958);
nor UO_491 (O_491,N_2965,N_2960);
or UO_492 (O_492,N_2996,N_2999);
and UO_493 (O_493,N_2974,N_2973);
nor UO_494 (O_494,N_2973,N_2967);
or UO_495 (O_495,N_2981,N_2982);
nor UO_496 (O_496,N_2966,N_2979);
and UO_497 (O_497,N_2986,N_2992);
nand UO_498 (O_498,N_2989,N_2987);
nor UO_499 (O_499,N_2973,N_2988);
endmodule