module basic_3000_30000_3500_6_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
and U0 (N_0,In_2452,In_664);
or U1 (N_1,In_1270,In_1069);
and U2 (N_2,In_114,In_1908);
nand U3 (N_3,In_1884,In_1202);
nand U4 (N_4,In_1470,In_1435);
or U5 (N_5,In_915,In_2504);
nor U6 (N_6,In_2316,In_183);
nand U7 (N_7,In_1028,In_1813);
xor U8 (N_8,In_1379,In_2361);
nand U9 (N_9,In_1366,In_916);
nand U10 (N_10,In_2978,In_2917);
nand U11 (N_11,In_105,In_2516);
nor U12 (N_12,In_1231,In_1117);
nor U13 (N_13,In_2616,In_2598);
nor U14 (N_14,In_2337,In_185);
and U15 (N_15,In_2165,In_2861);
xor U16 (N_16,In_1878,In_1585);
nand U17 (N_17,In_2623,In_2354);
and U18 (N_18,In_2118,In_961);
nor U19 (N_19,In_2432,In_1133);
or U20 (N_20,In_315,In_543);
and U21 (N_21,In_1049,In_2517);
nor U22 (N_22,In_1009,In_2735);
nand U23 (N_23,In_1960,In_53);
nand U24 (N_24,In_880,In_608);
nor U25 (N_25,In_1811,In_28);
nor U26 (N_26,In_1828,In_1809);
or U27 (N_27,In_2307,In_485);
or U28 (N_28,In_2987,In_856);
xor U29 (N_29,In_2343,In_2239);
and U30 (N_30,In_1510,In_2017);
or U31 (N_31,In_303,In_1038);
nand U32 (N_32,In_120,In_1999);
and U33 (N_33,In_2761,In_1974);
nor U34 (N_34,In_1113,In_1667);
or U35 (N_35,In_2026,In_2215);
nand U36 (N_36,In_1371,In_513);
and U37 (N_37,In_2086,In_2665);
and U38 (N_38,In_1940,In_1046);
xor U39 (N_39,In_2393,In_907);
nor U40 (N_40,In_1325,In_1968);
or U41 (N_41,In_2711,In_2588);
nor U42 (N_42,In_2553,In_2229);
nor U43 (N_43,In_1319,In_1831);
nand U44 (N_44,In_579,In_1862);
nor U45 (N_45,In_2336,In_1775);
and U46 (N_46,In_2357,In_2374);
or U47 (N_47,In_2851,In_1692);
nor U48 (N_48,In_230,In_1223);
and U49 (N_49,In_770,In_2119);
and U50 (N_50,In_10,In_2944);
nand U51 (N_51,In_1500,In_1336);
and U52 (N_52,In_2673,In_953);
and U53 (N_53,In_1305,In_2403);
nor U54 (N_54,In_2314,In_734);
nor U55 (N_55,In_1750,In_2322);
and U56 (N_56,In_693,In_602);
or U57 (N_57,In_2899,In_470);
nand U58 (N_58,In_1622,In_2979);
and U59 (N_59,In_1827,In_1674);
nor U60 (N_60,In_2214,In_1027);
nand U61 (N_61,In_1715,In_1335);
nor U62 (N_62,In_993,In_1506);
or U63 (N_63,In_2845,In_686);
nor U64 (N_64,In_2089,In_301);
or U65 (N_65,In_223,In_2750);
nor U66 (N_66,In_1517,In_1227);
and U67 (N_67,In_2746,In_1372);
nor U68 (N_68,In_330,In_2100);
nor U69 (N_69,In_2643,In_2251);
and U70 (N_70,In_1147,In_2160);
nor U71 (N_71,In_563,In_591);
and U72 (N_72,In_132,In_595);
nand U73 (N_73,In_2270,In_2480);
nor U74 (N_74,In_86,In_455);
or U75 (N_75,In_1271,In_610);
and U76 (N_76,In_1568,In_827);
xnor U77 (N_77,In_2843,In_932);
nand U78 (N_78,In_2346,In_2727);
nor U79 (N_79,In_1266,In_1785);
and U80 (N_80,In_190,In_484);
nand U81 (N_81,In_1485,In_2953);
and U82 (N_82,In_1628,In_1386);
or U83 (N_83,In_759,In_2175);
and U84 (N_84,In_556,In_2105);
and U85 (N_85,In_2339,In_2684);
or U86 (N_86,In_1612,In_2363);
nand U87 (N_87,In_14,In_1846);
and U88 (N_88,In_1053,In_2454);
nand U89 (N_89,In_1977,In_716);
nand U90 (N_90,In_784,In_2332);
xnor U91 (N_91,In_913,In_531);
or U92 (N_92,In_2325,In_1840);
nand U93 (N_93,In_2563,In_363);
nor U94 (N_94,In_2326,In_1912);
and U95 (N_95,In_2042,In_319);
or U96 (N_96,In_1368,In_1108);
nor U97 (N_97,In_1898,In_831);
nand U98 (N_98,In_722,In_2262);
nand U99 (N_99,In_2341,In_402);
nor U100 (N_100,In_1703,In_769);
and U101 (N_101,In_2369,In_2707);
nor U102 (N_102,In_754,In_1419);
or U103 (N_103,In_2434,In_195);
and U104 (N_104,In_1183,In_701);
and U105 (N_105,In_1519,In_238);
nor U106 (N_106,In_2168,In_1820);
xor U107 (N_107,In_1748,In_1592);
nor U108 (N_108,In_321,In_2367);
and U109 (N_109,In_2744,In_1440);
nand U110 (N_110,In_505,In_2417);
nand U111 (N_111,In_2779,In_72);
and U112 (N_112,In_950,In_518);
nor U113 (N_113,In_1007,In_440);
nand U114 (N_114,In_2862,In_66);
or U115 (N_115,In_903,In_265);
nand U116 (N_116,In_2660,In_1497);
xnor U117 (N_117,In_2968,In_2904);
nand U118 (N_118,In_1173,In_157);
xnor U119 (N_119,In_1758,In_540);
or U120 (N_120,In_1219,In_158);
nand U121 (N_121,In_2304,In_2308);
and U122 (N_122,In_752,In_525);
nor U123 (N_123,In_1503,In_2437);
and U124 (N_124,In_1641,In_2152);
and U125 (N_125,In_963,In_519);
nand U126 (N_126,In_729,In_820);
and U127 (N_127,In_2558,In_2064);
and U128 (N_128,In_1926,In_788);
nor U129 (N_129,In_2489,In_2948);
nand U130 (N_130,In_355,In_925);
and U131 (N_131,In_2267,In_2181);
xor U132 (N_132,In_1545,In_2859);
and U133 (N_133,In_978,In_497);
nand U134 (N_134,In_76,In_351);
nand U135 (N_135,In_2651,In_1561);
and U136 (N_136,In_1239,In_51);
xnor U137 (N_137,In_605,In_1719);
nor U138 (N_138,In_578,In_2233);
nor U139 (N_139,In_2083,In_1670);
or U140 (N_140,In_429,In_109);
nand U141 (N_141,In_2294,In_1559);
nor U142 (N_142,In_2220,In_2219);
nand U143 (N_143,In_2685,In_2945);
or U144 (N_144,In_584,In_1626);
or U145 (N_145,In_1122,In_2209);
nor U146 (N_146,In_1534,In_2018);
and U147 (N_147,In_278,In_30);
or U148 (N_148,In_2578,In_611);
or U149 (N_149,In_302,In_1537);
nor U150 (N_150,In_370,In_914);
nor U151 (N_151,In_2694,In_1564);
nand U152 (N_152,In_457,In_2283);
xor U153 (N_153,In_1005,In_1013);
nand U154 (N_154,In_1983,In_2524);
or U155 (N_155,In_2876,In_273);
nand U156 (N_156,In_2222,In_1552);
and U157 (N_157,In_2533,In_1967);
nor U158 (N_158,In_2221,In_2640);
or U159 (N_159,In_982,In_2243);
and U160 (N_160,In_1502,In_947);
nand U161 (N_161,In_1567,In_2344);
xnor U162 (N_162,In_1839,In_593);
nand U163 (N_163,In_1581,In_1932);
or U164 (N_164,In_1892,In_2523);
and U165 (N_165,In_205,In_1529);
xor U166 (N_166,In_2693,In_361);
nor U167 (N_167,In_2176,In_1041);
nand U168 (N_168,In_821,In_795);
and U169 (N_169,In_1315,In_2531);
or U170 (N_170,In_377,In_2666);
or U171 (N_171,In_2617,In_2129);
xor U172 (N_172,In_1776,In_2249);
nand U173 (N_173,In_755,In_2846);
nor U174 (N_174,In_991,In_1613);
nand U175 (N_175,In_946,In_847);
and U176 (N_176,In_1411,In_2914);
or U177 (N_177,In_168,In_2292);
or U178 (N_178,In_2298,In_2061);
and U179 (N_179,In_2500,In_727);
nand U180 (N_180,In_1021,In_456);
or U181 (N_181,In_2203,In_275);
and U182 (N_182,In_1997,In_2824);
xor U183 (N_183,In_1444,In_150);
nand U184 (N_184,In_2264,In_910);
nand U185 (N_185,In_1420,In_1521);
or U186 (N_186,In_1754,In_2002);
and U187 (N_187,In_1618,In_1237);
and U188 (N_188,In_2498,In_78);
and U189 (N_189,In_2228,In_2946);
and U190 (N_190,In_1321,In_311);
nor U191 (N_191,In_960,In_2592);
or U192 (N_192,In_1658,In_2244);
or U193 (N_193,In_1439,In_1787);
and U194 (N_194,In_433,In_1085);
and U195 (N_195,In_2891,In_2584);
and U196 (N_196,In_2802,In_104);
xnor U197 (N_197,In_804,In_2457);
nand U198 (N_198,In_2536,In_2658);
xor U199 (N_199,In_1701,In_2526);
or U200 (N_200,In_2476,In_2545);
xnor U201 (N_201,In_2525,In_2765);
or U202 (N_202,In_2556,In_2762);
nor U203 (N_203,In_2059,In_2335);
xor U204 (N_204,In_699,In_2225);
nand U205 (N_205,In_994,In_2163);
nor U206 (N_206,In_2712,In_1152);
nor U207 (N_207,In_794,In_2557);
and U208 (N_208,In_1140,In_1904);
or U209 (N_209,In_1697,In_776);
or U210 (N_210,In_622,In_2466);
or U211 (N_211,In_2108,In_706);
nand U212 (N_212,In_1621,In_498);
nand U213 (N_213,In_88,In_2029);
or U214 (N_214,In_1723,In_2157);
or U215 (N_215,In_1128,In_2519);
nand U216 (N_216,In_892,In_2187);
nor U217 (N_217,In_1914,In_121);
and U218 (N_218,In_951,In_1337);
nor U219 (N_219,In_1969,In_1812);
xor U220 (N_220,In_862,In_1412);
or U221 (N_221,In_906,In_2252);
nand U222 (N_222,In_940,In_477);
or U223 (N_223,In_2459,In_669);
and U224 (N_224,In_1293,In_620);
and U225 (N_225,In_1184,In_2966);
xor U226 (N_226,In_1316,In_1415);
or U227 (N_227,In_2709,In_502);
and U228 (N_228,In_1334,In_672);
nand U229 (N_229,In_1851,In_2513);
and U230 (N_230,In_1744,In_1106);
nor U231 (N_231,In_1285,In_1734);
or U232 (N_232,In_2133,In_186);
nand U233 (N_233,In_1772,In_2226);
nor U234 (N_234,In_2759,In_1396);
nor U235 (N_235,In_652,In_170);
nand U236 (N_236,In_1866,In_641);
xor U237 (N_237,In_1931,In_1243);
nand U238 (N_238,In_2833,In_1425);
or U239 (N_239,In_447,In_2716);
xor U240 (N_240,In_550,In_597);
or U241 (N_241,In_2784,In_2602);
nand U242 (N_242,In_472,In_1937);
nand U243 (N_243,In_801,In_1432);
or U244 (N_244,In_825,In_790);
or U245 (N_245,In_735,In_1905);
or U246 (N_246,In_1036,In_1409);
xnor U247 (N_247,In_1845,In_1741);
or U248 (N_248,In_1197,In_2491);
nor U249 (N_249,In_252,In_974);
nor U250 (N_250,In_2079,In_1003);
nor U251 (N_251,In_1870,In_1685);
and U252 (N_252,In_2528,In_2907);
or U253 (N_253,In_2004,In_2241);
nand U254 (N_254,In_2472,In_2597);
nor U255 (N_255,In_2421,In_2412);
nand U256 (N_256,In_2601,In_1076);
nand U257 (N_257,In_852,In_865);
nand U258 (N_258,In_1193,In_352);
or U259 (N_259,In_2991,In_1964);
or U260 (N_260,In_2530,In_1797);
xor U261 (N_261,In_2227,In_2719);
or U262 (N_262,In_1297,In_2134);
or U263 (N_263,In_1201,In_332);
nor U264 (N_264,In_492,In_177);
and U265 (N_265,In_2586,In_684);
nor U266 (N_266,In_182,In_935);
and U267 (N_267,In_2303,In_1216);
nor U268 (N_268,In_2150,In_2806);
or U269 (N_269,In_2698,In_131);
or U270 (N_270,In_399,In_1022);
and U271 (N_271,In_1576,In_1527);
nand U272 (N_272,In_337,In_681);
nand U273 (N_273,In_491,In_2781);
and U274 (N_274,In_524,In_1856);
nor U275 (N_275,In_2425,In_1404);
nor U276 (N_276,In_586,In_341);
xnor U277 (N_277,In_1952,In_692);
nand U278 (N_278,In_1678,In_333);
or U279 (N_279,In_2951,In_860);
nor U280 (N_280,In_1917,In_863);
nor U281 (N_281,In_154,In_1413);
and U282 (N_282,In_1570,In_2136);
nor U283 (N_283,In_2447,In_8);
xnor U284 (N_284,In_1406,In_2723);
nand U285 (N_285,In_79,In_1228);
or U286 (N_286,In_2096,In_743);
or U287 (N_287,In_1338,In_1381);
or U288 (N_288,In_2115,In_2003);
nand U289 (N_289,In_2677,In_115);
and U290 (N_290,In_926,In_1033);
and U291 (N_291,In_165,In_475);
nand U292 (N_292,In_1910,In_2474);
xor U293 (N_293,In_2826,In_1661);
or U294 (N_294,In_589,In_973);
nor U295 (N_295,In_2509,In_1683);
xor U296 (N_296,In_2894,In_738);
xor U297 (N_297,In_1680,In_384);
nand U298 (N_298,In_2844,In_489);
and U299 (N_299,In_680,In_2320);
nand U300 (N_300,In_689,In_2143);
nand U301 (N_301,In_2921,In_313);
and U302 (N_302,In_626,In_2722);
nor U303 (N_303,In_2767,In_2177);
nand U304 (N_304,In_1269,In_293);
xnor U305 (N_305,In_2025,In_2236);
and U306 (N_306,In_1248,In_1345);
nor U307 (N_307,In_2319,In_1669);
and U308 (N_308,In_1764,In_306);
nand U309 (N_309,In_739,In_493);
nand U310 (N_310,In_2550,In_842);
nand U311 (N_311,In_1416,In_1536);
or U312 (N_312,In_2999,In_241);
nand U313 (N_313,In_25,In_2925);
and U314 (N_314,In_1452,In_1948);
xor U315 (N_315,In_1233,In_2928);
or U316 (N_316,In_350,In_221);
nor U317 (N_317,In_1308,In_515);
or U318 (N_318,In_1781,In_733);
nor U319 (N_319,In_2077,In_2200);
nand U320 (N_320,In_836,In_709);
or U321 (N_321,In_2007,In_2488);
or U322 (N_322,In_2146,In_151);
nand U323 (N_323,In_198,In_1126);
nand U324 (N_324,In_2075,In_818);
nand U325 (N_325,In_1720,In_2934);
and U326 (N_326,In_1290,In_1804);
nor U327 (N_327,In_1982,In_31);
nor U328 (N_328,In_69,In_1829);
nor U329 (N_329,In_1174,In_1639);
nor U330 (N_330,In_703,In_685);
nor U331 (N_331,In_425,In_2629);
or U332 (N_332,In_1098,In_1312);
nand U333 (N_333,In_2608,In_335);
nor U334 (N_334,In_232,In_2376);
and U335 (N_335,In_1816,In_2331);
or U336 (N_336,In_812,In_1401);
nor U337 (N_337,In_222,In_2065);
nor U338 (N_338,In_294,In_2382);
xnor U339 (N_339,In_2178,In_2699);
nor U340 (N_340,In_2552,In_172);
nand U341 (N_341,In_799,In_2404);
nand U342 (N_342,In_1916,In_2208);
or U343 (N_343,In_2739,In_2475);
nor U344 (N_344,In_1479,In_928);
nor U345 (N_345,In_2300,In_592);
and U346 (N_346,In_2713,In_1455);
nor U347 (N_347,In_2258,In_1946);
or U348 (N_348,In_676,In_704);
and U349 (N_349,In_412,In_2293);
nor U350 (N_350,In_718,In_126);
xnor U351 (N_351,In_750,In_1257);
nor U352 (N_352,In_1358,In_2099);
nor U353 (N_353,In_1066,In_2855);
nand U354 (N_354,In_854,In_1498);
nor U355 (N_355,In_682,In_2734);
and U356 (N_356,In_828,In_2144);
or U357 (N_357,In_1978,In_869);
and U358 (N_358,In_886,In_1705);
xnor U359 (N_359,In_2772,In_1687);
and U360 (N_360,In_545,In_2755);
and U361 (N_361,In_1189,In_1252);
nor U362 (N_362,In_2438,In_1491);
and U363 (N_363,In_1694,In_2285);
nand U364 (N_364,In_2377,In_1737);
and U365 (N_365,In_1528,In_1514);
nor U366 (N_366,In_103,In_1625);
nor U367 (N_367,In_1708,In_1175);
nand U368 (N_368,In_258,In_1407);
or U369 (N_369,In_2095,In_380);
nand U370 (N_370,In_1143,In_2691);
and U371 (N_371,In_775,In_119);
xnor U372 (N_372,In_1543,In_898);
and U373 (N_373,In_838,In_1588);
and U374 (N_374,In_1689,In_1282);
nor U375 (N_375,In_1422,In_1087);
or U376 (N_376,In_2768,In_2248);
nor U377 (N_377,In_2555,In_145);
xnor U378 (N_378,In_253,In_964);
nand U379 (N_379,In_726,In_1725);
and U380 (N_380,In_1902,In_1918);
nor U381 (N_381,In_1499,In_2675);
nand U382 (N_382,In_1647,In_1037);
nand U383 (N_383,In_1794,In_39);
nand U384 (N_384,In_2977,In_2903);
nand U385 (N_385,In_829,In_127);
or U386 (N_386,In_2047,In_2565);
or U387 (N_387,In_320,In_1774);
nor U388 (N_388,In_2918,In_2170);
nand U389 (N_389,In_1645,In_2471);
and U390 (N_390,In_19,In_647);
or U391 (N_391,In_371,In_582);
nand U392 (N_392,In_1889,In_149);
and U393 (N_393,In_1648,In_2153);
nand U394 (N_394,In_2253,In_1151);
or U395 (N_395,In_2378,In_2192);
nand U396 (N_396,In_290,In_1329);
or U397 (N_397,In_988,In_2087);
nand U398 (N_398,In_958,In_1127);
nor U399 (N_399,In_878,In_1464);
nand U400 (N_400,In_1373,In_1949);
nor U401 (N_401,In_2638,In_1919);
xnor U402 (N_402,In_2439,In_712);
or U403 (N_403,In_2373,In_2287);
xnor U404 (N_404,In_1642,In_2009);
and U405 (N_405,In_437,In_1808);
and U406 (N_406,In_2091,In_1861);
and U407 (N_407,In_503,In_542);
and U408 (N_408,In_888,In_2821);
and U409 (N_409,In_2518,In_2246);
or U410 (N_410,In_2024,In_623);
nand U411 (N_411,In_75,In_2756);
nor U412 (N_412,In_2785,In_1300);
or U413 (N_413,In_2481,In_277);
and U414 (N_414,In_286,In_52);
nand U415 (N_415,In_448,In_378);
nor U416 (N_416,In_1102,In_872);
nor U417 (N_417,In_1991,In_1600);
nor U418 (N_418,In_2700,In_1075);
and U419 (N_419,In_129,In_1759);
and U420 (N_420,In_1296,In_917);
and U421 (N_421,In_1255,In_803);
and U422 (N_422,In_305,In_2281);
nor U423 (N_423,In_264,In_454);
and U424 (N_424,In_1099,In_1939);
or U425 (N_425,In_213,In_34);
nor U426 (N_426,In_336,In_1751);
or U427 (N_427,In_2897,In_1864);
nor U428 (N_428,In_1178,In_1560);
and U429 (N_429,In_67,In_2604);
or U430 (N_430,In_1032,In_2621);
and U431 (N_431,In_1509,In_783);
and U432 (N_432,In_1417,In_1154);
or U433 (N_433,In_668,In_2186);
nor U434 (N_434,In_331,In_1872);
nor U435 (N_435,In_1602,In_97);
nor U436 (N_436,In_2231,In_235);
nand U437 (N_437,In_1801,In_2360);
nand U438 (N_438,In_2841,In_1852);
xnor U439 (N_439,In_2986,In_508);
xnor U440 (N_440,In_632,In_2433);
nand U441 (N_441,In_1765,In_224);
and U442 (N_442,In_1225,In_2541);
or U443 (N_443,In_2884,In_533);
and U444 (N_444,In_816,In_1847);
nand U445 (N_445,In_1520,In_546);
nor U446 (N_446,In_1657,In_662);
and U447 (N_447,In_1426,In_1906);
or U448 (N_448,In_2872,In_1224);
or U449 (N_449,In_2803,In_1617);
nand U450 (N_450,In_2503,In_1267);
nor U451 (N_451,In_259,In_2793);
and U452 (N_452,In_717,In_1100);
xor U453 (N_453,In_102,In_1462);
xor U454 (N_454,In_1798,In_2174);
and U455 (N_455,In_1875,In_1250);
nand U456 (N_456,In_902,In_1788);
and U457 (N_457,In_468,In_1105);
or U458 (N_458,In_2005,In_1465);
nand U459 (N_459,In_2540,In_2817);
nand U460 (N_460,In_857,In_2858);
and U461 (N_461,In_583,In_1273);
xor U462 (N_462,In_1547,In_2849);
xnor U463 (N_463,In_1577,In_1888);
xor U464 (N_464,In_2706,In_2413);
and U465 (N_465,In_389,In_987);
and U466 (N_466,In_547,In_101);
nor U467 (N_467,In_2151,In_2235);
or U468 (N_468,In_2295,In_1423);
and U469 (N_469,In_1103,In_1476);
and U470 (N_470,In_110,In_587);
and U471 (N_471,In_1763,In_1821);
nor U472 (N_472,In_580,In_1504);
and U473 (N_473,In_2166,In_2692);
xor U474 (N_474,In_1256,In_1211);
nand U475 (N_475,In_748,In_562);
or U476 (N_476,In_1015,In_2868);
and U477 (N_477,In_1313,In_61);
or U478 (N_478,In_1574,In_2131);
nor U479 (N_479,In_787,In_2733);
or U480 (N_480,In_2196,In_2291);
xnor U481 (N_481,In_1124,In_2142);
nand U482 (N_482,In_921,In_231);
nor U483 (N_483,In_2959,In_4);
nand U484 (N_484,In_1930,In_713);
and U485 (N_485,In_1850,In_2280);
xor U486 (N_486,In_777,In_1383);
nor U487 (N_487,In_1921,In_488);
nand U488 (N_488,In_809,In_2593);
nor U489 (N_489,In_135,In_2538);
or U490 (N_490,In_1704,In_2139);
or U491 (N_491,In_2266,In_506);
and U492 (N_492,In_1299,In_553);
nand U493 (N_493,In_1279,In_2380);
nand U494 (N_494,In_832,In_1477);
and U495 (N_495,In_1058,In_2050);
and U496 (N_496,In_58,In_873);
nand U497 (N_497,In_2132,In_2112);
xor U498 (N_498,In_141,In_1323);
and U499 (N_499,In_2683,In_2937);
or U500 (N_500,In_1281,In_572);
xor U501 (N_501,In_2282,In_2853);
nor U502 (N_502,In_1017,In_2747);
nand U503 (N_503,In_2117,In_469);
and U504 (N_504,In_939,In_1168);
nor U505 (N_505,In_785,In_1572);
nor U506 (N_506,In_1145,In_723);
and U507 (N_507,In_2269,In_390);
and U508 (N_508,In_2865,In_1164);
nand U509 (N_509,In_1405,In_209);
nand U510 (N_510,In_250,In_1773);
or U511 (N_511,In_99,In_2599);
or U512 (N_512,In_882,In_1);
nor U513 (N_513,In_864,In_6);
xnor U514 (N_514,In_890,In_48);
or U515 (N_515,In_767,In_965);
and U516 (N_516,In_1238,In_1088);
nand U517 (N_517,In_2456,In_1729);
nor U518 (N_518,In_1752,In_683);
or U519 (N_519,In_616,In_366);
or U520 (N_520,In_1011,In_1749);
nor U521 (N_521,In_2027,In_408);
and U522 (N_522,In_54,In_1546);
and U523 (N_523,In_2109,In_2121);
and U524 (N_524,In_539,In_938);
nand U525 (N_525,In_2328,In_2068);
nor U526 (N_526,In_1943,In_1830);
or U527 (N_527,In_522,In_146);
xnor U528 (N_528,In_487,In_1261);
xor U529 (N_529,In_1994,In_202);
nand U530 (N_530,In_2482,In_2909);
nor U531 (N_531,In_2010,In_218);
and U532 (N_532,In_1649,In_1717);
nand U533 (N_533,In_2085,In_871);
nand U534 (N_534,In_1691,In_2532);
and U535 (N_535,In_2276,In_1495);
nand U536 (N_536,In_2169,In_1784);
nor U537 (N_537,In_2547,In_217);
nand U538 (N_538,In_1688,In_1276);
nor U539 (N_539,In_1077,In_2372);
nand U540 (N_540,In_1792,In_160);
and U541 (N_541,In_1258,In_1414);
nand U542 (N_542,In_1540,In_2633);
nor U543 (N_543,In_581,In_2468);
and U544 (N_544,In_382,In_1408);
or U545 (N_545,In_1778,In_2620);
and U546 (N_546,In_1832,In_1031);
nand U547 (N_547,In_206,In_2649);
nand U548 (N_548,In_276,In_240);
or U549 (N_549,In_173,In_283);
nand U550 (N_550,In_523,In_521);
and U551 (N_551,In_1001,In_257);
nor U552 (N_552,In_1180,In_1842);
and U553 (N_553,In_1885,In_2265);
xnor U554 (N_554,In_2093,In_819);
and U555 (N_555,In_2183,In_823);
xor U556 (N_556,In_1179,In_1911);
or U557 (N_557,In_2522,In_2880);
nor U558 (N_558,In_1160,In_77);
xnor U559 (N_559,In_1090,In_811);
nand U560 (N_560,In_687,In_1735);
nor U561 (N_561,In_143,In_1938);
and U562 (N_562,In_248,In_1277);
or U563 (N_563,In_2223,In_1818);
xor U564 (N_564,In_1865,In_2795);
and U565 (N_565,In_1165,In_2458);
nand U566 (N_566,In_2695,In_29);
and U567 (N_567,In_1843,In_648);
nor U568 (N_568,In_2615,In_2247);
nand U569 (N_569,In_596,In_269);
and U570 (N_570,In_949,In_1883);
nor U571 (N_571,In_1361,In_1993);
or U572 (N_572,In_270,In_1591);
or U573 (N_573,In_1125,In_100);
or U574 (N_574,In_1402,In_2901);
and U575 (N_575,In_1466,In_2272);
xnor U576 (N_576,In_2070,In_435);
or U577 (N_577,In_694,In_2687);
or U578 (N_578,In_1437,In_1490);
nand U579 (N_579,In_995,In_2780);
nor U580 (N_580,In_2888,In_1599);
nor U581 (N_581,In_555,In_2063);
and U582 (N_582,In_800,In_1101);
xnor U583 (N_583,In_698,In_1220);
or U584 (N_584,In_374,In_483);
and U585 (N_585,In_601,In_2051);
nor U586 (N_586,In_2981,In_866);
xor U587 (N_587,In_2864,In_2385);
or U588 (N_588,In_2539,In_243);
or U589 (N_589,In_225,In_2053);
or U590 (N_590,In_2783,In_1841);
and U591 (N_591,In_287,In_1284);
or U592 (N_592,In_1632,In_1799);
and U593 (N_593,In_590,In_2232);
or U594 (N_594,In_444,In_1453);
or U595 (N_595,In_20,In_2758);
nand U596 (N_596,In_1215,In_1002);
nor U597 (N_597,In_482,In_334);
nor U598 (N_598,In_895,In_364);
xnor U599 (N_599,In_2958,In_2867);
nand U600 (N_600,In_1615,In_1471);
nand U601 (N_601,In_1153,In_629);
xor U602 (N_602,In_1263,In_2870);
or U603 (N_603,In_1278,In_1218);
nand U604 (N_604,In_2679,In_207);
nor U605 (N_605,In_635,In_2440);
nand U606 (N_606,In_2881,In_2015);
or U607 (N_607,In_308,In_1431);
nor U608 (N_608,In_2568,In_1159);
nand U609 (N_609,In_1403,In_1352);
xor U610 (N_610,In_1182,In_1129);
nor U611 (N_611,In_2313,In_1294);
and U612 (N_612,In_1998,In_233);
and U613 (N_613,In_1320,In_227);
or U614 (N_614,In_708,In_1132);
nand U615 (N_615,In_445,In_1112);
and U616 (N_616,In_1023,In_822);
nand U617 (N_617,In_945,In_354);
xnor U618 (N_618,In_2741,In_1109);
xnor U619 (N_619,In_1695,In_2348);
or U620 (N_620,In_1020,In_1398);
or U621 (N_621,In_244,In_2652);
or U622 (N_622,In_1486,In_2842);
or U623 (N_623,In_2995,In_1962);
and U624 (N_624,In_338,In_2573);
or U625 (N_625,In_1390,In_481);
xor U626 (N_626,In_1586,In_541);
and U627 (N_627,In_2033,In_2329);
or U628 (N_628,In_2081,In_2672);
and U629 (N_629,In_710,In_1945);
nand U630 (N_630,In_397,In_897);
and U631 (N_631,In_242,In_123);
and U632 (N_632,In_343,In_2769);
or U633 (N_633,In_1457,In_2820);
nand U634 (N_634,In_1929,In_2715);
xor U635 (N_635,In_2147,In_296);
and U636 (N_636,In_2238,In_1934);
and U637 (N_637,In_1614,In_1897);
and U638 (N_638,In_1206,In_272);
nor U639 (N_639,In_2705,In_1731);
or U640 (N_640,In_414,In_2794);
and U641 (N_641,In_1474,In_969);
nand U642 (N_642,In_1035,In_310);
and U643 (N_643,In_1530,In_0);
and U644 (N_644,In_2159,In_1721);
nor U645 (N_645,In_849,In_2502);
and U646 (N_646,In_1896,In_1019);
nor U647 (N_647,In_1240,In_2837);
nor U648 (N_648,In_1569,In_730);
and U649 (N_649,In_1927,In_464);
nand U650 (N_650,In_2646,In_2305);
nor U651 (N_651,In_1666,In_2310);
xnor U652 (N_652,In_400,In_1274);
nor U653 (N_653,In_2816,In_2799);
and U654 (N_654,In_430,In_2819);
nand U655 (N_655,In_1200,In_2848);
nand U656 (N_656,In_1803,In_658);
and U657 (N_657,In_1242,In_2364);
xor U658 (N_658,In_46,In_309);
nor U659 (N_659,In_1275,In_317);
and U660 (N_660,In_2688,In_1024);
nand U661 (N_661,In_1635,In_466);
or U662 (N_662,In_298,In_2016);
or U663 (N_663,In_1235,In_657);
nor U664 (N_664,In_2071,In_924);
or U665 (N_665,In_1484,In_1871);
nor U666 (N_666,In_85,In_944);
nor U667 (N_667,In_1631,In_2571);
and U668 (N_668,In_1056,In_1360);
nand U669 (N_669,In_2240,In_1859);
nand U670 (N_670,In_2704,In_1824);
xor U671 (N_671,In_2409,In_2605);
nand U672 (N_672,In_2993,In_2829);
nand U673 (N_673,In_1566,In_574);
or U674 (N_674,In_1149,In_2366);
nand U675 (N_675,In_247,In_2321);
nor U676 (N_676,In_1819,In_1711);
nand U677 (N_677,In_2340,In_1739);
nor U678 (N_678,In_1693,In_1682);
nor U679 (N_679,In_1611,In_2427);
nor U680 (N_680,In_2742,In_1668);
or U681 (N_681,In_383,In_260);
and U682 (N_682,In_1706,In_2642);
nand U683 (N_683,In_1607,In_2575);
or U684 (N_684,In_2965,In_1890);
or U685 (N_685,In_1039,In_87);
or U686 (N_686,In_2537,In_281);
or U687 (N_687,In_1378,In_1782);
or U688 (N_688,In_955,In_2606);
or U689 (N_689,In_1679,In_405);
xor U690 (N_690,In_347,In_2771);
or U691 (N_691,In_1810,In_1137);
and U692 (N_692,In_2299,In_2943);
nand U693 (N_693,In_2044,In_2967);
or U694 (N_694,In_1699,In_2450);
nand U695 (N_695,In_2358,In_901);
and U696 (N_696,In_1768,In_295);
and U697 (N_697,In_2097,In_1887);
or U698 (N_698,In_765,In_291);
and U699 (N_699,In_1262,In_2603);
nor U700 (N_700,In_2499,In_751);
nor U701 (N_701,In_191,In_2034);
nand U702 (N_702,In_2469,In_200);
nor U703 (N_703,In_203,In_1971);
or U704 (N_704,In_2006,In_638);
or U705 (N_705,In_998,In_2952);
xor U706 (N_706,In_2543,In_636);
nand U707 (N_707,In_2527,In_107);
and U708 (N_708,In_74,In_1860);
nor U709 (N_709,In_1393,In_728);
and U710 (N_710,In_426,In_2647);
and U711 (N_711,In_1671,In_2428);
nand U712 (N_712,In_654,In_845);
and U713 (N_713,In_1207,In_2721);
nand U714 (N_714,In_2923,In_2738);
and U715 (N_715,In_867,In_1191);
nand U716 (N_716,In_1760,In_174);
xor U717 (N_717,In_1289,In_2634);
and U718 (N_718,In_975,In_2838);
and U719 (N_719,In_1079,In_2193);
and U720 (N_720,In_2777,In_325);
and U721 (N_721,In_1121,In_47);
or U722 (N_722,In_1924,In_1554);
nand U723 (N_723,In_1777,In_667);
or U724 (N_724,In_2612,In_2743);
and U725 (N_725,In_1447,In_621);
nor U726 (N_726,In_2074,In_2866);
xnor U727 (N_727,In_1186,In_2749);
nor U728 (N_728,In_2317,In_1008);
nor U729 (N_729,In_806,In_288);
and U730 (N_730,In_1374,In_837);
nor U731 (N_731,In_1761,In_2414);
or U732 (N_732,In_2149,In_2435);
and U733 (N_733,In_884,In_1551);
nor U734 (N_734,In_798,In_1014);
and U735 (N_735,In_280,In_416);
nand U736 (N_736,In_2,In_1150);
nand U737 (N_737,In_2514,In_1709);
nor U738 (N_738,In_644,In_1448);
xnor U739 (N_739,In_1060,In_954);
nor U740 (N_740,In_478,In_2912);
nor U741 (N_741,In_1295,In_1583);
or U742 (N_742,In_1340,In_266);
nand U743 (N_743,In_91,In_1791);
nor U744 (N_744,In_360,In_1523);
nor U745 (N_745,In_1283,In_2455);
nor U746 (N_746,In_1226,In_566);
and U747 (N_747,In_1272,In_1139);
nor U748 (N_748,In_2760,In_2137);
xor U749 (N_749,In_614,In_516);
nor U750 (N_750,In_142,In_1196);
nand U751 (N_751,In_2655,In_153);
nor U752 (N_752,In_2818,In_1553);
and U753 (N_753,In_2073,In_479);
and U754 (N_754,In_673,In_81);
and U755 (N_755,In_1728,In_1166);
and U756 (N_756,In_1185,In_1487);
or U757 (N_757,In_741,In_1260);
or U758 (N_758,In_2141,In_2508);
nor U759 (N_759,In_2082,In_2882);
nand U760 (N_760,In_1584,In_1399);
or U761 (N_761,In_212,In_2290);
nor U762 (N_762,In_2878,In_2257);
and U763 (N_763,In_2989,In_2237);
nor U764 (N_764,In_744,In_1610);
or U765 (N_765,In_2678,In_2383);
and U766 (N_766,In_2391,In_688);
xnor U767 (N_767,In_1740,In_1082);
nor U768 (N_768,In_342,In_2449);
xnor U769 (N_769,In_473,In_1347);
nor U770 (N_770,In_1876,In_2521);
nor U771 (N_771,In_453,In_1868);
and U772 (N_772,In_2822,In_889);
nand U773 (N_773,In_1571,In_1446);
nor U774 (N_774,In_2852,In_2906);
nor U775 (N_775,In_2396,In_136);
nor U776 (N_776,In_976,In_1589);
nand U777 (N_777,In_1086,In_781);
or U778 (N_778,In_570,In_2976);
and U779 (N_779,In_322,In_1643);
xnor U780 (N_780,In_677,In_2875);
nor U781 (N_781,In_510,In_1078);
and U782 (N_782,In_284,In_82);
nand U783 (N_783,In_1458,In_1073);
or U784 (N_784,In_1933,In_1306);
or U785 (N_785,In_624,In_2309);
and U786 (N_786,In_627,In_2052);
and U787 (N_787,In_2182,In_1941);
nand U788 (N_788,In_50,In_1430);
and U789 (N_789,In_2839,In_2446);
xor U790 (N_790,In_2873,In_858);
nor U791 (N_791,In_1071,In_1384);
or U792 (N_792,In_2090,In_2473);
or U793 (N_793,In_11,In_1686);
nor U794 (N_794,In_766,In_386);
nand U795 (N_795,In_376,In_984);
or U796 (N_796,In_362,In_1310);
nand U797 (N_797,In_797,In_369);
nor U798 (N_798,In_1606,In_1061);
and U799 (N_799,In_922,In_2037);
or U800 (N_800,In_1972,In_2697);
nor U801 (N_801,In_874,In_1006);
nand U802 (N_802,In_326,In_771);
nor U803 (N_803,In_2072,In_2036);
and U804 (N_804,In_651,In_2056);
xor U805 (N_805,In_2210,In_2128);
or U806 (N_806,In_559,In_1234);
and U807 (N_807,In_2542,In_1526);
nand U808 (N_808,In_1210,In_2400);
or U809 (N_809,In_1314,In_1989);
nor U810 (N_810,In_345,In_2792);
or U811 (N_811,In_1535,In_918);
and U812 (N_812,In_2094,In_853);
and U813 (N_813,In_1767,In_56);
nor U814 (N_814,In_1652,In_2854);
and U815 (N_815,In_2407,In_2708);
nand U816 (N_816,In_1755,In_1059);
and U817 (N_817,In_2885,In_1963);
nand U818 (N_818,In_817,In_2342);
and U819 (N_819,In_1494,In_1629);
xor U820 (N_820,In_714,In_637);
and U821 (N_821,In_2426,In_40);
nor U822 (N_822,In_396,In_1042);
or U823 (N_823,In_2289,In_1080);
nand U824 (N_824,In_2351,In_2814);
nand U825 (N_825,In_2167,In_2668);
and U826 (N_826,In_2120,In_972);
nor U827 (N_827,In_501,In_1550);
and U828 (N_828,In_653,In_42);
or U829 (N_829,In_1783,In_431);
xor U830 (N_830,In_719,In_2012);
nand U831 (N_831,In_1575,In_1833);
nand U832 (N_832,In_249,In_731);
or U833 (N_833,In_885,In_2825);
nor U834 (N_834,In_2830,In_707);
xor U835 (N_835,In_1475,In_2263);
and U836 (N_836,In_118,In_375);
nor U837 (N_837,In_2301,In_2980);
nand U838 (N_838,In_1397,In_1442);
nor U839 (N_839,In_2355,In_1726);
or U840 (N_840,In_1249,In_826);
and U841 (N_841,In_1241,In_931);
xnor U842 (N_842,In_2485,In_2390);
or U843 (N_843,In_2940,In_1304);
nor U844 (N_844,In_2730,In_1873);
or U845 (N_845,In_1331,In_1054);
nand U846 (N_846,In_2669,In_2049);
xor U847 (N_847,In_2286,In_600);
nor U848 (N_848,In_329,In_1247);
nor U849 (N_849,In_465,In_2985);
nor U850 (N_850,In_655,In_511);
nor U851 (N_851,In_1505,In_2431);
nor U852 (N_852,In_2577,In_2497);
and U853 (N_853,In_835,In_894);
xnor U854 (N_854,In_2856,In_2871);
nand U855 (N_855,In_2627,In_1188);
nand U856 (N_856,In_2388,In_2080);
nand U857 (N_857,In_1886,In_1493);
nor U858 (N_858,In_1084,In_499);
nor U859 (N_859,In_1970,In_970);
xor U860 (N_860,In_2302,In_2318);
or U861 (N_861,In_2624,In_2234);
nand U862 (N_862,In_1318,In_2614);
or U863 (N_863,In_2515,In_764);
or U864 (N_864,In_2202,In_2613);
and U865 (N_865,In_65,In_1595);
xor U866 (N_866,In_1795,In_879);
nor U867 (N_867,In_565,In_2467);
and U868 (N_868,In_1973,In_1727);
nor U869 (N_869,In_2113,In_2040);
nand U870 (N_870,In_1395,In_1656);
nand U871 (N_871,In_2496,In_2576);
and U872 (N_872,In_2356,In_1640);
and U873 (N_873,In_2420,In_1724);
and U874 (N_874,In_877,In_1880);
nor U875 (N_875,In_1951,In_2883);
nand U876 (N_876,In_167,In_147);
xnor U877 (N_877,In_2936,In_2353);
or U878 (N_878,In_1330,In_1045);
or U879 (N_879,In_2926,In_786);
or U880 (N_880,In_229,In_2371);
or U881 (N_881,In_2023,In_2256);
or U882 (N_882,In_679,In_1141);
and U883 (N_883,In_2058,In_2230);
nand U884 (N_884,In_615,In_606);
nand U885 (N_885,In_304,In_138);
nor U886 (N_886,In_93,In_1513);
xnor U887 (N_887,In_1891,In_2860);
and U888 (N_888,In_2123,In_2835);
or U889 (N_889,In_887,In_959);
or U890 (N_890,In_2156,In_2478);
or U891 (N_891,In_1436,In_2110);
or U892 (N_892,In_1743,In_1736);
or U893 (N_893,In_388,In_844);
and U894 (N_894,In_792,In_633);
nand U895 (N_895,In_2465,In_2375);
nand U896 (N_896,In_2984,In_2067);
nand U897 (N_897,In_2218,In_1232);
nor U898 (N_898,In_2046,In_2104);
nand U899 (N_899,In_38,In_2436);
and U900 (N_900,In_1573,In_463);
and U901 (N_901,In_2689,In_1148);
nand U902 (N_902,In_1454,In_179);
nor U903 (N_903,In_612,In_94);
and U904 (N_904,In_2998,In_2205);
nor U905 (N_905,In_859,In_1822);
and U906 (N_906,In_1332,In_2288);
nand U907 (N_907,In_2828,In_2964);
xor U908 (N_908,In_933,In_256);
nor U909 (N_909,In_194,In_2661);
and U910 (N_910,In_1603,In_55);
nand U911 (N_911,In_2847,In_1893);
and U912 (N_912,In_2778,In_22);
nor U913 (N_913,In_2941,In_1555);
and U914 (N_914,In_971,In_1745);
nand U915 (N_915,In_2663,In_1700);
or U916 (N_916,In_1222,In_474);
nor U917 (N_917,In_896,In_2338);
or U918 (N_918,In_387,In_1244);
nor U919 (N_919,In_757,In_1988);
or U920 (N_920,In_1903,In_2657);
nand U921 (N_921,In_2635,In_920);
nand U922 (N_922,In_1676,In_1770);
and U923 (N_923,In_2535,In_45);
nand U924 (N_924,In_2461,In_908);
and U925 (N_925,In_619,In_2786);
and U926 (N_926,In_494,In_1217);
and U927 (N_927,In_1565,In_2626);
and U928 (N_928,In_557,In_49);
and U929 (N_929,In_89,In_449);
or U930 (N_930,In_1429,In_1958);
nor U931 (N_931,In_1093,In_2879);
or U932 (N_932,In_2561,In_358);
or U933 (N_933,In_2782,In_323);
nand U934 (N_934,In_2445,In_2933);
or U935 (N_935,In_300,In_1311);
and U936 (N_936,In_193,In_1212);
xnor U937 (N_937,In_36,In_2680);
nor U938 (N_938,In_117,In_228);
nor U939 (N_939,In_1531,In_299);
or U940 (N_940,In_980,In_631);
nand U941 (N_941,In_1604,In_1194);
nor U942 (N_942,In_1327,In_349);
and U943 (N_943,In_2127,In_1044);
or U944 (N_944,In_2800,In_2126);
nor U945 (N_945,In_649,In_2392);
nand U946 (N_946,In_1236,In_780);
nand U947 (N_947,In_1083,In_2441);
nand U948 (N_948,In_665,In_452);
and U949 (N_949,In_1480,In_1245);
nor U950 (N_950,In_155,In_598);
nor U951 (N_951,In_1805,In_2916);
xor U952 (N_952,In_2148,In_1392);
xnor U953 (N_953,In_2639,In_2992);
and U954 (N_954,In_43,In_415);
nand U955 (N_955,In_2832,In_32);
and U956 (N_956,In_937,In_990);
nand U957 (N_957,In_796,In_2020);
nor U958 (N_958,In_2330,In_2368);
nand U959 (N_959,In_1280,In_2994);
or U960 (N_960,In_2924,In_2278);
xnor U961 (N_961,In_2564,In_1638);
nand U962 (N_962,In_1877,In_1155);
nand U963 (N_963,In_2949,In_824);
nand U964 (N_964,In_62,In_1339);
nand U965 (N_965,In_1209,In_2549);
xnor U966 (N_966,In_2625,In_1135);
nand U967 (N_967,In_1662,In_1713);
xor U968 (N_968,In_791,In_2982);
or U969 (N_969,In_732,In_215);
and U970 (N_970,In_930,In_929);
nand U971 (N_971,In_927,In_2805);
and U972 (N_972,In_666,In_201);
nor U973 (N_973,In_1230,In_2405);
and U974 (N_974,In_1070,In_496);
nor U975 (N_975,In_83,In_318);
nand U976 (N_976,In_1010,In_2312);
and U977 (N_977,In_549,In_2619);
nor U978 (N_978,In_3,In_981);
or U979 (N_979,In_1291,In_2197);
or U980 (N_980,In_1771,In_18);
nand U981 (N_981,In_758,In_2242);
or U982 (N_982,In_2581,In_216);
nor U983 (N_983,In_122,In_116);
xor U984 (N_984,In_1203,In_1463);
xor U985 (N_985,In_1134,In_2788);
nor U986 (N_986,In_2011,In_2415);
or U987 (N_987,In_2731,In_1198);
nand U988 (N_988,In_1853,In_1097);
and U989 (N_989,In_2511,In_1817);
nand U990 (N_990,In_802,In_2430);
or U991 (N_991,In_1492,In_1204);
and U992 (N_992,In_1064,In_577);
or U993 (N_993,In_2107,In_446);
nor U994 (N_994,In_2546,In_851);
nand U995 (N_995,In_1172,In_2823);
xnor U996 (N_996,In_2815,In_1512);
nor U997 (N_997,In_1556,In_1460);
nor U998 (N_998,In_2969,In_2483);
and U999 (N_999,In_900,In_1169);
nand U1000 (N_1000,In_1650,In_2632);
nand U1001 (N_1001,In_236,In_2102);
or U1002 (N_1002,In_1909,In_534);
or U1003 (N_1003,In_2324,In_660);
or U1004 (N_1004,In_893,In_1992);
or U1005 (N_1005,In_2729,In_2443);
xor U1006 (N_1006,In_1984,In_171);
and U1007 (N_1007,In_1636,In_561);
nor U1008 (N_1008,In_2350,In_13);
nor U1009 (N_1009,In_106,In_983);
nor U1010 (N_1010,In_720,In_529);
and U1011 (N_1011,In_1156,In_2790);
and U1012 (N_1012,In_1298,In_2585);
or U1013 (N_1013,In_2424,In_2349);
and U1014 (N_1014,In_2955,In_1507);
nand U1015 (N_1015,In_2323,In_166);
nand U1016 (N_1016,In_1953,In_2554);
and U1017 (N_1017,In_1367,In_923);
nand U1018 (N_1018,In_1986,In_353);
xnor U1019 (N_1019,In_443,In_26);
and U1020 (N_1020,In_2211,In_1052);
and U1021 (N_1021,In_1286,In_1433);
or U1022 (N_1022,In_41,In_2644);
xnor U1023 (N_1023,In_1634,In_1815);
and U1024 (N_1024,In_1074,In_2195);
and U1025 (N_1025,In_285,In_772);
or U1026 (N_1026,In_404,In_2664);
or U1027 (N_1027,In_2559,In_1040);
or U1028 (N_1028,In_2740,In_1627);
nor U1029 (N_1029,In_2701,In_702);
and U1030 (N_1030,In_2935,In_1707);
or U1031 (N_1031,In_2775,In_527);
xnor U1032 (N_1032,In_139,In_2448);
and U1033 (N_1033,In_1394,In_1181);
nor U1034 (N_1034,In_2055,In_1254);
or U1035 (N_1035,In_1637,In_90);
nand U1036 (N_1036,In_2770,In_2493);
nand U1037 (N_1037,In_379,In_2970);
nor U1038 (N_1038,In_1115,In_2352);
nor U1039 (N_1039,In_1094,In_942);
or U1040 (N_1040,In_2567,In_2919);
xor U1041 (N_1041,In_573,In_1710);
nand U1042 (N_1042,In_1114,In_1501);
or U1043 (N_1043,In_986,In_2589);
and U1044 (N_1044,In_2035,In_2185);
and U1045 (N_1045,In_344,In_2031);
and U1046 (N_1046,In_613,In_1672);
or U1047 (N_1047,In_2737,In_2184);
nor U1048 (N_1048,In_314,In_2279);
nor U1049 (N_1049,In_1483,In_1370);
nand U1050 (N_1050,In_2732,In_721);
nand U1051 (N_1051,In_2130,In_2451);
and U1052 (N_1052,In_1987,In_2610);
nand U1053 (N_1053,In_1533,In_1144);
or U1054 (N_1054,In_1660,In_537);
or U1055 (N_1055,In_2929,In_1582);
xor U1056 (N_1056,In_711,In_2911);
and U1057 (N_1057,In_2764,In_815);
and U1058 (N_1058,In_163,In_746);
or U1059 (N_1059,In_1353,In_2327);
nand U1060 (N_1060,In_2101,In_936);
or U1061 (N_1061,In_96,In_108);
nor U1062 (N_1062,In_1580,In_2505);
nand U1063 (N_1063,In_2676,In_2194);
and U1064 (N_1064,In_2972,In_254);
or U1065 (N_1065,In_2950,In_1995);
nor U1066 (N_1066,In_467,In_1955);
xnor U1067 (N_1067,In_1593,In_2534);
nand U1068 (N_1068,In_528,In_2406);
nor U1069 (N_1069,In_211,In_1246);
nand U1070 (N_1070,In_695,In_912);
or U1071 (N_1071,In_2720,In_2060);
or U1072 (N_1072,In_1063,In_187);
xnor U1073 (N_1073,In_419,In_462);
and U1074 (N_1074,In_1920,In_490);
or U1075 (N_1075,In_2510,In_1326);
or U1076 (N_1076,In_1539,In_2628);
xnor U1077 (N_1077,In_2548,In_548);
nor U1078 (N_1078,In_2297,In_2600);
and U1079 (N_1079,In_2188,In_159);
nor U1080 (N_1080,In_1095,In_292);
and U1081 (N_1081,In_1959,In_675);
or U1082 (N_1082,In_1363,In_60);
or U1083 (N_1083,In_2947,In_1459);
or U1084 (N_1084,In_2863,In_2114);
or U1085 (N_1085,In_2703,In_175);
nand U1086 (N_1086,In_999,In_1322);
nor U1087 (N_1087,In_64,In_148);
nor U1088 (N_1088,In_2670,In_2365);
or U1089 (N_1089,In_2395,In_373);
nor U1090 (N_1090,In_1659,In_2908);
and U1091 (N_1091,In_2748,In_2032);
nand U1092 (N_1092,In_671,In_2754);
nand U1093 (N_1093,In_1359,In_1264);
nor U1094 (N_1094,In_2198,In_2850);
nand U1095 (N_1095,In_2591,In_1450);
and U1096 (N_1096,In_156,In_943);
nand U1097 (N_1097,In_1107,In_2442);
nand U1098 (N_1098,In_948,In_2718);
nand U1099 (N_1099,In_1328,In_599);
nor U1100 (N_1100,In_2334,In_1468);
nor U1101 (N_1101,In_328,In_471);
nor U1102 (N_1102,In_1663,In_1104);
or U1103 (N_1103,In_1511,In_1489);
or U1104 (N_1104,In_742,In_1950);
nor U1105 (N_1105,In_968,In_2962);
xor U1106 (N_1106,In_1762,In_1525);
xor U1107 (N_1107,In_451,In_749);
and U1108 (N_1108,In_1522,In_760);
or U1109 (N_1109,In_2207,In_2887);
and U1110 (N_1110,In_2656,In_162);
nor U1111 (N_1111,In_1769,In_1400);
nand U1112 (N_1112,In_459,In_1655);
and U1113 (N_1113,In_372,In_855);
nand U1114 (N_1114,In_1116,In_2997);
nor U1115 (N_1115,In_2990,In_2066);
or U1116 (N_1116,In_271,In_1515);
or U1117 (N_1117,In_1633,In_609);
nand U1118 (N_1118,In_1790,In_2913);
xnor U1119 (N_1119,In_989,In_848);
nand U1120 (N_1120,In_2594,In_2590);
nand U1121 (N_1121,In_1848,In_1548);
xor U1122 (N_1122,In_27,In_2736);
and U1123 (N_1123,In_674,In_2892);
nor U1124 (N_1124,In_1789,In_2507);
nor U1125 (N_1125,In_255,In_316);
nand U1126 (N_1126,In_2429,In_643);
or U1127 (N_1127,In_2580,In_16);
or U1128 (N_1128,In_2915,In_1157);
or U1129 (N_1129,In_1834,In_134);
xnor U1130 (N_1130,In_1380,In_2834);
xnor U1131 (N_1131,In_1854,In_432);
xnor U1132 (N_1132,In_128,In_327);
and U1133 (N_1133,In_1355,In_1138);
and U1134 (N_1134,In_846,In_409);
nand U1135 (N_1135,In_1590,In_571);
and U1136 (N_1136,In_2164,In_1026);
nor U1137 (N_1137,In_1609,In_1354);
nor U1138 (N_1138,In_297,In_1684);
or U1139 (N_1139,In_2787,In_1449);
and U1140 (N_1140,In_560,In_2710);
nor U1141 (N_1141,In_762,In_909);
or U1142 (N_1142,In_1915,In_2213);
xor U1143 (N_1143,In_2889,In_196);
or U1144 (N_1144,In_2766,In_1844);
or U1145 (N_1145,In_1786,In_2877);
nor U1146 (N_1146,In_2572,In_830);
nand U1147 (N_1147,In_1608,In_423);
nand U1148 (N_1148,In_705,In_1542);
nor U1149 (N_1149,In_2569,In_2895);
and U1150 (N_1150,In_2813,In_282);
nand U1151 (N_1151,In_401,In_2008);
or U1152 (N_1152,In_1944,In_1434);
nand U1153 (N_1153,In_1170,In_1857);
or U1154 (N_1154,In_1562,In_1597);
and U1155 (N_1155,In_1524,In_1482);
or U1156 (N_1156,In_192,In_881);
nor U1157 (N_1157,In_1451,In_646);
or U1158 (N_1158,In_1935,In_2810);
nor U1159 (N_1159,In_2836,In_1623);
and U1160 (N_1160,In_2587,In_1979);
or U1161 (N_1161,In_2667,In_1142);
or U1162 (N_1162,In_696,In_1301);
nand U1163 (N_1163,In_538,In_663);
nor U1164 (N_1164,In_2869,In_966);
and U1165 (N_1165,In_1177,In_2359);
nor U1166 (N_1166,In_289,In_176);
xnor U1167 (N_1167,In_868,In_1377);
nor U1168 (N_1168,In_1901,In_92);
and U1169 (N_1169,In_1780,In_2796);
and U1170 (N_1170,In_2384,In_2386);
nor U1171 (N_1171,In_779,In_152);
and U1172 (N_1172,In_71,In_413);
nor U1173 (N_1173,In_997,In_2974);
nor U1174 (N_1174,In_12,In_2398);
or U1175 (N_1175,In_2345,In_2831);
nor U1176 (N_1176,In_169,In_2389);
and U1177 (N_1177,In_2650,In_2444);
and U1178 (N_1178,In_2690,In_1835);
and U1179 (N_1179,In_2495,In_1895);
or U1180 (N_1180,In_1161,In_1424);
nor U1181 (N_1181,In_1532,In_691);
nand U1182 (N_1182,In_1516,In_967);
or U1183 (N_1183,In_1990,In_2347);
or U1184 (N_1184,In_2622,In_2726);
or U1185 (N_1185,In_1796,In_312);
nor U1186 (N_1186,In_2387,In_2717);
nand U1187 (N_1187,In_1802,In_1746);
nor U1188 (N_1188,In_1136,In_2757);
xnor U1189 (N_1189,In_1391,In_2492);
nor U1190 (N_1190,In_2724,In_2191);
nand U1191 (N_1191,In_1333,In_438);
or U1192 (N_1192,In_1461,In_2271);
nand U1193 (N_1193,In_2103,In_977);
nand U1194 (N_1194,In_625,In_2224);
nor U1195 (N_1195,In_339,In_2596);
nor U1196 (N_1196,In_1779,In_2057);
nor U1197 (N_1197,In_57,In_891);
nand U1198 (N_1198,In_1619,In_348);
nor U1199 (N_1199,In_2145,In_161);
and U1200 (N_1200,In_1601,In_1012);
nor U1201 (N_1201,In_1048,In_1146);
and U1202 (N_1202,In_1214,In_2045);
nand U1203 (N_1203,In_460,In_1324);
nand U1204 (N_1204,In_1620,In_1208);
and U1205 (N_1205,In_9,In_1922);
nor U1206 (N_1206,In_2274,In_2939);
and U1207 (N_1207,In_1265,In_911);
and U1208 (N_1208,In_181,In_1346);
xor U1209 (N_1209,In_1738,In_2486);
and U1210 (N_1210,In_532,In_678);
and U1211 (N_1211,In_2725,In_1730);
xnor U1212 (N_1212,In_2014,In_992);
and U1213 (N_1213,In_2048,In_1557);
or U1214 (N_1214,In_2574,In_2857);
nor U1215 (N_1215,In_219,In_1348);
xor U1216 (N_1216,In_1823,In_941);
and U1217 (N_1217,In_68,In_23);
and U1218 (N_1218,In_368,In_1441);
or U1219 (N_1219,In_1051,In_558);
nor U1220 (N_1220,In_406,In_365);
xor U1221 (N_1221,In_2954,In_1624);
nand U1222 (N_1222,In_1081,In_520);
nand U1223 (N_1223,In_1030,In_1382);
nand U1224 (N_1224,In_526,In_164);
nand U1225 (N_1225,In_630,In_1287);
nor U1226 (N_1226,In_778,In_2648);
or U1227 (N_1227,In_450,In_810);
nor U1228 (N_1228,In_1445,In_1605);
or U1229 (N_1229,In_2260,In_2791);
and U1230 (N_1230,In_410,In_919);
nor U1231 (N_1231,In_2696,In_2674);
nand U1232 (N_1232,In_2030,In_2277);
nor U1233 (N_1233,In_1594,In_1163);
nor U1234 (N_1234,In_1518,In_307);
and U1235 (N_1235,In_1096,In_700);
and U1236 (N_1236,In_1881,In_2682);
and U1237 (N_1237,In_2311,In_1867);
nand U1238 (N_1238,In_1837,In_2938);
xnor U1239 (N_1239,In_2000,In_2942);
or U1240 (N_1240,In_2529,In_661);
nor U1241 (N_1241,In_514,In_1357);
xor U1242 (N_1242,In_1110,In_1913);
or U1243 (N_1243,In_1966,In_552);
and U1244 (N_1244,In_2896,In_850);
and U1245 (N_1245,In_180,In_486);
xnor U1246 (N_1246,In_1472,In_2062);
nor U1247 (N_1247,In_2840,In_761);
or U1248 (N_1248,In_2416,In_628);
or U1249 (N_1249,In_1317,In_1675);
nand U1250 (N_1250,In_2125,In_24);
and U1251 (N_1251,In_1119,In_111);
or U1252 (N_1252,In_2190,In_2971);
or U1253 (N_1253,In_656,In_1253);
nand U1254 (N_1254,In_204,In_697);
or U1255 (N_1255,In_381,In_736);
nand U1256 (N_1256,In_1428,In_2402);
and U1257 (N_1257,In_208,In_112);
nor U1258 (N_1258,In_642,In_1980);
xnor U1259 (N_1259,In_2204,In_37);
and U1260 (N_1260,In_1732,In_2370);
xor U1261 (N_1261,In_952,In_393);
and U1262 (N_1262,In_188,In_789);
and U1263 (N_1263,In_2920,In_2463);
or U1264 (N_1264,In_98,In_2618);
xor U1265 (N_1265,In_2001,In_745);
xnor U1266 (N_1266,In_1793,In_1549);
and U1267 (N_1267,In_2886,In_2179);
xor U1268 (N_1268,In_2013,In_1563);
or U1269 (N_1269,In_1288,In_2135);
and U1270 (N_1270,In_1579,In_267);
nand U1271 (N_1271,In_220,In_1690);
nand U1272 (N_1272,In_725,In_1016);
nand U1273 (N_1273,In_507,In_2039);
and U1274 (N_1274,In_1091,In_2653);
xnor U1275 (N_1275,In_504,In_2199);
nor U1276 (N_1276,In_2702,In_398);
and U1277 (N_1277,In_357,In_2686);
or U1278 (N_1278,In_2162,In_367);
nor U1279 (N_1279,In_1753,In_2418);
and U1280 (N_1280,In_575,In_1696);
or U1281 (N_1281,In_1385,In_1251);
and U1282 (N_1282,In_1712,In_833);
xor U1283 (N_1283,In_1644,In_199);
xor U1284 (N_1284,In_2078,In_442);
or U1285 (N_1285,In_1443,In_2092);
nor U1286 (N_1286,In_2512,In_1369);
nor U1287 (N_1287,In_2381,In_420);
and U1288 (N_1288,In_640,In_2811);
or U1289 (N_1289,In_1055,In_137);
and U1290 (N_1290,In_2122,In_1167);
and U1291 (N_1291,In_1928,In_2076);
and U1292 (N_1292,In_2022,In_1616);
and U1293 (N_1293,In_2983,In_1654);
nor U1294 (N_1294,In_2106,In_1421);
nor U1295 (N_1295,In_793,In_1538);
or U1296 (N_1296,In_2453,In_500);
nand U1297 (N_1297,In_979,In_1467);
nand U1298 (N_1298,In_2041,In_63);
or U1299 (N_1299,In_394,In_1558);
nand U1300 (N_1300,In_44,In_1757);
and U1301 (N_1301,In_1307,In_2801);
or U1302 (N_1302,In_2021,In_2410);
or U1303 (N_1303,In_618,In_1747);
xnor U1304 (N_1304,In_1365,In_1742);
or U1305 (N_1305,In_2216,In_476);
nand U1306 (N_1306,In_1034,In_517);
nor U1307 (N_1307,In_645,In_2630);
and U1308 (N_1308,In_690,In_2607);
and U1309 (N_1309,In_2583,In_2773);
and U1310 (N_1310,In_2579,In_1195);
nor U1311 (N_1311,In_395,In_1544);
or U1312 (N_1312,In_2069,In_2098);
nand U1313 (N_1313,In_2963,In_340);
nand U1314 (N_1314,In_814,In_805);
nand U1315 (N_1315,In_1673,In_1192);
xor U1316 (N_1316,In_1923,In_2957);
or U1317 (N_1317,In_2189,In_2776);
nor U1318 (N_1318,In_2752,In_1578);
nand U1319 (N_1319,In_567,In_1162);
or U1320 (N_1320,In_1954,In_346);
and U1321 (N_1321,In_2054,In_1942);
nand U1322 (N_1322,In_1229,In_551);
and U1323 (N_1323,In_2470,In_1714);
and U1324 (N_1324,In_359,In_2462);
and U1325 (N_1325,In_418,In_1481);
xor U1326 (N_1326,In_2595,In_1961);
or U1327 (N_1327,In_870,In_585);
nand U1328 (N_1328,In_1598,In_2172);
and U1329 (N_1329,In_2206,In_985);
nor U1330 (N_1330,In_356,In_2261);
nor U1331 (N_1331,In_1981,In_1187);
and U1332 (N_1332,In_782,In_1389);
and U1333 (N_1333,In_197,In_594);
nor U1334 (N_1334,In_1350,In_2487);
nand U1335 (N_1335,In_1427,In_2161);
nor U1336 (N_1336,In_536,In_392);
xnor U1337 (N_1337,In_2960,In_2201);
nor U1338 (N_1338,In_1176,In_59);
nor U1339 (N_1339,In_2217,In_1068);
xnor U1340 (N_1340,In_417,In_2140);
and U1341 (N_1341,In_80,In_1806);
nor U1342 (N_1342,In_1387,In_617);
nand U1343 (N_1343,In_1047,In_768);
or U1344 (N_1344,In_2544,In_1388);
nand U1345 (N_1345,In_407,In_1342);
and U1346 (N_1346,In_2671,In_184);
and U1347 (N_1347,In_753,In_33);
nor U1348 (N_1348,In_1677,In_210);
nand U1349 (N_1349,In_424,In_2930);
xnor U1350 (N_1350,In_2551,In_2662);
nor U1351 (N_1351,In_1343,In_2807);
or U1352 (N_1352,In_813,In_2315);
or U1353 (N_1353,In_1362,In_1947);
xnor U1354 (N_1354,In_2804,In_1089);
or U1355 (N_1355,In_2422,In_1869);
and U1356 (N_1356,In_1018,In_1478);
and U1357 (N_1357,In_740,In_1807);
and U1358 (N_1358,In_905,In_458);
nor U1359 (N_1359,In_670,In_461);
xnor U1360 (N_1360,In_1356,In_403);
and U1361 (N_1361,In_1718,In_2408);
nand U1362 (N_1362,In_35,In_2975);
and U1363 (N_1363,In_512,In_962);
and U1364 (N_1364,In_1456,In_634);
or U1365 (N_1365,In_1716,In_1508);
nand U1366 (N_1366,In_2306,In_1653);
nand U1367 (N_1367,In_2259,In_1349);
nor U1368 (N_1368,In_899,In_2333);
and U1369 (N_1369,In_480,In_1072);
nand U1370 (N_1370,In_1587,In_904);
nor U1371 (N_1371,In_1651,In_2611);
xor U1372 (N_1372,In_274,In_1702);
nand U1373 (N_1373,In_1376,In_530);
nand U1374 (N_1374,In_1303,In_1488);
xnor U1375 (N_1375,In_2931,In_2124);
and U1376 (N_1376,In_2609,In_2812);
nand U1377 (N_1377,In_2973,In_2910);
xnor U1378 (N_1378,In_133,In_441);
and U1379 (N_1379,In_1199,In_841);
nand U1380 (N_1380,In_2111,In_724);
nand U1381 (N_1381,In_1665,In_1630);
nand U1382 (N_1382,In_934,In_1814);
or U1383 (N_1383,In_2362,In_763);
nor U1384 (N_1384,In_2419,In_2490);
or U1385 (N_1385,In_144,In_650);
and U1386 (N_1386,In_1302,In_1722);
nand U1387 (N_1387,In_1057,In_639);
xnor U1388 (N_1388,In_1375,In_1292);
xor U1389 (N_1389,In_1541,In_1473);
nor U1390 (N_1390,In_1025,In_1836);
or U1391 (N_1391,In_234,In_1123);
and U1392 (N_1392,In_226,In_807);
nor U1393 (N_1393,In_2774,In_2753);
and U1394 (N_1394,In_1838,In_5);
and U1395 (N_1395,In_1130,In_2173);
and U1396 (N_1396,In_1863,In_140);
nand U1397 (N_1397,In_2254,In_1858);
and U1398 (N_1398,In_2212,In_7);
and U1399 (N_1399,In_2394,In_2637);
nand U1400 (N_1400,In_1894,In_1855);
or U1401 (N_1401,In_875,In_434);
nor U1402 (N_1402,In_245,In_715);
nor U1403 (N_1403,In_2154,In_251);
nor U1404 (N_1404,In_2900,In_439);
nor U1405 (N_1405,In_2028,In_130);
nor U1406 (N_1406,In_576,In_385);
and U1407 (N_1407,In_2641,In_544);
and U1408 (N_1408,In_2827,In_2479);
nand U1409 (N_1409,In_2268,In_2180);
or U1410 (N_1410,In_1190,In_2961);
xor U1411 (N_1411,In_428,In_2088);
or U1412 (N_1412,In_1936,In_2560);
nor U1413 (N_1413,In_391,In_808);
or U1414 (N_1414,In_2789,In_1158);
and U1415 (N_1415,In_2654,In_839);
and U1416 (N_1416,In_2927,In_2155);
xor U1417 (N_1417,In_1205,In_2808);
nor U1418 (N_1418,In_564,In_2275);
and U1419 (N_1419,In_737,In_2506);
or U1420 (N_1420,In_2477,In_1849);
nor U1421 (N_1421,In_1825,In_422);
xnor U1422 (N_1422,In_1065,In_84);
or U1423 (N_1423,In_2116,In_957);
nor U1424 (N_1424,In_2681,In_263);
and U1425 (N_1425,In_21,In_2171);
nor U1426 (N_1426,In_95,In_1092);
and U1427 (N_1427,In_1496,In_2631);
nand U1428 (N_1428,In_604,In_1956);
or U1429 (N_1429,In_73,In_2636);
nand U1430 (N_1430,In_588,In_659);
xor U1431 (N_1431,In_2401,In_214);
and U1432 (N_1432,In_261,In_569);
nor U1433 (N_1433,In_883,In_189);
or U1434 (N_1434,In_2423,In_2570);
xnor U1435 (N_1435,In_1469,In_2809);
xor U1436 (N_1436,In_773,In_1000);
xnor U1437 (N_1437,In_1111,In_1800);
nor U1438 (N_1438,In_246,In_1975);
or U1439 (N_1439,In_603,In_70);
and U1440 (N_1440,In_2397,In_1120);
nand U1441 (N_1441,In_1050,In_2996);
and U1442 (N_1442,In_607,In_2893);
nor U1443 (N_1443,In_1268,In_113);
xnor U1444 (N_1444,In_1899,In_2562);
nor U1445 (N_1445,In_124,In_2797);
nand U1446 (N_1446,In_2245,In_411);
and U1447 (N_1447,In_1698,In_2379);
nor U1448 (N_1448,In_2898,In_1976);
nor U1449 (N_1449,In_1756,In_509);
and U1450 (N_1450,In_2566,In_1351);
nor U1451 (N_1451,In_2399,In_1221);
or U1452 (N_1452,In_1259,In_1344);
and U1453 (N_1453,In_1879,In_268);
nand U1454 (N_1454,In_2043,In_436);
nand U1455 (N_1455,In_861,In_125);
and U1456 (N_1456,In_2890,In_1062);
nor U1457 (N_1457,In_2460,In_1213);
nor U1458 (N_1458,In_1996,In_2284);
nor U1459 (N_1459,In_1664,In_1364);
or U1460 (N_1460,In_2988,In_2798);
and U1461 (N_1461,In_2501,In_1733);
and U1462 (N_1462,In_15,In_1067);
xnor U1463 (N_1463,In_956,In_1309);
nand U1464 (N_1464,In_2902,In_2763);
nor U1465 (N_1465,In_1766,In_2250);
nand U1466 (N_1466,In_1043,In_535);
or U1467 (N_1467,In_2494,In_1131);
nand U1468 (N_1468,In_1965,In_568);
nor U1469 (N_1469,In_1925,In_1171);
nor U1470 (N_1470,In_2464,In_2745);
and U1471 (N_1471,In_279,In_262);
nor U1472 (N_1472,In_427,In_2932);
nor U1473 (N_1473,In_1681,In_2158);
nor U1474 (N_1474,In_1882,In_2751);
nor U1475 (N_1475,In_421,In_774);
or U1476 (N_1476,In_1826,In_1029);
or U1477 (N_1477,In_1418,In_2645);
nand U1478 (N_1478,In_843,In_1907);
or U1479 (N_1479,In_2874,In_2922);
or U1480 (N_1480,In_1438,In_2255);
and U1481 (N_1481,In_1118,In_17);
nand U1482 (N_1482,In_2956,In_495);
and U1483 (N_1483,In_2714,In_1874);
nand U1484 (N_1484,In_2296,In_2084);
nor U1485 (N_1485,In_840,In_2582);
nor U1486 (N_1486,In_876,In_747);
nand U1487 (N_1487,In_554,In_2138);
nand U1488 (N_1488,In_996,In_2273);
and U1489 (N_1489,In_1341,In_2905);
or U1490 (N_1490,In_1646,In_1596);
nand U1491 (N_1491,In_834,In_1900);
nor U1492 (N_1492,In_2019,In_2728);
and U1493 (N_1493,In_2411,In_1957);
nor U1494 (N_1494,In_237,In_2484);
or U1495 (N_1495,In_1410,In_2659);
and U1496 (N_1496,In_324,In_2038);
or U1497 (N_1497,In_2520,In_178);
or U1498 (N_1498,In_756,In_1985);
and U1499 (N_1499,In_1004,In_239);
nor U1500 (N_1500,In_2588,In_540);
nor U1501 (N_1501,In_297,In_2246);
and U1502 (N_1502,In_962,In_1098);
and U1503 (N_1503,In_32,In_2300);
xnor U1504 (N_1504,In_549,In_1186);
or U1505 (N_1505,In_245,In_813);
and U1506 (N_1506,In_2534,In_2445);
or U1507 (N_1507,In_836,In_2088);
or U1508 (N_1508,In_2030,In_232);
nand U1509 (N_1509,In_2843,In_1364);
nor U1510 (N_1510,In_2810,In_2896);
nand U1511 (N_1511,In_213,In_1458);
or U1512 (N_1512,In_903,In_2127);
nor U1513 (N_1513,In_2856,In_313);
nand U1514 (N_1514,In_465,In_174);
or U1515 (N_1515,In_741,In_35);
nor U1516 (N_1516,In_1716,In_2900);
or U1517 (N_1517,In_404,In_587);
and U1518 (N_1518,In_171,In_1667);
nor U1519 (N_1519,In_2453,In_26);
nor U1520 (N_1520,In_1484,In_1269);
xor U1521 (N_1521,In_1938,In_786);
nor U1522 (N_1522,In_1447,In_1863);
or U1523 (N_1523,In_1589,In_1696);
xor U1524 (N_1524,In_2701,In_2956);
nand U1525 (N_1525,In_2643,In_334);
and U1526 (N_1526,In_2538,In_132);
xnor U1527 (N_1527,In_2709,In_1595);
or U1528 (N_1528,In_1851,In_1806);
xnor U1529 (N_1529,In_210,In_1033);
xnor U1530 (N_1530,In_757,In_956);
and U1531 (N_1531,In_34,In_354);
nor U1532 (N_1532,In_862,In_724);
nand U1533 (N_1533,In_2730,In_326);
and U1534 (N_1534,In_2969,In_2019);
or U1535 (N_1535,In_1629,In_917);
or U1536 (N_1536,In_995,In_668);
nor U1537 (N_1537,In_262,In_2427);
nor U1538 (N_1538,In_1664,In_2234);
nor U1539 (N_1539,In_1802,In_182);
or U1540 (N_1540,In_2415,In_247);
or U1541 (N_1541,In_644,In_1906);
nor U1542 (N_1542,In_595,In_2751);
nor U1543 (N_1543,In_626,In_277);
nor U1544 (N_1544,In_1053,In_1519);
and U1545 (N_1545,In_2793,In_534);
nand U1546 (N_1546,In_2927,In_1383);
and U1547 (N_1547,In_1157,In_1824);
nor U1548 (N_1548,In_1205,In_893);
or U1549 (N_1549,In_1916,In_1655);
nor U1550 (N_1550,In_1111,In_2650);
nor U1551 (N_1551,In_2199,In_1203);
and U1552 (N_1552,In_2918,In_1370);
and U1553 (N_1553,In_1204,In_1089);
nor U1554 (N_1554,In_732,In_2550);
or U1555 (N_1555,In_658,In_1631);
nand U1556 (N_1556,In_1587,In_2575);
nand U1557 (N_1557,In_2513,In_206);
nand U1558 (N_1558,In_67,In_3);
nand U1559 (N_1559,In_47,In_2075);
or U1560 (N_1560,In_893,In_2786);
xnor U1561 (N_1561,In_1051,In_611);
nand U1562 (N_1562,In_1036,In_934);
and U1563 (N_1563,In_2625,In_1104);
and U1564 (N_1564,In_2676,In_779);
xnor U1565 (N_1565,In_1034,In_888);
and U1566 (N_1566,In_1646,In_2090);
xor U1567 (N_1567,In_209,In_2930);
xor U1568 (N_1568,In_2200,In_2542);
nor U1569 (N_1569,In_792,In_1055);
nor U1570 (N_1570,In_2993,In_86);
and U1571 (N_1571,In_2364,In_2887);
nand U1572 (N_1572,In_2131,In_2588);
or U1573 (N_1573,In_1604,In_1450);
or U1574 (N_1574,In_500,In_812);
and U1575 (N_1575,In_2816,In_1574);
or U1576 (N_1576,In_935,In_1491);
nor U1577 (N_1577,In_471,In_272);
nand U1578 (N_1578,In_152,In_300);
or U1579 (N_1579,In_713,In_2528);
or U1580 (N_1580,In_2715,In_2763);
nor U1581 (N_1581,In_2607,In_2097);
nand U1582 (N_1582,In_2636,In_1462);
and U1583 (N_1583,In_604,In_212);
nand U1584 (N_1584,In_2579,In_1167);
nor U1585 (N_1585,In_709,In_1301);
and U1586 (N_1586,In_845,In_1515);
nor U1587 (N_1587,In_1028,In_1711);
nand U1588 (N_1588,In_1382,In_395);
or U1589 (N_1589,In_1870,In_502);
or U1590 (N_1590,In_322,In_194);
nor U1591 (N_1591,In_368,In_1017);
or U1592 (N_1592,In_1440,In_1417);
or U1593 (N_1593,In_779,In_2878);
nor U1594 (N_1594,In_688,In_2640);
or U1595 (N_1595,In_594,In_2265);
or U1596 (N_1596,In_221,In_2404);
or U1597 (N_1597,In_513,In_1286);
nand U1598 (N_1598,In_1261,In_2168);
and U1599 (N_1599,In_1017,In_2575);
nor U1600 (N_1600,In_297,In_1468);
nand U1601 (N_1601,In_41,In_2841);
and U1602 (N_1602,In_2736,In_2371);
nand U1603 (N_1603,In_2456,In_1601);
and U1604 (N_1604,In_2786,In_1116);
and U1605 (N_1605,In_2759,In_431);
or U1606 (N_1606,In_2855,In_1293);
or U1607 (N_1607,In_1220,In_1828);
or U1608 (N_1608,In_2272,In_253);
nor U1609 (N_1609,In_1282,In_820);
or U1610 (N_1610,In_1872,In_19);
nor U1611 (N_1611,In_2056,In_215);
or U1612 (N_1612,In_1267,In_2754);
and U1613 (N_1613,In_224,In_1323);
or U1614 (N_1614,In_2546,In_1978);
xor U1615 (N_1615,In_99,In_1896);
nand U1616 (N_1616,In_2815,In_509);
nand U1617 (N_1617,In_1403,In_1250);
and U1618 (N_1618,In_677,In_1044);
xor U1619 (N_1619,In_1374,In_1925);
nor U1620 (N_1620,In_1047,In_227);
and U1621 (N_1621,In_1646,In_1430);
or U1622 (N_1622,In_2216,In_151);
or U1623 (N_1623,In_1886,In_1530);
xnor U1624 (N_1624,In_2805,In_231);
and U1625 (N_1625,In_2198,In_2053);
or U1626 (N_1626,In_267,In_2687);
or U1627 (N_1627,In_1094,In_1549);
nand U1628 (N_1628,In_163,In_1666);
nand U1629 (N_1629,In_1174,In_2204);
or U1630 (N_1630,In_2367,In_598);
or U1631 (N_1631,In_678,In_1673);
nor U1632 (N_1632,In_2841,In_1315);
or U1633 (N_1633,In_595,In_914);
nand U1634 (N_1634,In_2099,In_2753);
and U1635 (N_1635,In_2521,In_1274);
nand U1636 (N_1636,In_1789,In_2794);
or U1637 (N_1637,In_196,In_2368);
nor U1638 (N_1638,In_525,In_1658);
nor U1639 (N_1639,In_2378,In_2508);
or U1640 (N_1640,In_2075,In_2413);
or U1641 (N_1641,In_418,In_1786);
nand U1642 (N_1642,In_1249,In_1824);
nor U1643 (N_1643,In_1941,In_384);
nand U1644 (N_1644,In_2720,In_2696);
or U1645 (N_1645,In_1464,In_67);
or U1646 (N_1646,In_2606,In_1426);
or U1647 (N_1647,In_2958,In_1993);
nand U1648 (N_1648,In_1279,In_2915);
nand U1649 (N_1649,In_1250,In_1012);
and U1650 (N_1650,In_2121,In_2982);
or U1651 (N_1651,In_182,In_339);
or U1652 (N_1652,In_1660,In_203);
xnor U1653 (N_1653,In_347,In_2292);
nand U1654 (N_1654,In_30,In_1523);
or U1655 (N_1655,In_999,In_11);
xor U1656 (N_1656,In_1315,In_2944);
nor U1657 (N_1657,In_2326,In_381);
xnor U1658 (N_1658,In_2914,In_1526);
nor U1659 (N_1659,In_1233,In_350);
or U1660 (N_1660,In_280,In_256);
xnor U1661 (N_1661,In_327,In_1290);
or U1662 (N_1662,In_2128,In_1315);
and U1663 (N_1663,In_2586,In_397);
and U1664 (N_1664,In_1153,In_903);
and U1665 (N_1665,In_1393,In_579);
nor U1666 (N_1666,In_1103,In_2779);
nand U1667 (N_1667,In_376,In_852);
nor U1668 (N_1668,In_1469,In_2038);
nand U1669 (N_1669,In_1934,In_1033);
nor U1670 (N_1670,In_2478,In_478);
nand U1671 (N_1671,In_2454,In_2582);
xnor U1672 (N_1672,In_1250,In_2024);
nor U1673 (N_1673,In_156,In_1458);
or U1674 (N_1674,In_1969,In_1461);
and U1675 (N_1675,In_1873,In_260);
nor U1676 (N_1676,In_578,In_1395);
nand U1677 (N_1677,In_458,In_2334);
nand U1678 (N_1678,In_1209,In_1872);
nand U1679 (N_1679,In_1979,In_1726);
and U1680 (N_1680,In_842,In_1581);
nand U1681 (N_1681,In_1144,In_85);
and U1682 (N_1682,In_2989,In_2011);
nor U1683 (N_1683,In_1039,In_1011);
nor U1684 (N_1684,In_1233,In_856);
nor U1685 (N_1685,In_7,In_1262);
or U1686 (N_1686,In_890,In_2672);
and U1687 (N_1687,In_2463,In_527);
and U1688 (N_1688,In_1241,In_993);
or U1689 (N_1689,In_487,In_2701);
nand U1690 (N_1690,In_1650,In_743);
or U1691 (N_1691,In_2292,In_1683);
nand U1692 (N_1692,In_883,In_1568);
and U1693 (N_1693,In_628,In_2935);
xor U1694 (N_1694,In_2393,In_259);
or U1695 (N_1695,In_1265,In_457);
and U1696 (N_1696,In_386,In_2567);
and U1697 (N_1697,In_2280,In_1190);
or U1698 (N_1698,In_2197,In_2407);
nor U1699 (N_1699,In_660,In_2508);
and U1700 (N_1700,In_1887,In_1227);
nand U1701 (N_1701,In_131,In_1219);
nor U1702 (N_1702,In_1189,In_884);
or U1703 (N_1703,In_139,In_291);
and U1704 (N_1704,In_82,In_1729);
nand U1705 (N_1705,In_2142,In_1787);
nor U1706 (N_1706,In_1834,In_515);
or U1707 (N_1707,In_1378,In_263);
nor U1708 (N_1708,In_871,In_1875);
nor U1709 (N_1709,In_2561,In_2665);
nor U1710 (N_1710,In_2225,In_430);
and U1711 (N_1711,In_387,In_2099);
xor U1712 (N_1712,In_1389,In_2366);
nand U1713 (N_1713,In_980,In_2805);
nor U1714 (N_1714,In_2905,In_1436);
nor U1715 (N_1715,In_1145,In_1792);
or U1716 (N_1716,In_738,In_946);
nand U1717 (N_1717,In_163,In_672);
nand U1718 (N_1718,In_2166,In_2087);
or U1719 (N_1719,In_1725,In_2835);
or U1720 (N_1720,In_1465,In_1056);
nand U1721 (N_1721,In_911,In_441);
and U1722 (N_1722,In_1743,In_1591);
nand U1723 (N_1723,In_1152,In_1601);
xor U1724 (N_1724,In_696,In_535);
and U1725 (N_1725,In_702,In_2106);
nor U1726 (N_1726,In_547,In_1930);
or U1727 (N_1727,In_514,In_1959);
nand U1728 (N_1728,In_1434,In_1435);
nor U1729 (N_1729,In_2919,In_2726);
nor U1730 (N_1730,In_2601,In_1423);
nor U1731 (N_1731,In_1762,In_2128);
nor U1732 (N_1732,In_2637,In_156);
and U1733 (N_1733,In_2721,In_2218);
xnor U1734 (N_1734,In_786,In_1990);
and U1735 (N_1735,In_446,In_2599);
xnor U1736 (N_1736,In_901,In_2334);
nor U1737 (N_1737,In_1748,In_1660);
or U1738 (N_1738,In_1,In_52);
nor U1739 (N_1739,In_891,In_1889);
nor U1740 (N_1740,In_762,In_1222);
and U1741 (N_1741,In_83,In_2095);
or U1742 (N_1742,In_2733,In_795);
or U1743 (N_1743,In_424,In_1622);
nand U1744 (N_1744,In_2826,In_1239);
xor U1745 (N_1745,In_1353,In_1677);
or U1746 (N_1746,In_2368,In_2861);
nand U1747 (N_1747,In_1997,In_2052);
nor U1748 (N_1748,In_446,In_2141);
or U1749 (N_1749,In_2116,In_1163);
nand U1750 (N_1750,In_2738,In_2763);
nand U1751 (N_1751,In_1376,In_1488);
nand U1752 (N_1752,In_1660,In_801);
nor U1753 (N_1753,In_1231,In_1069);
and U1754 (N_1754,In_1263,In_787);
or U1755 (N_1755,In_2905,In_551);
or U1756 (N_1756,In_79,In_1368);
nor U1757 (N_1757,In_2575,In_1533);
or U1758 (N_1758,In_2658,In_51);
xnor U1759 (N_1759,In_1332,In_370);
and U1760 (N_1760,In_1585,In_1729);
or U1761 (N_1761,In_1722,In_2590);
or U1762 (N_1762,In_2720,In_2952);
xor U1763 (N_1763,In_2530,In_1795);
or U1764 (N_1764,In_2358,In_1695);
or U1765 (N_1765,In_121,In_2348);
and U1766 (N_1766,In_192,In_2847);
nor U1767 (N_1767,In_1957,In_489);
nand U1768 (N_1768,In_679,In_2911);
and U1769 (N_1769,In_1568,In_56);
and U1770 (N_1770,In_190,In_827);
and U1771 (N_1771,In_2366,In_1623);
nand U1772 (N_1772,In_2798,In_2199);
nand U1773 (N_1773,In_448,In_1108);
or U1774 (N_1774,In_1146,In_1847);
nor U1775 (N_1775,In_16,In_28);
and U1776 (N_1776,In_2479,In_1688);
nor U1777 (N_1777,In_2914,In_2399);
nor U1778 (N_1778,In_2468,In_1514);
nor U1779 (N_1779,In_1407,In_1078);
xnor U1780 (N_1780,In_1177,In_2363);
xor U1781 (N_1781,In_1299,In_1637);
and U1782 (N_1782,In_344,In_496);
or U1783 (N_1783,In_78,In_2895);
and U1784 (N_1784,In_1762,In_2505);
and U1785 (N_1785,In_1223,In_213);
nand U1786 (N_1786,In_184,In_118);
xnor U1787 (N_1787,In_2611,In_1546);
or U1788 (N_1788,In_2362,In_1301);
xnor U1789 (N_1789,In_1981,In_2937);
or U1790 (N_1790,In_2526,In_1970);
nand U1791 (N_1791,In_2785,In_2009);
xor U1792 (N_1792,In_39,In_2785);
nor U1793 (N_1793,In_38,In_2964);
and U1794 (N_1794,In_405,In_335);
nor U1795 (N_1795,In_1422,In_2910);
or U1796 (N_1796,In_1827,In_2503);
nor U1797 (N_1797,In_2884,In_977);
or U1798 (N_1798,In_129,In_2341);
or U1799 (N_1799,In_771,In_1937);
nand U1800 (N_1800,In_2788,In_2285);
nor U1801 (N_1801,In_1108,In_199);
nand U1802 (N_1802,In_1280,In_685);
nor U1803 (N_1803,In_2376,In_2628);
and U1804 (N_1804,In_762,In_542);
nor U1805 (N_1805,In_1238,In_489);
nor U1806 (N_1806,In_1286,In_2389);
nor U1807 (N_1807,In_2053,In_378);
xor U1808 (N_1808,In_1139,In_2180);
and U1809 (N_1809,In_189,In_730);
and U1810 (N_1810,In_1626,In_2215);
nand U1811 (N_1811,In_1063,In_2626);
xnor U1812 (N_1812,In_236,In_1442);
xnor U1813 (N_1813,In_1425,In_2296);
and U1814 (N_1814,In_1471,In_457);
nand U1815 (N_1815,In_902,In_2650);
nor U1816 (N_1816,In_2390,In_877);
nor U1817 (N_1817,In_404,In_1668);
nor U1818 (N_1818,In_1671,In_1215);
nand U1819 (N_1819,In_2759,In_303);
xnor U1820 (N_1820,In_1454,In_802);
and U1821 (N_1821,In_10,In_2209);
nor U1822 (N_1822,In_2010,In_1091);
nand U1823 (N_1823,In_1130,In_2768);
nand U1824 (N_1824,In_767,In_173);
or U1825 (N_1825,In_1836,In_1341);
or U1826 (N_1826,In_837,In_921);
nor U1827 (N_1827,In_1088,In_2858);
and U1828 (N_1828,In_818,In_824);
nor U1829 (N_1829,In_1269,In_1886);
nor U1830 (N_1830,In_1123,In_2491);
and U1831 (N_1831,In_2654,In_788);
and U1832 (N_1832,In_2181,In_315);
nand U1833 (N_1833,In_1869,In_2619);
and U1834 (N_1834,In_2119,In_1168);
nand U1835 (N_1835,In_2719,In_2182);
nor U1836 (N_1836,In_254,In_1717);
nor U1837 (N_1837,In_1102,In_726);
nor U1838 (N_1838,In_1830,In_2791);
or U1839 (N_1839,In_2076,In_1082);
or U1840 (N_1840,In_1222,In_990);
or U1841 (N_1841,In_1988,In_2097);
nand U1842 (N_1842,In_2144,In_608);
or U1843 (N_1843,In_1,In_2012);
xnor U1844 (N_1844,In_1857,In_2528);
and U1845 (N_1845,In_1520,In_2386);
nor U1846 (N_1846,In_464,In_2184);
nand U1847 (N_1847,In_2599,In_1370);
and U1848 (N_1848,In_2391,In_1012);
nor U1849 (N_1849,In_1874,In_2094);
or U1850 (N_1850,In_1855,In_2809);
and U1851 (N_1851,In_1447,In_2977);
and U1852 (N_1852,In_2922,In_826);
nor U1853 (N_1853,In_1897,In_204);
xnor U1854 (N_1854,In_620,In_2823);
nor U1855 (N_1855,In_1220,In_834);
and U1856 (N_1856,In_579,In_2238);
nor U1857 (N_1857,In_993,In_367);
and U1858 (N_1858,In_1774,In_1523);
or U1859 (N_1859,In_2196,In_1994);
nand U1860 (N_1860,In_1293,In_2513);
xor U1861 (N_1861,In_2228,In_2507);
nor U1862 (N_1862,In_2270,In_2301);
nand U1863 (N_1863,In_2133,In_686);
and U1864 (N_1864,In_2202,In_2673);
and U1865 (N_1865,In_1757,In_293);
nor U1866 (N_1866,In_859,In_729);
or U1867 (N_1867,In_1232,In_2272);
and U1868 (N_1868,In_348,In_865);
and U1869 (N_1869,In_474,In_1259);
nand U1870 (N_1870,In_501,In_2677);
and U1871 (N_1871,In_156,In_1921);
and U1872 (N_1872,In_1125,In_58);
or U1873 (N_1873,In_1853,In_2619);
or U1874 (N_1874,In_1099,In_1747);
or U1875 (N_1875,In_961,In_419);
or U1876 (N_1876,In_2072,In_302);
or U1877 (N_1877,In_1834,In_2285);
or U1878 (N_1878,In_2016,In_2963);
and U1879 (N_1879,In_340,In_1552);
nor U1880 (N_1880,In_2654,In_444);
or U1881 (N_1881,In_2762,In_1145);
nor U1882 (N_1882,In_1285,In_1890);
and U1883 (N_1883,In_1878,In_903);
and U1884 (N_1884,In_2886,In_1172);
nand U1885 (N_1885,In_2166,In_1640);
nand U1886 (N_1886,In_2887,In_1603);
and U1887 (N_1887,In_591,In_787);
nand U1888 (N_1888,In_2250,In_2919);
or U1889 (N_1889,In_1040,In_1501);
nand U1890 (N_1890,In_543,In_1078);
and U1891 (N_1891,In_2734,In_1298);
or U1892 (N_1892,In_2723,In_1595);
and U1893 (N_1893,In_1594,In_380);
nand U1894 (N_1894,In_1210,In_2919);
or U1895 (N_1895,In_1834,In_2272);
and U1896 (N_1896,In_1695,In_383);
nor U1897 (N_1897,In_1177,In_2134);
or U1898 (N_1898,In_1635,In_1369);
or U1899 (N_1899,In_1438,In_1497);
and U1900 (N_1900,In_2180,In_1072);
nand U1901 (N_1901,In_1034,In_2944);
nand U1902 (N_1902,In_2016,In_1551);
or U1903 (N_1903,In_2416,In_1756);
nor U1904 (N_1904,In_2206,In_414);
xor U1905 (N_1905,In_880,In_2873);
nor U1906 (N_1906,In_2146,In_1040);
and U1907 (N_1907,In_40,In_453);
and U1908 (N_1908,In_2021,In_1505);
nand U1909 (N_1909,In_1738,In_192);
nand U1910 (N_1910,In_1843,In_1500);
and U1911 (N_1911,In_140,In_2512);
nor U1912 (N_1912,In_1410,In_2497);
nor U1913 (N_1913,In_2202,In_1941);
and U1914 (N_1914,In_237,In_2664);
and U1915 (N_1915,In_500,In_286);
nand U1916 (N_1916,In_729,In_649);
nand U1917 (N_1917,In_1101,In_2753);
or U1918 (N_1918,In_1247,In_2159);
xnor U1919 (N_1919,In_107,In_2626);
or U1920 (N_1920,In_2773,In_2660);
nand U1921 (N_1921,In_2612,In_2635);
nor U1922 (N_1922,In_1483,In_10);
nand U1923 (N_1923,In_920,In_1089);
nand U1924 (N_1924,In_2143,In_571);
or U1925 (N_1925,In_197,In_1027);
and U1926 (N_1926,In_2198,In_1373);
xnor U1927 (N_1927,In_818,In_354);
nor U1928 (N_1928,In_2421,In_2885);
nand U1929 (N_1929,In_2656,In_2407);
nor U1930 (N_1930,In_2681,In_1974);
xnor U1931 (N_1931,In_1556,In_618);
nand U1932 (N_1932,In_728,In_1789);
xnor U1933 (N_1933,In_1431,In_2339);
or U1934 (N_1934,In_1551,In_526);
and U1935 (N_1935,In_118,In_956);
and U1936 (N_1936,In_384,In_37);
and U1937 (N_1937,In_2722,In_1938);
nor U1938 (N_1938,In_1604,In_516);
xnor U1939 (N_1939,In_2574,In_125);
and U1940 (N_1940,In_1791,In_2874);
or U1941 (N_1941,In_480,In_2371);
nand U1942 (N_1942,In_468,In_357);
nand U1943 (N_1943,In_1571,In_2858);
nor U1944 (N_1944,In_838,In_557);
nand U1945 (N_1945,In_415,In_774);
or U1946 (N_1946,In_812,In_1111);
nor U1947 (N_1947,In_538,In_2521);
xnor U1948 (N_1948,In_2569,In_596);
nor U1949 (N_1949,In_1627,In_1798);
nor U1950 (N_1950,In_2578,In_1542);
and U1951 (N_1951,In_2330,In_448);
nand U1952 (N_1952,In_144,In_858);
and U1953 (N_1953,In_1645,In_1504);
or U1954 (N_1954,In_2779,In_1546);
nand U1955 (N_1955,In_128,In_2917);
xor U1956 (N_1956,In_801,In_477);
and U1957 (N_1957,In_363,In_2103);
nand U1958 (N_1958,In_2328,In_1821);
nand U1959 (N_1959,In_750,In_984);
nor U1960 (N_1960,In_1376,In_2641);
and U1961 (N_1961,In_2809,In_2948);
or U1962 (N_1962,In_1492,In_1658);
or U1963 (N_1963,In_908,In_1947);
nor U1964 (N_1964,In_61,In_1852);
xnor U1965 (N_1965,In_362,In_106);
and U1966 (N_1966,In_2204,In_828);
nor U1967 (N_1967,In_2821,In_2857);
and U1968 (N_1968,In_2654,In_913);
nor U1969 (N_1969,In_2328,In_2935);
and U1970 (N_1970,In_933,In_1757);
nor U1971 (N_1971,In_573,In_349);
or U1972 (N_1972,In_2653,In_2454);
and U1973 (N_1973,In_922,In_434);
nor U1974 (N_1974,In_2478,In_925);
or U1975 (N_1975,In_2828,In_121);
nand U1976 (N_1976,In_672,In_2640);
and U1977 (N_1977,In_491,In_1220);
and U1978 (N_1978,In_2016,In_1710);
and U1979 (N_1979,In_1438,In_411);
nor U1980 (N_1980,In_1156,In_165);
nor U1981 (N_1981,In_666,In_2551);
nand U1982 (N_1982,In_2284,In_2622);
xnor U1983 (N_1983,In_44,In_1141);
xor U1984 (N_1984,In_223,In_909);
and U1985 (N_1985,In_797,In_891);
nor U1986 (N_1986,In_454,In_1740);
xor U1987 (N_1987,In_1640,In_1684);
nor U1988 (N_1988,In_1210,In_541);
or U1989 (N_1989,In_2199,In_2423);
nor U1990 (N_1990,In_1257,In_1112);
or U1991 (N_1991,In_293,In_1072);
or U1992 (N_1992,In_192,In_1000);
and U1993 (N_1993,In_1684,In_2480);
and U1994 (N_1994,In_312,In_1139);
and U1995 (N_1995,In_2101,In_1712);
nand U1996 (N_1996,In_2585,In_2948);
nand U1997 (N_1997,In_554,In_2154);
nor U1998 (N_1998,In_1136,In_584);
nand U1999 (N_1999,In_1837,In_2193);
nor U2000 (N_2000,In_993,In_418);
xor U2001 (N_2001,In_2674,In_1683);
nor U2002 (N_2002,In_188,In_2029);
xor U2003 (N_2003,In_1842,In_1049);
xor U2004 (N_2004,In_1603,In_2069);
nand U2005 (N_2005,In_1594,In_307);
nand U2006 (N_2006,In_1539,In_2018);
or U2007 (N_2007,In_762,In_2221);
or U2008 (N_2008,In_2326,In_2172);
xnor U2009 (N_2009,In_913,In_2311);
nor U2010 (N_2010,In_607,In_1708);
and U2011 (N_2011,In_1406,In_715);
nor U2012 (N_2012,In_625,In_2964);
and U2013 (N_2013,In_1279,In_2901);
or U2014 (N_2014,In_1612,In_250);
nor U2015 (N_2015,In_309,In_336);
or U2016 (N_2016,In_2663,In_552);
nand U2017 (N_2017,In_1362,In_2778);
nor U2018 (N_2018,In_2545,In_1863);
or U2019 (N_2019,In_1647,In_1111);
or U2020 (N_2020,In_595,In_1870);
or U2021 (N_2021,In_1866,In_1009);
or U2022 (N_2022,In_107,In_2715);
nor U2023 (N_2023,In_2735,In_2942);
nor U2024 (N_2024,In_1630,In_2287);
nand U2025 (N_2025,In_1409,In_2319);
or U2026 (N_2026,In_204,In_2819);
nor U2027 (N_2027,In_337,In_657);
nor U2028 (N_2028,In_2212,In_372);
and U2029 (N_2029,In_344,In_429);
and U2030 (N_2030,In_791,In_539);
nor U2031 (N_2031,In_2842,In_1475);
nor U2032 (N_2032,In_845,In_1193);
or U2033 (N_2033,In_1546,In_852);
or U2034 (N_2034,In_877,In_1165);
or U2035 (N_2035,In_1964,In_650);
nor U2036 (N_2036,In_796,In_1383);
nand U2037 (N_2037,In_66,In_1119);
nand U2038 (N_2038,In_855,In_2509);
nand U2039 (N_2039,In_377,In_1238);
xnor U2040 (N_2040,In_2503,In_712);
or U2041 (N_2041,In_2413,In_2665);
nand U2042 (N_2042,In_1374,In_2207);
and U2043 (N_2043,In_129,In_295);
nor U2044 (N_2044,In_214,In_2846);
and U2045 (N_2045,In_2579,In_2746);
nand U2046 (N_2046,In_320,In_1584);
and U2047 (N_2047,In_2643,In_16);
nand U2048 (N_2048,In_2009,In_2120);
nand U2049 (N_2049,In_1355,In_330);
and U2050 (N_2050,In_456,In_1581);
nand U2051 (N_2051,In_1558,In_2315);
and U2052 (N_2052,In_1916,In_1495);
nor U2053 (N_2053,In_2255,In_916);
nor U2054 (N_2054,In_1101,In_309);
or U2055 (N_2055,In_2162,In_1003);
and U2056 (N_2056,In_2440,In_2723);
and U2057 (N_2057,In_1294,In_2307);
and U2058 (N_2058,In_973,In_2097);
or U2059 (N_2059,In_375,In_1021);
or U2060 (N_2060,In_1640,In_2246);
or U2061 (N_2061,In_1447,In_581);
and U2062 (N_2062,In_900,In_1011);
or U2063 (N_2063,In_1280,In_1434);
and U2064 (N_2064,In_2882,In_1506);
nand U2065 (N_2065,In_1383,In_2165);
and U2066 (N_2066,In_13,In_2287);
or U2067 (N_2067,In_1479,In_1584);
nand U2068 (N_2068,In_2187,In_582);
nand U2069 (N_2069,In_2975,In_1658);
or U2070 (N_2070,In_64,In_1721);
and U2071 (N_2071,In_1158,In_2007);
nor U2072 (N_2072,In_2437,In_1570);
or U2073 (N_2073,In_2822,In_2296);
xnor U2074 (N_2074,In_1562,In_162);
nand U2075 (N_2075,In_1748,In_1001);
nor U2076 (N_2076,In_2262,In_177);
nand U2077 (N_2077,In_1456,In_148);
nand U2078 (N_2078,In_2521,In_2343);
nor U2079 (N_2079,In_2760,In_2841);
or U2080 (N_2080,In_1482,In_2936);
and U2081 (N_2081,In_103,In_1247);
nor U2082 (N_2082,In_2413,In_1666);
nand U2083 (N_2083,In_2060,In_498);
and U2084 (N_2084,In_1727,In_2215);
nor U2085 (N_2085,In_695,In_522);
or U2086 (N_2086,In_1971,In_2552);
or U2087 (N_2087,In_2467,In_1255);
or U2088 (N_2088,In_106,In_826);
nor U2089 (N_2089,In_1152,In_1432);
nand U2090 (N_2090,In_1532,In_781);
xnor U2091 (N_2091,In_612,In_1433);
or U2092 (N_2092,In_2299,In_1589);
nand U2093 (N_2093,In_1722,In_1964);
or U2094 (N_2094,In_2747,In_2767);
xnor U2095 (N_2095,In_2109,In_2236);
nand U2096 (N_2096,In_2794,In_2427);
and U2097 (N_2097,In_1845,In_2332);
nand U2098 (N_2098,In_2221,In_40);
nor U2099 (N_2099,In_1977,In_657);
nor U2100 (N_2100,In_920,In_1859);
nand U2101 (N_2101,In_1935,In_2718);
nor U2102 (N_2102,In_1527,In_2173);
xnor U2103 (N_2103,In_399,In_277);
xor U2104 (N_2104,In_2794,In_727);
and U2105 (N_2105,In_584,In_2046);
nand U2106 (N_2106,In_1118,In_1723);
nand U2107 (N_2107,In_2657,In_2483);
nand U2108 (N_2108,In_171,In_89);
or U2109 (N_2109,In_2655,In_404);
xor U2110 (N_2110,In_690,In_1589);
or U2111 (N_2111,In_1178,In_1252);
and U2112 (N_2112,In_301,In_1517);
or U2113 (N_2113,In_2570,In_1365);
xor U2114 (N_2114,In_1912,In_2513);
or U2115 (N_2115,In_1914,In_1432);
or U2116 (N_2116,In_1266,In_2004);
nand U2117 (N_2117,In_1266,In_1638);
and U2118 (N_2118,In_2199,In_1010);
or U2119 (N_2119,In_2489,In_2757);
nand U2120 (N_2120,In_1206,In_258);
or U2121 (N_2121,In_92,In_287);
nand U2122 (N_2122,In_2432,In_888);
nand U2123 (N_2123,In_2303,In_2288);
nand U2124 (N_2124,In_2760,In_2047);
or U2125 (N_2125,In_1718,In_432);
nand U2126 (N_2126,In_1561,In_1319);
nor U2127 (N_2127,In_1558,In_2607);
and U2128 (N_2128,In_502,In_2732);
nand U2129 (N_2129,In_1472,In_1583);
nor U2130 (N_2130,In_2223,In_1072);
nor U2131 (N_2131,In_113,In_2908);
nand U2132 (N_2132,In_2536,In_2033);
nor U2133 (N_2133,In_1016,In_2600);
or U2134 (N_2134,In_2793,In_1596);
nand U2135 (N_2135,In_494,In_1809);
xnor U2136 (N_2136,In_923,In_1891);
nand U2137 (N_2137,In_1640,In_1883);
and U2138 (N_2138,In_2222,In_1173);
nor U2139 (N_2139,In_869,In_2791);
nor U2140 (N_2140,In_583,In_751);
nand U2141 (N_2141,In_1593,In_2343);
or U2142 (N_2142,In_1359,In_1473);
nor U2143 (N_2143,In_2279,In_1321);
or U2144 (N_2144,In_597,In_2699);
nor U2145 (N_2145,In_1551,In_2428);
nor U2146 (N_2146,In_2056,In_2419);
nand U2147 (N_2147,In_361,In_2812);
nor U2148 (N_2148,In_2284,In_226);
nor U2149 (N_2149,In_1607,In_1572);
or U2150 (N_2150,In_2472,In_127);
nand U2151 (N_2151,In_630,In_134);
nand U2152 (N_2152,In_996,In_131);
and U2153 (N_2153,In_28,In_1994);
and U2154 (N_2154,In_21,In_363);
nor U2155 (N_2155,In_2558,In_330);
and U2156 (N_2156,In_1059,In_2587);
nor U2157 (N_2157,In_1671,In_1367);
nor U2158 (N_2158,In_708,In_2863);
nor U2159 (N_2159,In_1320,In_822);
or U2160 (N_2160,In_991,In_1988);
nand U2161 (N_2161,In_2840,In_1563);
nand U2162 (N_2162,In_1922,In_911);
or U2163 (N_2163,In_34,In_2789);
or U2164 (N_2164,In_54,In_2439);
nor U2165 (N_2165,In_1863,In_145);
or U2166 (N_2166,In_1598,In_1866);
nor U2167 (N_2167,In_17,In_329);
or U2168 (N_2168,In_2924,In_734);
nor U2169 (N_2169,In_998,In_2849);
nor U2170 (N_2170,In_1513,In_1314);
nor U2171 (N_2171,In_1961,In_710);
nor U2172 (N_2172,In_2133,In_536);
nor U2173 (N_2173,In_1397,In_531);
nor U2174 (N_2174,In_2462,In_70);
nor U2175 (N_2175,In_2715,In_2575);
nand U2176 (N_2176,In_211,In_304);
nor U2177 (N_2177,In_150,In_493);
nor U2178 (N_2178,In_1694,In_2965);
and U2179 (N_2179,In_2092,In_143);
nor U2180 (N_2180,In_2212,In_1584);
nand U2181 (N_2181,In_1685,In_455);
or U2182 (N_2182,In_120,In_952);
nand U2183 (N_2183,In_1406,In_1458);
nor U2184 (N_2184,In_1565,In_1288);
nand U2185 (N_2185,In_2848,In_2943);
and U2186 (N_2186,In_881,In_525);
or U2187 (N_2187,In_1404,In_2225);
nand U2188 (N_2188,In_2075,In_875);
and U2189 (N_2189,In_260,In_1919);
nand U2190 (N_2190,In_839,In_951);
nand U2191 (N_2191,In_784,In_1645);
nor U2192 (N_2192,In_531,In_2095);
or U2193 (N_2193,In_2555,In_1093);
nor U2194 (N_2194,In_2227,In_913);
xnor U2195 (N_2195,In_902,In_1076);
nor U2196 (N_2196,In_1919,In_1708);
and U2197 (N_2197,In_662,In_1238);
and U2198 (N_2198,In_1998,In_241);
or U2199 (N_2199,In_2597,In_339);
nand U2200 (N_2200,In_607,In_2091);
nand U2201 (N_2201,In_1261,In_2727);
nand U2202 (N_2202,In_1910,In_1924);
and U2203 (N_2203,In_507,In_523);
or U2204 (N_2204,In_1303,In_74);
xor U2205 (N_2205,In_277,In_2064);
and U2206 (N_2206,In_1229,In_2986);
or U2207 (N_2207,In_1574,In_309);
nand U2208 (N_2208,In_2108,In_2517);
nor U2209 (N_2209,In_2939,In_2049);
nand U2210 (N_2210,In_2624,In_2177);
or U2211 (N_2211,In_1264,In_263);
nand U2212 (N_2212,In_2254,In_1174);
nor U2213 (N_2213,In_2219,In_2202);
xor U2214 (N_2214,In_812,In_301);
or U2215 (N_2215,In_467,In_1457);
xnor U2216 (N_2216,In_2621,In_1579);
and U2217 (N_2217,In_1668,In_1732);
or U2218 (N_2218,In_1019,In_756);
nor U2219 (N_2219,In_959,In_1104);
nand U2220 (N_2220,In_1007,In_813);
nand U2221 (N_2221,In_2856,In_2885);
nand U2222 (N_2222,In_1968,In_2756);
nor U2223 (N_2223,In_2336,In_134);
xor U2224 (N_2224,In_2073,In_2397);
or U2225 (N_2225,In_1758,In_1217);
xor U2226 (N_2226,In_1908,In_2553);
or U2227 (N_2227,In_2320,In_1725);
nor U2228 (N_2228,In_2756,In_135);
nand U2229 (N_2229,In_719,In_755);
and U2230 (N_2230,In_565,In_1008);
nand U2231 (N_2231,In_2665,In_2485);
and U2232 (N_2232,In_2603,In_1060);
nand U2233 (N_2233,In_590,In_4);
or U2234 (N_2234,In_104,In_146);
nand U2235 (N_2235,In_872,In_825);
xor U2236 (N_2236,In_1735,In_2395);
nand U2237 (N_2237,In_833,In_2995);
or U2238 (N_2238,In_1230,In_2666);
nor U2239 (N_2239,In_576,In_304);
nand U2240 (N_2240,In_1906,In_1620);
and U2241 (N_2241,In_198,In_2256);
nor U2242 (N_2242,In_2667,In_99);
nand U2243 (N_2243,In_455,In_2187);
or U2244 (N_2244,In_689,In_514);
xor U2245 (N_2245,In_2204,In_2288);
xnor U2246 (N_2246,In_2308,In_1334);
nor U2247 (N_2247,In_1701,In_1011);
or U2248 (N_2248,In_1902,In_570);
xor U2249 (N_2249,In_2305,In_1066);
nor U2250 (N_2250,In_321,In_324);
nor U2251 (N_2251,In_1001,In_1275);
nand U2252 (N_2252,In_126,In_1420);
and U2253 (N_2253,In_2843,In_1017);
and U2254 (N_2254,In_1158,In_26);
nor U2255 (N_2255,In_2529,In_972);
nor U2256 (N_2256,In_2925,In_1368);
and U2257 (N_2257,In_1384,In_311);
xnor U2258 (N_2258,In_2361,In_1049);
or U2259 (N_2259,In_967,In_19);
and U2260 (N_2260,In_2510,In_2957);
or U2261 (N_2261,In_1563,In_672);
nand U2262 (N_2262,In_2000,In_760);
nand U2263 (N_2263,In_1779,In_46);
nor U2264 (N_2264,In_5,In_368);
or U2265 (N_2265,In_1265,In_498);
and U2266 (N_2266,In_1772,In_50);
and U2267 (N_2267,In_1044,In_710);
nor U2268 (N_2268,In_2167,In_788);
and U2269 (N_2269,In_1472,In_2499);
nand U2270 (N_2270,In_1612,In_2018);
nand U2271 (N_2271,In_633,In_1048);
nor U2272 (N_2272,In_2067,In_2329);
nand U2273 (N_2273,In_366,In_422);
nor U2274 (N_2274,In_2939,In_1346);
and U2275 (N_2275,In_2569,In_462);
and U2276 (N_2276,In_2994,In_1671);
nand U2277 (N_2277,In_1058,In_1928);
or U2278 (N_2278,In_1510,In_768);
nand U2279 (N_2279,In_2557,In_287);
nand U2280 (N_2280,In_790,In_1668);
or U2281 (N_2281,In_1588,In_1469);
nand U2282 (N_2282,In_1197,In_620);
or U2283 (N_2283,In_2971,In_1029);
nor U2284 (N_2284,In_2824,In_1000);
nand U2285 (N_2285,In_1626,In_181);
nor U2286 (N_2286,In_1620,In_2646);
and U2287 (N_2287,In_2089,In_2820);
nand U2288 (N_2288,In_1662,In_2377);
nand U2289 (N_2289,In_2589,In_74);
nand U2290 (N_2290,In_687,In_246);
nand U2291 (N_2291,In_2076,In_1771);
xor U2292 (N_2292,In_1210,In_2362);
and U2293 (N_2293,In_458,In_762);
or U2294 (N_2294,In_2432,In_2305);
nor U2295 (N_2295,In_1002,In_199);
nor U2296 (N_2296,In_931,In_1646);
nand U2297 (N_2297,In_686,In_2191);
nor U2298 (N_2298,In_1668,In_1993);
or U2299 (N_2299,In_196,In_1439);
or U2300 (N_2300,In_549,In_152);
or U2301 (N_2301,In_594,In_2197);
nand U2302 (N_2302,In_760,In_2830);
nor U2303 (N_2303,In_2811,In_2999);
nand U2304 (N_2304,In_2085,In_648);
xor U2305 (N_2305,In_1792,In_1990);
and U2306 (N_2306,In_1139,In_1775);
or U2307 (N_2307,In_1970,In_1547);
or U2308 (N_2308,In_721,In_2833);
nand U2309 (N_2309,In_2410,In_1703);
nor U2310 (N_2310,In_2363,In_251);
nor U2311 (N_2311,In_156,In_210);
or U2312 (N_2312,In_1297,In_2409);
or U2313 (N_2313,In_1095,In_2365);
nor U2314 (N_2314,In_2896,In_1541);
and U2315 (N_2315,In_656,In_2728);
nor U2316 (N_2316,In_62,In_1255);
and U2317 (N_2317,In_127,In_226);
or U2318 (N_2318,In_2730,In_1115);
nor U2319 (N_2319,In_2875,In_2192);
nor U2320 (N_2320,In_870,In_810);
nand U2321 (N_2321,In_2678,In_828);
xor U2322 (N_2322,In_1755,In_1642);
nor U2323 (N_2323,In_1058,In_1120);
and U2324 (N_2324,In_1263,In_1172);
nor U2325 (N_2325,In_146,In_1160);
or U2326 (N_2326,In_1175,In_1341);
nor U2327 (N_2327,In_1819,In_2640);
nand U2328 (N_2328,In_2837,In_499);
or U2329 (N_2329,In_1877,In_263);
and U2330 (N_2330,In_1373,In_2646);
nor U2331 (N_2331,In_1640,In_1715);
nand U2332 (N_2332,In_1150,In_2270);
and U2333 (N_2333,In_2712,In_523);
and U2334 (N_2334,In_1064,In_2828);
and U2335 (N_2335,In_1769,In_1893);
nand U2336 (N_2336,In_1342,In_2569);
nor U2337 (N_2337,In_194,In_2224);
nor U2338 (N_2338,In_1224,In_2060);
xnor U2339 (N_2339,In_2373,In_1297);
or U2340 (N_2340,In_1457,In_84);
nand U2341 (N_2341,In_203,In_1885);
nand U2342 (N_2342,In_1221,In_1129);
or U2343 (N_2343,In_1003,In_1325);
nor U2344 (N_2344,In_2726,In_2489);
nand U2345 (N_2345,In_2536,In_2773);
nor U2346 (N_2346,In_972,In_1122);
and U2347 (N_2347,In_274,In_2789);
and U2348 (N_2348,In_1132,In_693);
and U2349 (N_2349,In_968,In_1519);
or U2350 (N_2350,In_2280,In_2934);
xor U2351 (N_2351,In_973,In_1839);
and U2352 (N_2352,In_110,In_894);
and U2353 (N_2353,In_1297,In_274);
or U2354 (N_2354,In_147,In_1932);
and U2355 (N_2355,In_3,In_2253);
xnor U2356 (N_2356,In_341,In_349);
or U2357 (N_2357,In_2175,In_2082);
nand U2358 (N_2358,In_646,In_2897);
and U2359 (N_2359,In_1523,In_1701);
nor U2360 (N_2360,In_2878,In_705);
nor U2361 (N_2361,In_300,In_2314);
nor U2362 (N_2362,In_42,In_2957);
and U2363 (N_2363,In_1285,In_2353);
and U2364 (N_2364,In_2383,In_1869);
nand U2365 (N_2365,In_328,In_1248);
and U2366 (N_2366,In_2770,In_1507);
xor U2367 (N_2367,In_2481,In_1661);
xnor U2368 (N_2368,In_743,In_1459);
or U2369 (N_2369,In_973,In_579);
nand U2370 (N_2370,In_1712,In_2159);
nor U2371 (N_2371,In_2076,In_1600);
nor U2372 (N_2372,In_1728,In_552);
nor U2373 (N_2373,In_634,In_843);
or U2374 (N_2374,In_2318,In_339);
nor U2375 (N_2375,In_1314,In_2955);
and U2376 (N_2376,In_2683,In_59);
or U2377 (N_2377,In_2197,In_1245);
and U2378 (N_2378,In_120,In_1807);
or U2379 (N_2379,In_2707,In_463);
nand U2380 (N_2380,In_1042,In_2516);
or U2381 (N_2381,In_2077,In_384);
or U2382 (N_2382,In_1560,In_1563);
nand U2383 (N_2383,In_943,In_2216);
nor U2384 (N_2384,In_586,In_814);
nand U2385 (N_2385,In_2412,In_1186);
and U2386 (N_2386,In_138,In_2562);
or U2387 (N_2387,In_910,In_698);
nor U2388 (N_2388,In_297,In_1671);
and U2389 (N_2389,In_612,In_1205);
nand U2390 (N_2390,In_2333,In_2229);
or U2391 (N_2391,In_367,In_1307);
nor U2392 (N_2392,In_572,In_1483);
or U2393 (N_2393,In_2671,In_1471);
nor U2394 (N_2394,In_416,In_1094);
nor U2395 (N_2395,In_2015,In_454);
nand U2396 (N_2396,In_1573,In_227);
nand U2397 (N_2397,In_914,In_2673);
nand U2398 (N_2398,In_1857,In_1716);
or U2399 (N_2399,In_1901,In_2849);
nand U2400 (N_2400,In_55,In_2173);
and U2401 (N_2401,In_2592,In_79);
nand U2402 (N_2402,In_2024,In_1362);
nand U2403 (N_2403,In_2720,In_424);
nor U2404 (N_2404,In_2683,In_163);
nand U2405 (N_2405,In_879,In_1240);
and U2406 (N_2406,In_2931,In_1784);
and U2407 (N_2407,In_2968,In_2250);
or U2408 (N_2408,In_2104,In_2723);
or U2409 (N_2409,In_628,In_2833);
nor U2410 (N_2410,In_2110,In_775);
or U2411 (N_2411,In_1091,In_417);
nand U2412 (N_2412,In_596,In_2307);
and U2413 (N_2413,In_1171,In_2796);
or U2414 (N_2414,In_1540,In_1507);
and U2415 (N_2415,In_826,In_1217);
nand U2416 (N_2416,In_1739,In_629);
nand U2417 (N_2417,In_2163,In_2833);
xnor U2418 (N_2418,In_419,In_58);
or U2419 (N_2419,In_1165,In_984);
nor U2420 (N_2420,In_2534,In_1983);
or U2421 (N_2421,In_1985,In_631);
nor U2422 (N_2422,In_959,In_336);
nor U2423 (N_2423,In_1409,In_235);
nor U2424 (N_2424,In_2914,In_904);
nand U2425 (N_2425,In_612,In_2105);
nand U2426 (N_2426,In_265,In_131);
or U2427 (N_2427,In_2283,In_1281);
nand U2428 (N_2428,In_2331,In_1078);
or U2429 (N_2429,In_804,In_1676);
and U2430 (N_2430,In_2665,In_134);
nor U2431 (N_2431,In_1066,In_176);
nor U2432 (N_2432,In_604,In_1615);
or U2433 (N_2433,In_2664,In_1866);
or U2434 (N_2434,In_1593,In_1504);
nor U2435 (N_2435,In_2557,In_77);
xor U2436 (N_2436,In_519,In_2181);
nor U2437 (N_2437,In_2557,In_29);
nor U2438 (N_2438,In_1489,In_586);
and U2439 (N_2439,In_2982,In_2487);
nand U2440 (N_2440,In_2054,In_1298);
and U2441 (N_2441,In_2224,In_614);
nor U2442 (N_2442,In_1597,In_490);
and U2443 (N_2443,In_2489,In_1037);
xnor U2444 (N_2444,In_2407,In_2657);
xnor U2445 (N_2445,In_857,In_582);
nor U2446 (N_2446,In_1656,In_2036);
xnor U2447 (N_2447,In_454,In_996);
and U2448 (N_2448,In_1755,In_2842);
or U2449 (N_2449,In_2969,In_2056);
nor U2450 (N_2450,In_833,In_964);
or U2451 (N_2451,In_2384,In_127);
nor U2452 (N_2452,In_1647,In_895);
and U2453 (N_2453,In_1910,In_2782);
nor U2454 (N_2454,In_65,In_2436);
nor U2455 (N_2455,In_1155,In_971);
nand U2456 (N_2456,In_2957,In_1335);
or U2457 (N_2457,In_1765,In_1734);
nor U2458 (N_2458,In_1599,In_214);
or U2459 (N_2459,In_274,In_183);
nand U2460 (N_2460,In_2248,In_2843);
xor U2461 (N_2461,In_686,In_6);
nor U2462 (N_2462,In_257,In_426);
nand U2463 (N_2463,In_2163,In_875);
nor U2464 (N_2464,In_650,In_647);
xor U2465 (N_2465,In_1233,In_400);
nand U2466 (N_2466,In_470,In_2891);
nand U2467 (N_2467,In_2547,In_625);
nor U2468 (N_2468,In_1620,In_218);
nor U2469 (N_2469,In_1392,In_2377);
xor U2470 (N_2470,In_205,In_1959);
nand U2471 (N_2471,In_588,In_1577);
and U2472 (N_2472,In_513,In_2580);
and U2473 (N_2473,In_2427,In_1429);
and U2474 (N_2474,In_2671,In_852);
nand U2475 (N_2475,In_1985,In_75);
nand U2476 (N_2476,In_1800,In_1270);
or U2477 (N_2477,In_211,In_2266);
nand U2478 (N_2478,In_86,In_1498);
nor U2479 (N_2479,In_1443,In_2786);
nor U2480 (N_2480,In_549,In_2471);
nor U2481 (N_2481,In_1496,In_1342);
or U2482 (N_2482,In_653,In_1399);
nor U2483 (N_2483,In_258,In_1362);
nor U2484 (N_2484,In_392,In_798);
nor U2485 (N_2485,In_166,In_1129);
or U2486 (N_2486,In_1625,In_743);
or U2487 (N_2487,In_334,In_2764);
nand U2488 (N_2488,In_37,In_1996);
nor U2489 (N_2489,In_1467,In_2944);
and U2490 (N_2490,In_2761,In_717);
or U2491 (N_2491,In_144,In_600);
nor U2492 (N_2492,In_710,In_929);
or U2493 (N_2493,In_1049,In_371);
or U2494 (N_2494,In_99,In_796);
nand U2495 (N_2495,In_2722,In_398);
xor U2496 (N_2496,In_1850,In_1374);
or U2497 (N_2497,In_965,In_2257);
or U2498 (N_2498,In_2441,In_601);
and U2499 (N_2499,In_927,In_876);
nor U2500 (N_2500,In_1111,In_1073);
and U2501 (N_2501,In_336,In_1703);
and U2502 (N_2502,In_1209,In_1709);
or U2503 (N_2503,In_1065,In_2488);
nor U2504 (N_2504,In_2114,In_1841);
nand U2505 (N_2505,In_440,In_2924);
nand U2506 (N_2506,In_1283,In_364);
or U2507 (N_2507,In_2056,In_1878);
nor U2508 (N_2508,In_145,In_898);
or U2509 (N_2509,In_69,In_1185);
nor U2510 (N_2510,In_1866,In_2558);
nand U2511 (N_2511,In_1183,In_2260);
nand U2512 (N_2512,In_723,In_160);
and U2513 (N_2513,In_1312,In_2592);
nand U2514 (N_2514,In_1009,In_1051);
xor U2515 (N_2515,In_988,In_5);
nor U2516 (N_2516,In_2732,In_2181);
and U2517 (N_2517,In_677,In_77);
nor U2518 (N_2518,In_1621,In_948);
or U2519 (N_2519,In_2955,In_13);
nand U2520 (N_2520,In_1639,In_1469);
and U2521 (N_2521,In_1630,In_905);
or U2522 (N_2522,In_1340,In_2368);
and U2523 (N_2523,In_1653,In_2670);
or U2524 (N_2524,In_1708,In_2468);
nor U2525 (N_2525,In_1346,In_1101);
nor U2526 (N_2526,In_324,In_1537);
nand U2527 (N_2527,In_831,In_186);
nand U2528 (N_2528,In_1158,In_2001);
nand U2529 (N_2529,In_176,In_1138);
and U2530 (N_2530,In_870,In_1986);
xnor U2531 (N_2531,In_2458,In_2010);
and U2532 (N_2532,In_2245,In_2814);
nor U2533 (N_2533,In_2102,In_2948);
nor U2534 (N_2534,In_1873,In_1335);
or U2535 (N_2535,In_1664,In_1901);
nor U2536 (N_2536,In_2556,In_1624);
and U2537 (N_2537,In_320,In_2734);
nand U2538 (N_2538,In_1446,In_2730);
or U2539 (N_2539,In_1881,In_380);
nor U2540 (N_2540,In_2168,In_2003);
and U2541 (N_2541,In_2118,In_2952);
nand U2542 (N_2542,In_632,In_1742);
nor U2543 (N_2543,In_1674,In_2697);
nor U2544 (N_2544,In_161,In_244);
and U2545 (N_2545,In_315,In_1378);
or U2546 (N_2546,In_532,In_2626);
nor U2547 (N_2547,In_2501,In_2562);
or U2548 (N_2548,In_2083,In_2066);
nand U2549 (N_2549,In_771,In_2636);
or U2550 (N_2550,In_822,In_2328);
or U2551 (N_2551,In_2496,In_1594);
nor U2552 (N_2552,In_1374,In_753);
nand U2553 (N_2553,In_1376,In_1403);
nor U2554 (N_2554,In_2069,In_2492);
nor U2555 (N_2555,In_2975,In_296);
nand U2556 (N_2556,In_205,In_1195);
nand U2557 (N_2557,In_2439,In_1731);
nor U2558 (N_2558,In_371,In_2534);
xnor U2559 (N_2559,In_1390,In_98);
nand U2560 (N_2560,In_1940,In_234);
nor U2561 (N_2561,In_904,In_1013);
nand U2562 (N_2562,In_1963,In_1833);
nand U2563 (N_2563,In_924,In_2258);
or U2564 (N_2564,In_2919,In_1490);
xnor U2565 (N_2565,In_2298,In_1330);
and U2566 (N_2566,In_165,In_791);
xor U2567 (N_2567,In_1504,In_1728);
and U2568 (N_2568,In_2968,In_777);
nor U2569 (N_2569,In_968,In_1879);
or U2570 (N_2570,In_492,In_493);
or U2571 (N_2571,In_2496,In_1362);
and U2572 (N_2572,In_93,In_2608);
and U2573 (N_2573,In_1981,In_1943);
and U2574 (N_2574,In_2658,In_580);
nand U2575 (N_2575,In_2240,In_2420);
or U2576 (N_2576,In_1908,In_2361);
xor U2577 (N_2577,In_1214,In_523);
nor U2578 (N_2578,In_2730,In_680);
nor U2579 (N_2579,In_1649,In_1305);
nand U2580 (N_2580,In_1926,In_2995);
and U2581 (N_2581,In_1726,In_2124);
nor U2582 (N_2582,In_2450,In_2752);
and U2583 (N_2583,In_111,In_2378);
nand U2584 (N_2584,In_111,In_794);
nand U2585 (N_2585,In_2298,In_700);
nor U2586 (N_2586,In_2001,In_1075);
nor U2587 (N_2587,In_2681,In_370);
nand U2588 (N_2588,In_2090,In_2354);
and U2589 (N_2589,In_2440,In_2245);
or U2590 (N_2590,In_2603,In_2178);
and U2591 (N_2591,In_1659,In_2753);
nor U2592 (N_2592,In_1226,In_2406);
nor U2593 (N_2593,In_710,In_1881);
nor U2594 (N_2594,In_2527,In_1971);
or U2595 (N_2595,In_1956,In_1801);
or U2596 (N_2596,In_1061,In_1529);
and U2597 (N_2597,In_2594,In_1562);
nor U2598 (N_2598,In_2676,In_2700);
xnor U2599 (N_2599,In_1798,In_2216);
and U2600 (N_2600,In_684,In_1868);
nor U2601 (N_2601,In_164,In_804);
or U2602 (N_2602,In_148,In_2903);
or U2603 (N_2603,In_2341,In_1008);
nor U2604 (N_2604,In_935,In_381);
nor U2605 (N_2605,In_791,In_2201);
nor U2606 (N_2606,In_969,In_2952);
nor U2607 (N_2607,In_1262,In_2209);
nor U2608 (N_2608,In_1273,In_2303);
nor U2609 (N_2609,In_1413,In_97);
or U2610 (N_2610,In_486,In_1148);
and U2611 (N_2611,In_2231,In_520);
nand U2612 (N_2612,In_1369,In_1005);
nand U2613 (N_2613,In_130,In_948);
nand U2614 (N_2614,In_2111,In_1076);
or U2615 (N_2615,In_1519,In_1976);
nor U2616 (N_2616,In_1625,In_393);
and U2617 (N_2617,In_2934,In_1922);
or U2618 (N_2618,In_2245,In_2655);
nand U2619 (N_2619,In_789,In_1366);
or U2620 (N_2620,In_562,In_805);
nor U2621 (N_2621,In_1375,In_1833);
and U2622 (N_2622,In_752,In_346);
nand U2623 (N_2623,In_2462,In_1370);
xnor U2624 (N_2624,In_1675,In_416);
and U2625 (N_2625,In_1409,In_2797);
or U2626 (N_2626,In_2464,In_1372);
nor U2627 (N_2627,In_99,In_2835);
and U2628 (N_2628,In_968,In_119);
and U2629 (N_2629,In_2082,In_1973);
or U2630 (N_2630,In_2321,In_2234);
nand U2631 (N_2631,In_1812,In_1623);
or U2632 (N_2632,In_2791,In_2998);
nand U2633 (N_2633,In_219,In_2577);
and U2634 (N_2634,In_467,In_1344);
nand U2635 (N_2635,In_1285,In_411);
nand U2636 (N_2636,In_983,In_803);
or U2637 (N_2637,In_2938,In_2089);
or U2638 (N_2638,In_727,In_2474);
nor U2639 (N_2639,In_2100,In_30);
nand U2640 (N_2640,In_2656,In_1009);
and U2641 (N_2641,In_1688,In_2115);
or U2642 (N_2642,In_615,In_1220);
or U2643 (N_2643,In_2583,In_371);
nand U2644 (N_2644,In_2014,In_1520);
and U2645 (N_2645,In_2828,In_1234);
or U2646 (N_2646,In_1059,In_2635);
nand U2647 (N_2647,In_2172,In_1276);
nor U2648 (N_2648,In_66,In_2994);
or U2649 (N_2649,In_794,In_156);
nand U2650 (N_2650,In_2793,In_64);
xnor U2651 (N_2651,In_1215,In_2883);
and U2652 (N_2652,In_2745,In_1113);
and U2653 (N_2653,In_2038,In_328);
nand U2654 (N_2654,In_763,In_400);
and U2655 (N_2655,In_328,In_1712);
and U2656 (N_2656,In_2909,In_1655);
and U2657 (N_2657,In_2542,In_311);
or U2658 (N_2658,In_1902,In_1678);
nand U2659 (N_2659,In_2806,In_188);
nand U2660 (N_2660,In_1581,In_2541);
or U2661 (N_2661,In_158,In_1994);
nand U2662 (N_2662,In_29,In_2233);
or U2663 (N_2663,In_1844,In_2038);
or U2664 (N_2664,In_2790,In_521);
nor U2665 (N_2665,In_2877,In_441);
xnor U2666 (N_2666,In_2391,In_93);
xor U2667 (N_2667,In_2071,In_1415);
or U2668 (N_2668,In_302,In_749);
and U2669 (N_2669,In_1917,In_2891);
nand U2670 (N_2670,In_1059,In_2684);
nor U2671 (N_2671,In_365,In_620);
nand U2672 (N_2672,In_2338,In_2874);
or U2673 (N_2673,In_1429,In_222);
and U2674 (N_2674,In_2772,In_2357);
and U2675 (N_2675,In_2990,In_775);
nand U2676 (N_2676,In_29,In_2473);
nand U2677 (N_2677,In_2737,In_1979);
nand U2678 (N_2678,In_81,In_2531);
and U2679 (N_2679,In_1673,In_552);
or U2680 (N_2680,In_93,In_2417);
nand U2681 (N_2681,In_2822,In_1679);
xor U2682 (N_2682,In_50,In_1080);
nor U2683 (N_2683,In_2476,In_1776);
nor U2684 (N_2684,In_1707,In_358);
and U2685 (N_2685,In_427,In_1150);
xnor U2686 (N_2686,In_723,In_981);
nand U2687 (N_2687,In_846,In_2535);
or U2688 (N_2688,In_754,In_1694);
and U2689 (N_2689,In_2355,In_1593);
nand U2690 (N_2690,In_1299,In_2778);
and U2691 (N_2691,In_1431,In_538);
or U2692 (N_2692,In_1424,In_2111);
xor U2693 (N_2693,In_1019,In_2394);
and U2694 (N_2694,In_540,In_2869);
nand U2695 (N_2695,In_1995,In_2952);
or U2696 (N_2696,In_2193,In_1353);
or U2697 (N_2697,In_1251,In_2960);
and U2698 (N_2698,In_2988,In_345);
and U2699 (N_2699,In_260,In_2286);
and U2700 (N_2700,In_860,In_59);
or U2701 (N_2701,In_1176,In_989);
nand U2702 (N_2702,In_1131,In_424);
nor U2703 (N_2703,In_322,In_1099);
or U2704 (N_2704,In_93,In_2460);
nand U2705 (N_2705,In_2933,In_2012);
xor U2706 (N_2706,In_776,In_366);
or U2707 (N_2707,In_1744,In_445);
nand U2708 (N_2708,In_1633,In_2827);
nor U2709 (N_2709,In_1971,In_1784);
or U2710 (N_2710,In_1739,In_2817);
nand U2711 (N_2711,In_1920,In_1307);
or U2712 (N_2712,In_1362,In_222);
nor U2713 (N_2713,In_1126,In_1726);
nor U2714 (N_2714,In_1585,In_425);
and U2715 (N_2715,In_1445,In_2605);
nor U2716 (N_2716,In_1590,In_1840);
nand U2717 (N_2717,In_2766,In_2777);
and U2718 (N_2718,In_2963,In_2140);
and U2719 (N_2719,In_962,In_1219);
nand U2720 (N_2720,In_1886,In_1636);
nand U2721 (N_2721,In_1191,In_1405);
nor U2722 (N_2722,In_992,In_863);
or U2723 (N_2723,In_962,In_723);
or U2724 (N_2724,In_2653,In_664);
nand U2725 (N_2725,In_846,In_2398);
or U2726 (N_2726,In_975,In_2420);
nand U2727 (N_2727,In_779,In_984);
xnor U2728 (N_2728,In_407,In_2138);
or U2729 (N_2729,In_1554,In_1689);
nand U2730 (N_2730,In_1824,In_2395);
and U2731 (N_2731,In_2124,In_1705);
nor U2732 (N_2732,In_2588,In_2277);
and U2733 (N_2733,In_2832,In_1802);
nand U2734 (N_2734,In_350,In_34);
nor U2735 (N_2735,In_2155,In_2830);
nand U2736 (N_2736,In_2374,In_2191);
nor U2737 (N_2737,In_2930,In_2057);
nand U2738 (N_2738,In_1134,In_1532);
nand U2739 (N_2739,In_1320,In_2938);
xor U2740 (N_2740,In_333,In_2679);
xnor U2741 (N_2741,In_2784,In_619);
xnor U2742 (N_2742,In_2559,In_2037);
nor U2743 (N_2743,In_2997,In_502);
nand U2744 (N_2744,In_2843,In_393);
nor U2745 (N_2745,In_484,In_2114);
and U2746 (N_2746,In_1289,In_2153);
nand U2747 (N_2747,In_173,In_991);
or U2748 (N_2748,In_1446,In_2328);
nand U2749 (N_2749,In_2246,In_2738);
and U2750 (N_2750,In_1479,In_1995);
nor U2751 (N_2751,In_2764,In_908);
nand U2752 (N_2752,In_276,In_2652);
nor U2753 (N_2753,In_186,In_1740);
or U2754 (N_2754,In_690,In_852);
or U2755 (N_2755,In_557,In_156);
xnor U2756 (N_2756,In_1911,In_939);
nand U2757 (N_2757,In_14,In_2518);
xor U2758 (N_2758,In_778,In_1633);
and U2759 (N_2759,In_2442,In_2891);
nor U2760 (N_2760,In_1237,In_2099);
nand U2761 (N_2761,In_467,In_619);
and U2762 (N_2762,In_1655,In_2770);
nand U2763 (N_2763,In_1694,In_20);
or U2764 (N_2764,In_2807,In_2310);
and U2765 (N_2765,In_1773,In_1415);
and U2766 (N_2766,In_1961,In_993);
or U2767 (N_2767,In_381,In_2637);
nor U2768 (N_2768,In_845,In_667);
and U2769 (N_2769,In_2284,In_1587);
or U2770 (N_2770,In_989,In_456);
nand U2771 (N_2771,In_1943,In_1666);
nor U2772 (N_2772,In_2657,In_931);
and U2773 (N_2773,In_2909,In_1035);
nor U2774 (N_2774,In_828,In_887);
or U2775 (N_2775,In_2957,In_1908);
or U2776 (N_2776,In_2083,In_1549);
nor U2777 (N_2777,In_79,In_980);
and U2778 (N_2778,In_1711,In_2444);
and U2779 (N_2779,In_592,In_2215);
and U2780 (N_2780,In_1504,In_2462);
or U2781 (N_2781,In_1161,In_369);
and U2782 (N_2782,In_955,In_334);
or U2783 (N_2783,In_725,In_477);
nor U2784 (N_2784,In_1634,In_659);
or U2785 (N_2785,In_1139,In_389);
or U2786 (N_2786,In_1486,In_194);
nand U2787 (N_2787,In_701,In_2603);
and U2788 (N_2788,In_1864,In_134);
and U2789 (N_2789,In_1725,In_1344);
or U2790 (N_2790,In_1818,In_2762);
and U2791 (N_2791,In_885,In_258);
xnor U2792 (N_2792,In_759,In_236);
nor U2793 (N_2793,In_2251,In_2721);
nand U2794 (N_2794,In_1964,In_1921);
and U2795 (N_2795,In_644,In_1383);
or U2796 (N_2796,In_732,In_2876);
and U2797 (N_2797,In_2204,In_197);
and U2798 (N_2798,In_2203,In_2184);
or U2799 (N_2799,In_686,In_2214);
or U2800 (N_2800,In_441,In_1260);
nor U2801 (N_2801,In_2331,In_2716);
nor U2802 (N_2802,In_562,In_532);
or U2803 (N_2803,In_1055,In_1429);
nor U2804 (N_2804,In_2218,In_1033);
nor U2805 (N_2805,In_577,In_2788);
xor U2806 (N_2806,In_566,In_1133);
and U2807 (N_2807,In_1114,In_2895);
and U2808 (N_2808,In_2843,In_2194);
nor U2809 (N_2809,In_1887,In_384);
nor U2810 (N_2810,In_1523,In_2532);
xnor U2811 (N_2811,In_2157,In_2619);
and U2812 (N_2812,In_112,In_1925);
nor U2813 (N_2813,In_984,In_1161);
nor U2814 (N_2814,In_2561,In_1750);
nor U2815 (N_2815,In_2529,In_1488);
or U2816 (N_2816,In_1074,In_2750);
or U2817 (N_2817,In_263,In_2387);
nor U2818 (N_2818,In_1214,In_505);
nand U2819 (N_2819,In_2376,In_1097);
or U2820 (N_2820,In_1274,In_2534);
xnor U2821 (N_2821,In_134,In_1259);
nand U2822 (N_2822,In_2737,In_1609);
or U2823 (N_2823,In_2667,In_748);
and U2824 (N_2824,In_1702,In_2109);
nor U2825 (N_2825,In_2159,In_358);
and U2826 (N_2826,In_2330,In_1857);
or U2827 (N_2827,In_1655,In_654);
and U2828 (N_2828,In_299,In_1308);
xnor U2829 (N_2829,In_2345,In_2623);
nand U2830 (N_2830,In_1604,In_2824);
and U2831 (N_2831,In_1943,In_1299);
or U2832 (N_2832,In_1986,In_787);
or U2833 (N_2833,In_226,In_641);
nor U2834 (N_2834,In_1596,In_1416);
and U2835 (N_2835,In_1264,In_2175);
nand U2836 (N_2836,In_1463,In_986);
nor U2837 (N_2837,In_1643,In_1554);
and U2838 (N_2838,In_2091,In_1190);
or U2839 (N_2839,In_797,In_2257);
nor U2840 (N_2840,In_2719,In_2468);
or U2841 (N_2841,In_1947,In_1714);
nor U2842 (N_2842,In_2423,In_776);
and U2843 (N_2843,In_315,In_2458);
nand U2844 (N_2844,In_1739,In_795);
nand U2845 (N_2845,In_319,In_2166);
nor U2846 (N_2846,In_779,In_666);
and U2847 (N_2847,In_1417,In_1256);
xor U2848 (N_2848,In_1290,In_1);
or U2849 (N_2849,In_2185,In_1342);
xor U2850 (N_2850,In_539,In_1536);
nor U2851 (N_2851,In_263,In_318);
and U2852 (N_2852,In_1704,In_2850);
nand U2853 (N_2853,In_2421,In_1325);
nor U2854 (N_2854,In_208,In_2880);
nand U2855 (N_2855,In_1129,In_2033);
xnor U2856 (N_2856,In_764,In_2098);
or U2857 (N_2857,In_1949,In_2687);
or U2858 (N_2858,In_2435,In_107);
nor U2859 (N_2859,In_670,In_932);
nand U2860 (N_2860,In_330,In_510);
and U2861 (N_2861,In_1907,In_367);
or U2862 (N_2862,In_2171,In_196);
and U2863 (N_2863,In_2783,In_2352);
or U2864 (N_2864,In_2186,In_2637);
nand U2865 (N_2865,In_1201,In_351);
xnor U2866 (N_2866,In_78,In_307);
nand U2867 (N_2867,In_1849,In_797);
or U2868 (N_2868,In_1643,In_1904);
and U2869 (N_2869,In_1142,In_325);
xnor U2870 (N_2870,In_616,In_596);
or U2871 (N_2871,In_267,In_953);
or U2872 (N_2872,In_2934,In_224);
or U2873 (N_2873,In_13,In_2187);
or U2874 (N_2874,In_2526,In_917);
and U2875 (N_2875,In_2440,In_2692);
xor U2876 (N_2876,In_2678,In_1744);
nand U2877 (N_2877,In_2837,In_849);
or U2878 (N_2878,In_2228,In_1955);
or U2879 (N_2879,In_1659,In_2565);
or U2880 (N_2880,In_1615,In_960);
nor U2881 (N_2881,In_1489,In_864);
nor U2882 (N_2882,In_82,In_1616);
and U2883 (N_2883,In_771,In_130);
or U2884 (N_2884,In_417,In_795);
or U2885 (N_2885,In_1509,In_1693);
nor U2886 (N_2886,In_2914,In_1382);
nor U2887 (N_2887,In_62,In_2850);
nor U2888 (N_2888,In_815,In_2724);
xnor U2889 (N_2889,In_2896,In_2476);
and U2890 (N_2890,In_159,In_2052);
nand U2891 (N_2891,In_1882,In_2457);
nand U2892 (N_2892,In_1515,In_613);
nor U2893 (N_2893,In_562,In_1363);
and U2894 (N_2894,In_2264,In_1627);
nor U2895 (N_2895,In_2415,In_1554);
or U2896 (N_2896,In_2283,In_1263);
nor U2897 (N_2897,In_831,In_2433);
nor U2898 (N_2898,In_1464,In_1605);
or U2899 (N_2899,In_447,In_1861);
or U2900 (N_2900,In_954,In_2332);
and U2901 (N_2901,In_827,In_144);
nand U2902 (N_2902,In_2934,In_860);
nor U2903 (N_2903,In_2404,In_453);
nor U2904 (N_2904,In_757,In_899);
or U2905 (N_2905,In_2337,In_858);
nor U2906 (N_2906,In_97,In_954);
or U2907 (N_2907,In_2702,In_1718);
or U2908 (N_2908,In_1713,In_933);
or U2909 (N_2909,In_1060,In_2373);
xor U2910 (N_2910,In_564,In_1528);
or U2911 (N_2911,In_1665,In_1955);
nor U2912 (N_2912,In_1968,In_1980);
nor U2913 (N_2913,In_1839,In_1505);
nand U2914 (N_2914,In_524,In_1758);
and U2915 (N_2915,In_2364,In_220);
or U2916 (N_2916,In_2324,In_1440);
nor U2917 (N_2917,In_1937,In_2973);
or U2918 (N_2918,In_2086,In_1758);
xor U2919 (N_2919,In_460,In_1462);
or U2920 (N_2920,In_420,In_2558);
nor U2921 (N_2921,In_1606,In_2133);
or U2922 (N_2922,In_2089,In_47);
nand U2923 (N_2923,In_36,In_1158);
nor U2924 (N_2924,In_2211,In_1557);
nand U2925 (N_2925,In_2185,In_1048);
nor U2926 (N_2926,In_2655,In_1316);
nand U2927 (N_2927,In_2674,In_2021);
or U2928 (N_2928,In_2599,In_1596);
nand U2929 (N_2929,In_2273,In_2349);
and U2930 (N_2930,In_2850,In_1034);
and U2931 (N_2931,In_2376,In_541);
or U2932 (N_2932,In_2766,In_2929);
or U2933 (N_2933,In_184,In_25);
and U2934 (N_2934,In_2287,In_1134);
xor U2935 (N_2935,In_2739,In_2854);
or U2936 (N_2936,In_6,In_906);
or U2937 (N_2937,In_2635,In_2818);
or U2938 (N_2938,In_1998,In_2238);
nor U2939 (N_2939,In_2391,In_466);
nand U2940 (N_2940,In_2319,In_1759);
and U2941 (N_2941,In_838,In_2554);
and U2942 (N_2942,In_1459,In_1599);
xnor U2943 (N_2943,In_2510,In_556);
xor U2944 (N_2944,In_372,In_357);
and U2945 (N_2945,In_1273,In_2266);
nor U2946 (N_2946,In_2998,In_2594);
or U2947 (N_2947,In_723,In_2016);
and U2948 (N_2948,In_1842,In_2254);
xnor U2949 (N_2949,In_361,In_2774);
or U2950 (N_2950,In_838,In_1515);
nand U2951 (N_2951,In_2160,In_844);
and U2952 (N_2952,In_2422,In_2342);
nand U2953 (N_2953,In_2000,In_361);
nand U2954 (N_2954,In_1986,In_370);
and U2955 (N_2955,In_1300,In_1051);
xor U2956 (N_2956,In_2163,In_1754);
nor U2957 (N_2957,In_551,In_2086);
nor U2958 (N_2958,In_2365,In_1930);
xor U2959 (N_2959,In_1892,In_1298);
or U2960 (N_2960,In_204,In_2965);
nand U2961 (N_2961,In_2033,In_443);
and U2962 (N_2962,In_2491,In_2917);
nand U2963 (N_2963,In_984,In_995);
xor U2964 (N_2964,In_565,In_1360);
nand U2965 (N_2965,In_1213,In_2438);
nand U2966 (N_2966,In_946,In_2473);
or U2967 (N_2967,In_1844,In_1838);
xor U2968 (N_2968,In_2286,In_1464);
nor U2969 (N_2969,In_1663,In_947);
nor U2970 (N_2970,In_2932,In_544);
nor U2971 (N_2971,In_1195,In_678);
or U2972 (N_2972,In_239,In_1204);
and U2973 (N_2973,In_2662,In_2304);
and U2974 (N_2974,In_1086,In_2720);
or U2975 (N_2975,In_2887,In_2217);
nand U2976 (N_2976,In_408,In_2077);
nand U2977 (N_2977,In_104,In_1092);
or U2978 (N_2978,In_1451,In_1928);
nor U2979 (N_2979,In_1336,In_2847);
or U2980 (N_2980,In_1255,In_2892);
nor U2981 (N_2981,In_2192,In_423);
nand U2982 (N_2982,In_2447,In_1594);
nor U2983 (N_2983,In_2219,In_908);
or U2984 (N_2984,In_1695,In_419);
or U2985 (N_2985,In_2946,In_330);
nor U2986 (N_2986,In_342,In_1921);
and U2987 (N_2987,In_624,In_1317);
nor U2988 (N_2988,In_2831,In_1523);
nand U2989 (N_2989,In_1519,In_1631);
nand U2990 (N_2990,In_682,In_1561);
and U2991 (N_2991,In_1316,In_352);
xnor U2992 (N_2992,In_2132,In_2595);
nor U2993 (N_2993,In_2497,In_1700);
nor U2994 (N_2994,In_572,In_346);
nor U2995 (N_2995,In_949,In_2057);
and U2996 (N_2996,In_1423,In_1110);
or U2997 (N_2997,In_116,In_57);
and U2998 (N_2998,In_2521,In_971);
nand U2999 (N_2999,In_2155,In_1471);
and U3000 (N_3000,In_2713,In_103);
nand U3001 (N_3001,In_1127,In_1437);
or U3002 (N_3002,In_207,In_2433);
nor U3003 (N_3003,In_1753,In_2457);
xnor U3004 (N_3004,In_1573,In_2060);
nor U3005 (N_3005,In_1513,In_766);
nand U3006 (N_3006,In_1315,In_90);
or U3007 (N_3007,In_2115,In_952);
nand U3008 (N_3008,In_720,In_341);
or U3009 (N_3009,In_976,In_2060);
nand U3010 (N_3010,In_1428,In_2724);
nand U3011 (N_3011,In_2914,In_680);
nor U3012 (N_3012,In_610,In_1072);
nor U3013 (N_3013,In_2705,In_1430);
nand U3014 (N_3014,In_2877,In_209);
nor U3015 (N_3015,In_1042,In_2190);
nand U3016 (N_3016,In_971,In_2182);
and U3017 (N_3017,In_36,In_2063);
nand U3018 (N_3018,In_2200,In_1551);
or U3019 (N_3019,In_1293,In_251);
or U3020 (N_3020,In_1663,In_241);
nand U3021 (N_3021,In_1513,In_2124);
nand U3022 (N_3022,In_2651,In_2378);
xor U3023 (N_3023,In_345,In_2557);
nor U3024 (N_3024,In_321,In_2984);
and U3025 (N_3025,In_551,In_453);
xor U3026 (N_3026,In_2144,In_2383);
nand U3027 (N_3027,In_1966,In_1977);
or U3028 (N_3028,In_416,In_1789);
nor U3029 (N_3029,In_1562,In_2801);
or U3030 (N_3030,In_948,In_1866);
nor U3031 (N_3031,In_802,In_819);
and U3032 (N_3032,In_1022,In_2290);
nand U3033 (N_3033,In_2244,In_2329);
and U3034 (N_3034,In_977,In_1576);
xnor U3035 (N_3035,In_2594,In_1114);
or U3036 (N_3036,In_1675,In_660);
and U3037 (N_3037,In_674,In_2192);
xor U3038 (N_3038,In_557,In_739);
and U3039 (N_3039,In_1857,In_47);
xor U3040 (N_3040,In_2544,In_2674);
nor U3041 (N_3041,In_107,In_1249);
and U3042 (N_3042,In_2518,In_1093);
or U3043 (N_3043,In_2125,In_782);
nand U3044 (N_3044,In_439,In_2823);
and U3045 (N_3045,In_1524,In_412);
and U3046 (N_3046,In_661,In_49);
nor U3047 (N_3047,In_1825,In_743);
and U3048 (N_3048,In_1533,In_1140);
and U3049 (N_3049,In_804,In_1346);
and U3050 (N_3050,In_2226,In_2022);
nor U3051 (N_3051,In_700,In_2780);
nand U3052 (N_3052,In_1761,In_771);
and U3053 (N_3053,In_2965,In_1012);
nand U3054 (N_3054,In_2606,In_854);
nor U3055 (N_3055,In_2696,In_1356);
nand U3056 (N_3056,In_451,In_2373);
or U3057 (N_3057,In_2045,In_2291);
nor U3058 (N_3058,In_1780,In_1808);
or U3059 (N_3059,In_1105,In_673);
nor U3060 (N_3060,In_26,In_573);
or U3061 (N_3061,In_359,In_1348);
and U3062 (N_3062,In_2130,In_186);
nor U3063 (N_3063,In_882,In_502);
nor U3064 (N_3064,In_1486,In_682);
and U3065 (N_3065,In_318,In_1381);
nor U3066 (N_3066,In_1578,In_1022);
and U3067 (N_3067,In_188,In_462);
or U3068 (N_3068,In_1653,In_1807);
nand U3069 (N_3069,In_2244,In_868);
xnor U3070 (N_3070,In_845,In_709);
nor U3071 (N_3071,In_2263,In_446);
or U3072 (N_3072,In_120,In_2217);
or U3073 (N_3073,In_920,In_2061);
nor U3074 (N_3074,In_2792,In_2371);
nor U3075 (N_3075,In_1644,In_1392);
xnor U3076 (N_3076,In_767,In_900);
nand U3077 (N_3077,In_2250,In_549);
nor U3078 (N_3078,In_1733,In_1722);
nor U3079 (N_3079,In_1372,In_1771);
or U3080 (N_3080,In_2997,In_2145);
nand U3081 (N_3081,In_181,In_455);
and U3082 (N_3082,In_1979,In_1056);
nand U3083 (N_3083,In_986,In_404);
and U3084 (N_3084,In_2257,In_1804);
and U3085 (N_3085,In_2032,In_1524);
and U3086 (N_3086,In_506,In_2689);
and U3087 (N_3087,In_1698,In_343);
nor U3088 (N_3088,In_176,In_2455);
nor U3089 (N_3089,In_1300,In_2865);
nor U3090 (N_3090,In_2254,In_226);
nor U3091 (N_3091,In_1436,In_781);
or U3092 (N_3092,In_697,In_93);
nand U3093 (N_3093,In_2555,In_780);
or U3094 (N_3094,In_2630,In_1517);
nand U3095 (N_3095,In_1063,In_851);
and U3096 (N_3096,In_442,In_930);
nor U3097 (N_3097,In_1961,In_835);
and U3098 (N_3098,In_1381,In_410);
xnor U3099 (N_3099,In_2614,In_526);
and U3100 (N_3100,In_436,In_352);
nand U3101 (N_3101,In_1353,In_2900);
and U3102 (N_3102,In_883,In_2294);
and U3103 (N_3103,In_1156,In_1142);
or U3104 (N_3104,In_612,In_1802);
or U3105 (N_3105,In_12,In_1508);
or U3106 (N_3106,In_2072,In_2176);
xnor U3107 (N_3107,In_327,In_2092);
or U3108 (N_3108,In_1288,In_182);
nor U3109 (N_3109,In_756,In_620);
nor U3110 (N_3110,In_2946,In_880);
and U3111 (N_3111,In_1117,In_2202);
nand U3112 (N_3112,In_2861,In_145);
or U3113 (N_3113,In_2679,In_2593);
or U3114 (N_3114,In_1891,In_527);
xor U3115 (N_3115,In_1054,In_1777);
or U3116 (N_3116,In_2486,In_301);
or U3117 (N_3117,In_2888,In_506);
nor U3118 (N_3118,In_642,In_2442);
and U3119 (N_3119,In_329,In_2962);
xnor U3120 (N_3120,In_2818,In_666);
nor U3121 (N_3121,In_439,In_287);
and U3122 (N_3122,In_2410,In_2487);
and U3123 (N_3123,In_2431,In_2523);
xor U3124 (N_3124,In_2374,In_2623);
or U3125 (N_3125,In_682,In_710);
and U3126 (N_3126,In_1206,In_813);
and U3127 (N_3127,In_2869,In_115);
nor U3128 (N_3128,In_2145,In_903);
xor U3129 (N_3129,In_915,In_2854);
nor U3130 (N_3130,In_979,In_920);
nand U3131 (N_3131,In_122,In_1816);
nand U3132 (N_3132,In_1067,In_1689);
nand U3133 (N_3133,In_2082,In_2906);
nand U3134 (N_3134,In_201,In_1349);
and U3135 (N_3135,In_2935,In_1652);
or U3136 (N_3136,In_1887,In_61);
or U3137 (N_3137,In_523,In_1957);
nand U3138 (N_3138,In_2051,In_1264);
nand U3139 (N_3139,In_432,In_837);
and U3140 (N_3140,In_411,In_759);
and U3141 (N_3141,In_1423,In_2834);
and U3142 (N_3142,In_1383,In_2827);
and U3143 (N_3143,In_751,In_776);
xor U3144 (N_3144,In_1240,In_1283);
nand U3145 (N_3145,In_1890,In_417);
or U3146 (N_3146,In_215,In_48);
nand U3147 (N_3147,In_1840,In_2716);
or U3148 (N_3148,In_1693,In_2892);
and U3149 (N_3149,In_1725,In_2433);
and U3150 (N_3150,In_649,In_1599);
or U3151 (N_3151,In_1352,In_2829);
xnor U3152 (N_3152,In_1087,In_601);
nand U3153 (N_3153,In_2519,In_243);
and U3154 (N_3154,In_1397,In_1971);
or U3155 (N_3155,In_2315,In_957);
or U3156 (N_3156,In_1780,In_2638);
xnor U3157 (N_3157,In_286,In_1275);
nor U3158 (N_3158,In_2782,In_563);
or U3159 (N_3159,In_254,In_211);
nor U3160 (N_3160,In_2151,In_422);
nand U3161 (N_3161,In_1612,In_1205);
and U3162 (N_3162,In_2076,In_2914);
xor U3163 (N_3163,In_2580,In_1783);
nand U3164 (N_3164,In_255,In_2107);
xnor U3165 (N_3165,In_1183,In_1799);
nand U3166 (N_3166,In_952,In_1105);
xor U3167 (N_3167,In_1988,In_275);
and U3168 (N_3168,In_2113,In_1775);
nand U3169 (N_3169,In_2548,In_1545);
nand U3170 (N_3170,In_944,In_2515);
and U3171 (N_3171,In_647,In_2047);
or U3172 (N_3172,In_2997,In_102);
nand U3173 (N_3173,In_1256,In_1894);
nor U3174 (N_3174,In_2530,In_79);
and U3175 (N_3175,In_1267,In_1470);
and U3176 (N_3176,In_909,In_886);
or U3177 (N_3177,In_1819,In_144);
nor U3178 (N_3178,In_2782,In_2231);
or U3179 (N_3179,In_980,In_2322);
and U3180 (N_3180,In_2259,In_1182);
or U3181 (N_3181,In_160,In_2913);
or U3182 (N_3182,In_2296,In_403);
nand U3183 (N_3183,In_2108,In_119);
xnor U3184 (N_3184,In_1877,In_1115);
nand U3185 (N_3185,In_2932,In_1804);
and U3186 (N_3186,In_1576,In_2495);
nand U3187 (N_3187,In_1808,In_2004);
nor U3188 (N_3188,In_719,In_1416);
nor U3189 (N_3189,In_700,In_2741);
nand U3190 (N_3190,In_160,In_1764);
nand U3191 (N_3191,In_591,In_538);
nand U3192 (N_3192,In_1580,In_914);
or U3193 (N_3193,In_599,In_1270);
nand U3194 (N_3194,In_1459,In_311);
or U3195 (N_3195,In_1814,In_2224);
and U3196 (N_3196,In_1515,In_1035);
and U3197 (N_3197,In_978,In_2836);
and U3198 (N_3198,In_1574,In_1151);
and U3199 (N_3199,In_1033,In_2207);
or U3200 (N_3200,In_2513,In_985);
nand U3201 (N_3201,In_21,In_1371);
or U3202 (N_3202,In_2921,In_2122);
or U3203 (N_3203,In_1105,In_2732);
and U3204 (N_3204,In_1907,In_1631);
nor U3205 (N_3205,In_2987,In_2467);
nor U3206 (N_3206,In_78,In_821);
nand U3207 (N_3207,In_657,In_2060);
and U3208 (N_3208,In_928,In_2693);
nand U3209 (N_3209,In_2436,In_1233);
nor U3210 (N_3210,In_95,In_1226);
nor U3211 (N_3211,In_218,In_564);
xnor U3212 (N_3212,In_2381,In_311);
nor U3213 (N_3213,In_1699,In_2013);
xor U3214 (N_3214,In_2055,In_2748);
xor U3215 (N_3215,In_1525,In_781);
and U3216 (N_3216,In_2425,In_1853);
nor U3217 (N_3217,In_724,In_2978);
or U3218 (N_3218,In_1260,In_1753);
and U3219 (N_3219,In_869,In_1026);
nand U3220 (N_3220,In_2334,In_2872);
or U3221 (N_3221,In_2381,In_1370);
or U3222 (N_3222,In_792,In_1953);
nand U3223 (N_3223,In_2535,In_2655);
nor U3224 (N_3224,In_1445,In_383);
nand U3225 (N_3225,In_372,In_328);
nor U3226 (N_3226,In_1988,In_767);
nor U3227 (N_3227,In_141,In_982);
and U3228 (N_3228,In_2250,In_695);
or U3229 (N_3229,In_1611,In_2842);
and U3230 (N_3230,In_2485,In_763);
or U3231 (N_3231,In_620,In_2663);
and U3232 (N_3232,In_2328,In_684);
or U3233 (N_3233,In_1941,In_2590);
nand U3234 (N_3234,In_744,In_1341);
or U3235 (N_3235,In_1274,In_1518);
nor U3236 (N_3236,In_986,In_1610);
nand U3237 (N_3237,In_2505,In_2934);
or U3238 (N_3238,In_2874,In_405);
nor U3239 (N_3239,In_1172,In_212);
nand U3240 (N_3240,In_1530,In_1953);
xnor U3241 (N_3241,In_2612,In_109);
nand U3242 (N_3242,In_1663,In_2331);
nand U3243 (N_3243,In_2984,In_1931);
nor U3244 (N_3244,In_2360,In_593);
and U3245 (N_3245,In_2351,In_1578);
and U3246 (N_3246,In_1287,In_1145);
and U3247 (N_3247,In_2918,In_434);
xor U3248 (N_3248,In_591,In_988);
and U3249 (N_3249,In_2365,In_2636);
nand U3250 (N_3250,In_545,In_260);
nor U3251 (N_3251,In_2389,In_1708);
and U3252 (N_3252,In_2560,In_865);
xor U3253 (N_3253,In_1106,In_2466);
or U3254 (N_3254,In_1791,In_463);
or U3255 (N_3255,In_2773,In_2687);
nor U3256 (N_3256,In_2487,In_2049);
or U3257 (N_3257,In_1066,In_1676);
and U3258 (N_3258,In_2110,In_1139);
nand U3259 (N_3259,In_1407,In_458);
nand U3260 (N_3260,In_2554,In_1434);
and U3261 (N_3261,In_2707,In_1661);
xor U3262 (N_3262,In_2332,In_2128);
nand U3263 (N_3263,In_2238,In_1807);
and U3264 (N_3264,In_200,In_1051);
nand U3265 (N_3265,In_988,In_76);
nor U3266 (N_3266,In_1027,In_2577);
nand U3267 (N_3267,In_2605,In_1252);
nor U3268 (N_3268,In_1558,In_868);
and U3269 (N_3269,In_2424,In_2177);
nor U3270 (N_3270,In_2177,In_2751);
or U3271 (N_3271,In_2150,In_2278);
or U3272 (N_3272,In_504,In_109);
xnor U3273 (N_3273,In_642,In_2511);
nand U3274 (N_3274,In_1847,In_2774);
nor U3275 (N_3275,In_1227,In_1735);
or U3276 (N_3276,In_1845,In_2194);
nand U3277 (N_3277,In_2123,In_2628);
or U3278 (N_3278,In_2550,In_2511);
or U3279 (N_3279,In_2385,In_1348);
or U3280 (N_3280,In_229,In_1399);
nand U3281 (N_3281,In_2854,In_1230);
and U3282 (N_3282,In_1698,In_1012);
nand U3283 (N_3283,In_183,In_1062);
nand U3284 (N_3284,In_2073,In_1344);
xor U3285 (N_3285,In_1288,In_1693);
nand U3286 (N_3286,In_583,In_1475);
nor U3287 (N_3287,In_2348,In_935);
or U3288 (N_3288,In_730,In_2460);
nand U3289 (N_3289,In_2695,In_766);
xnor U3290 (N_3290,In_1520,In_2472);
nand U3291 (N_3291,In_2876,In_2725);
xnor U3292 (N_3292,In_969,In_2791);
or U3293 (N_3293,In_2399,In_2085);
and U3294 (N_3294,In_989,In_2734);
and U3295 (N_3295,In_2572,In_2590);
or U3296 (N_3296,In_1778,In_2080);
or U3297 (N_3297,In_2038,In_1984);
or U3298 (N_3298,In_2473,In_16);
or U3299 (N_3299,In_2223,In_1651);
nand U3300 (N_3300,In_372,In_2102);
nand U3301 (N_3301,In_2891,In_359);
or U3302 (N_3302,In_1600,In_920);
nor U3303 (N_3303,In_1521,In_1978);
nand U3304 (N_3304,In_2447,In_76);
nor U3305 (N_3305,In_2062,In_2183);
and U3306 (N_3306,In_514,In_2599);
nand U3307 (N_3307,In_2795,In_996);
nor U3308 (N_3308,In_572,In_539);
xnor U3309 (N_3309,In_1570,In_1216);
and U3310 (N_3310,In_37,In_2401);
xnor U3311 (N_3311,In_1994,In_807);
and U3312 (N_3312,In_2677,In_1917);
or U3313 (N_3313,In_626,In_2055);
xnor U3314 (N_3314,In_1835,In_911);
or U3315 (N_3315,In_2186,In_10);
nand U3316 (N_3316,In_670,In_2786);
xnor U3317 (N_3317,In_1836,In_1281);
nor U3318 (N_3318,In_2713,In_624);
nand U3319 (N_3319,In_513,In_2410);
or U3320 (N_3320,In_671,In_2578);
nand U3321 (N_3321,In_552,In_905);
nand U3322 (N_3322,In_842,In_1464);
or U3323 (N_3323,In_946,In_1064);
nor U3324 (N_3324,In_2494,In_2416);
and U3325 (N_3325,In_2212,In_1567);
and U3326 (N_3326,In_602,In_407);
nor U3327 (N_3327,In_640,In_913);
or U3328 (N_3328,In_2086,In_1351);
nor U3329 (N_3329,In_749,In_2858);
and U3330 (N_3330,In_1891,In_2337);
and U3331 (N_3331,In_1,In_2712);
nor U3332 (N_3332,In_2428,In_215);
and U3333 (N_3333,In_2696,In_1937);
or U3334 (N_3334,In_2534,In_1079);
or U3335 (N_3335,In_1709,In_2998);
nor U3336 (N_3336,In_2567,In_2091);
nor U3337 (N_3337,In_554,In_1367);
and U3338 (N_3338,In_45,In_753);
and U3339 (N_3339,In_495,In_2688);
and U3340 (N_3340,In_1783,In_1842);
nand U3341 (N_3341,In_1946,In_2759);
or U3342 (N_3342,In_2211,In_957);
nor U3343 (N_3343,In_85,In_1747);
and U3344 (N_3344,In_1528,In_2129);
nor U3345 (N_3345,In_2173,In_2763);
nand U3346 (N_3346,In_1368,In_925);
nor U3347 (N_3347,In_59,In_693);
nor U3348 (N_3348,In_1034,In_2165);
and U3349 (N_3349,In_202,In_1311);
nand U3350 (N_3350,In_1032,In_424);
and U3351 (N_3351,In_1165,In_1433);
or U3352 (N_3352,In_2485,In_760);
nand U3353 (N_3353,In_781,In_636);
and U3354 (N_3354,In_1026,In_34);
and U3355 (N_3355,In_469,In_769);
nor U3356 (N_3356,In_2752,In_1631);
and U3357 (N_3357,In_15,In_553);
and U3358 (N_3358,In_2247,In_818);
and U3359 (N_3359,In_2254,In_1423);
nor U3360 (N_3360,In_241,In_749);
nor U3361 (N_3361,In_1220,In_116);
and U3362 (N_3362,In_746,In_1875);
nor U3363 (N_3363,In_1323,In_2424);
nor U3364 (N_3364,In_745,In_2878);
and U3365 (N_3365,In_2811,In_485);
or U3366 (N_3366,In_543,In_2406);
and U3367 (N_3367,In_1761,In_962);
nand U3368 (N_3368,In_2494,In_534);
nor U3369 (N_3369,In_1127,In_1489);
nor U3370 (N_3370,In_1247,In_2740);
and U3371 (N_3371,In_1642,In_2547);
and U3372 (N_3372,In_277,In_428);
and U3373 (N_3373,In_1778,In_1943);
and U3374 (N_3374,In_823,In_2563);
or U3375 (N_3375,In_279,In_91);
nand U3376 (N_3376,In_1351,In_1139);
nand U3377 (N_3377,In_2199,In_2200);
or U3378 (N_3378,In_1565,In_2116);
and U3379 (N_3379,In_2441,In_2717);
and U3380 (N_3380,In_2550,In_1604);
and U3381 (N_3381,In_355,In_2918);
or U3382 (N_3382,In_1472,In_2724);
or U3383 (N_3383,In_2999,In_2405);
nand U3384 (N_3384,In_552,In_70);
nand U3385 (N_3385,In_429,In_2551);
xnor U3386 (N_3386,In_165,In_159);
xor U3387 (N_3387,In_1270,In_1614);
nor U3388 (N_3388,In_654,In_1463);
xor U3389 (N_3389,In_1603,In_1298);
and U3390 (N_3390,In_2012,In_1948);
nor U3391 (N_3391,In_2608,In_1730);
nor U3392 (N_3392,In_1010,In_990);
nor U3393 (N_3393,In_226,In_744);
or U3394 (N_3394,In_1631,In_2931);
or U3395 (N_3395,In_229,In_1383);
or U3396 (N_3396,In_1134,In_2911);
nor U3397 (N_3397,In_2104,In_484);
nand U3398 (N_3398,In_1369,In_319);
nand U3399 (N_3399,In_2163,In_11);
and U3400 (N_3400,In_1816,In_887);
nor U3401 (N_3401,In_331,In_574);
nand U3402 (N_3402,In_552,In_771);
nand U3403 (N_3403,In_2324,In_1438);
nor U3404 (N_3404,In_1052,In_1861);
nand U3405 (N_3405,In_2438,In_2635);
and U3406 (N_3406,In_2709,In_237);
nor U3407 (N_3407,In_1738,In_1337);
xnor U3408 (N_3408,In_332,In_1344);
nor U3409 (N_3409,In_716,In_2765);
nand U3410 (N_3410,In_254,In_789);
nand U3411 (N_3411,In_2867,In_1441);
and U3412 (N_3412,In_1512,In_1976);
nand U3413 (N_3413,In_923,In_1203);
xnor U3414 (N_3414,In_1260,In_80);
nor U3415 (N_3415,In_1620,In_329);
nor U3416 (N_3416,In_2868,In_1732);
nor U3417 (N_3417,In_937,In_2854);
nor U3418 (N_3418,In_1872,In_1168);
nor U3419 (N_3419,In_2287,In_1977);
nand U3420 (N_3420,In_741,In_2842);
xnor U3421 (N_3421,In_710,In_92);
nor U3422 (N_3422,In_2062,In_92);
or U3423 (N_3423,In_990,In_2940);
and U3424 (N_3424,In_2703,In_1552);
or U3425 (N_3425,In_2570,In_743);
and U3426 (N_3426,In_184,In_755);
and U3427 (N_3427,In_877,In_2965);
nand U3428 (N_3428,In_948,In_1556);
nand U3429 (N_3429,In_2206,In_2401);
and U3430 (N_3430,In_1362,In_1911);
and U3431 (N_3431,In_1708,In_1367);
and U3432 (N_3432,In_1774,In_2692);
nor U3433 (N_3433,In_2625,In_1915);
nor U3434 (N_3434,In_2816,In_1454);
or U3435 (N_3435,In_2052,In_559);
or U3436 (N_3436,In_1283,In_848);
or U3437 (N_3437,In_662,In_1201);
or U3438 (N_3438,In_1500,In_2187);
and U3439 (N_3439,In_1154,In_482);
xor U3440 (N_3440,In_2009,In_2101);
or U3441 (N_3441,In_2526,In_1574);
nand U3442 (N_3442,In_1403,In_1964);
nor U3443 (N_3443,In_1773,In_442);
or U3444 (N_3444,In_615,In_363);
nor U3445 (N_3445,In_564,In_62);
xnor U3446 (N_3446,In_2674,In_309);
or U3447 (N_3447,In_2890,In_1671);
xor U3448 (N_3448,In_4,In_1667);
nand U3449 (N_3449,In_1044,In_2276);
nand U3450 (N_3450,In_1183,In_2511);
xnor U3451 (N_3451,In_1933,In_2594);
or U3452 (N_3452,In_2527,In_1020);
nor U3453 (N_3453,In_956,In_1894);
or U3454 (N_3454,In_2294,In_1350);
or U3455 (N_3455,In_1860,In_899);
nand U3456 (N_3456,In_2077,In_253);
nor U3457 (N_3457,In_212,In_739);
nand U3458 (N_3458,In_2807,In_2611);
or U3459 (N_3459,In_1783,In_1649);
nand U3460 (N_3460,In_753,In_2343);
or U3461 (N_3461,In_2068,In_1770);
xnor U3462 (N_3462,In_26,In_1294);
and U3463 (N_3463,In_2385,In_2490);
nand U3464 (N_3464,In_537,In_812);
and U3465 (N_3465,In_290,In_2699);
or U3466 (N_3466,In_309,In_24);
nand U3467 (N_3467,In_2401,In_1606);
xnor U3468 (N_3468,In_122,In_244);
or U3469 (N_3469,In_1775,In_904);
and U3470 (N_3470,In_1065,In_2730);
and U3471 (N_3471,In_1324,In_666);
nor U3472 (N_3472,In_264,In_2808);
and U3473 (N_3473,In_2827,In_1290);
nand U3474 (N_3474,In_1162,In_1366);
nor U3475 (N_3475,In_502,In_974);
nor U3476 (N_3476,In_553,In_1614);
nand U3477 (N_3477,In_1446,In_288);
or U3478 (N_3478,In_988,In_2798);
nor U3479 (N_3479,In_979,In_332);
and U3480 (N_3480,In_2254,In_2353);
and U3481 (N_3481,In_943,In_1758);
or U3482 (N_3482,In_2648,In_2297);
xnor U3483 (N_3483,In_2061,In_150);
and U3484 (N_3484,In_1874,In_2843);
or U3485 (N_3485,In_1874,In_1863);
and U3486 (N_3486,In_2360,In_2641);
nand U3487 (N_3487,In_2979,In_1770);
nand U3488 (N_3488,In_1762,In_1568);
nor U3489 (N_3489,In_2504,In_577);
nand U3490 (N_3490,In_2701,In_1049);
and U3491 (N_3491,In_2367,In_1140);
or U3492 (N_3492,In_2245,In_2422);
xnor U3493 (N_3493,In_2671,In_1182);
and U3494 (N_3494,In_2527,In_2916);
xor U3495 (N_3495,In_1235,In_801);
and U3496 (N_3496,In_2821,In_532);
nor U3497 (N_3497,In_2584,In_425);
or U3498 (N_3498,In_2368,In_2795);
nand U3499 (N_3499,In_678,In_1215);
nor U3500 (N_3500,In_479,In_1980);
nor U3501 (N_3501,In_540,In_2491);
or U3502 (N_3502,In_1196,In_2893);
nand U3503 (N_3503,In_2228,In_1148);
or U3504 (N_3504,In_1615,In_838);
and U3505 (N_3505,In_795,In_129);
and U3506 (N_3506,In_2057,In_1013);
nor U3507 (N_3507,In_2262,In_1818);
or U3508 (N_3508,In_2321,In_838);
nor U3509 (N_3509,In_1794,In_586);
or U3510 (N_3510,In_2563,In_955);
nand U3511 (N_3511,In_662,In_199);
xnor U3512 (N_3512,In_1079,In_1468);
nor U3513 (N_3513,In_907,In_2746);
or U3514 (N_3514,In_1853,In_2283);
and U3515 (N_3515,In_2558,In_1598);
nor U3516 (N_3516,In_694,In_1042);
xor U3517 (N_3517,In_1818,In_1058);
xnor U3518 (N_3518,In_748,In_1843);
nor U3519 (N_3519,In_2035,In_148);
nand U3520 (N_3520,In_1835,In_1276);
nor U3521 (N_3521,In_1750,In_2669);
and U3522 (N_3522,In_771,In_1508);
nor U3523 (N_3523,In_2986,In_687);
and U3524 (N_3524,In_2732,In_1687);
or U3525 (N_3525,In_121,In_2458);
nand U3526 (N_3526,In_218,In_1748);
nand U3527 (N_3527,In_2744,In_1531);
nor U3528 (N_3528,In_388,In_2343);
and U3529 (N_3529,In_2016,In_2754);
xnor U3530 (N_3530,In_258,In_1032);
nand U3531 (N_3531,In_1161,In_911);
or U3532 (N_3532,In_1056,In_2836);
and U3533 (N_3533,In_2988,In_477);
or U3534 (N_3534,In_666,In_2861);
xor U3535 (N_3535,In_1105,In_1530);
nand U3536 (N_3536,In_2488,In_2717);
and U3537 (N_3537,In_2143,In_1800);
and U3538 (N_3538,In_2908,In_2887);
nand U3539 (N_3539,In_2289,In_2631);
and U3540 (N_3540,In_2226,In_81);
xor U3541 (N_3541,In_2795,In_1331);
and U3542 (N_3542,In_1133,In_2624);
and U3543 (N_3543,In_2902,In_1549);
nand U3544 (N_3544,In_2409,In_430);
and U3545 (N_3545,In_2194,In_1762);
xnor U3546 (N_3546,In_2879,In_236);
nand U3547 (N_3547,In_210,In_1550);
xor U3548 (N_3548,In_467,In_2200);
or U3549 (N_3549,In_1838,In_199);
nor U3550 (N_3550,In_1828,In_1361);
nor U3551 (N_3551,In_1615,In_1142);
and U3552 (N_3552,In_1111,In_372);
nor U3553 (N_3553,In_2549,In_996);
nand U3554 (N_3554,In_1951,In_337);
nand U3555 (N_3555,In_1363,In_830);
or U3556 (N_3556,In_1539,In_301);
nor U3557 (N_3557,In_1804,In_2837);
xor U3558 (N_3558,In_2786,In_1096);
xnor U3559 (N_3559,In_2567,In_2428);
nor U3560 (N_3560,In_636,In_1425);
xnor U3561 (N_3561,In_1726,In_507);
nor U3562 (N_3562,In_1641,In_2081);
or U3563 (N_3563,In_1097,In_2134);
and U3564 (N_3564,In_2594,In_2005);
nand U3565 (N_3565,In_2034,In_1861);
nand U3566 (N_3566,In_1603,In_1881);
or U3567 (N_3567,In_56,In_1625);
nor U3568 (N_3568,In_2687,In_2846);
and U3569 (N_3569,In_1659,In_2960);
nand U3570 (N_3570,In_2452,In_2681);
xnor U3571 (N_3571,In_2442,In_1392);
nand U3572 (N_3572,In_2131,In_455);
or U3573 (N_3573,In_705,In_2252);
and U3574 (N_3574,In_1436,In_118);
nor U3575 (N_3575,In_2699,In_2921);
or U3576 (N_3576,In_1937,In_628);
nor U3577 (N_3577,In_2161,In_1662);
nand U3578 (N_3578,In_2278,In_2555);
nand U3579 (N_3579,In_2897,In_2268);
nor U3580 (N_3580,In_1524,In_2436);
xnor U3581 (N_3581,In_1396,In_593);
or U3582 (N_3582,In_2265,In_604);
or U3583 (N_3583,In_805,In_1788);
nand U3584 (N_3584,In_2210,In_1398);
and U3585 (N_3585,In_2655,In_1406);
xor U3586 (N_3586,In_1774,In_210);
and U3587 (N_3587,In_1705,In_1326);
nand U3588 (N_3588,In_2669,In_2829);
nand U3589 (N_3589,In_2506,In_1129);
or U3590 (N_3590,In_641,In_1133);
xnor U3591 (N_3591,In_1955,In_1637);
or U3592 (N_3592,In_468,In_1);
and U3593 (N_3593,In_127,In_2695);
and U3594 (N_3594,In_43,In_2846);
nor U3595 (N_3595,In_1434,In_1013);
and U3596 (N_3596,In_603,In_2619);
xor U3597 (N_3597,In_1,In_2220);
nor U3598 (N_3598,In_2030,In_984);
and U3599 (N_3599,In_1755,In_892);
or U3600 (N_3600,In_1496,In_1366);
nor U3601 (N_3601,In_2562,In_452);
and U3602 (N_3602,In_216,In_1170);
nor U3603 (N_3603,In_2151,In_2987);
nand U3604 (N_3604,In_1641,In_104);
and U3605 (N_3605,In_533,In_1445);
or U3606 (N_3606,In_2805,In_2581);
xnor U3607 (N_3607,In_2180,In_841);
and U3608 (N_3608,In_2724,In_999);
and U3609 (N_3609,In_1037,In_546);
and U3610 (N_3610,In_1354,In_860);
and U3611 (N_3611,In_2688,In_2031);
or U3612 (N_3612,In_908,In_1404);
nand U3613 (N_3613,In_389,In_225);
nor U3614 (N_3614,In_413,In_2356);
xor U3615 (N_3615,In_2556,In_2990);
and U3616 (N_3616,In_1042,In_91);
and U3617 (N_3617,In_136,In_1475);
xnor U3618 (N_3618,In_619,In_1923);
nand U3619 (N_3619,In_2587,In_1793);
or U3620 (N_3620,In_1762,In_1059);
and U3621 (N_3621,In_1456,In_1532);
nand U3622 (N_3622,In_287,In_545);
nand U3623 (N_3623,In_1002,In_1081);
or U3624 (N_3624,In_1966,In_1082);
and U3625 (N_3625,In_1917,In_2230);
nand U3626 (N_3626,In_408,In_1614);
nor U3627 (N_3627,In_155,In_2731);
and U3628 (N_3628,In_1683,In_68);
or U3629 (N_3629,In_2669,In_2313);
nand U3630 (N_3630,In_2918,In_1695);
xnor U3631 (N_3631,In_1228,In_1191);
nand U3632 (N_3632,In_354,In_2980);
and U3633 (N_3633,In_2089,In_1277);
nand U3634 (N_3634,In_2125,In_795);
or U3635 (N_3635,In_360,In_1086);
and U3636 (N_3636,In_2998,In_1882);
and U3637 (N_3637,In_2282,In_1549);
nand U3638 (N_3638,In_2164,In_535);
nand U3639 (N_3639,In_1018,In_474);
and U3640 (N_3640,In_2936,In_532);
xnor U3641 (N_3641,In_2445,In_1938);
nor U3642 (N_3642,In_2505,In_2727);
nand U3643 (N_3643,In_597,In_841);
nor U3644 (N_3644,In_155,In_1830);
xor U3645 (N_3645,In_430,In_1616);
or U3646 (N_3646,In_737,In_1775);
nand U3647 (N_3647,In_876,In_1765);
nor U3648 (N_3648,In_2635,In_1047);
nor U3649 (N_3649,In_1146,In_798);
nand U3650 (N_3650,In_2198,In_2541);
and U3651 (N_3651,In_561,In_964);
xor U3652 (N_3652,In_233,In_640);
and U3653 (N_3653,In_1915,In_1854);
nand U3654 (N_3654,In_900,In_1595);
or U3655 (N_3655,In_120,In_2930);
nor U3656 (N_3656,In_2823,In_2662);
or U3657 (N_3657,In_2878,In_647);
or U3658 (N_3658,In_1912,In_2822);
or U3659 (N_3659,In_1366,In_501);
or U3660 (N_3660,In_461,In_1024);
xnor U3661 (N_3661,In_122,In_2855);
xnor U3662 (N_3662,In_1602,In_349);
and U3663 (N_3663,In_1198,In_661);
and U3664 (N_3664,In_288,In_2815);
xnor U3665 (N_3665,In_1885,In_2178);
and U3666 (N_3666,In_2517,In_1483);
or U3667 (N_3667,In_342,In_998);
xor U3668 (N_3668,In_133,In_2199);
nor U3669 (N_3669,In_888,In_1843);
or U3670 (N_3670,In_1519,In_2317);
and U3671 (N_3671,In_377,In_739);
and U3672 (N_3672,In_2637,In_97);
xnor U3673 (N_3673,In_612,In_1659);
nand U3674 (N_3674,In_238,In_1738);
nor U3675 (N_3675,In_2220,In_2483);
nor U3676 (N_3676,In_1444,In_2178);
nand U3677 (N_3677,In_334,In_1446);
xor U3678 (N_3678,In_2454,In_987);
or U3679 (N_3679,In_469,In_817);
and U3680 (N_3680,In_39,In_2060);
xnor U3681 (N_3681,In_2910,In_2623);
nor U3682 (N_3682,In_1059,In_1196);
nor U3683 (N_3683,In_1422,In_1995);
or U3684 (N_3684,In_685,In_1607);
nor U3685 (N_3685,In_2510,In_1295);
xor U3686 (N_3686,In_1339,In_1890);
nand U3687 (N_3687,In_1862,In_2288);
nor U3688 (N_3688,In_1476,In_417);
xor U3689 (N_3689,In_2642,In_358);
nand U3690 (N_3690,In_2070,In_2811);
nand U3691 (N_3691,In_2217,In_1092);
and U3692 (N_3692,In_2978,In_2146);
nand U3693 (N_3693,In_2790,In_2752);
nand U3694 (N_3694,In_2540,In_349);
nor U3695 (N_3695,In_582,In_1801);
or U3696 (N_3696,In_282,In_2859);
or U3697 (N_3697,In_1785,In_518);
nand U3698 (N_3698,In_2839,In_1899);
nand U3699 (N_3699,In_66,In_2043);
nand U3700 (N_3700,In_1388,In_2157);
nor U3701 (N_3701,In_2179,In_1754);
nor U3702 (N_3702,In_115,In_2115);
and U3703 (N_3703,In_2745,In_2935);
or U3704 (N_3704,In_1218,In_1140);
nand U3705 (N_3705,In_1359,In_1603);
nand U3706 (N_3706,In_24,In_290);
and U3707 (N_3707,In_2171,In_1344);
nand U3708 (N_3708,In_2642,In_2676);
and U3709 (N_3709,In_2629,In_2084);
nand U3710 (N_3710,In_705,In_1109);
or U3711 (N_3711,In_466,In_2676);
nand U3712 (N_3712,In_1983,In_2441);
and U3713 (N_3713,In_2590,In_2209);
or U3714 (N_3714,In_1181,In_207);
nor U3715 (N_3715,In_2137,In_2592);
nor U3716 (N_3716,In_1515,In_1491);
or U3717 (N_3717,In_2536,In_2190);
or U3718 (N_3718,In_491,In_78);
nand U3719 (N_3719,In_2050,In_1538);
and U3720 (N_3720,In_1868,In_1032);
or U3721 (N_3721,In_2920,In_413);
or U3722 (N_3722,In_59,In_2129);
and U3723 (N_3723,In_610,In_2186);
or U3724 (N_3724,In_1880,In_2397);
nand U3725 (N_3725,In_255,In_90);
or U3726 (N_3726,In_2529,In_2161);
and U3727 (N_3727,In_2516,In_415);
nand U3728 (N_3728,In_2985,In_256);
and U3729 (N_3729,In_2593,In_1980);
nand U3730 (N_3730,In_388,In_1742);
or U3731 (N_3731,In_908,In_2304);
and U3732 (N_3732,In_777,In_795);
or U3733 (N_3733,In_2999,In_2822);
nor U3734 (N_3734,In_700,In_1300);
nand U3735 (N_3735,In_151,In_2489);
nand U3736 (N_3736,In_2303,In_2588);
nand U3737 (N_3737,In_941,In_2613);
xor U3738 (N_3738,In_3,In_1987);
or U3739 (N_3739,In_22,In_861);
nand U3740 (N_3740,In_1634,In_1097);
nand U3741 (N_3741,In_1511,In_847);
or U3742 (N_3742,In_1183,In_1430);
nand U3743 (N_3743,In_600,In_499);
and U3744 (N_3744,In_323,In_603);
nor U3745 (N_3745,In_219,In_2929);
nand U3746 (N_3746,In_2795,In_2222);
nand U3747 (N_3747,In_1570,In_2996);
nor U3748 (N_3748,In_44,In_581);
and U3749 (N_3749,In_140,In_2121);
nand U3750 (N_3750,In_1115,In_1736);
nor U3751 (N_3751,In_914,In_31);
nand U3752 (N_3752,In_340,In_2143);
and U3753 (N_3753,In_1237,In_2171);
or U3754 (N_3754,In_239,In_241);
nor U3755 (N_3755,In_354,In_1247);
nor U3756 (N_3756,In_2551,In_623);
nand U3757 (N_3757,In_1369,In_2905);
xor U3758 (N_3758,In_2870,In_1548);
nor U3759 (N_3759,In_71,In_1019);
and U3760 (N_3760,In_2024,In_293);
and U3761 (N_3761,In_2898,In_1649);
and U3762 (N_3762,In_447,In_1343);
and U3763 (N_3763,In_358,In_2516);
nor U3764 (N_3764,In_104,In_2386);
and U3765 (N_3765,In_1049,In_2593);
nand U3766 (N_3766,In_1663,In_794);
nand U3767 (N_3767,In_2827,In_1512);
nor U3768 (N_3768,In_2727,In_2353);
and U3769 (N_3769,In_213,In_1144);
nor U3770 (N_3770,In_640,In_2681);
nor U3771 (N_3771,In_875,In_2317);
and U3772 (N_3772,In_1587,In_2878);
nand U3773 (N_3773,In_2385,In_565);
or U3774 (N_3774,In_1735,In_2087);
nand U3775 (N_3775,In_419,In_867);
or U3776 (N_3776,In_2412,In_50);
and U3777 (N_3777,In_2310,In_1074);
or U3778 (N_3778,In_2576,In_665);
xor U3779 (N_3779,In_1765,In_2607);
and U3780 (N_3780,In_2055,In_1933);
nor U3781 (N_3781,In_488,In_992);
or U3782 (N_3782,In_121,In_599);
nor U3783 (N_3783,In_2,In_1115);
nand U3784 (N_3784,In_185,In_881);
nand U3785 (N_3785,In_725,In_680);
nor U3786 (N_3786,In_158,In_2469);
and U3787 (N_3787,In_1522,In_935);
and U3788 (N_3788,In_1681,In_1106);
nand U3789 (N_3789,In_84,In_1181);
and U3790 (N_3790,In_826,In_2963);
nor U3791 (N_3791,In_2707,In_1035);
nand U3792 (N_3792,In_2223,In_2050);
nand U3793 (N_3793,In_964,In_1346);
and U3794 (N_3794,In_2301,In_1546);
and U3795 (N_3795,In_278,In_485);
nand U3796 (N_3796,In_2796,In_680);
and U3797 (N_3797,In_824,In_2084);
and U3798 (N_3798,In_2681,In_2355);
or U3799 (N_3799,In_1842,In_748);
nand U3800 (N_3800,In_533,In_721);
nand U3801 (N_3801,In_11,In_2251);
nand U3802 (N_3802,In_576,In_2845);
nor U3803 (N_3803,In_1547,In_2679);
nand U3804 (N_3804,In_746,In_1697);
nor U3805 (N_3805,In_1556,In_2190);
xor U3806 (N_3806,In_859,In_1284);
or U3807 (N_3807,In_2461,In_1668);
and U3808 (N_3808,In_2899,In_2910);
or U3809 (N_3809,In_775,In_680);
nor U3810 (N_3810,In_1798,In_339);
nor U3811 (N_3811,In_595,In_1526);
nor U3812 (N_3812,In_1095,In_2240);
or U3813 (N_3813,In_2043,In_305);
nor U3814 (N_3814,In_1937,In_1538);
xnor U3815 (N_3815,In_1737,In_1676);
or U3816 (N_3816,In_501,In_3);
or U3817 (N_3817,In_1357,In_419);
or U3818 (N_3818,In_1526,In_1017);
and U3819 (N_3819,In_1147,In_2433);
or U3820 (N_3820,In_2621,In_1400);
nand U3821 (N_3821,In_827,In_2173);
or U3822 (N_3822,In_149,In_519);
nand U3823 (N_3823,In_2939,In_1385);
nand U3824 (N_3824,In_1427,In_1225);
or U3825 (N_3825,In_1727,In_1287);
nor U3826 (N_3826,In_1818,In_1573);
or U3827 (N_3827,In_2788,In_1847);
nand U3828 (N_3828,In_2448,In_215);
xnor U3829 (N_3829,In_2940,In_461);
nand U3830 (N_3830,In_2992,In_1760);
or U3831 (N_3831,In_1423,In_784);
and U3832 (N_3832,In_36,In_2480);
xor U3833 (N_3833,In_2376,In_2096);
nand U3834 (N_3834,In_179,In_87);
xor U3835 (N_3835,In_1439,In_2273);
nand U3836 (N_3836,In_1217,In_1716);
or U3837 (N_3837,In_587,In_1176);
and U3838 (N_3838,In_2475,In_2255);
nand U3839 (N_3839,In_1816,In_2105);
and U3840 (N_3840,In_1348,In_2999);
nand U3841 (N_3841,In_2074,In_2417);
or U3842 (N_3842,In_1878,In_1598);
and U3843 (N_3843,In_831,In_548);
or U3844 (N_3844,In_1510,In_1225);
and U3845 (N_3845,In_1989,In_2303);
or U3846 (N_3846,In_1402,In_351);
nor U3847 (N_3847,In_405,In_2507);
nor U3848 (N_3848,In_2026,In_340);
xnor U3849 (N_3849,In_409,In_2994);
nor U3850 (N_3850,In_1055,In_2100);
and U3851 (N_3851,In_1578,In_370);
and U3852 (N_3852,In_1770,In_2796);
or U3853 (N_3853,In_1826,In_2621);
and U3854 (N_3854,In_1905,In_1988);
xor U3855 (N_3855,In_1477,In_1744);
or U3856 (N_3856,In_1822,In_2763);
nand U3857 (N_3857,In_1857,In_533);
nand U3858 (N_3858,In_748,In_1202);
nor U3859 (N_3859,In_1502,In_2856);
and U3860 (N_3860,In_1841,In_190);
and U3861 (N_3861,In_1350,In_2129);
nor U3862 (N_3862,In_2989,In_51);
and U3863 (N_3863,In_691,In_884);
and U3864 (N_3864,In_1510,In_845);
nor U3865 (N_3865,In_2540,In_2712);
or U3866 (N_3866,In_756,In_2116);
or U3867 (N_3867,In_42,In_827);
nand U3868 (N_3868,In_2349,In_570);
nor U3869 (N_3869,In_1972,In_1754);
nand U3870 (N_3870,In_1464,In_2022);
nand U3871 (N_3871,In_1740,In_1975);
and U3872 (N_3872,In_2721,In_2718);
and U3873 (N_3873,In_1765,In_1600);
xor U3874 (N_3874,In_2510,In_2434);
and U3875 (N_3875,In_1211,In_953);
and U3876 (N_3876,In_1874,In_1175);
nand U3877 (N_3877,In_2814,In_704);
nor U3878 (N_3878,In_305,In_693);
nand U3879 (N_3879,In_1971,In_179);
nor U3880 (N_3880,In_349,In_1584);
nor U3881 (N_3881,In_413,In_653);
nor U3882 (N_3882,In_2116,In_2028);
xnor U3883 (N_3883,In_2921,In_680);
and U3884 (N_3884,In_648,In_961);
nor U3885 (N_3885,In_1564,In_369);
or U3886 (N_3886,In_750,In_1797);
or U3887 (N_3887,In_2671,In_1494);
nor U3888 (N_3888,In_1353,In_2923);
or U3889 (N_3889,In_1950,In_2437);
and U3890 (N_3890,In_763,In_915);
nand U3891 (N_3891,In_238,In_820);
nand U3892 (N_3892,In_2372,In_1519);
xnor U3893 (N_3893,In_1627,In_1205);
nor U3894 (N_3894,In_1978,In_1205);
or U3895 (N_3895,In_949,In_1353);
nand U3896 (N_3896,In_1751,In_84);
nor U3897 (N_3897,In_2715,In_589);
nand U3898 (N_3898,In_1997,In_1277);
or U3899 (N_3899,In_597,In_423);
nand U3900 (N_3900,In_806,In_451);
nand U3901 (N_3901,In_2433,In_655);
or U3902 (N_3902,In_2948,In_751);
nor U3903 (N_3903,In_2337,In_425);
nand U3904 (N_3904,In_1869,In_749);
nand U3905 (N_3905,In_2614,In_1947);
nor U3906 (N_3906,In_1800,In_1970);
or U3907 (N_3907,In_1498,In_1610);
nand U3908 (N_3908,In_965,In_2474);
xnor U3909 (N_3909,In_1524,In_379);
and U3910 (N_3910,In_2142,In_2944);
and U3911 (N_3911,In_1054,In_1531);
nand U3912 (N_3912,In_2352,In_2258);
or U3913 (N_3913,In_1415,In_2527);
nand U3914 (N_3914,In_2395,In_664);
nand U3915 (N_3915,In_875,In_330);
and U3916 (N_3916,In_566,In_2749);
xnor U3917 (N_3917,In_1578,In_2265);
nand U3918 (N_3918,In_2102,In_519);
or U3919 (N_3919,In_2043,In_426);
nand U3920 (N_3920,In_91,In_2425);
nor U3921 (N_3921,In_484,In_2157);
nor U3922 (N_3922,In_649,In_2377);
xor U3923 (N_3923,In_2770,In_1481);
nor U3924 (N_3924,In_1834,In_2503);
and U3925 (N_3925,In_2124,In_490);
or U3926 (N_3926,In_2698,In_141);
or U3927 (N_3927,In_192,In_1660);
xnor U3928 (N_3928,In_1645,In_412);
nor U3929 (N_3929,In_877,In_176);
nand U3930 (N_3930,In_29,In_2389);
nor U3931 (N_3931,In_419,In_2521);
and U3932 (N_3932,In_1031,In_2016);
or U3933 (N_3933,In_436,In_34);
and U3934 (N_3934,In_1431,In_2044);
nor U3935 (N_3935,In_2188,In_716);
and U3936 (N_3936,In_2649,In_2302);
xnor U3937 (N_3937,In_2680,In_2754);
or U3938 (N_3938,In_1333,In_1250);
nor U3939 (N_3939,In_1267,In_1135);
nor U3940 (N_3940,In_736,In_288);
or U3941 (N_3941,In_2610,In_164);
nand U3942 (N_3942,In_450,In_273);
xnor U3943 (N_3943,In_1407,In_2221);
and U3944 (N_3944,In_2999,In_1072);
and U3945 (N_3945,In_450,In_845);
and U3946 (N_3946,In_1712,In_893);
or U3947 (N_3947,In_1412,In_435);
and U3948 (N_3948,In_2975,In_136);
and U3949 (N_3949,In_2163,In_1781);
nor U3950 (N_3950,In_2951,In_543);
nand U3951 (N_3951,In_1837,In_2444);
nand U3952 (N_3952,In_2783,In_1190);
nor U3953 (N_3953,In_342,In_1728);
nor U3954 (N_3954,In_382,In_2232);
xnor U3955 (N_3955,In_1096,In_682);
nand U3956 (N_3956,In_161,In_1414);
or U3957 (N_3957,In_1697,In_2294);
and U3958 (N_3958,In_1553,In_1969);
nand U3959 (N_3959,In_1281,In_609);
nand U3960 (N_3960,In_589,In_957);
nand U3961 (N_3961,In_1112,In_1585);
nor U3962 (N_3962,In_904,In_2645);
nor U3963 (N_3963,In_2264,In_1281);
or U3964 (N_3964,In_1266,In_8);
or U3965 (N_3965,In_2738,In_2129);
and U3966 (N_3966,In_2320,In_893);
nor U3967 (N_3967,In_1975,In_416);
nand U3968 (N_3968,In_1170,In_36);
or U3969 (N_3969,In_1078,In_277);
nor U3970 (N_3970,In_353,In_2584);
nor U3971 (N_3971,In_1896,In_1950);
and U3972 (N_3972,In_1481,In_1368);
nor U3973 (N_3973,In_267,In_1939);
nand U3974 (N_3974,In_639,In_982);
nand U3975 (N_3975,In_2033,In_287);
xnor U3976 (N_3976,In_565,In_2976);
and U3977 (N_3977,In_2848,In_2834);
xor U3978 (N_3978,In_169,In_419);
xnor U3979 (N_3979,In_1131,In_503);
nand U3980 (N_3980,In_2280,In_1508);
and U3981 (N_3981,In_1746,In_596);
nor U3982 (N_3982,In_2210,In_675);
nor U3983 (N_3983,In_1165,In_2893);
or U3984 (N_3984,In_1875,In_819);
nor U3985 (N_3985,In_1965,In_1838);
nor U3986 (N_3986,In_2286,In_1209);
nor U3987 (N_3987,In_1399,In_2821);
nor U3988 (N_3988,In_1164,In_1647);
and U3989 (N_3989,In_566,In_154);
and U3990 (N_3990,In_789,In_2609);
or U3991 (N_3991,In_2465,In_26);
and U3992 (N_3992,In_853,In_152);
or U3993 (N_3993,In_1781,In_997);
or U3994 (N_3994,In_2706,In_1102);
nand U3995 (N_3995,In_866,In_1598);
and U3996 (N_3996,In_1206,In_713);
and U3997 (N_3997,In_1407,In_133);
and U3998 (N_3998,In_2726,In_1541);
nand U3999 (N_3999,In_2241,In_1959);
nor U4000 (N_4000,In_2632,In_1102);
or U4001 (N_4001,In_1819,In_311);
or U4002 (N_4002,In_233,In_2700);
and U4003 (N_4003,In_1547,In_545);
xor U4004 (N_4004,In_1601,In_2037);
nor U4005 (N_4005,In_201,In_742);
nand U4006 (N_4006,In_2153,In_2577);
or U4007 (N_4007,In_2145,In_2663);
nand U4008 (N_4008,In_1346,In_2279);
nor U4009 (N_4009,In_270,In_2176);
nor U4010 (N_4010,In_495,In_1595);
nor U4011 (N_4011,In_2268,In_2051);
nor U4012 (N_4012,In_1117,In_1338);
and U4013 (N_4013,In_1074,In_1126);
nand U4014 (N_4014,In_1966,In_2921);
nand U4015 (N_4015,In_1632,In_1881);
or U4016 (N_4016,In_2420,In_1719);
xor U4017 (N_4017,In_215,In_2147);
nand U4018 (N_4018,In_837,In_986);
nand U4019 (N_4019,In_2218,In_1635);
or U4020 (N_4020,In_239,In_161);
or U4021 (N_4021,In_319,In_91);
xnor U4022 (N_4022,In_178,In_1092);
xnor U4023 (N_4023,In_2752,In_2145);
nand U4024 (N_4024,In_1122,In_2548);
xor U4025 (N_4025,In_1256,In_1397);
nor U4026 (N_4026,In_2709,In_2079);
nor U4027 (N_4027,In_2991,In_2304);
nor U4028 (N_4028,In_1440,In_390);
or U4029 (N_4029,In_2103,In_2329);
and U4030 (N_4030,In_695,In_2945);
xnor U4031 (N_4031,In_18,In_676);
nand U4032 (N_4032,In_612,In_130);
nand U4033 (N_4033,In_209,In_1827);
nor U4034 (N_4034,In_183,In_1597);
xnor U4035 (N_4035,In_698,In_2947);
nor U4036 (N_4036,In_6,In_135);
nand U4037 (N_4037,In_2324,In_1434);
nand U4038 (N_4038,In_331,In_16);
or U4039 (N_4039,In_962,In_2533);
or U4040 (N_4040,In_376,In_2575);
and U4041 (N_4041,In_685,In_2471);
nand U4042 (N_4042,In_2520,In_1368);
nor U4043 (N_4043,In_236,In_990);
xnor U4044 (N_4044,In_2715,In_264);
nand U4045 (N_4045,In_1177,In_1527);
nand U4046 (N_4046,In_2347,In_2993);
nor U4047 (N_4047,In_2145,In_2417);
nor U4048 (N_4048,In_2147,In_1463);
nor U4049 (N_4049,In_1027,In_226);
and U4050 (N_4050,In_285,In_2458);
and U4051 (N_4051,In_1513,In_1886);
nor U4052 (N_4052,In_1859,In_1750);
nand U4053 (N_4053,In_2968,In_1813);
nor U4054 (N_4054,In_563,In_1429);
nor U4055 (N_4055,In_2756,In_1200);
or U4056 (N_4056,In_1334,In_1373);
and U4057 (N_4057,In_66,In_1496);
nand U4058 (N_4058,In_1938,In_1796);
or U4059 (N_4059,In_898,In_2611);
nand U4060 (N_4060,In_954,In_2776);
and U4061 (N_4061,In_935,In_2556);
nand U4062 (N_4062,In_2243,In_1489);
nand U4063 (N_4063,In_1047,In_2633);
and U4064 (N_4064,In_1447,In_1926);
nand U4065 (N_4065,In_1533,In_2109);
or U4066 (N_4066,In_1301,In_2633);
or U4067 (N_4067,In_1230,In_1271);
nor U4068 (N_4068,In_1812,In_393);
xnor U4069 (N_4069,In_1731,In_2489);
and U4070 (N_4070,In_1602,In_2516);
and U4071 (N_4071,In_2299,In_2957);
nor U4072 (N_4072,In_2746,In_1455);
xor U4073 (N_4073,In_2349,In_1384);
or U4074 (N_4074,In_2807,In_523);
xor U4075 (N_4075,In_1233,In_1615);
nor U4076 (N_4076,In_141,In_2140);
nand U4077 (N_4077,In_1384,In_1218);
and U4078 (N_4078,In_928,In_1333);
nand U4079 (N_4079,In_1367,In_1308);
nor U4080 (N_4080,In_2583,In_1313);
or U4081 (N_4081,In_1616,In_1688);
nand U4082 (N_4082,In_999,In_2908);
and U4083 (N_4083,In_107,In_1764);
and U4084 (N_4084,In_627,In_2175);
or U4085 (N_4085,In_2215,In_422);
nand U4086 (N_4086,In_2135,In_1295);
and U4087 (N_4087,In_2267,In_797);
nor U4088 (N_4088,In_464,In_678);
nor U4089 (N_4089,In_2653,In_83);
or U4090 (N_4090,In_553,In_2635);
nor U4091 (N_4091,In_1568,In_2367);
nand U4092 (N_4092,In_2539,In_1304);
nor U4093 (N_4093,In_2517,In_1891);
nand U4094 (N_4094,In_560,In_2167);
nor U4095 (N_4095,In_2366,In_262);
nor U4096 (N_4096,In_2795,In_1321);
nand U4097 (N_4097,In_2502,In_160);
xor U4098 (N_4098,In_2,In_2470);
nand U4099 (N_4099,In_638,In_1448);
nand U4100 (N_4100,In_2822,In_2640);
or U4101 (N_4101,In_520,In_1354);
xnor U4102 (N_4102,In_2951,In_109);
nand U4103 (N_4103,In_2866,In_2840);
nor U4104 (N_4104,In_2922,In_250);
or U4105 (N_4105,In_1036,In_2103);
and U4106 (N_4106,In_778,In_1007);
xnor U4107 (N_4107,In_1775,In_2342);
and U4108 (N_4108,In_2846,In_1326);
nand U4109 (N_4109,In_1255,In_1003);
and U4110 (N_4110,In_2713,In_233);
nand U4111 (N_4111,In_1364,In_619);
xnor U4112 (N_4112,In_2927,In_2658);
and U4113 (N_4113,In_2068,In_339);
xnor U4114 (N_4114,In_2370,In_559);
or U4115 (N_4115,In_426,In_1677);
or U4116 (N_4116,In_1105,In_2538);
or U4117 (N_4117,In_1771,In_964);
nor U4118 (N_4118,In_2377,In_2144);
and U4119 (N_4119,In_1501,In_542);
nand U4120 (N_4120,In_1515,In_2549);
nand U4121 (N_4121,In_1496,In_2269);
or U4122 (N_4122,In_2818,In_453);
or U4123 (N_4123,In_2501,In_2581);
or U4124 (N_4124,In_368,In_2041);
or U4125 (N_4125,In_2503,In_1352);
nor U4126 (N_4126,In_643,In_652);
and U4127 (N_4127,In_1421,In_266);
and U4128 (N_4128,In_539,In_2056);
nor U4129 (N_4129,In_1309,In_1485);
and U4130 (N_4130,In_1281,In_2230);
and U4131 (N_4131,In_2049,In_1551);
and U4132 (N_4132,In_224,In_333);
and U4133 (N_4133,In_1906,In_1524);
xor U4134 (N_4134,In_2615,In_2187);
or U4135 (N_4135,In_943,In_2668);
and U4136 (N_4136,In_1535,In_2865);
and U4137 (N_4137,In_2124,In_2421);
or U4138 (N_4138,In_1962,In_1863);
nand U4139 (N_4139,In_1998,In_773);
and U4140 (N_4140,In_2650,In_1285);
nor U4141 (N_4141,In_648,In_169);
or U4142 (N_4142,In_1712,In_2264);
nor U4143 (N_4143,In_1773,In_1950);
or U4144 (N_4144,In_1729,In_144);
nor U4145 (N_4145,In_400,In_1679);
nor U4146 (N_4146,In_1693,In_2349);
nor U4147 (N_4147,In_865,In_2482);
or U4148 (N_4148,In_652,In_656);
or U4149 (N_4149,In_348,In_382);
nor U4150 (N_4150,In_1462,In_1346);
nor U4151 (N_4151,In_597,In_2753);
xor U4152 (N_4152,In_2645,In_2604);
xor U4153 (N_4153,In_5,In_1191);
and U4154 (N_4154,In_1440,In_679);
nor U4155 (N_4155,In_1796,In_2530);
or U4156 (N_4156,In_243,In_2140);
nor U4157 (N_4157,In_1533,In_2604);
or U4158 (N_4158,In_1831,In_931);
nand U4159 (N_4159,In_1284,In_1871);
or U4160 (N_4160,In_402,In_2968);
or U4161 (N_4161,In_82,In_1376);
and U4162 (N_4162,In_1970,In_2082);
and U4163 (N_4163,In_2599,In_1105);
or U4164 (N_4164,In_24,In_893);
nor U4165 (N_4165,In_421,In_2254);
or U4166 (N_4166,In_148,In_363);
and U4167 (N_4167,In_2527,In_345);
nand U4168 (N_4168,In_1468,In_2781);
nor U4169 (N_4169,In_469,In_2095);
or U4170 (N_4170,In_2022,In_121);
and U4171 (N_4171,In_1388,In_1026);
and U4172 (N_4172,In_1156,In_1361);
and U4173 (N_4173,In_1971,In_1531);
and U4174 (N_4174,In_1209,In_643);
nand U4175 (N_4175,In_189,In_2275);
nor U4176 (N_4176,In_2581,In_2248);
nand U4177 (N_4177,In_344,In_2816);
or U4178 (N_4178,In_2348,In_526);
or U4179 (N_4179,In_681,In_2936);
nor U4180 (N_4180,In_1260,In_366);
nand U4181 (N_4181,In_2351,In_2830);
or U4182 (N_4182,In_2600,In_1305);
nand U4183 (N_4183,In_2025,In_461);
nor U4184 (N_4184,In_2399,In_592);
and U4185 (N_4185,In_2790,In_592);
nand U4186 (N_4186,In_382,In_2893);
nor U4187 (N_4187,In_105,In_110);
and U4188 (N_4188,In_2522,In_1066);
and U4189 (N_4189,In_2549,In_1899);
nor U4190 (N_4190,In_2674,In_2340);
xor U4191 (N_4191,In_2283,In_2930);
nor U4192 (N_4192,In_489,In_2261);
and U4193 (N_4193,In_2325,In_294);
nor U4194 (N_4194,In_497,In_2988);
and U4195 (N_4195,In_2029,In_1913);
and U4196 (N_4196,In_728,In_2600);
nor U4197 (N_4197,In_2861,In_294);
or U4198 (N_4198,In_29,In_388);
xor U4199 (N_4199,In_577,In_1469);
nor U4200 (N_4200,In_933,In_1556);
or U4201 (N_4201,In_2030,In_74);
nor U4202 (N_4202,In_1476,In_714);
and U4203 (N_4203,In_1200,In_2018);
nor U4204 (N_4204,In_2260,In_1910);
nand U4205 (N_4205,In_2435,In_2199);
or U4206 (N_4206,In_1240,In_11);
nor U4207 (N_4207,In_2834,In_2420);
nor U4208 (N_4208,In_1152,In_2143);
and U4209 (N_4209,In_1309,In_2771);
or U4210 (N_4210,In_1256,In_1629);
and U4211 (N_4211,In_2961,In_100);
and U4212 (N_4212,In_2362,In_779);
nand U4213 (N_4213,In_1615,In_1854);
nand U4214 (N_4214,In_2197,In_2269);
nand U4215 (N_4215,In_45,In_1897);
nor U4216 (N_4216,In_2732,In_702);
nand U4217 (N_4217,In_1698,In_674);
nor U4218 (N_4218,In_514,In_2613);
nor U4219 (N_4219,In_610,In_525);
nor U4220 (N_4220,In_395,In_928);
or U4221 (N_4221,In_340,In_1258);
nand U4222 (N_4222,In_2082,In_681);
and U4223 (N_4223,In_887,In_745);
or U4224 (N_4224,In_1979,In_1408);
nand U4225 (N_4225,In_2559,In_472);
or U4226 (N_4226,In_1766,In_543);
nand U4227 (N_4227,In_1051,In_1229);
nor U4228 (N_4228,In_788,In_2385);
nand U4229 (N_4229,In_210,In_1528);
nand U4230 (N_4230,In_1120,In_2390);
nor U4231 (N_4231,In_1835,In_2504);
nor U4232 (N_4232,In_1184,In_385);
or U4233 (N_4233,In_1054,In_812);
or U4234 (N_4234,In_2811,In_2075);
nand U4235 (N_4235,In_2820,In_2079);
nand U4236 (N_4236,In_332,In_1194);
xor U4237 (N_4237,In_2528,In_1530);
nor U4238 (N_4238,In_466,In_825);
and U4239 (N_4239,In_2448,In_584);
nand U4240 (N_4240,In_1852,In_801);
xor U4241 (N_4241,In_2120,In_1452);
nand U4242 (N_4242,In_197,In_1842);
or U4243 (N_4243,In_2164,In_998);
xor U4244 (N_4244,In_2271,In_2820);
and U4245 (N_4245,In_1696,In_1072);
nor U4246 (N_4246,In_2384,In_430);
and U4247 (N_4247,In_1663,In_2802);
nand U4248 (N_4248,In_2780,In_1399);
nand U4249 (N_4249,In_32,In_1326);
nand U4250 (N_4250,In_2810,In_758);
xnor U4251 (N_4251,In_1149,In_284);
and U4252 (N_4252,In_1335,In_820);
nor U4253 (N_4253,In_1432,In_879);
nand U4254 (N_4254,In_1476,In_358);
nor U4255 (N_4255,In_8,In_2697);
nand U4256 (N_4256,In_2141,In_426);
xor U4257 (N_4257,In_331,In_1649);
nor U4258 (N_4258,In_1457,In_2588);
and U4259 (N_4259,In_1458,In_284);
nor U4260 (N_4260,In_1415,In_2723);
nor U4261 (N_4261,In_625,In_1512);
and U4262 (N_4262,In_2797,In_1790);
nor U4263 (N_4263,In_2115,In_1799);
and U4264 (N_4264,In_2582,In_534);
or U4265 (N_4265,In_481,In_1218);
nor U4266 (N_4266,In_941,In_2898);
nand U4267 (N_4267,In_890,In_2236);
xor U4268 (N_4268,In_503,In_305);
and U4269 (N_4269,In_1349,In_380);
or U4270 (N_4270,In_2988,In_181);
nand U4271 (N_4271,In_48,In_2967);
nor U4272 (N_4272,In_1097,In_4);
and U4273 (N_4273,In_385,In_355);
nand U4274 (N_4274,In_269,In_713);
or U4275 (N_4275,In_2256,In_2880);
nor U4276 (N_4276,In_2021,In_2217);
nand U4277 (N_4277,In_2410,In_1032);
xor U4278 (N_4278,In_1506,In_451);
or U4279 (N_4279,In_316,In_604);
and U4280 (N_4280,In_2540,In_37);
and U4281 (N_4281,In_1188,In_172);
nor U4282 (N_4282,In_1184,In_555);
nor U4283 (N_4283,In_1408,In_2563);
nand U4284 (N_4284,In_2743,In_2526);
and U4285 (N_4285,In_108,In_935);
and U4286 (N_4286,In_2157,In_2353);
nor U4287 (N_4287,In_2202,In_925);
nand U4288 (N_4288,In_2682,In_396);
and U4289 (N_4289,In_131,In_134);
and U4290 (N_4290,In_1203,In_688);
nand U4291 (N_4291,In_1902,In_2721);
nand U4292 (N_4292,In_2970,In_1813);
nand U4293 (N_4293,In_2599,In_1920);
nor U4294 (N_4294,In_1909,In_246);
or U4295 (N_4295,In_2682,In_2846);
nand U4296 (N_4296,In_2082,In_285);
xnor U4297 (N_4297,In_819,In_2889);
nor U4298 (N_4298,In_643,In_1447);
nand U4299 (N_4299,In_449,In_2029);
nand U4300 (N_4300,In_214,In_327);
nand U4301 (N_4301,In_2552,In_2098);
nand U4302 (N_4302,In_2156,In_2402);
and U4303 (N_4303,In_848,In_1279);
or U4304 (N_4304,In_331,In_928);
nand U4305 (N_4305,In_217,In_362);
nor U4306 (N_4306,In_2633,In_1690);
nor U4307 (N_4307,In_2004,In_1016);
or U4308 (N_4308,In_1233,In_1699);
nor U4309 (N_4309,In_2549,In_295);
nand U4310 (N_4310,In_2734,In_1268);
nor U4311 (N_4311,In_2918,In_2573);
nand U4312 (N_4312,In_1928,In_1626);
nand U4313 (N_4313,In_1226,In_2960);
and U4314 (N_4314,In_1024,In_1876);
or U4315 (N_4315,In_2823,In_722);
xnor U4316 (N_4316,In_850,In_705);
and U4317 (N_4317,In_1273,In_2083);
nand U4318 (N_4318,In_1115,In_2087);
nor U4319 (N_4319,In_2210,In_2263);
xnor U4320 (N_4320,In_218,In_705);
and U4321 (N_4321,In_1820,In_1785);
and U4322 (N_4322,In_170,In_345);
nor U4323 (N_4323,In_1234,In_1869);
or U4324 (N_4324,In_2405,In_1755);
nor U4325 (N_4325,In_1309,In_974);
xor U4326 (N_4326,In_2791,In_2602);
and U4327 (N_4327,In_1601,In_2315);
and U4328 (N_4328,In_1527,In_585);
xor U4329 (N_4329,In_2439,In_1770);
nor U4330 (N_4330,In_2003,In_1444);
or U4331 (N_4331,In_1778,In_1949);
xnor U4332 (N_4332,In_1912,In_423);
or U4333 (N_4333,In_25,In_2476);
and U4334 (N_4334,In_2403,In_1652);
nand U4335 (N_4335,In_1809,In_1099);
and U4336 (N_4336,In_99,In_113);
or U4337 (N_4337,In_1719,In_880);
and U4338 (N_4338,In_1182,In_378);
nor U4339 (N_4339,In_558,In_1676);
or U4340 (N_4340,In_470,In_782);
and U4341 (N_4341,In_2589,In_2923);
or U4342 (N_4342,In_2674,In_1856);
nand U4343 (N_4343,In_716,In_2888);
and U4344 (N_4344,In_2144,In_687);
nand U4345 (N_4345,In_916,In_991);
and U4346 (N_4346,In_459,In_2658);
nor U4347 (N_4347,In_121,In_1553);
or U4348 (N_4348,In_352,In_1496);
or U4349 (N_4349,In_1249,In_751);
or U4350 (N_4350,In_2756,In_2080);
or U4351 (N_4351,In_2404,In_2029);
and U4352 (N_4352,In_901,In_772);
or U4353 (N_4353,In_1762,In_2292);
nand U4354 (N_4354,In_1838,In_22);
and U4355 (N_4355,In_2441,In_2923);
and U4356 (N_4356,In_733,In_2452);
nand U4357 (N_4357,In_696,In_2447);
and U4358 (N_4358,In_900,In_119);
and U4359 (N_4359,In_746,In_805);
nor U4360 (N_4360,In_1578,In_740);
or U4361 (N_4361,In_197,In_1978);
nor U4362 (N_4362,In_1078,In_705);
nor U4363 (N_4363,In_2197,In_1121);
nor U4364 (N_4364,In_1298,In_1879);
nor U4365 (N_4365,In_103,In_2998);
or U4366 (N_4366,In_844,In_1557);
nand U4367 (N_4367,In_2404,In_598);
and U4368 (N_4368,In_427,In_739);
or U4369 (N_4369,In_843,In_797);
and U4370 (N_4370,In_591,In_2006);
or U4371 (N_4371,In_966,In_1983);
nor U4372 (N_4372,In_1227,In_1939);
nand U4373 (N_4373,In_569,In_2741);
xor U4374 (N_4374,In_2448,In_505);
nor U4375 (N_4375,In_2601,In_1149);
nor U4376 (N_4376,In_2266,In_1055);
and U4377 (N_4377,In_662,In_131);
and U4378 (N_4378,In_468,In_2638);
and U4379 (N_4379,In_2566,In_1076);
nand U4380 (N_4380,In_1502,In_379);
nand U4381 (N_4381,In_1280,In_260);
or U4382 (N_4382,In_392,In_283);
nand U4383 (N_4383,In_519,In_2105);
or U4384 (N_4384,In_1379,In_1278);
xor U4385 (N_4385,In_610,In_2034);
nand U4386 (N_4386,In_1032,In_2704);
xor U4387 (N_4387,In_1982,In_2485);
and U4388 (N_4388,In_493,In_2904);
and U4389 (N_4389,In_2749,In_2700);
nor U4390 (N_4390,In_133,In_804);
or U4391 (N_4391,In_990,In_1605);
or U4392 (N_4392,In_0,In_2969);
nor U4393 (N_4393,In_1752,In_1082);
nor U4394 (N_4394,In_1298,In_888);
or U4395 (N_4395,In_2660,In_612);
or U4396 (N_4396,In_2245,In_1904);
and U4397 (N_4397,In_2633,In_1773);
or U4398 (N_4398,In_2402,In_1421);
nand U4399 (N_4399,In_2637,In_679);
or U4400 (N_4400,In_2719,In_2411);
or U4401 (N_4401,In_2031,In_2033);
or U4402 (N_4402,In_935,In_1360);
nand U4403 (N_4403,In_116,In_1713);
or U4404 (N_4404,In_241,In_1537);
nand U4405 (N_4405,In_514,In_1694);
nor U4406 (N_4406,In_844,In_365);
xnor U4407 (N_4407,In_1981,In_119);
or U4408 (N_4408,In_237,In_283);
and U4409 (N_4409,In_377,In_1820);
and U4410 (N_4410,In_851,In_2268);
nand U4411 (N_4411,In_1402,In_1039);
xor U4412 (N_4412,In_962,In_1826);
and U4413 (N_4413,In_2262,In_2796);
or U4414 (N_4414,In_2687,In_2017);
and U4415 (N_4415,In_2904,In_2462);
nand U4416 (N_4416,In_792,In_2886);
xor U4417 (N_4417,In_2034,In_1177);
nor U4418 (N_4418,In_1117,In_2145);
or U4419 (N_4419,In_2860,In_999);
nor U4420 (N_4420,In_442,In_463);
and U4421 (N_4421,In_1876,In_1291);
and U4422 (N_4422,In_2291,In_1395);
nor U4423 (N_4423,In_45,In_1481);
and U4424 (N_4424,In_1017,In_505);
and U4425 (N_4425,In_2237,In_2427);
nor U4426 (N_4426,In_1365,In_2136);
and U4427 (N_4427,In_1613,In_2978);
or U4428 (N_4428,In_1287,In_2871);
or U4429 (N_4429,In_2709,In_2749);
and U4430 (N_4430,In_1203,In_90);
or U4431 (N_4431,In_593,In_58);
or U4432 (N_4432,In_1115,In_1089);
and U4433 (N_4433,In_2489,In_1583);
nor U4434 (N_4434,In_43,In_1307);
or U4435 (N_4435,In_267,In_2290);
nor U4436 (N_4436,In_1883,In_544);
nand U4437 (N_4437,In_2771,In_2289);
nor U4438 (N_4438,In_2205,In_2093);
nor U4439 (N_4439,In_1125,In_2544);
nor U4440 (N_4440,In_871,In_1978);
nand U4441 (N_4441,In_54,In_1941);
nor U4442 (N_4442,In_2154,In_399);
or U4443 (N_4443,In_895,In_1480);
nand U4444 (N_4444,In_400,In_2741);
or U4445 (N_4445,In_2659,In_549);
and U4446 (N_4446,In_195,In_1700);
or U4447 (N_4447,In_666,In_2644);
nand U4448 (N_4448,In_252,In_439);
nand U4449 (N_4449,In_1464,In_1730);
nor U4450 (N_4450,In_2772,In_1515);
nor U4451 (N_4451,In_2949,In_189);
nor U4452 (N_4452,In_2049,In_2883);
or U4453 (N_4453,In_1168,In_2368);
and U4454 (N_4454,In_2690,In_2333);
nand U4455 (N_4455,In_2643,In_1037);
nor U4456 (N_4456,In_635,In_2678);
nor U4457 (N_4457,In_919,In_689);
and U4458 (N_4458,In_2610,In_1345);
nor U4459 (N_4459,In_1974,In_407);
or U4460 (N_4460,In_1261,In_282);
and U4461 (N_4461,In_2371,In_1230);
or U4462 (N_4462,In_1851,In_2117);
and U4463 (N_4463,In_1978,In_1503);
or U4464 (N_4464,In_1932,In_2739);
nand U4465 (N_4465,In_919,In_176);
nor U4466 (N_4466,In_150,In_2081);
nand U4467 (N_4467,In_1625,In_2295);
nor U4468 (N_4468,In_2516,In_0);
or U4469 (N_4469,In_618,In_1188);
nand U4470 (N_4470,In_367,In_2420);
nand U4471 (N_4471,In_160,In_915);
or U4472 (N_4472,In_1688,In_2589);
xor U4473 (N_4473,In_1801,In_697);
or U4474 (N_4474,In_73,In_1432);
nor U4475 (N_4475,In_1327,In_1139);
and U4476 (N_4476,In_711,In_1299);
xnor U4477 (N_4477,In_2601,In_270);
nand U4478 (N_4478,In_979,In_167);
nor U4479 (N_4479,In_2555,In_1906);
or U4480 (N_4480,In_51,In_887);
and U4481 (N_4481,In_1383,In_1359);
nor U4482 (N_4482,In_806,In_2599);
nor U4483 (N_4483,In_1812,In_2327);
and U4484 (N_4484,In_2599,In_1164);
nand U4485 (N_4485,In_1157,In_197);
and U4486 (N_4486,In_1332,In_766);
nand U4487 (N_4487,In_1770,In_820);
or U4488 (N_4488,In_59,In_997);
nor U4489 (N_4489,In_740,In_675);
nor U4490 (N_4490,In_913,In_2671);
nand U4491 (N_4491,In_2297,In_401);
or U4492 (N_4492,In_138,In_799);
xor U4493 (N_4493,In_817,In_2706);
xnor U4494 (N_4494,In_129,In_814);
nor U4495 (N_4495,In_1640,In_2236);
or U4496 (N_4496,In_1804,In_288);
and U4497 (N_4497,In_1447,In_2663);
and U4498 (N_4498,In_1786,In_1673);
nand U4499 (N_4499,In_1796,In_2787);
or U4500 (N_4500,In_827,In_2715);
nand U4501 (N_4501,In_2033,In_2992);
or U4502 (N_4502,In_2634,In_1848);
and U4503 (N_4503,In_1108,In_567);
and U4504 (N_4504,In_2605,In_2331);
and U4505 (N_4505,In_2755,In_2823);
or U4506 (N_4506,In_588,In_902);
or U4507 (N_4507,In_2851,In_2273);
and U4508 (N_4508,In_1974,In_709);
nand U4509 (N_4509,In_2620,In_1748);
nor U4510 (N_4510,In_2352,In_1268);
nor U4511 (N_4511,In_1738,In_1162);
and U4512 (N_4512,In_1860,In_1902);
and U4513 (N_4513,In_1149,In_1356);
nand U4514 (N_4514,In_1383,In_555);
and U4515 (N_4515,In_1179,In_158);
xor U4516 (N_4516,In_1668,In_1255);
and U4517 (N_4517,In_305,In_1430);
and U4518 (N_4518,In_2278,In_1798);
or U4519 (N_4519,In_837,In_2163);
or U4520 (N_4520,In_58,In_1091);
nand U4521 (N_4521,In_160,In_1418);
nor U4522 (N_4522,In_917,In_2161);
or U4523 (N_4523,In_1720,In_2721);
nand U4524 (N_4524,In_1354,In_2917);
xor U4525 (N_4525,In_1916,In_1582);
xor U4526 (N_4526,In_2823,In_2288);
or U4527 (N_4527,In_1213,In_1397);
and U4528 (N_4528,In_1585,In_803);
or U4529 (N_4529,In_1074,In_2655);
nand U4530 (N_4530,In_755,In_534);
nand U4531 (N_4531,In_2868,In_2948);
nand U4532 (N_4532,In_826,In_456);
nand U4533 (N_4533,In_1895,In_1400);
or U4534 (N_4534,In_314,In_825);
nand U4535 (N_4535,In_1660,In_1675);
or U4536 (N_4536,In_2411,In_33);
xor U4537 (N_4537,In_930,In_1574);
nand U4538 (N_4538,In_2885,In_2530);
nand U4539 (N_4539,In_2326,In_793);
and U4540 (N_4540,In_33,In_2179);
xor U4541 (N_4541,In_1078,In_2670);
and U4542 (N_4542,In_1858,In_2859);
nor U4543 (N_4543,In_449,In_212);
nand U4544 (N_4544,In_1289,In_1125);
nand U4545 (N_4545,In_2194,In_823);
nand U4546 (N_4546,In_515,In_1424);
or U4547 (N_4547,In_2176,In_2596);
xor U4548 (N_4548,In_428,In_2138);
nand U4549 (N_4549,In_695,In_985);
and U4550 (N_4550,In_2055,In_188);
nor U4551 (N_4551,In_2421,In_644);
or U4552 (N_4552,In_1271,In_2568);
nand U4553 (N_4553,In_517,In_2147);
or U4554 (N_4554,In_4,In_1298);
xor U4555 (N_4555,In_2771,In_714);
and U4556 (N_4556,In_2374,In_377);
xnor U4557 (N_4557,In_1201,In_148);
and U4558 (N_4558,In_2102,In_2718);
and U4559 (N_4559,In_1750,In_48);
or U4560 (N_4560,In_2024,In_1806);
nand U4561 (N_4561,In_2801,In_1734);
nor U4562 (N_4562,In_358,In_124);
or U4563 (N_4563,In_2692,In_2577);
xnor U4564 (N_4564,In_2741,In_2213);
xor U4565 (N_4565,In_1545,In_400);
nand U4566 (N_4566,In_1690,In_157);
or U4567 (N_4567,In_2157,In_1009);
nand U4568 (N_4568,In_1178,In_2341);
or U4569 (N_4569,In_325,In_2863);
xor U4570 (N_4570,In_759,In_125);
nor U4571 (N_4571,In_239,In_2972);
xnor U4572 (N_4572,In_1306,In_1241);
xor U4573 (N_4573,In_914,In_586);
nor U4574 (N_4574,In_1849,In_1490);
or U4575 (N_4575,In_2477,In_465);
nor U4576 (N_4576,In_2275,In_2501);
nor U4577 (N_4577,In_2064,In_7);
or U4578 (N_4578,In_2657,In_1715);
nor U4579 (N_4579,In_2796,In_1191);
nor U4580 (N_4580,In_631,In_2497);
nor U4581 (N_4581,In_1869,In_1501);
xor U4582 (N_4582,In_494,In_1281);
nand U4583 (N_4583,In_2366,In_717);
nor U4584 (N_4584,In_333,In_213);
nand U4585 (N_4585,In_1127,In_566);
xnor U4586 (N_4586,In_71,In_2618);
nand U4587 (N_4587,In_1067,In_406);
or U4588 (N_4588,In_2388,In_137);
or U4589 (N_4589,In_2976,In_2066);
and U4590 (N_4590,In_1139,In_2181);
nand U4591 (N_4591,In_692,In_2074);
nor U4592 (N_4592,In_691,In_1341);
or U4593 (N_4593,In_1517,In_719);
nor U4594 (N_4594,In_1213,In_1339);
and U4595 (N_4595,In_2967,In_334);
and U4596 (N_4596,In_381,In_442);
and U4597 (N_4597,In_398,In_499);
nand U4598 (N_4598,In_772,In_409);
nand U4599 (N_4599,In_41,In_2749);
or U4600 (N_4600,In_1690,In_74);
nand U4601 (N_4601,In_2319,In_1263);
nand U4602 (N_4602,In_2172,In_164);
and U4603 (N_4603,In_151,In_2689);
nand U4604 (N_4604,In_427,In_1974);
nand U4605 (N_4605,In_1590,In_2394);
nor U4606 (N_4606,In_2034,In_257);
nand U4607 (N_4607,In_815,In_807);
or U4608 (N_4608,In_2625,In_1651);
nand U4609 (N_4609,In_2979,In_1698);
and U4610 (N_4610,In_1212,In_2044);
xnor U4611 (N_4611,In_852,In_1953);
xor U4612 (N_4612,In_1536,In_1902);
or U4613 (N_4613,In_1670,In_1496);
and U4614 (N_4614,In_1434,In_1671);
and U4615 (N_4615,In_2426,In_790);
or U4616 (N_4616,In_2249,In_1945);
nand U4617 (N_4617,In_1791,In_104);
nand U4618 (N_4618,In_2500,In_540);
nor U4619 (N_4619,In_1909,In_2440);
or U4620 (N_4620,In_1254,In_1521);
nand U4621 (N_4621,In_934,In_186);
nand U4622 (N_4622,In_2411,In_1224);
or U4623 (N_4623,In_286,In_2844);
and U4624 (N_4624,In_2505,In_786);
and U4625 (N_4625,In_254,In_1175);
nand U4626 (N_4626,In_2227,In_2750);
and U4627 (N_4627,In_1697,In_974);
nor U4628 (N_4628,In_2647,In_2336);
nor U4629 (N_4629,In_1224,In_1384);
nand U4630 (N_4630,In_1959,In_2885);
or U4631 (N_4631,In_2931,In_226);
nand U4632 (N_4632,In_1991,In_1895);
and U4633 (N_4633,In_2408,In_596);
or U4634 (N_4634,In_1776,In_736);
nor U4635 (N_4635,In_875,In_738);
and U4636 (N_4636,In_2962,In_860);
and U4637 (N_4637,In_2364,In_153);
nor U4638 (N_4638,In_2451,In_2971);
xor U4639 (N_4639,In_809,In_507);
nor U4640 (N_4640,In_2642,In_2344);
nand U4641 (N_4641,In_1397,In_2092);
and U4642 (N_4642,In_22,In_114);
xor U4643 (N_4643,In_926,In_1569);
xor U4644 (N_4644,In_868,In_1894);
or U4645 (N_4645,In_2832,In_838);
or U4646 (N_4646,In_2294,In_896);
nor U4647 (N_4647,In_2028,In_2166);
and U4648 (N_4648,In_2474,In_2780);
and U4649 (N_4649,In_2911,In_2795);
nor U4650 (N_4650,In_126,In_2527);
nand U4651 (N_4651,In_454,In_497);
xnor U4652 (N_4652,In_2772,In_192);
nor U4653 (N_4653,In_1292,In_1502);
or U4654 (N_4654,In_2327,In_2483);
nor U4655 (N_4655,In_1191,In_1328);
nor U4656 (N_4656,In_2146,In_495);
nor U4657 (N_4657,In_1234,In_2945);
nand U4658 (N_4658,In_1471,In_103);
or U4659 (N_4659,In_494,In_412);
xnor U4660 (N_4660,In_2786,In_2092);
nor U4661 (N_4661,In_1635,In_1840);
nand U4662 (N_4662,In_509,In_282);
and U4663 (N_4663,In_1275,In_2188);
and U4664 (N_4664,In_2495,In_2491);
nor U4665 (N_4665,In_1811,In_949);
xnor U4666 (N_4666,In_1605,In_1233);
nand U4667 (N_4667,In_652,In_1156);
nor U4668 (N_4668,In_2938,In_1048);
nand U4669 (N_4669,In_992,In_1992);
nand U4670 (N_4670,In_1090,In_1012);
or U4671 (N_4671,In_508,In_2556);
xor U4672 (N_4672,In_2054,In_233);
and U4673 (N_4673,In_2883,In_138);
nand U4674 (N_4674,In_1732,In_981);
nor U4675 (N_4675,In_2050,In_1465);
nand U4676 (N_4676,In_1156,In_1929);
and U4677 (N_4677,In_1059,In_2878);
or U4678 (N_4678,In_2325,In_1309);
nor U4679 (N_4679,In_447,In_2154);
and U4680 (N_4680,In_1444,In_887);
nor U4681 (N_4681,In_2651,In_2773);
and U4682 (N_4682,In_520,In_1094);
or U4683 (N_4683,In_1715,In_1308);
nor U4684 (N_4684,In_2378,In_734);
or U4685 (N_4685,In_1896,In_1279);
or U4686 (N_4686,In_2820,In_1477);
nor U4687 (N_4687,In_1210,In_225);
xor U4688 (N_4688,In_2033,In_1358);
and U4689 (N_4689,In_179,In_67);
nor U4690 (N_4690,In_1381,In_2353);
or U4691 (N_4691,In_2197,In_2704);
nand U4692 (N_4692,In_2198,In_2938);
nor U4693 (N_4693,In_1459,In_1405);
and U4694 (N_4694,In_724,In_1138);
and U4695 (N_4695,In_526,In_643);
and U4696 (N_4696,In_2577,In_1241);
nand U4697 (N_4697,In_1549,In_2460);
nor U4698 (N_4698,In_2061,In_1654);
and U4699 (N_4699,In_2296,In_2213);
nand U4700 (N_4700,In_332,In_1872);
nand U4701 (N_4701,In_2029,In_1959);
nand U4702 (N_4702,In_1028,In_1226);
xnor U4703 (N_4703,In_1014,In_2842);
nor U4704 (N_4704,In_788,In_147);
or U4705 (N_4705,In_2105,In_853);
or U4706 (N_4706,In_1680,In_2957);
xnor U4707 (N_4707,In_2162,In_1053);
or U4708 (N_4708,In_189,In_428);
or U4709 (N_4709,In_399,In_1989);
nor U4710 (N_4710,In_151,In_2368);
nor U4711 (N_4711,In_2048,In_2770);
nand U4712 (N_4712,In_17,In_1923);
nor U4713 (N_4713,In_2724,In_1261);
nand U4714 (N_4714,In_838,In_2849);
or U4715 (N_4715,In_1503,In_798);
nor U4716 (N_4716,In_2669,In_650);
or U4717 (N_4717,In_2794,In_295);
and U4718 (N_4718,In_1435,In_1478);
and U4719 (N_4719,In_2530,In_1945);
and U4720 (N_4720,In_2766,In_304);
or U4721 (N_4721,In_2750,In_1561);
and U4722 (N_4722,In_2142,In_355);
and U4723 (N_4723,In_1726,In_2306);
nor U4724 (N_4724,In_1051,In_1940);
and U4725 (N_4725,In_994,In_1839);
or U4726 (N_4726,In_2133,In_2400);
or U4727 (N_4727,In_1110,In_2277);
and U4728 (N_4728,In_1687,In_405);
or U4729 (N_4729,In_783,In_273);
xnor U4730 (N_4730,In_2616,In_2636);
or U4731 (N_4731,In_1463,In_729);
nand U4732 (N_4732,In_1178,In_2084);
nor U4733 (N_4733,In_320,In_2262);
or U4734 (N_4734,In_676,In_684);
nor U4735 (N_4735,In_1665,In_1925);
nor U4736 (N_4736,In_461,In_1469);
nor U4737 (N_4737,In_892,In_1533);
nor U4738 (N_4738,In_22,In_713);
and U4739 (N_4739,In_977,In_119);
nand U4740 (N_4740,In_2299,In_1926);
or U4741 (N_4741,In_1667,In_425);
nand U4742 (N_4742,In_2178,In_2905);
and U4743 (N_4743,In_2592,In_339);
nand U4744 (N_4744,In_399,In_2533);
or U4745 (N_4745,In_1069,In_1022);
nor U4746 (N_4746,In_711,In_1760);
nor U4747 (N_4747,In_2566,In_399);
and U4748 (N_4748,In_767,In_606);
nor U4749 (N_4749,In_2700,In_574);
and U4750 (N_4750,In_2321,In_986);
or U4751 (N_4751,In_2939,In_1376);
and U4752 (N_4752,In_2319,In_2371);
and U4753 (N_4753,In_2872,In_558);
nor U4754 (N_4754,In_996,In_1567);
and U4755 (N_4755,In_466,In_2601);
and U4756 (N_4756,In_999,In_2871);
nor U4757 (N_4757,In_1641,In_1061);
or U4758 (N_4758,In_2609,In_2733);
or U4759 (N_4759,In_1386,In_2656);
xnor U4760 (N_4760,In_325,In_2876);
nand U4761 (N_4761,In_675,In_1585);
or U4762 (N_4762,In_1996,In_2332);
or U4763 (N_4763,In_1343,In_2462);
or U4764 (N_4764,In_208,In_1079);
nand U4765 (N_4765,In_2172,In_1213);
and U4766 (N_4766,In_2735,In_2325);
or U4767 (N_4767,In_1712,In_1833);
xnor U4768 (N_4768,In_1972,In_2326);
nor U4769 (N_4769,In_1624,In_2376);
nand U4770 (N_4770,In_2121,In_1119);
nand U4771 (N_4771,In_555,In_1049);
nor U4772 (N_4772,In_1893,In_1120);
nor U4773 (N_4773,In_1867,In_1891);
nand U4774 (N_4774,In_1787,In_2303);
nand U4775 (N_4775,In_2370,In_2359);
nor U4776 (N_4776,In_1,In_357);
and U4777 (N_4777,In_2828,In_246);
nor U4778 (N_4778,In_2161,In_2729);
nand U4779 (N_4779,In_504,In_1856);
xor U4780 (N_4780,In_126,In_1461);
nor U4781 (N_4781,In_1298,In_2920);
nand U4782 (N_4782,In_1471,In_1394);
nand U4783 (N_4783,In_957,In_1623);
and U4784 (N_4784,In_284,In_2488);
nor U4785 (N_4785,In_524,In_30);
and U4786 (N_4786,In_2513,In_493);
nand U4787 (N_4787,In_563,In_1065);
nor U4788 (N_4788,In_2218,In_1582);
and U4789 (N_4789,In_2171,In_2690);
nor U4790 (N_4790,In_2983,In_2211);
nor U4791 (N_4791,In_1404,In_2645);
nor U4792 (N_4792,In_1191,In_1239);
and U4793 (N_4793,In_2709,In_1312);
and U4794 (N_4794,In_1091,In_1269);
or U4795 (N_4795,In_398,In_2447);
nand U4796 (N_4796,In_1248,In_656);
nor U4797 (N_4797,In_1154,In_2780);
or U4798 (N_4798,In_1971,In_100);
nor U4799 (N_4799,In_1009,In_2885);
and U4800 (N_4800,In_2969,In_1518);
or U4801 (N_4801,In_1647,In_2363);
nor U4802 (N_4802,In_2343,In_2233);
nor U4803 (N_4803,In_996,In_962);
or U4804 (N_4804,In_2871,In_1966);
and U4805 (N_4805,In_1768,In_1103);
xor U4806 (N_4806,In_2835,In_1025);
or U4807 (N_4807,In_1346,In_1913);
and U4808 (N_4808,In_897,In_1745);
nand U4809 (N_4809,In_2403,In_2187);
nand U4810 (N_4810,In_470,In_1229);
and U4811 (N_4811,In_2063,In_516);
nand U4812 (N_4812,In_913,In_1506);
and U4813 (N_4813,In_371,In_809);
nand U4814 (N_4814,In_1297,In_1561);
nor U4815 (N_4815,In_1251,In_2415);
nand U4816 (N_4816,In_2962,In_2596);
or U4817 (N_4817,In_2111,In_2751);
nand U4818 (N_4818,In_229,In_2778);
or U4819 (N_4819,In_1984,In_1407);
xnor U4820 (N_4820,In_2069,In_1908);
nand U4821 (N_4821,In_763,In_1844);
and U4822 (N_4822,In_1903,In_776);
or U4823 (N_4823,In_2013,In_2668);
or U4824 (N_4824,In_811,In_1488);
and U4825 (N_4825,In_1221,In_2043);
xor U4826 (N_4826,In_2540,In_2927);
nand U4827 (N_4827,In_674,In_565);
nor U4828 (N_4828,In_1162,In_1398);
and U4829 (N_4829,In_2731,In_747);
or U4830 (N_4830,In_19,In_606);
nor U4831 (N_4831,In_1193,In_502);
and U4832 (N_4832,In_1344,In_1536);
xnor U4833 (N_4833,In_823,In_2645);
nor U4834 (N_4834,In_1933,In_1526);
nor U4835 (N_4835,In_2197,In_720);
nor U4836 (N_4836,In_122,In_2243);
nor U4837 (N_4837,In_2269,In_996);
or U4838 (N_4838,In_2885,In_2874);
nand U4839 (N_4839,In_1271,In_317);
nor U4840 (N_4840,In_2945,In_1352);
xor U4841 (N_4841,In_1307,In_1401);
or U4842 (N_4842,In_1775,In_2064);
and U4843 (N_4843,In_2329,In_2510);
and U4844 (N_4844,In_1681,In_1070);
and U4845 (N_4845,In_1181,In_1235);
nand U4846 (N_4846,In_2169,In_2677);
or U4847 (N_4847,In_1682,In_2735);
nand U4848 (N_4848,In_189,In_634);
and U4849 (N_4849,In_1248,In_2770);
and U4850 (N_4850,In_767,In_226);
nand U4851 (N_4851,In_1440,In_1173);
or U4852 (N_4852,In_2741,In_174);
nor U4853 (N_4853,In_831,In_1671);
nor U4854 (N_4854,In_932,In_856);
xor U4855 (N_4855,In_1267,In_1870);
xnor U4856 (N_4856,In_1914,In_986);
or U4857 (N_4857,In_1927,In_92);
and U4858 (N_4858,In_2837,In_2402);
nand U4859 (N_4859,In_2654,In_1292);
nor U4860 (N_4860,In_1323,In_887);
nor U4861 (N_4861,In_2930,In_1519);
and U4862 (N_4862,In_2311,In_2211);
xor U4863 (N_4863,In_49,In_2014);
and U4864 (N_4864,In_2672,In_2928);
and U4865 (N_4865,In_1457,In_2878);
or U4866 (N_4866,In_2229,In_1168);
nand U4867 (N_4867,In_189,In_1681);
or U4868 (N_4868,In_754,In_2659);
nand U4869 (N_4869,In_1601,In_2850);
nand U4870 (N_4870,In_794,In_1100);
nor U4871 (N_4871,In_422,In_28);
nor U4872 (N_4872,In_769,In_313);
and U4873 (N_4873,In_2955,In_212);
and U4874 (N_4874,In_1376,In_1013);
nand U4875 (N_4875,In_266,In_306);
nor U4876 (N_4876,In_1035,In_377);
and U4877 (N_4877,In_2648,In_2577);
or U4878 (N_4878,In_2193,In_8);
and U4879 (N_4879,In_684,In_1256);
and U4880 (N_4880,In_2434,In_1346);
nor U4881 (N_4881,In_1823,In_2472);
or U4882 (N_4882,In_1771,In_2091);
and U4883 (N_4883,In_753,In_1658);
and U4884 (N_4884,In_67,In_1053);
and U4885 (N_4885,In_2047,In_1521);
and U4886 (N_4886,In_1965,In_1825);
and U4887 (N_4887,In_2079,In_1987);
nand U4888 (N_4888,In_2247,In_2358);
nand U4889 (N_4889,In_1771,In_505);
nand U4890 (N_4890,In_2167,In_2606);
or U4891 (N_4891,In_1687,In_323);
xnor U4892 (N_4892,In_854,In_1207);
nor U4893 (N_4893,In_2967,In_1871);
or U4894 (N_4894,In_1510,In_103);
nand U4895 (N_4895,In_1802,In_2185);
and U4896 (N_4896,In_2310,In_166);
nor U4897 (N_4897,In_2113,In_2531);
and U4898 (N_4898,In_1543,In_1701);
nor U4899 (N_4899,In_1966,In_2663);
nand U4900 (N_4900,In_2963,In_2023);
and U4901 (N_4901,In_2030,In_302);
and U4902 (N_4902,In_284,In_2535);
nor U4903 (N_4903,In_2597,In_835);
nor U4904 (N_4904,In_933,In_2401);
nand U4905 (N_4905,In_2159,In_508);
nor U4906 (N_4906,In_1515,In_1186);
nand U4907 (N_4907,In_1612,In_1512);
or U4908 (N_4908,In_1688,In_1318);
and U4909 (N_4909,In_2250,In_539);
nand U4910 (N_4910,In_1493,In_272);
nor U4911 (N_4911,In_1667,In_557);
or U4912 (N_4912,In_2507,In_1643);
nor U4913 (N_4913,In_654,In_1199);
nand U4914 (N_4914,In_844,In_1168);
and U4915 (N_4915,In_725,In_2008);
or U4916 (N_4916,In_1611,In_841);
or U4917 (N_4917,In_2647,In_139);
and U4918 (N_4918,In_1066,In_1893);
nand U4919 (N_4919,In_1470,In_794);
nor U4920 (N_4920,In_2879,In_178);
and U4921 (N_4921,In_420,In_1885);
nor U4922 (N_4922,In_1922,In_339);
nor U4923 (N_4923,In_1133,In_2169);
and U4924 (N_4924,In_2930,In_2344);
or U4925 (N_4925,In_2567,In_1981);
and U4926 (N_4926,In_131,In_1474);
nand U4927 (N_4927,In_2538,In_126);
or U4928 (N_4928,In_903,In_2894);
nor U4929 (N_4929,In_595,In_1466);
nor U4930 (N_4930,In_1175,In_101);
nand U4931 (N_4931,In_1825,In_1661);
xor U4932 (N_4932,In_2269,In_230);
or U4933 (N_4933,In_1091,In_2023);
nor U4934 (N_4934,In_288,In_2266);
nand U4935 (N_4935,In_2867,In_353);
or U4936 (N_4936,In_1517,In_2722);
or U4937 (N_4937,In_390,In_681);
nor U4938 (N_4938,In_350,In_2264);
and U4939 (N_4939,In_1263,In_1280);
nor U4940 (N_4940,In_15,In_148);
and U4941 (N_4941,In_1809,In_1049);
or U4942 (N_4942,In_2288,In_258);
and U4943 (N_4943,In_2431,In_703);
xnor U4944 (N_4944,In_2938,In_741);
xor U4945 (N_4945,In_1692,In_2132);
and U4946 (N_4946,In_519,In_1964);
xor U4947 (N_4947,In_1979,In_2745);
xnor U4948 (N_4948,In_919,In_2197);
nand U4949 (N_4949,In_67,In_1874);
nand U4950 (N_4950,In_906,In_1011);
nor U4951 (N_4951,In_1972,In_1836);
nor U4952 (N_4952,In_1451,In_403);
and U4953 (N_4953,In_1977,In_1210);
nand U4954 (N_4954,In_1450,In_1931);
nand U4955 (N_4955,In_1169,In_137);
nand U4956 (N_4956,In_2352,In_1330);
nand U4957 (N_4957,In_57,In_1127);
and U4958 (N_4958,In_1066,In_986);
nand U4959 (N_4959,In_1322,In_2614);
or U4960 (N_4960,In_653,In_0);
or U4961 (N_4961,In_1508,In_2467);
nand U4962 (N_4962,In_832,In_24);
or U4963 (N_4963,In_1564,In_876);
or U4964 (N_4964,In_2366,In_66);
nand U4965 (N_4965,In_2618,In_2292);
nor U4966 (N_4966,In_1671,In_786);
or U4967 (N_4967,In_1540,In_2893);
nand U4968 (N_4968,In_1293,In_2483);
nand U4969 (N_4969,In_2405,In_1900);
and U4970 (N_4970,In_492,In_1365);
xnor U4971 (N_4971,In_737,In_2350);
nand U4972 (N_4972,In_110,In_2394);
nand U4973 (N_4973,In_322,In_2193);
nand U4974 (N_4974,In_1179,In_1656);
and U4975 (N_4975,In_2118,In_1154);
nor U4976 (N_4976,In_1540,In_2032);
or U4977 (N_4977,In_1807,In_1165);
nand U4978 (N_4978,In_2443,In_2627);
or U4979 (N_4979,In_1416,In_2156);
or U4980 (N_4980,In_1447,In_2381);
nor U4981 (N_4981,In_2019,In_477);
and U4982 (N_4982,In_2762,In_1439);
nor U4983 (N_4983,In_1585,In_770);
nor U4984 (N_4984,In_293,In_2349);
xor U4985 (N_4985,In_788,In_731);
and U4986 (N_4986,In_2662,In_1645);
nor U4987 (N_4987,In_170,In_2895);
nand U4988 (N_4988,In_2720,In_1774);
or U4989 (N_4989,In_444,In_237);
and U4990 (N_4990,In_2653,In_2159);
nand U4991 (N_4991,In_2213,In_2669);
nand U4992 (N_4992,In_1214,In_2487);
and U4993 (N_4993,In_358,In_1853);
or U4994 (N_4994,In_2283,In_1600);
or U4995 (N_4995,In_1852,In_2019);
nand U4996 (N_4996,In_1805,In_1459);
or U4997 (N_4997,In_2509,In_1844);
nand U4998 (N_4998,In_1607,In_1552);
and U4999 (N_4999,In_1845,In_2980);
nor U5000 (N_5000,N_238,N_2777);
xnor U5001 (N_5001,N_150,N_4495);
and U5002 (N_5002,N_74,N_1990);
nor U5003 (N_5003,N_3855,N_2240);
nor U5004 (N_5004,N_2960,N_2161);
and U5005 (N_5005,N_3453,N_3669);
or U5006 (N_5006,N_4548,N_947);
and U5007 (N_5007,N_2404,N_4456);
or U5008 (N_5008,N_580,N_1505);
nand U5009 (N_5009,N_1174,N_3745);
nand U5010 (N_5010,N_4022,N_1290);
nor U5011 (N_5011,N_1999,N_4887);
and U5012 (N_5012,N_4466,N_789);
or U5013 (N_5013,N_3771,N_3873);
nand U5014 (N_5014,N_1477,N_2130);
nor U5015 (N_5015,N_3552,N_4742);
and U5016 (N_5016,N_889,N_4347);
nor U5017 (N_5017,N_1099,N_4025);
or U5018 (N_5018,N_3235,N_4473);
nand U5019 (N_5019,N_1620,N_3211);
and U5020 (N_5020,N_1448,N_87);
nor U5021 (N_5021,N_3338,N_1413);
nor U5022 (N_5022,N_2,N_405);
nand U5023 (N_5023,N_1892,N_1901);
or U5024 (N_5024,N_1974,N_1707);
or U5025 (N_5025,N_1077,N_2359);
nor U5026 (N_5026,N_2854,N_1383);
and U5027 (N_5027,N_1617,N_983);
nand U5028 (N_5028,N_2050,N_3147);
nor U5029 (N_5029,N_641,N_3471);
nor U5030 (N_5030,N_4723,N_1557);
or U5031 (N_5031,N_4203,N_3094);
nand U5032 (N_5032,N_934,N_1754);
and U5033 (N_5033,N_831,N_3410);
nor U5034 (N_5034,N_463,N_3291);
nand U5035 (N_5035,N_1391,N_4610);
or U5036 (N_5036,N_3396,N_1865);
or U5037 (N_5037,N_2316,N_1381);
or U5038 (N_5038,N_921,N_1136);
or U5039 (N_5039,N_155,N_3017);
and U5040 (N_5040,N_1071,N_2298);
or U5041 (N_5041,N_2906,N_3937);
nor U5042 (N_5042,N_712,N_648);
and U5043 (N_5043,N_3934,N_3014);
or U5044 (N_5044,N_1926,N_1576);
and U5045 (N_5045,N_2734,N_1186);
or U5046 (N_5046,N_3616,N_3695);
nor U5047 (N_5047,N_1273,N_3899);
or U5048 (N_5048,N_4690,N_1335);
and U5049 (N_5049,N_2063,N_474);
or U5050 (N_5050,N_2141,N_1291);
and U5051 (N_5051,N_1514,N_1729);
and U5052 (N_5052,N_1217,N_3470);
and U5053 (N_5053,N_630,N_4844);
nand U5054 (N_5054,N_703,N_970);
and U5055 (N_5055,N_1629,N_2055);
and U5056 (N_5056,N_3778,N_117);
or U5057 (N_5057,N_795,N_3007);
nor U5058 (N_5058,N_1899,N_4178);
and U5059 (N_5059,N_2225,N_1386);
nor U5060 (N_5060,N_2422,N_4101);
and U5061 (N_5061,N_2746,N_3436);
or U5062 (N_5062,N_4926,N_2750);
or U5063 (N_5063,N_1327,N_683);
or U5064 (N_5064,N_2958,N_1221);
xor U5065 (N_5065,N_3395,N_1703);
and U5066 (N_5066,N_4241,N_1666);
or U5067 (N_5067,N_4269,N_215);
nor U5068 (N_5068,N_3943,N_2855);
nor U5069 (N_5069,N_1789,N_1472);
and U5070 (N_5070,N_179,N_2711);
nor U5071 (N_5071,N_3402,N_1758);
and U5072 (N_5072,N_1047,N_4807);
nor U5073 (N_5073,N_4051,N_3723);
and U5074 (N_5074,N_4044,N_3203);
or U5075 (N_5075,N_3596,N_2506);
xor U5076 (N_5076,N_3348,N_2226);
and U5077 (N_5077,N_1971,N_4502);
or U5078 (N_5078,N_1195,N_1496);
nor U5079 (N_5079,N_1839,N_2542);
nor U5080 (N_5080,N_1018,N_930);
nor U5081 (N_5081,N_444,N_239);
or U5082 (N_5082,N_2637,N_4881);
and U5083 (N_5083,N_633,N_543);
nor U5084 (N_5084,N_643,N_2816);
and U5085 (N_5085,N_4719,N_4527);
and U5086 (N_5086,N_450,N_2448);
xor U5087 (N_5087,N_385,N_3123);
or U5088 (N_5088,N_752,N_4820);
or U5089 (N_5089,N_1852,N_3859);
nand U5090 (N_5090,N_1346,N_1267);
or U5091 (N_5091,N_4970,N_692);
xor U5092 (N_5092,N_3202,N_4131);
or U5093 (N_5093,N_2527,N_993);
and U5094 (N_5094,N_3084,N_3566);
nor U5095 (N_5095,N_2718,N_4087);
nor U5096 (N_5096,N_2019,N_121);
or U5097 (N_5097,N_4383,N_2940);
and U5098 (N_5098,N_2454,N_70);
and U5099 (N_5099,N_3406,N_2307);
or U5100 (N_5100,N_3642,N_2852);
xnor U5101 (N_5101,N_1627,N_3274);
and U5102 (N_5102,N_307,N_2368);
or U5103 (N_5103,N_4315,N_659);
nand U5104 (N_5104,N_4000,N_2531);
and U5105 (N_5105,N_4598,N_2179);
and U5106 (N_5106,N_1821,N_3414);
or U5107 (N_5107,N_1203,N_1907);
and U5108 (N_5108,N_4179,N_2065);
nand U5109 (N_5109,N_4592,N_1139);
or U5110 (N_5110,N_4065,N_2467);
and U5111 (N_5111,N_1604,N_2492);
and U5112 (N_5112,N_2285,N_2670);
nand U5113 (N_5113,N_1919,N_3521);
nor U5114 (N_5114,N_3105,N_4954);
nor U5115 (N_5115,N_1495,N_4830);
nand U5116 (N_5116,N_613,N_1403);
nor U5117 (N_5117,N_25,N_4270);
nor U5118 (N_5118,N_3482,N_3843);
nor U5119 (N_5119,N_1605,N_4867);
or U5120 (N_5120,N_3854,N_1868);
and U5121 (N_5121,N_2710,N_60);
and U5122 (N_5122,N_3887,N_284);
nand U5123 (N_5123,N_3604,N_3823);
or U5124 (N_5124,N_2767,N_2132);
nor U5125 (N_5125,N_3961,N_1224);
and U5126 (N_5126,N_26,N_1694);
nor U5127 (N_5127,N_2614,N_422);
or U5128 (N_5128,N_3364,N_3038);
or U5129 (N_5129,N_3654,N_4666);
and U5130 (N_5130,N_3412,N_4721);
xnor U5131 (N_5131,N_4018,N_1841);
or U5132 (N_5132,N_2441,N_491);
or U5133 (N_5133,N_4083,N_2952);
nor U5134 (N_5134,N_913,N_1750);
nor U5135 (N_5135,N_4217,N_180);
nand U5136 (N_5136,N_2021,N_72);
nor U5137 (N_5137,N_2461,N_3583);
nor U5138 (N_5138,N_177,N_3045);
nand U5139 (N_5139,N_2231,N_3390);
or U5140 (N_5140,N_478,N_4019);
nor U5141 (N_5141,N_2624,N_1575);
nand U5142 (N_5142,N_527,N_1281);
nor U5143 (N_5143,N_4826,N_2210);
nor U5144 (N_5144,N_539,N_4906);
nand U5145 (N_5145,N_4584,N_4528);
and U5146 (N_5146,N_2214,N_4379);
and U5147 (N_5147,N_971,N_2831);
xor U5148 (N_5148,N_669,N_2223);
nand U5149 (N_5149,N_635,N_3064);
nand U5150 (N_5150,N_3181,N_1471);
nor U5151 (N_5151,N_4498,N_4378);
and U5152 (N_5152,N_3413,N_2388);
nor U5153 (N_5153,N_829,N_47);
nand U5154 (N_5154,N_1688,N_2679);
or U5155 (N_5155,N_340,N_1511);
or U5156 (N_5156,N_2269,N_3120);
and U5157 (N_5157,N_2337,N_3356);
or U5158 (N_5158,N_1051,N_1888);
nand U5159 (N_5159,N_3747,N_1902);
and U5160 (N_5160,N_2957,N_4869);
nand U5161 (N_5161,N_1458,N_2053);
nand U5162 (N_5162,N_4218,N_287);
nand U5163 (N_5163,N_1669,N_479);
nor U5164 (N_5164,N_3391,N_3861);
nor U5165 (N_5165,N_547,N_2631);
or U5166 (N_5166,N_3144,N_420);
nand U5167 (N_5167,N_2197,N_4306);
nand U5168 (N_5168,N_3688,N_4095);
or U5169 (N_5169,N_2686,N_476);
and U5170 (N_5170,N_3136,N_3459);
or U5171 (N_5171,N_4901,N_3733);
nand U5172 (N_5172,N_4911,N_251);
nand U5173 (N_5173,N_3044,N_732);
nand U5174 (N_5174,N_1998,N_3025);
nand U5175 (N_5175,N_1583,N_1460);
or U5176 (N_5176,N_326,N_4432);
nand U5177 (N_5177,N_4030,N_3739);
and U5178 (N_5178,N_345,N_1134);
nand U5179 (N_5179,N_1776,N_3568);
or U5180 (N_5180,N_745,N_1987);
nor U5181 (N_5181,N_3306,N_2829);
or U5182 (N_5182,N_4920,N_2083);
nand U5183 (N_5183,N_2523,N_4145);
and U5184 (N_5184,N_3134,N_3193);
or U5185 (N_5185,N_4789,N_1096);
nor U5186 (N_5186,N_4801,N_438);
xor U5187 (N_5187,N_2724,N_520);
or U5188 (N_5188,N_974,N_4727);
and U5189 (N_5189,N_4490,N_3247);
and U5190 (N_5190,N_556,N_1793);
or U5191 (N_5191,N_3290,N_4258);
xnor U5192 (N_5192,N_1469,N_1979);
xnor U5193 (N_5193,N_4056,N_226);
nor U5194 (N_5194,N_38,N_246);
nand U5195 (N_5195,N_2970,N_1023);
nor U5196 (N_5196,N_1034,N_4272);
or U5197 (N_5197,N_2294,N_1531);
or U5198 (N_5198,N_3791,N_1442);
nand U5199 (N_5199,N_4447,N_3539);
xnor U5200 (N_5200,N_440,N_3909);
nand U5201 (N_5201,N_595,N_24);
xnor U5202 (N_5202,N_3848,N_4851);
and U5203 (N_5203,N_4791,N_877);
xnor U5204 (N_5204,N_4261,N_2607);
nor U5205 (N_5205,N_3154,N_574);
nand U5206 (N_5206,N_3982,N_3159);
or U5207 (N_5207,N_3085,N_2039);
xor U5208 (N_5208,N_4591,N_1059);
or U5209 (N_5209,N_2856,N_3576);
nor U5210 (N_5210,N_571,N_2348);
xor U5211 (N_5211,N_1851,N_1169);
nor U5212 (N_5212,N_3016,N_780);
and U5213 (N_5213,N_548,N_408);
or U5214 (N_5214,N_1570,N_4698);
xor U5215 (N_5215,N_2598,N_3834);
or U5216 (N_5216,N_2204,N_2097);
and U5217 (N_5217,N_576,N_4989);
or U5218 (N_5218,N_3927,N_1211);
or U5219 (N_5219,N_189,N_1184);
and U5220 (N_5220,N_4641,N_4012);
or U5221 (N_5221,N_1352,N_4945);
nand U5222 (N_5222,N_4084,N_4667);
or U5223 (N_5223,N_1615,N_2255);
or U5224 (N_5224,N_1866,N_699);
nor U5225 (N_5225,N_2364,N_4219);
nand U5226 (N_5226,N_404,N_4180);
and U5227 (N_5227,N_1972,N_1554);
and U5228 (N_5228,N_2375,N_3868);
xnor U5229 (N_5229,N_174,N_3199);
or U5230 (N_5230,N_1479,N_3169);
or U5231 (N_5231,N_1407,N_710);
and U5232 (N_5232,N_3703,N_2478);
and U5233 (N_5233,N_288,N_4171);
nand U5234 (N_5234,N_3884,N_2773);
nor U5235 (N_5235,N_2923,N_66);
nor U5236 (N_5236,N_4054,N_1056);
nand U5237 (N_5237,N_4784,N_1229);
xor U5238 (N_5238,N_280,N_1264);
or U5239 (N_5239,N_3667,N_4023);
xnor U5240 (N_5240,N_4385,N_2213);
and U5241 (N_5241,N_2626,N_494);
or U5242 (N_5242,N_2653,N_3630);
or U5243 (N_5243,N_1968,N_868);
or U5244 (N_5244,N_335,N_3842);
nand U5245 (N_5245,N_3832,N_2826);
or U5246 (N_5246,N_3644,N_3717);
nand U5247 (N_5247,N_2172,N_4366);
and U5248 (N_5248,N_1643,N_20);
xnor U5249 (N_5249,N_1539,N_2191);
xor U5250 (N_5250,N_4015,N_1263);
nor U5251 (N_5251,N_636,N_859);
and U5252 (N_5252,N_1146,N_4158);
nor U5253 (N_5253,N_1421,N_862);
nand U5254 (N_5254,N_689,N_2599);
and U5255 (N_5255,N_461,N_3115);
or U5256 (N_5256,N_2124,N_1510);
nand U5257 (N_5257,N_101,N_267);
xor U5258 (N_5258,N_826,N_4156);
nor U5259 (N_5259,N_4511,N_4799);
xnor U5260 (N_5260,N_3359,N_3003);
and U5261 (N_5261,N_3598,N_456);
nor U5262 (N_5262,N_3039,N_4988);
and U5263 (N_5263,N_1395,N_65);
or U5264 (N_5264,N_260,N_1220);
or U5265 (N_5265,N_3592,N_2028);
nand U5266 (N_5266,N_2980,N_4738);
and U5267 (N_5267,N_757,N_3789);
and U5268 (N_5268,N_4759,N_4505);
or U5269 (N_5269,N_4750,N_979);
xor U5270 (N_5270,N_2801,N_902);
nor U5271 (N_5271,N_841,N_4872);
and U5272 (N_5272,N_4835,N_3300);
xor U5273 (N_5273,N_4333,N_2840);
nor U5274 (N_5274,N_4724,N_1553);
or U5275 (N_5275,N_1388,N_1131);
xnor U5276 (N_5276,N_52,N_3536);
nor U5277 (N_5277,N_235,N_2592);
or U5278 (N_5278,N_1020,N_2543);
nor U5279 (N_5279,N_2372,N_1844);
nand U5280 (N_5280,N_509,N_2575);
xnor U5281 (N_5281,N_4681,N_3740);
or U5282 (N_5282,N_4341,N_49);
nand U5283 (N_5283,N_3691,N_906);
xor U5284 (N_5284,N_4129,N_1188);
nand U5285 (N_5285,N_1302,N_4668);
xor U5286 (N_5286,N_338,N_1538);
and U5287 (N_5287,N_2744,N_4031);
or U5288 (N_5288,N_4337,N_3495);
nand U5289 (N_5289,N_223,N_171);
nor U5290 (N_5290,N_3462,N_2396);
and U5291 (N_5291,N_172,N_2431);
xnor U5292 (N_5292,N_803,N_2815);
and U5293 (N_5293,N_1813,N_3297);
nand U5294 (N_5294,N_2100,N_1027);
nor U5295 (N_5295,N_655,N_378);
or U5296 (N_5296,N_426,N_533);
nand U5297 (N_5297,N_1587,N_3784);
and U5298 (N_5298,N_3191,N_1040);
nand U5299 (N_5299,N_103,N_2150);
nand U5300 (N_5300,N_2456,N_3265);
nand U5301 (N_5301,N_4705,N_3780);
nor U5302 (N_5302,N_4188,N_2689);
and U5303 (N_5303,N_2500,N_995);
and U5304 (N_5304,N_2459,N_4543);
nor U5305 (N_5305,N_2555,N_3097);
nand U5306 (N_5306,N_733,N_744);
nor U5307 (N_5307,N_3239,N_2520);
nor U5308 (N_5308,N_1426,N_6);
nand U5309 (N_5309,N_516,N_4318);
nand U5310 (N_5310,N_2703,N_1678);
or U5311 (N_5311,N_4144,N_2182);
nor U5312 (N_5312,N_4141,N_4434);
nor U5313 (N_5313,N_471,N_3368);
nand U5314 (N_5314,N_4783,N_4580);
xnor U5315 (N_5315,N_2630,N_4961);
or U5316 (N_5316,N_3903,N_883);
nor U5317 (N_5317,N_3153,N_3376);
nor U5318 (N_5318,N_2414,N_4104);
nand U5319 (N_5319,N_4355,N_412);
and U5320 (N_5320,N_381,N_2962);
nand U5321 (N_5321,N_4174,N_4903);
nand U5322 (N_5322,N_2695,N_4134);
nand U5323 (N_5323,N_14,N_923);
nand U5324 (N_5324,N_4577,N_3183);
and U5325 (N_5325,N_3342,N_3629);
nor U5326 (N_5326,N_2878,N_3807);
or U5327 (N_5327,N_3641,N_858);
and U5328 (N_5328,N_2338,N_4530);
xor U5329 (N_5329,N_4718,N_484);
nand U5330 (N_5330,N_2705,N_4990);
or U5331 (N_5331,N_3768,N_3006);
nor U5332 (N_5332,N_4944,N_394);
nor U5333 (N_5333,N_4863,N_950);
nor U5334 (N_5334,N_1070,N_4068);
and U5335 (N_5335,N_4800,N_1348);
nor U5336 (N_5336,N_2419,N_4972);
nor U5337 (N_5337,N_2989,N_447);
and U5338 (N_5338,N_2099,N_871);
and U5339 (N_5339,N_4557,N_4574);
nand U5340 (N_5340,N_3430,N_996);
xor U5341 (N_5341,N_3036,N_4417);
or U5342 (N_5342,N_4613,N_946);
nand U5343 (N_5343,N_3009,N_4332);
nor U5344 (N_5344,N_29,N_2249);
nand U5345 (N_5345,N_4778,N_1054);
nor U5346 (N_5346,N_122,N_1949);
or U5347 (N_5347,N_4623,N_1248);
and U5348 (N_5348,N_662,N_978);
nand U5349 (N_5349,N_3333,N_4137);
xnor U5350 (N_5350,N_4387,N_214);
nor U5351 (N_5351,N_2888,N_608);
nand U5352 (N_5352,N_1529,N_4462);
nand U5353 (N_5353,N_3912,N_1624);
nand U5354 (N_5354,N_842,N_1751);
or U5355 (N_5355,N_3046,N_904);
nand U5356 (N_5356,N_1385,N_4121);
nand U5357 (N_5357,N_2200,N_646);
nor U5358 (N_5358,N_3323,N_4411);
and U5359 (N_5359,N_2810,N_3200);
and U5360 (N_5360,N_2739,N_1761);
and U5361 (N_5361,N_567,N_2822);
nand U5362 (N_5362,N_4986,N_4150);
or U5363 (N_5363,N_1832,N_4079);
nor U5364 (N_5364,N_4561,N_2691);
or U5365 (N_5365,N_3969,N_4371);
or U5366 (N_5366,N_1631,N_3091);
nand U5367 (N_5367,N_2574,N_3053);
nor U5368 (N_5368,N_1645,N_3070);
and U5369 (N_5369,N_3224,N_1760);
nor U5370 (N_5370,N_1494,N_151);
nor U5371 (N_5371,N_71,N_3653);
and U5372 (N_5372,N_1743,N_1341);
or U5373 (N_5373,N_2433,N_4397);
nand U5374 (N_5374,N_4532,N_2146);
nor U5375 (N_5375,N_835,N_4248);
nor U5376 (N_5376,N_2262,N_106);
or U5377 (N_5377,N_2205,N_1245);
or U5378 (N_5378,N_227,N_2511);
and U5379 (N_5379,N_3916,N_3540);
nor U5380 (N_5380,N_4879,N_2743);
and U5381 (N_5381,N_4080,N_207);
or U5382 (N_5382,N_1815,N_455);
and U5383 (N_5383,N_2343,N_660);
and U5384 (N_5384,N_3614,N_4660);
or U5385 (N_5385,N_4856,N_1796);
nand U5386 (N_5386,N_3978,N_4740);
or U5387 (N_5387,N_3004,N_4702);
and U5388 (N_5388,N_1317,N_2408);
or U5389 (N_5389,N_2060,N_442);
and U5390 (N_5390,N_671,N_4951);
nor U5391 (N_5391,N_4883,N_4227);
or U5392 (N_5392,N_1745,N_1487);
nand U5393 (N_5393,N_1853,N_2881);
and U5394 (N_5394,N_41,N_1820);
nor U5395 (N_5395,N_1614,N_1996);
nor U5396 (N_5396,N_222,N_3894);
nand U5397 (N_5397,N_468,N_2830);
nand U5398 (N_5398,N_285,N_406);
nor U5399 (N_5399,N_3748,N_2407);
nand U5400 (N_5400,N_3093,N_3424);
or U5401 (N_5401,N_3151,N_1827);
nor U5402 (N_5402,N_54,N_4028);
or U5403 (N_5403,N_4207,N_3057);
nor U5404 (N_5404,N_2257,N_593);
and U5405 (N_5405,N_1915,N_1118);
nand U5406 (N_5406,N_2891,N_658);
xor U5407 (N_5407,N_1166,N_1321);
xor U5408 (N_5408,N_421,N_2514);
or U5409 (N_5409,N_1602,N_4253);
and U5410 (N_5410,N_770,N_2254);
and U5411 (N_5411,N_903,N_1490);
xnor U5412 (N_5412,N_3829,N_4496);
and U5413 (N_5413,N_2473,N_2863);
and U5414 (N_5414,N_791,N_1013);
xnor U5415 (N_5415,N_321,N_3956);
or U5416 (N_5416,N_1149,N_1507);
and U5417 (N_5417,N_2608,N_1209);
nor U5418 (N_5418,N_2975,N_1406);
nand U5419 (N_5419,N_1970,N_3194);
or U5420 (N_5420,N_2532,N_3026);
or U5421 (N_5421,N_4302,N_4374);
nor U5422 (N_5422,N_2893,N_1778);
nor U5423 (N_5423,N_1055,N_2636);
and U5424 (N_5424,N_2518,N_3821);
or U5425 (N_5425,N_3643,N_1016);
nor U5426 (N_5426,N_3312,N_2236);
or U5427 (N_5427,N_2963,N_2234);
xnor U5428 (N_5428,N_4110,N_1331);
nand U5429 (N_5429,N_1228,N_4984);
nor U5430 (N_5430,N_4695,N_1986);
and U5431 (N_5431,N_4324,N_1767);
nor U5432 (N_5432,N_4402,N_97);
xor U5433 (N_5433,N_2722,N_1097);
nor U5434 (N_5434,N_4890,N_2698);
xnor U5435 (N_5435,N_3732,N_1953);
nand U5436 (N_5436,N_4524,N_358);
nor U5437 (N_5437,N_2074,N_316);
nor U5438 (N_5438,N_2838,N_4624);
nand U5439 (N_5439,N_1294,N_1359);
nand U5440 (N_5440,N_2499,N_1452);
nor U5441 (N_5441,N_3959,N_459);
or U5442 (N_5442,N_1464,N_687);
and U5443 (N_5443,N_960,N_977);
nand U5444 (N_5444,N_742,N_1912);
or U5445 (N_5445,N_2727,N_4818);
or U5446 (N_5446,N_1503,N_629);
nand U5447 (N_5447,N_573,N_1213);
xnor U5448 (N_5448,N_399,N_2241);
or U5449 (N_5449,N_2044,N_1581);
and U5450 (N_5450,N_4653,N_875);
and U5451 (N_5451,N_2468,N_3606);
and U5452 (N_5452,N_1176,N_1590);
nor U5453 (N_5453,N_3002,N_4772);
or U5454 (N_5454,N_1345,N_283);
nand U5455 (N_5455,N_1417,N_1873);
or U5456 (N_5456,N_175,N_3742);
and U5457 (N_5457,N_3981,N_4865);
or U5458 (N_5458,N_688,N_4657);
and U5459 (N_5459,N_3569,N_3129);
or U5460 (N_5460,N_1400,N_728);
and U5461 (N_5461,N_2105,N_1394);
nor U5462 (N_5462,N_765,N_1342);
xor U5463 (N_5463,N_3163,N_2983);
or U5464 (N_5464,N_99,N_2786);
and U5465 (N_5465,N_236,N_4857);
and U5466 (N_5466,N_1914,N_1940);
xnor U5467 (N_5467,N_581,N_1903);
and U5468 (N_5468,N_3697,N_4788);
nand U5469 (N_5469,N_2004,N_2535);
or U5470 (N_5470,N_1679,N_1655);
nand U5471 (N_5471,N_716,N_1123);
nand U5472 (N_5472,N_3634,N_2713);
nand U5473 (N_5473,N_1115,N_4436);
xor U5474 (N_5474,N_1584,N_2358);
and U5475 (N_5475,N_1547,N_4293);
xor U5476 (N_5476,N_2858,N_1946);
or U5477 (N_5477,N_1162,N_96);
nand U5478 (N_5478,N_1112,N_2998);
xnor U5479 (N_5479,N_1684,N_1886);
or U5480 (N_5480,N_1043,N_3920);
nor U5481 (N_5481,N_2319,N_93);
or U5482 (N_5482,N_2618,N_4190);
nor U5483 (N_5483,N_4255,N_4935);
nand U5484 (N_5484,N_3901,N_4655);
nor U5485 (N_5485,N_4157,N_1328);
or U5486 (N_5486,N_2832,N_2190);
and U5487 (N_5487,N_4161,N_4929);
or U5488 (N_5488,N_4922,N_1171);
nand U5489 (N_5489,N_1696,N_2103);
nor U5490 (N_5490,N_1208,N_2026);
nand U5491 (N_5491,N_2658,N_2803);
and U5492 (N_5492,N_3130,N_3836);
and U5493 (N_5493,N_2651,N_2273);
or U5494 (N_5494,N_1764,N_4215);
nor U5495 (N_5495,N_2024,N_514);
nand U5496 (N_5496,N_4413,N_3062);
nor U5497 (N_5497,N_4554,N_397);
or U5498 (N_5498,N_3892,N_583);
and U5499 (N_5499,N_1323,N_2095);
xor U5500 (N_5500,N_1781,N_156);
nand U5501 (N_5501,N_4100,N_1768);
nor U5502 (N_5502,N_1113,N_2509);
nand U5503 (N_5503,N_4981,N_4136);
or U5504 (N_5504,N_768,N_928);
or U5505 (N_5505,N_4349,N_3964);
or U5506 (N_5506,N_589,N_1623);
nand U5507 (N_5507,N_297,N_4766);
and U5508 (N_5508,N_178,N_256);
and U5509 (N_5509,N_1238,N_2308);
xnor U5510 (N_5510,N_2187,N_938);
or U5511 (N_5511,N_2462,N_3336);
and U5512 (N_5512,N_1715,N_3446);
nand U5513 (N_5513,N_2418,N_2859);
or U5514 (N_5514,N_3493,N_1958);
or U5515 (N_5515,N_4089,N_3050);
nand U5516 (N_5516,N_4898,N_4811);
or U5517 (N_5517,N_3468,N_3702);
nand U5518 (N_5518,N_1261,N_1984);
nor U5519 (N_5519,N_3767,N_1157);
nand U5520 (N_5520,N_2367,N_4825);
or U5521 (N_5521,N_116,N_2127);
xor U5522 (N_5522,N_125,N_2096);
nor U5523 (N_5523,N_873,N_882);
and U5524 (N_5524,N_4888,N_1089);
and U5525 (N_5525,N_102,N_2495);
or U5526 (N_5526,N_2147,N_4192);
or U5527 (N_5527,N_129,N_880);
and U5528 (N_5528,N_4427,N_3535);
or U5529 (N_5529,N_2613,N_2799);
nor U5530 (N_5530,N_4751,N_254);
or U5531 (N_5531,N_4870,N_2279);
nor U5532 (N_5532,N_4454,N_1068);
and U5533 (N_5533,N_2895,N_3879);
and U5534 (N_5534,N_336,N_1226);
nor U5535 (N_5535,N_1433,N_1787);
nand U5536 (N_5536,N_4534,N_4457);
or U5537 (N_5537,N_764,N_3551);
nor U5538 (N_5538,N_2755,N_901);
and U5539 (N_5539,N_4982,N_3143);
and U5540 (N_5540,N_3423,N_1526);
nand U5541 (N_5541,N_3806,N_1461);
xor U5542 (N_5542,N_4757,N_3437);
and U5543 (N_5543,N_1755,N_2278);
nand U5544 (N_5544,N_2339,N_4388);
nor U5545 (N_5545,N_2993,N_1925);
nand U5546 (N_5546,N_2916,N_107);
nand U5547 (N_5547,N_465,N_3700);
or U5548 (N_5548,N_137,N_820);
xor U5549 (N_5549,N_551,N_4829);
nand U5550 (N_5550,N_1742,N_1324);
and U5551 (N_5551,N_198,N_4334);
nand U5552 (N_5552,N_2175,N_242);
and U5553 (N_5553,N_2335,N_1731);
or U5554 (N_5554,N_1164,N_4633);
xor U5555 (N_5555,N_4590,N_3562);
and U5556 (N_5556,N_2978,N_2046);
or U5557 (N_5557,N_4686,N_1389);
nor U5558 (N_5558,N_4563,N_3435);
nor U5559 (N_5559,N_3197,N_511);
nor U5560 (N_5560,N_1716,N_2969);
xnor U5561 (N_5561,N_799,N_4047);
and U5562 (N_5562,N_4679,N_1600);
nor U5563 (N_5563,N_4481,N_4312);
nand U5564 (N_5564,N_1869,N_1181);
xor U5565 (N_5565,N_1897,N_1648);
or U5566 (N_5566,N_1548,N_1610);
or U5567 (N_5567,N_4866,N_4514);
and U5568 (N_5568,N_2391,N_4221);
or U5569 (N_5569,N_2112,N_2550);
or U5570 (N_5570,N_801,N_1777);
nor U5571 (N_5571,N_3358,N_460);
xor U5572 (N_5572,N_1029,N_1465);
nor U5573 (N_5573,N_2541,N_4350);
nand U5574 (N_5574,N_276,N_948);
and U5575 (N_5575,N_4339,N_502);
and U5576 (N_5576,N_4905,N_1775);
and U5577 (N_5577,N_932,N_1922);
nand U5578 (N_5578,N_1863,N_4250);
xor U5579 (N_5579,N_3883,N_1364);
or U5580 (N_5580,N_651,N_1630);
and U5581 (N_5581,N_4572,N_1725);
and U5582 (N_5582,N_839,N_2483);
nor U5583 (N_5583,N_3941,N_330);
nand U5584 (N_5584,N_2845,N_1735);
and U5585 (N_5585,N_2157,N_3525);
nor U5586 (N_5586,N_3819,N_2802);
or U5587 (N_5587,N_4037,N_3207);
nand U5588 (N_5588,N_3609,N_985);
nor U5589 (N_5589,N_2807,N_4072);
and U5590 (N_5590,N_2051,N_88);
nand U5591 (N_5591,N_2497,N_2005);
xor U5592 (N_5592,N_2688,N_4014);
xnor U5593 (N_5593,N_746,N_3830);
nor U5594 (N_5594,N_4478,N_1022);
nand U5595 (N_5595,N_834,N_3337);
nor U5596 (N_5596,N_2558,N_317);
nor U5597 (N_5597,N_3264,N_4882);
nor U5598 (N_5598,N_771,N_143);
nor U5599 (N_5599,N_2111,N_3258);
or U5600 (N_5600,N_3958,N_467);
or U5601 (N_5601,N_4112,N_1824);
or U5602 (N_5602,N_353,N_2318);
nor U5603 (N_5603,N_4435,N_3035);
nand U5604 (N_5604,N_4586,N_587);
nand U5605 (N_5605,N_333,N_2030);
xnor U5606 (N_5606,N_856,N_2284);
or U5607 (N_5607,N_1565,N_2672);
nor U5608 (N_5608,N_159,N_2745);
or U5609 (N_5609,N_1031,N_1524);
and U5610 (N_5610,N_3213,N_1197);
nor U5611 (N_5611,N_3914,N_193);
or U5612 (N_5612,N_1689,N_2489);
nor U5613 (N_5613,N_695,N_3165);
nor U5614 (N_5614,N_2549,N_1991);
nor U5615 (N_5615,N_1858,N_4077);
nor U5616 (N_5616,N_482,N_623);
or U5617 (N_5617,N_2602,N_4235);
xor U5618 (N_5618,N_3340,N_3067);
nand U5619 (N_5619,N_1661,N_1508);
nor U5620 (N_5620,N_4564,N_1804);
nand U5621 (N_5621,N_1478,N_1921);
or U5622 (N_5622,N_935,N_4186);
xor U5623 (N_5623,N_2475,N_1235);
xor U5624 (N_5624,N_16,N_909);
and U5625 (N_5625,N_4717,N_418);
and U5626 (N_5626,N_833,N_4353);
or U5627 (N_5627,N_3550,N_2457);
or U5628 (N_5628,N_3309,N_631);
and U5629 (N_5629,N_1376,N_4310);
nand U5630 (N_5630,N_4117,N_3828);
nand U5631 (N_5631,N_4980,N_2451);
or U5632 (N_5632,N_2933,N_4877);
nor U5633 (N_5633,N_3330,N_4670);
and U5634 (N_5634,N_3508,N_4519);
or U5635 (N_5635,N_1241,N_3081);
nand U5636 (N_5636,N_609,N_3987);
or U5637 (N_5637,N_1726,N_3079);
nor U5638 (N_5638,N_4729,N_3971);
or U5639 (N_5639,N_2524,N_1005);
xnor U5640 (N_5640,N_3314,N_987);
or U5641 (N_5641,N_1085,N_1288);
and U5642 (N_5642,N_3709,N_3824);
and U5643 (N_5643,N_570,N_879);
nand U5644 (N_5644,N_3974,N_2272);
nand U5645 (N_5645,N_3318,N_1582);
or U5646 (N_5646,N_2181,N_3710);
nor U5647 (N_5647,N_1215,N_3405);
xnor U5648 (N_5648,N_4966,N_4295);
or U5649 (N_5649,N_2329,N_3687);
nand U5650 (N_5650,N_3113,N_2392);
xnor U5651 (N_5651,N_794,N_1652);
and U5652 (N_5652,N_4438,N_2776);
and U5653 (N_5653,N_264,N_644);
and U5654 (N_5654,N_1957,N_4222);
and U5655 (N_5655,N_4787,N_2665);
or U5656 (N_5656,N_2061,N_1806);
xor U5657 (N_5657,N_206,N_4322);
nor U5658 (N_5658,N_1882,N_118);
nand U5659 (N_5659,N_3587,N_1560);
and U5660 (N_5660,N_1240,N_2460);
nand U5661 (N_5661,N_4064,N_3394);
nand U5662 (N_5662,N_3638,N_3505);
xnor U5663 (N_5663,N_1561,N_3195);
nor U5664 (N_5664,N_391,N_3474);
xnor U5665 (N_5665,N_2296,N_638);
and U5666 (N_5666,N_320,N_2440);
nor U5667 (N_5667,N_3012,N_1462);
nor U5668 (N_5668,N_1913,N_259);
nand U5669 (N_5669,N_4604,N_1773);
nand U5670 (N_5670,N_62,N_4834);
nor U5671 (N_5671,N_2333,N_2351);
xnor U5672 (N_5672,N_3727,N_27);
and U5673 (N_5673,N_1431,N_615);
or U5674 (N_5674,N_3532,N_3433);
xor U5675 (N_5675,N_1673,N_187);
nor U5676 (N_5676,N_245,N_2529);
nor U5677 (N_5677,N_4619,N_4793);
or U5678 (N_5678,N_942,N_1314);
nand U5679 (N_5679,N_3760,N_3296);
xnor U5680 (N_5680,N_1145,N_3870);
or U5681 (N_5681,N_2640,N_1938);
nor U5682 (N_5682,N_216,N_1320);
nand U5683 (N_5683,N_4340,N_250);
xnor U5684 (N_5684,N_36,N_4209);
xnor U5685 (N_5685,N_4964,N_1765);
nand U5686 (N_5686,N_209,N_3098);
xnor U5687 (N_5687,N_2270,N_3549);
and U5688 (N_5688,N_797,N_2153);
and U5689 (N_5689,N_2972,N_2932);
nor U5690 (N_5690,N_4176,N_3610);
nand U5691 (N_5691,N_4468,N_2821);
or U5692 (N_5692,N_810,N_1435);
nand U5693 (N_5693,N_4822,N_2870);
nand U5694 (N_5694,N_4075,N_2864);
and U5695 (N_5695,N_1790,N_3219);
nor U5696 (N_5696,N_3988,N_1419);
nor U5697 (N_5697,N_1399,N_1920);
nand U5698 (N_5698,N_2874,N_1295);
or U5699 (N_5699,N_1147,N_2450);
nor U5700 (N_5700,N_2844,N_3287);
nor U5701 (N_5701,N_2808,N_4429);
nand U5702 (N_5702,N_337,N_3250);
and U5703 (N_5703,N_1429,N_3302);
nand U5704 (N_5704,N_4162,N_416);
or U5705 (N_5705,N_4257,N_3858);
and U5706 (N_5706,N_373,N_1607);
nor U5707 (N_5707,N_2346,N_2169);
xnor U5708 (N_5708,N_4821,N_3352);
nor U5709 (N_5709,N_881,N_558);
nor U5710 (N_5710,N_2399,N_4730);
xnor U5711 (N_5711,N_2759,N_4659);
nand U5712 (N_5712,N_2742,N_2753);
xor U5713 (N_5713,N_3381,N_2444);
nand U5714 (N_5714,N_1692,N_113);
nor U5715 (N_5715,N_3715,N_572);
nand U5716 (N_5716,N_3232,N_3387);
nand U5717 (N_5717,N_1423,N_4861);
nor U5718 (N_5718,N_1609,N_2397);
nor U5719 (N_5719,N_1336,N_3479);
or U5720 (N_5720,N_2068,N_4460);
or U5721 (N_5721,N_3872,N_410);
nor U5722 (N_5722,N_4798,N_2656);
nor U5723 (N_5723,N_3229,N_2820);
or U5724 (N_5724,N_2943,N_311);
and U5725 (N_5725,N_4754,N_2465);
xor U5726 (N_5726,N_4319,N_4953);
nand U5727 (N_5727,N_2081,N_76);
nor U5728 (N_5728,N_2345,N_1759);
or U5729 (N_5729,N_3478,N_1088);
or U5730 (N_5730,N_2259,N_653);
nor U5731 (N_5731,N_366,N_4497);
nand U5732 (N_5732,N_2944,N_650);
or U5733 (N_5733,N_3619,N_3220);
and U5734 (N_5734,N_4860,N_568);
and U5735 (N_5735,N_3416,N_4501);
or U5736 (N_5736,N_3327,N_3236);
nor U5737 (N_5737,N_3491,N_4424);
nand U5738 (N_5738,N_1243,N_1936);
nor U5739 (N_5739,N_1072,N_3172);
and U5740 (N_5740,N_3267,N_4407);
and U5741 (N_5741,N_679,N_1065);
and U5742 (N_5742,N_4370,N_3556);
and U5743 (N_5743,N_3976,N_1700);
nand U5744 (N_5744,N_2721,N_2305);
and U5745 (N_5745,N_544,N_1214);
nand U5746 (N_5746,N_1875,N_1449);
nor U5747 (N_5747,N_1492,N_696);
or U5748 (N_5748,N_1651,N_1063);
and U5749 (N_5749,N_4268,N_1880);
nand U5750 (N_5750,N_3089,N_2280);
nand U5751 (N_5751,N_329,N_497);
nand U5752 (N_5752,N_127,N_1207);
or U5753 (N_5753,N_1470,N_4938);
xnor U5754 (N_5754,N_2109,N_4841);
nor U5755 (N_5755,N_3719,N_3750);
or U5756 (N_5756,N_4626,N_314);
and U5757 (N_5757,N_2377,N_541);
nor U5758 (N_5758,N_4540,N_1838);
or U5759 (N_5759,N_3317,N_1316);
and U5760 (N_5760,N_4685,N_1216);
and U5761 (N_5761,N_4201,N_2619);
or U5762 (N_5762,N_84,N_3270);
nor U5763 (N_5763,N_451,N_3228);
nor U5764 (N_5764,N_1871,N_4256);
nand U5765 (N_5765,N_2108,N_3140);
nor U5766 (N_5766,N_1038,N_1812);
nor U5767 (N_5767,N_4063,N_4008);
nor U5768 (N_5768,N_2300,N_2498);
and U5769 (N_5769,N_4589,N_2684);
nand U5770 (N_5770,N_3362,N_3279);
nor U5771 (N_5771,N_2472,N_1380);
or U5772 (N_5772,N_4199,N_3938);
and U5773 (N_5773,N_4070,N_3503);
nand U5774 (N_5774,N_4646,N_4722);
nor U5775 (N_5775,N_40,N_3801);
or U5776 (N_5776,N_111,N_277);
or U5777 (N_5777,N_3242,N_2594);
xnor U5778 (N_5778,N_4151,N_1642);
xnor U5779 (N_5779,N_1597,N_1829);
and U5780 (N_5780,N_4208,N_1304);
and U5781 (N_5781,N_4296,N_4552);
nand U5782 (N_5782,N_4541,N_2827);
nand U5783 (N_5783,N_3253,N_3677);
nand U5784 (N_5784,N_1473,N_2413);
nor U5785 (N_5785,N_3355,N_4726);
or U5786 (N_5786,N_380,N_740);
xnor U5787 (N_5787,N_2453,N_1591);
xnor U5788 (N_5788,N_4600,N_1083);
or U5789 (N_5789,N_4393,N_3917);
nor U5790 (N_5790,N_1409,N_3180);
nand U5791 (N_5791,N_2540,N_4763);
nand U5792 (N_5792,N_4512,N_1732);
and U5793 (N_5793,N_4363,N_1486);
nand U5794 (N_5794,N_1111,N_602);
nor U5795 (N_5795,N_3255,N_1512);
xor U5796 (N_5796,N_1900,N_2894);
and U5797 (N_5797,N_706,N_1439);
or U5798 (N_5798,N_411,N_4430);
nor U5799 (N_5799,N_257,N_168);
nand U5800 (N_5800,N_4637,N_566);
nand U5801 (N_5801,N_2545,N_3989);
or U5802 (N_5802,N_1260,N_2747);
xor U5803 (N_5803,N_3531,N_4323);
and U5804 (N_5804,N_2471,N_4027);
nand U5805 (N_5805,N_2578,N_2117);
and U5806 (N_5806,N_2866,N_876);
nor U5807 (N_5807,N_4308,N_2295);
or U5808 (N_5808,N_4352,N_4937);
or U5809 (N_5809,N_2913,N_312);
or U5810 (N_5810,N_3121,N_1567);
nand U5811 (N_5811,N_3979,N_2922);
or U5812 (N_5812,N_428,N_409);
xnor U5813 (N_5813,N_2562,N_2726);
xnor U5814 (N_5814,N_140,N_490);
or U5815 (N_5815,N_3919,N_2737);
nor U5816 (N_5816,N_4040,N_3567);
nor U5817 (N_5817,N_4309,N_3243);
nand U5818 (N_5818,N_3999,N_1710);
or U5819 (N_5819,N_4260,N_3543);
nor U5820 (N_5820,N_2675,N_1373);
nor U5821 (N_5821,N_3365,N_2025);
and U5822 (N_5822,N_3846,N_4525);
or U5823 (N_5823,N_4683,N_937);
nand U5824 (N_5824,N_1222,N_2788);
nor U5825 (N_5825,N_3008,N_1939);
and U5826 (N_5826,N_4098,N_4983);
or U5827 (N_5827,N_4776,N_2842);
nor U5828 (N_5828,N_2964,N_1135);
nand U5829 (N_5829,N_1466,N_4958);
or U5830 (N_5830,N_4043,N_1864);
nand U5831 (N_5831,N_2770,N_4824);
nor U5832 (N_5832,N_2567,N_1682);
and U5833 (N_5833,N_281,N_773);
or U5834 (N_5834,N_3524,N_3117);
or U5835 (N_5835,N_2652,N_80);
or U5836 (N_5836,N_2800,N_940);
nor U5837 (N_5837,N_1646,N_4252);
xnor U5838 (N_5838,N_684,N_3484);
or U5839 (N_5839,N_2352,N_1231);
or U5840 (N_5840,N_4125,N_4106);
and U5841 (N_5841,N_4472,N_2765);
and U5842 (N_5842,N_4622,N_4288);
nand U5843 (N_5843,N_4392,N_4779);
nor U5844 (N_5844,N_4109,N_4381);
nor U5845 (N_5845,N_3166,N_4544);
or U5846 (N_5846,N_920,N_4896);
or U5847 (N_5847,N_4831,N_2162);
and U5848 (N_5848,N_990,N_915);
and U5849 (N_5849,N_905,N_1434);
nor U5850 (N_5850,N_1819,N_891);
nand U5851 (N_5851,N_4758,N_3114);
and U5852 (N_5852,N_4902,N_4616);
nand U5853 (N_5853,N_3972,N_3133);
xnor U5854 (N_5854,N_3452,N_2189);
nor U5855 (N_5855,N_1140,N_1129);
nand U5856 (N_5856,N_1444,N_3752);
or U5857 (N_5857,N_1931,N_4513);
nor U5858 (N_5858,N_4932,N_4752);
and U5859 (N_5859,N_2986,N_384);
nor U5860 (N_5860,N_2548,N_3623);
and U5861 (N_5861,N_4290,N_82);
and U5862 (N_5862,N_30,N_4939);
nor U5863 (N_5863,N_2163,N_407);
nand U5864 (N_5864,N_1885,N_2361);
nand U5865 (N_5865,N_792,N_3751);
nor U5866 (N_5866,N_1856,N_3363);
or U5867 (N_5867,N_1310,N_3640);
nor U5868 (N_5868,N_2967,N_1762);
or U5869 (N_5869,N_4819,N_1937);
or U5870 (N_5870,N_98,N_2668);
nor U5871 (N_5871,N_2380,N_4058);
or U5872 (N_5872,N_477,N_4569);
nand U5873 (N_5873,N_2323,N_980);
or U5874 (N_5874,N_3018,N_3595);
nand U5875 (N_5875,N_3108,N_1311);
nand U5876 (N_5876,N_2814,N_2570);
xnor U5877 (N_5877,N_3597,N_4635);
and U5878 (N_5878,N_3665,N_2627);
and U5879 (N_5879,N_1339,N_1480);
nor U5880 (N_5880,N_4691,N_1573);
and U5881 (N_5881,N_894,N_306);
nor U5882 (N_5882,N_2544,N_1189);
or U5883 (N_5883,N_1050,N_3285);
nand U5884 (N_5884,N_2415,N_3573);
or U5885 (N_5885,N_1484,N_1894);
nand U5886 (N_5886,N_1552,N_3838);
and U5887 (N_5887,N_2093,N_1287);
and U5888 (N_5888,N_3206,N_1906);
and U5889 (N_5889,N_1280,N_349);
or U5890 (N_5890,N_3347,N_1523);
and U5891 (N_5891,N_4712,N_2224);
nor U5892 (N_5892,N_4940,N_1143);
nor U5893 (N_5893,N_131,N_1279);
or U5894 (N_5894,N_2016,N_3523);
nor U5895 (N_5895,N_4596,N_4386);
nand U5896 (N_5896,N_273,N_667);
nand U5897 (N_5897,N_1095,N_4010);
nand U5898 (N_5898,N_13,N_1997);
or U5899 (N_5899,N_2794,N_1392);
and U5900 (N_5900,N_2644,N_4060);
nor U5901 (N_5901,N_1772,N_313);
nand U5902 (N_5902,N_3353,N_991);
or U5903 (N_5903,N_1330,N_2253);
nor U5904 (N_5904,N_2805,N_139);
nor U5905 (N_5905,N_4167,N_1542);
xor U5906 (N_5906,N_134,N_1862);
and U5907 (N_5907,N_2782,N_4020);
nand U5908 (N_5908,N_3944,N_2650);
and U5909 (N_5909,N_3966,N_462);
xnor U5910 (N_5910,N_4768,N_3179);
or U5911 (N_5911,N_2326,N_3585);
and U5912 (N_5912,N_1232,N_2819);
or U5913 (N_5913,N_3759,N_2884);
and U5914 (N_5914,N_4082,N_160);
xnor U5915 (N_5915,N_105,N_1599);
or U5916 (N_5916,N_61,N_3246);
xor U5917 (N_5917,N_100,N_3841);
nand U5918 (N_5918,N_3635,N_480);
nor U5919 (N_5919,N_1667,N_560);
nand U5920 (N_5920,N_46,N_3714);
or U5921 (N_5921,N_217,N_1923);
nor U5922 (N_5922,N_1141,N_1179);
nand U5923 (N_5923,N_2671,N_2945);
nor U5924 (N_5924,N_141,N_1687);
nand U5925 (N_5925,N_1369,N_293);
xor U5926 (N_5926,N_2677,N_2439);
nand U5927 (N_5927,N_3608,N_4605);
nor U5928 (N_5928,N_528,N_1117);
or U5929 (N_5929,N_584,N_4956);
nor U5930 (N_5930,N_1803,N_4645);
xnor U5931 (N_5931,N_3272,N_3839);
and U5932 (N_5932,N_1332,N_2950);
nor U5933 (N_5933,N_2787,N_4007);
and U5934 (N_5934,N_4587,N_3326);
nor U5935 (N_5935,N_2321,N_3563);
or U5936 (N_5936,N_3069,N_3582);
nor U5937 (N_5937,N_1896,N_4529);
or U5938 (N_5938,N_798,N_2791);
nand U5939 (N_5939,N_2194,N_19);
nand U5940 (N_5940,N_3188,N_2926);
nand U5941 (N_5941,N_1293,N_808);
nor U5942 (N_5942,N_2851,N_2889);
or U5943 (N_5943,N_488,N_3571);
nand U5944 (N_5944,N_4943,N_4704);
or U5945 (N_5945,N_931,N_3721);
nand U5946 (N_5946,N_3792,N_3787);
or U5947 (N_5947,N_2480,N_788);
nor U5948 (N_5948,N_3910,N_382);
nand U5949 (N_5949,N_2948,N_761);
xnor U5950 (N_5950,N_1062,N_2823);
and U5951 (N_5951,N_1424,N_1242);
nand U5952 (N_5952,N_2924,N_4336);
nand U5953 (N_5953,N_3581,N_165);
nand U5954 (N_5954,N_3156,N_1791);
nand U5955 (N_5955,N_4850,N_248);
or U5956 (N_5956,N_2166,N_4313);
or U5957 (N_5957,N_2306,N_1770);
nand U5958 (N_5958,N_3173,N_793);
nand U5959 (N_5959,N_2781,N_4455);
nor U5960 (N_5960,N_3725,N_292);
and U5961 (N_5961,N_3382,N_4515);
nor U5962 (N_5962,N_965,N_4843);
or U5963 (N_5963,N_4967,N_1504);
and U5964 (N_5964,N_4612,N_763);
xnor U5965 (N_5965,N_2736,N_2387);
nand U5966 (N_5966,N_3847,N_1497);
and U5967 (N_5967,N_3817,N_395);
and U5968 (N_5968,N_3320,N_2872);
nand U5969 (N_5969,N_2761,N_2085);
nand U5970 (N_5970,N_3170,N_3218);
or U5971 (N_5971,N_535,N_190);
and U5972 (N_5972,N_4755,N_2667);
xor U5973 (N_5973,N_1596,N_2310);
or U5974 (N_5974,N_561,N_800);
nand U5975 (N_5975,N_3448,N_1148);
nand U5976 (N_5976,N_3805,N_690);
nand U5977 (N_5977,N_3322,N_4917);
or U5978 (N_5978,N_3284,N_3699);
nor U5979 (N_5979,N_1275,N_1076);
nand U5980 (N_5980,N_1955,N_4437);
or U5981 (N_5981,N_4244,N_2075);
or U5982 (N_5982,N_823,N_4606);
and U5983 (N_5983,N_4195,N_4976);
or U5984 (N_5984,N_3730,N_665);
nor U5985 (N_5985,N_2873,N_331);
nand U5986 (N_5986,N_356,N_3705);
and U5987 (N_5987,N_302,N_3548);
nor U5988 (N_5988,N_4401,N_4632);
nand U5989 (N_5989,N_3731,N_3871);
or U5990 (N_5990,N_1606,N_929);
or U5991 (N_5991,N_1911,N_2771);
nor U5992 (N_5992,N_443,N_4828);
nor U5993 (N_5993,N_2693,N_2027);
or U5994 (N_5994,N_1021,N_2647);
nand U5995 (N_5995,N_2427,N_3073);
or U5996 (N_5996,N_3686,N_4573);
or U5997 (N_5997,N_575,N_4996);
nor U5998 (N_5998,N_2229,N_1299);
or U5999 (N_5999,N_3456,N_3074);
nor U6000 (N_6000,N_811,N_1825);
and U6001 (N_6001,N_2638,N_63);
or U6002 (N_6002,N_4274,N_1995);
or U6003 (N_6003,N_4878,N_3579);
or U6004 (N_6004,N_4484,N_1265);
and U6005 (N_6005,N_4425,N_4231);
nand U6006 (N_6006,N_2871,N_4959);
nor U6007 (N_6007,N_755,N_202);
nand U6008 (N_6008,N_617,N_1717);
nor U6009 (N_6009,N_981,N_4708);
nand U6010 (N_6010,N_3794,N_2988);
nor U6011 (N_6011,N_4204,N_4278);
nor U6012 (N_6012,N_1002,N_727);
nor U6013 (N_6013,N_4267,N_4187);
and U6014 (N_6014,N_448,N_91);
and U6015 (N_6015,N_224,N_3056);
or U6016 (N_6016,N_3119,N_1259);
nor U6017 (N_6017,N_1626,N_57);
xor U6018 (N_6018,N_2757,N_3385);
nand U6019 (N_6019,N_3889,N_908);
or U6020 (N_6020,N_1313,N_386);
nor U6021 (N_6021,N_4461,N_3160);
nor U6022 (N_6022,N_3458,N_1253);
and U6023 (N_6023,N_4648,N_360);
nand U6024 (N_6024,N_1137,N_1551);
nand U6025 (N_6025,N_3252,N_3704);
nand U6026 (N_6026,N_3380,N_3465);
and U6027 (N_6027,N_3935,N_3496);
or U6028 (N_6028,N_2701,N_4423);
or U6029 (N_6029,N_1881,N_1127);
nor U6030 (N_6030,N_4016,N_1210);
nand U6031 (N_6031,N_708,N_2836);
nand U6032 (N_6032,N_2131,N_1660);
nand U6033 (N_6033,N_2156,N_999);
and U6034 (N_6034,N_821,N_3417);
nor U6035 (N_6035,N_4949,N_1680);
nand U6036 (N_6036,N_1109,N_1467);
or U6037 (N_6037,N_2861,N_4999);
nor U6038 (N_6038,N_1183,N_3015);
nor U6039 (N_6039,N_2707,N_3449);
nand U6040 (N_6040,N_4553,N_4431);
nand U6041 (N_6041,N_3231,N_2942);
xor U6042 (N_6042,N_621,N_1225);
or U6043 (N_6043,N_837,N_1325);
and U6044 (N_6044,N_2052,N_4226);
nand U6045 (N_6045,N_676,N_2379);
nor U6046 (N_6046,N_3663,N_3223);
and U6047 (N_6047,N_184,N_1167);
nor U6048 (N_6048,N_3782,N_3116);
and U6049 (N_6049,N_1393,N_1244);
or U6050 (N_6050,N_2617,N_4671);
or U6051 (N_6051,N_1082,N_1746);
or U6052 (N_6052,N_2428,N_3948);
and U6053 (N_6053,N_2857,N_1121);
and U6054 (N_6054,N_2900,N_3779);
nor U6055 (N_6055,N_2612,N_2579);
or U6056 (N_6056,N_2195,N_1278);
or U6057 (N_6057,N_2571,N_845);
and U6058 (N_6058,N_4725,N_4479);
nand U6059 (N_6059,N_984,N_2216);
and U6060 (N_6060,N_2968,N_3698);
or U6061 (N_6061,N_4418,N_1738);
or U6062 (N_6062,N_1110,N_3351);
nand U6063 (N_6063,N_1779,N_3346);
nand U6064 (N_6064,N_4168,N_3560);
nor U6065 (N_6065,N_483,N_2949);
and U6066 (N_6066,N_2033,N_2519);
or U6067 (N_6067,N_2717,N_515);
or U6068 (N_6068,N_3485,N_4409);
nor U6069 (N_6069,N_4526,N_3620);
xor U6070 (N_6070,N_2029,N_2775);
xnor U6071 (N_6071,N_778,N_4506);
or U6072 (N_6072,N_4111,N_3621);
and U6073 (N_6073,N_3386,N_3537);
and U6074 (N_6074,N_682,N_2148);
nor U6075 (N_6075,N_2432,N_3500);
nand U6076 (N_6076,N_4582,N_2809);
nor U6077 (N_6077,N_2606,N_1518);
or U6078 (N_6078,N_2293,N_4701);
nand U6079 (N_6079,N_1049,N_2078);
nand U6080 (N_6080,N_3564,N_3230);
and U6081 (N_6081,N_1985,N_4404);
nor U6082 (N_6082,N_2655,N_3626);
xnor U6083 (N_6083,N_310,N_4774);
and U6084 (N_6084,N_81,N_1425);
or U6085 (N_6085,N_3349,N_3921);
nor U6086 (N_6086,N_1568,N_2299);
xor U6087 (N_6087,N_645,N_654);
and U6088 (N_6088,N_377,N_1909);
nand U6089 (N_6089,N_870,N_749);
and U6090 (N_6090,N_3149,N_3426);
or U6091 (N_6091,N_975,N_208);
and U6092 (N_6092,N_2155,N_3343);
nand U6093 (N_6093,N_2072,N_3590);
xor U6094 (N_6094,N_3096,N_3087);
and U6095 (N_6095,N_153,N_3924);
nand U6096 (N_6096,N_2525,N_2569);
and U6097 (N_6097,N_3692,N_3301);
and U6098 (N_6098,N_3796,N_278);
nor U6099 (N_6099,N_2754,N_606);
or U6100 (N_6100,N_2825,N_3820);
nand U6101 (N_6101,N_4790,N_1904);
nor U6102 (N_6102,N_2090,N_1516);
nor U6103 (N_6103,N_1037,N_357);
nor U6104 (N_6104,N_4504,N_3632);
xnor U6105 (N_6105,N_3615,N_2828);
or U6106 (N_6106,N_4921,N_1223);
nand U6107 (N_6107,N_3591,N_1855);
or U6108 (N_6108,N_186,N_1879);
nand U6109 (N_6109,N_2546,N_4568);
or U6110 (N_6110,N_2360,N_4469);
xor U6111 (N_6111,N_1133,N_2381);
nand U6112 (N_6112,N_3882,N_3182);
or U6113 (N_6113,N_4827,N_1705);
and U6114 (N_6114,N_4345,N_1783);
and U6115 (N_6115,N_3915,N_503);
nor U6116 (N_6116,N_3530,N_4963);
and U6117 (N_6117,N_3954,N_4709);
nand U6118 (N_6118,N_219,N_2817);
and U6119 (N_6119,N_3904,N_588);
or U6120 (N_6120,N_4126,N_3481);
or U6121 (N_6121,N_2288,N_3881);
nand U6122 (N_6122,N_3772,N_531);
nand U6123 (N_6123,N_1572,N_3607);
nand U6124 (N_6124,N_199,N_693);
nor U6125 (N_6125,N_4678,N_3315);
or U6126 (N_6126,N_523,N_2265);
nor U6127 (N_6127,N_2811,N_3450);
or U6128 (N_6128,N_1502,N_334);
nor U6129 (N_6129,N_3464,N_2905);
or U6130 (N_6130,N_846,N_4785);
nor U6131 (N_6131,N_4283,N_618);
or U6132 (N_6132,N_4415,N_369);
xnor U6133 (N_6133,N_2632,N_579);
or U6134 (N_6134,N_1941,N_3262);
nor U6135 (N_6135,N_110,N_2604);
or U6136 (N_6136,N_3221,N_767);
nand U6137 (N_6137,N_4749,N_3029);
or U6138 (N_6138,N_3126,N_4128);
or U6139 (N_6139,N_4485,N_3357);
and U6140 (N_6140,N_888,N_3898);
nor U6141 (N_6141,N_872,N_2589);
xnor U6142 (N_6142,N_50,N_1491);
nand U6143 (N_6143,N_709,N_657);
or U6144 (N_6144,N_2896,N_4038);
and U6145 (N_6145,N_1367,N_4094);
or U6146 (N_6146,N_475,N_1436);
nand U6147 (N_6147,N_2186,N_3652);
nor U6148 (N_6148,N_4463,N_1665);
xor U6149 (N_6149,N_649,N_4663);
nor U6150 (N_6150,N_1657,N_1802);
nor U6151 (N_6151,N_1541,N_4647);
nor U6152 (N_6152,N_2729,N_3256);
and U6153 (N_6153,N_603,N_212);
or U6154 (N_6154,N_836,N_3980);
nor U6155 (N_6155,N_4049,N_4842);
or U6156 (N_6156,N_3208,N_355);
nand U6157 (N_6157,N_2769,N_3065);
nand U6158 (N_6158,N_1427,N_4546);
nor U6159 (N_6159,N_3659,N_4955);
nor U6160 (N_6160,N_2158,N_4078);
nor U6161 (N_6161,N_3321,N_741);
and U6162 (N_6162,N_704,N_0);
and U6163 (N_6163,N_3867,N_2374);
xnor U6164 (N_6164,N_8,N_3454);
nor U6165 (N_6165,N_3455,N_4808);
nor U6166 (N_6166,N_4975,N_668);
or U6167 (N_6167,N_1847,N_3472);
nor U6168 (N_6168,N_2043,N_1598);
nor U6169 (N_6169,N_1358,N_3925);
xor U6170 (N_6170,N_2869,N_1586);
nor U6171 (N_6171,N_2446,N_637);
and U6172 (N_6172,N_3370,N_4459);
nand U6173 (N_6173,N_1004,N_4780);
or U6174 (N_6174,N_352,N_2212);
or U6175 (N_6175,N_2720,N_2642);
nor U6176 (N_6176,N_3837,N_2464);
nor U6177 (N_6177,N_2066,N_492);
or U6178 (N_6178,N_3204,N_678);
xnor U6179 (N_6179,N_2057,N_325);
or U6180 (N_6180,N_4467,N_3289);
or U6181 (N_6181,N_3150,N_4035);
nor U6182 (N_6182,N_3251,N_1711);
or U6183 (N_6183,N_865,N_3690);
nor U6184 (N_6184,N_917,N_1411);
or U6185 (N_6185,N_1437,N_1613);
nand U6186 (N_6186,N_1835,N_4689);
or U6187 (N_6187,N_1366,N_2600);
or U6188 (N_6188,N_530,N_2185);
xnor U6189 (N_6189,N_2354,N_1060);
and U6190 (N_6190,N_4331,N_3940);
nor U6191 (N_6191,N_3457,N_2314);
or U6192 (N_6192,N_2171,N_4651);
or U6193 (N_6193,N_3000,N_3707);
xnor U6194 (N_6194,N_1784,N_3800);
or U6195 (N_6195,N_1451,N_1347);
nor U6196 (N_6196,N_4714,N_3685);
xnor U6197 (N_6197,N_3403,N_1962);
or U6198 (N_6198,N_1654,N_376);
nor U6199 (N_6199,N_1633,N_4895);
nor U6200 (N_6200,N_2512,N_149);
xnor U6201 (N_6201,N_3480,N_1747);
nand U6202 (N_6202,N_2740,N_3167);
or U6203 (N_6203,N_4487,N_4855);
and U6204 (N_6204,N_2059,N_639);
nand U6205 (N_6205,N_735,N_1154);
and U6206 (N_6206,N_2267,N_1334);
nand U6207 (N_6207,N_3711,N_1365);
or U6208 (N_6208,N_1816,N_1315);
nand U6209 (N_6209,N_1305,N_941);
and U6210 (N_6210,N_1165,N_4802);
xnor U6211 (N_6211,N_2738,N_15);
or U6212 (N_6212,N_4522,N_2247);
nand U6213 (N_6213,N_532,N_414);
or U6214 (N_6214,N_564,N_4033);
nor U6215 (N_6215,N_286,N_3803);
nand U6216 (N_6216,N_363,N_2142);
and U6217 (N_6217,N_796,N_3810);
nand U6218 (N_6218,N_726,N_4127);
or U6219 (N_6219,N_1786,N_3655);
nand U6220 (N_6220,N_3973,N_2002);
nand U6221 (N_6221,N_166,N_3773);
nand U6222 (N_6222,N_4453,N_2917);
or U6223 (N_6223,N_3557,N_2315);
and U6224 (N_6224,N_907,N_89);
or U6225 (N_6225,N_4232,N_1030);
and U6226 (N_6226,N_1410,N_1093);
or U6227 (N_6227,N_2564,N_2452);
or U6228 (N_6228,N_2233,N_878);
xor U6229 (N_6229,N_4942,N_4669);
and U6230 (N_6230,N_396,N_2286);
and U6231 (N_6231,N_1739,N_4021);
or U6232 (N_6232,N_1319,N_1601);
and U6233 (N_6233,N_2394,N_3955);
nor U6234 (N_6234,N_4464,N_4581);
nor U6235 (N_6235,N_3,N_3546);
nand U6236 (N_6236,N_4412,N_1530);
nor U6237 (N_6237,N_4159,N_1890);
nor U6238 (N_6238,N_2850,N_1535);
xnor U6239 (N_6239,N_3694,N_1010);
or U6240 (N_6240,N_4836,N_275);
nand U6241 (N_6241,N_37,N_1632);
nor U6242 (N_6242,N_956,N_371);
nand U6243 (N_6243,N_2356,N_1521);
nor U6244 (N_6244,N_270,N_1622);
and U6245 (N_6245,N_1954,N_4741);
or U6246 (N_6246,N_624,N_2384);
or U6247 (N_6247,N_2011,N_2330);
and U6248 (N_6248,N_375,N_966);
nand U6249 (N_6249,N_1025,N_2484);
nor U6250 (N_6250,N_213,N_2768);
and U6251 (N_6251,N_884,N_389);
xor U6252 (N_6252,N_4421,N_4971);
or U6253 (N_6253,N_1268,N_3645);
or U6254 (N_6254,N_961,N_1849);
xnor U6255 (N_6255,N_1447,N_4191);
or U6256 (N_6256,N_852,N_3055);
and U6257 (N_6257,N_1036,N_2401);
or U6258 (N_6258,N_3486,N_1370);
or U6259 (N_6259,N_963,N_1635);
and U6260 (N_6260,N_4936,N_4833);
xnor U6261 (N_6261,N_3555,N_3826);
nor U6262 (N_6262,N_4864,N_4711);
xor U6263 (N_6263,N_4852,N_2493);
nand U6264 (N_6264,N_1155,N_3729);
and U6265 (N_6265,N_1405,N_1282);
nand U6266 (N_6266,N_1908,N_4523);
nand U6267 (N_6267,N_164,N_4280);
and U6268 (N_6268,N_988,N_3628);
nand U6269 (N_6269,N_3234,N_4771);
nor U6270 (N_6270,N_549,N_4500);
nand U6271 (N_6271,N_3186,N_269);
xnor U6272 (N_6272,N_4001,N_22);
nor U6273 (N_6273,N_4155,N_807);
xor U6274 (N_6274,N_804,N_2110);
nor U6275 (N_6275,N_4303,N_3292);
and U6276 (N_6276,N_3764,N_900);
or U6277 (N_6277,N_3895,N_4991);
nor U6278 (N_6278,N_1126,N_3506);
and U6279 (N_6279,N_1905,N_2661);
and U6280 (N_6280,N_1788,N_2366);
nor U6281 (N_6281,N_4287,N_1150);
xor U6282 (N_6282,N_2463,N_2954);
nor U6283 (N_6283,N_1161,N_2340);
nand U6284 (N_6284,N_12,N_7);
and U6285 (N_6285,N_2778,N_1522);
nand U6286 (N_6286,N_4642,N_1736);
nand U6287 (N_6287,N_2429,N_3877);
or U6288 (N_6288,N_3722,N_2521);
xnor U6289 (N_6289,N_3011,N_2357);
and U6290 (N_6290,N_1580,N_109);
nor U6291 (N_6291,N_429,N_2076);
nor U6292 (N_6292,N_182,N_3962);
nor U6293 (N_6293,N_3196,N_736);
nand U6294 (N_6294,N_3515,N_756);
or U6295 (N_6295,N_4672,N_968);
or U6296 (N_6296,N_1309,N_4200);
and U6297 (N_6297,N_4452,N_1658);
xor U6298 (N_6298,N_1308,N_59);
and U6299 (N_6299,N_2344,N_1556);
and U6300 (N_6300,N_3215,N_4551);
xnor U6301 (N_6301,N_612,N_3570);
nor U6302 (N_6302,N_4284,N_2875);
or U6303 (N_6303,N_3137,N_4521);
and U6304 (N_6304,N_4753,N_4947);
nand U6305 (N_6305,N_4291,N_3075);
or U6306 (N_6306,N_3650,N_1052);
and U6307 (N_6307,N_1916,N_3101);
or U6308 (N_6308,N_271,N_3795);
nand U6309 (N_6309,N_4139,N_3128);
and U6310 (N_6310,N_3030,N_1296);
nand U6311 (N_6311,N_4542,N_3092);
xnor U6312 (N_6312,N_1420,N_1517);
or U6313 (N_6313,N_3519,N_2196);
or U6314 (N_6314,N_1675,N_4809);
nor U6315 (N_6315,N_747,N_2756);
nand U6316 (N_6316,N_3103,N_4848);
nor U6317 (N_6317,N_3276,N_784);
and U6318 (N_6318,N_1817,N_1719);
nor U6319 (N_6319,N_3497,N_128);
nor U6320 (N_6320,N_3275,N_1084);
and U6321 (N_6321,N_2276,N_782);
nand U6322 (N_6322,N_2048,N_1081);
or U6323 (N_6323,N_3047,N_4045);
and U6324 (N_6324,N_619,N_1618);
nor U6325 (N_6325,N_4475,N_717);
nor U6326 (N_6326,N_1515,N_1706);
or U6327 (N_6327,N_3658,N_522);
nor U6328 (N_6328,N_3888,N_1659);
and U6329 (N_6329,N_3293,N_1540);
nand U6330 (N_6330,N_3048,N_3822);
and U6331 (N_6331,N_2134,N_3422);
or U6332 (N_6332,N_2035,N_1105);
nand U6333 (N_6333,N_4728,N_92);
nand U6334 (N_6334,N_1848,N_4184);
and U6335 (N_6335,N_3544,N_3398);
nand U6336 (N_6336,N_4535,N_4);
and U6337 (N_6337,N_1073,N_986);
nand U6338 (N_6338,N_4476,N_4298);
nand U6339 (N_6339,N_3078,N_4662);
and U6340 (N_6340,N_1934,N_58);
nor U6341 (N_6341,N_2797,N_2192);
nand U6342 (N_6342,N_4846,N_4533);
nor U6343 (N_6343,N_4182,N_3492);
or U6344 (N_6344,N_2266,N_3313);
and U6345 (N_6345,N_525,N_3005);
xor U6346 (N_6346,N_4545,N_3975);
or U6347 (N_6347,N_4118,N_449);
nand U6348 (N_6348,N_2222,N_2714);
xnor U6349 (N_6349,N_157,N_3397);
nand U6350 (N_6350,N_2199,N_3668);
nor U6351 (N_6351,N_2504,N_3401);
nor U6352 (N_6352,N_430,N_1379);
nor U6353 (N_6353,N_1046,N_3400);
nand U6354 (N_6354,N_3845,N_4364);
or U6355 (N_6355,N_562,N_4720);
or U6356 (N_6356,N_2410,N_2119);
and U6357 (N_6357,N_4815,N_890);
and U6358 (N_6358,N_2961,N_4599);
xnor U6359 (N_6359,N_1122,N_1967);
and U6360 (N_6360,N_1983,N_4733);
xnor U6361 (N_6361,N_1206,N_4113);
nand U6362 (N_6362,N_1701,N_4286);
nand U6363 (N_6363,N_4814,N_1357);
and U6364 (N_6364,N_322,N_783);
nand U6365 (N_6365,N_144,N_4316);
nand U6366 (N_6366,N_3268,N_2089);
nand U6367 (N_6367,N_258,N_4471);
or U6368 (N_6368,N_3054,N_319);
nand U6369 (N_6369,N_1239,N_2683);
nand U6370 (N_6370,N_3696,N_2238);
nand U6371 (N_6371,N_4794,N_4675);
and U6372 (N_6372,N_4797,N_4301);
xor U6373 (N_6373,N_4899,N_2517);
and U6374 (N_6374,N_4305,N_813);
nand U6375 (N_6375,N_1254,N_1656);
or U6376 (N_6376,N_2994,N_3680);
nand U6377 (N_6377,N_136,N_2751);
and U6378 (N_6378,N_4169,N_3432);
and U6379 (N_6379,N_3415,N_3950);
and U6380 (N_6380,N_3646,N_3371);
or U6381 (N_6381,N_4214,N_724);
xnor U6382 (N_6382,N_115,N_4562);
nand U6383 (N_6383,N_2657,N_83);
nor U6384 (N_6384,N_3577,N_3923);
nand U6385 (N_6385,N_2173,N_1948);
or U6386 (N_6386,N_681,N_1513);
nor U6387 (N_6387,N_347,N_4416);
or U6388 (N_6388,N_2251,N_3734);
nand U6389 (N_6389,N_1676,N_2416);
nor U6390 (N_6390,N_2622,N_255);
or U6391 (N_6391,N_452,N_1500);
nor U6392 (N_6392,N_1454,N_3090);
and U6393 (N_6393,N_4859,N_112);
nand U6394 (N_6394,N_4997,N_1019);
nand U6395 (N_6395,N_3814,N_3063);
and U6396 (N_6396,N_1843,N_3781);
and U6397 (N_6397,N_4713,N_3527);
xor U6398 (N_6398,N_1830,N_1975);
and U6399 (N_6399,N_3280,N_4968);
nor U6400 (N_6400,N_2748,N_200);
and U6401 (N_6401,N_90,N_4539);
or U6402 (N_6402,N_2143,N_769);
or U6403 (N_6403,N_1422,N_2252);
and U6404 (N_6404,N_2708,N_2193);
or U6405 (N_6405,N_4731,N_3404);
or U6406 (N_6406,N_2890,N_4744);
and U6407 (N_6407,N_4615,N_2577);
or U6408 (N_6408,N_3443,N_723);
nand U6409 (N_6409,N_3713,N_4395);
nor U6410 (N_6410,N_3701,N_1639);
or U6411 (N_6411,N_2248,N_1453);
nand U6412 (N_6412,N_3636,N_424);
and U6413 (N_6413,N_1674,N_2008);
and U6414 (N_6414,N_4952,N_3613);
nor U6415 (N_6415,N_844,N_2436);
xnor U6416 (N_6416,N_2763,N_4369);
nor U6417 (N_6417,N_2398,N_2659);
nand U6418 (N_6418,N_501,N_4644);
and U6419 (N_6419,N_1307,N_4146);
nand U6420 (N_6420,N_2122,N_3507);
nor U6421 (N_6421,N_3706,N_1102);
nor U6422 (N_6422,N_3766,N_3802);
nor U6423 (N_6423,N_425,N_634);
nand U6424 (N_6424,N_2201,N_2220);
nor U6425 (N_6425,N_3758,N_2128);
and U6426 (N_6426,N_2702,N_2928);
and U6427 (N_6427,N_181,N_3936);
xnor U6428 (N_6428,N_2435,N_1956);
nand U6429 (N_6429,N_1445,N_1961);
xnor U6430 (N_6430,N_104,N_3184);
nor U6431 (N_6431,N_1298,N_4948);
and U6432 (N_6432,N_2551,N_4583);
or U6433 (N_6433,N_4088,N_4361);
nand U6434 (N_6434,N_1180,N_2145);
and U6435 (N_6435,N_1251,N_3897);
and U6436 (N_6436,N_4228,N_914);
or U6437 (N_6437,N_4342,N_2014);
nor U6438 (N_6438,N_819,N_4914);
nor U6439 (N_6439,N_3148,N_2731);
nor U6440 (N_6440,N_2383,N_2243);
or U6441 (N_6441,N_3350,N_3798);
and U6442 (N_6442,N_3905,N_4344);
and U6443 (N_6443,N_2327,N_3517);
and U6444 (N_6444,N_504,N_4153);
nor U6445 (N_6445,N_1930,N_1362);
and U6446 (N_6446,N_324,N_2426);
or U6447 (N_6447,N_1266,N_4053);
nor U6448 (N_6448,N_766,N_2245);
and U6449 (N_6449,N_569,N_2218);
nand U6450 (N_6450,N_779,N_1326);
xnor U6451 (N_6451,N_673,N_2332);
xnor U6452 (N_6452,N_485,N_95);
nor U6453 (N_6453,N_2621,N_4132);
or U6454 (N_6454,N_1638,N_2581);
or U6455 (N_6455,N_433,N_758);
nand U6456 (N_6456,N_2373,N_830);
xnor U6457 (N_6457,N_1125,N_3375);
nor U6458 (N_6458,N_2959,N_2673);
xor U6459 (N_6459,N_4558,N_3673);
or U6460 (N_6460,N_4643,N_2915);
nand U6461 (N_6461,N_3051,N_3360);
and U6462 (N_6462,N_487,N_1857);
nand U6463 (N_6463,N_3603,N_3460);
and U6464 (N_6464,N_2037,N_225);
or U6465 (N_6465,N_1933,N_578);
xnor U6466 (N_6466,N_3311,N_4048);
and U6467 (N_6467,N_3319,N_1555);
nand U6468 (N_6468,N_2209,N_3862);
nand U6469 (N_6469,N_3886,N_3857);
xor U6470 (N_6470,N_2430,N_4451);
or U6471 (N_6471,N_197,N_1559);
nand U6472 (N_6472,N_2580,N_2159);
xor U6473 (N_6473,N_205,N_4042);
nand U6474 (N_6474,N_3718,N_4494);
and U6475 (N_6475,N_2862,N_1200);
nor U6476 (N_6476,N_2590,N_4489);
nor U6477 (N_6477,N_1374,N_1270);
and U6478 (N_6478,N_2984,N_1124);
and U6479 (N_6479,N_2073,N_1306);
nand U6480 (N_6480,N_2114,N_1712);
or U6481 (N_6481,N_2139,N_4046);
nand U6482 (N_6482,N_1446,N_2045);
or U6483 (N_6483,N_3261,N_3518);
and U6484 (N_6484,N_354,N_4764);
nand U6485 (N_6485,N_2062,N_3142);
nand U6486 (N_6486,N_4503,N_4628);
nand U6487 (N_6487,N_2596,N_2144);
nor U6488 (N_6488,N_308,N_4775);
nand U6489 (N_6489,N_1861,N_1416);
nor U6490 (N_6490,N_1,N_4254);
and U6491 (N_6491,N_1752,N_1686);
nand U6492 (N_6492,N_3248,N_814);
or U6493 (N_6493,N_3797,N_298);
and U6494 (N_6494,N_3295,N_1927);
nor U6495 (N_6495,N_2914,N_69);
nor U6496 (N_6496,N_1343,N_2712);
nand U6497 (N_6497,N_1981,N_2287);
or U6498 (N_6498,N_2908,N_2516);
xnor U6499 (N_6499,N_230,N_1303);
nand U6500 (N_6500,N_1441,N_4262);
and U6501 (N_6501,N_2302,N_3392);
nand U6502 (N_6502,N_403,N_234);
or U6503 (N_6503,N_3602,N_866);
nor U6504 (N_6504,N_1172,N_3171);
nor U6505 (N_6505,N_2137,N_952);
nand U6506 (N_6506,N_1982,N_2406);
nor U6507 (N_6507,N_4410,N_2882);
nor U6508 (N_6508,N_857,N_237);
or U6509 (N_6509,N_4477,N_2682);
nand U6510 (N_6510,N_2140,N_119);
nor U6511 (N_6511,N_2219,N_4102);
or U6512 (N_6512,N_1269,N_4359);
nor U6513 (N_6513,N_4993,N_1636);
and U6514 (N_6514,N_510,N_3086);
and U6515 (N_6515,N_4631,N_4946);
and U6516 (N_6516,N_1205,N_3178);
nor U6517 (N_6517,N_3428,N_628);
and U6518 (N_6518,N_1766,N_3384);
and U6519 (N_6519,N_3997,N_3080);
nand U6520 (N_6520,N_3674,N_266);
nand U6521 (N_6521,N_2586,N_994);
nand U6522 (N_6522,N_2363,N_1549);
and U6523 (N_6523,N_2547,N_2991);
or U6524 (N_6524,N_4266,N_4576);
xnor U6525 (N_6525,N_2496,N_1872);
nor U6526 (N_6526,N_1428,N_4148);
and U6527 (N_6527,N_3088,N_3451);
nand U6528 (N_6528,N_698,N_2215);
and U6529 (N_6529,N_4840,N_2867);
nand U6530 (N_6530,N_3174,N_2040);
and U6531 (N_6531,N_3647,N_4398);
or U6532 (N_6532,N_2779,N_4682);
nand U6533 (N_6533,N_2573,N_2289);
nand U6534 (N_6534,N_4916,N_1818);
nand U6535 (N_6535,N_274,N_348);
and U6536 (N_6536,N_2897,N_263);
nand U6537 (N_6537,N_3019,N_1333);
nor U6538 (N_6538,N_3777,N_953);
or U6539 (N_6539,N_2206,N_1893);
and U6540 (N_6540,N_2920,N_3467);
nand U6541 (N_6541,N_1107,N_4594);
nand U6542 (N_6542,N_863,N_1763);
nand U6543 (N_6543,N_1588,N_3325);
nor U6544 (N_6544,N_605,N_2977);
nand U6545 (N_6545,N_123,N_4213);
nor U6546 (N_6546,N_4874,N_1061);
or U6547 (N_6547,N_218,N_781);
and U6548 (N_6548,N_4193,N_3844);
nand U6549 (N_6549,N_232,N_1152);
and U6550 (N_6550,N_855,N_4716);
xor U6551 (N_6551,N_1672,N_3034);
nor U6552 (N_6552,N_1756,N_4230);
nand U6553 (N_6553,N_4338,N_2009);
nand U6554 (N_6554,N_3724,N_3960);
and U6555 (N_6555,N_725,N_718);
and U6556 (N_6556,N_1489,N_2741);
or U6557 (N_6557,N_4871,N_3502);
nor U6558 (N_6558,N_2951,N_2001);
nand U6559 (N_6559,N_627,N_2690);
nor U6560 (N_6560,N_786,N_3444);
nor U6561 (N_6561,N_3804,N_4181);
xnor U6562 (N_6562,N_1233,N_2421);
and U6563 (N_6563,N_1300,N_1650);
nor U6564 (N_6564,N_632,N_910);
or U6565 (N_6565,N_4142,N_3911);
and U6566 (N_6566,N_4693,N_2946);
xnor U6567 (N_6567,N_3605,N_3305);
nor U6568 (N_6568,N_2764,N_2237);
and U6569 (N_6569,N_3554,N_3354);
and U6570 (N_6570,N_493,N_1867);
nor U6571 (N_6571,N_3588,N_2000);
xor U6572 (N_6572,N_1175,N_4609);
or U6573 (N_6573,N_3970,N_1408);
and U6574 (N_6574,N_4081,N_4391);
and U6575 (N_6575,N_2402,N_1785);
nand U6576 (N_6576,N_1826,N_2244);
nor U6577 (N_6577,N_2843,N_1693);
nand U6578 (N_6578,N_3678,N_2966);
or U6579 (N_6579,N_1671,N_2591);
nand U6580 (N_6580,N_2833,N_4706);
nor U6581 (N_6581,N_3192,N_1952);
and U6582 (N_6582,N_922,N_2999);
and U6583 (N_6583,N_1159,N_816);
nor U6584 (N_6584,N_4565,N_3152);
nor U6585 (N_6585,N_1569,N_1641);
nor U6586 (N_6586,N_1724,N_713);
or U6587 (N_6587,N_4205,N_4925);
nand U6588 (N_6588,N_1488,N_2609);
or U6589 (N_6589,N_3853,N_1621);
nand U6590 (N_6590,N_393,N_1011);
nor U6591 (N_6591,N_3880,N_2469);
xnor U6592 (N_6592,N_4703,N_720);
or U6593 (N_6593,N_555,N_4120);
and U6594 (N_6594,N_3177,N_3864);
or U6595 (N_6595,N_4279,N_2938);
or U6596 (N_6596,N_3769,N_2595);
and U6597 (N_6597,N_2538,N_1430);
or U6598 (N_6598,N_2113,N_4039);
nand U6599 (N_6599,N_1262,N_3378);
xnor U6600 (N_6600,N_1574,N_2576);
nor U6601 (N_6601,N_1086,N_3612);
xor U6602 (N_6602,N_3099,N_1670);
nor U6603 (N_6603,N_3077,N_772);
and U6604 (N_6604,N_4510,N_4223);
or U6605 (N_6605,N_2301,N_4367);
xnor U6606 (N_6606,N_3765,N_677);
and U6607 (N_6607,N_2982,N_4024);
and U6608 (N_6608,N_3775,N_4354);
or U6609 (N_6609,N_828,N_4891);
or U6610 (N_6610,N_2676,N_1697);
or U6611 (N_6611,N_4847,N_1969);
or U6612 (N_6612,N_108,N_3466);
nor U6613 (N_6613,N_498,N_2510);
or U6614 (N_6614,N_3849,N_2981);
and U6615 (N_6615,N_860,N_4002);
or U6616 (N_6616,N_3254,N_899);
nor U6617 (N_6617,N_4773,N_705);
nand U6618 (N_6618,N_1257,N_4483);
nor U6619 (N_6619,N_2507,N_1249);
xnor U6620 (N_6620,N_2979,N_3865);
nand U6621 (N_6621,N_3445,N_1151);
and U6622 (N_6622,N_183,N_3021);
and U6623 (N_6623,N_1284,N_2084);
nor U6624 (N_6624,N_3263,N_4210);
nor U6625 (N_6625,N_4913,N_3209);
nor U6626 (N_6626,N_2762,N_1230);
xnor U6627 (N_6627,N_4737,N_2395);
and U6628 (N_6628,N_2350,N_3520);
and U6629 (N_6629,N_4152,N_4380);
and U6630 (N_6630,N_2885,N_1509);
and U6631 (N_6631,N_4734,N_2965);
nand U6632 (N_6632,N_3127,N_1690);
nand U6633 (N_6633,N_1537,N_4602);
nor U6634 (N_6634,N_4249,N_1681);
and U6635 (N_6635,N_3024,N_2625);
or U6636 (N_6636,N_4076,N_3138);
nand U6637 (N_6637,N_4238,N_1318);
and U6638 (N_6638,N_4026,N_4650);
nand U6639 (N_6639,N_1977,N_1069);
xnor U6640 (N_6640,N_3869,N_3145);
nor U6641 (N_6641,N_1965,N_344);
or U6642 (N_6642,N_721,N_3271);
or U6643 (N_6643,N_787,N_2907);
or U6644 (N_6644,N_626,N_4629);
nand U6645 (N_6645,N_4735,N_383);
nor U6646 (N_6646,N_3689,N_3913);
nand U6647 (N_6647,N_545,N_4924);
nor U6648 (N_6648,N_4368,N_1234);
or U6649 (N_6649,N_4185,N_3176);
and U6650 (N_6650,N_812,N_4508);
and U6651 (N_6651,N_252,N_2125);
xnor U6652 (N_6652,N_552,N_3929);
nor U6653 (N_6653,N_3189,N_4320);
and U6654 (N_6654,N_1625,N_3908);
nor U6655 (N_6655,N_4908,N_3509);
and U6656 (N_6656,N_2886,N_2013);
nor U6657 (N_6657,N_457,N_2438);
and U6658 (N_6658,N_3490,N_3932);
nand U6659 (N_6659,N_3146,N_3790);
nand U6660 (N_6660,N_4492,N_3023);
nand U6661 (N_6661,N_685,N_4237);
or U6662 (N_6662,N_4977,N_1468);
or U6663 (N_6663,N_3672,N_1810);
nand U6664 (N_6664,N_3100,N_4491);
and U6665 (N_6665,N_4408,N_2490);
or U6666 (N_6666,N_481,N_3072);
and U6667 (N_6667,N_2115,N_3162);
or U6668 (N_6668,N_818,N_4428);
and U6669 (N_6669,N_3545,N_3222);
or U6670 (N_6670,N_44,N_519);
nor U6671 (N_6671,N_2054,N_4326);
nand U6672 (N_6672,N_469,N_4216);
nor U6673 (N_6673,N_2371,N_2458);
nand U6674 (N_6674,N_1481,N_2587);
xor U6675 (N_6675,N_2056,N_4837);
and U6676 (N_6676,N_4130,N_1644);
nand U6677 (N_6677,N_4531,N_992);
nor U6678 (N_6678,N_176,N_4520);
nand U6679 (N_6679,N_2641,N_2620);
and U6680 (N_6680,N_3625,N_454);
nand U6681 (N_6681,N_1845,N_3942);
or U6682 (N_6682,N_4055,N_1120);
nand U6683 (N_6683,N_3083,N_4995);
nand U6684 (N_6684,N_2303,N_3257);
nand U6685 (N_6685,N_1090,N_739);
and U6686 (N_6686,N_2116,N_832);
or U6687 (N_6687,N_700,N_1173);
or U6688 (N_6688,N_4289,N_534);
and U6689 (N_6689,N_4197,N_2275);
nor U6690 (N_6690,N_1372,N_3662);
or U6691 (N_6691,N_4918,N_927);
nand U6692 (N_6692,N_4327,N_827);
or U6693 (N_6693,N_4618,N_1976);
nor U6694 (N_6694,N_4123,N_1190);
xor U6695 (N_6695,N_4069,N_39);
nor U6696 (N_6696,N_402,N_1884);
nand U6697 (N_6697,N_3949,N_702);
xor U6698 (N_6698,N_1525,N_4630);
nor U6699 (N_6699,N_4697,N_3902);
and U6700 (N_6700,N_3735,N_2985);
nand U6701 (N_6701,N_85,N_1014);
and U6702 (N_6702,N_4245,N_4206);
nor U6703 (N_6703,N_4517,N_1823);
nor U6704 (N_6704,N_1344,N_1564);
xnor U6705 (N_6705,N_2921,N_4061);
nor U6706 (N_6706,N_1138,N_3377);
nand U6707 (N_6707,N_1836,N_2118);
and U6708 (N_6708,N_4236,N_4904);
nand U6709 (N_6709,N_2868,N_304);
nand U6710 (N_6710,N_2304,N_4006);
and U6711 (N_6711,N_2783,N_554);
xnor U6712 (N_6712,N_2554,N_2038);
or U6713 (N_6713,N_126,N_4930);
or U6714 (N_6714,N_3542,N_3984);
or U6715 (N_6715,N_2841,N_1015);
nand U6716 (N_6716,N_2798,N_3373);
xnor U6717 (N_6717,N_1842,N_2560);
nor U6718 (N_6718,N_1252,N_1876);
nor U6719 (N_6719,N_2094,N_2784);
nor U6720 (N_6720,N_315,N_1349);
and U6721 (N_6721,N_4441,N_824);
xnor U6722 (N_6722,N_4636,N_4897);
and U6723 (N_6723,N_2481,N_3589);
nand U6724 (N_6724,N_339,N_3835);
nand U6725 (N_6725,N_196,N_3068);
and U6726 (N_6726,N_4143,N_1698);
or U6727 (N_6727,N_1771,N_3240);
nand U6728 (N_6728,N_1571,N_3131);
nor U6729 (N_6729,N_247,N_869);
nor U6730 (N_6730,N_3475,N_1831);
xnor U6731 (N_6731,N_730,N_1053);
and U6732 (N_6732,N_1008,N_2643);
or U6733 (N_6733,N_4998,N_3308);
nor U6734 (N_6734,N_3335,N_2931);
and U6735 (N_6735,N_1415,N_2501);
nor U6736 (N_6736,N_4360,N_4567);
and U6737 (N_6737,N_2420,N_537);
or U6738 (N_6738,N_4634,N_192);
or U6739 (N_6739,N_3198,N_3875);
nand U6740 (N_6740,N_1611,N_3408);
and U6741 (N_6741,N_4013,N_622);
nor U6742 (N_6742,N_2793,N_4242);
and U6743 (N_6743,N_374,N_2849);
or U6744 (N_6744,N_3190,N_2349);
and U6745 (N_6745,N_435,N_3393);
nand U6746 (N_6746,N_2860,N_4894);
or U6747 (N_6747,N_1592,N_2256);
and U6748 (N_6748,N_2796,N_2939);
or U6749 (N_6749,N_1080,N_496);
or U6750 (N_6750,N_1000,N_4373);
nor U6751 (N_6751,N_3028,N_1116);
xor U6752 (N_6752,N_2733,N_513);
or U6753 (N_6753,N_670,N_1006);
nand U6754 (N_6754,N_2669,N_305);
or U6755 (N_6755,N_1048,N_4707);
and U6756 (N_6756,N_3332,N_1246);
or U6757 (N_6757,N_822,N_701);
xnor U6758 (N_6758,N_1945,N_2217);
nor U6759 (N_6759,N_4011,N_2645);
and U6760 (N_6760,N_3896,N_1026);
and U6761 (N_6761,N_1702,N_3534);
nor U6762 (N_6762,N_2031,N_4091);
nand U6763 (N_6763,N_53,N_4299);
or U6764 (N_6764,N_1558,N_3633);
nor U6765 (N_6765,N_2423,N_2079);
xor U6766 (N_6766,N_3726,N_1536);
or U6767 (N_6767,N_4909,N_1794);
or U6768 (N_6768,N_4732,N_936);
or U6769 (N_6769,N_4676,N_1039);
and U6770 (N_6770,N_362,N_1255);
nand U6771 (N_6771,N_815,N_138);
nand U6772 (N_6772,N_542,N_4419);
nor U6773 (N_6773,N_3157,N_1870);
nor U6774 (N_6774,N_1079,N_4957);
and U6775 (N_6775,N_3957,N_919);
and U6776 (N_6776,N_2615,N_3238);
nor U6777 (N_6777,N_4578,N_3922);
xnor U6778 (N_6778,N_3411,N_4621);
or U6779 (N_6779,N_642,N_4034);
and U6780 (N_6780,N_499,N_4096);
nor U6781 (N_6781,N_1833,N_4858);
nor U6782 (N_6782,N_4862,N_3681);
nor U6783 (N_6783,N_2136,N_2382);
or U6784 (N_6784,N_4934,N_261);
nand U6785 (N_6785,N_557,N_1709);
or U6786 (N_6786,N_2839,N_2772);
and U6787 (N_6787,N_191,N_1356);
nand U6788 (N_6788,N_2646,N_1595);
or U6789 (N_6789,N_4516,N_1404);
nand U6790 (N_6790,N_2976,N_686);
nand U6791 (N_6791,N_2334,N_3558);
and U6792 (N_6792,N_2309,N_1993);
xnor U6793 (N_6793,N_4661,N_423);
nor U6794 (N_6794,N_4271,N_2987);
or U6795 (N_6795,N_4694,N_4770);
or U6796 (N_6796,N_3060,N_4692);
nor U6797 (N_6797,N_3027,N_2165);
nand U6798 (N_6798,N_3985,N_2385);
and U6799 (N_6799,N_228,N_3891);
and U6800 (N_6800,N_3298,N_2188);
nor U6801 (N_6801,N_4579,N_4114);
nor U6802 (N_6802,N_4739,N_3001);
nand U6803 (N_6803,N_958,N_1272);
xnor U6804 (N_6804,N_436,N_1483);
nand U6805 (N_6805,N_3013,N_3052);
and U6806 (N_6806,N_2455,N_4743);
nand U6807 (N_6807,N_3618,N_318);
or U6808 (N_6808,N_512,N_1322);
and U6809 (N_6809,N_3283,N_1928);
and U6810 (N_6810,N_4965,N_3890);
nand U6811 (N_6811,N_1989,N_4372);
xor U6812 (N_6812,N_2092,N_473);
nor U6813 (N_6813,N_4154,N_4234);
or U6814 (N_6814,N_2552,N_272);
nor U6815 (N_6815,N_3528,N_4987);
xnor U6816 (N_6816,N_1722,N_1456);
and U6817 (N_6817,N_3575,N_4507);
and U6818 (N_6818,N_585,N_672);
nand U6819 (N_6819,N_3906,N_2539);
or U6820 (N_6820,N_2412,N_4547);
nand U6821 (N_6821,N_2202,N_694);
or U6822 (N_6822,N_3513,N_4803);
nand U6823 (N_6823,N_722,N_43);
and U6824 (N_6824,N_1236,N_3676);
and U6825 (N_6825,N_1355,N_2470);
or U6826 (N_6826,N_3399,N_2474);
or U6827 (N_6827,N_1463,N_2837);
nand U6828 (N_6828,N_1704,N_3161);
nor U6829 (N_6829,N_1528,N_132);
nor U6830 (N_6830,N_3850,N_1532);
nand U6831 (N_6831,N_4224,N_933);
xnor U6832 (N_6832,N_2102,N_4617);
nor U6833 (N_6833,N_4458,N_4873);
nand U6834 (N_6834,N_843,N_4443);
or U6835 (N_6835,N_387,N_1450);
and U6836 (N_6836,N_432,N_1476);
nand U6837 (N_6837,N_2522,N_3856);
xor U6838 (N_6838,N_1506,N_4875);
nand U6839 (N_6839,N_3671,N_1727);
nand U6840 (N_6840,N_56,N_1774);
or U6841 (N_6841,N_1078,N_2071);
or U6842 (N_6842,N_77,N_1978);
nand U6843 (N_6843,N_2883,N_2947);
xor U6844 (N_6844,N_3288,N_4173);
and U6845 (N_6845,N_4115,N_4108);
nor U6846 (N_6846,N_3774,N_2559);
nor U6847 (N_6847,N_2996,N_1577);
or U6848 (N_6848,N_2700,N_2036);
nand U6849 (N_6849,N_3770,N_4927);
and U6850 (N_6850,N_3339,N_3031);
and U6851 (N_6851,N_2974,N_1695);
and U6852 (N_6852,N_2322,N_1274);
nor U6853 (N_6853,N_2434,N_4017);
nand U6854 (N_6854,N_3815,N_2929);
or U6855 (N_6855,N_3744,N_4960);
or U6856 (N_6856,N_4499,N_4950);
and U6857 (N_6857,N_4979,N_2639);
and U6858 (N_6858,N_1563,N_972);
nor U6859 (N_6859,N_1218,N_4105);
nand U6860 (N_6860,N_3559,N_4680);
nand U6861 (N_6861,N_1094,N_3637);
nor U6862 (N_6862,N_2728,N_1647);
and U6863 (N_6863,N_4396,N_2221);
nand U6864 (N_6864,N_3061,N_896);
or U6865 (N_6865,N_4059,N_3995);
nand U6866 (N_6866,N_1895,N_4384);
and U6867 (N_6867,N_2263,N_3786);
nand U6868 (N_6868,N_4382,N_2834);
nand U6869 (N_6869,N_1130,N_4769);
and U6870 (N_6870,N_4066,N_3331);
nor U6871 (N_6871,N_4710,N_4317);
or U6872 (N_6872,N_4116,N_505);
or U6873 (N_6873,N_625,N_3746);
and U6874 (N_6874,N_582,N_4390);
nand U6875 (N_6875,N_892,N_1723);
nand U6876 (N_6876,N_2442,N_2320);
and U6877 (N_6877,N_4314,N_2034);
or U6878 (N_6878,N_4889,N_2533);
or U6879 (N_6879,N_3440,N_94);
or U6880 (N_6880,N_957,N_290);
nor U6881 (N_6881,N_3851,N_4394);
nor U6882 (N_6882,N_1276,N_1874);
nor U6883 (N_6883,N_4052,N_73);
and U6884 (N_6884,N_1045,N_553);
nand U6885 (N_6885,N_188,N_210);
nand U6886 (N_6886,N_3372,N_897);
nor U6887 (N_6887,N_4595,N_2086);
nor U6888 (N_6888,N_3463,N_78);
xor U6889 (N_6889,N_4325,N_973);
nand U6890 (N_6890,N_2912,N_847);
nand U6891 (N_6891,N_4292,N_2106);
nand U6892 (N_6892,N_244,N_3278);
nor U6893 (N_6893,N_3593,N_145);
and U6894 (N_6894,N_3388,N_3993);
nor U6895 (N_6895,N_4760,N_4941);
and U6896 (N_6896,N_2719,N_1003);
or U6897 (N_6897,N_1329,N_893);
nor U6898 (N_6898,N_4845,N_79);
xor U6899 (N_6899,N_3282,N_3082);
nand U6900 (N_6900,N_1545,N_2411);
nand U6901 (N_6901,N_2324,N_3344);
and U6902 (N_6902,N_4962,N_4804);
nand U6903 (N_6903,N_805,N_2795);
nand U6904 (N_6904,N_2502,N_4806);
or U6905 (N_6905,N_3514,N_3939);
nand U6906 (N_6906,N_3827,N_3226);
and U6907 (N_6907,N_4480,N_4910);
nand U6908 (N_6908,N_2818,N_2887);
xor U6909 (N_6909,N_1959,N_1527);
or U6910 (N_6910,N_1361,N_3816);
nand U6911 (N_6911,N_2378,N_753);
or U6912 (N_6912,N_1128,N_838);
or U6913 (N_6913,N_2232,N_2292);
nor U6914 (N_6914,N_2342,N_1924);
nand U6915 (N_6915,N_3307,N_2935);
and U6916 (N_6916,N_3237,N_3561);
or U6917 (N_6917,N_3447,N_4978);
or U6918 (N_6918,N_303,N_3754);
or U6919 (N_6919,N_4239,N_1809);
nor U6920 (N_6920,N_4782,N_777);
or U6921 (N_6921,N_762,N_2069);
and U6922 (N_6922,N_1170,N_4086);
and U6923 (N_6923,N_4005,N_3429);
and U6924 (N_6924,N_2120,N_2425);
and U6925 (N_6925,N_1075,N_146);
or U6926 (N_6926,N_1721,N_1634);
nand U6927 (N_6927,N_392,N_2466);
and U6928 (N_6928,N_350,N_675);
nand U6929 (N_6929,N_4149,N_3983);
nand U6930 (N_6930,N_1387,N_2865);
and U6931 (N_6931,N_4677,N_774);
or U6932 (N_6932,N_4688,N_413);
nand U6933 (N_6933,N_3205,N_2154);
and U6934 (N_6934,N_2605,N_4885);
xor U6935 (N_6935,N_3304,N_2282);
and U6936 (N_6936,N_3158,N_2121);
nand U6937 (N_6937,N_233,N_2716);
nor U6938 (N_6938,N_3811,N_3639);
nor U6939 (N_6939,N_124,N_2064);
and U6940 (N_6940,N_3095,N_1685);
or U6941 (N_6941,N_2235,N_4400);
nand U6942 (N_6942,N_2047,N_4923);
and U6943 (N_6943,N_301,N_1033);
or U6944 (N_6944,N_4973,N_4399);
xnor U6945 (N_6945,N_2941,N_3963);
and U6946 (N_6946,N_1384,N_4928);
nor U6947 (N_6947,N_3757,N_715);
nand U6948 (N_6948,N_4198,N_4796);
or U6949 (N_6949,N_2536,N_1744);
or U6950 (N_6950,N_1947,N_2242);
xor U6951 (N_6951,N_3245,N_4212);
or U6952 (N_6952,N_2405,N_4931);
nand U6953 (N_6953,N_2919,N_1219);
nand U6954 (N_6954,N_4537,N_4486);
nor U6955 (N_6955,N_419,N_599);
nor U6956 (N_6956,N_911,N_1932);
and U6957 (N_6957,N_495,N_1378);
xor U6958 (N_6958,N_3541,N_1440);
nor U6959 (N_6959,N_4607,N_4140);
xnor U6960 (N_6960,N_327,N_3419);
or U6961 (N_6961,N_4620,N_3833);
or U6962 (N_6962,N_2934,N_2835);
nand U6963 (N_6963,N_4994,N_1741);
and U6964 (N_6964,N_2341,N_691);
nand U6965 (N_6965,N_1012,N_2903);
or U6966 (N_6966,N_895,N_594);
and U6967 (N_6967,N_1951,N_3799);
or U6968 (N_6968,N_4164,N_1898);
or U6969 (N_6969,N_3345,N_2530);
or U6970 (N_6970,N_734,N_4658);
nor U6971 (N_6971,N_291,N_4465);
nand U6972 (N_6972,N_2067,N_2176);
or U6973 (N_6973,N_3175,N_2930);
xor U6974 (N_6974,N_1256,N_4854);
and U6975 (N_6975,N_1156,N_3900);
xnor U6976 (N_6976,N_3498,N_2277);
or U6977 (N_6977,N_1891,N_1132);
nand U6978 (N_6978,N_4781,N_4839);
and U6979 (N_6979,N_4422,N_3860);
and U6980 (N_6980,N_3683,N_203);
nand U6981 (N_6981,N_4493,N_4919);
and U6982 (N_6982,N_3049,N_1350);
or U6983 (N_6983,N_3737,N_3041);
nor U6984 (N_6984,N_114,N_3107);
nand U6985 (N_6985,N_294,N_776);
xnor U6986 (N_6986,N_2611,N_23);
nand U6987 (N_6987,N_2291,N_68);
and U6988 (N_6988,N_2328,N_2892);
nand U6989 (N_6989,N_4085,N_1757);
xor U6990 (N_6990,N_1182,N_4488);
and U6991 (N_6991,N_1713,N_147);
and U6992 (N_6992,N_1457,N_3991);
and U6993 (N_6993,N_2515,N_924);
and U6994 (N_6994,N_1485,N_169);
or U6995 (N_6995,N_86,N_4335);
nand U6996 (N_6996,N_2561,N_664);
and U6997 (N_6997,N_4233,N_2792);
xnor U6998 (N_6998,N_4649,N_2164);
nor U6999 (N_6999,N_4240,N_51);
or U7000 (N_7000,N_295,N_4183);
nand U7001 (N_7001,N_1546,N_2723);
and U7002 (N_7002,N_372,N_2758);
nand U7003 (N_7003,N_959,N_2585);
xor U7004 (N_7004,N_989,N_3788);
and U7005 (N_7005,N_2813,N_4550);
nand U7006 (N_7006,N_3572,N_750);
or U7007 (N_7007,N_4915,N_3809);
or U7008 (N_7008,N_3442,N_268);
nor U7009 (N_7009,N_2393,N_4362);
nand U7010 (N_7010,N_945,N_3930);
xor U7011 (N_7011,N_4138,N_2785);
or U7012 (N_7012,N_2508,N_850);
and U7013 (N_7013,N_2623,N_1114);
and U7014 (N_7014,N_67,N_4673);
nor U7015 (N_7015,N_142,N_3931);
or U7016 (N_7016,N_4251,N_3516);
xnor U7017 (N_7017,N_1163,N_359);
nand U7018 (N_7018,N_2697,N_3756);
nand U7019 (N_7019,N_3968,N_370);
and U7020 (N_7020,N_2648,N_592);
nor U7021 (N_7021,N_4351,N_1883);
nand U7022 (N_7022,N_1973,N_1142);
nor U7023 (N_7023,N_3185,N_2601);
nor U7024 (N_7024,N_4765,N_75);
or U7025 (N_7025,N_4285,N_1092);
nor U7026 (N_7026,N_3743,N_1740);
nand U7027 (N_7027,N_4093,N_2780);
and U7028 (N_7028,N_2271,N_825);
nand U7029 (N_7029,N_364,N_4107);
and U7030 (N_7030,N_1035,N_3379);
nor U7031 (N_7031,N_2486,N_2879);
nand U7032 (N_7032,N_507,N_3998);
nor U7033 (N_7033,N_2058,N_3785);
nand U7034 (N_7034,N_611,N_3664);
nor U7035 (N_7035,N_4761,N_4684);
nor U7036 (N_7036,N_864,N_3361);
and U7037 (N_7037,N_2752,N_4912);
nand U7038 (N_7038,N_1699,N_1799);
or U7039 (N_7039,N_3761,N_3965);
and U7040 (N_7040,N_2732,N_3273);
and U7041 (N_7041,N_3216,N_674);
or U7042 (N_7042,N_133,N_949);
nand U7043 (N_7043,N_4805,N_3033);
and U7044 (N_7044,N_3617,N_2281);
xnor U7045 (N_7045,N_997,N_4664);
nor U7046 (N_7046,N_2806,N_2568);
and U7047 (N_7047,N_886,N_415);
xor U7048 (N_7048,N_3720,N_4795);
and U7049 (N_7049,N_3648,N_2654);
xnor U7050 (N_7050,N_4817,N_4608);
nand U7051 (N_7051,N_3874,N_1859);
or U7052 (N_7052,N_2207,N_346);
or U7053 (N_7053,N_743,N_1289);
nor U7054 (N_7054,N_3928,N_3529);
nor U7055 (N_7055,N_4003,N_2104);
or U7056 (N_7056,N_361,N_4311);
nand U7057 (N_7057,N_3499,N_4652);
nand U7058 (N_7058,N_3201,N_663);
xor U7059 (N_7059,N_4196,N_707);
nor U7060 (N_7060,N_3511,N_3299);
nor U7061 (N_7061,N_42,N_289);
nand U7062 (N_7062,N_4099,N_4699);
nand U7063 (N_7063,N_3793,N_3494);
xor U7064 (N_7064,N_3601,N_2297);
or U7065 (N_7065,N_3310,N_2902);
and U7066 (N_7066,N_2766,N_4745);
or U7067 (N_7067,N_1714,N_3421);
and U7068 (N_7068,N_2012,N_3244);
and U7069 (N_7069,N_1199,N_4009);
and U7070 (N_7070,N_1935,N_1811);
and U7071 (N_7071,N_1455,N_2022);
nand U7072 (N_7072,N_3040,N_4172);
or U7073 (N_7073,N_2936,N_2997);
nor U7074 (N_7074,N_3303,N_2010);
and U7075 (N_7075,N_1185,N_1363);
nand U7076 (N_7076,N_2312,N_4588);
and U7077 (N_7077,N_17,N_28);
xor U7078 (N_7078,N_3580,N_4566);
or U7079 (N_7079,N_4813,N_1668);
nor U7080 (N_7080,N_1087,N_1337);
and U7081 (N_7081,N_3227,N_1566);
nor U7082 (N_7082,N_163,N_4474);
nand U7083 (N_7083,N_3753,N_2687);
xor U7084 (N_7084,N_2901,N_4639);
nand U7085 (N_7085,N_4133,N_2910);
nand U7086 (N_7086,N_1193,N_2749);
and U7087 (N_7087,N_1354,N_4041);
xor U7088 (N_7088,N_1753,N_4985);
or U7089 (N_7089,N_379,N_3316);
or U7090 (N_7090,N_1283,N_854);
nor U7091 (N_7091,N_458,N_4243);
or U7092 (N_7092,N_3656,N_964);
or U7093 (N_7093,N_2258,N_851);
and U7094 (N_7094,N_3578,N_2437);
nor U7095 (N_7095,N_185,N_4538);
and U7096 (N_7096,N_4868,N_4147);
or U7097 (N_7097,N_1360,N_3599);
and U7098 (N_7098,N_3366,N_1578);
nor U7099 (N_7099,N_2880,N_2488);
nor U7100 (N_7100,N_300,N_2167);
nor U7101 (N_7101,N_204,N_4603);
nand U7102 (N_7102,N_2082,N_3553);
or U7103 (N_7103,N_48,N_3210);
and U7104 (N_7104,N_3329,N_4907);
and U7105 (N_7105,N_3679,N_1158);
and U7106 (N_7106,N_3547,N_2006);
nand U7107 (N_7107,N_4211,N_173);
nor U7108 (N_7108,N_4356,N_4654);
nand U7109 (N_7109,N_4449,N_1042);
or U7110 (N_7110,N_737,N_445);
or U7111 (N_7111,N_2503,N_351);
and U7112 (N_7112,N_3241,N_2664);
and U7113 (N_7113,N_1009,N_4036);
or U7114 (N_7114,N_1277,N_2534);
xnor U7115 (N_7115,N_342,N_2123);
nor U7116 (N_7116,N_1589,N_4536);
nand U7117 (N_7117,N_3533,N_64);
nor U7118 (N_7118,N_2389,N_4405);
nand U7119 (N_7119,N_2160,N_4119);
xor U7120 (N_7120,N_3657,N_661);
nand U7121 (N_7121,N_3135,N_3996);
nand U7122 (N_7122,N_1562,N_1153);
nand U7123 (N_7123,N_1877,N_4259);
xor U7124 (N_7124,N_2400,N_4446);
and U7125 (N_7125,N_1247,N_3584);
nand U7126 (N_7126,N_4426,N_4067);
and U7127 (N_7127,N_2513,N_3483);
nor U7128 (N_7128,N_2260,N_4062);
nand U7129 (N_7129,N_2909,N_1950);
and U7130 (N_7130,N_1846,N_785);
and U7131 (N_7131,N_2715,N_4177);
and U7132 (N_7132,N_2482,N_3586);
or U7133 (N_7133,N_1805,N_2077);
and U7134 (N_7134,N_2853,N_2583);
and U7135 (N_7135,N_1860,N_3476);
nand U7136 (N_7136,N_719,N_2847);
nand U7137 (N_7137,N_1312,N_4057);
or U7138 (N_7138,N_2603,N_34);
nand U7139 (N_7139,N_332,N_1204);
or U7140 (N_7140,N_2566,N_158);
nand U7141 (N_7141,N_2584,N_464);
xor U7142 (N_7142,N_2362,N_2898);
or U7143 (N_7143,N_802,N_2662);
or U7144 (N_7144,N_3818,N_1196);
nand U7145 (N_7145,N_1683,N_4220);
nor U7146 (N_7146,N_4556,N_666);
or U7147 (N_7147,N_1798,N_3281);
nand U7148 (N_7148,N_3155,N_3660);
and U7149 (N_7149,N_3728,N_1474);
nor U7150 (N_7150,N_120,N_760);
or U7151 (N_7151,N_3058,N_2973);
or U7152 (N_7152,N_1637,N_243);
or U7153 (N_7153,N_323,N_1007);
nand U7154 (N_7154,N_2476,N_3977);
or U7155 (N_7155,N_912,N_1301);
nand U7156 (N_7156,N_365,N_4403);
nand U7157 (N_7157,N_2152,N_1653);
nand U7158 (N_7158,N_3139,N_3831);
or U7159 (N_7159,N_4614,N_431);
nand U7160 (N_7160,N_3992,N_2582);
xor U7161 (N_7161,N_2877,N_2990);
nand U7162 (N_7162,N_2563,N_229);
xnor U7163 (N_7163,N_2449,N_601);
nand U7164 (N_7164,N_1616,N_201);
nand U7165 (N_7165,N_4611,N_2610);
or U7166 (N_7166,N_1285,N_4004);
nand U7167 (N_7167,N_1603,N_3649);
nand U7168 (N_7168,N_1619,N_1402);
nor U7169 (N_7169,N_3104,N_2424);
and U7170 (N_7170,N_565,N_614);
nor U7171 (N_7171,N_195,N_1103);
or U7172 (N_7172,N_1942,N_680);
or U7173 (N_7173,N_951,N_1664);
or U7174 (N_7174,N_3666,N_3124);
nor U7175 (N_7175,N_2003,N_3594);
or U7176 (N_7176,N_2041,N_563);
and U7177 (N_7177,N_1286,N_299);
nor U7178 (N_7178,N_2634,N_1718);
and U7179 (N_7179,N_2088,N_4810);
xor U7180 (N_7180,N_1064,N_1074);
nand U7181 (N_7181,N_2804,N_4687);
nand U7182 (N_7182,N_1980,N_3565);
and U7183 (N_7183,N_1878,N_2704);
xor U7184 (N_7184,N_898,N_3217);
or U7185 (N_7185,N_343,N_2184);
nor U7186 (N_7186,N_2699,N_4414);
and U7187 (N_7187,N_4275,N_4297);
nor U7188 (N_7188,N_2678,N_1066);
nand U7189 (N_7189,N_3783,N_559);
or U7190 (N_7190,N_154,N_656);
nand U7191 (N_7191,N_2616,N_21);
and U7192 (N_7192,N_1297,N_135);
nor U7193 (N_7193,N_3420,N_887);
nand U7194 (N_7194,N_2628,N_874);
and U7195 (N_7195,N_939,N_3425);
nor U7196 (N_7196,N_4969,N_241);
and U7197 (N_7197,N_45,N_529);
xor U7198 (N_7198,N_4073,N_3526);
nand U7199 (N_7199,N_170,N_1910);
nand U7200 (N_7200,N_4601,N_4518);
nor U7201 (N_7201,N_2317,N_1992);
nand U7202 (N_7202,N_1663,N_600);
and U7203 (N_7203,N_2824,N_4767);
nand U7204 (N_7204,N_4165,N_1737);
nand U7205 (N_7205,N_4482,N_590);
xor U7206 (N_7206,N_2918,N_4263);
nor U7207 (N_7207,N_4700,N_4389);
or U7208 (N_7208,N_604,N_524);
nand U7209 (N_7209,N_4816,N_711);
nand U7210 (N_7210,N_538,N_2250);
nor U7211 (N_7211,N_4365,N_4440);
nor U7212 (N_7212,N_1187,N_1834);
nand U7213 (N_7213,N_3622,N_3812);
nand U7214 (N_7214,N_328,N_1382);
nand U7215 (N_7215,N_1579,N_1840);
nand U7216 (N_7216,N_4282,N_3488);
nor U7217 (N_7217,N_1533,N_3885);
xnor U7218 (N_7218,N_1733,N_2725);
or U7219 (N_7219,N_2706,N_806);
and U7220 (N_7220,N_3106,N_1100);
or U7221 (N_7221,N_194,N_3125);
and U7222 (N_7222,N_3233,N_1044);
and U7223 (N_7223,N_2042,N_265);
nand U7224 (N_7224,N_4328,N_152);
nand U7225 (N_7225,N_4715,N_1963);
and U7226 (N_7226,N_969,N_2261);
or U7227 (N_7227,N_3813,N_4376);
and U7228 (N_7228,N_3407,N_220);
nand U7229 (N_7229,N_4656,N_1988);
or U7230 (N_7230,N_2635,N_1351);
nand U7231 (N_7231,N_4853,N_3102);
nand U7232 (N_7232,N_3374,N_4560);
nor U7233 (N_7233,N_620,N_916);
or U7234 (N_7234,N_4509,N_2177);
and U7235 (N_7235,N_4786,N_2494);
xnor U7236 (N_7236,N_3522,N_591);
nor U7237 (N_7237,N_3776,N_597);
or U7238 (N_7238,N_18,N_31);
or U7239 (N_7239,N_4892,N_885);
and U7240 (N_7240,N_3762,N_2203);
nand U7241 (N_7241,N_550,N_2403);
and U7242 (N_7242,N_1828,N_4330);
nor U7243 (N_7243,N_962,N_998);
nand U7244 (N_7244,N_4886,N_2848);
or U7245 (N_7245,N_3893,N_4265);
nand U7246 (N_7246,N_3438,N_4357);
xnor U7247 (N_7247,N_4163,N_4585);
nor U7248 (N_7248,N_3324,N_2557);
xnor U7249 (N_7249,N_3708,N_398);
nor U7250 (N_7250,N_1807,N_861);
or U7251 (N_7251,N_1258,N_2696);
nand U7252 (N_7252,N_3141,N_3418);
nand U7253 (N_7253,N_1108,N_3294);
nand U7254 (N_7254,N_2760,N_1482);
and U7255 (N_7255,N_2135,N_2790);
nor U7256 (N_7256,N_3693,N_3367);
nand U7257 (N_7257,N_2674,N_506);
nand U7258 (N_7258,N_262,N_4638);
nor U7259 (N_7259,N_3389,N_4135);
nand U7260 (N_7260,N_3225,N_3212);
nor U7261 (N_7261,N_4097,N_2170);
and U7262 (N_7262,N_925,N_967);
nor U7263 (N_7263,N_610,N_1944);
or U7264 (N_7264,N_1227,N_417);
or U7265 (N_7265,N_1749,N_3986);
nor U7266 (N_7266,N_1390,N_1800);
nand U7267 (N_7267,N_2313,N_2937);
or U7268 (N_7268,N_1091,N_231);
or U7269 (N_7269,N_517,N_390);
or U7270 (N_7270,N_2812,N_2180);
nand U7271 (N_7271,N_3504,N_817);
nand U7272 (N_7272,N_3876,N_4640);
and U7273 (N_7273,N_1041,N_1202);
or U7274 (N_7274,N_4597,N_1119);
or U7275 (N_7275,N_2274,N_1192);
nand U7276 (N_7276,N_1438,N_1917);
or U7277 (N_7277,N_9,N_466);
nor U7278 (N_7278,N_1338,N_1691);
xor U7279 (N_7279,N_2956,N_2138);
or U7280 (N_7280,N_3286,N_2198);
nor U7281 (N_7281,N_4229,N_775);
and U7282 (N_7282,N_1377,N_3110);
or U7283 (N_7283,N_400,N_3738);
nor U7284 (N_7284,N_1271,N_1943);
nand U7285 (N_7285,N_3951,N_4570);
xor U7286 (N_7286,N_1966,N_3441);
nor U7287 (N_7287,N_729,N_2876);
and U7288 (N_7288,N_840,N_3341);
or U7289 (N_7289,N_4974,N_441);
nand U7290 (N_7290,N_1795,N_2556);
nor U7291 (N_7291,N_3489,N_3763);
or U7292 (N_7292,N_148,N_1104);
and U7293 (N_7293,N_4090,N_2174);
or U7294 (N_7294,N_1191,N_640);
nor U7295 (N_7295,N_5,N_3037);
or U7296 (N_7296,N_2376,N_2417);
nand U7297 (N_7297,N_2070,N_1519);
and U7298 (N_7298,N_4880,N_2528);
nor U7299 (N_7299,N_540,N_1929);
and U7300 (N_7300,N_714,N_2443);
nand U7301 (N_7301,N_472,N_3741);
or U7302 (N_7302,N_521,N_446);
and U7303 (N_7303,N_918,N_2597);
and U7304 (N_7304,N_4103,N_2208);
xnor U7305 (N_7305,N_4122,N_3260);
xnor U7306 (N_7306,N_1544,N_3409);
nand U7307 (N_7307,N_4032,N_4549);
nor U7308 (N_7308,N_3164,N_4448);
xnor U7309 (N_7309,N_2126,N_3675);
or U7310 (N_7310,N_2227,N_2846);
nand U7311 (N_7311,N_55,N_586);
and U7312 (N_7312,N_211,N_2331);
nor U7313 (N_7313,N_1608,N_10);
or U7314 (N_7314,N_853,N_2694);
xnor U7315 (N_7315,N_3661,N_2087);
or U7316 (N_7316,N_367,N_1960);
and U7317 (N_7317,N_1640,N_4900);
nor U7318 (N_7318,N_2526,N_3122);
or U7319 (N_7319,N_341,N_926);
or U7320 (N_7320,N_2049,N_3852);
nand U7321 (N_7321,N_809,N_2264);
and U7322 (N_7322,N_2680,N_1501);
nor U7323 (N_7323,N_2774,N_1594);
nand U7324 (N_7324,N_3755,N_1292);
nor U7325 (N_7325,N_2953,N_4823);
and U7326 (N_7326,N_296,N_4375);
nor U7327 (N_7327,N_1534,N_3334);
nand U7328 (N_7328,N_1649,N_2709);
or U7329 (N_7329,N_4377,N_1024);
xnor U7330 (N_7330,N_4442,N_3383);
or U7331 (N_7331,N_652,N_1493);
nand U7332 (N_7332,N_3431,N_4555);
or U7333 (N_7333,N_2386,N_4777);
and U7334 (N_7334,N_3032,N_1432);
nor U7335 (N_7335,N_1708,N_3670);
or U7336 (N_7336,N_3510,N_1001);
or U7337 (N_7337,N_4202,N_3736);
nand U7338 (N_7338,N_1106,N_1677);
nor U7339 (N_7339,N_4812,N_1837);
nand U7340 (N_7340,N_3187,N_4124);
xnor U7341 (N_7341,N_1475,N_1887);
or U7342 (N_7342,N_4420,N_4277);
and U7343 (N_7343,N_2178,N_976);
and U7344 (N_7344,N_3109,N_2649);
or U7345 (N_7345,N_2666,N_2151);
nor U7346 (N_7346,N_1017,N_2633);
and U7347 (N_7347,N_3020,N_4992);
nor U7348 (N_7348,N_3947,N_2007);
or U7349 (N_7349,N_2325,N_11);
xor U7350 (N_7350,N_470,N_4884);
or U7351 (N_7351,N_2477,N_3168);
or U7352 (N_7352,N_4674,N_790);
or U7353 (N_7353,N_32,N_3631);
or U7354 (N_7354,N_1067,N_3866);
or U7355 (N_7355,N_253,N_3749);
or U7356 (N_7356,N_2660,N_3266);
nand U7357 (N_7357,N_489,N_4593);
or U7358 (N_7358,N_3967,N_536);
and U7359 (N_7359,N_3022,N_2133);
or U7360 (N_7360,N_4246,N_1662);
and U7361 (N_7361,N_4166,N_3574);
and U7362 (N_7362,N_1850,N_1720);
or U7363 (N_7363,N_4346,N_3945);
nand U7364 (N_7364,N_1593,N_1994);
xor U7365 (N_7365,N_1543,N_2168);
nor U7366 (N_7366,N_486,N_4746);
and U7367 (N_7367,N_1353,N_1250);
nor U7368 (N_7368,N_161,N_3439);
nor U7369 (N_7369,N_388,N_3132);
nand U7370 (N_7370,N_4273,N_4348);
and U7371 (N_7371,N_4736,N_221);
nand U7372 (N_7372,N_3249,N_3066);
and U7373 (N_7373,N_4225,N_4358);
and U7374 (N_7374,N_282,N_3118);
nor U7375 (N_7375,N_2390,N_4050);
or U7376 (N_7376,N_2369,N_4439);
or U7377 (N_7377,N_3512,N_1628);
nand U7378 (N_7378,N_1198,N_1178);
nand U7379 (N_7379,N_3863,N_3042);
or U7380 (N_7380,N_616,N_2409);
or U7381 (N_7381,N_1201,N_1340);
nor U7382 (N_7382,N_867,N_1144);
nand U7383 (N_7383,N_1160,N_3214);
or U7384 (N_7384,N_240,N_2355);
nand U7385 (N_7385,N_4575,N_2098);
and U7386 (N_7386,N_4748,N_427);
and U7387 (N_7387,N_2663,N_848);
nand U7388 (N_7388,N_1412,N_4747);
and U7389 (N_7389,N_4792,N_849);
nor U7390 (N_7390,N_1212,N_500);
nor U7391 (N_7391,N_4175,N_3918);
and U7392 (N_7392,N_4304,N_1375);
and U7393 (N_7393,N_1028,N_3611);
xor U7394 (N_7394,N_1550,N_3369);
xnor U7395 (N_7395,N_2080,N_2239);
nor U7396 (N_7396,N_2023,N_4696);
nor U7397 (N_7397,N_3269,N_2904);
nand U7398 (N_7398,N_35,N_1520);
or U7399 (N_7399,N_3624,N_759);
and U7400 (N_7400,N_1782,N_2681);
nor U7401 (N_7401,N_2107,N_4665);
xor U7402 (N_7402,N_4893,N_3473);
and U7403 (N_7403,N_4329,N_4838);
nand U7404 (N_7404,N_3926,N_607);
nand U7405 (N_7405,N_2992,N_3878);
or U7406 (N_7406,N_3538,N_1748);
nand U7407 (N_7407,N_2971,N_3907);
or U7408 (N_7408,N_2899,N_1769);
xnor U7409 (N_7409,N_4470,N_453);
and U7410 (N_7410,N_3277,N_33);
or U7411 (N_7411,N_2347,N_1797);
xnor U7412 (N_7412,N_1964,N_3501);
nor U7413 (N_7413,N_249,N_598);
or U7414 (N_7414,N_1237,N_4832);
xnor U7415 (N_7415,N_4160,N_3010);
nand U7416 (N_7416,N_2553,N_1371);
and U7417 (N_7417,N_596,N_1101);
or U7418 (N_7418,N_4264,N_3994);
nor U7419 (N_7419,N_944,N_4321);
nand U7420 (N_7420,N_3933,N_2353);
or U7421 (N_7421,N_2370,N_3684);
and U7422 (N_7422,N_1792,N_2911);
and U7423 (N_7423,N_1414,N_2995);
nand U7424 (N_7424,N_3461,N_4300);
nor U7425 (N_7425,N_1418,N_2479);
nand U7426 (N_7426,N_4756,N_2445);
or U7427 (N_7427,N_4444,N_4194);
and U7428 (N_7428,N_748,N_731);
xor U7429 (N_7429,N_4170,N_1889);
nand U7430 (N_7430,N_738,N_3600);
xor U7431 (N_7431,N_3825,N_2485);
xnor U7432 (N_7432,N_2228,N_1822);
or U7433 (N_7433,N_4074,N_647);
nand U7434 (N_7434,N_3651,N_4343);
nor U7435 (N_7435,N_2692,N_2927);
or U7436 (N_7436,N_4029,N_2487);
nand U7437 (N_7437,N_3071,N_3682);
nand U7438 (N_7438,N_546,N_3990);
nand U7439 (N_7439,N_4627,N_162);
nand U7440 (N_7440,N_4433,N_1032);
nor U7441 (N_7441,N_2149,N_3043);
or U7442 (N_7442,N_401,N_3627);
nand U7443 (N_7443,N_4294,N_1780);
and U7444 (N_7444,N_1443,N_2290);
nand U7445 (N_7445,N_2565,N_1734);
or U7446 (N_7446,N_577,N_1808);
nor U7447 (N_7447,N_2789,N_955);
and U7448 (N_7448,N_3076,N_1730);
and U7449 (N_7449,N_1459,N_2505);
and U7450 (N_7450,N_3259,N_1168);
or U7451 (N_7451,N_3946,N_437);
or U7452 (N_7452,N_1194,N_2593);
or U7453 (N_7453,N_1368,N_1398);
or U7454 (N_7454,N_2537,N_3487);
xnor U7455 (N_7455,N_2129,N_2283);
nor U7456 (N_7456,N_1854,N_954);
or U7457 (N_7457,N_2246,N_434);
and U7458 (N_7458,N_1397,N_2020);
nor U7459 (N_7459,N_2015,N_2447);
or U7460 (N_7460,N_2336,N_1801);
nor U7461 (N_7461,N_3477,N_4189);
xor U7462 (N_7462,N_1058,N_1057);
xnor U7463 (N_7463,N_2588,N_982);
nand U7464 (N_7464,N_2268,N_518);
nand U7465 (N_7465,N_3328,N_279);
nand U7466 (N_7466,N_2735,N_508);
nor U7467 (N_7467,N_4281,N_754);
and U7468 (N_7468,N_1098,N_2101);
or U7469 (N_7469,N_4571,N_4762);
nand U7470 (N_7470,N_1612,N_1728);
nor U7471 (N_7471,N_309,N_3953);
nor U7472 (N_7472,N_2311,N_2685);
xnor U7473 (N_7473,N_1401,N_526);
and U7474 (N_7474,N_3469,N_4406);
nand U7475 (N_7475,N_2183,N_1498);
or U7476 (N_7476,N_2365,N_3111);
and U7477 (N_7477,N_4625,N_2730);
nand U7478 (N_7478,N_943,N_3716);
or U7479 (N_7479,N_3808,N_4307);
nor U7480 (N_7480,N_751,N_2925);
or U7481 (N_7481,N_4933,N_3712);
nand U7482 (N_7482,N_2572,N_3952);
nor U7483 (N_7483,N_4445,N_2211);
nand U7484 (N_7484,N_1499,N_3112);
nor U7485 (N_7485,N_4849,N_3840);
nor U7486 (N_7486,N_2955,N_439);
or U7487 (N_7487,N_3434,N_130);
xor U7488 (N_7488,N_2018,N_2491);
xnor U7489 (N_7489,N_1177,N_3059);
and U7490 (N_7490,N_4876,N_4092);
nand U7491 (N_7491,N_697,N_2017);
or U7492 (N_7492,N_4559,N_368);
and U7493 (N_7493,N_1585,N_2032);
or U7494 (N_7494,N_1396,N_4247);
nor U7495 (N_7495,N_4276,N_167);
and U7496 (N_7496,N_1918,N_4071);
xor U7497 (N_7497,N_2091,N_4450);
and U7498 (N_7498,N_2629,N_3427);
nor U7499 (N_7499,N_1814,N_2230);
and U7500 (N_7500,N_3651,N_3383);
nor U7501 (N_7501,N_3839,N_1190);
and U7502 (N_7502,N_1124,N_4354);
nor U7503 (N_7503,N_3110,N_2878);
and U7504 (N_7504,N_1201,N_4392);
nor U7505 (N_7505,N_4663,N_3024);
or U7506 (N_7506,N_2543,N_750);
or U7507 (N_7507,N_2616,N_3294);
nand U7508 (N_7508,N_1623,N_4145);
or U7509 (N_7509,N_404,N_3068);
or U7510 (N_7510,N_3653,N_1425);
and U7511 (N_7511,N_232,N_2541);
nor U7512 (N_7512,N_1171,N_3281);
or U7513 (N_7513,N_3669,N_349);
or U7514 (N_7514,N_1668,N_1671);
nand U7515 (N_7515,N_2184,N_3767);
or U7516 (N_7516,N_1801,N_904);
or U7517 (N_7517,N_3739,N_1976);
nand U7518 (N_7518,N_4653,N_2783);
nor U7519 (N_7519,N_2441,N_3736);
nand U7520 (N_7520,N_2792,N_4005);
and U7521 (N_7521,N_4864,N_856);
nand U7522 (N_7522,N_1759,N_1314);
nor U7523 (N_7523,N_2216,N_1094);
and U7524 (N_7524,N_669,N_3657);
or U7525 (N_7525,N_3541,N_2627);
nand U7526 (N_7526,N_2984,N_43);
and U7527 (N_7527,N_3791,N_891);
nand U7528 (N_7528,N_1695,N_2574);
nor U7529 (N_7529,N_549,N_176);
nor U7530 (N_7530,N_4035,N_3954);
or U7531 (N_7531,N_4000,N_2009);
nor U7532 (N_7532,N_620,N_4849);
or U7533 (N_7533,N_3701,N_2872);
or U7534 (N_7534,N_3678,N_4459);
and U7535 (N_7535,N_886,N_259);
nor U7536 (N_7536,N_4157,N_3558);
and U7537 (N_7537,N_2930,N_2833);
nand U7538 (N_7538,N_2426,N_3255);
nand U7539 (N_7539,N_4225,N_1936);
nand U7540 (N_7540,N_4399,N_4069);
xnor U7541 (N_7541,N_4427,N_1183);
or U7542 (N_7542,N_746,N_4571);
nand U7543 (N_7543,N_4491,N_4843);
nor U7544 (N_7544,N_3490,N_1330);
nand U7545 (N_7545,N_3622,N_2293);
nand U7546 (N_7546,N_4358,N_4135);
or U7547 (N_7547,N_770,N_1027);
and U7548 (N_7548,N_4903,N_2395);
nand U7549 (N_7549,N_4740,N_3176);
and U7550 (N_7550,N_4360,N_950);
nand U7551 (N_7551,N_3435,N_4634);
nor U7552 (N_7552,N_2056,N_1589);
nor U7553 (N_7553,N_2397,N_739);
or U7554 (N_7554,N_2238,N_2618);
nand U7555 (N_7555,N_1239,N_1161);
or U7556 (N_7556,N_3405,N_1163);
nand U7557 (N_7557,N_3774,N_199);
xnor U7558 (N_7558,N_4768,N_2570);
or U7559 (N_7559,N_1553,N_1380);
and U7560 (N_7560,N_2035,N_4409);
or U7561 (N_7561,N_4529,N_637);
nor U7562 (N_7562,N_2607,N_438);
and U7563 (N_7563,N_112,N_2276);
xnor U7564 (N_7564,N_2240,N_1503);
nand U7565 (N_7565,N_1906,N_2243);
nor U7566 (N_7566,N_1958,N_2520);
nand U7567 (N_7567,N_1997,N_2326);
or U7568 (N_7568,N_3458,N_4835);
and U7569 (N_7569,N_4632,N_3522);
and U7570 (N_7570,N_4373,N_776);
and U7571 (N_7571,N_3093,N_3774);
nor U7572 (N_7572,N_1884,N_81);
nand U7573 (N_7573,N_2187,N_4791);
and U7574 (N_7574,N_1309,N_1948);
nand U7575 (N_7575,N_1682,N_1224);
and U7576 (N_7576,N_3394,N_4866);
nor U7577 (N_7577,N_1781,N_1918);
or U7578 (N_7578,N_1754,N_663);
or U7579 (N_7579,N_3484,N_69);
nand U7580 (N_7580,N_590,N_3234);
or U7581 (N_7581,N_588,N_1550);
or U7582 (N_7582,N_2391,N_1622);
and U7583 (N_7583,N_2360,N_1428);
or U7584 (N_7584,N_1736,N_221);
and U7585 (N_7585,N_662,N_517);
and U7586 (N_7586,N_4063,N_2898);
nand U7587 (N_7587,N_3700,N_2150);
nand U7588 (N_7588,N_3010,N_2194);
nand U7589 (N_7589,N_2145,N_1855);
nand U7590 (N_7590,N_606,N_256);
nor U7591 (N_7591,N_3437,N_968);
and U7592 (N_7592,N_3992,N_3588);
or U7593 (N_7593,N_2032,N_1686);
or U7594 (N_7594,N_1780,N_2948);
nor U7595 (N_7595,N_4059,N_2594);
and U7596 (N_7596,N_1870,N_942);
and U7597 (N_7597,N_3755,N_2494);
and U7598 (N_7598,N_4965,N_4617);
and U7599 (N_7599,N_16,N_1712);
nand U7600 (N_7600,N_4253,N_3037);
and U7601 (N_7601,N_2106,N_2090);
or U7602 (N_7602,N_2692,N_4096);
nor U7603 (N_7603,N_2250,N_2773);
and U7604 (N_7604,N_4988,N_2478);
or U7605 (N_7605,N_983,N_4037);
and U7606 (N_7606,N_3270,N_3714);
and U7607 (N_7607,N_3623,N_2494);
and U7608 (N_7608,N_986,N_1348);
or U7609 (N_7609,N_3898,N_3664);
and U7610 (N_7610,N_1547,N_4435);
or U7611 (N_7611,N_1133,N_3048);
nor U7612 (N_7612,N_489,N_1935);
and U7613 (N_7613,N_2100,N_2443);
nand U7614 (N_7614,N_4936,N_2207);
nor U7615 (N_7615,N_2983,N_2931);
and U7616 (N_7616,N_3718,N_479);
and U7617 (N_7617,N_1909,N_1908);
nand U7618 (N_7618,N_3080,N_826);
xor U7619 (N_7619,N_2778,N_1933);
nor U7620 (N_7620,N_4213,N_4556);
nand U7621 (N_7621,N_1023,N_887);
and U7622 (N_7622,N_3751,N_2430);
nand U7623 (N_7623,N_3531,N_2104);
nand U7624 (N_7624,N_4214,N_3082);
xnor U7625 (N_7625,N_1892,N_3501);
or U7626 (N_7626,N_1277,N_2553);
nor U7627 (N_7627,N_4980,N_4105);
nand U7628 (N_7628,N_4657,N_1605);
nor U7629 (N_7629,N_3302,N_263);
and U7630 (N_7630,N_304,N_3371);
xnor U7631 (N_7631,N_3802,N_2801);
nor U7632 (N_7632,N_3789,N_3924);
nor U7633 (N_7633,N_4954,N_1289);
nor U7634 (N_7634,N_1898,N_3878);
xor U7635 (N_7635,N_3480,N_62);
and U7636 (N_7636,N_3065,N_928);
nand U7637 (N_7637,N_4691,N_1823);
xnor U7638 (N_7638,N_4678,N_5);
nor U7639 (N_7639,N_2402,N_2996);
and U7640 (N_7640,N_1478,N_2202);
or U7641 (N_7641,N_4841,N_620);
and U7642 (N_7642,N_4278,N_2070);
or U7643 (N_7643,N_4725,N_702);
nor U7644 (N_7644,N_2627,N_3840);
nor U7645 (N_7645,N_1744,N_729);
or U7646 (N_7646,N_662,N_3785);
or U7647 (N_7647,N_2453,N_4835);
nor U7648 (N_7648,N_2655,N_1331);
nand U7649 (N_7649,N_3984,N_3146);
xor U7650 (N_7650,N_982,N_1794);
nor U7651 (N_7651,N_4202,N_1224);
and U7652 (N_7652,N_1805,N_3200);
or U7653 (N_7653,N_3879,N_1159);
xor U7654 (N_7654,N_3268,N_2576);
and U7655 (N_7655,N_3465,N_1183);
nor U7656 (N_7656,N_3361,N_107);
or U7657 (N_7657,N_3883,N_3854);
or U7658 (N_7658,N_2518,N_3210);
and U7659 (N_7659,N_2152,N_592);
or U7660 (N_7660,N_4696,N_19);
nor U7661 (N_7661,N_565,N_4817);
and U7662 (N_7662,N_415,N_1279);
or U7663 (N_7663,N_640,N_1152);
nor U7664 (N_7664,N_1371,N_3042);
nor U7665 (N_7665,N_2457,N_4261);
nand U7666 (N_7666,N_1401,N_4159);
and U7667 (N_7667,N_2172,N_1858);
and U7668 (N_7668,N_4278,N_4574);
nor U7669 (N_7669,N_2691,N_2810);
or U7670 (N_7670,N_811,N_2315);
xor U7671 (N_7671,N_4808,N_3381);
nor U7672 (N_7672,N_443,N_1665);
and U7673 (N_7673,N_2755,N_4621);
or U7674 (N_7674,N_3087,N_179);
xor U7675 (N_7675,N_4505,N_3943);
or U7676 (N_7676,N_3291,N_1130);
nand U7677 (N_7677,N_3176,N_1868);
or U7678 (N_7678,N_1131,N_1851);
nand U7679 (N_7679,N_3914,N_2225);
and U7680 (N_7680,N_2786,N_793);
nor U7681 (N_7681,N_180,N_4046);
nand U7682 (N_7682,N_1783,N_4725);
and U7683 (N_7683,N_4493,N_1039);
nor U7684 (N_7684,N_621,N_2654);
nand U7685 (N_7685,N_441,N_254);
xnor U7686 (N_7686,N_449,N_2718);
xnor U7687 (N_7687,N_4926,N_549);
or U7688 (N_7688,N_944,N_1265);
and U7689 (N_7689,N_2579,N_3226);
nor U7690 (N_7690,N_556,N_1059);
or U7691 (N_7691,N_1413,N_161);
nand U7692 (N_7692,N_3857,N_4904);
nor U7693 (N_7693,N_2090,N_602);
nand U7694 (N_7694,N_2073,N_2289);
xnor U7695 (N_7695,N_2146,N_4072);
or U7696 (N_7696,N_234,N_4630);
and U7697 (N_7697,N_3920,N_2913);
xor U7698 (N_7698,N_625,N_2364);
nor U7699 (N_7699,N_3342,N_2366);
and U7700 (N_7700,N_914,N_4);
nor U7701 (N_7701,N_1515,N_400);
nand U7702 (N_7702,N_3769,N_3121);
nand U7703 (N_7703,N_4374,N_2913);
and U7704 (N_7704,N_2637,N_441);
or U7705 (N_7705,N_3998,N_2688);
or U7706 (N_7706,N_1055,N_2099);
nand U7707 (N_7707,N_1245,N_4052);
nand U7708 (N_7708,N_1538,N_3896);
or U7709 (N_7709,N_2412,N_1659);
or U7710 (N_7710,N_660,N_2968);
and U7711 (N_7711,N_3396,N_1360);
xor U7712 (N_7712,N_2138,N_712);
nand U7713 (N_7713,N_3503,N_4050);
nor U7714 (N_7714,N_3623,N_3483);
or U7715 (N_7715,N_2770,N_2218);
or U7716 (N_7716,N_4240,N_2555);
and U7717 (N_7717,N_3079,N_3318);
nand U7718 (N_7718,N_4552,N_3004);
nand U7719 (N_7719,N_4484,N_2461);
nand U7720 (N_7720,N_4599,N_3240);
or U7721 (N_7721,N_1167,N_3984);
nor U7722 (N_7722,N_4954,N_4162);
nand U7723 (N_7723,N_1751,N_1314);
nor U7724 (N_7724,N_3015,N_4028);
nor U7725 (N_7725,N_3823,N_1980);
nor U7726 (N_7726,N_706,N_4236);
or U7727 (N_7727,N_2027,N_4597);
and U7728 (N_7728,N_560,N_617);
nand U7729 (N_7729,N_4127,N_3886);
nand U7730 (N_7730,N_3698,N_2440);
xnor U7731 (N_7731,N_4772,N_3888);
nand U7732 (N_7732,N_109,N_3743);
or U7733 (N_7733,N_4000,N_4462);
xor U7734 (N_7734,N_4212,N_2948);
nor U7735 (N_7735,N_1536,N_3073);
and U7736 (N_7736,N_2536,N_2439);
and U7737 (N_7737,N_178,N_3408);
nand U7738 (N_7738,N_3707,N_2178);
xnor U7739 (N_7739,N_1077,N_2481);
xor U7740 (N_7740,N_4439,N_3096);
nand U7741 (N_7741,N_1721,N_2582);
and U7742 (N_7742,N_1397,N_4398);
xnor U7743 (N_7743,N_901,N_1639);
and U7744 (N_7744,N_3437,N_100);
and U7745 (N_7745,N_2359,N_4750);
nor U7746 (N_7746,N_3648,N_3359);
and U7747 (N_7747,N_691,N_1571);
nand U7748 (N_7748,N_3865,N_1403);
and U7749 (N_7749,N_3762,N_3994);
nor U7750 (N_7750,N_4906,N_3936);
or U7751 (N_7751,N_4639,N_588);
nor U7752 (N_7752,N_4227,N_2643);
or U7753 (N_7753,N_4768,N_4945);
nand U7754 (N_7754,N_4645,N_3947);
or U7755 (N_7755,N_546,N_1554);
nand U7756 (N_7756,N_4926,N_4009);
or U7757 (N_7757,N_1370,N_684);
and U7758 (N_7758,N_2468,N_1863);
or U7759 (N_7759,N_1324,N_2150);
nand U7760 (N_7760,N_3886,N_2822);
or U7761 (N_7761,N_2262,N_2486);
nor U7762 (N_7762,N_2000,N_21);
or U7763 (N_7763,N_4311,N_531);
and U7764 (N_7764,N_4227,N_3839);
xnor U7765 (N_7765,N_3472,N_1263);
or U7766 (N_7766,N_2734,N_4453);
nor U7767 (N_7767,N_3178,N_2658);
nand U7768 (N_7768,N_3554,N_503);
and U7769 (N_7769,N_261,N_4108);
or U7770 (N_7770,N_938,N_1848);
or U7771 (N_7771,N_1373,N_598);
xnor U7772 (N_7772,N_3493,N_1039);
nor U7773 (N_7773,N_1446,N_4025);
and U7774 (N_7774,N_197,N_4559);
and U7775 (N_7775,N_2908,N_3449);
nand U7776 (N_7776,N_962,N_3367);
or U7777 (N_7777,N_22,N_65);
or U7778 (N_7778,N_3347,N_2017);
nor U7779 (N_7779,N_1411,N_3338);
and U7780 (N_7780,N_327,N_2847);
or U7781 (N_7781,N_3548,N_2403);
and U7782 (N_7782,N_4617,N_3755);
and U7783 (N_7783,N_2861,N_1675);
and U7784 (N_7784,N_979,N_1201);
or U7785 (N_7785,N_4899,N_3645);
nand U7786 (N_7786,N_2679,N_791);
and U7787 (N_7787,N_72,N_4115);
nand U7788 (N_7788,N_3286,N_2020);
nor U7789 (N_7789,N_2493,N_1322);
nor U7790 (N_7790,N_3587,N_756);
nor U7791 (N_7791,N_4421,N_3117);
xnor U7792 (N_7792,N_2939,N_624);
or U7793 (N_7793,N_3789,N_3664);
nor U7794 (N_7794,N_345,N_4834);
and U7795 (N_7795,N_2842,N_555);
nand U7796 (N_7796,N_4863,N_3872);
and U7797 (N_7797,N_3100,N_727);
nor U7798 (N_7798,N_4938,N_3079);
or U7799 (N_7799,N_1095,N_4482);
xnor U7800 (N_7800,N_3371,N_239);
and U7801 (N_7801,N_2207,N_535);
nand U7802 (N_7802,N_3231,N_4963);
xnor U7803 (N_7803,N_33,N_1308);
nor U7804 (N_7804,N_1315,N_1120);
and U7805 (N_7805,N_4727,N_4722);
or U7806 (N_7806,N_3539,N_3248);
nand U7807 (N_7807,N_340,N_3384);
nand U7808 (N_7808,N_329,N_3671);
xor U7809 (N_7809,N_3127,N_3774);
nor U7810 (N_7810,N_845,N_387);
nand U7811 (N_7811,N_4953,N_1123);
and U7812 (N_7812,N_3226,N_4496);
nand U7813 (N_7813,N_988,N_1687);
nor U7814 (N_7814,N_44,N_1373);
nor U7815 (N_7815,N_4441,N_254);
xnor U7816 (N_7816,N_4925,N_1980);
nor U7817 (N_7817,N_1799,N_186);
nor U7818 (N_7818,N_877,N_1992);
and U7819 (N_7819,N_2716,N_1758);
nor U7820 (N_7820,N_1230,N_583);
or U7821 (N_7821,N_3887,N_3187);
or U7822 (N_7822,N_247,N_611);
and U7823 (N_7823,N_4645,N_3228);
or U7824 (N_7824,N_1389,N_3836);
xnor U7825 (N_7825,N_1265,N_4221);
or U7826 (N_7826,N_4367,N_2791);
nand U7827 (N_7827,N_3727,N_2722);
xnor U7828 (N_7828,N_3196,N_4003);
or U7829 (N_7829,N_4132,N_4795);
and U7830 (N_7830,N_1236,N_3028);
or U7831 (N_7831,N_3249,N_1645);
or U7832 (N_7832,N_1570,N_1341);
nor U7833 (N_7833,N_3045,N_1125);
and U7834 (N_7834,N_2096,N_4512);
nand U7835 (N_7835,N_2590,N_2501);
nand U7836 (N_7836,N_1811,N_1577);
nor U7837 (N_7837,N_2077,N_2804);
xnor U7838 (N_7838,N_3672,N_1609);
nand U7839 (N_7839,N_1364,N_440);
or U7840 (N_7840,N_3766,N_4121);
or U7841 (N_7841,N_4071,N_3575);
xor U7842 (N_7842,N_2319,N_1113);
or U7843 (N_7843,N_99,N_1144);
nand U7844 (N_7844,N_2981,N_117);
nor U7845 (N_7845,N_2918,N_4671);
nand U7846 (N_7846,N_4728,N_3610);
nor U7847 (N_7847,N_4065,N_1584);
nor U7848 (N_7848,N_4051,N_2130);
or U7849 (N_7849,N_2952,N_2015);
and U7850 (N_7850,N_245,N_4459);
nand U7851 (N_7851,N_1000,N_1732);
or U7852 (N_7852,N_590,N_3747);
nand U7853 (N_7853,N_3092,N_3695);
nor U7854 (N_7854,N_422,N_1576);
nand U7855 (N_7855,N_2488,N_1226);
or U7856 (N_7856,N_924,N_677);
nand U7857 (N_7857,N_4985,N_1894);
xor U7858 (N_7858,N_463,N_4453);
or U7859 (N_7859,N_3764,N_4411);
xor U7860 (N_7860,N_1890,N_805);
nor U7861 (N_7861,N_3543,N_2916);
nand U7862 (N_7862,N_2300,N_1347);
and U7863 (N_7863,N_3752,N_4069);
nor U7864 (N_7864,N_4112,N_4541);
xor U7865 (N_7865,N_4241,N_4745);
or U7866 (N_7866,N_4924,N_1945);
nand U7867 (N_7867,N_4156,N_1439);
nand U7868 (N_7868,N_3862,N_1748);
nand U7869 (N_7869,N_3779,N_4252);
nand U7870 (N_7870,N_4540,N_2395);
nor U7871 (N_7871,N_2041,N_1004);
and U7872 (N_7872,N_1747,N_3640);
nand U7873 (N_7873,N_2054,N_1996);
nor U7874 (N_7874,N_4789,N_4936);
nand U7875 (N_7875,N_103,N_2433);
or U7876 (N_7876,N_3283,N_259);
nand U7877 (N_7877,N_4354,N_3431);
and U7878 (N_7878,N_2905,N_668);
or U7879 (N_7879,N_4887,N_4386);
or U7880 (N_7880,N_4789,N_3446);
and U7881 (N_7881,N_1099,N_3980);
or U7882 (N_7882,N_2461,N_2335);
nand U7883 (N_7883,N_3207,N_4818);
or U7884 (N_7884,N_235,N_2753);
or U7885 (N_7885,N_3282,N_1401);
nor U7886 (N_7886,N_617,N_71);
nand U7887 (N_7887,N_3268,N_2825);
or U7888 (N_7888,N_2587,N_2387);
or U7889 (N_7889,N_1043,N_3139);
or U7890 (N_7890,N_3531,N_106);
nor U7891 (N_7891,N_744,N_4320);
nand U7892 (N_7892,N_3912,N_3061);
nor U7893 (N_7893,N_2462,N_2894);
or U7894 (N_7894,N_3223,N_1207);
or U7895 (N_7895,N_2902,N_4007);
nand U7896 (N_7896,N_1677,N_540);
nor U7897 (N_7897,N_1500,N_1335);
and U7898 (N_7898,N_1042,N_4502);
nor U7899 (N_7899,N_2234,N_2711);
nor U7900 (N_7900,N_2223,N_1421);
nand U7901 (N_7901,N_2936,N_2070);
xor U7902 (N_7902,N_3276,N_3248);
and U7903 (N_7903,N_924,N_4425);
nor U7904 (N_7904,N_3360,N_4911);
and U7905 (N_7905,N_437,N_3401);
and U7906 (N_7906,N_3586,N_885);
and U7907 (N_7907,N_4638,N_2774);
nor U7908 (N_7908,N_4765,N_3588);
nor U7909 (N_7909,N_596,N_1930);
nand U7910 (N_7910,N_3445,N_4149);
nand U7911 (N_7911,N_4905,N_2055);
and U7912 (N_7912,N_1173,N_3043);
nor U7913 (N_7913,N_2089,N_391);
nand U7914 (N_7914,N_367,N_2984);
and U7915 (N_7915,N_897,N_2954);
nor U7916 (N_7916,N_4076,N_2985);
or U7917 (N_7917,N_4132,N_1358);
nor U7918 (N_7918,N_4643,N_245);
or U7919 (N_7919,N_2673,N_2821);
or U7920 (N_7920,N_3164,N_201);
nor U7921 (N_7921,N_662,N_4822);
nand U7922 (N_7922,N_4010,N_4205);
or U7923 (N_7923,N_451,N_3773);
nor U7924 (N_7924,N_907,N_1909);
and U7925 (N_7925,N_3124,N_2537);
nand U7926 (N_7926,N_3149,N_2997);
nor U7927 (N_7927,N_4123,N_1005);
xnor U7928 (N_7928,N_2542,N_2298);
and U7929 (N_7929,N_494,N_2543);
and U7930 (N_7930,N_2771,N_2592);
and U7931 (N_7931,N_2813,N_2199);
and U7932 (N_7932,N_3648,N_856);
and U7933 (N_7933,N_2839,N_1050);
and U7934 (N_7934,N_4430,N_1626);
nor U7935 (N_7935,N_4090,N_630);
or U7936 (N_7936,N_488,N_2048);
and U7937 (N_7937,N_2871,N_905);
nand U7938 (N_7938,N_4111,N_952);
nand U7939 (N_7939,N_1428,N_4969);
xnor U7940 (N_7940,N_227,N_4611);
nor U7941 (N_7941,N_762,N_4242);
nand U7942 (N_7942,N_4483,N_33);
nor U7943 (N_7943,N_4969,N_1118);
and U7944 (N_7944,N_2209,N_543);
nor U7945 (N_7945,N_2592,N_3374);
or U7946 (N_7946,N_3756,N_4845);
xor U7947 (N_7947,N_1667,N_2658);
or U7948 (N_7948,N_947,N_1766);
nand U7949 (N_7949,N_2048,N_816);
or U7950 (N_7950,N_1751,N_3069);
nand U7951 (N_7951,N_4816,N_1176);
nand U7952 (N_7952,N_1449,N_488);
nor U7953 (N_7953,N_3192,N_3656);
or U7954 (N_7954,N_3946,N_3352);
nand U7955 (N_7955,N_1608,N_3606);
nor U7956 (N_7956,N_293,N_1506);
and U7957 (N_7957,N_3422,N_1887);
xnor U7958 (N_7958,N_12,N_4855);
and U7959 (N_7959,N_1167,N_2318);
nand U7960 (N_7960,N_816,N_1566);
nand U7961 (N_7961,N_3347,N_62);
nor U7962 (N_7962,N_4284,N_4893);
and U7963 (N_7963,N_1619,N_4594);
nor U7964 (N_7964,N_3983,N_1399);
nand U7965 (N_7965,N_1461,N_2555);
nand U7966 (N_7966,N_2322,N_2039);
or U7967 (N_7967,N_1296,N_2568);
and U7968 (N_7968,N_3237,N_2146);
or U7969 (N_7969,N_3814,N_4505);
nor U7970 (N_7970,N_4780,N_594);
nand U7971 (N_7971,N_4675,N_3925);
nand U7972 (N_7972,N_3844,N_1115);
nor U7973 (N_7973,N_3474,N_2933);
and U7974 (N_7974,N_941,N_1430);
nor U7975 (N_7975,N_2554,N_3456);
and U7976 (N_7976,N_508,N_4798);
or U7977 (N_7977,N_2741,N_1563);
nand U7978 (N_7978,N_2562,N_428);
and U7979 (N_7979,N_718,N_4663);
nand U7980 (N_7980,N_2097,N_4312);
and U7981 (N_7981,N_3549,N_1802);
nor U7982 (N_7982,N_2779,N_3585);
nand U7983 (N_7983,N_3087,N_4936);
or U7984 (N_7984,N_320,N_112);
and U7985 (N_7985,N_2475,N_481);
xnor U7986 (N_7986,N_372,N_1807);
nor U7987 (N_7987,N_4732,N_312);
xnor U7988 (N_7988,N_3988,N_590);
nor U7989 (N_7989,N_282,N_2472);
nand U7990 (N_7990,N_1948,N_423);
nor U7991 (N_7991,N_3398,N_1425);
and U7992 (N_7992,N_173,N_3870);
and U7993 (N_7993,N_2905,N_4611);
nor U7994 (N_7994,N_4667,N_3251);
and U7995 (N_7995,N_2672,N_1114);
or U7996 (N_7996,N_1426,N_3696);
nand U7997 (N_7997,N_2836,N_355);
nand U7998 (N_7998,N_3422,N_1353);
nor U7999 (N_7999,N_1735,N_172);
nand U8000 (N_8000,N_4387,N_3938);
nor U8001 (N_8001,N_909,N_39);
or U8002 (N_8002,N_1016,N_750);
and U8003 (N_8003,N_640,N_1292);
or U8004 (N_8004,N_2049,N_2084);
or U8005 (N_8005,N_1086,N_1664);
nor U8006 (N_8006,N_2901,N_1710);
xnor U8007 (N_8007,N_1416,N_3216);
nor U8008 (N_8008,N_2335,N_3489);
and U8009 (N_8009,N_1551,N_1603);
or U8010 (N_8010,N_3672,N_3938);
nand U8011 (N_8011,N_525,N_3912);
nor U8012 (N_8012,N_2026,N_1973);
and U8013 (N_8013,N_3336,N_1610);
and U8014 (N_8014,N_2791,N_4117);
or U8015 (N_8015,N_917,N_910);
nor U8016 (N_8016,N_2163,N_1477);
nor U8017 (N_8017,N_1464,N_252);
xor U8018 (N_8018,N_932,N_3945);
nor U8019 (N_8019,N_1058,N_176);
nor U8020 (N_8020,N_1532,N_2742);
and U8021 (N_8021,N_3902,N_1372);
xnor U8022 (N_8022,N_3337,N_66);
xnor U8023 (N_8023,N_4997,N_101);
or U8024 (N_8024,N_155,N_4075);
nand U8025 (N_8025,N_2825,N_3063);
nor U8026 (N_8026,N_4827,N_2514);
nor U8027 (N_8027,N_31,N_697);
or U8028 (N_8028,N_1045,N_3323);
nand U8029 (N_8029,N_4741,N_1296);
nor U8030 (N_8030,N_63,N_4161);
and U8031 (N_8031,N_2853,N_3031);
or U8032 (N_8032,N_3764,N_2459);
or U8033 (N_8033,N_2661,N_3750);
and U8034 (N_8034,N_1591,N_3115);
xnor U8035 (N_8035,N_2975,N_54);
xnor U8036 (N_8036,N_4377,N_3643);
and U8037 (N_8037,N_3550,N_4053);
or U8038 (N_8038,N_1381,N_3912);
nor U8039 (N_8039,N_292,N_2853);
nor U8040 (N_8040,N_2879,N_4351);
or U8041 (N_8041,N_3022,N_4551);
xnor U8042 (N_8042,N_1383,N_2576);
nor U8043 (N_8043,N_2008,N_1678);
nor U8044 (N_8044,N_3414,N_1751);
and U8045 (N_8045,N_2488,N_4843);
or U8046 (N_8046,N_1704,N_4037);
and U8047 (N_8047,N_1620,N_2855);
or U8048 (N_8048,N_1635,N_965);
nor U8049 (N_8049,N_2520,N_4951);
nor U8050 (N_8050,N_4141,N_4053);
and U8051 (N_8051,N_3977,N_691);
nand U8052 (N_8052,N_3224,N_840);
and U8053 (N_8053,N_206,N_4249);
nor U8054 (N_8054,N_4635,N_4791);
and U8055 (N_8055,N_880,N_3435);
or U8056 (N_8056,N_4950,N_3643);
or U8057 (N_8057,N_3882,N_1233);
and U8058 (N_8058,N_3827,N_2003);
nand U8059 (N_8059,N_2320,N_40);
or U8060 (N_8060,N_1358,N_1203);
and U8061 (N_8061,N_2948,N_1325);
nor U8062 (N_8062,N_2361,N_3695);
nor U8063 (N_8063,N_3964,N_1872);
or U8064 (N_8064,N_1726,N_4904);
or U8065 (N_8065,N_297,N_1609);
nor U8066 (N_8066,N_1074,N_2864);
nor U8067 (N_8067,N_4348,N_488);
and U8068 (N_8068,N_1531,N_155);
nand U8069 (N_8069,N_2746,N_3801);
or U8070 (N_8070,N_2237,N_4921);
nor U8071 (N_8071,N_2966,N_2361);
xor U8072 (N_8072,N_244,N_4345);
nor U8073 (N_8073,N_4045,N_1898);
and U8074 (N_8074,N_709,N_3970);
or U8075 (N_8075,N_230,N_3861);
or U8076 (N_8076,N_2401,N_3393);
or U8077 (N_8077,N_4554,N_365);
nor U8078 (N_8078,N_756,N_4553);
and U8079 (N_8079,N_3876,N_4588);
nor U8080 (N_8080,N_1800,N_2365);
nor U8081 (N_8081,N_1217,N_142);
nand U8082 (N_8082,N_4174,N_3810);
and U8083 (N_8083,N_2794,N_3820);
or U8084 (N_8084,N_1767,N_2065);
or U8085 (N_8085,N_4916,N_3321);
or U8086 (N_8086,N_3490,N_3227);
and U8087 (N_8087,N_103,N_2231);
or U8088 (N_8088,N_4868,N_3432);
nand U8089 (N_8089,N_3955,N_699);
or U8090 (N_8090,N_4933,N_799);
or U8091 (N_8091,N_3706,N_2171);
or U8092 (N_8092,N_445,N_460);
xor U8093 (N_8093,N_3107,N_2454);
or U8094 (N_8094,N_1018,N_4627);
and U8095 (N_8095,N_2153,N_3800);
or U8096 (N_8096,N_3582,N_670);
or U8097 (N_8097,N_97,N_4480);
nand U8098 (N_8098,N_1215,N_808);
or U8099 (N_8099,N_1908,N_124);
and U8100 (N_8100,N_4099,N_634);
nand U8101 (N_8101,N_3515,N_4268);
nor U8102 (N_8102,N_117,N_4563);
xnor U8103 (N_8103,N_3600,N_1745);
nand U8104 (N_8104,N_2283,N_3259);
nand U8105 (N_8105,N_3728,N_913);
xor U8106 (N_8106,N_1540,N_2255);
nor U8107 (N_8107,N_214,N_3663);
and U8108 (N_8108,N_1198,N_3986);
nand U8109 (N_8109,N_832,N_3555);
or U8110 (N_8110,N_3802,N_3753);
nor U8111 (N_8111,N_889,N_3876);
nor U8112 (N_8112,N_3142,N_1201);
and U8113 (N_8113,N_2195,N_3176);
nor U8114 (N_8114,N_4931,N_886);
nand U8115 (N_8115,N_4513,N_4117);
nand U8116 (N_8116,N_3635,N_1807);
xnor U8117 (N_8117,N_3660,N_2600);
nand U8118 (N_8118,N_266,N_2441);
xor U8119 (N_8119,N_1575,N_2726);
or U8120 (N_8120,N_1365,N_3409);
or U8121 (N_8121,N_505,N_4631);
or U8122 (N_8122,N_1759,N_2489);
nand U8123 (N_8123,N_1463,N_4003);
xnor U8124 (N_8124,N_1079,N_522);
nand U8125 (N_8125,N_2142,N_1178);
or U8126 (N_8126,N_4214,N_3731);
or U8127 (N_8127,N_4181,N_1385);
nor U8128 (N_8128,N_3334,N_4449);
or U8129 (N_8129,N_497,N_1685);
nand U8130 (N_8130,N_878,N_125);
or U8131 (N_8131,N_241,N_1157);
and U8132 (N_8132,N_4940,N_4471);
and U8133 (N_8133,N_4269,N_3746);
nor U8134 (N_8134,N_64,N_2757);
xnor U8135 (N_8135,N_3101,N_193);
and U8136 (N_8136,N_2334,N_4066);
xor U8137 (N_8137,N_13,N_2672);
xnor U8138 (N_8138,N_1917,N_3465);
and U8139 (N_8139,N_2222,N_59);
and U8140 (N_8140,N_4630,N_876);
xnor U8141 (N_8141,N_1976,N_954);
or U8142 (N_8142,N_1538,N_2611);
and U8143 (N_8143,N_2442,N_4315);
and U8144 (N_8144,N_1204,N_2435);
xnor U8145 (N_8145,N_2196,N_105);
nor U8146 (N_8146,N_361,N_3674);
and U8147 (N_8147,N_4679,N_2586);
nand U8148 (N_8148,N_1399,N_3754);
or U8149 (N_8149,N_4839,N_1893);
nand U8150 (N_8150,N_1536,N_3098);
nor U8151 (N_8151,N_1405,N_2693);
nand U8152 (N_8152,N_3686,N_1897);
xnor U8153 (N_8153,N_3169,N_743);
nand U8154 (N_8154,N_3256,N_3012);
nor U8155 (N_8155,N_2014,N_4424);
or U8156 (N_8156,N_2854,N_3150);
nor U8157 (N_8157,N_4200,N_3777);
nor U8158 (N_8158,N_568,N_2993);
xor U8159 (N_8159,N_801,N_2627);
nor U8160 (N_8160,N_185,N_2739);
and U8161 (N_8161,N_1721,N_4784);
or U8162 (N_8162,N_2904,N_639);
or U8163 (N_8163,N_2611,N_3076);
nor U8164 (N_8164,N_3763,N_2238);
or U8165 (N_8165,N_4396,N_213);
and U8166 (N_8166,N_3042,N_148);
nor U8167 (N_8167,N_1538,N_3077);
and U8168 (N_8168,N_4163,N_4298);
or U8169 (N_8169,N_4252,N_1948);
xnor U8170 (N_8170,N_4702,N_2202);
nor U8171 (N_8171,N_3836,N_1453);
xnor U8172 (N_8172,N_4272,N_1665);
and U8173 (N_8173,N_4551,N_2817);
or U8174 (N_8174,N_1282,N_1032);
or U8175 (N_8175,N_2218,N_4595);
nand U8176 (N_8176,N_3984,N_1412);
and U8177 (N_8177,N_1162,N_4056);
nand U8178 (N_8178,N_1289,N_1859);
nand U8179 (N_8179,N_3484,N_2038);
nand U8180 (N_8180,N_2748,N_2896);
or U8181 (N_8181,N_3163,N_1750);
xor U8182 (N_8182,N_1336,N_3195);
xor U8183 (N_8183,N_341,N_442);
nand U8184 (N_8184,N_2410,N_3646);
nor U8185 (N_8185,N_4638,N_2131);
nand U8186 (N_8186,N_617,N_1311);
nor U8187 (N_8187,N_3113,N_3775);
nor U8188 (N_8188,N_2209,N_3510);
nand U8189 (N_8189,N_1602,N_3102);
and U8190 (N_8190,N_3574,N_612);
or U8191 (N_8191,N_129,N_3254);
or U8192 (N_8192,N_3457,N_982);
and U8193 (N_8193,N_1005,N_2067);
nor U8194 (N_8194,N_434,N_717);
nand U8195 (N_8195,N_166,N_3266);
and U8196 (N_8196,N_206,N_4091);
nand U8197 (N_8197,N_3413,N_3838);
xnor U8198 (N_8198,N_2648,N_2422);
nand U8199 (N_8199,N_2153,N_3696);
nor U8200 (N_8200,N_3070,N_2164);
nor U8201 (N_8201,N_523,N_3489);
and U8202 (N_8202,N_335,N_4400);
or U8203 (N_8203,N_1887,N_792);
or U8204 (N_8204,N_1923,N_401);
and U8205 (N_8205,N_879,N_4645);
and U8206 (N_8206,N_774,N_2455);
nor U8207 (N_8207,N_927,N_1341);
nor U8208 (N_8208,N_2838,N_2572);
and U8209 (N_8209,N_4633,N_493);
nor U8210 (N_8210,N_1798,N_3696);
and U8211 (N_8211,N_1074,N_3384);
or U8212 (N_8212,N_2104,N_4016);
and U8213 (N_8213,N_4390,N_1957);
nor U8214 (N_8214,N_949,N_2122);
and U8215 (N_8215,N_4517,N_2586);
xor U8216 (N_8216,N_1125,N_3988);
nand U8217 (N_8217,N_2336,N_4843);
and U8218 (N_8218,N_1734,N_2071);
nor U8219 (N_8219,N_3294,N_4495);
nand U8220 (N_8220,N_4110,N_3639);
and U8221 (N_8221,N_1188,N_4436);
nand U8222 (N_8222,N_2101,N_2836);
xnor U8223 (N_8223,N_3189,N_2874);
nand U8224 (N_8224,N_3803,N_914);
or U8225 (N_8225,N_1281,N_3613);
or U8226 (N_8226,N_2041,N_1679);
or U8227 (N_8227,N_46,N_2126);
nand U8228 (N_8228,N_4888,N_4438);
or U8229 (N_8229,N_4965,N_4010);
or U8230 (N_8230,N_3408,N_513);
nor U8231 (N_8231,N_1216,N_967);
nor U8232 (N_8232,N_2117,N_2705);
nand U8233 (N_8233,N_1148,N_3937);
xor U8234 (N_8234,N_3489,N_1244);
nand U8235 (N_8235,N_529,N_1932);
and U8236 (N_8236,N_3456,N_1612);
and U8237 (N_8237,N_4599,N_143);
nor U8238 (N_8238,N_1765,N_2980);
nand U8239 (N_8239,N_2034,N_1358);
nor U8240 (N_8240,N_4903,N_717);
xor U8241 (N_8241,N_686,N_2071);
and U8242 (N_8242,N_3319,N_179);
nand U8243 (N_8243,N_2166,N_2840);
nand U8244 (N_8244,N_2869,N_2394);
nor U8245 (N_8245,N_4099,N_502);
nand U8246 (N_8246,N_4028,N_206);
and U8247 (N_8247,N_1143,N_1799);
nand U8248 (N_8248,N_1144,N_103);
nand U8249 (N_8249,N_2409,N_1803);
nand U8250 (N_8250,N_3047,N_775);
nand U8251 (N_8251,N_4502,N_4155);
and U8252 (N_8252,N_2268,N_3470);
and U8253 (N_8253,N_565,N_1802);
nand U8254 (N_8254,N_4856,N_1027);
nand U8255 (N_8255,N_4616,N_371);
and U8256 (N_8256,N_448,N_3390);
nand U8257 (N_8257,N_1552,N_1537);
and U8258 (N_8258,N_385,N_1661);
nand U8259 (N_8259,N_3038,N_1874);
and U8260 (N_8260,N_3301,N_2948);
and U8261 (N_8261,N_4475,N_832);
and U8262 (N_8262,N_4661,N_2986);
and U8263 (N_8263,N_2458,N_3872);
and U8264 (N_8264,N_512,N_924);
and U8265 (N_8265,N_1232,N_4313);
nor U8266 (N_8266,N_1978,N_2943);
or U8267 (N_8267,N_4987,N_1367);
nor U8268 (N_8268,N_170,N_3271);
xnor U8269 (N_8269,N_3091,N_2264);
nor U8270 (N_8270,N_4003,N_1573);
nor U8271 (N_8271,N_1332,N_3299);
or U8272 (N_8272,N_1771,N_3160);
or U8273 (N_8273,N_2413,N_3788);
nor U8274 (N_8274,N_2227,N_2092);
xnor U8275 (N_8275,N_4404,N_2013);
and U8276 (N_8276,N_2009,N_1354);
nand U8277 (N_8277,N_3003,N_711);
nor U8278 (N_8278,N_4896,N_3466);
nand U8279 (N_8279,N_2712,N_3295);
or U8280 (N_8280,N_2762,N_894);
xnor U8281 (N_8281,N_967,N_67);
and U8282 (N_8282,N_2953,N_4708);
nor U8283 (N_8283,N_2000,N_2938);
and U8284 (N_8284,N_3221,N_886);
xor U8285 (N_8285,N_4507,N_1124);
nor U8286 (N_8286,N_3142,N_229);
and U8287 (N_8287,N_3112,N_454);
or U8288 (N_8288,N_3671,N_3992);
and U8289 (N_8289,N_3844,N_3101);
or U8290 (N_8290,N_4818,N_3620);
and U8291 (N_8291,N_3917,N_3705);
and U8292 (N_8292,N_4542,N_246);
or U8293 (N_8293,N_3367,N_1345);
and U8294 (N_8294,N_2996,N_101);
xnor U8295 (N_8295,N_811,N_580);
or U8296 (N_8296,N_3521,N_971);
or U8297 (N_8297,N_3703,N_2013);
and U8298 (N_8298,N_4362,N_3941);
or U8299 (N_8299,N_3814,N_2299);
or U8300 (N_8300,N_4077,N_1263);
or U8301 (N_8301,N_2929,N_1614);
nand U8302 (N_8302,N_2173,N_828);
or U8303 (N_8303,N_62,N_164);
or U8304 (N_8304,N_2523,N_1112);
or U8305 (N_8305,N_3180,N_4004);
or U8306 (N_8306,N_84,N_798);
nand U8307 (N_8307,N_235,N_2601);
nand U8308 (N_8308,N_96,N_1613);
nand U8309 (N_8309,N_4302,N_4382);
nor U8310 (N_8310,N_4382,N_2490);
or U8311 (N_8311,N_2096,N_1963);
and U8312 (N_8312,N_3991,N_1537);
nor U8313 (N_8313,N_1078,N_690);
and U8314 (N_8314,N_1473,N_674);
nand U8315 (N_8315,N_2673,N_2886);
nand U8316 (N_8316,N_903,N_4649);
and U8317 (N_8317,N_1129,N_495);
nand U8318 (N_8318,N_2091,N_749);
xor U8319 (N_8319,N_4266,N_1507);
nor U8320 (N_8320,N_1676,N_3840);
or U8321 (N_8321,N_831,N_4211);
nor U8322 (N_8322,N_1460,N_2696);
and U8323 (N_8323,N_1216,N_322);
or U8324 (N_8324,N_589,N_2962);
and U8325 (N_8325,N_348,N_954);
nor U8326 (N_8326,N_4863,N_4995);
xor U8327 (N_8327,N_4006,N_4215);
or U8328 (N_8328,N_286,N_4999);
or U8329 (N_8329,N_2566,N_4893);
nor U8330 (N_8330,N_3070,N_4074);
xor U8331 (N_8331,N_1106,N_2344);
or U8332 (N_8332,N_2721,N_2469);
and U8333 (N_8333,N_4311,N_4666);
and U8334 (N_8334,N_3385,N_1034);
nand U8335 (N_8335,N_999,N_228);
xor U8336 (N_8336,N_1819,N_2616);
nor U8337 (N_8337,N_1902,N_4622);
nand U8338 (N_8338,N_3607,N_3313);
or U8339 (N_8339,N_2235,N_3855);
xor U8340 (N_8340,N_2111,N_3764);
nand U8341 (N_8341,N_2954,N_4963);
nand U8342 (N_8342,N_2819,N_3627);
nand U8343 (N_8343,N_1314,N_2077);
and U8344 (N_8344,N_4393,N_4200);
and U8345 (N_8345,N_3427,N_2759);
nand U8346 (N_8346,N_1364,N_4256);
and U8347 (N_8347,N_2517,N_1594);
nand U8348 (N_8348,N_3599,N_2642);
or U8349 (N_8349,N_2235,N_581);
or U8350 (N_8350,N_1036,N_363);
nand U8351 (N_8351,N_1612,N_4827);
nand U8352 (N_8352,N_2713,N_3335);
nor U8353 (N_8353,N_2619,N_2014);
xor U8354 (N_8354,N_2681,N_3328);
or U8355 (N_8355,N_3254,N_953);
nand U8356 (N_8356,N_2157,N_3585);
xor U8357 (N_8357,N_4005,N_4003);
nand U8358 (N_8358,N_1186,N_1760);
nand U8359 (N_8359,N_3175,N_680);
and U8360 (N_8360,N_409,N_1900);
and U8361 (N_8361,N_3705,N_3135);
nor U8362 (N_8362,N_3527,N_3152);
nor U8363 (N_8363,N_2870,N_2960);
or U8364 (N_8364,N_851,N_937);
nand U8365 (N_8365,N_4977,N_775);
xnor U8366 (N_8366,N_4846,N_3716);
or U8367 (N_8367,N_418,N_3648);
nand U8368 (N_8368,N_981,N_1157);
and U8369 (N_8369,N_1268,N_4183);
or U8370 (N_8370,N_157,N_2535);
nand U8371 (N_8371,N_832,N_3872);
nor U8372 (N_8372,N_2830,N_4030);
or U8373 (N_8373,N_120,N_1579);
or U8374 (N_8374,N_3993,N_4092);
or U8375 (N_8375,N_4370,N_2956);
nor U8376 (N_8376,N_2685,N_1988);
and U8377 (N_8377,N_630,N_2902);
or U8378 (N_8378,N_2167,N_1204);
xnor U8379 (N_8379,N_3326,N_3743);
nor U8380 (N_8380,N_1829,N_184);
or U8381 (N_8381,N_2140,N_3630);
nor U8382 (N_8382,N_1835,N_145);
nand U8383 (N_8383,N_562,N_314);
or U8384 (N_8384,N_87,N_2758);
or U8385 (N_8385,N_1951,N_643);
and U8386 (N_8386,N_788,N_122);
and U8387 (N_8387,N_4898,N_202);
nand U8388 (N_8388,N_1334,N_1182);
nand U8389 (N_8389,N_1152,N_4820);
nand U8390 (N_8390,N_4327,N_4656);
nand U8391 (N_8391,N_4047,N_3813);
or U8392 (N_8392,N_3838,N_3039);
nand U8393 (N_8393,N_1389,N_4904);
or U8394 (N_8394,N_1713,N_2234);
and U8395 (N_8395,N_2405,N_1524);
and U8396 (N_8396,N_4725,N_717);
or U8397 (N_8397,N_4048,N_398);
xor U8398 (N_8398,N_2815,N_3206);
or U8399 (N_8399,N_1790,N_2102);
and U8400 (N_8400,N_2155,N_3465);
nor U8401 (N_8401,N_4203,N_2025);
or U8402 (N_8402,N_4994,N_3102);
nand U8403 (N_8403,N_4054,N_727);
xnor U8404 (N_8404,N_3607,N_2283);
or U8405 (N_8405,N_3876,N_4379);
or U8406 (N_8406,N_2785,N_4073);
or U8407 (N_8407,N_3920,N_130);
nand U8408 (N_8408,N_2620,N_2338);
or U8409 (N_8409,N_781,N_4015);
nor U8410 (N_8410,N_4452,N_552);
or U8411 (N_8411,N_2861,N_3930);
nor U8412 (N_8412,N_4288,N_2120);
or U8413 (N_8413,N_128,N_4397);
nand U8414 (N_8414,N_3807,N_3991);
and U8415 (N_8415,N_3342,N_2813);
and U8416 (N_8416,N_4085,N_3406);
or U8417 (N_8417,N_763,N_3251);
xor U8418 (N_8418,N_3714,N_939);
and U8419 (N_8419,N_4056,N_3735);
or U8420 (N_8420,N_1528,N_1844);
and U8421 (N_8421,N_3974,N_533);
and U8422 (N_8422,N_358,N_2022);
and U8423 (N_8423,N_4593,N_1138);
nor U8424 (N_8424,N_945,N_1258);
nand U8425 (N_8425,N_4415,N_4722);
nand U8426 (N_8426,N_3721,N_989);
and U8427 (N_8427,N_3619,N_2562);
nand U8428 (N_8428,N_1743,N_501);
nand U8429 (N_8429,N_4594,N_3209);
nand U8430 (N_8430,N_2108,N_90);
nor U8431 (N_8431,N_829,N_885);
nor U8432 (N_8432,N_2605,N_2250);
nor U8433 (N_8433,N_114,N_489);
and U8434 (N_8434,N_1957,N_2600);
xor U8435 (N_8435,N_1690,N_1738);
and U8436 (N_8436,N_14,N_4887);
nand U8437 (N_8437,N_1124,N_235);
and U8438 (N_8438,N_3917,N_2795);
nand U8439 (N_8439,N_2137,N_4749);
and U8440 (N_8440,N_2524,N_2922);
or U8441 (N_8441,N_3026,N_4340);
and U8442 (N_8442,N_427,N_4684);
xor U8443 (N_8443,N_895,N_3367);
xor U8444 (N_8444,N_755,N_2890);
or U8445 (N_8445,N_2957,N_1518);
and U8446 (N_8446,N_3662,N_3532);
xnor U8447 (N_8447,N_2868,N_2749);
or U8448 (N_8448,N_3645,N_799);
nor U8449 (N_8449,N_4507,N_2512);
or U8450 (N_8450,N_1682,N_4819);
and U8451 (N_8451,N_1479,N_2298);
nand U8452 (N_8452,N_3663,N_2522);
nor U8453 (N_8453,N_1405,N_649);
and U8454 (N_8454,N_4350,N_416);
nor U8455 (N_8455,N_995,N_4569);
and U8456 (N_8456,N_203,N_4929);
nor U8457 (N_8457,N_4395,N_1227);
nand U8458 (N_8458,N_4305,N_4895);
and U8459 (N_8459,N_2663,N_2892);
xnor U8460 (N_8460,N_4617,N_4112);
xor U8461 (N_8461,N_2618,N_48);
nand U8462 (N_8462,N_4615,N_3514);
or U8463 (N_8463,N_753,N_787);
nor U8464 (N_8464,N_559,N_4970);
nand U8465 (N_8465,N_604,N_4060);
or U8466 (N_8466,N_286,N_882);
xnor U8467 (N_8467,N_3556,N_1598);
nor U8468 (N_8468,N_4797,N_2730);
and U8469 (N_8469,N_1492,N_282);
and U8470 (N_8470,N_2731,N_3573);
nand U8471 (N_8471,N_251,N_1643);
nor U8472 (N_8472,N_2411,N_3064);
or U8473 (N_8473,N_2047,N_4083);
or U8474 (N_8474,N_4456,N_189);
nand U8475 (N_8475,N_88,N_4245);
xor U8476 (N_8476,N_2708,N_4247);
and U8477 (N_8477,N_2631,N_878);
and U8478 (N_8478,N_3058,N_4786);
nand U8479 (N_8479,N_1300,N_514);
or U8480 (N_8480,N_2265,N_3736);
and U8481 (N_8481,N_169,N_1238);
or U8482 (N_8482,N_1172,N_2638);
and U8483 (N_8483,N_891,N_3647);
nor U8484 (N_8484,N_1113,N_2783);
and U8485 (N_8485,N_4809,N_3368);
nand U8486 (N_8486,N_1957,N_4752);
nand U8487 (N_8487,N_290,N_438);
nor U8488 (N_8488,N_4512,N_3810);
nor U8489 (N_8489,N_1551,N_1634);
xor U8490 (N_8490,N_2193,N_3730);
or U8491 (N_8491,N_2801,N_4030);
and U8492 (N_8492,N_2099,N_4292);
and U8493 (N_8493,N_4353,N_1977);
xor U8494 (N_8494,N_2004,N_1069);
nor U8495 (N_8495,N_2616,N_1703);
xnor U8496 (N_8496,N_2114,N_270);
xor U8497 (N_8497,N_2633,N_646);
nor U8498 (N_8498,N_3025,N_4306);
or U8499 (N_8499,N_2975,N_228);
nand U8500 (N_8500,N_1278,N_1564);
nand U8501 (N_8501,N_345,N_4079);
nor U8502 (N_8502,N_3013,N_2255);
nand U8503 (N_8503,N_3472,N_4455);
and U8504 (N_8504,N_2608,N_4270);
nor U8505 (N_8505,N_1624,N_1432);
and U8506 (N_8506,N_1506,N_1020);
or U8507 (N_8507,N_4811,N_1405);
and U8508 (N_8508,N_3046,N_1289);
nand U8509 (N_8509,N_2248,N_1551);
xor U8510 (N_8510,N_924,N_3419);
or U8511 (N_8511,N_737,N_425);
nand U8512 (N_8512,N_4696,N_3270);
nand U8513 (N_8513,N_1554,N_2088);
and U8514 (N_8514,N_1663,N_3575);
nor U8515 (N_8515,N_4291,N_1353);
or U8516 (N_8516,N_1938,N_2534);
nand U8517 (N_8517,N_4625,N_2277);
nor U8518 (N_8518,N_4319,N_4991);
xnor U8519 (N_8519,N_1533,N_1272);
or U8520 (N_8520,N_4572,N_3410);
or U8521 (N_8521,N_1721,N_1968);
nor U8522 (N_8522,N_519,N_4045);
and U8523 (N_8523,N_2700,N_1627);
or U8524 (N_8524,N_734,N_2935);
nand U8525 (N_8525,N_1861,N_4770);
nor U8526 (N_8526,N_4486,N_1253);
nor U8527 (N_8527,N_3651,N_3207);
xor U8528 (N_8528,N_243,N_899);
and U8529 (N_8529,N_2124,N_3262);
and U8530 (N_8530,N_1454,N_2066);
xnor U8531 (N_8531,N_2109,N_1008);
nand U8532 (N_8532,N_3524,N_3868);
nor U8533 (N_8533,N_3134,N_2135);
nand U8534 (N_8534,N_4188,N_3529);
nor U8535 (N_8535,N_947,N_195);
and U8536 (N_8536,N_4492,N_2627);
and U8537 (N_8537,N_93,N_3763);
nand U8538 (N_8538,N_999,N_2715);
nand U8539 (N_8539,N_673,N_2947);
or U8540 (N_8540,N_3645,N_800);
nand U8541 (N_8541,N_3967,N_4792);
xnor U8542 (N_8542,N_1477,N_3522);
or U8543 (N_8543,N_203,N_3272);
nor U8544 (N_8544,N_290,N_3131);
nor U8545 (N_8545,N_1537,N_3645);
nand U8546 (N_8546,N_3467,N_381);
and U8547 (N_8547,N_4323,N_4374);
and U8548 (N_8548,N_4053,N_1029);
nor U8549 (N_8549,N_2980,N_1792);
nor U8550 (N_8550,N_2167,N_4223);
xor U8551 (N_8551,N_4338,N_3074);
and U8552 (N_8552,N_1938,N_2250);
or U8553 (N_8553,N_4668,N_4006);
nor U8554 (N_8554,N_4296,N_4700);
and U8555 (N_8555,N_855,N_1565);
and U8556 (N_8556,N_2209,N_1072);
nor U8557 (N_8557,N_2865,N_2237);
nor U8558 (N_8558,N_4951,N_3180);
or U8559 (N_8559,N_2167,N_3915);
and U8560 (N_8560,N_2698,N_2847);
nor U8561 (N_8561,N_1647,N_1369);
nand U8562 (N_8562,N_2136,N_899);
xor U8563 (N_8563,N_1847,N_469);
nor U8564 (N_8564,N_1132,N_2769);
and U8565 (N_8565,N_2247,N_540);
or U8566 (N_8566,N_1981,N_2964);
or U8567 (N_8567,N_1806,N_1573);
and U8568 (N_8568,N_388,N_3232);
or U8569 (N_8569,N_1904,N_2863);
and U8570 (N_8570,N_2951,N_3526);
and U8571 (N_8571,N_161,N_3185);
or U8572 (N_8572,N_4206,N_2425);
nand U8573 (N_8573,N_3365,N_2908);
or U8574 (N_8574,N_4733,N_1947);
nor U8575 (N_8575,N_3730,N_562);
or U8576 (N_8576,N_1262,N_3238);
nor U8577 (N_8577,N_1042,N_2510);
or U8578 (N_8578,N_3349,N_1239);
or U8579 (N_8579,N_1934,N_966);
and U8580 (N_8580,N_2707,N_913);
nor U8581 (N_8581,N_2221,N_3247);
nand U8582 (N_8582,N_2074,N_1671);
and U8583 (N_8583,N_4014,N_3804);
or U8584 (N_8584,N_652,N_1821);
nand U8585 (N_8585,N_479,N_3541);
or U8586 (N_8586,N_1699,N_1530);
and U8587 (N_8587,N_4579,N_1406);
and U8588 (N_8588,N_4325,N_2035);
nor U8589 (N_8589,N_1818,N_4364);
nor U8590 (N_8590,N_3175,N_810);
xnor U8591 (N_8591,N_3570,N_3245);
or U8592 (N_8592,N_3239,N_2067);
and U8593 (N_8593,N_952,N_542);
nand U8594 (N_8594,N_4851,N_147);
or U8595 (N_8595,N_663,N_4547);
xnor U8596 (N_8596,N_223,N_886);
nand U8597 (N_8597,N_4775,N_2952);
or U8598 (N_8598,N_3844,N_1926);
nor U8599 (N_8599,N_1420,N_2913);
xor U8600 (N_8600,N_2863,N_3256);
or U8601 (N_8601,N_3380,N_2856);
nor U8602 (N_8602,N_4879,N_3900);
nand U8603 (N_8603,N_436,N_2018);
or U8604 (N_8604,N_687,N_3903);
nor U8605 (N_8605,N_4045,N_941);
or U8606 (N_8606,N_1988,N_4455);
and U8607 (N_8607,N_560,N_1437);
nor U8608 (N_8608,N_2464,N_2775);
nand U8609 (N_8609,N_4467,N_2629);
and U8610 (N_8610,N_709,N_3831);
and U8611 (N_8611,N_2785,N_2468);
nand U8612 (N_8612,N_1178,N_4830);
or U8613 (N_8613,N_2515,N_2130);
nand U8614 (N_8614,N_255,N_421);
and U8615 (N_8615,N_1401,N_3950);
nand U8616 (N_8616,N_3863,N_2161);
and U8617 (N_8617,N_2513,N_449);
or U8618 (N_8618,N_1213,N_2415);
nor U8619 (N_8619,N_3686,N_4638);
or U8620 (N_8620,N_567,N_1000);
and U8621 (N_8621,N_4354,N_4767);
or U8622 (N_8622,N_663,N_4721);
nand U8623 (N_8623,N_4125,N_2770);
nand U8624 (N_8624,N_3882,N_4313);
or U8625 (N_8625,N_1620,N_1928);
and U8626 (N_8626,N_3816,N_2989);
xnor U8627 (N_8627,N_1291,N_2801);
or U8628 (N_8628,N_2890,N_11);
nand U8629 (N_8629,N_4661,N_431);
nor U8630 (N_8630,N_4547,N_2004);
nor U8631 (N_8631,N_3047,N_1438);
nor U8632 (N_8632,N_231,N_856);
nand U8633 (N_8633,N_2916,N_3159);
nor U8634 (N_8634,N_1102,N_4248);
or U8635 (N_8635,N_4289,N_4525);
nor U8636 (N_8636,N_728,N_1996);
nor U8637 (N_8637,N_2475,N_1535);
and U8638 (N_8638,N_3005,N_4508);
and U8639 (N_8639,N_4534,N_3010);
nand U8640 (N_8640,N_618,N_3189);
nor U8641 (N_8641,N_2618,N_1670);
and U8642 (N_8642,N_1514,N_2682);
nor U8643 (N_8643,N_2520,N_36);
nand U8644 (N_8644,N_4686,N_2116);
or U8645 (N_8645,N_2670,N_2410);
nand U8646 (N_8646,N_1759,N_1682);
xnor U8647 (N_8647,N_3664,N_3816);
nor U8648 (N_8648,N_2852,N_1792);
or U8649 (N_8649,N_4377,N_2675);
or U8650 (N_8650,N_1601,N_4471);
or U8651 (N_8651,N_1524,N_105);
or U8652 (N_8652,N_3231,N_1679);
nand U8653 (N_8653,N_1199,N_4457);
xor U8654 (N_8654,N_893,N_1972);
nand U8655 (N_8655,N_243,N_2696);
nor U8656 (N_8656,N_2914,N_3148);
or U8657 (N_8657,N_4622,N_2945);
nand U8658 (N_8658,N_4983,N_3164);
or U8659 (N_8659,N_3926,N_3405);
xor U8660 (N_8660,N_315,N_3439);
or U8661 (N_8661,N_2960,N_4888);
and U8662 (N_8662,N_690,N_2286);
xnor U8663 (N_8663,N_4325,N_2637);
nand U8664 (N_8664,N_2416,N_4292);
nand U8665 (N_8665,N_4677,N_1186);
nor U8666 (N_8666,N_17,N_4984);
and U8667 (N_8667,N_151,N_3708);
nand U8668 (N_8668,N_3926,N_4317);
nand U8669 (N_8669,N_3882,N_3279);
nand U8670 (N_8670,N_454,N_4516);
and U8671 (N_8671,N_1476,N_1290);
and U8672 (N_8672,N_177,N_2968);
xnor U8673 (N_8673,N_4846,N_2631);
or U8674 (N_8674,N_1282,N_3642);
or U8675 (N_8675,N_3633,N_4977);
xor U8676 (N_8676,N_4547,N_3298);
or U8677 (N_8677,N_4189,N_3399);
xnor U8678 (N_8678,N_2377,N_1209);
or U8679 (N_8679,N_2202,N_640);
or U8680 (N_8680,N_2294,N_3867);
nor U8681 (N_8681,N_2604,N_3627);
xor U8682 (N_8682,N_4668,N_2267);
nor U8683 (N_8683,N_4135,N_1091);
nor U8684 (N_8684,N_4499,N_3007);
and U8685 (N_8685,N_4981,N_2023);
or U8686 (N_8686,N_932,N_3661);
nand U8687 (N_8687,N_1410,N_3633);
and U8688 (N_8688,N_2348,N_2300);
nor U8689 (N_8689,N_2613,N_3818);
xor U8690 (N_8690,N_3756,N_3373);
nand U8691 (N_8691,N_1461,N_66);
or U8692 (N_8692,N_4766,N_1999);
nand U8693 (N_8693,N_688,N_4268);
xor U8694 (N_8694,N_3158,N_742);
or U8695 (N_8695,N_683,N_4426);
nor U8696 (N_8696,N_3679,N_1441);
nor U8697 (N_8697,N_4445,N_3156);
xor U8698 (N_8698,N_4547,N_1616);
nor U8699 (N_8699,N_4895,N_1914);
and U8700 (N_8700,N_720,N_3891);
xor U8701 (N_8701,N_2278,N_2642);
nand U8702 (N_8702,N_2160,N_2106);
nor U8703 (N_8703,N_2118,N_4541);
nand U8704 (N_8704,N_3019,N_496);
nand U8705 (N_8705,N_1307,N_2676);
or U8706 (N_8706,N_3226,N_4427);
and U8707 (N_8707,N_2885,N_3794);
nor U8708 (N_8708,N_3999,N_4742);
nor U8709 (N_8709,N_2837,N_2851);
nor U8710 (N_8710,N_4306,N_4710);
nand U8711 (N_8711,N_1448,N_352);
xnor U8712 (N_8712,N_3893,N_652);
nand U8713 (N_8713,N_2592,N_4505);
and U8714 (N_8714,N_58,N_4170);
nor U8715 (N_8715,N_4805,N_4085);
xnor U8716 (N_8716,N_4787,N_4859);
nor U8717 (N_8717,N_3204,N_3686);
and U8718 (N_8718,N_244,N_3443);
and U8719 (N_8719,N_4204,N_4723);
and U8720 (N_8720,N_3510,N_3839);
nand U8721 (N_8721,N_3063,N_3067);
and U8722 (N_8722,N_4729,N_4877);
or U8723 (N_8723,N_925,N_61);
nor U8724 (N_8724,N_849,N_2300);
or U8725 (N_8725,N_2496,N_516);
nor U8726 (N_8726,N_2145,N_1335);
or U8727 (N_8727,N_1131,N_2729);
and U8728 (N_8728,N_3447,N_1698);
and U8729 (N_8729,N_2937,N_112);
and U8730 (N_8730,N_4700,N_4797);
and U8731 (N_8731,N_4936,N_32);
and U8732 (N_8732,N_4774,N_3021);
xnor U8733 (N_8733,N_884,N_4712);
and U8734 (N_8734,N_4462,N_2771);
nand U8735 (N_8735,N_4581,N_2642);
or U8736 (N_8736,N_4092,N_3914);
nor U8737 (N_8737,N_4483,N_2724);
nand U8738 (N_8738,N_2798,N_49);
or U8739 (N_8739,N_4270,N_2647);
nand U8740 (N_8740,N_514,N_1590);
or U8741 (N_8741,N_3074,N_4472);
xnor U8742 (N_8742,N_2209,N_4584);
and U8743 (N_8743,N_3257,N_3111);
nor U8744 (N_8744,N_3608,N_1701);
or U8745 (N_8745,N_4034,N_4258);
and U8746 (N_8746,N_152,N_4487);
and U8747 (N_8747,N_2842,N_1965);
nor U8748 (N_8748,N_2995,N_2090);
nor U8749 (N_8749,N_4858,N_4107);
nor U8750 (N_8750,N_1866,N_4387);
and U8751 (N_8751,N_1846,N_3764);
or U8752 (N_8752,N_510,N_3333);
and U8753 (N_8753,N_4169,N_3359);
nand U8754 (N_8754,N_3630,N_1034);
and U8755 (N_8755,N_3913,N_1837);
or U8756 (N_8756,N_2303,N_3532);
and U8757 (N_8757,N_2830,N_2893);
or U8758 (N_8758,N_4702,N_1759);
xor U8759 (N_8759,N_4835,N_3967);
nand U8760 (N_8760,N_1083,N_3161);
nand U8761 (N_8761,N_3388,N_2335);
nor U8762 (N_8762,N_3156,N_1931);
nand U8763 (N_8763,N_3938,N_2334);
and U8764 (N_8764,N_3064,N_99);
nand U8765 (N_8765,N_3256,N_3384);
nand U8766 (N_8766,N_4345,N_2210);
nand U8767 (N_8767,N_1354,N_2191);
and U8768 (N_8768,N_2830,N_3999);
and U8769 (N_8769,N_3296,N_38);
xnor U8770 (N_8770,N_580,N_421);
nor U8771 (N_8771,N_1973,N_3639);
xnor U8772 (N_8772,N_4362,N_373);
nor U8773 (N_8773,N_736,N_479);
nand U8774 (N_8774,N_721,N_1533);
nor U8775 (N_8775,N_2906,N_3536);
or U8776 (N_8776,N_192,N_1171);
and U8777 (N_8777,N_1176,N_1102);
nor U8778 (N_8778,N_2132,N_4315);
nand U8779 (N_8779,N_4313,N_1187);
and U8780 (N_8780,N_3277,N_2744);
or U8781 (N_8781,N_2078,N_4846);
or U8782 (N_8782,N_1064,N_3749);
nor U8783 (N_8783,N_878,N_3980);
and U8784 (N_8784,N_3957,N_2555);
and U8785 (N_8785,N_3401,N_4685);
or U8786 (N_8786,N_119,N_3497);
or U8787 (N_8787,N_3977,N_2486);
and U8788 (N_8788,N_4772,N_1684);
nand U8789 (N_8789,N_1,N_149);
or U8790 (N_8790,N_3942,N_2629);
nand U8791 (N_8791,N_1662,N_2498);
and U8792 (N_8792,N_2035,N_1716);
nor U8793 (N_8793,N_4040,N_602);
nor U8794 (N_8794,N_1035,N_4557);
nand U8795 (N_8795,N_1689,N_2670);
or U8796 (N_8796,N_3596,N_4005);
nor U8797 (N_8797,N_3525,N_2053);
nor U8798 (N_8798,N_141,N_3384);
and U8799 (N_8799,N_4846,N_1664);
or U8800 (N_8800,N_4010,N_3719);
nand U8801 (N_8801,N_488,N_4534);
nand U8802 (N_8802,N_2936,N_1575);
nor U8803 (N_8803,N_4319,N_2057);
and U8804 (N_8804,N_765,N_1302);
or U8805 (N_8805,N_2080,N_2594);
or U8806 (N_8806,N_4895,N_234);
or U8807 (N_8807,N_4267,N_1197);
and U8808 (N_8808,N_1585,N_2457);
and U8809 (N_8809,N_195,N_2151);
nor U8810 (N_8810,N_1234,N_2087);
and U8811 (N_8811,N_1111,N_1008);
nor U8812 (N_8812,N_2277,N_1238);
or U8813 (N_8813,N_4129,N_1447);
or U8814 (N_8814,N_2239,N_631);
nand U8815 (N_8815,N_2756,N_1911);
and U8816 (N_8816,N_1072,N_2339);
and U8817 (N_8817,N_1302,N_497);
and U8818 (N_8818,N_3760,N_2864);
nand U8819 (N_8819,N_4642,N_3560);
xor U8820 (N_8820,N_469,N_4805);
or U8821 (N_8821,N_3889,N_170);
and U8822 (N_8822,N_1661,N_3707);
nand U8823 (N_8823,N_643,N_4097);
nor U8824 (N_8824,N_69,N_2798);
and U8825 (N_8825,N_84,N_1414);
nor U8826 (N_8826,N_2661,N_2863);
and U8827 (N_8827,N_2128,N_836);
or U8828 (N_8828,N_2896,N_1310);
and U8829 (N_8829,N_3314,N_1025);
nor U8830 (N_8830,N_2251,N_3990);
nand U8831 (N_8831,N_1240,N_100);
nand U8832 (N_8832,N_3684,N_822);
or U8833 (N_8833,N_4235,N_3941);
nor U8834 (N_8834,N_1014,N_687);
xor U8835 (N_8835,N_2002,N_1443);
and U8836 (N_8836,N_4349,N_2849);
or U8837 (N_8837,N_116,N_3552);
and U8838 (N_8838,N_1941,N_1776);
nor U8839 (N_8839,N_515,N_4863);
or U8840 (N_8840,N_2262,N_1443);
nor U8841 (N_8841,N_1303,N_2421);
or U8842 (N_8842,N_4790,N_2378);
xor U8843 (N_8843,N_4696,N_4816);
nand U8844 (N_8844,N_126,N_4133);
and U8845 (N_8845,N_3864,N_3902);
nor U8846 (N_8846,N_778,N_1583);
or U8847 (N_8847,N_2649,N_1157);
xnor U8848 (N_8848,N_736,N_4167);
or U8849 (N_8849,N_2274,N_3064);
nand U8850 (N_8850,N_3234,N_3474);
nand U8851 (N_8851,N_3291,N_4220);
nor U8852 (N_8852,N_4968,N_4034);
nor U8853 (N_8853,N_1531,N_2527);
nand U8854 (N_8854,N_1523,N_2267);
nand U8855 (N_8855,N_2304,N_429);
nand U8856 (N_8856,N_257,N_2763);
nor U8857 (N_8857,N_1789,N_4748);
nor U8858 (N_8858,N_3842,N_4190);
or U8859 (N_8859,N_3759,N_4764);
nand U8860 (N_8860,N_1538,N_1532);
and U8861 (N_8861,N_638,N_276);
or U8862 (N_8862,N_2068,N_2332);
nor U8863 (N_8863,N_3685,N_2593);
xnor U8864 (N_8864,N_2645,N_2992);
nand U8865 (N_8865,N_591,N_4438);
nor U8866 (N_8866,N_1018,N_2903);
nand U8867 (N_8867,N_705,N_4697);
or U8868 (N_8868,N_2571,N_2501);
nor U8869 (N_8869,N_1879,N_316);
nand U8870 (N_8870,N_2207,N_4866);
or U8871 (N_8871,N_3095,N_415);
nor U8872 (N_8872,N_1668,N_4658);
and U8873 (N_8873,N_3426,N_3262);
nand U8874 (N_8874,N_1800,N_1839);
nor U8875 (N_8875,N_1381,N_4956);
nand U8876 (N_8876,N_3722,N_2706);
nor U8877 (N_8877,N_4415,N_1119);
nand U8878 (N_8878,N_4581,N_3814);
nor U8879 (N_8879,N_4915,N_4181);
xnor U8880 (N_8880,N_1531,N_4698);
xor U8881 (N_8881,N_4363,N_4948);
or U8882 (N_8882,N_2392,N_3643);
nand U8883 (N_8883,N_4586,N_2782);
nor U8884 (N_8884,N_1980,N_512);
xor U8885 (N_8885,N_4669,N_933);
or U8886 (N_8886,N_4662,N_507);
nand U8887 (N_8887,N_4457,N_1867);
and U8888 (N_8888,N_2898,N_4283);
and U8889 (N_8889,N_3189,N_2007);
nor U8890 (N_8890,N_499,N_1005);
or U8891 (N_8891,N_1795,N_4695);
nand U8892 (N_8892,N_4650,N_2183);
nand U8893 (N_8893,N_4633,N_3886);
nand U8894 (N_8894,N_2145,N_2938);
or U8895 (N_8895,N_3616,N_1693);
and U8896 (N_8896,N_1706,N_4641);
nor U8897 (N_8897,N_2339,N_671);
nor U8898 (N_8898,N_3023,N_3729);
and U8899 (N_8899,N_2496,N_3369);
xor U8900 (N_8900,N_1604,N_4292);
nor U8901 (N_8901,N_1845,N_3569);
and U8902 (N_8902,N_3653,N_2503);
or U8903 (N_8903,N_579,N_2771);
nand U8904 (N_8904,N_156,N_2278);
nor U8905 (N_8905,N_2831,N_3956);
or U8906 (N_8906,N_4215,N_1723);
or U8907 (N_8907,N_3270,N_1960);
xor U8908 (N_8908,N_1412,N_4899);
and U8909 (N_8909,N_4962,N_1007);
or U8910 (N_8910,N_2148,N_575);
xor U8911 (N_8911,N_2224,N_3554);
and U8912 (N_8912,N_4825,N_1057);
or U8913 (N_8913,N_2309,N_1352);
or U8914 (N_8914,N_2871,N_2405);
and U8915 (N_8915,N_1081,N_4707);
and U8916 (N_8916,N_3414,N_4280);
or U8917 (N_8917,N_404,N_4142);
nor U8918 (N_8918,N_4279,N_1948);
xnor U8919 (N_8919,N_4023,N_4239);
and U8920 (N_8920,N_88,N_1518);
and U8921 (N_8921,N_4278,N_3977);
nand U8922 (N_8922,N_3481,N_3857);
nor U8923 (N_8923,N_2947,N_2043);
and U8924 (N_8924,N_2165,N_1514);
nand U8925 (N_8925,N_4914,N_1322);
xor U8926 (N_8926,N_1901,N_2601);
and U8927 (N_8927,N_3892,N_989);
and U8928 (N_8928,N_2231,N_3933);
or U8929 (N_8929,N_1283,N_394);
nand U8930 (N_8930,N_1915,N_4402);
nand U8931 (N_8931,N_3310,N_315);
nor U8932 (N_8932,N_1705,N_1684);
and U8933 (N_8933,N_599,N_1488);
and U8934 (N_8934,N_181,N_2231);
or U8935 (N_8935,N_1094,N_3509);
nor U8936 (N_8936,N_1457,N_253);
nor U8937 (N_8937,N_864,N_4708);
nand U8938 (N_8938,N_1140,N_2340);
nand U8939 (N_8939,N_2400,N_562);
and U8940 (N_8940,N_3544,N_4167);
or U8941 (N_8941,N_2389,N_4771);
nor U8942 (N_8942,N_1320,N_3884);
and U8943 (N_8943,N_4703,N_4478);
xor U8944 (N_8944,N_1661,N_2410);
or U8945 (N_8945,N_2614,N_2195);
nand U8946 (N_8946,N_4946,N_1067);
xnor U8947 (N_8947,N_4332,N_4783);
or U8948 (N_8948,N_3761,N_3994);
and U8949 (N_8949,N_4433,N_83);
and U8950 (N_8950,N_3586,N_856);
nand U8951 (N_8951,N_4892,N_3305);
and U8952 (N_8952,N_3779,N_4755);
nand U8953 (N_8953,N_2665,N_2131);
xor U8954 (N_8954,N_4231,N_1064);
nand U8955 (N_8955,N_1338,N_281);
xor U8956 (N_8956,N_2416,N_4751);
and U8957 (N_8957,N_2106,N_1530);
and U8958 (N_8958,N_624,N_4286);
and U8959 (N_8959,N_1347,N_4576);
nand U8960 (N_8960,N_2358,N_2858);
and U8961 (N_8961,N_1196,N_2993);
nand U8962 (N_8962,N_2643,N_204);
nand U8963 (N_8963,N_2814,N_2446);
or U8964 (N_8964,N_987,N_233);
nor U8965 (N_8965,N_4365,N_1060);
or U8966 (N_8966,N_357,N_3175);
nor U8967 (N_8967,N_2140,N_772);
and U8968 (N_8968,N_4717,N_994);
nand U8969 (N_8969,N_4656,N_400);
xor U8970 (N_8970,N_3143,N_1637);
nor U8971 (N_8971,N_2958,N_516);
and U8972 (N_8972,N_1638,N_3106);
nor U8973 (N_8973,N_3593,N_4940);
nor U8974 (N_8974,N_4379,N_3936);
nor U8975 (N_8975,N_50,N_3596);
nand U8976 (N_8976,N_4214,N_2056);
or U8977 (N_8977,N_1901,N_1085);
nor U8978 (N_8978,N_2679,N_1274);
or U8979 (N_8979,N_1534,N_2247);
or U8980 (N_8980,N_3043,N_3716);
and U8981 (N_8981,N_2991,N_4727);
or U8982 (N_8982,N_206,N_324);
nor U8983 (N_8983,N_726,N_124);
and U8984 (N_8984,N_2413,N_995);
and U8985 (N_8985,N_2330,N_2042);
and U8986 (N_8986,N_548,N_213);
and U8987 (N_8987,N_4922,N_4851);
nor U8988 (N_8988,N_3090,N_1326);
and U8989 (N_8989,N_4340,N_1221);
or U8990 (N_8990,N_4263,N_2548);
xnor U8991 (N_8991,N_4316,N_2246);
or U8992 (N_8992,N_397,N_14);
nor U8993 (N_8993,N_2355,N_4190);
or U8994 (N_8994,N_1970,N_1049);
and U8995 (N_8995,N_1494,N_146);
nand U8996 (N_8996,N_1751,N_2582);
nand U8997 (N_8997,N_928,N_3569);
and U8998 (N_8998,N_4487,N_289);
or U8999 (N_8999,N_427,N_3172);
or U9000 (N_9000,N_55,N_869);
or U9001 (N_9001,N_3348,N_1628);
nor U9002 (N_9002,N_4686,N_1905);
or U9003 (N_9003,N_172,N_1503);
and U9004 (N_9004,N_1872,N_833);
nor U9005 (N_9005,N_1488,N_2419);
nor U9006 (N_9006,N_2711,N_2383);
nand U9007 (N_9007,N_1961,N_655);
or U9008 (N_9008,N_588,N_2598);
and U9009 (N_9009,N_4796,N_2146);
nor U9010 (N_9010,N_640,N_2240);
or U9011 (N_9011,N_758,N_312);
nor U9012 (N_9012,N_2231,N_592);
and U9013 (N_9013,N_3296,N_4317);
and U9014 (N_9014,N_2057,N_2720);
nor U9015 (N_9015,N_3527,N_1337);
nand U9016 (N_9016,N_1404,N_1750);
nor U9017 (N_9017,N_13,N_226);
or U9018 (N_9018,N_1706,N_3151);
and U9019 (N_9019,N_1475,N_2157);
nand U9020 (N_9020,N_4259,N_2323);
or U9021 (N_9021,N_3782,N_230);
and U9022 (N_9022,N_4270,N_635);
or U9023 (N_9023,N_3118,N_460);
nor U9024 (N_9024,N_658,N_127);
xnor U9025 (N_9025,N_4056,N_514);
or U9026 (N_9026,N_3424,N_4928);
nor U9027 (N_9027,N_3888,N_4394);
nand U9028 (N_9028,N_2600,N_2747);
and U9029 (N_9029,N_3621,N_3985);
or U9030 (N_9030,N_2513,N_4561);
xor U9031 (N_9031,N_895,N_1501);
and U9032 (N_9032,N_716,N_4493);
nand U9033 (N_9033,N_1663,N_33);
nor U9034 (N_9034,N_2150,N_4113);
nor U9035 (N_9035,N_981,N_1319);
and U9036 (N_9036,N_3537,N_2929);
and U9037 (N_9037,N_1278,N_823);
nor U9038 (N_9038,N_2347,N_4521);
or U9039 (N_9039,N_4887,N_1800);
nand U9040 (N_9040,N_3297,N_174);
or U9041 (N_9041,N_3620,N_1736);
and U9042 (N_9042,N_1626,N_1129);
and U9043 (N_9043,N_2955,N_2242);
nand U9044 (N_9044,N_2096,N_1923);
and U9045 (N_9045,N_2926,N_3186);
nor U9046 (N_9046,N_1716,N_387);
nand U9047 (N_9047,N_684,N_4464);
nor U9048 (N_9048,N_3479,N_1615);
or U9049 (N_9049,N_2500,N_751);
or U9050 (N_9050,N_4807,N_279);
xnor U9051 (N_9051,N_1453,N_3361);
xnor U9052 (N_9052,N_2656,N_4630);
or U9053 (N_9053,N_3572,N_4702);
xor U9054 (N_9054,N_2820,N_3416);
and U9055 (N_9055,N_3847,N_4750);
and U9056 (N_9056,N_2993,N_3295);
nor U9057 (N_9057,N_139,N_3281);
or U9058 (N_9058,N_1186,N_941);
and U9059 (N_9059,N_3003,N_1370);
nand U9060 (N_9060,N_1908,N_2650);
and U9061 (N_9061,N_900,N_242);
nand U9062 (N_9062,N_4407,N_3662);
or U9063 (N_9063,N_4419,N_1411);
nand U9064 (N_9064,N_4809,N_2914);
nand U9065 (N_9065,N_4145,N_3929);
or U9066 (N_9066,N_3070,N_2839);
nor U9067 (N_9067,N_2,N_767);
nor U9068 (N_9068,N_2079,N_3501);
nor U9069 (N_9069,N_1804,N_4363);
nand U9070 (N_9070,N_3915,N_976);
nor U9071 (N_9071,N_3385,N_534);
and U9072 (N_9072,N_4603,N_1002);
xor U9073 (N_9073,N_2188,N_724);
or U9074 (N_9074,N_1715,N_4917);
nand U9075 (N_9075,N_2925,N_4053);
nand U9076 (N_9076,N_4967,N_296);
nor U9077 (N_9077,N_3915,N_1413);
nand U9078 (N_9078,N_1964,N_4704);
nor U9079 (N_9079,N_4863,N_3449);
nor U9080 (N_9080,N_36,N_28);
nand U9081 (N_9081,N_4407,N_4561);
nand U9082 (N_9082,N_1950,N_2649);
and U9083 (N_9083,N_844,N_1341);
or U9084 (N_9084,N_3301,N_674);
xor U9085 (N_9085,N_2754,N_1342);
nor U9086 (N_9086,N_291,N_2558);
nand U9087 (N_9087,N_3072,N_1741);
xor U9088 (N_9088,N_4667,N_4697);
or U9089 (N_9089,N_2492,N_746);
nand U9090 (N_9090,N_4108,N_4922);
and U9091 (N_9091,N_4197,N_3739);
or U9092 (N_9092,N_4069,N_3219);
nand U9093 (N_9093,N_2663,N_2984);
nand U9094 (N_9094,N_4308,N_1360);
and U9095 (N_9095,N_3213,N_1749);
or U9096 (N_9096,N_2965,N_3305);
and U9097 (N_9097,N_1409,N_1741);
nor U9098 (N_9098,N_647,N_3809);
nor U9099 (N_9099,N_3449,N_4798);
nor U9100 (N_9100,N_1345,N_1957);
and U9101 (N_9101,N_2836,N_3045);
xnor U9102 (N_9102,N_2034,N_4116);
xnor U9103 (N_9103,N_1444,N_393);
nand U9104 (N_9104,N_3844,N_1278);
nor U9105 (N_9105,N_3159,N_1644);
and U9106 (N_9106,N_822,N_2745);
or U9107 (N_9107,N_2721,N_2163);
nor U9108 (N_9108,N_1125,N_4264);
nor U9109 (N_9109,N_2221,N_3888);
and U9110 (N_9110,N_4749,N_2795);
nand U9111 (N_9111,N_4871,N_3753);
or U9112 (N_9112,N_3204,N_4456);
and U9113 (N_9113,N_3735,N_3603);
nor U9114 (N_9114,N_2049,N_1384);
nor U9115 (N_9115,N_897,N_96);
nor U9116 (N_9116,N_4447,N_1426);
or U9117 (N_9117,N_2844,N_3132);
nor U9118 (N_9118,N_3341,N_3409);
and U9119 (N_9119,N_66,N_1274);
nor U9120 (N_9120,N_3474,N_560);
and U9121 (N_9121,N_4433,N_2514);
xor U9122 (N_9122,N_1657,N_2086);
nor U9123 (N_9123,N_57,N_1192);
xor U9124 (N_9124,N_4301,N_1551);
and U9125 (N_9125,N_251,N_131);
nand U9126 (N_9126,N_4491,N_2904);
and U9127 (N_9127,N_3479,N_1630);
nand U9128 (N_9128,N_172,N_1268);
or U9129 (N_9129,N_81,N_3429);
or U9130 (N_9130,N_4427,N_3408);
or U9131 (N_9131,N_1080,N_468);
or U9132 (N_9132,N_1258,N_4071);
xor U9133 (N_9133,N_304,N_1785);
nand U9134 (N_9134,N_1650,N_4619);
nand U9135 (N_9135,N_2655,N_2460);
nand U9136 (N_9136,N_3024,N_816);
nor U9137 (N_9137,N_1101,N_3883);
or U9138 (N_9138,N_2774,N_4174);
or U9139 (N_9139,N_567,N_3535);
nor U9140 (N_9140,N_2273,N_2448);
nand U9141 (N_9141,N_1626,N_1210);
nand U9142 (N_9142,N_4971,N_4943);
nor U9143 (N_9143,N_30,N_291);
or U9144 (N_9144,N_93,N_3205);
or U9145 (N_9145,N_3015,N_3794);
or U9146 (N_9146,N_1474,N_1848);
or U9147 (N_9147,N_491,N_1797);
and U9148 (N_9148,N_1037,N_2462);
nor U9149 (N_9149,N_2266,N_568);
xor U9150 (N_9150,N_4450,N_641);
nor U9151 (N_9151,N_4466,N_2433);
and U9152 (N_9152,N_473,N_3510);
or U9153 (N_9153,N_2235,N_742);
nand U9154 (N_9154,N_900,N_4968);
or U9155 (N_9155,N_1781,N_3162);
or U9156 (N_9156,N_3504,N_266);
nand U9157 (N_9157,N_4603,N_3800);
or U9158 (N_9158,N_602,N_3919);
nand U9159 (N_9159,N_1606,N_1877);
or U9160 (N_9160,N_1642,N_4024);
nand U9161 (N_9161,N_3052,N_3812);
xor U9162 (N_9162,N_1263,N_3221);
nand U9163 (N_9163,N_3476,N_2134);
or U9164 (N_9164,N_2051,N_1361);
nor U9165 (N_9165,N_4895,N_1230);
nand U9166 (N_9166,N_2530,N_2641);
or U9167 (N_9167,N_597,N_4872);
nand U9168 (N_9168,N_157,N_1453);
and U9169 (N_9169,N_4545,N_4150);
nor U9170 (N_9170,N_1493,N_1089);
nor U9171 (N_9171,N_3484,N_2286);
or U9172 (N_9172,N_2466,N_2775);
xor U9173 (N_9173,N_2786,N_1503);
nor U9174 (N_9174,N_2357,N_2529);
nor U9175 (N_9175,N_4406,N_2707);
xnor U9176 (N_9176,N_3583,N_2430);
xor U9177 (N_9177,N_1712,N_238);
or U9178 (N_9178,N_2720,N_628);
nand U9179 (N_9179,N_418,N_1224);
nor U9180 (N_9180,N_2760,N_2873);
or U9181 (N_9181,N_3046,N_4445);
nand U9182 (N_9182,N_3105,N_1133);
or U9183 (N_9183,N_4900,N_3114);
xor U9184 (N_9184,N_1353,N_2163);
or U9185 (N_9185,N_4731,N_3241);
nor U9186 (N_9186,N_3974,N_2675);
nor U9187 (N_9187,N_1301,N_360);
and U9188 (N_9188,N_421,N_4927);
and U9189 (N_9189,N_1854,N_1058);
and U9190 (N_9190,N_1508,N_4808);
or U9191 (N_9191,N_3231,N_1366);
and U9192 (N_9192,N_4059,N_81);
nor U9193 (N_9193,N_3520,N_999);
and U9194 (N_9194,N_1711,N_230);
nor U9195 (N_9195,N_2672,N_1989);
and U9196 (N_9196,N_2403,N_2209);
xor U9197 (N_9197,N_1840,N_2227);
or U9198 (N_9198,N_1728,N_836);
nor U9199 (N_9199,N_649,N_661);
and U9200 (N_9200,N_896,N_2221);
and U9201 (N_9201,N_4240,N_2128);
nor U9202 (N_9202,N_1710,N_935);
and U9203 (N_9203,N_2507,N_3915);
nor U9204 (N_9204,N_4572,N_4147);
xor U9205 (N_9205,N_2011,N_3547);
and U9206 (N_9206,N_891,N_2537);
or U9207 (N_9207,N_1074,N_3959);
and U9208 (N_9208,N_3234,N_2720);
nor U9209 (N_9209,N_773,N_2073);
nor U9210 (N_9210,N_2714,N_1038);
nor U9211 (N_9211,N_1842,N_75);
xnor U9212 (N_9212,N_796,N_2476);
nor U9213 (N_9213,N_3149,N_171);
or U9214 (N_9214,N_3734,N_2938);
nor U9215 (N_9215,N_3896,N_4312);
or U9216 (N_9216,N_148,N_2155);
nand U9217 (N_9217,N_3786,N_2519);
xnor U9218 (N_9218,N_1708,N_4852);
nand U9219 (N_9219,N_3608,N_2387);
nand U9220 (N_9220,N_4014,N_1086);
nand U9221 (N_9221,N_3144,N_3985);
xnor U9222 (N_9222,N_3399,N_4747);
and U9223 (N_9223,N_3309,N_3606);
or U9224 (N_9224,N_4176,N_2319);
nor U9225 (N_9225,N_2101,N_2939);
nor U9226 (N_9226,N_1111,N_823);
nand U9227 (N_9227,N_2817,N_3979);
and U9228 (N_9228,N_794,N_956);
nor U9229 (N_9229,N_38,N_1789);
and U9230 (N_9230,N_2016,N_565);
or U9231 (N_9231,N_4738,N_4945);
nand U9232 (N_9232,N_1815,N_1178);
or U9233 (N_9233,N_3346,N_4285);
nand U9234 (N_9234,N_294,N_1258);
and U9235 (N_9235,N_4525,N_3450);
or U9236 (N_9236,N_2285,N_658);
or U9237 (N_9237,N_690,N_1780);
nor U9238 (N_9238,N_4745,N_986);
or U9239 (N_9239,N_1095,N_1234);
and U9240 (N_9240,N_3893,N_2334);
nor U9241 (N_9241,N_3884,N_1180);
or U9242 (N_9242,N_1469,N_798);
nor U9243 (N_9243,N_4773,N_1347);
or U9244 (N_9244,N_1359,N_1684);
and U9245 (N_9245,N_4863,N_3765);
and U9246 (N_9246,N_1992,N_2981);
or U9247 (N_9247,N_3186,N_4235);
xor U9248 (N_9248,N_2652,N_4490);
or U9249 (N_9249,N_4059,N_921);
nand U9250 (N_9250,N_3169,N_2413);
nor U9251 (N_9251,N_3844,N_3890);
nand U9252 (N_9252,N_2275,N_4771);
and U9253 (N_9253,N_2518,N_3485);
nor U9254 (N_9254,N_1225,N_725);
or U9255 (N_9255,N_3187,N_2645);
nor U9256 (N_9256,N_2034,N_4827);
nor U9257 (N_9257,N_1820,N_1069);
nor U9258 (N_9258,N_3721,N_1441);
and U9259 (N_9259,N_421,N_1285);
nand U9260 (N_9260,N_4794,N_1244);
nand U9261 (N_9261,N_1168,N_4757);
nor U9262 (N_9262,N_4195,N_594);
or U9263 (N_9263,N_42,N_489);
xor U9264 (N_9264,N_861,N_645);
nor U9265 (N_9265,N_4978,N_403);
and U9266 (N_9266,N_3609,N_293);
and U9267 (N_9267,N_3289,N_4533);
nor U9268 (N_9268,N_3700,N_3199);
or U9269 (N_9269,N_1653,N_4204);
or U9270 (N_9270,N_4413,N_671);
nor U9271 (N_9271,N_964,N_4319);
nor U9272 (N_9272,N_564,N_1643);
nor U9273 (N_9273,N_369,N_384);
nor U9274 (N_9274,N_4425,N_4694);
nor U9275 (N_9275,N_3407,N_1691);
or U9276 (N_9276,N_2013,N_404);
nand U9277 (N_9277,N_3203,N_1674);
nor U9278 (N_9278,N_194,N_1854);
or U9279 (N_9279,N_4540,N_909);
nand U9280 (N_9280,N_4493,N_1005);
xor U9281 (N_9281,N_4059,N_115);
nand U9282 (N_9282,N_2702,N_819);
nand U9283 (N_9283,N_979,N_3442);
nand U9284 (N_9284,N_177,N_3071);
or U9285 (N_9285,N_1540,N_2327);
nand U9286 (N_9286,N_3371,N_2824);
nand U9287 (N_9287,N_268,N_1890);
and U9288 (N_9288,N_3403,N_3875);
nand U9289 (N_9289,N_1298,N_4100);
or U9290 (N_9290,N_2166,N_2367);
nor U9291 (N_9291,N_1230,N_2971);
and U9292 (N_9292,N_2729,N_3777);
nor U9293 (N_9293,N_4365,N_4650);
nor U9294 (N_9294,N_4820,N_1214);
nand U9295 (N_9295,N_4033,N_563);
xnor U9296 (N_9296,N_4400,N_3797);
nand U9297 (N_9297,N_1529,N_4126);
or U9298 (N_9298,N_4148,N_1197);
nand U9299 (N_9299,N_1392,N_2251);
nor U9300 (N_9300,N_1626,N_2649);
or U9301 (N_9301,N_3889,N_4253);
and U9302 (N_9302,N_1868,N_3075);
and U9303 (N_9303,N_3717,N_2416);
or U9304 (N_9304,N_3074,N_3418);
xnor U9305 (N_9305,N_1972,N_3113);
and U9306 (N_9306,N_2489,N_1664);
nor U9307 (N_9307,N_1114,N_4472);
nand U9308 (N_9308,N_159,N_828);
xnor U9309 (N_9309,N_1716,N_232);
xor U9310 (N_9310,N_1292,N_4424);
nand U9311 (N_9311,N_4376,N_1791);
and U9312 (N_9312,N_2449,N_401);
nor U9313 (N_9313,N_4699,N_4923);
nor U9314 (N_9314,N_4450,N_4700);
and U9315 (N_9315,N_3093,N_4368);
nand U9316 (N_9316,N_635,N_2952);
xnor U9317 (N_9317,N_3965,N_1004);
and U9318 (N_9318,N_23,N_3814);
and U9319 (N_9319,N_1368,N_4440);
nor U9320 (N_9320,N_2782,N_2832);
nand U9321 (N_9321,N_4459,N_127);
nor U9322 (N_9322,N_4577,N_4783);
and U9323 (N_9323,N_2161,N_1592);
and U9324 (N_9324,N_3577,N_1787);
nor U9325 (N_9325,N_1009,N_1144);
nor U9326 (N_9326,N_9,N_1741);
or U9327 (N_9327,N_2661,N_1555);
nor U9328 (N_9328,N_3217,N_603);
or U9329 (N_9329,N_2380,N_1760);
nor U9330 (N_9330,N_2156,N_309);
and U9331 (N_9331,N_1306,N_1780);
nor U9332 (N_9332,N_2278,N_1029);
nand U9333 (N_9333,N_1570,N_4983);
nor U9334 (N_9334,N_2327,N_764);
nand U9335 (N_9335,N_199,N_2807);
nor U9336 (N_9336,N_939,N_3734);
and U9337 (N_9337,N_4692,N_3167);
nand U9338 (N_9338,N_1003,N_4890);
and U9339 (N_9339,N_3947,N_2624);
and U9340 (N_9340,N_3538,N_1363);
nand U9341 (N_9341,N_992,N_41);
or U9342 (N_9342,N_2695,N_4662);
or U9343 (N_9343,N_4081,N_4539);
or U9344 (N_9344,N_2693,N_4644);
nand U9345 (N_9345,N_3632,N_2720);
nand U9346 (N_9346,N_3039,N_1651);
or U9347 (N_9347,N_4048,N_146);
or U9348 (N_9348,N_408,N_4233);
nand U9349 (N_9349,N_2070,N_1195);
xnor U9350 (N_9350,N_2070,N_2576);
nor U9351 (N_9351,N_3524,N_87);
nand U9352 (N_9352,N_2062,N_4100);
nor U9353 (N_9353,N_3300,N_38);
nor U9354 (N_9354,N_2132,N_1610);
and U9355 (N_9355,N_330,N_3866);
nand U9356 (N_9356,N_793,N_2866);
and U9357 (N_9357,N_3908,N_4061);
nand U9358 (N_9358,N_3502,N_4771);
xnor U9359 (N_9359,N_363,N_2048);
or U9360 (N_9360,N_2498,N_1803);
nand U9361 (N_9361,N_771,N_4102);
or U9362 (N_9362,N_3700,N_4443);
nand U9363 (N_9363,N_4477,N_115);
nand U9364 (N_9364,N_3084,N_1784);
and U9365 (N_9365,N_371,N_2196);
nand U9366 (N_9366,N_3873,N_2880);
and U9367 (N_9367,N_935,N_3370);
or U9368 (N_9368,N_1895,N_4980);
nor U9369 (N_9369,N_1125,N_4625);
nand U9370 (N_9370,N_75,N_2282);
xnor U9371 (N_9371,N_2340,N_900);
xor U9372 (N_9372,N_4942,N_820);
nand U9373 (N_9373,N_1542,N_4146);
nand U9374 (N_9374,N_1741,N_1838);
or U9375 (N_9375,N_2280,N_220);
and U9376 (N_9376,N_549,N_3479);
nand U9377 (N_9377,N_3072,N_4138);
and U9378 (N_9378,N_1666,N_1964);
and U9379 (N_9379,N_4093,N_3667);
xor U9380 (N_9380,N_684,N_1906);
nand U9381 (N_9381,N_3804,N_3405);
and U9382 (N_9382,N_3901,N_3042);
and U9383 (N_9383,N_4182,N_4029);
nand U9384 (N_9384,N_3364,N_1114);
nor U9385 (N_9385,N_1805,N_582);
xnor U9386 (N_9386,N_4539,N_2859);
nand U9387 (N_9387,N_121,N_4173);
or U9388 (N_9388,N_2775,N_774);
nand U9389 (N_9389,N_1955,N_2047);
or U9390 (N_9390,N_3227,N_2293);
or U9391 (N_9391,N_1926,N_2709);
nand U9392 (N_9392,N_788,N_3963);
or U9393 (N_9393,N_4210,N_3047);
nor U9394 (N_9394,N_675,N_3175);
or U9395 (N_9395,N_1469,N_3259);
nand U9396 (N_9396,N_4993,N_3693);
and U9397 (N_9397,N_289,N_177);
nand U9398 (N_9398,N_2395,N_2941);
nor U9399 (N_9399,N_1188,N_4666);
nor U9400 (N_9400,N_4561,N_802);
nand U9401 (N_9401,N_3939,N_4584);
or U9402 (N_9402,N_3839,N_639);
and U9403 (N_9403,N_1008,N_1689);
and U9404 (N_9404,N_210,N_1601);
nor U9405 (N_9405,N_847,N_2641);
and U9406 (N_9406,N_4715,N_2654);
or U9407 (N_9407,N_2640,N_3276);
xnor U9408 (N_9408,N_2436,N_992);
xnor U9409 (N_9409,N_1505,N_1022);
xnor U9410 (N_9410,N_1629,N_3204);
or U9411 (N_9411,N_3355,N_2337);
nor U9412 (N_9412,N_4099,N_4979);
nor U9413 (N_9413,N_4799,N_1280);
nand U9414 (N_9414,N_3929,N_381);
nor U9415 (N_9415,N_3468,N_1467);
nor U9416 (N_9416,N_2198,N_273);
nor U9417 (N_9417,N_616,N_4308);
and U9418 (N_9418,N_2496,N_2075);
or U9419 (N_9419,N_1173,N_155);
nand U9420 (N_9420,N_3890,N_3224);
or U9421 (N_9421,N_233,N_982);
or U9422 (N_9422,N_232,N_3025);
nor U9423 (N_9423,N_608,N_2936);
nor U9424 (N_9424,N_1933,N_4369);
and U9425 (N_9425,N_3905,N_459);
nor U9426 (N_9426,N_4271,N_1028);
or U9427 (N_9427,N_2353,N_531);
nand U9428 (N_9428,N_3680,N_3102);
or U9429 (N_9429,N_4945,N_860);
nor U9430 (N_9430,N_3796,N_1969);
and U9431 (N_9431,N_851,N_3726);
xor U9432 (N_9432,N_3335,N_1399);
and U9433 (N_9433,N_3510,N_4246);
nand U9434 (N_9434,N_2582,N_4681);
or U9435 (N_9435,N_4370,N_437);
nor U9436 (N_9436,N_2236,N_2764);
and U9437 (N_9437,N_1098,N_2948);
or U9438 (N_9438,N_3089,N_2758);
or U9439 (N_9439,N_2785,N_2335);
nor U9440 (N_9440,N_1474,N_4521);
nand U9441 (N_9441,N_3409,N_175);
and U9442 (N_9442,N_4601,N_3392);
nor U9443 (N_9443,N_4799,N_2664);
nor U9444 (N_9444,N_105,N_182);
xor U9445 (N_9445,N_196,N_2930);
or U9446 (N_9446,N_829,N_1985);
xnor U9447 (N_9447,N_927,N_3867);
nand U9448 (N_9448,N_631,N_156);
or U9449 (N_9449,N_2178,N_944);
nor U9450 (N_9450,N_4451,N_303);
and U9451 (N_9451,N_2926,N_4633);
and U9452 (N_9452,N_4484,N_3983);
nand U9453 (N_9453,N_4934,N_1036);
and U9454 (N_9454,N_3051,N_4790);
nand U9455 (N_9455,N_182,N_4694);
nor U9456 (N_9456,N_4715,N_704);
nor U9457 (N_9457,N_1504,N_809);
nand U9458 (N_9458,N_4282,N_2911);
nand U9459 (N_9459,N_4639,N_11);
and U9460 (N_9460,N_977,N_1025);
and U9461 (N_9461,N_1543,N_3003);
or U9462 (N_9462,N_190,N_2232);
xor U9463 (N_9463,N_3872,N_4250);
nor U9464 (N_9464,N_4781,N_3429);
nand U9465 (N_9465,N_1124,N_3697);
nor U9466 (N_9466,N_3053,N_2600);
and U9467 (N_9467,N_4621,N_309);
nand U9468 (N_9468,N_328,N_628);
or U9469 (N_9469,N_828,N_475);
and U9470 (N_9470,N_4989,N_4981);
nand U9471 (N_9471,N_3714,N_503);
nor U9472 (N_9472,N_489,N_2330);
or U9473 (N_9473,N_163,N_1017);
or U9474 (N_9474,N_877,N_3732);
nor U9475 (N_9475,N_567,N_239);
nand U9476 (N_9476,N_2503,N_1693);
nor U9477 (N_9477,N_1273,N_2526);
nor U9478 (N_9478,N_2164,N_393);
or U9479 (N_9479,N_4810,N_2385);
and U9480 (N_9480,N_711,N_875);
and U9481 (N_9481,N_3174,N_2193);
and U9482 (N_9482,N_1162,N_4181);
nand U9483 (N_9483,N_823,N_1697);
nor U9484 (N_9484,N_3795,N_2678);
nand U9485 (N_9485,N_3099,N_3444);
nand U9486 (N_9486,N_2595,N_4159);
xor U9487 (N_9487,N_1859,N_4365);
nand U9488 (N_9488,N_4983,N_3644);
and U9489 (N_9489,N_195,N_2341);
or U9490 (N_9490,N_491,N_2483);
nand U9491 (N_9491,N_2301,N_3278);
nand U9492 (N_9492,N_1063,N_1713);
and U9493 (N_9493,N_2624,N_3678);
xor U9494 (N_9494,N_2256,N_1991);
or U9495 (N_9495,N_546,N_3988);
nor U9496 (N_9496,N_1921,N_1206);
xor U9497 (N_9497,N_4018,N_237);
nor U9498 (N_9498,N_3896,N_718);
and U9499 (N_9499,N_2643,N_4401);
or U9500 (N_9500,N_4752,N_1935);
nand U9501 (N_9501,N_2727,N_3413);
nand U9502 (N_9502,N_261,N_3595);
nand U9503 (N_9503,N_395,N_4022);
nand U9504 (N_9504,N_1751,N_1598);
xor U9505 (N_9505,N_879,N_521);
nor U9506 (N_9506,N_2633,N_349);
and U9507 (N_9507,N_3329,N_2881);
and U9508 (N_9508,N_2876,N_4443);
nand U9509 (N_9509,N_3633,N_1911);
and U9510 (N_9510,N_3888,N_203);
nor U9511 (N_9511,N_2442,N_4611);
nor U9512 (N_9512,N_2866,N_931);
and U9513 (N_9513,N_3576,N_668);
nand U9514 (N_9514,N_1784,N_1589);
nor U9515 (N_9515,N_2733,N_1563);
xnor U9516 (N_9516,N_4828,N_116);
nand U9517 (N_9517,N_1121,N_3383);
and U9518 (N_9518,N_1960,N_3702);
xor U9519 (N_9519,N_2369,N_2836);
nand U9520 (N_9520,N_570,N_2289);
or U9521 (N_9521,N_4676,N_2755);
nand U9522 (N_9522,N_3465,N_3767);
nor U9523 (N_9523,N_4809,N_3699);
nor U9524 (N_9524,N_4952,N_2421);
nor U9525 (N_9525,N_1246,N_3010);
nor U9526 (N_9526,N_4325,N_4800);
nand U9527 (N_9527,N_1146,N_57);
nor U9528 (N_9528,N_3978,N_4996);
nor U9529 (N_9529,N_4478,N_1040);
nand U9530 (N_9530,N_1896,N_3827);
nand U9531 (N_9531,N_1856,N_1608);
nor U9532 (N_9532,N_4865,N_4748);
nand U9533 (N_9533,N_1787,N_2392);
nor U9534 (N_9534,N_2315,N_46);
nand U9535 (N_9535,N_3404,N_3259);
nor U9536 (N_9536,N_3902,N_669);
nand U9537 (N_9537,N_3,N_3436);
nor U9538 (N_9538,N_4849,N_422);
and U9539 (N_9539,N_2883,N_2446);
and U9540 (N_9540,N_2346,N_2416);
or U9541 (N_9541,N_2701,N_1622);
and U9542 (N_9542,N_1309,N_2535);
or U9543 (N_9543,N_66,N_3652);
nor U9544 (N_9544,N_752,N_2863);
nand U9545 (N_9545,N_791,N_507);
nand U9546 (N_9546,N_1181,N_2815);
nand U9547 (N_9547,N_4525,N_3130);
nand U9548 (N_9548,N_2733,N_4359);
nand U9549 (N_9549,N_2187,N_4206);
nor U9550 (N_9550,N_2670,N_1497);
nand U9551 (N_9551,N_3818,N_4152);
or U9552 (N_9552,N_3026,N_2339);
nor U9553 (N_9553,N_1320,N_1918);
and U9554 (N_9554,N_2426,N_451);
or U9555 (N_9555,N_4468,N_59);
or U9556 (N_9556,N_446,N_2605);
or U9557 (N_9557,N_3813,N_2543);
nor U9558 (N_9558,N_2436,N_545);
or U9559 (N_9559,N_944,N_308);
nor U9560 (N_9560,N_1256,N_905);
or U9561 (N_9561,N_955,N_4989);
nor U9562 (N_9562,N_759,N_4890);
and U9563 (N_9563,N_2400,N_3505);
nand U9564 (N_9564,N_4487,N_3795);
nand U9565 (N_9565,N_3364,N_1441);
nand U9566 (N_9566,N_2054,N_2021);
and U9567 (N_9567,N_669,N_4543);
and U9568 (N_9568,N_4530,N_4654);
and U9569 (N_9569,N_484,N_145);
nand U9570 (N_9570,N_343,N_4647);
xor U9571 (N_9571,N_1960,N_3414);
or U9572 (N_9572,N_3452,N_4889);
nand U9573 (N_9573,N_3552,N_337);
nand U9574 (N_9574,N_4848,N_1261);
xor U9575 (N_9575,N_2400,N_3463);
nand U9576 (N_9576,N_1870,N_259);
or U9577 (N_9577,N_4864,N_1178);
nand U9578 (N_9578,N_4654,N_135);
and U9579 (N_9579,N_2610,N_2589);
nor U9580 (N_9580,N_4723,N_349);
nor U9581 (N_9581,N_1205,N_127);
or U9582 (N_9582,N_68,N_3959);
xor U9583 (N_9583,N_4330,N_4628);
and U9584 (N_9584,N_2104,N_1994);
nand U9585 (N_9585,N_2853,N_433);
or U9586 (N_9586,N_2502,N_2932);
and U9587 (N_9587,N_4765,N_1464);
nor U9588 (N_9588,N_1830,N_3799);
nand U9589 (N_9589,N_3006,N_1070);
nor U9590 (N_9590,N_1199,N_3128);
or U9591 (N_9591,N_3584,N_1566);
nor U9592 (N_9592,N_1928,N_4429);
and U9593 (N_9593,N_3270,N_1860);
and U9594 (N_9594,N_939,N_3813);
or U9595 (N_9595,N_2220,N_1610);
or U9596 (N_9596,N_2567,N_3185);
or U9597 (N_9597,N_142,N_4055);
nand U9598 (N_9598,N_2826,N_2440);
nand U9599 (N_9599,N_4609,N_291);
nand U9600 (N_9600,N_1903,N_1857);
or U9601 (N_9601,N_470,N_676);
and U9602 (N_9602,N_1090,N_1258);
and U9603 (N_9603,N_2432,N_3449);
nand U9604 (N_9604,N_3253,N_2984);
and U9605 (N_9605,N_2476,N_4545);
nand U9606 (N_9606,N_422,N_1478);
nor U9607 (N_9607,N_3285,N_1237);
or U9608 (N_9608,N_4123,N_2033);
nor U9609 (N_9609,N_2740,N_3247);
and U9610 (N_9610,N_4380,N_1101);
and U9611 (N_9611,N_1284,N_658);
nor U9612 (N_9612,N_1710,N_1753);
nand U9613 (N_9613,N_2589,N_525);
nand U9614 (N_9614,N_290,N_4517);
nor U9615 (N_9615,N_4364,N_3535);
and U9616 (N_9616,N_4738,N_2640);
nor U9617 (N_9617,N_3564,N_678);
nand U9618 (N_9618,N_2186,N_3221);
nor U9619 (N_9619,N_1684,N_1961);
xnor U9620 (N_9620,N_4154,N_4955);
or U9621 (N_9621,N_3599,N_1799);
nor U9622 (N_9622,N_648,N_3609);
nor U9623 (N_9623,N_2887,N_1085);
and U9624 (N_9624,N_3093,N_974);
or U9625 (N_9625,N_4467,N_2479);
or U9626 (N_9626,N_155,N_1186);
nor U9627 (N_9627,N_3969,N_1912);
nand U9628 (N_9628,N_683,N_374);
and U9629 (N_9629,N_920,N_935);
or U9630 (N_9630,N_4494,N_4261);
or U9631 (N_9631,N_1116,N_4525);
nor U9632 (N_9632,N_3749,N_3259);
xnor U9633 (N_9633,N_1230,N_1962);
and U9634 (N_9634,N_4330,N_1422);
or U9635 (N_9635,N_1026,N_3136);
nor U9636 (N_9636,N_3459,N_451);
nor U9637 (N_9637,N_1227,N_3109);
or U9638 (N_9638,N_1379,N_1210);
and U9639 (N_9639,N_4801,N_1627);
xnor U9640 (N_9640,N_2484,N_252);
and U9641 (N_9641,N_4007,N_1948);
and U9642 (N_9642,N_4543,N_173);
nor U9643 (N_9643,N_2999,N_200);
or U9644 (N_9644,N_1658,N_2639);
xnor U9645 (N_9645,N_1837,N_1548);
or U9646 (N_9646,N_2364,N_1724);
nand U9647 (N_9647,N_144,N_3837);
nand U9648 (N_9648,N_3046,N_2680);
or U9649 (N_9649,N_3958,N_2784);
and U9650 (N_9650,N_1502,N_1071);
nor U9651 (N_9651,N_2197,N_4398);
and U9652 (N_9652,N_1925,N_1966);
or U9653 (N_9653,N_2178,N_281);
nand U9654 (N_9654,N_3071,N_175);
or U9655 (N_9655,N_275,N_361);
nor U9656 (N_9656,N_515,N_4866);
nand U9657 (N_9657,N_1644,N_4739);
xnor U9658 (N_9658,N_1209,N_181);
or U9659 (N_9659,N_2082,N_4744);
nor U9660 (N_9660,N_2799,N_3290);
or U9661 (N_9661,N_4442,N_2946);
or U9662 (N_9662,N_789,N_2337);
xor U9663 (N_9663,N_429,N_786);
xor U9664 (N_9664,N_2134,N_2636);
or U9665 (N_9665,N_2630,N_3926);
nand U9666 (N_9666,N_2170,N_3201);
nor U9667 (N_9667,N_2080,N_1455);
nand U9668 (N_9668,N_488,N_363);
and U9669 (N_9669,N_3412,N_695);
nand U9670 (N_9670,N_2594,N_1378);
nor U9671 (N_9671,N_2761,N_4250);
and U9672 (N_9672,N_1811,N_4893);
xnor U9673 (N_9673,N_4507,N_4729);
and U9674 (N_9674,N_1468,N_214);
and U9675 (N_9675,N_2544,N_3632);
nor U9676 (N_9676,N_639,N_4844);
and U9677 (N_9677,N_2116,N_4657);
and U9678 (N_9678,N_966,N_1249);
nor U9679 (N_9679,N_4450,N_3215);
nor U9680 (N_9680,N_2205,N_2630);
nand U9681 (N_9681,N_1400,N_441);
or U9682 (N_9682,N_2762,N_1117);
nand U9683 (N_9683,N_4147,N_2314);
nand U9684 (N_9684,N_2142,N_4083);
nand U9685 (N_9685,N_3641,N_925);
nand U9686 (N_9686,N_1289,N_627);
and U9687 (N_9687,N_2578,N_2726);
nand U9688 (N_9688,N_3693,N_2740);
and U9689 (N_9689,N_156,N_2671);
or U9690 (N_9690,N_1202,N_455);
nand U9691 (N_9691,N_3144,N_3645);
nor U9692 (N_9692,N_2407,N_499);
and U9693 (N_9693,N_4842,N_4920);
nor U9694 (N_9694,N_3986,N_3597);
and U9695 (N_9695,N_4732,N_4430);
xnor U9696 (N_9696,N_3392,N_3038);
xor U9697 (N_9697,N_2647,N_2);
nor U9698 (N_9698,N_3281,N_2575);
xor U9699 (N_9699,N_4274,N_3879);
xor U9700 (N_9700,N_2708,N_3390);
nor U9701 (N_9701,N_1155,N_35);
and U9702 (N_9702,N_3536,N_2088);
and U9703 (N_9703,N_3695,N_1350);
nor U9704 (N_9704,N_1744,N_1495);
or U9705 (N_9705,N_4142,N_836);
and U9706 (N_9706,N_2691,N_2466);
and U9707 (N_9707,N_2285,N_3882);
and U9708 (N_9708,N_792,N_3616);
nand U9709 (N_9709,N_3497,N_700);
nand U9710 (N_9710,N_4887,N_2822);
or U9711 (N_9711,N_447,N_1321);
and U9712 (N_9712,N_4663,N_379);
and U9713 (N_9713,N_4475,N_3268);
and U9714 (N_9714,N_1979,N_2373);
or U9715 (N_9715,N_1513,N_3165);
and U9716 (N_9716,N_3579,N_4150);
nor U9717 (N_9717,N_2501,N_4490);
nand U9718 (N_9718,N_3856,N_3866);
and U9719 (N_9719,N_3308,N_3924);
and U9720 (N_9720,N_407,N_4636);
or U9721 (N_9721,N_853,N_2491);
and U9722 (N_9722,N_525,N_3386);
nand U9723 (N_9723,N_928,N_4006);
nand U9724 (N_9724,N_4684,N_663);
and U9725 (N_9725,N_4420,N_2207);
or U9726 (N_9726,N_2744,N_4214);
or U9727 (N_9727,N_2328,N_3366);
and U9728 (N_9728,N_1590,N_4065);
nand U9729 (N_9729,N_1012,N_3732);
or U9730 (N_9730,N_3753,N_1152);
or U9731 (N_9731,N_81,N_21);
nand U9732 (N_9732,N_4513,N_285);
nor U9733 (N_9733,N_1589,N_4554);
and U9734 (N_9734,N_4611,N_1677);
nor U9735 (N_9735,N_3961,N_2143);
and U9736 (N_9736,N_2048,N_4765);
or U9737 (N_9737,N_3179,N_1962);
and U9738 (N_9738,N_3781,N_4957);
and U9739 (N_9739,N_4321,N_1883);
nor U9740 (N_9740,N_2070,N_2984);
or U9741 (N_9741,N_2752,N_2318);
nand U9742 (N_9742,N_4624,N_440);
nor U9743 (N_9743,N_1174,N_1385);
and U9744 (N_9744,N_1686,N_2802);
nand U9745 (N_9745,N_1423,N_4190);
or U9746 (N_9746,N_1691,N_721);
nor U9747 (N_9747,N_1108,N_3221);
and U9748 (N_9748,N_4535,N_796);
nor U9749 (N_9749,N_1356,N_3380);
nor U9750 (N_9750,N_1890,N_2894);
nand U9751 (N_9751,N_4323,N_4707);
nand U9752 (N_9752,N_2296,N_3437);
and U9753 (N_9753,N_2107,N_1965);
or U9754 (N_9754,N_4912,N_2039);
nand U9755 (N_9755,N_2827,N_2495);
nand U9756 (N_9756,N_1458,N_1520);
xor U9757 (N_9757,N_4988,N_3398);
nand U9758 (N_9758,N_1774,N_1519);
xor U9759 (N_9759,N_778,N_1455);
and U9760 (N_9760,N_2383,N_4128);
and U9761 (N_9761,N_3385,N_2119);
nand U9762 (N_9762,N_630,N_32);
or U9763 (N_9763,N_4562,N_950);
and U9764 (N_9764,N_1356,N_1688);
nor U9765 (N_9765,N_2151,N_961);
or U9766 (N_9766,N_1335,N_1617);
or U9767 (N_9767,N_3557,N_4746);
nor U9768 (N_9768,N_993,N_3996);
nand U9769 (N_9769,N_2941,N_1471);
or U9770 (N_9770,N_756,N_2804);
nand U9771 (N_9771,N_4337,N_728);
nor U9772 (N_9772,N_76,N_3357);
and U9773 (N_9773,N_4760,N_4470);
nand U9774 (N_9774,N_582,N_2594);
and U9775 (N_9775,N_1290,N_1700);
or U9776 (N_9776,N_1842,N_2809);
or U9777 (N_9777,N_3978,N_2160);
and U9778 (N_9778,N_4741,N_3993);
nand U9779 (N_9779,N_2458,N_4600);
or U9780 (N_9780,N_3676,N_1234);
and U9781 (N_9781,N_2156,N_3290);
or U9782 (N_9782,N_3653,N_2109);
nor U9783 (N_9783,N_3180,N_2948);
nor U9784 (N_9784,N_4524,N_4388);
or U9785 (N_9785,N_4597,N_636);
nand U9786 (N_9786,N_2448,N_738);
nand U9787 (N_9787,N_3087,N_4686);
or U9788 (N_9788,N_2379,N_624);
xnor U9789 (N_9789,N_3584,N_44);
or U9790 (N_9790,N_310,N_1775);
nor U9791 (N_9791,N_4191,N_3889);
xnor U9792 (N_9792,N_908,N_3595);
nand U9793 (N_9793,N_4346,N_3982);
nor U9794 (N_9794,N_990,N_1758);
xnor U9795 (N_9795,N_1627,N_512);
nand U9796 (N_9796,N_3720,N_3367);
nand U9797 (N_9797,N_1540,N_619);
nor U9798 (N_9798,N_3645,N_384);
and U9799 (N_9799,N_266,N_2356);
nor U9800 (N_9800,N_3686,N_3636);
nand U9801 (N_9801,N_2202,N_4938);
nand U9802 (N_9802,N_302,N_2911);
and U9803 (N_9803,N_1914,N_1287);
or U9804 (N_9804,N_4521,N_1158);
nor U9805 (N_9805,N_3235,N_1072);
xor U9806 (N_9806,N_4568,N_2266);
nor U9807 (N_9807,N_2996,N_3542);
xnor U9808 (N_9808,N_1753,N_4569);
nor U9809 (N_9809,N_3900,N_2643);
nor U9810 (N_9810,N_1359,N_3429);
or U9811 (N_9811,N_1129,N_2359);
nor U9812 (N_9812,N_1193,N_85);
nor U9813 (N_9813,N_872,N_4823);
nand U9814 (N_9814,N_2366,N_1987);
nor U9815 (N_9815,N_189,N_862);
nand U9816 (N_9816,N_1107,N_2555);
nand U9817 (N_9817,N_3865,N_1129);
nor U9818 (N_9818,N_1927,N_3012);
nor U9819 (N_9819,N_4493,N_14);
xnor U9820 (N_9820,N_1019,N_4718);
nor U9821 (N_9821,N_2225,N_677);
nand U9822 (N_9822,N_3496,N_455);
and U9823 (N_9823,N_441,N_2201);
nand U9824 (N_9824,N_316,N_3989);
and U9825 (N_9825,N_1233,N_2941);
nand U9826 (N_9826,N_840,N_4622);
or U9827 (N_9827,N_3520,N_669);
xor U9828 (N_9828,N_4614,N_2044);
and U9829 (N_9829,N_3632,N_3376);
nor U9830 (N_9830,N_1386,N_558);
nand U9831 (N_9831,N_4119,N_278);
nor U9832 (N_9832,N_4960,N_4692);
or U9833 (N_9833,N_3342,N_2043);
nand U9834 (N_9834,N_4726,N_1540);
and U9835 (N_9835,N_554,N_1084);
or U9836 (N_9836,N_2167,N_3959);
or U9837 (N_9837,N_656,N_2644);
nand U9838 (N_9838,N_2059,N_1535);
nor U9839 (N_9839,N_4010,N_3347);
xor U9840 (N_9840,N_719,N_4996);
and U9841 (N_9841,N_520,N_3234);
or U9842 (N_9842,N_3688,N_2853);
and U9843 (N_9843,N_2222,N_2870);
xnor U9844 (N_9844,N_3605,N_3341);
nand U9845 (N_9845,N_3416,N_2135);
and U9846 (N_9846,N_4765,N_2703);
or U9847 (N_9847,N_1635,N_3944);
xor U9848 (N_9848,N_741,N_4128);
and U9849 (N_9849,N_3724,N_2291);
nor U9850 (N_9850,N_818,N_2696);
or U9851 (N_9851,N_2977,N_2188);
nor U9852 (N_9852,N_3243,N_4176);
nand U9853 (N_9853,N_2728,N_362);
and U9854 (N_9854,N_890,N_4393);
or U9855 (N_9855,N_3240,N_2608);
nand U9856 (N_9856,N_3519,N_690);
and U9857 (N_9857,N_2652,N_3717);
nor U9858 (N_9858,N_4330,N_3411);
or U9859 (N_9859,N_3938,N_350);
nand U9860 (N_9860,N_4370,N_3199);
nor U9861 (N_9861,N_3148,N_5);
nand U9862 (N_9862,N_3423,N_2950);
nor U9863 (N_9863,N_1820,N_4521);
or U9864 (N_9864,N_2366,N_2212);
xor U9865 (N_9865,N_2666,N_950);
nor U9866 (N_9866,N_4909,N_4040);
and U9867 (N_9867,N_1257,N_632);
nand U9868 (N_9868,N_2683,N_4315);
and U9869 (N_9869,N_2686,N_2406);
nor U9870 (N_9870,N_4417,N_630);
nor U9871 (N_9871,N_1256,N_647);
or U9872 (N_9872,N_2435,N_3853);
and U9873 (N_9873,N_4913,N_3429);
or U9874 (N_9874,N_3914,N_2821);
and U9875 (N_9875,N_1192,N_1423);
and U9876 (N_9876,N_3564,N_3658);
nor U9877 (N_9877,N_4761,N_2089);
nand U9878 (N_9878,N_134,N_135);
and U9879 (N_9879,N_4174,N_2244);
and U9880 (N_9880,N_327,N_3309);
or U9881 (N_9881,N_1627,N_3522);
and U9882 (N_9882,N_2568,N_3548);
nor U9883 (N_9883,N_741,N_3838);
nand U9884 (N_9884,N_2611,N_2333);
or U9885 (N_9885,N_91,N_2683);
nand U9886 (N_9886,N_2008,N_4436);
nand U9887 (N_9887,N_724,N_1014);
xnor U9888 (N_9888,N_4786,N_2464);
or U9889 (N_9889,N_3804,N_4897);
nor U9890 (N_9890,N_1754,N_1808);
or U9891 (N_9891,N_1500,N_3877);
nor U9892 (N_9892,N_846,N_2137);
and U9893 (N_9893,N_2900,N_1266);
and U9894 (N_9894,N_2258,N_1745);
and U9895 (N_9895,N_542,N_318);
and U9896 (N_9896,N_2809,N_4271);
nand U9897 (N_9897,N_3481,N_4592);
and U9898 (N_9898,N_4478,N_3788);
nor U9899 (N_9899,N_1383,N_284);
nand U9900 (N_9900,N_3789,N_0);
nor U9901 (N_9901,N_1043,N_1790);
and U9902 (N_9902,N_4619,N_4450);
nor U9903 (N_9903,N_3923,N_1944);
nor U9904 (N_9904,N_3283,N_1550);
nand U9905 (N_9905,N_2457,N_2966);
nor U9906 (N_9906,N_4841,N_3524);
nand U9907 (N_9907,N_2173,N_1033);
xor U9908 (N_9908,N_4628,N_188);
nand U9909 (N_9909,N_3446,N_1710);
xnor U9910 (N_9910,N_538,N_2144);
and U9911 (N_9911,N_2468,N_1109);
or U9912 (N_9912,N_787,N_4434);
and U9913 (N_9913,N_3984,N_2020);
or U9914 (N_9914,N_2027,N_4729);
nor U9915 (N_9915,N_1433,N_3470);
and U9916 (N_9916,N_807,N_2798);
or U9917 (N_9917,N_2515,N_4264);
and U9918 (N_9918,N_547,N_681);
xnor U9919 (N_9919,N_4101,N_1101);
nand U9920 (N_9920,N_1901,N_1722);
and U9921 (N_9921,N_2280,N_3167);
nor U9922 (N_9922,N_2306,N_3468);
or U9923 (N_9923,N_1313,N_4530);
nor U9924 (N_9924,N_640,N_1821);
or U9925 (N_9925,N_1601,N_2804);
and U9926 (N_9926,N_2585,N_2793);
or U9927 (N_9927,N_4914,N_4033);
and U9928 (N_9928,N_378,N_1152);
and U9929 (N_9929,N_4426,N_4988);
nor U9930 (N_9930,N_4831,N_3225);
and U9931 (N_9931,N_3521,N_115);
or U9932 (N_9932,N_2023,N_605);
xor U9933 (N_9933,N_37,N_3391);
or U9934 (N_9934,N_337,N_3291);
and U9935 (N_9935,N_4122,N_1651);
xor U9936 (N_9936,N_4553,N_86);
or U9937 (N_9937,N_4080,N_4226);
or U9938 (N_9938,N_110,N_1564);
or U9939 (N_9939,N_3004,N_4540);
or U9940 (N_9940,N_3988,N_2273);
nor U9941 (N_9941,N_1566,N_4204);
nor U9942 (N_9942,N_3003,N_3940);
xnor U9943 (N_9943,N_3704,N_1452);
nor U9944 (N_9944,N_2109,N_4472);
nor U9945 (N_9945,N_4211,N_3642);
nand U9946 (N_9946,N_1852,N_2815);
or U9947 (N_9947,N_1094,N_1777);
or U9948 (N_9948,N_1068,N_1283);
nor U9949 (N_9949,N_1793,N_3073);
and U9950 (N_9950,N_893,N_293);
and U9951 (N_9951,N_617,N_3450);
nand U9952 (N_9952,N_2194,N_157);
or U9953 (N_9953,N_3007,N_3142);
or U9954 (N_9954,N_4918,N_276);
or U9955 (N_9955,N_2790,N_1192);
and U9956 (N_9956,N_1429,N_2505);
or U9957 (N_9957,N_1949,N_599);
nor U9958 (N_9958,N_2600,N_1966);
nand U9959 (N_9959,N_631,N_2681);
or U9960 (N_9960,N_40,N_4059);
nor U9961 (N_9961,N_2126,N_723);
and U9962 (N_9962,N_3425,N_1486);
and U9963 (N_9963,N_3535,N_3872);
nand U9964 (N_9964,N_4241,N_2304);
or U9965 (N_9965,N_802,N_3745);
or U9966 (N_9966,N_1307,N_461);
nand U9967 (N_9967,N_2852,N_4450);
nand U9968 (N_9968,N_4344,N_2825);
nand U9969 (N_9969,N_3093,N_2662);
nor U9970 (N_9970,N_3386,N_255);
nor U9971 (N_9971,N_2679,N_2797);
or U9972 (N_9972,N_587,N_2807);
nor U9973 (N_9973,N_2498,N_890);
nand U9974 (N_9974,N_933,N_441);
or U9975 (N_9975,N_4861,N_1801);
nor U9976 (N_9976,N_4890,N_2140);
nand U9977 (N_9977,N_4710,N_4783);
or U9978 (N_9978,N_4248,N_2756);
xnor U9979 (N_9979,N_2677,N_1567);
xnor U9980 (N_9980,N_228,N_3641);
or U9981 (N_9981,N_4688,N_3410);
nand U9982 (N_9982,N_3881,N_3415);
or U9983 (N_9983,N_2795,N_4500);
nor U9984 (N_9984,N_4009,N_5);
and U9985 (N_9985,N_3081,N_2515);
or U9986 (N_9986,N_764,N_3472);
nand U9987 (N_9987,N_3183,N_4088);
or U9988 (N_9988,N_766,N_2294);
and U9989 (N_9989,N_4409,N_94);
and U9990 (N_9990,N_447,N_2641);
or U9991 (N_9991,N_188,N_3292);
and U9992 (N_9992,N_243,N_607);
nor U9993 (N_9993,N_4236,N_876);
and U9994 (N_9994,N_4604,N_2881);
nand U9995 (N_9995,N_1626,N_2704);
and U9996 (N_9996,N_3741,N_2995);
and U9997 (N_9997,N_3553,N_2653);
and U9998 (N_9998,N_3201,N_3724);
nand U9999 (N_9999,N_1101,N_1013);
nand U10000 (N_10000,N_5751,N_8297);
nand U10001 (N_10001,N_6635,N_8996);
and U10002 (N_10002,N_8257,N_6638);
nand U10003 (N_10003,N_6913,N_6428);
and U10004 (N_10004,N_6055,N_9779);
nor U10005 (N_10005,N_9584,N_7971);
or U10006 (N_10006,N_8531,N_9268);
or U10007 (N_10007,N_9259,N_6271);
and U10008 (N_10008,N_6975,N_7657);
nor U10009 (N_10009,N_5274,N_9233);
nand U10010 (N_10010,N_9652,N_5135);
or U10011 (N_10011,N_7054,N_9859);
or U10012 (N_10012,N_6468,N_6640);
and U10013 (N_10013,N_9301,N_8960);
and U10014 (N_10014,N_6714,N_7361);
nor U10015 (N_10015,N_8057,N_5610);
and U10016 (N_10016,N_9730,N_9458);
or U10017 (N_10017,N_5053,N_9134);
nor U10018 (N_10018,N_9346,N_7681);
nand U10019 (N_10019,N_9451,N_5999);
nand U10020 (N_10020,N_9060,N_5073);
nand U10021 (N_10021,N_8185,N_9315);
nor U10022 (N_10022,N_9772,N_9917);
or U10023 (N_10023,N_7650,N_9115);
or U10024 (N_10024,N_7660,N_9701);
nand U10025 (N_10025,N_5229,N_9628);
or U10026 (N_10026,N_6399,N_8303);
and U10027 (N_10027,N_5338,N_9365);
nand U10028 (N_10028,N_5567,N_7093);
and U10029 (N_10029,N_5572,N_8671);
nand U10030 (N_10030,N_9207,N_5235);
nand U10031 (N_10031,N_9804,N_9444);
and U10032 (N_10032,N_9837,N_7744);
or U10033 (N_10033,N_7796,N_9025);
nand U10034 (N_10034,N_5617,N_9799);
and U10035 (N_10035,N_7258,N_6406);
nor U10036 (N_10036,N_5790,N_7221);
and U10037 (N_10037,N_5444,N_9145);
xnor U10038 (N_10038,N_6583,N_7570);
and U10039 (N_10039,N_8172,N_9682);
xor U10040 (N_10040,N_8628,N_7763);
or U10041 (N_10041,N_8553,N_9503);
and U10042 (N_10042,N_7242,N_6636);
nand U10043 (N_10043,N_6404,N_6286);
nor U10044 (N_10044,N_9291,N_8326);
nand U10045 (N_10045,N_6022,N_6459);
and U10046 (N_10046,N_9431,N_6996);
xnor U10047 (N_10047,N_5194,N_5876);
or U10048 (N_10048,N_5223,N_6113);
nor U10049 (N_10049,N_7263,N_7463);
xor U10050 (N_10050,N_7939,N_7889);
nand U10051 (N_10051,N_6655,N_7278);
xor U10052 (N_10052,N_8699,N_6709);
nor U10053 (N_10053,N_7789,N_5022);
nor U10054 (N_10054,N_5388,N_5689);
or U10055 (N_10055,N_8800,N_7643);
nor U10056 (N_10056,N_7536,N_6494);
nand U10057 (N_10057,N_6748,N_8871);
and U10058 (N_10058,N_7662,N_6212);
nand U10059 (N_10059,N_6499,N_6799);
and U10060 (N_10060,N_8486,N_5735);
and U10061 (N_10061,N_6992,N_7052);
xor U10062 (N_10062,N_8028,N_9508);
and U10063 (N_10063,N_7609,N_7251);
nor U10064 (N_10064,N_8092,N_8764);
nor U10065 (N_10065,N_5769,N_8272);
xor U10066 (N_10066,N_6859,N_7422);
nor U10067 (N_10067,N_6018,N_5827);
nor U10068 (N_10068,N_5351,N_5519);
nand U10069 (N_10069,N_9513,N_8851);
nor U10070 (N_10070,N_5347,N_7351);
xor U10071 (N_10071,N_8350,N_5342);
nand U10072 (N_10072,N_9852,N_7511);
and U10073 (N_10073,N_6521,N_7893);
and U10074 (N_10074,N_6962,N_9337);
and U10075 (N_10075,N_7821,N_5512);
xnor U10076 (N_10076,N_8448,N_9063);
nand U10077 (N_10077,N_9775,N_7767);
and U10078 (N_10078,N_9718,N_5178);
and U10079 (N_10079,N_5740,N_5973);
nand U10080 (N_10080,N_9320,N_5279);
and U10081 (N_10081,N_6054,N_6949);
nand U10082 (N_10082,N_5034,N_5111);
and U10083 (N_10083,N_8418,N_8314);
nand U10084 (N_10084,N_5280,N_9965);
and U10085 (N_10085,N_6519,N_5115);
and U10086 (N_10086,N_5492,N_6878);
or U10087 (N_10087,N_6110,N_7017);
nand U10088 (N_10088,N_5545,N_8682);
and U10089 (N_10089,N_9553,N_7369);
and U10090 (N_10090,N_8070,N_8374);
nand U10091 (N_10091,N_8902,N_6745);
xnor U10092 (N_10092,N_6316,N_9971);
and U10093 (N_10093,N_9987,N_7768);
nand U10094 (N_10094,N_6605,N_5171);
and U10095 (N_10095,N_5216,N_8889);
or U10096 (N_10096,N_5291,N_6674);
nand U10097 (N_10097,N_9362,N_8280);
nand U10098 (N_10098,N_5142,N_6074);
nand U10099 (N_10099,N_9177,N_7718);
nor U10100 (N_10100,N_9782,N_9057);
nor U10101 (N_10101,N_5190,N_5088);
nand U10102 (N_10102,N_7720,N_7780);
or U10103 (N_10103,N_6136,N_9831);
nor U10104 (N_10104,N_6001,N_9323);
nor U10105 (N_10105,N_8945,N_9022);
nand U10106 (N_10106,N_8860,N_8051);
nor U10107 (N_10107,N_5932,N_9281);
or U10108 (N_10108,N_6080,N_9729);
or U10109 (N_10109,N_6908,N_8719);
or U10110 (N_10110,N_9140,N_6780);
nor U10111 (N_10111,N_8982,N_9264);
and U10112 (N_10112,N_7310,N_5882);
xor U10113 (N_10113,N_7959,N_6105);
or U10114 (N_10114,N_5359,N_5843);
nor U10115 (N_10115,N_9146,N_8457);
and U10116 (N_10116,N_5303,N_8333);
or U10117 (N_10117,N_9582,N_9892);
and U10118 (N_10118,N_7595,N_9974);
xor U10119 (N_10119,N_9549,N_5813);
nor U10120 (N_10120,N_9119,N_9302);
xor U10121 (N_10121,N_5158,N_8766);
or U10122 (N_10122,N_7740,N_8406);
nor U10123 (N_10123,N_5426,N_8214);
and U10124 (N_10124,N_8342,N_9750);
or U10125 (N_10125,N_6269,N_6888);
and U10126 (N_10126,N_5160,N_6164);
nand U10127 (N_10127,N_7309,N_9869);
nand U10128 (N_10128,N_5753,N_7528);
and U10129 (N_10129,N_9690,N_6585);
nand U10130 (N_10130,N_9252,N_5316);
and U10131 (N_10131,N_7498,N_8515);
or U10132 (N_10132,N_5252,N_8141);
and U10133 (N_10133,N_8569,N_5634);
nor U10134 (N_10134,N_6569,N_7848);
xor U10135 (N_10135,N_7065,N_7013);
and U10136 (N_10136,N_6033,N_5383);
or U10137 (N_10137,N_8327,N_7653);
nand U10138 (N_10138,N_5715,N_8987);
nand U10139 (N_10139,N_7342,N_8991);
nor U10140 (N_10140,N_9941,N_9490);
and U10141 (N_10141,N_9762,N_5871);
nor U10142 (N_10142,N_7901,N_9183);
and U10143 (N_10143,N_9350,N_5148);
and U10144 (N_10144,N_6845,N_8095);
nand U10145 (N_10145,N_7073,N_9578);
or U10146 (N_10146,N_5393,N_5227);
nand U10147 (N_10147,N_5380,N_6787);
or U10148 (N_10148,N_7487,N_6615);
nand U10149 (N_10149,N_5570,N_5786);
and U10150 (N_10150,N_6012,N_8736);
nand U10151 (N_10151,N_9858,N_6296);
nand U10152 (N_10152,N_6434,N_6265);
or U10153 (N_10153,N_5513,N_8271);
or U10154 (N_10154,N_7910,N_9216);
or U10155 (N_10155,N_8485,N_8198);
nand U10156 (N_10156,N_8565,N_5612);
nor U10157 (N_10157,N_6790,N_6551);
xor U10158 (N_10158,N_7236,N_9904);
nand U10159 (N_10159,N_9052,N_9817);
and U10160 (N_10160,N_7717,N_5119);
nand U10161 (N_10161,N_9231,N_9910);
nor U10162 (N_10162,N_7521,N_5846);
or U10163 (N_10163,N_7230,N_8887);
or U10164 (N_10164,N_7173,N_6174);
nand U10165 (N_10165,N_8311,N_8029);
or U10166 (N_10166,N_9844,N_5661);
nand U10167 (N_10167,N_6960,N_8423);
xor U10168 (N_10168,N_6506,N_7390);
xor U10169 (N_10169,N_8165,N_5077);
nor U10170 (N_10170,N_7820,N_7854);
xnor U10171 (N_10171,N_5446,N_6972);
nand U10172 (N_10172,N_6612,N_7620);
and U10173 (N_10173,N_5348,N_7563);
or U10174 (N_10174,N_6108,N_9939);
and U10175 (N_10175,N_7007,N_8261);
or U10176 (N_10176,N_8601,N_5470);
and U10177 (N_10177,N_6393,N_6870);
or U10178 (N_10178,N_8263,N_5367);
or U10179 (N_10179,N_9055,N_9998);
nand U10180 (N_10180,N_7524,N_9012);
xnor U10181 (N_10181,N_5991,N_6232);
nand U10182 (N_10182,N_8109,N_8455);
nand U10183 (N_10183,N_6043,N_9442);
and U10184 (N_10184,N_6059,N_8684);
and U10185 (N_10185,N_7691,N_7082);
and U10186 (N_10186,N_5861,N_5020);
and U10187 (N_10187,N_7966,N_9737);
or U10188 (N_10188,N_6994,N_8433);
nand U10189 (N_10189,N_8016,N_6096);
or U10190 (N_10190,N_8420,N_8644);
and U10191 (N_10191,N_7492,N_8742);
xor U10192 (N_10192,N_8838,N_5533);
nor U10193 (N_10193,N_6090,N_8648);
and U10194 (N_10194,N_5980,N_7348);
or U10195 (N_10195,N_9861,N_6119);
xor U10196 (N_10196,N_9678,N_7738);
nor U10197 (N_10197,N_8778,N_8478);
and U10198 (N_10198,N_5177,N_6210);
or U10199 (N_10199,N_8909,N_8576);
and U10200 (N_10200,N_6221,N_7191);
or U10201 (N_10201,N_8679,N_9615);
nand U10202 (N_10202,N_5797,N_5820);
nor U10203 (N_10203,N_8662,N_7765);
nor U10204 (N_10204,N_9573,N_8425);
nand U10205 (N_10205,N_8290,N_5441);
nor U10206 (N_10206,N_9656,N_9129);
and U10207 (N_10207,N_6207,N_5702);
or U10208 (N_10208,N_8654,N_9091);
and U10209 (N_10209,N_8949,N_8842);
nand U10210 (N_10210,N_6518,N_9441);
or U10211 (N_10211,N_8950,N_7379);
and U10212 (N_10212,N_9843,N_9499);
or U10213 (N_10213,N_5575,N_6394);
nand U10214 (N_10214,N_5754,N_8431);
and U10215 (N_10215,N_9469,N_7053);
nand U10216 (N_10216,N_7917,N_6535);
nor U10217 (N_10217,N_8089,N_8846);
nor U10218 (N_10218,N_7514,N_7749);
nand U10219 (N_10219,N_8351,N_7575);
or U10220 (N_10220,N_8988,N_8504);
or U10221 (N_10221,N_8927,N_7862);
xnor U10222 (N_10222,N_9120,N_5319);
nand U10223 (N_10223,N_8843,N_6284);
or U10224 (N_10224,N_7518,N_9007);
or U10225 (N_10225,N_5568,N_6458);
nand U10226 (N_10226,N_7790,N_7205);
and U10227 (N_10227,N_6941,N_5560);
nor U10228 (N_10228,N_9169,N_6503);
nand U10229 (N_10229,N_6758,N_7285);
nor U10230 (N_10230,N_9866,N_6673);
and U10231 (N_10231,N_7911,N_5556);
or U10232 (N_10232,N_9871,N_9369);
xor U10233 (N_10233,N_7688,N_9933);
or U10234 (N_10234,N_6883,N_5681);
nor U10235 (N_10235,N_8331,N_8204);
nor U10236 (N_10236,N_7861,N_8560);
nand U10237 (N_10237,N_7014,N_8564);
xor U10238 (N_10238,N_8244,N_9112);
or U10239 (N_10239,N_5576,N_7571);
and U10240 (N_10240,N_6133,N_9520);
nand U10241 (N_10241,N_8220,N_8735);
nand U10242 (N_10242,N_5208,N_7193);
or U10243 (N_10243,N_8266,N_7297);
nand U10244 (N_10244,N_9793,N_9480);
or U10245 (N_10245,N_8824,N_6000);
nor U10246 (N_10246,N_6175,N_9605);
nor U10247 (N_10247,N_7211,N_5228);
and U10248 (N_10248,N_7454,N_8558);
nor U10249 (N_10249,N_7299,N_5648);
or U10250 (N_10250,N_5130,N_9377);
nand U10251 (N_10251,N_5995,N_5543);
nand U10252 (N_10252,N_5495,N_9897);
nand U10253 (N_10253,N_9398,N_9905);
and U10254 (N_10254,N_6131,N_8424);
and U10255 (N_10255,N_9955,N_6408);
nor U10256 (N_10256,N_5801,N_6733);
nor U10257 (N_10257,N_6849,N_9746);
and U10258 (N_10258,N_5231,N_6923);
nor U10259 (N_10259,N_6484,N_9461);
nand U10260 (N_10260,N_6047,N_9251);
xnor U10261 (N_10261,N_5749,N_8864);
nand U10262 (N_10262,N_6282,N_9238);
nand U10263 (N_10263,N_5738,N_5660);
or U10264 (N_10264,N_9215,N_9133);
nor U10265 (N_10265,N_6556,N_7470);
xor U10266 (N_10266,N_7408,N_5925);
or U10267 (N_10267,N_6141,N_5840);
nor U10268 (N_10268,N_6129,N_7644);
nor U10269 (N_10269,N_5816,N_6144);
nand U10270 (N_10270,N_5870,N_5241);
nand U10271 (N_10271,N_9211,N_9415);
nor U10272 (N_10272,N_9594,N_5105);
xnor U10273 (N_10273,N_6313,N_6301);
or U10274 (N_10274,N_9953,N_5984);
nor U10275 (N_10275,N_7494,N_9368);
and U10276 (N_10276,N_5003,N_6645);
nor U10277 (N_10277,N_8482,N_9295);
nand U10278 (N_10278,N_6092,N_7144);
and U10279 (N_10279,N_5427,N_9827);
xor U10280 (N_10280,N_7277,N_5972);
nor U10281 (N_10281,N_9631,N_5036);
xnor U10282 (N_10282,N_5919,N_5116);
or U10283 (N_10283,N_8337,N_6168);
nand U10284 (N_10284,N_8335,N_7851);
or U10285 (N_10285,N_5478,N_9943);
or U10286 (N_10286,N_7812,N_8316);
or U10287 (N_10287,N_8543,N_8677);
or U10288 (N_10288,N_6021,N_8470);
nor U10289 (N_10289,N_7261,N_5086);
or U10290 (N_10290,N_9994,N_5466);
or U10291 (N_10291,N_7976,N_8875);
and U10292 (N_10292,N_6087,N_9443);
nor U10293 (N_10293,N_8313,N_8075);
or U10294 (N_10294,N_9769,N_7421);
nand U10295 (N_10295,N_5480,N_6100);
nor U10296 (N_10296,N_5764,N_5888);
nand U10297 (N_10297,N_5578,N_5154);
and U10298 (N_10298,N_5079,N_8940);
and U10299 (N_10299,N_6875,N_5015);
xnor U10300 (N_10300,N_7220,N_6153);
and U10301 (N_10301,N_5454,N_6999);
nor U10302 (N_10302,N_6628,N_6006);
nor U10303 (N_10303,N_7884,N_5185);
nand U10304 (N_10304,N_7909,N_6017);
xor U10305 (N_10305,N_9414,N_8366);
nor U10306 (N_10306,N_9764,N_9358);
or U10307 (N_10307,N_9370,N_6738);
or U10308 (N_10308,N_9988,N_5708);
xnor U10309 (N_10309,N_7604,N_6671);
nand U10310 (N_10310,N_7329,N_6151);
and U10311 (N_10311,N_9585,N_8994);
and U10312 (N_10312,N_9657,N_6249);
and U10313 (N_10313,N_7493,N_5561);
or U10314 (N_10314,N_6598,N_8779);
and U10315 (N_10315,N_9072,N_8700);
nor U10316 (N_10316,N_8099,N_5355);
xnor U10317 (N_10317,N_6186,N_9670);
nand U10318 (N_10318,N_8215,N_9946);
nor U10319 (N_10319,N_9253,N_5908);
nor U10320 (N_10320,N_9335,N_8462);
or U10321 (N_10321,N_6348,N_5777);
nand U10322 (N_10322,N_9900,N_5161);
xnor U10323 (N_10323,N_9452,N_6602);
nand U10324 (N_10324,N_7464,N_8043);
and U10325 (N_10325,N_8008,N_6031);
nor U10326 (N_10326,N_6810,N_9921);
xor U10327 (N_10327,N_8390,N_7206);
nor U10328 (N_10328,N_9039,N_5627);
or U10329 (N_10329,N_7313,N_7872);
or U10330 (N_10330,N_9166,N_8783);
nand U10331 (N_10331,N_9621,N_8893);
and U10332 (N_10332,N_5395,N_9633);
nor U10333 (N_10333,N_6582,N_8378);
or U10334 (N_10334,N_7453,N_5633);
or U10335 (N_10335,N_6101,N_9317);
nand U10336 (N_10336,N_9136,N_7430);
and U10337 (N_10337,N_8498,N_7811);
or U10338 (N_10338,N_8487,N_9884);
nand U10339 (N_10339,N_5944,N_5254);
or U10340 (N_10340,N_7702,N_7920);
nor U10341 (N_10341,N_9828,N_9898);
xnor U10342 (N_10342,N_5437,N_9363);
nand U10343 (N_10343,N_6217,N_6209);
nand U10344 (N_10344,N_7476,N_5831);
or U10345 (N_10345,N_6725,N_9926);
xor U10346 (N_10346,N_5093,N_8753);
or U10347 (N_10347,N_6202,N_5173);
or U10348 (N_10348,N_8072,N_5039);
nand U10349 (N_10349,N_5907,N_9567);
and U10350 (N_10350,N_8655,N_7724);
nor U10351 (N_10351,N_5686,N_6690);
xnor U10352 (N_10352,N_7307,N_6872);
nor U10353 (N_10353,N_5181,N_6173);
or U10354 (N_10354,N_9061,N_9371);
nor U10355 (N_10355,N_7015,N_6976);
or U10356 (N_10356,N_7735,N_6631);
and U10357 (N_10357,N_6233,N_9526);
or U10358 (N_10358,N_9913,N_9402);
and U10359 (N_10359,N_5268,N_9922);
and U10360 (N_10360,N_5784,N_5849);
nand U10361 (N_10361,N_9367,N_6824);
or U10362 (N_10362,N_9803,N_9294);
and U10363 (N_10363,N_5089,N_7786);
and U10364 (N_10364,N_5821,N_6050);
or U10365 (N_10365,N_6679,N_8422);
or U10366 (N_10366,N_8046,N_5169);
and U10367 (N_10367,N_7537,N_5425);
nand U10368 (N_10368,N_5134,N_5082);
nand U10369 (N_10369,N_8652,N_7881);
xor U10370 (N_10370,N_8923,N_7896);
or U10371 (N_10371,N_7341,N_6425);
and U10372 (N_10372,N_8617,N_6653);
nor U10373 (N_10373,N_6085,N_8001);
nor U10374 (N_10374,N_5957,N_7141);
nand U10375 (N_10375,N_6794,N_6201);
and U10376 (N_10376,N_6698,N_8449);
nor U10377 (N_10377,N_8722,N_9767);
nor U10378 (N_10378,N_7535,N_7068);
xor U10379 (N_10379,N_6188,N_8222);
and U10380 (N_10380,N_8630,N_6646);
nor U10381 (N_10381,N_5853,N_6658);
nor U10382 (N_10382,N_8835,N_7835);
nor U10383 (N_10383,N_5051,N_9620);
xor U10384 (N_10384,N_8038,N_7356);
and U10385 (N_10385,N_6150,N_5547);
or U10386 (N_10386,N_8398,N_5654);
nand U10387 (N_10387,N_6364,N_7830);
xnor U10388 (N_10388,N_8759,N_6135);
and U10389 (N_10389,N_5737,N_5673);
xor U10390 (N_10390,N_5858,N_5700);
and U10391 (N_10391,N_8855,N_8101);
xor U10392 (N_10392,N_9272,N_8445);
or U10393 (N_10393,N_9357,N_5885);
nor U10394 (N_10394,N_9054,N_6586);
nand U10395 (N_10395,N_5284,N_7257);
nor U10396 (N_10396,N_7226,N_6116);
xor U10397 (N_10397,N_5270,N_6412);
and U10398 (N_10398,N_7246,N_9588);
xnor U10399 (N_10399,N_9604,N_9204);
or U10400 (N_10400,N_6732,N_7364);
nand U10401 (N_10401,N_5954,N_6804);
nor U10402 (N_10402,N_8407,N_6125);
xnor U10403 (N_10403,N_9839,N_9122);
nand U10404 (N_10404,N_6040,N_6678);
nand U10405 (N_10405,N_5360,N_7044);
nor U10406 (N_10406,N_6270,N_5792);
nand U10407 (N_10407,N_7371,N_7184);
nor U10408 (N_10408,N_9161,N_6061);
xnor U10409 (N_10409,N_6846,N_7160);
or U10410 (N_10410,N_6389,N_9606);
or U10411 (N_10411,N_7636,N_9805);
xnor U10412 (N_10412,N_6597,N_9962);
nor U10413 (N_10413,N_7047,N_7166);
or U10414 (N_10414,N_7346,N_6410);
xor U10415 (N_10415,N_8414,N_6239);
or U10416 (N_10416,N_5330,N_8248);
nand U10417 (N_10417,N_7087,N_6114);
xor U10418 (N_10418,N_9395,N_8627);
or U10419 (N_10419,N_5474,N_7446);
nand U10420 (N_10420,N_6199,N_5323);
nand U10421 (N_10421,N_7664,N_9524);
or U10422 (N_10422,N_9305,N_6662);
or U10423 (N_10423,N_5256,N_8287);
nor U10424 (N_10424,N_9986,N_7244);
and U10425 (N_10425,N_7782,N_7879);
or U10426 (N_10426,N_8749,N_5406);
nand U10427 (N_10427,N_7965,N_5676);
xor U10428 (N_10428,N_8530,N_5156);
and U10429 (N_10429,N_6600,N_5057);
nor U10430 (N_10430,N_9945,N_9430);
nand U10431 (N_10431,N_9372,N_6895);
nand U10432 (N_10432,N_7953,N_7898);
and U10433 (N_10433,N_5828,N_7713);
xnor U10434 (N_10434,N_8953,N_5065);
nand U10435 (N_10435,N_8738,N_9653);
or U10436 (N_10436,N_9507,N_9096);
or U10437 (N_10437,N_8154,N_6327);
nand U10438 (N_10438,N_9798,N_7292);
or U10439 (N_10439,N_5971,N_5193);
nand U10440 (N_10440,N_5799,N_6718);
and U10441 (N_10441,N_6250,N_8148);
nand U10442 (N_10442,N_9464,N_5449);
nor U10443 (N_10443,N_7810,N_5940);
and U10444 (N_10444,N_8968,N_6401);
and U10445 (N_10445,N_9245,N_7363);
nor U10446 (N_10446,N_5489,N_6487);
and U10447 (N_10447,N_5191,N_6587);
nand U10448 (N_10448,N_8724,N_8288);
or U10449 (N_10449,N_5485,N_9515);
and U10450 (N_10450,N_5421,N_6007);
and U10451 (N_10451,N_6044,N_5428);
nand U10452 (N_10452,N_9059,N_6966);
nor U10453 (N_10453,N_8917,N_6300);
or U10454 (N_10454,N_9593,N_9961);
and U10455 (N_10455,N_6456,N_9246);
and U10456 (N_10456,N_7525,N_6366);
or U10457 (N_10457,N_5997,N_7995);
or U10458 (N_10458,N_7598,N_9279);
or U10459 (N_10459,N_7723,N_5486);
and U10460 (N_10460,N_6413,N_8834);
xor U10461 (N_10461,N_8415,N_5796);
nand U10462 (N_10462,N_6553,N_6609);
and U10463 (N_10463,N_5329,N_6692);
or U10464 (N_10464,N_7926,N_6332);
or U10465 (N_10465,N_7585,N_7129);
nand U10466 (N_10466,N_9448,N_7937);
nand U10467 (N_10467,N_5933,N_5856);
nand U10468 (N_10468,N_5027,N_8421);
xor U10469 (N_10469,N_7034,N_5320);
nor U10470 (N_10470,N_6591,N_5264);
or U10471 (N_10471,N_7151,N_5195);
or U10472 (N_10472,N_5747,N_9102);
or U10473 (N_10473,N_8419,N_5601);
and U10474 (N_10474,N_7389,N_7955);
and U10475 (N_10475,N_8392,N_6034);
or U10476 (N_10476,N_6915,N_7481);
nand U10477 (N_10477,N_9247,N_7661);
and U10478 (N_10478,N_9044,N_6037);
xnor U10479 (N_10479,N_6418,N_8368);
and U10480 (N_10480,N_5565,N_5061);
or U10481 (N_10481,N_5211,N_7725);
nor U10482 (N_10482,N_6937,N_7085);
nand U10483 (N_10483,N_9608,N_8899);
and U10484 (N_10484,N_9568,N_8646);
nand U10485 (N_10485,N_9812,N_5356);
nor U10486 (N_10486,N_9031,N_7336);
nand U10487 (N_10487,N_5372,N_7549);
and U10488 (N_10488,N_5324,N_7042);
nand U10489 (N_10489,N_8795,N_6689);
xor U10490 (N_10490,N_5436,N_5746);
nor U10491 (N_10491,N_8026,N_7900);
nor U10492 (N_10492,N_6371,N_8323);
nand U10493 (N_10493,N_5021,N_6633);
and U10494 (N_10494,N_6978,N_5418);
or U10495 (N_10495,N_7274,N_7846);
xor U10496 (N_10496,N_6053,N_8884);
or U10497 (N_10497,N_6734,N_7097);
and U10498 (N_10498,N_8301,N_7663);
nor U10499 (N_10499,N_8750,N_8709);
nand U10500 (N_10500,N_8439,N_8258);
or U10501 (N_10501,N_9168,N_7283);
and U10502 (N_10502,N_5705,N_7935);
xnor U10503 (N_10503,N_8547,N_5203);
or U10504 (N_10504,N_8136,N_7026);
or U10505 (N_10505,N_9570,N_5910);
nor U10506 (N_10506,N_8508,N_7704);
xnor U10507 (N_10507,N_9648,N_9819);
nand U10508 (N_10508,N_5852,N_7589);
or U10509 (N_10509,N_5236,N_8355);
or U10510 (N_10510,N_8955,N_7000);
nand U10511 (N_10511,N_6281,N_5423);
and U10512 (N_10512,N_7709,N_5929);
nand U10513 (N_10513,N_5528,N_6392);
xor U10514 (N_10514,N_7472,N_6853);
and U10515 (N_10515,N_5687,N_8745);
and U10516 (N_10516,N_8133,N_6324);
nor U10517 (N_10517,N_6343,N_5780);
nor U10518 (N_10518,N_5918,N_7868);
and U10519 (N_10519,N_8752,N_5920);
or U10520 (N_10520,N_8509,N_6681);
and U10521 (N_10521,N_9047,N_6063);
nand U10522 (N_10522,N_9062,N_7385);
xnor U10523 (N_10523,N_5206,N_6789);
or U10524 (N_10524,N_6561,N_5832);
nor U10525 (N_10525,N_9539,N_6524);
nand U10526 (N_10526,N_6420,N_7647);
nor U10527 (N_10527,N_6383,N_7186);
or U10528 (N_10528,N_8264,N_5672);
or U10529 (N_10529,N_5394,N_6912);
and U10530 (N_10530,N_8118,N_5362);
and U10531 (N_10531,N_8389,N_6278);
or U10532 (N_10532,N_7947,N_6179);
or U10533 (N_10533,N_9356,N_7367);
and U10534 (N_10534,N_5664,N_8624);
or U10535 (N_10535,N_9824,N_9777);
nor U10536 (N_10536,N_8080,N_7886);
nor U10537 (N_10537,N_5354,N_5864);
nand U10538 (N_10538,N_8224,N_8036);
and U10539 (N_10539,N_7024,N_6122);
and U10540 (N_10540,N_6821,N_9822);
and U10541 (N_10541,N_6158,N_6608);
and U10542 (N_10542,N_7077,N_5433);
or U10543 (N_10543,N_8245,N_7096);
and U10544 (N_10544,N_5677,N_6685);
nand U10545 (N_10545,N_9713,N_9037);
or U10546 (N_10546,N_5107,N_7412);
xnor U10547 (N_10547,N_5233,N_6925);
xor U10548 (N_10548,N_7316,N_6099);
or U10549 (N_10549,N_5987,N_6581);
xnor U10550 (N_10550,N_7816,N_7652);
nand U10551 (N_10551,N_8079,N_5043);
or U10552 (N_10552,N_6137,N_5887);
or U10553 (N_10553,N_6502,N_7582);
xnor U10554 (N_10554,N_5642,N_9419);
xor U10555 (N_10555,N_5392,N_8194);
or U10556 (N_10556,N_9382,N_5787);
nor U10557 (N_10557,N_9410,N_9867);
xnor U10558 (N_10558,N_9327,N_6384);
nor U10559 (N_10559,N_6419,N_9486);
or U10560 (N_10560,N_9589,N_8395);
or U10561 (N_10561,N_5155,N_8488);
nor U10562 (N_10562,N_6455,N_5373);
nor U10563 (N_10563,N_6065,N_5479);
and U10564 (N_10564,N_7400,N_5122);
nor U10565 (N_10565,N_8456,N_8317);
xnor U10566 (N_10566,N_5458,N_7303);
and U10567 (N_10567,N_8166,N_8022);
nor U10568 (N_10568,N_6702,N_6058);
nand U10569 (N_10569,N_5090,N_5609);
nor U10570 (N_10570,N_7269,N_5793);
and U10571 (N_10571,N_9344,N_6840);
and U10572 (N_10572,N_8659,N_7225);
nand U10573 (N_10573,N_9113,N_5978);
and U10574 (N_10574,N_9139,N_8361);
or U10575 (N_10575,N_8649,N_5766);
or U10576 (N_10576,N_8437,N_9651);
nor U10577 (N_10577,N_5331,N_7940);
nand U10578 (N_10578,N_6548,N_8039);
or U10579 (N_10579,N_6884,N_8501);
xor U10580 (N_10580,N_5584,N_5144);
nand U10581 (N_10581,N_6924,N_9538);
or U10582 (N_10582,N_5285,N_5725);
nand U10583 (N_10583,N_9680,N_5742);
nand U10584 (N_10584,N_9616,N_8053);
or U10585 (N_10585,N_8634,N_6590);
nor U10586 (N_10586,N_5299,N_7908);
xnor U10587 (N_10587,N_6985,N_6549);
nor U10588 (N_10588,N_8202,N_5847);
nand U10589 (N_10589,N_5200,N_7117);
nand U10590 (N_10590,N_9456,N_7132);
nand U10591 (N_10591,N_8920,N_9887);
xor U10592 (N_10592,N_5838,N_8359);
xnor U10593 (N_10593,N_8471,N_9535);
or U10594 (N_10594,N_5443,N_7495);
or U10595 (N_10595,N_7880,N_5237);
or U10596 (N_10596,N_9413,N_5639);
and U10597 (N_10597,N_6532,N_6936);
nand U10598 (N_10598,N_7506,N_5774);
and U10599 (N_10599,N_8004,N_7587);
nor U10600 (N_10600,N_9927,N_8663);
xor U10601 (N_10601,N_7807,N_8117);
or U10602 (N_10602,N_9438,N_6340);
nand U10603 (N_10603,N_8971,N_8306);
or U10604 (N_10604,N_9347,N_8242);
or U10605 (N_10605,N_9242,N_8256);
nand U10606 (N_10606,N_9796,N_9278);
and U10607 (N_10607,N_7509,N_8977);
and U10608 (N_10608,N_8123,N_9649);
xor U10609 (N_10609,N_6650,N_8382);
nand U10610 (N_10610,N_5247,N_8055);
nand U10611 (N_10611,N_9227,N_9542);
or U10612 (N_10612,N_8796,N_7547);
nand U10613 (N_10613,N_9514,N_7593);
and U10614 (N_10614,N_8744,N_7154);
nor U10615 (N_10615,N_8083,N_9277);
nor U10616 (N_10616,N_5432,N_6084);
and U10617 (N_10617,N_5187,N_5912);
nand U10618 (N_10618,N_6907,N_9848);
or U10619 (N_10619,N_8718,N_9200);
nand U10620 (N_10620,N_6437,N_5698);
and U10621 (N_10621,N_7974,N_6857);
nor U10622 (N_10622,N_8223,N_7200);
nand U10623 (N_10623,N_9065,N_8237);
nor U10624 (N_10624,N_8477,N_6365);
or U10625 (N_10625,N_9896,N_9420);
or U10626 (N_10626,N_5151,N_6112);
or U10627 (N_10627,N_6664,N_8566);
nor U10628 (N_10628,N_8743,N_7771);
nand U10629 (N_10629,N_8153,N_6495);
nor U10630 (N_10630,N_6139,N_5720);
nor U10631 (N_10631,N_5622,N_7510);
or U10632 (N_10632,N_7115,N_6191);
nor U10633 (N_10633,N_5692,N_9153);
and U10634 (N_10634,N_7216,N_6862);
nand U10635 (N_10635,N_7311,N_7705);
nand U10636 (N_10636,N_5260,N_9256);
nand U10637 (N_10637,N_6776,N_7195);
or U10638 (N_10638,N_6305,N_5614);
and U10639 (N_10639,N_5234,N_7669);
nor U10640 (N_10640,N_5251,N_8033);
and U10641 (N_10641,N_8751,N_5949);
nand U10642 (N_10642,N_8841,N_8144);
or U10643 (N_10643,N_5894,N_5170);
nor U10644 (N_10644,N_8519,N_8938);
xor U10645 (N_10645,N_7625,N_7583);
or U10646 (N_10646,N_8265,N_6352);
nand U10647 (N_10647,N_6388,N_5397);
nor U10648 (N_10648,N_9250,N_7546);
and U10649 (N_10649,N_7322,N_7066);
and U10650 (N_10650,N_9555,N_5240);
nand U10651 (N_10651,N_9689,N_6312);
and U10652 (N_10652,N_8728,N_5651);
nand U10653 (N_10653,N_6356,N_9041);
nand U10654 (N_10654,N_5238,N_5294);
or U10655 (N_10655,N_5129,N_5300);
nor U10656 (N_10656,N_9712,N_9985);
nor U10657 (N_10657,N_5457,N_9661);
and U10658 (N_10658,N_7164,N_5098);
nand U10659 (N_10659,N_9586,N_7301);
and U10660 (N_10660,N_8733,N_6684);
or U10661 (N_10661,N_9034,N_6930);
xor U10662 (N_10662,N_5523,N_5647);
xnor U10663 (N_10663,N_7388,N_5950);
and U10664 (N_10664,N_6334,N_6905);
or U10665 (N_10665,N_8771,N_5631);
and U10666 (N_10666,N_7870,N_7071);
nor U10667 (N_10667,N_7451,N_9809);
or U10668 (N_10668,N_8936,N_5970);
and U10669 (N_10669,N_6363,N_6130);
or U10670 (N_10670,N_6539,N_7212);
or U10671 (N_10671,N_8583,N_7635);
nand U10672 (N_10672,N_6956,N_6808);
nor U10673 (N_10673,N_9138,N_5490);
and U10674 (N_10674,N_8364,N_9181);
nor U10675 (N_10675,N_9422,N_9557);
nand U10676 (N_10676,N_5807,N_8236);
xnor U10677 (N_10677,N_7805,N_6911);
xnor U10678 (N_10678,N_5249,N_7847);
nand U10679 (N_10679,N_9773,N_5253);
and U10680 (N_10680,N_5398,N_7473);
or U10681 (N_10681,N_5464,N_5721);
nand U10682 (N_10682,N_5382,N_7475);
nand U10683 (N_10683,N_5340,N_7479);
or U10684 (N_10684,N_5183,N_8551);
nor U10685 (N_10685,N_9095,N_9383);
or U10686 (N_10686,N_9303,N_7183);
nor U10687 (N_10687,N_8786,N_7420);
and U10688 (N_10688,N_8358,N_8027);
or U10689 (N_10689,N_8465,N_5966);
or U10690 (N_10690,N_9957,N_8836);
nor U10691 (N_10691,N_6754,N_6731);
nor U10692 (N_10692,N_5671,N_8259);
or U10693 (N_10693,N_6450,N_7832);
or U10694 (N_10694,N_9468,N_7877);
xnor U10695 (N_10695,N_5198,N_7733);
nor U10696 (N_10696,N_8676,N_8961);
nor U10697 (N_10697,N_9708,N_6496);
and U10698 (N_10698,N_6082,N_7519);
nand U10699 (N_10699,N_8349,N_9976);
and U10700 (N_10700,N_9009,N_5955);
xnor U10701 (N_10701,N_8391,N_7452);
xor U10702 (N_10702,N_6563,N_6274);
and U10703 (N_10703,N_8707,N_5782);
nand U10704 (N_10704,N_7444,N_6051);
nand U10705 (N_10705,N_8436,N_8691);
nand U10706 (N_10706,N_8320,N_9212);
nand U10707 (N_10707,N_7804,N_5945);
and U10708 (N_10708,N_9190,N_6020);
nor U10709 (N_10709,N_9088,N_8912);
and U10710 (N_10710,N_7951,N_7057);
nand U10711 (N_10711,N_8712,N_7590);
nand U10712 (N_10712,N_6023,N_9877);
nand U10713 (N_10713,N_6329,N_7787);
nand U10714 (N_10714,N_8307,N_8792);
and U10715 (N_10715,N_8458,N_6118);
nand U10716 (N_10716,N_5308,N_8403);
or U10717 (N_10717,N_7486,N_8908);
nor U10718 (N_10718,N_8605,N_7373);
nand U10719 (N_10719,N_8523,N_9220);
nand U10720 (N_10720,N_9266,N_7445);
and U10721 (N_10721,N_9330,N_5327);
nand U10722 (N_10722,N_7354,N_7060);
and U10723 (N_10723,N_9667,N_8516);
nor U10724 (N_10724,N_8068,N_9048);
nor U10725 (N_10725,N_7443,N_9956);
nor U10726 (N_10726,N_5292,N_9263);
or U10727 (N_10727,N_6945,N_7646);
or U10728 (N_10728,N_5960,N_8108);
nor U10729 (N_10729,N_8963,N_8348);
nand U10730 (N_10730,N_8665,N_8717);
or U10731 (N_10731,N_5164,N_9101);
nand U10732 (N_10732,N_8623,N_5370);
or U10733 (N_10733,N_5520,N_9029);
and U10734 (N_10734,N_6064,N_6438);
and U10735 (N_10735,N_5410,N_7335);
xor U10736 (N_10736,N_8370,N_6656);
nor U10737 (N_10737,N_9384,N_9085);
nand U10738 (N_10738,N_8643,N_6863);
nor U10739 (N_10739,N_8734,N_6740);
or U10740 (N_10740,N_8492,N_5325);
and U10741 (N_10741,N_8042,N_5958);
and U10742 (N_10742,N_7078,N_6185);
nor U10743 (N_10743,N_5791,N_6288);
nand U10744 (N_10744,N_6783,N_6255);
or U10745 (N_10745,N_6355,N_9308);
or U10746 (N_10746,N_9719,N_6747);
nand U10747 (N_10747,N_6347,N_9321);
nand U10748 (N_10748,N_9487,N_9610);
nor U10749 (N_10749,N_5555,N_7442);
nand U10750 (N_10750,N_7596,N_9396);
or U10751 (N_10751,N_8822,N_5808);
nand U10752 (N_10752,N_6529,N_7676);
or U10753 (N_10753,N_8339,N_9355);
nor U10754 (N_10754,N_8828,N_7932);
nor U10755 (N_10755,N_5346,N_9106);
and U10756 (N_10756,N_9477,N_6169);
and U10757 (N_10757,N_9100,N_7760);
and U10758 (N_10758,N_7070,N_8460);
and U10759 (N_10759,N_7394,N_8704);
nand U10760 (N_10760,N_5069,N_5445);
and U10761 (N_10761,N_5350,N_6596);
or U10762 (N_10762,N_5875,N_7152);
nand U10763 (N_10763,N_8119,N_6323);
nand U10764 (N_10764,N_6604,N_8522);
nor U10765 (N_10765,N_8737,N_9262);
nor U10766 (N_10766,N_6893,N_5152);
nand U10767 (N_10767,N_5594,N_9574);
or U10768 (N_10768,N_6917,N_6617);
nor U10769 (N_10769,N_7127,N_9533);
or U10770 (N_10770,N_8239,N_5953);
nand U10771 (N_10771,N_9647,N_7623);
and U10772 (N_10772,N_8702,N_9160);
nor U10773 (N_10773,N_6042,N_8594);
nor U10774 (N_10774,N_7123,N_9951);
xor U10775 (N_10775,N_6947,N_7883);
and U10776 (N_10776,N_5364,N_9879);
or U10777 (N_10777,N_8690,N_5804);
nand U10778 (N_10778,N_9625,N_6801);
or U10779 (N_10779,N_7762,N_8451);
nand U10780 (N_10780,N_6474,N_5220);
and U10781 (N_10781,N_9173,N_9600);
and U10782 (N_10782,N_9747,N_9254);
nor U10783 (N_10783,N_8739,N_7368);
and U10784 (N_10784,N_8096,N_5931);
and U10785 (N_10785,N_7137,N_5739);
or U10786 (N_10786,N_6190,N_5608);
or U10787 (N_10787,N_7801,N_8073);
and U10788 (N_10788,N_9494,N_9450);
nand U10789 (N_10789,N_8464,N_6676);
nand U10790 (N_10790,N_6926,N_5851);
xor U10791 (N_10791,N_6592,N_6796);
nand U10792 (N_10792,N_9092,N_7290);
nor U10793 (N_10793,N_5046,N_7856);
xnor U10794 (N_10794,N_9340,N_8911);
nand U10795 (N_10795,N_6973,N_5289);
nor U10796 (N_10796,N_7375,N_7276);
or U10797 (N_10797,N_9741,N_5625);
nor U10798 (N_10798,N_7923,N_5055);
and U10799 (N_10799,N_8620,N_7120);
and U10800 (N_10800,N_5499,N_5312);
and U10801 (N_10801,N_9361,N_9624);
nand U10802 (N_10802,N_5854,N_8050);
or U10803 (N_10803,N_8791,N_7360);
nor U10804 (N_10804,N_7980,N_6237);
and U10805 (N_10805,N_7496,N_5509);
or U10806 (N_10806,N_5538,N_7009);
or U10807 (N_10807,N_7243,N_7680);
and U10808 (N_10808,N_6766,N_8010);
or U10809 (N_10809,N_7860,N_8638);
or U10810 (N_10810,N_8435,N_7973);
nor U10811 (N_10811,N_6786,N_5730);
nor U10812 (N_10812,N_6928,N_9425);
or U10813 (N_10813,N_6387,N_6573);
nor U10814 (N_10814,N_5515,N_8510);
and U10815 (N_10815,N_9757,N_9863);
nor U10816 (N_10816,N_7404,N_5494);
nand U10817 (N_10817,N_8705,N_7559);
or U10818 (N_10818,N_8625,N_9995);
nand U10819 (N_10819,N_5075,N_5343);
and U10820 (N_10820,N_5045,N_5371);
and U10821 (N_10821,N_8180,N_6854);
nor U10822 (N_10822,N_5716,N_7095);
or U10823 (N_10823,N_9918,N_9375);
and U10824 (N_10824,N_9966,N_7130);
and U10825 (N_10825,N_9182,N_9436);
xnor U10826 (N_10826,N_6453,N_9825);
nand U10827 (N_10827,N_8472,N_6555);
or U10828 (N_10828,N_8060,N_8972);
and U10829 (N_10829,N_5465,N_9171);
nand U10830 (N_10830,N_6855,N_6086);
or U10831 (N_10831,N_8896,N_7640);
or U10832 (N_10832,N_5983,N_5969);
nand U10833 (N_10833,N_5785,N_5047);
or U10834 (N_10834,N_7172,N_8467);
or U10835 (N_10835,N_6093,N_9580);
nand U10836 (N_10836,N_6176,N_8003);
and U10837 (N_10837,N_6154,N_7672);
and U10838 (N_10838,N_6195,N_6381);
or U10839 (N_10839,N_6367,N_9217);
nor U10840 (N_10840,N_6253,N_9845);
or U10841 (N_10841,N_5696,N_5463);
xnor U10842 (N_10842,N_9269,N_6847);
and U10843 (N_10843,N_8847,N_7284);
and U10844 (N_10844,N_6198,N_5638);
xnor U10845 (N_10845,N_6688,N_9437);
nand U10846 (N_10846,N_8171,N_9528);
nor U10847 (N_10847,N_9203,N_8524);
or U10848 (N_10848,N_7149,N_7169);
xnor U10849 (N_10849,N_6665,N_9108);
nor U10850 (N_10850,N_5099,N_6225);
or U10851 (N_10851,N_7891,N_7701);
nand U10852 (N_10852,N_8120,N_8243);
nand U10853 (N_10853,N_8495,N_6686);
nand U10854 (N_10854,N_9783,N_6358);
nand U10855 (N_10855,N_7708,N_8189);
xnor U10856 (N_10856,N_8127,N_9270);
and U10857 (N_10857,N_5301,N_9944);
or U10858 (N_10858,N_8116,N_7401);
nand U10859 (N_10859,N_5915,N_9293);
and U10860 (N_10860,N_6626,N_9908);
xnor U10861 (N_10861,N_9332,N_6998);
and U10862 (N_10862,N_8255,N_9491);
xor U10863 (N_10863,N_6501,N_9885);
xor U10864 (N_10864,N_5834,N_7428);
nor U10865 (N_10865,N_8169,N_9067);
xnor U10866 (N_10866,N_6431,N_6891);
and U10867 (N_10867,N_7692,N_6874);
and U10868 (N_10868,N_5605,N_8365);
nor U10869 (N_10869,N_6443,N_7797);
or U10870 (N_10870,N_7707,N_6687);
or U10871 (N_10871,N_9928,N_8696);
and U10872 (N_10872,N_6142,N_8078);
and U10873 (N_10873,N_9607,N_7437);
or U10874 (N_10874,N_8085,N_5013);
nor U10875 (N_10875,N_7942,N_7668);
and U10876 (N_10876,N_5491,N_9675);
nand U10877 (N_10877,N_9935,N_5653);
nor U10878 (N_10878,N_6830,N_5723);
nor U10879 (N_10879,N_5345,N_9659);
nor U10880 (N_10880,N_5145,N_8754);
and U10881 (N_10881,N_5508,N_5488);
or U10882 (N_10882,N_6951,N_6767);
nor U10883 (N_10883,N_9732,N_5563);
and U10884 (N_10884,N_6869,N_5332);
and U10885 (N_10885,N_8859,N_7300);
nor U10886 (N_10886,N_5736,N_7259);
nor U10887 (N_10887,N_7038,N_6070);
or U10888 (N_10888,N_7779,N_5817);
or U10889 (N_10889,N_5452,N_5298);
nand U10890 (N_10890,N_5504,N_7075);
nor U10891 (N_10891,N_8268,N_5789);
nand U10892 (N_10892,N_6030,N_5822);
xor U10893 (N_10893,N_6511,N_9042);
or U10894 (N_10894,N_5182,N_7192);
or U10895 (N_10895,N_7802,N_9802);
xor U10896 (N_10896,N_6102,N_7266);
xor U10897 (N_10897,N_6864,N_7381);
nand U10898 (N_10898,N_9942,N_6803);
xnor U10899 (N_10899,N_8137,N_8310);
or U10900 (N_10900,N_8546,N_5031);
nor U10901 (N_10901,N_7597,N_5008);
or U10902 (N_10902,N_5839,N_9709);
or U10903 (N_10903,N_5682,N_8305);
and U10904 (N_10904,N_6104,N_6557);
or U10905 (N_10905,N_8808,N_5399);
xnor U10906 (N_10906,N_7349,N_6273);
or U10907 (N_10907,N_6811,N_8746);
xor U10908 (N_10908,N_8035,N_5546);
and U10909 (N_10909,N_5591,N_8815);
nor U10910 (N_10910,N_8241,N_7887);
xor U10911 (N_10911,N_6823,N_6703);
xnor U10912 (N_10912,N_5936,N_6261);
nor U10913 (N_10913,N_8219,N_6374);
and U10914 (N_10914,N_8253,N_7731);
and U10915 (N_10915,N_5775,N_5172);
and U10916 (N_10916,N_8726,N_8973);
nand U10917 (N_10917,N_9751,N_6156);
nand U10918 (N_10918,N_9470,N_7700);
xnor U10919 (N_10919,N_9407,N_8084);
and U10920 (N_10920,N_7116,N_8132);
xnor U10921 (N_10921,N_7051,N_9745);
nor U10922 (N_10922,N_6422,N_9851);
nand U10923 (N_10923,N_8755,N_7392);
and U10924 (N_10924,N_7675,N_8344);
nor U10925 (N_10925,N_5108,N_5934);
or U10926 (N_10926,N_9338,N_9849);
nor U10927 (N_10927,N_8329,N_5848);
or U10928 (N_10928,N_8232,N_5818);
and U10929 (N_10929,N_8044,N_7921);
nor U10930 (N_10930,N_7655,N_6739);
nor U10931 (N_10931,N_7090,N_9142);
and U10932 (N_10932,N_7545,N_6016);
and U10933 (N_10933,N_9766,N_9596);
nand U10934 (N_10934,N_7238,N_7397);
and U10935 (N_10935,N_6660,N_5536);
and U10936 (N_10936,N_7618,N_7544);
and U10937 (N_10937,N_7148,N_6536);
nand U10938 (N_10938,N_6331,N_7055);
nand U10939 (N_10939,N_9336,N_9237);
nand U10940 (N_10940,N_8094,N_5377);
xnor U10941 (N_10941,N_6552,N_6264);
or U10942 (N_10942,N_6326,N_9516);
or U10943 (N_10943,N_6710,N_8430);
or U10944 (N_10944,N_5400,N_7383);
nor U10945 (N_10945,N_5976,N_5307);
or U10946 (N_10946,N_5756,N_9916);
or U10947 (N_10947,N_9306,N_7433);
xnor U10948 (N_10948,N_6781,N_6873);
xor U10949 (N_10949,N_8586,N_5462);
or U10950 (N_10950,N_6713,N_8396);
or U10951 (N_10951,N_7606,N_8694);
and U10952 (N_10952,N_7605,N_8499);
or U10953 (N_10953,N_7438,N_9639);
nor U10954 (N_10954,N_8381,N_7619);
nor U10955 (N_10955,N_7712,N_6815);
or U10956 (N_10956,N_7916,N_8103);
or U10957 (N_10957,N_5054,N_8538);
nand U10958 (N_10958,N_9763,N_9816);
and U10959 (N_10959,N_7319,N_6385);
or U10960 (N_10960,N_5023,N_8393);
or U10961 (N_10961,N_8913,N_9716);
xor U10962 (N_10962,N_6648,N_7822);
nand U10963 (N_10963,N_9333,N_7305);
nor U10964 (N_10964,N_5599,N_8830);
nor U10965 (N_10965,N_6229,N_9475);
and U10966 (N_10966,N_9202,N_8186);
nand U10967 (N_10967,N_9360,N_5262);
nor U10968 (N_10968,N_8632,N_8635);
nor U10969 (N_10969,N_6868,N_6248);
nand U10970 (N_10970,N_7350,N_6957);
nand U10971 (N_10971,N_9733,N_6677);
nor U10972 (N_10972,N_7331,N_7323);
nor U10973 (N_10973,N_8801,N_6814);
nand U10974 (N_10974,N_6041,N_6400);
nor U10975 (N_10975,N_6756,N_7108);
nand U10976 (N_10976,N_6497,N_8227);
or U10977 (N_10977,N_9114,N_9239);
and U10978 (N_10978,N_6952,N_5674);
nor U10979 (N_10979,N_7960,N_9018);
nand U10980 (N_10980,N_9569,N_9127);
and U10981 (N_10981,N_5131,N_6470);
nor U10982 (N_10982,N_7809,N_6230);
or U10983 (N_10983,N_7330,N_7584);
and U10984 (N_10984,N_5798,N_5524);
and U10985 (N_10985,N_9550,N_5527);
xnor U10986 (N_10986,N_8191,N_7869);
nand U10987 (N_10987,N_5018,N_9937);
nor U10988 (N_10988,N_7776,N_8765);
nand U10989 (N_10989,N_7189,N_9068);
or U10990 (N_10990,N_7954,N_9298);
nand U10991 (N_10991,N_9658,N_6170);
xor U10992 (N_10992,N_9665,N_8862);
nand U10993 (N_10993,N_9838,N_9449);
nand U10994 (N_10994,N_7970,N_8581);
or U10995 (N_10995,N_7831,N_7045);
or U10996 (N_10996,N_9005,N_8030);
or U10997 (N_10997,N_8517,N_5829);
nor U10998 (N_10998,N_6362,N_7098);
nor U10999 (N_10999,N_9792,N_5419);
nand U11000 (N_11000,N_9969,N_8701);
nor U11001 (N_11001,N_6222,N_6753);
nand U11002 (N_11002,N_8545,N_5697);
nor U11003 (N_11003,N_7698,N_5092);
and U11004 (N_11004,N_9975,N_5909);
nor U11005 (N_11005,N_8681,N_5892);
or U11006 (N_11006,N_8397,N_8575);
nand U11007 (N_11007,N_9189,N_9187);
nor U11008 (N_11008,N_6293,N_8591);
and U11009 (N_11009,N_9500,N_5196);
or U11010 (N_11010,N_9137,N_5007);
xnor U11011 (N_11011,N_7834,N_8775);
xnor U11012 (N_11012,N_7981,N_8376);
or U11013 (N_11013,N_7111,N_8897);
nor U11014 (N_11014,N_6537,N_5311);
nor U11015 (N_11015,N_5123,N_9739);
nor U11016 (N_11016,N_5710,N_7777);
and U11017 (N_11017,N_7424,N_7987);
nor U11018 (N_11018,N_7118,N_7062);
nand U11019 (N_11019,N_5558,N_5091);
and U11020 (N_11020,N_6935,N_7222);
nor U11021 (N_11021,N_5040,N_6126);
or U11022 (N_11022,N_7304,N_9454);
nor U11023 (N_11023,N_8593,N_8983);
and U11024 (N_11024,N_7499,N_7656);
nand U11025 (N_11025,N_7912,N_9929);
and U11026 (N_11026,N_9043,N_9109);
nor U11027 (N_11027,N_9014,N_8685);
nand U11028 (N_11028,N_8826,N_8071);
or U11029 (N_11029,N_8503,N_7288);
and U11030 (N_11030,N_6206,N_9786);
or U11031 (N_11031,N_9010,N_8134);
and U11032 (N_11032,N_9213,N_9143);
and U11033 (N_11033,N_5941,N_8429);
nand U11034 (N_11034,N_5002,N_9053);
and U11035 (N_11035,N_6782,N_9434);
nand U11036 (N_11036,N_6887,N_8947);
nand U11037 (N_11037,N_9706,N_5531);
and U11038 (N_11038,N_9681,N_5810);
nand U11039 (N_11039,N_5243,N_6995);
or U11040 (N_11040,N_6876,N_6193);
and U11041 (N_11041,N_7434,N_8805);
or U11042 (N_11042,N_9260,N_5244);
xor U11043 (N_11043,N_7699,N_7199);
xnor U11044 (N_11044,N_7948,N_6321);
nand U11045 (N_11045,N_5179,N_5094);
or U11046 (N_11046,N_8559,N_6881);
nor U11047 (N_11047,N_9290,N_5577);
nand U11048 (N_11048,N_6062,N_7750);
nor U11049 (N_11049,N_9880,N_9479);
and U11050 (N_11050,N_8476,N_7721);
and U11051 (N_11051,N_9679,N_6471);
xnor U11052 (N_11052,N_5776,N_9023);
nand U11053 (N_11053,N_5379,N_5004);
and U11054 (N_11054,N_8494,N_8781);
nor U11055 (N_11055,N_9423,N_8164);
or U11056 (N_11056,N_7142,N_7930);
nor U11057 (N_11057,N_8636,N_8000);
or U11058 (N_11058,N_7988,N_9309);
or U11059 (N_11059,N_8572,N_6641);
or U11060 (N_11060,N_8631,N_5943);
or U11061 (N_11061,N_6219,N_8895);
or U11062 (N_11062,N_8854,N_8357);
or U11063 (N_11063,N_9673,N_9522);
nor U11064 (N_11064,N_9248,N_9416);
nor U11065 (N_11065,N_6115,N_7986);
and U11066 (N_11066,N_9780,N_9519);
and U11067 (N_11067,N_6318,N_5559);
nand U11068 (N_11068,N_5212,N_6792);
nand U11069 (N_11069,N_5012,N_7020);
and U11070 (N_11070,N_8557,N_7531);
or U11071 (N_11071,N_5201,N_8725);
nand U11072 (N_11072,N_7906,N_8544);
nand U11073 (N_11073,N_9498,N_8880);
nand U11074 (N_11074,N_8925,N_9463);
and U11075 (N_11075,N_6769,N_5693);
and U11076 (N_11076,N_9353,N_5146);
nand U11077 (N_11077,N_7435,N_9104);
and U11078 (N_11078,N_9155,N_5352);
or U11079 (N_11079,N_8343,N_5286);
or U11080 (N_11080,N_7441,N_7334);
and U11081 (N_11081,N_6069,N_9552);
and U11082 (N_11082,N_9165,N_9148);
or U11083 (N_11083,N_6896,N_5707);
nor U11084 (N_11084,N_7512,N_9640);
nor U11085 (N_11085,N_9341,N_6432);
or U11086 (N_11086,N_8703,N_7234);
or U11087 (N_11087,N_7806,N_5472);
xor U11088 (N_11088,N_8024,N_5511);
or U11089 (N_11089,N_5120,N_6512);
and U11090 (N_11090,N_8058,N_8216);
nand U11091 (N_11091,N_7067,N_9768);
xor U11092 (N_11092,N_7772,N_8450);
nand U11093 (N_11093,N_9963,N_5361);
or U11094 (N_11094,N_7059,N_7677);
and U11095 (N_11095,N_7092,N_8262);
or U11096 (N_11096,N_5409,N_8334);
nand U11097 (N_11097,N_6308,N_8621);
nor U11098 (N_11098,N_9990,N_7275);
nor U11099 (N_11099,N_6184,N_5313);
and U11100 (N_11100,N_5962,N_7658);
nand U11101 (N_11101,N_9011,N_5760);
and U11102 (N_11102,N_7962,N_8549);
or U11103 (N_11103,N_7781,N_5613);
nand U11104 (N_11104,N_7485,N_7550);
nor U11105 (N_11105,N_7576,N_7344);
or U11106 (N_11106,N_5217,N_5522);
nor U11107 (N_11107,N_6066,N_7748);
and U11108 (N_11108,N_9972,N_9020);
and U11109 (N_11109,N_7818,N_7482);
xor U11110 (N_11110,N_6829,N_9725);
and U11111 (N_11111,N_9855,N_6802);
or U11112 (N_11112,N_7240,N_8731);
or U11113 (N_11113,N_7508,N_5722);
xnor U11114 (N_11114,N_6886,N_8542);
nand U11115 (N_11115,N_6466,N_6304);
or U11116 (N_11116,N_5453,N_6675);
nor U11117 (N_11117,N_9147,N_6889);
xnor U11118 (N_11118,N_6299,N_8025);
nor U11119 (N_11119,N_7788,N_7248);
and U11120 (N_11120,N_5706,N_9565);
xor U11121 (N_11121,N_6990,N_8906);
nor U11122 (N_11122,N_5842,N_8229);
nor U11123 (N_11123,N_9591,N_7188);
and U11124 (N_11124,N_6325,N_7850);
or U11125 (N_11125,N_9646,N_7915);
nand U11126 (N_11126,N_6545,N_8907);
nand U11127 (N_11127,N_7600,N_6696);
and U11128 (N_11128,N_7573,N_5597);
or U11129 (N_11129,N_6311,N_7894);
and U11130 (N_11130,N_7841,N_5935);
nand U11131 (N_11131,N_9219,N_9485);
or U11132 (N_11132,N_6706,N_6028);
nor U11133 (N_11133,N_7196,N_7808);
nand U11134 (N_11134,N_7197,N_9352);
and U11135 (N_11135,N_8974,N_6670);
or U11136 (N_11136,N_5205,N_5175);
and U11137 (N_11137,N_9292,N_9222);
and U11138 (N_11138,N_5024,N_7791);
and U11139 (N_11139,N_7280,N_6447);
nor U11140 (N_11140,N_8124,N_7377);
and U11141 (N_11141,N_9643,N_7610);
nand U11142 (N_11142,N_9388,N_8138);
and U11143 (N_11143,N_9090,N_6968);
and U11144 (N_11144,N_5153,N_8577);
or U11145 (N_11145,N_8341,N_9693);
and U11146 (N_11146,N_8683,N_9979);
or U11147 (N_11147,N_5986,N_6942);
nand U11148 (N_11148,N_9167,N_8205);
xnor U11149 (N_11149,N_6482,N_7224);
nor U11150 (N_11150,N_9506,N_5431);
xor U11151 (N_11151,N_6463,N_9705);
and U11152 (N_11152,N_8818,N_7515);
or U11153 (N_11153,N_6644,N_9810);
and U11154 (N_11154,N_9504,N_7030);
or U11155 (N_11155,N_7202,N_8642);
nor U11156 (N_11156,N_5557,N_8757);
nand U11157 (N_11157,N_8233,N_6531);
or U11158 (N_11158,N_5481,N_6353);
nand U11159 (N_11159,N_6077,N_6621);
nand U11160 (N_11160,N_8900,N_5768);
nor U11161 (N_11161,N_8770,N_9645);
or U11162 (N_11162,N_9787,N_5544);
nor U11163 (N_11163,N_7648,N_5101);
nand U11164 (N_11164,N_8105,N_6205);
and U11165 (N_11165,N_6610,N_9467);
nand U11166 (N_11166,N_9465,N_9205);
or U11167 (N_11167,N_6128,N_9544);
or U11168 (N_11168,N_9981,N_7396);
nand U11169 (N_11169,N_5757,N_5017);
nand U11170 (N_11170,N_6541,N_7063);
nand U11171 (N_11171,N_9723,N_5403);
and U11172 (N_11172,N_8090,N_9532);
or U11173 (N_11173,N_7651,N_6791);
nor U11174 (N_11174,N_8408,N_5025);
nor U11175 (N_11175,N_7857,N_5109);
and U11176 (N_11176,N_5071,N_8254);
and U11177 (N_11177,N_7382,N_8161);
nand U11178 (N_11178,N_8208,N_9774);
or U11179 (N_11179,N_5525,N_7179);
xor U11180 (N_11180,N_6564,N_5823);
nor U11181 (N_11181,N_9334,N_5469);
nor U11182 (N_11182,N_6832,N_9984);
nor U11183 (N_11183,N_8179,N_8785);
and U11184 (N_11184,N_9401,N_9752);
xor U11185 (N_11185,N_5275,N_5679);
and U11186 (N_11186,N_6510,N_5662);
xor U11187 (N_11187,N_6015,N_5880);
nand U11188 (N_11188,N_5138,N_8597);
nand U11189 (N_11189,N_8891,N_6533);
nand U11190 (N_11190,N_8135,N_8345);
xnor U11191 (N_11191,N_5214,N_8790);
or U11192 (N_11192,N_9460,N_7716);
nor U11193 (N_11193,N_6196,N_8608);
nand U11194 (N_11194,N_8432,N_7190);
and U11195 (N_11195,N_9249,N_7761);
and U11196 (N_11196,N_7633,N_6989);
nor U11197 (N_11197,N_8484,N_7569);
xor U11198 (N_11198,N_5758,N_7187);
nand U11199 (N_11199,N_7425,N_9151);
nand U11200 (N_11200,N_6252,N_9525);
xor U11201 (N_11201,N_8298,N_8063);
or U11202 (N_11202,N_6728,N_6622);
nor U11203 (N_11203,N_8066,N_5202);
or U11204 (N_11204,N_7612,N_8459);
nand U11205 (N_11205,N_7561,N_6398);
xor U11206 (N_11206,N_6950,N_9027);
or U11207 (N_11207,N_8534,N_9394);
and U11208 (N_11208,N_8152,N_7502);
and U11209 (N_11209,N_7752,N_9870);
and U11210 (N_11210,N_8338,N_7890);
nand U11211 (N_11211,N_5083,N_6386);
and U11212 (N_11212,N_5293,N_8162);
xor U11213 (N_11213,N_9936,N_5140);
nand U11214 (N_11214,N_7448,N_6048);
xnor U11215 (N_11215,N_6619,N_8689);
nand U11216 (N_11216,N_9331,N_9244);
and U11217 (N_11217,N_7175,N_7865);
and U11218 (N_11218,N_9577,N_5385);
nor U11219 (N_11219,N_6380,N_8400);
nor U11220 (N_11220,N_5981,N_9273);
nand U11221 (N_11221,N_6761,N_5952);
nand U11222 (N_11222,N_9597,N_6593);
or U11223 (N_11223,N_5717,N_7048);
nand U11224 (N_11224,N_9743,N_8740);
and U11225 (N_11225,N_8916,N_5422);
and U11226 (N_11226,N_5815,N_6272);
or U11227 (N_11227,N_9864,N_7632);
or U11228 (N_11228,N_8535,N_5304);
nor U11229 (N_11229,N_8797,N_6800);
and U11230 (N_11230,N_7295,N_8282);
and U11231 (N_11231,N_7756,N_9130);
xnor U11232 (N_11232,N_9016,N_9890);
or U11233 (N_11233,N_5974,N_5032);
and U11234 (N_11234,N_9888,N_8037);
xnor U11235 (N_11235,N_5503,N_8082);
or U11236 (N_11236,N_6026,N_8986);
or U11237 (N_11237,N_9373,N_6457);
nand U11238 (N_11238,N_5219,N_8756);
nor U11239 (N_11239,N_8438,N_6649);
nand U11240 (N_11240,N_5914,N_5897);
and U11241 (N_11241,N_9257,N_6838);
xnor U11242 (N_11242,N_7468,N_5569);
or U11243 (N_11243,N_6958,N_7866);
and U11244 (N_11244,N_8175,N_9912);
or U11245 (N_11245,N_6492,N_7649);
nand U11246 (N_11246,N_6448,N_7602);
nand U11247 (N_11247,N_5295,N_9176);
and U11248 (N_11248,N_5128,N_8892);
or U11249 (N_11249,N_8588,N_5517);
and U11250 (N_11250,N_8555,N_5964);
nand U11251 (N_11251,N_7080,N_7945);
and U11252 (N_11252,N_8990,N_8195);
nor U11253 (N_11253,N_6208,N_5442);
or U11254 (N_11254,N_9077,N_7774);
nand U11255 (N_11255,N_8997,N_5042);
or U11256 (N_11256,N_6236,N_9691);
nor U11257 (N_11257,N_8556,N_6760);
and U11258 (N_11258,N_5117,N_5963);
xor U11259 (N_11259,N_6345,N_8468);
nor U11260 (N_11260,N_5632,N_7215);
xor U11261 (N_11261,N_7010,N_6056);
or U11262 (N_11262,N_8469,N_8443);
nand U11263 (N_11263,N_6871,N_8730);
or U11264 (N_11264,N_7177,N_6460);
xor U11265 (N_11265,N_9391,N_6430);
nor U11266 (N_11266,N_8613,N_7918);
nand U11267 (N_11267,N_6974,N_6542);
nor U11268 (N_11268,N_7270,N_7427);
nand U11269 (N_11269,N_6454,N_7568);
or U11270 (N_11270,N_8697,N_8009);
or U11271 (N_11271,N_7384,N_5288);
nor U11272 (N_11272,N_8163,N_5141);
and U11273 (N_11273,N_9894,N_8273);
or U11274 (N_11274,N_7941,N_8656);
and U11275 (N_11275,N_8809,N_9399);
nand U11276 (N_11276,N_7209,N_6906);
nand U11277 (N_11277,N_9814,N_6291);
nor U11278 (N_11278,N_6354,N_6120);
or U11279 (N_11279,N_7091,N_6493);
or U11280 (N_11280,N_6509,N_5593);
or U11281 (N_11281,N_6280,N_5127);
nor U11282 (N_11282,N_8747,N_5636);
and U11283 (N_11283,N_8100,N_7003);
and U11284 (N_11284,N_6577,N_5795);
nand U11285 (N_11285,N_5484,N_6625);
xnor U11286 (N_11286,N_7783,N_6839);
or U11287 (N_11287,N_9626,N_5937);
nand U11288 (N_11288,N_6427,N_9907);
nand U11289 (N_11289,N_6513,N_9287);
nor U11290 (N_11290,N_5921,N_5835);
nor U11291 (N_11291,N_6558,N_9381);
nor U11292 (N_11292,N_7302,N_9197);
or U11293 (N_11293,N_9758,N_6651);
and U11294 (N_11294,N_6475,N_9923);
or U11295 (N_11295,N_8356,N_7046);
nand U11296 (N_11296,N_7287,N_7256);
nand U11297 (N_11297,N_9800,N_7198);
or U11298 (N_11298,N_6121,N_8196);
nor U11299 (N_11299,N_6032,N_6319);
and U11300 (N_11300,N_9857,N_8650);
or U11301 (N_11301,N_5150,N_8489);
nand U11302 (N_11302,N_9603,N_8537);
nor U11303 (N_11303,N_7836,N_6490);
xor U11304 (N_11304,N_5434,N_7228);
and U11305 (N_11305,N_9483,N_7370);
or U11306 (N_11306,N_8567,N_8054);
nand U11307 (N_11307,N_8325,N_5930);
nor U11308 (N_11308,N_5913,N_9744);
or U11309 (N_11309,N_9070,N_7174);
or U11310 (N_11310,N_9996,N_9424);
and U11311 (N_11311,N_6719,N_8768);
nor U11312 (N_11312,N_6963,N_7161);
or U11313 (N_11313,N_7892,N_8061);
nand U11314 (N_11314,N_7491,N_8005);
and U11315 (N_11315,N_7875,N_6446);
nor U11316 (N_11316,N_6699,N_6700);
or U11317 (N_11317,N_6982,N_8931);
and U11318 (N_11318,N_7002,N_6224);
xor U11319 (N_11319,N_9958,N_6771);
nand U11320 (N_11320,N_7722,N_6570);
nor U11321 (N_11321,N_6423,N_9821);
nor U11322 (N_11322,N_6166,N_6228);
xnor U11323 (N_11323,N_7944,N_9313);
nand U11324 (N_11324,N_7432,N_6724);
nand U11325 (N_11325,N_8976,N_5258);
and U11326 (N_11326,N_8668,N_7439);
nand U11327 (N_11327,N_5564,N_5248);
and U11328 (N_11328,N_5865,N_5475);
nand U11329 (N_11329,N_7961,N_7314);
nor U11330 (N_11330,N_6473,N_7084);
and U11331 (N_11331,N_6981,N_5589);
and U11332 (N_11332,N_8647,N_8139);
or U11333 (N_11333,N_8156,N_5640);
and U11334 (N_11334,N_6971,N_5535);
and U11335 (N_11335,N_6944,N_7631);
and U11336 (N_11336,N_9299,N_9150);
or U11337 (N_11337,N_5133,N_6819);
or U11338 (N_11338,N_6616,N_8610);
and U11339 (N_11339,N_6180,N_7497);
and U11340 (N_11340,N_7325,N_7565);
nor U11341 (N_11341,N_8964,N_5590);
nand U11342 (N_11342,N_7128,N_9125);
and U11343 (N_11343,N_6752,N_6902);
and U11344 (N_11344,N_9496,N_8049);
nand U11345 (N_11345,N_5084,N_8529);
nor U11346 (N_11346,N_8729,N_7773);
or U11347 (N_11347,N_7969,N_5946);
nand U11348 (N_11348,N_6167,N_6723);
or U11349 (N_11349,N_9271,N_6843);
nand U11350 (N_11350,N_9914,N_7426);
or U11351 (N_11351,N_9495,N_7719);
or U11352 (N_11352,N_6433,N_8598);
or U11353 (N_11353,N_5246,N_7758);
xor U11354 (N_11354,N_9132,N_9466);
xnor U11355 (N_11355,N_9889,N_9518);
nor U11356 (N_11356,N_9641,N_7012);
xor U11357 (N_11357,N_6680,N_6370);
nor U11358 (N_11358,N_6297,N_6663);
and U11359 (N_11359,N_5811,N_5166);
or U11360 (N_11360,N_5762,N_6088);
or U11361 (N_11361,N_7402,N_9614);
and U11362 (N_11362,N_6480,N_8394);
nor U11363 (N_11363,N_7102,N_9432);
nor U11364 (N_11364,N_9004,N_6231);
nor U11365 (N_11365,N_7897,N_7703);
or U11366 (N_11366,N_9234,N_7667);
nand U11367 (N_11367,N_9613,N_7904);
and U11368 (N_11368,N_9684,N_8970);
xnor U11369 (N_11369,N_6349,N_6708);
xor U11370 (N_11370,N_7327,N_8388);
nand U11371 (N_11371,N_7146,N_9076);
or U11372 (N_11372,N_6107,N_7754);
and U11373 (N_11373,N_5337,N_5213);
xor U11374 (N_11374,N_5948,N_8225);
nor U11375 (N_11375,N_5886,N_9531);
nand U11376 (N_11376,N_9511,N_5322);
nand U11377 (N_11377,N_8032,N_7946);
nor U11378 (N_11378,N_7253,N_8732);
or U11379 (N_11379,N_5334,N_6797);
or U11380 (N_11380,N_5879,N_9223);
and U11381 (N_11381,N_6727,N_5889);
nand U11382 (N_11382,N_7372,N_9380);
and U11383 (N_11383,N_9056,N_9778);
xor U11384 (N_11384,N_7358,N_8274);
or U11385 (N_11385,N_9702,N_5657);
nor U11386 (N_11386,N_7109,N_9811);
xnor U11387 (N_11387,N_8045,N_8787);
nand U11388 (N_11388,N_7409,N_5540);
xor U11389 (N_11389,N_5860,N_9179);
and U11390 (N_11390,N_5459,N_6900);
nor U11391 (N_11391,N_8857,N_8769);
nand U11392 (N_11392,N_8536,N_9566);
nand U11393 (N_11393,N_9724,N_7913);
nand U11394 (N_11394,N_7267,N_9058);
or U11395 (N_11395,N_8506,N_8590);
and U11396 (N_11396,N_8595,N_5990);
nor U11397 (N_11397,N_9540,N_5667);
or U11398 (N_11398,N_7124,N_7534);
and U11399 (N_11399,N_6507,N_7686);
or U11400 (N_11400,N_6959,N_8918);
or U11401 (N_11401,N_8012,N_9771);
nor U11402 (N_11402,N_7714,N_7025);
and U11403 (N_11403,N_5803,N_8966);
and U11404 (N_11404,N_7232,N_8269);
xor U11405 (N_11405,N_8182,N_8935);
nor U11406 (N_11406,N_9351,N_8578);
nand U11407 (N_11407,N_8570,N_5665);
or U11408 (N_11408,N_7040,N_5143);
nor U11409 (N_11409,N_7227,N_5942);
nor U11410 (N_11410,N_9924,N_8521);
nor U11411 (N_11411,N_9875,N_9948);
nor U11412 (N_11412,N_5845,N_9300);
or U11413 (N_11413,N_8853,N_6279);
nand U11414 (N_11414,N_5863,N_5694);
and U11415 (N_11415,N_9571,N_9697);
nor U11416 (N_11416,N_9717,N_8527);
nand U11417 (N_11417,N_5606,N_6469);
or U11418 (N_11418,N_6472,N_7099);
xor U11419 (N_11419,N_9696,N_9038);
or U11420 (N_11420,N_8873,N_8914);
nor U11421 (N_11421,N_9715,N_6187);
or U11422 (N_11422,N_9770,N_6784);
nand U11423 (N_11423,N_8284,N_7449);
nand U11424 (N_11424,N_8939,N_7119);
nand U11425 (N_11425,N_8799,N_5663);
and U11426 (N_11426,N_8574,N_9834);
nor U11427 (N_11427,N_8299,N_7332);
nand U11428 (N_11428,N_8428,N_5439);
or U11429 (N_11429,N_9390,N_6337);
nand U11430 (N_11430,N_7543,N_9478);
nand U11431 (N_11431,N_8967,N_6140);
or U11432 (N_11432,N_8416,N_8692);
nor U11433 (N_11433,N_7201,N_7823);
nor U11434 (N_11434,N_8675,N_6189);
and U11435 (N_11435,N_8286,N_7143);
nand U11436 (N_11436,N_6132,N_6289);
xnor U11437 (N_11437,N_7134,N_5005);
nor U11438 (N_11438,N_7058,N_6540);
nand U11439 (N_11439,N_6328,N_7182);
xnor U11440 (N_11440,N_8140,N_9840);
and U11441 (N_11441,N_5276,N_8142);
nand U11442 (N_11442,N_8217,N_5650);
or U11443 (N_11443,N_8856,N_7006);
and U11444 (N_11444,N_8881,N_5884);
or U11445 (N_11445,N_8571,N_9359);
xor U11446 (N_11446,N_5825,N_6477);
or U11447 (N_11447,N_5272,N_5477);
or U11448 (N_11448,N_5389,N_7471);
or U11449 (N_11449,N_7522,N_6817);
or U11450 (N_11450,N_5658,N_9699);
or U11451 (N_11451,N_5080,N_8463);
and U11452 (N_11452,N_7800,N_6376);
xnor U11453 (N_11453,N_7218,N_5635);
xor U11454 (N_11454,N_5649,N_9674);
xor U11455 (N_11455,N_5988,N_9258);
nor U11456 (N_11456,N_6440,N_6836);
and U11457 (N_11457,N_9529,N_9662);
or U11458 (N_11458,N_6378,N_9878);
nor U11459 (N_11459,N_9453,N_8664);
and U11460 (N_11460,N_9201,N_6916);
nor U11461 (N_11461,N_9280,N_9446);
and U11462 (N_11462,N_5314,N_8780);
nor U11463 (N_11463,N_7679,N_7567);
and U11464 (N_11464,N_5727,N_9546);
nand U11465 (N_11465,N_5374,N_7983);
and U11466 (N_11466,N_7586,N_5438);
and U11467 (N_11467,N_8944,N_8989);
nor U11468 (N_11468,N_7613,N_7043);
nor U11469 (N_11469,N_8788,N_5759);
or U11470 (N_11470,N_5841,N_6618);
and U11471 (N_11471,N_8579,N_7975);
or U11472 (N_11472,N_8928,N_6964);
xnor U11473 (N_11473,N_5923,N_5743);
nor U11474 (N_11474,N_8760,N_9074);
or U11475 (N_11475,N_8324,N_8480);
nand U11476 (N_11476,N_6652,N_9186);
nand U11477 (N_11477,N_8720,N_9319);
nor U11478 (N_11478,N_8249,N_9635);
xnor U11479 (N_11479,N_8539,N_8965);
nand U11480 (N_11480,N_6828,N_5770);
nand U11481 (N_11481,N_6500,N_6036);
nand U11482 (N_11482,N_8183,N_8192);
or U11483 (N_11483,N_5552,N_8104);
nor U11484 (N_11484,N_7027,N_8867);
nor U11485 (N_11485,N_5404,N_7081);
nor U11486 (N_11486,N_9920,N_8713);
nand U11487 (N_11487,N_9938,N_6922);
nand U11488 (N_11488,N_7588,N_6525);
nor U11489 (N_11489,N_9472,N_8943);
nor U11490 (N_11490,N_8372,N_5985);
nor U11491 (N_11491,N_8115,N_5030);
or U11492 (N_11492,N_7785,N_6160);
or U11493 (N_11493,N_9627,N_5222);
nor U11494 (N_11494,N_7952,N_9081);
nand U11495 (N_11495,N_8672,N_6005);
and U11496 (N_11496,N_8886,N_8087);
or U11497 (N_11497,N_5959,N_8295);
nor U11498 (N_11498,N_7147,N_6921);
or U11499 (N_11499,N_8762,N_5336);
xor U11500 (N_11500,N_7555,N_6009);
and U11501 (N_11501,N_6268,N_8776);
or U11502 (N_11502,N_8505,N_5184);
nand U11503 (N_11503,N_7645,N_8014);
nand U11504 (N_11504,N_5267,N_7365);
or U11505 (N_11505,N_6302,N_5624);
and U11506 (N_11506,N_7607,N_8252);
nor U11507 (N_11507,N_8387,N_5009);
or U11508 (N_11508,N_9123,N_7355);
or U11509 (N_11509,N_5619,N_8377);
or U11510 (N_11510,N_6213,N_6220);
and U11511 (N_11511,N_9808,N_5596);
nor U11512 (N_11512,N_5502,N_7079);
nor U11513 (N_11513,N_5271,N_6897);
xnor U11514 (N_11514,N_7578,N_5659);
or U11515 (N_11515,N_5623,N_9275);
and U11516 (N_11516,N_5901,N_5407);
nor U11517 (N_11517,N_5956,N_6517);
and U11518 (N_11518,N_7178,N_5902);
nand U11519 (N_11519,N_9791,N_6027);
nor U11520 (N_11520,N_8924,N_9899);
nand U11521 (N_11521,N_5232,N_7386);
and U11522 (N_11522,N_8277,N_6263);
nand U11523 (N_11523,N_5505,N_7963);
or U11524 (N_11524,N_8619,N_5898);
nor U11525 (N_11525,N_9886,N_6614);
xor U11526 (N_11526,N_8904,N_8065);
and U11527 (N_11527,N_7033,N_8452);
and U11528 (N_11528,N_7687,N_5019);
nand U11529 (N_11529,N_9736,N_5476);
and U11530 (N_11530,N_8688,N_7126);
and U11531 (N_11531,N_9619,N_6095);
and U11532 (N_11532,N_9749,N_5765);
nand U11533 (N_11533,N_6931,N_9761);
and U11534 (N_11534,N_7419,N_5016);
or U11535 (N_11535,N_5186,N_9083);
nand U11536 (N_11536,N_7429,N_9180);
and U11537 (N_11537,N_9748,N_7089);
nand U11538 (N_11538,N_5507,N_7417);
and U11539 (N_11539,N_9274,N_6478);
xnor U11540 (N_11540,N_7289,N_6514);
nor U11541 (N_11541,N_6826,N_9082);
nand U11542 (N_11542,N_5905,N_5060);
or U11543 (N_11543,N_8992,N_5044);
or U11544 (N_11544,N_7159,N_5402);
or U11545 (N_11545,N_5781,N_5750);
and U11546 (N_11546,N_6705,N_9668);
or U11547 (N_11547,N_6565,N_9324);
or U11548 (N_11548,N_9439,N_7031);
nor U11549 (N_11549,N_8741,N_6067);
nor U11550 (N_11550,N_8145,N_9704);
nor U11551 (N_11551,N_5711,N_5586);
nand U11552 (N_11552,N_5174,N_5440);
nor U11553 (N_11553,N_8491,N_7694);
xor U11554 (N_11554,N_5562,N_6218);
or U11555 (N_11555,N_6127,N_5467);
or U11556 (N_11556,N_5626,N_8863);
or U11557 (N_11557,N_6620,N_5225);
and U11558 (N_11558,N_8603,N_7405);
nand U11559 (N_11559,N_6736,N_9548);
or U11560 (N_11560,N_6266,N_5224);
or U11561 (N_11561,N_6711,N_5226);
nor U11562 (N_11562,N_8708,N_5620);
or U11563 (N_11563,N_7828,N_5779);
and U11564 (N_11564,N_8221,N_5139);
nor U11565 (N_11565,N_6254,N_5387);
nor U11566 (N_11566,N_7467,N_6589);
or U11567 (N_11567,N_5772,N_7393);
nor U11568 (N_11568,N_5056,N_8716);
or U11569 (N_11569,N_8512,N_8006);
xor U11570 (N_11570,N_6953,N_5850);
or U11571 (N_11571,N_6943,N_8328);
or U11572 (N_11572,N_7943,N_8399);
nand U11573 (N_11573,N_8187,N_6436);
nand U11574 (N_11574,N_8278,N_5001);
xnor U11575 (N_11575,N_7011,N_8260);
nand U11576 (N_11576,N_5412,N_9644);
nor U11577 (N_11577,N_5878,N_9196);
nand U11578 (N_11578,N_6580,N_6865);
nand U11579 (N_11579,N_9069,N_8763);
xnor U11580 (N_11580,N_5369,N_9312);
and U11581 (N_11581,N_8199,N_8367);
xor U11582 (N_11582,N_8174,N_8074);
or U11583 (N_11583,N_5927,N_6143);
nand U11584 (N_11584,N_6722,N_9731);
or U11585 (N_11585,N_6008,N_7004);
xnor U11586 (N_11586,N_8081,N_8059);
nand U11587 (N_11587,N_7135,N_6416);
nor U11588 (N_11588,N_6003,N_9343);
or U11589 (N_11589,N_6576,N_8874);
or U11590 (N_11590,N_6647,N_5773);
or U11591 (N_11591,N_5867,N_7440);
nor U11592 (N_11592,N_6276,N_8666);
xnor U11593 (N_11593,N_8794,N_5645);
nand U11594 (N_11594,N_5550,N_8810);
nor U11595 (N_11595,N_9554,N_7819);
and U11596 (N_11596,N_6743,N_9497);
or U11597 (N_11597,N_7611,N_6629);
nor U11598 (N_11598,N_6146,N_7803);
and U11599 (N_11599,N_9008,N_8052);
xnor U11600 (N_11600,N_9408,N_6234);
or U11601 (N_11601,N_7317,N_5539);
xnor U11602 (N_11602,N_6073,N_5473);
nand U11603 (N_11603,N_6818,N_9692);
nor U11604 (N_11604,N_5868,N_7414);
and U11605 (N_11605,N_9144,N_6898);
nor U11606 (N_11606,N_6417,N_5384);
nor U11607 (N_11607,N_7778,N_8479);
nand U11608 (N_11608,N_9874,N_5514);
nor U11609 (N_11609,N_9818,N_6860);
nor U11610 (N_11610,N_7933,N_9185);
nand U11611 (N_11611,N_5926,N_6991);
nand U11612 (N_11612,N_8302,N_9868);
nand U11613 (N_11613,N_6657,N_7484);
nand U11614 (N_11614,N_9118,N_9872);
nor U11615 (N_11615,N_5911,N_5549);
nand U11616 (N_11616,N_6547,N_6599);
or U11617 (N_11617,N_6317,N_8883);
and U11618 (N_11618,N_6894,N_5363);
nor U11619 (N_11619,N_9208,N_5067);
and U11620 (N_11620,N_5405,N_8193);
nor U11621 (N_11621,N_8600,N_5670);
nor U11622 (N_11622,N_5050,N_5487);
nand U11623 (N_11623,N_8878,N_7345);
and U11624 (N_11624,N_8279,N_5386);
nand U11625 (N_11625,N_8850,N_9241);
or U11626 (N_11626,N_5691,N_8336);
and U11627 (N_11627,N_5728,N_8568);
and U11628 (N_11628,N_6277,N_8497);
and U11629 (N_11629,N_8870,N_6165);
nor U11630 (N_11630,N_7167,N_8444);
nor U11631 (N_11631,N_6295,N_5448);
and U11632 (N_11632,N_7387,N_8446);
and U11633 (N_11633,N_5112,N_7139);
and U11634 (N_11634,N_5390,N_6965);
or U11635 (N_11635,N_7577,N_7775);
and U11636 (N_11636,N_6607,N_7905);
nand U11637 (N_11637,N_5310,N_9760);
or U11638 (N_11638,N_8582,N_6751);
nand U11639 (N_11639,N_9230,N_9911);
nand U11640 (N_11640,N_5287,N_8375);
and U11641 (N_11641,N_7008,N_8200);
and U11642 (N_11642,N_5333,N_6257);
nand U11643 (N_11643,N_6820,N_7403);
and U11644 (N_11644,N_5318,N_6373);
nand U11645 (N_11645,N_6567,N_9562);
and U11646 (N_11646,N_9517,N_6227);
or U11647 (N_11647,N_8294,N_9595);
nand U11648 (N_11648,N_6488,N_6594);
nor U11649 (N_11649,N_6405,N_8434);
nor U11650 (N_11650,N_8957,N_9235);
or U11651 (N_11651,N_6691,N_6850);
and U11652 (N_11652,N_9999,N_6426);
nand U11653 (N_11653,N_7730,N_6320);
or U11654 (N_11654,N_6948,N_8113);
or U11655 (N_11655,N_5328,N_9240);
nor U11656 (N_11656,N_9296,N_5207);
nand U11657 (N_11657,N_9510,N_6258);
xnor U11658 (N_11658,N_6075,N_9387);
nand U11659 (N_11659,N_5581,N_7194);
and U11660 (N_11660,N_7347,N_6049);
or U11661 (N_11661,N_9374,N_7554);
or U11662 (N_11662,N_6929,N_6933);
and U11663 (N_11663,N_9194,N_7979);
xor U11664 (N_11664,N_7673,N_7359);
xor U11665 (N_11665,N_7674,N_8541);
nor U11666 (N_11666,N_9949,N_6613);
nor U11667 (N_11667,N_7728,N_9790);
and U11668 (N_11668,N_5468,N_5209);
nand U11669 (N_11669,N_9206,N_5026);
and U11670 (N_11670,N_9873,N_7250);
and U11671 (N_11671,N_8234,N_9973);
nor U11672 (N_11672,N_9530,N_5814);
nand U11673 (N_11673,N_6588,N_7231);
nor U11674 (N_11674,N_6403,N_6867);
nor U11675 (N_11675,N_6997,N_8110);
nor U11676 (N_11676,N_5994,N_9906);
xnor U11677 (N_11677,N_5102,N_8150);
or U11678 (N_11678,N_9032,N_7500);
xnor U11679 (N_11679,N_9882,N_5713);
and U11680 (N_11680,N_7957,N_8848);
or U11681 (N_11681,N_7855,N_7260);
nand U11682 (N_11682,N_7626,N_7320);
or U11683 (N_11683,N_7615,N_5669);
nand U11684 (N_11684,N_9853,N_5059);
nand U11685 (N_11685,N_5455,N_5763);
and U11686 (N_11686,N_8832,N_7406);
and U11687 (N_11687,N_8959,N_6368);
xor U11688 (N_11688,N_6939,N_5592);
nand U11689 (N_11689,N_9447,N_8554);
and U11690 (N_11690,N_7312,N_8767);
xnor U11691 (N_11691,N_6571,N_8340);
nor U11692 (N_11692,N_8802,N_8226);
and U11693 (N_11693,N_6932,N_7978);
nor U11694 (N_11694,N_7964,N_6806);
nand U11695 (N_11695,N_6785,N_6081);
nor U11696 (N_11696,N_7977,N_8660);
and U11697 (N_11697,N_7542,N_7907);
or U11698 (N_11698,N_7352,N_8958);
and U11699 (N_11699,N_8270,N_6361);
xor U11700 (N_11700,N_7001,N_8157);
or U11701 (N_11701,N_5684,N_6837);
nor U11702 (N_11702,N_7516,N_5521);
nand U11703 (N_11703,N_7241,N_7591);
nor U11704 (N_11704,N_9983,N_5114);
or U11705 (N_11705,N_8507,N_5574);
and U11706 (N_11706,N_8240,N_7794);
nor U11707 (N_11707,N_7556,N_9722);
nor U11708 (N_11708,N_6177,N_7603);
nand U11709 (N_11709,N_8626,N_5893);
and U11710 (N_11710,N_8607,N_8817);
or U11711 (N_11711,N_7291,N_8784);
or U11712 (N_11712,N_8980,N_9826);
and U11713 (N_11713,N_8411,N_7608);
or U11714 (N_11714,N_9404,N_6669);
or U11715 (N_11715,N_8292,N_8615);
or U11716 (N_11716,N_8159,N_9992);
or U11717 (N_11717,N_7150,N_8276);
nand U11718 (N_11718,N_7751,N_5644);
nor U11719 (N_11719,N_5603,N_8789);
nand U11720 (N_11720,N_8064,N_5277);
and U11721 (N_11721,N_6986,N_7564);
nand U11722 (N_11722,N_9455,N_5890);
and U11723 (N_11723,N_8405,N_9110);
or U11724 (N_11724,N_5551,N_9634);
or U11725 (N_11725,N_7690,N_9026);
or U11726 (N_11726,N_6983,N_8203);
xnor U11727 (N_11727,N_7138,N_7715);
nand U11728 (N_11728,N_5326,N_8686);
nor U11729 (N_11729,N_6462,N_9013);
xor U11730 (N_11730,N_5266,N_9820);
or U11731 (N_11731,N_7029,N_9727);
and U11732 (N_11732,N_7764,N_5526);
xnor U11733 (N_11733,N_7968,N_8748);
or U11734 (N_11734,N_7447,N_5497);
and U11735 (N_11735,N_7539,N_8806);
and U11736 (N_11736,N_7741,N_5726);
nor U11737 (N_11737,N_7982,N_9107);
xor U11738 (N_11738,N_7814,N_9989);
nor U11739 (N_11739,N_8385,N_6223);
nor U11740 (N_11740,N_8131,N_8250);
nor U11741 (N_11741,N_5037,N_8930);
nand U11742 (N_11742,N_7163,N_7637);
or U11743 (N_11743,N_8481,N_8088);
nand U11744 (N_11744,N_8868,N_6415);
or U11745 (N_11745,N_6770,N_7924);
or U11746 (N_11746,N_5881,N_8951);
and U11747 (N_11747,N_7925,N_7465);
and U11748 (N_11748,N_9141,N_5358);
nor U11749 (N_11749,N_5998,N_7670);
nand U11750 (N_11750,N_7922,N_8289);
nand U11751 (N_11751,N_9036,N_5257);
nor U11752 (N_11752,N_9505,N_9630);
nand U11753 (N_11753,N_6467,N_8147);
xnor U11754 (N_11754,N_9563,N_8910);
nand U11755 (N_11755,N_7252,N_7460);
and U11756 (N_11756,N_9664,N_8309);
nor U11757 (N_11757,N_7938,N_5416);
or U11758 (N_11758,N_8901,N_7553);
and U11759 (N_11759,N_5656,N_7732);
nor U11760 (N_11760,N_5230,N_5583);
or U11761 (N_11761,N_5302,N_8651);
nor U11762 (N_11762,N_7529,N_5149);
or U11763 (N_11763,N_9225,N_7064);
and U11764 (N_11764,N_9835,N_6750);
and U11765 (N_11765,N_8475,N_7697);
and U11766 (N_11766,N_6759,N_5812);
nor U11767 (N_11767,N_9654,N_9086);
nand U11768 (N_11768,N_8383,N_7407);
nand U11769 (N_11769,N_7255,N_6508);
nand U11770 (N_11770,N_7461,N_9930);
or U11771 (N_11771,N_6094,N_5366);
nand U11772 (N_11772,N_9405,N_8954);
xor U11773 (N_11773,N_9738,N_9671);
nand U11774 (N_11774,N_7378,N_7028);
nor U11775 (N_11775,N_7624,N_5542);
or U11776 (N_11776,N_6375,N_5695);
and U11777 (N_11777,N_8698,N_8894);
and U11778 (N_11778,N_9255,N_7639);
xor U11779 (N_11779,N_9655,N_9993);
and U11780 (N_11780,N_8319,N_9154);
nand U11781 (N_11781,N_7181,N_8130);
nor U11782 (N_11782,N_5975,N_9688);
xor U11783 (N_11783,N_6562,N_5451);
or U11784 (N_11784,N_6025,N_5493);
or U11785 (N_11785,N_9282,N_6559);
nand U11786 (N_11786,N_9349,N_5529);
xor U11787 (N_11787,N_5263,N_7876);
and U11788 (N_11788,N_7736,N_6409);
xor U11789 (N_11789,N_7308,N_6147);
and U11790 (N_11790,N_5553,N_7530);
or U11791 (N_11791,N_5068,N_5450);
nand U11792 (N_11792,N_7706,N_5085);
xor U11793 (N_11793,N_8173,N_7103);
or U11794 (N_11794,N_8143,N_8798);
and U11795 (N_11795,N_9547,N_8111);
nand U11796 (N_11796,N_5375,N_7362);
nor U11797 (N_11797,N_9714,N_7153);
nand U11798 (N_11798,N_8807,N_8596);
xor U11799 (N_11799,N_5460,N_6479);
nand U11800 (N_11800,N_9172,N_9881);
and U11801 (N_11801,N_7503,N_9035);
nor U11802 (N_11802,N_7829,N_7457);
or U11803 (N_11803,N_7729,N_7107);
and U11804 (N_11804,N_8839,N_5573);
nor U11805 (N_11805,N_7235,N_9400);
or U11806 (N_11806,N_9599,N_8814);
xor U11807 (N_11807,N_7505,N_6910);
nor U11808 (N_11808,N_6449,N_9493);
nor U11809 (N_11809,N_8573,N_7353);
nor U11810 (N_11810,N_8811,N_9754);
nor U11811 (N_11811,N_7214,N_6741);
and U11812 (N_11812,N_8181,N_9666);
nor U11813 (N_11813,N_9421,N_5113);
or U11814 (N_11814,N_7140,N_6089);
or U11815 (N_11815,N_7469,N_7592);
xor U11816 (N_11816,N_9559,N_6011);
or U11817 (N_11817,N_9891,N_8409);
xor U11818 (N_11818,N_5078,N_5643);
and U11819 (N_11819,N_9105,N_5297);
nand U11820 (N_11820,N_6285,N_6835);
xnor U11821 (N_11821,N_6262,N_9162);
and U11822 (N_11822,N_8017,N_7168);
or U11823 (N_11823,N_7041,N_9841);
or U11824 (N_11824,N_7852,N_8849);
and U11825 (N_11825,N_7994,N_9226);
and U11826 (N_11826,N_9807,N_9318);
xor U11827 (N_11827,N_5456,N_5501);
or U11828 (N_11828,N_6351,N_9551);
nor U11829 (N_11829,N_6575,N_9191);
or U11830 (N_11830,N_6338,N_8318);
or U11831 (N_11831,N_6775,N_8937);
and U11832 (N_11832,N_8687,N_8715);
nand U11833 (N_11833,N_8401,N_6451);
xor U11834 (N_11834,N_9175,N_7793);
nand U11835 (N_11835,N_7271,N_7264);
nor U11836 (N_11836,N_9228,N_9940);
nand U11837 (N_11837,N_5058,N_5611);
nand U11838 (N_11838,N_5778,N_8584);
or U11839 (N_11839,N_8168,N_7513);
nor U11840 (N_11840,N_5683,N_7950);
and U11841 (N_11841,N_5744,N_6346);
or U11842 (N_11842,N_7863,N_9019);
nand U11843 (N_11843,N_6369,N_9364);
nand U11844 (N_11844,N_7813,N_6919);
or U11845 (N_11845,N_7210,N_5261);
nor U11846 (N_11846,N_8332,N_5239);
nor U11847 (N_11847,N_6442,N_9934);
xor U11848 (N_11848,N_5305,N_6918);
xnor U11849 (N_11849,N_6666,N_9209);
and U11850 (N_11850,N_6159,N_6729);
and U11851 (N_11851,N_9099,N_5996);
nand U11852 (N_11852,N_5939,N_9721);
and U11853 (N_11853,N_5498,N_6831);
xor U11854 (N_11854,N_9543,N_6955);
and U11855 (N_11855,N_5221,N_8473);
xor U11856 (N_11856,N_7480,N_7984);
xor U11857 (N_11857,N_5391,N_7121);
and U11858 (N_11858,N_7638,N_9765);
or U11859 (N_11859,N_7410,N_5430);
nand U11860 (N_11860,N_7991,N_7122);
and U11861 (N_11861,N_5176,N_9094);
xnor U11862 (N_11862,N_9049,N_7039);
and U11863 (N_11863,N_6171,N_9968);
nor U11864 (N_11864,N_8599,N_5168);
or U11865 (N_11865,N_7223,N_8525);
and U11866 (N_11866,N_9707,N_8102);
or U11867 (N_11867,N_9954,N_9103);
and U11868 (N_11868,N_5341,N_6530);
nand U11869 (N_11869,N_9726,N_5532);
xnor U11870 (N_11870,N_6333,N_8040);
nand U11871 (N_11871,N_6793,N_5396);
nand U11872 (N_11872,N_9734,N_6901);
and U11873 (N_11873,N_9322,N_9028);
nand U11874 (N_11874,N_5675,N_7458);
nor U11875 (N_11875,N_5435,N_5096);
or U11876 (N_11876,N_5049,N_7333);
and U11877 (N_11877,N_9289,N_6967);
nand U11878 (N_11878,N_8926,N_8833);
and U11879 (N_11879,N_7622,N_8373);
nand U11880 (N_11880,N_7858,N_9997);
nor U11881 (N_11881,N_5317,N_7849);
nand U11882 (N_11882,N_8490,N_5924);
or U11883 (N_11883,N_5951,N_5132);
or U11884 (N_11884,N_6161,N_5125);
nor U11885 (N_11885,N_9403,N_6068);
or U11886 (N_11886,N_6701,N_7997);
or U11887 (N_11887,N_8281,N_7678);
nor U11888 (N_11888,N_8048,N_5729);
and U11889 (N_11889,N_9006,N_7399);
or U11890 (N_11890,N_7203,N_6483);
xor U11891 (N_11891,N_5104,N_5510);
or U11892 (N_11892,N_6744,N_5041);
nand U11893 (N_11893,N_7035,N_9728);
nor U11894 (N_11894,N_5714,N_8125);
nand U11895 (N_11895,N_6885,N_6379);
and U11896 (N_11896,N_7037,N_8210);
nor U11897 (N_11897,N_5903,N_5724);
or U11898 (N_11898,N_5855,N_9813);
xor U11899 (N_11899,N_9071,N_6203);
and U11900 (N_11900,N_6637,N_6809);
xnor U11901 (N_11901,N_6192,N_8447);
nor U11902 (N_11902,N_6572,N_8637);
nor U11903 (N_11903,N_5704,N_6822);
nor U11904 (N_11904,N_6211,N_8877);
and U11905 (N_11905,N_9801,N_6396);
nand U11906 (N_11906,N_7826,N_9925);
or U11907 (N_11907,N_5461,N_7418);
and U11908 (N_11908,N_5471,N_7601);
or U11909 (N_11909,N_9629,N_9149);
and U11910 (N_11910,N_8251,N_5180);
and U11911 (N_11911,N_6024,N_8106);
nor U11912 (N_11912,N_6861,N_6851);
xnor U11913 (N_11913,N_7339,N_7474);
and U11914 (N_11914,N_6407,N_7710);
and U11915 (N_11915,N_6267,N_6072);
nand U11916 (N_11916,N_5197,N_7784);
or U11917 (N_11917,N_5628,N_8978);
and U11918 (N_11918,N_7641,N_9124);
nand U11919 (N_11919,N_8616,N_7366);
nand U11920 (N_11920,N_7391,N_9509);
xor U11921 (N_11921,N_7268,N_8606);
or U11922 (N_11922,N_8347,N_5518);
and U11923 (N_11923,N_9128,N_5917);
nor U11924 (N_11924,N_7998,N_6083);
or U11925 (N_11925,N_5874,N_6528);
nand U11926 (N_11926,N_6029,N_6214);
nor U11927 (N_11927,N_7104,N_6076);
or U11928 (N_11928,N_9066,N_8653);
nand U11929 (N_11929,N_6330,N_6882);
nor U11930 (N_11930,N_9265,N_7019);
and U11931 (N_11931,N_6988,N_9428);
and U11932 (N_11932,N_8176,N_8820);
nor U11933 (N_11933,N_6350,N_9471);
or U11934 (N_11934,N_7315,N_6152);
and U11935 (N_11935,N_5413,N_9915);
nor U11936 (N_11936,N_5652,N_8812);
and U11937 (N_11937,N_6444,N_9080);
nor U11938 (N_11938,N_9188,N_7526);
xnor U11939 (N_11939,N_8706,N_7666);
and U11940 (N_11940,N_7483,N_8453);
or U11941 (N_11941,N_8402,N_6642);
nand U11942 (N_11942,N_8585,N_7413);
or U11943 (N_11943,N_5982,N_8882);
xnor U11944 (N_11944,N_5752,N_7110);
and U11945 (N_11945,N_9564,N_6045);
or U11946 (N_11946,N_5866,N_5541);
nor U11947 (N_11947,N_7867,N_6402);
and U11948 (N_11948,N_8821,N_9602);
xnor U11949 (N_11949,N_7899,N_5678);
nor U11950 (N_11950,N_6489,N_9178);
nand U11951 (N_11951,N_5534,N_6788);
or U11952 (N_11952,N_7527,N_8612);
nor U11953 (N_11953,N_5000,N_7967);
nor U11954 (N_11954,N_5081,N_9192);
nor U11955 (N_11955,N_7069,N_7928);
xor U11956 (N_11956,N_7171,N_8354);
nand U11957 (N_11957,N_6543,N_5800);
xor U11958 (N_11958,N_7501,N_7076);
or U11959 (N_11959,N_9409,N_6841);
nand U11960 (N_11960,N_6624,N_8188);
nand U11961 (N_11961,N_6903,N_6294);
or U11962 (N_11962,N_5281,N_5836);
nand U11963 (N_11963,N_8283,N_9084);
or U11964 (N_11964,N_7523,N_9159);
nand U11965 (N_11965,N_7294,N_6623);
or U11966 (N_11966,N_8155,N_7380);
and U11967 (N_11967,N_5259,N_6078);
nand U11968 (N_11968,N_8304,N_7580);
nand U11969 (N_11969,N_5580,N_7958);
and U11970 (N_11970,N_6491,N_5095);
nand U11971 (N_11971,N_6157,N_6890);
or U11972 (N_11972,N_8674,N_7282);
xnor U11973 (N_11973,N_7936,N_7328);
and U11974 (N_11974,N_8511,N_7659);
nor U11975 (N_11975,N_9541,N_9325);
xor U11976 (N_11976,N_7281,N_7321);
xnor U11977 (N_11977,N_9850,N_7927);
nand U11978 (N_11978,N_5269,N_7853);
or U11979 (N_11979,N_9345,N_8993);
nor U11980 (N_11980,N_9788,N_9919);
nand U11981 (N_11981,N_9117,N_9459);
nand U11982 (N_11982,N_8589,N_7156);
nand U11983 (N_11983,N_5688,N_6485);
or U11984 (N_11984,N_8275,N_5703);
nor U11985 (N_11985,N_5805,N_7627);
and U11986 (N_11986,N_7885,N_6852);
xnor U11987 (N_11987,N_8034,N_6395);
and U11988 (N_11988,N_5376,N_9385);
and U11989 (N_11989,N_5794,N_6546);
nor U11990 (N_11990,N_9429,N_6038);
or U11991 (N_11991,N_6672,N_9756);
nand U11992 (N_11992,N_5506,N_6755);
or U11993 (N_11993,N_6938,N_5028);
or U11994 (N_11994,N_5607,N_8890);
and U11995 (N_11995,N_8658,N_7759);
and U11996 (N_11996,N_9243,N_8946);
nand U11997 (N_11997,N_8609,N_9184);
or U11998 (N_11998,N_6002,N_9195);
or U11999 (N_11999,N_7455,N_6961);
xnor U12000 (N_12000,N_9078,N_7989);
and U12001 (N_12001,N_5365,N_8773);
or U12002 (N_12002,N_7949,N_9903);
and U12003 (N_12003,N_6242,N_5255);
nor U12004 (N_12004,N_6946,N_9883);
nand U12005 (N_12005,N_9311,N_6601);
and U12006 (N_12006,N_6251,N_8190);
or U12007 (N_12007,N_9482,N_9156);
nor U12008 (N_12008,N_5646,N_8774);
nor U12009 (N_12009,N_8919,N_8442);
or U12010 (N_12010,N_6639,N_8293);
and U12011 (N_12011,N_7338,N_7795);
nor U12012 (N_12012,N_6879,N_5857);
nand U12013 (N_12013,N_7792,N_5070);
nand U12014 (N_12014,N_7617,N_5537);
nor U12015 (N_12015,N_5895,N_9481);
nand U12016 (N_12016,N_7996,N_5447);
nand U12017 (N_12017,N_8067,N_6632);
nor U12018 (N_12018,N_7840,N_6342);
or U12019 (N_12019,N_8346,N_9832);
xnor U12020 (N_12020,N_9660,N_9488);
nor U12021 (N_12021,N_9978,N_6181);
and U12022 (N_12022,N_7737,N_7170);
nor U12023 (N_12023,N_6726,N_5029);
or U12024 (N_12024,N_6520,N_7727);
or U12025 (N_12025,N_5582,N_9687);
nand U12026 (N_12026,N_6103,N_6357);
xor U12027 (N_12027,N_7155,N_6909);
or U12028 (N_12028,N_8831,N_6134);
nor U12029 (N_12029,N_6764,N_9521);
or U12030 (N_12030,N_9033,N_7157);
nor U12031 (N_12031,N_9611,N_9561);
nor U12032 (N_12032,N_9932,N_7306);
nor U12033 (N_12033,N_7272,N_6880);
nand U12034 (N_12034,N_8562,N_6019);
nand U12035 (N_12035,N_9199,N_9304);
nand U12036 (N_12036,N_9412,N_8879);
nand U12037 (N_12037,N_7265,N_6683);
xnor U12038 (N_12038,N_7086,N_7824);
xnor U12039 (N_12039,N_6807,N_8678);
nand U12040 (N_12040,N_9163,N_5163);
or U12041 (N_12041,N_6464,N_7560);
and U12042 (N_12042,N_8933,N_8670);
or U12043 (N_12043,N_8013,N_7574);
nor U12044 (N_12044,N_7757,N_9417);
xnor U12045 (N_12045,N_7343,N_8238);
nand U12046 (N_12046,N_9823,N_8903);
nor U12047 (N_12047,N_7233,N_9753);
or U12048 (N_12048,N_9030,N_7094);
nor U12049 (N_12049,N_8441,N_8540);
nor U12050 (N_12050,N_5124,N_8019);
nor U12051 (N_12051,N_6695,N_9366);
or U12052 (N_12052,N_8384,N_8865);
nand U12053 (N_12053,N_8548,N_7100);
nand U12054 (N_12054,N_6825,N_5718);
nand U12055 (N_12055,N_8956,N_7859);
nand U12056 (N_12056,N_6309,N_8804);
and U12057 (N_12057,N_5600,N_9683);
xor U12058 (N_12058,N_9376,N_6465);
or U12059 (N_12059,N_8823,N_5103);
or U12060 (N_12060,N_5872,N_9001);
xnor U12061 (N_12061,N_8921,N_5137);
nand U12062 (N_12062,N_7599,N_6060);
or U12063 (N_12063,N_5968,N_9073);
nand U12064 (N_12064,N_6452,N_8898);
nand U12065 (N_12065,N_9856,N_9617);
or U12066 (N_12066,N_8526,N_8984);
or U12067 (N_12067,N_9784,N_7864);
nand U12068 (N_12068,N_8018,N_6833);
and U12069 (N_12069,N_8952,N_8962);
nor U12070 (N_12070,N_9342,N_7061);
nor U12071 (N_12071,N_6079,N_8661);
and U12072 (N_12072,N_6290,N_6544);
nand U12073 (N_12073,N_8093,N_5064);
nor U12074 (N_12074,N_6805,N_6934);
or U12075 (N_12075,N_8312,N_9686);
or U12076 (N_12076,N_6720,N_7279);
and U12077 (N_12077,N_5837,N_5630);
xnor U12078 (N_12078,N_6256,N_7654);
or U12079 (N_12079,N_9794,N_5883);
nand U12080 (N_12080,N_5136,N_9601);
nor U12081 (N_12081,N_6216,N_5010);
xnor U12082 (N_12082,N_5087,N_7689);
nor U12083 (N_12083,N_6538,N_8772);
and U12084 (N_12084,N_9703,N_8170);
nand U12085 (N_12085,N_7579,N_8386);
nand U12086 (N_12086,N_8513,N_5602);
nand U12087 (N_12087,N_8829,N_6260);
and U12088 (N_12088,N_8669,N_6505);
nand U12089 (N_12089,N_9537,N_9126);
and U12090 (N_12090,N_9622,N_7551);
nor U12091 (N_12091,N_8047,N_6149);
or U12092 (N_12092,N_7533,N_7229);
and U12093 (N_12093,N_8167,N_7839);
nand U12094 (N_12094,N_8207,N_7815);
or U12095 (N_12095,N_6534,N_9210);
and U12096 (N_12096,N_6052,N_5321);
nor U12097 (N_12097,N_6226,N_5482);
xor U12098 (N_12098,N_8520,N_5192);
and U12099 (N_12099,N_6372,N_9759);
and U12100 (N_12100,N_8667,N_9740);
or U12101 (N_12101,N_6522,N_7136);
xor U12102 (N_12102,N_8710,N_9609);
or U12103 (N_12103,N_8532,N_9193);
nor U12104 (N_12104,N_8922,N_5159);
and U12105 (N_12105,N_5110,N_8714);
and U12106 (N_12106,N_9842,N_7318);
nand U12107 (N_12107,N_7972,N_7753);
and U12108 (N_12108,N_5961,N_7158);
nor U12109 (N_12109,N_6194,N_7874);
or U12110 (N_12110,N_6668,N_7766);
or U12111 (N_12111,N_8151,N_5188);
or U12112 (N_12112,N_7462,N_5167);
and U12113 (N_12113,N_5709,N_7882);
or U12114 (N_12114,N_9694,N_8177);
nand U12115 (N_12115,N_9592,N_7845);
nand U12116 (N_12116,N_9575,N_5483);
or U12117 (N_12117,N_6627,N_9642);
nand U12118 (N_12118,N_7683,N_5900);
or U12119 (N_12119,N_7871,N_9960);
nor U12120 (N_12120,N_8721,N_8861);
nand U12121 (N_12121,N_7745,N_8885);
and U12122 (N_12122,N_8015,N_5378);
nor U12123 (N_12123,N_8412,N_8941);
nand U12124 (N_12124,N_9435,N_8454);
nand U12125 (N_12125,N_8622,N_5424);
and U12126 (N_12126,N_9121,N_5097);
nor U12127 (N_12127,N_7376,N_6969);
or U12128 (N_12128,N_9310,N_8929);
and U12129 (N_12129,N_9909,N_6927);
nor U12130 (N_12130,N_8905,N_7088);
xor U12131 (N_12131,N_6178,N_6772);
or U12132 (N_12132,N_8761,N_8362);
nand U12133 (N_12133,N_6155,N_7931);
nand U12134 (N_12134,N_9512,N_6148);
and U12135 (N_12135,N_8352,N_6106);
nand U12136 (N_12136,N_8011,N_5734);
and U12137 (N_12137,N_9021,N_9079);
and U12138 (N_12138,N_9386,N_9623);
or U12139 (N_12139,N_6842,N_7696);
nor U12140 (N_12140,N_9854,N_9698);
or U12141 (N_12141,N_7340,N_6730);
and U12142 (N_12142,N_6568,N_6721);
nand U12143 (N_12143,N_9876,N_8845);
nand U12144 (N_12144,N_5690,N_6390);
nor U12145 (N_12145,N_7934,N_9236);
or U12146 (N_12146,N_9484,N_9776);
or U12147 (N_12147,N_9959,N_6183);
nand U12148 (N_12148,N_9002,N_7298);
nor U12149 (N_12149,N_6634,N_8296);
or U12150 (N_12150,N_5916,N_5162);
or U12151 (N_12151,N_8803,N_6182);
nand U12152 (N_12152,N_6812,N_7036);
nor U12153 (N_12153,N_9111,N_5595);
nand U12154 (N_12154,N_9116,N_9378);
or U12155 (N_12155,N_6247,N_5712);
or U12156 (N_12156,N_7101,N_5767);
xor U12157 (N_12157,N_7165,N_6795);
and U12158 (N_12158,N_8267,N_8866);
or U12159 (N_12159,N_9618,N_8158);
or U12160 (N_12160,N_9847,N_7914);
nand U12161 (N_12161,N_9502,N_7398);
and U12162 (N_12162,N_6762,N_8640);
nand U12163 (N_12163,N_9742,N_8410);
nand U12164 (N_12164,N_9710,N_7548);
xnor U12165 (N_12165,N_7628,N_5357);
xor U12166 (N_12166,N_6315,N_8211);
and U12167 (N_12167,N_9040,N_6097);
and U12168 (N_12168,N_7056,N_5052);
xnor U12169 (N_12169,N_6516,N_9576);
or U12170 (N_12170,N_6707,N_9131);
and U12171 (N_12171,N_5429,N_8371);
nor U12172 (N_12172,N_7204,N_8602);
or U12173 (N_12173,N_5349,N_6970);
nor U12174 (N_12174,N_6773,N_8888);
xor U12175 (N_12175,N_6643,N_5830);
and U12176 (N_12176,N_5306,N_8948);
xor U12177 (N_12177,N_5869,N_8819);
nand U12178 (N_12178,N_7532,N_6071);
or U12179 (N_12179,N_8496,N_7956);
xnor U12180 (N_12180,N_6848,N_6704);
or U12181 (N_12181,N_8528,N_8077);
or U12182 (N_12182,N_7357,N_6200);
nor U12183 (N_12183,N_9474,N_6314);
or U12184 (N_12184,N_7324,N_7985);
nand U12185 (N_12185,N_6414,N_8184);
nor U12186 (N_12186,N_8641,N_9229);
or U12187 (N_12187,N_5076,N_5862);
nor U12188 (N_12188,N_7990,N_9348);
or U12189 (N_12189,N_6694,N_6774);
or U12190 (N_12190,N_9785,N_7755);
nor U12191 (N_12191,N_5977,N_9836);
nand U12192 (N_12192,N_9379,N_9170);
nor U12193 (N_12193,N_9087,N_5618);
nand U12194 (N_12194,N_8518,N_5938);
nor U12195 (N_12195,N_8969,N_9830);
nor U12196 (N_12196,N_8680,N_8999);
nand U12197 (N_12197,N_8440,N_7742);
nand U12198 (N_12198,N_5877,N_5806);
nor U12199 (N_12199,N_9558,N_5411);
nand U12200 (N_12200,N_9098,N_5215);
nor U12201 (N_12201,N_8837,N_7239);
nand U12202 (N_12202,N_6899,N_9860);
nand U12203 (N_12203,N_9267,N_7827);
or U12204 (N_12204,N_7799,N_5906);
and U12205 (N_12205,N_7416,N_9545);
nand U12206 (N_12206,N_7262,N_6486);
or U12207 (N_12207,N_8230,N_8285);
xor U12208 (N_12208,N_6554,N_7490);
or U12209 (N_12209,N_8461,N_9328);
and U12210 (N_12210,N_8308,N_6145);
or U12211 (N_12211,N_8247,N_7074);
and U12212 (N_12212,N_6344,N_7423);
and U12213 (N_12213,N_9815,N_6566);
nand U12214 (N_12214,N_6445,N_7113);
or U12215 (N_12215,N_7798,N_5967);
xnor U12216 (N_12216,N_5824,N_6197);
xor U12217 (N_12217,N_7326,N_7746);
nor U12218 (N_12218,N_9000,N_9977);
nor U12219 (N_12219,N_6098,N_5282);
or U12220 (N_12220,N_8041,N_9663);
or U12221 (N_12221,N_9339,N_6439);
or U12222 (N_12222,N_8213,N_9833);
nor U12223 (N_12223,N_6035,N_8379);
and U12224 (N_12224,N_9024,N_7541);
or U12225 (N_12225,N_7286,N_7999);
nor U12226 (N_12226,N_8876,N_7902);
nand U12227 (N_12227,N_7436,N_5353);
nor U12228 (N_12228,N_8231,N_9329);
nor U12229 (N_12229,N_7337,N_6523);
nor U12230 (N_12230,N_8427,N_7833);
xor U12231 (N_12231,N_6697,N_5585);
or U12232 (N_12232,N_8816,N_8474);
nor U12233 (N_12233,N_7005,N_8493);
and U12234 (N_12234,N_9579,N_7888);
or U12235 (N_12235,N_8727,N_5719);
xor U12236 (N_12236,N_5218,N_9612);
or U12237 (N_12237,N_7770,N_8825);
nand U12238 (N_12238,N_7552,N_8852);
and U12239 (N_12239,N_6560,N_8128);
or U12240 (N_12240,N_5106,N_9051);
nand U12241 (N_12241,N_8563,N_8592);
or U12242 (N_12242,N_7083,N_5566);
and U12243 (N_12243,N_9286,N_8417);
nand U12244 (N_12244,N_8228,N_7695);
nand U12245 (N_12245,N_7023,N_9224);
and U12246 (N_12246,N_7665,N_5126);
nor U12247 (N_12247,N_6550,N_6241);
and U12248 (N_12248,N_7237,N_6235);
nor U12249 (N_12249,N_5420,N_8985);
and U12250 (N_12250,N_5121,N_9806);
and U12251 (N_12251,N_9982,N_9695);
xnor U12252 (N_12252,N_7992,N_6341);
or U12253 (N_12253,N_5731,N_6606);
nand U12254 (N_12254,N_6215,N_9157);
xor U12255 (N_12255,N_6579,N_9632);
and U12256 (N_12256,N_6977,N_6984);
nor U12257 (N_12257,N_5500,N_7520);
nand U12258 (N_12258,N_9931,N_6779);
and U12259 (N_12259,N_7072,N_5621);
or U12260 (N_12260,N_9964,N_9672);
and U12261 (N_12261,N_9755,N_8693);
nor U12262 (N_12262,N_5048,N_6954);
xnor U12263 (N_12263,N_8793,N_9473);
or U12264 (N_12264,N_5273,N_5165);
and U12265 (N_12265,N_7538,N_9476);
nor U12266 (N_12266,N_5074,N_7825);
and U12267 (N_12267,N_7572,N_8614);
xor U12268 (N_12268,N_6749,N_9406);
nand U12269 (N_12269,N_6424,N_9457);
and U12270 (N_12270,N_7247,N_7642);
and U12271 (N_12271,N_9064,N_7838);
nor U12272 (N_12272,N_8934,N_8975);
nor U12273 (N_12273,N_7634,N_6039);
or U12274 (N_12274,N_6661,N_7208);
xor U12275 (N_12275,N_8197,N_9426);
and U12276 (N_12276,N_7213,N_8178);
or U12277 (N_12277,N_8942,N_9846);
and U12278 (N_12278,N_6715,N_9392);
nand U12279 (N_12279,N_9556,N_8315);
nand U12280 (N_12280,N_9720,N_6339);
nor U12281 (N_12281,N_7671,N_6737);
xnor U12282 (N_12282,N_8206,N_5242);
nor U12283 (N_12283,N_5755,N_7219);
xor U12284 (N_12284,N_5699,N_5928);
nor U12285 (N_12285,N_9638,N_8840);
nand U12286 (N_12286,N_7614,N_7488);
nor U12287 (N_12287,N_7929,N_6798);
and U12288 (N_12288,N_7919,N_5947);
xor U12289 (N_12289,N_6504,N_6481);
xor U12290 (N_12290,N_8121,N_5199);
nor U12291 (N_12291,N_6163,N_9980);
and U12292 (N_12292,N_5245,N_5629);
nand U12293 (N_12293,N_7374,N_6742);
nand U12294 (N_12294,N_6287,N_8129);
nor U12295 (N_12295,N_9967,N_6091);
nand U12296 (N_12296,N_5641,N_5072);
nor U12297 (N_12297,N_5745,N_7517);
or U12298 (N_12298,N_6138,N_8069);
nand U12299 (N_12299,N_5011,N_9590);
nor U12300 (N_12300,N_9285,N_8618);
or U12301 (N_12301,N_8561,N_5309);
nand U12302 (N_12302,N_9685,N_7769);
nand U12303 (N_12303,N_5802,N_6360);
and U12304 (N_12304,N_7217,N_9316);
nand U12305 (N_12305,N_5896,N_7180);
and U12306 (N_12306,N_6292,N_7273);
xor U12307 (N_12307,N_9862,N_8122);
or U12308 (N_12308,N_9089,N_5335);
or U12309 (N_12309,N_7395,N_8872);
nor U12310 (N_12310,N_9587,N_5006);
or U12311 (N_12311,N_9789,N_6856);
nor U12312 (N_12312,N_5062,N_9411);
or U12313 (N_12313,N_7477,N_7621);
nand U12314 (N_12314,N_5833,N_6275);
xor U12315 (N_12315,N_5788,N_6717);
or U12316 (N_12316,N_8695,N_7743);
nor U12317 (N_12317,N_6244,N_8380);
or U12318 (N_12318,N_7993,N_7176);
nand U12319 (N_12319,N_7895,N_9901);
and U12320 (N_12320,N_8533,N_5014);
and U12321 (N_12321,N_9462,N_8330);
nand U12322 (N_12322,N_7842,N_5809);
nor U12323 (N_12323,N_6377,N_9389);
nand U12324 (N_12324,N_6298,N_7254);
and U12325 (N_12325,N_7456,N_8126);
nand U12326 (N_12326,N_9218,N_9534);
nand U12327 (N_12327,N_8201,N_7557);
and U12328 (N_12328,N_6987,N_5100);
nand U12329 (N_12329,N_6421,N_7105);
and U12330 (N_12330,N_7685,N_6858);
nor U12331 (N_12331,N_9669,N_6712);
or U12332 (N_12332,N_7844,N_7145);
or U12333 (N_12333,N_9902,N_8146);
or U12334 (N_12334,N_5118,N_7249);
xnor U12335 (N_12335,N_8363,N_7878);
and U12336 (N_12336,N_5265,N_9637);
or U12337 (N_12337,N_7478,N_5637);
or U12338 (N_12338,N_5587,N_9433);
or U12339 (N_12339,N_6310,N_9583);
and U12340 (N_12340,N_8160,N_6768);
xnor U12341 (N_12341,N_8322,N_5571);
and U12342 (N_12342,N_5554,N_6892);
nand U12343 (N_12343,N_9523,N_7207);
xnor U12344 (N_12344,N_7022,N_8149);
nand U12345 (N_12345,N_6527,N_9947);
nor U12346 (N_12346,N_7125,N_6716);
xor U12347 (N_12347,N_9492,N_8995);
nand U12348 (N_12348,N_5278,N_9046);
and U12349 (N_12349,N_7594,N_5417);
and U12350 (N_12350,N_6322,N_5250);
or U12351 (N_12351,N_9581,N_9093);
and U12352 (N_12352,N_8114,N_9865);
or U12353 (N_12353,N_8611,N_5904);
nand U12354 (N_12354,N_6245,N_6013);
or U12355 (N_12355,N_8629,N_7131);
and U12356 (N_12356,N_5038,N_9829);
xnor U12357 (N_12357,N_8514,N_5732);
nor U12358 (N_12358,N_6834,N_5548);
nand U12359 (N_12359,N_5579,N_6611);
and U12360 (N_12360,N_7726,N_5315);
xnor U12361 (N_12361,N_9164,N_9501);
or U12362 (N_12362,N_7558,N_6429);
nand U12363 (N_12363,N_7903,N_6014);
nor U12364 (N_12364,N_5204,N_8466);
nand U12365 (N_12365,N_5859,N_7581);
and U12366 (N_12366,N_5701,N_6057);
or U12367 (N_12367,N_5668,N_5655);
nor U12368 (N_12368,N_6526,N_5680);
nor U12369 (N_12369,N_8587,N_9427);
nand U12370 (N_12370,N_6777,N_6172);
nor U12371 (N_12371,N_8426,N_7411);
nor U12372 (N_12372,N_6763,N_5748);
or U12373 (N_12373,N_5530,N_8782);
xnor U12374 (N_12374,N_5401,N_6046);
nand U12375 (N_12375,N_8813,N_5993);
or U12376 (N_12376,N_7693,N_7114);
or U12377 (N_12377,N_7296,N_9174);
nand U12378 (N_12378,N_6816,N_6109);
or U12379 (N_12379,N_7873,N_8981);
nand U12380 (N_12380,N_5761,N_5414);
and U12381 (N_12381,N_8321,N_6498);
or U12382 (N_12382,N_7489,N_5989);
nand U12383 (N_12383,N_5666,N_9572);
nand U12384 (N_12384,N_8235,N_6461);
and U12385 (N_12385,N_6240,N_8580);
or U12386 (N_12386,N_8483,N_9952);
xor U12387 (N_12387,N_9097,N_6603);
or U12388 (N_12388,N_6654,N_9418);
nor U12389 (N_12389,N_6397,N_9261);
and U12390 (N_12390,N_6411,N_8998);
nand U12391 (N_12391,N_6246,N_7711);
nor U12392 (N_12392,N_9677,N_8112);
or U12393 (N_12393,N_5979,N_6476);
nor U12394 (N_12394,N_7684,N_5873);
nand U12395 (N_12395,N_5616,N_7630);
nand U12396 (N_12396,N_6595,N_8360);
nand U12397 (N_12397,N_9314,N_8645);
or U12398 (N_12398,N_8604,N_5339);
nor U12399 (N_12399,N_6765,N_8500);
nor U12400 (N_12400,N_8218,N_8777);
or U12401 (N_12401,N_9676,N_8300);
nand U12402 (N_12402,N_7162,N_6659);
or U12403 (N_12403,N_9393,N_8091);
xor U12404 (N_12404,N_5283,N_8369);
or U12405 (N_12405,N_9536,N_5733);
nand U12406 (N_12406,N_6435,N_9893);
nand U12407 (N_12407,N_6682,N_7504);
and U12408 (N_12408,N_5189,N_8086);
or U12409 (N_12409,N_5157,N_8076);
or U12410 (N_12410,N_8844,N_6746);
nand U12411 (N_12411,N_8062,N_6117);
or U12412 (N_12412,N_8023,N_9598);
nor U12413 (N_12413,N_7106,N_5891);
nand U12414 (N_12414,N_6844,N_6584);
nor U12415 (N_12415,N_6693,N_5368);
or U12416 (N_12416,N_5741,N_8827);
and U12417 (N_12417,N_9297,N_8633);
nand U12418 (N_12418,N_8021,N_6382);
and U12419 (N_12419,N_7682,N_5210);
xnor U12420 (N_12420,N_6336,N_9214);
nor U12421 (N_12421,N_9003,N_7293);
and U12422 (N_12422,N_9445,N_9560);
and U12423 (N_12423,N_6391,N_9158);
nand U12424 (N_12424,N_5604,N_8212);
nor U12425 (N_12425,N_9050,N_7032);
nand U12426 (N_12426,N_8031,N_6778);
nor U12427 (N_12427,N_6877,N_5296);
and U12428 (N_12428,N_8097,N_6283);
nand U12429 (N_12429,N_6993,N_7817);
nor U12430 (N_12430,N_9489,N_9283);
nor U12431 (N_12431,N_9015,N_5344);
and U12432 (N_12432,N_6735,N_6904);
xnor U12433 (N_12433,N_8107,N_9135);
nand U12434 (N_12434,N_5035,N_9276);
nor U12435 (N_12435,N_7133,N_6574);
and U12436 (N_12436,N_5147,N_7016);
and U12437 (N_12437,N_6813,N_5826);
xor U12438 (N_12438,N_7450,N_7112);
or U12439 (N_12439,N_6306,N_9440);
and U12440 (N_12440,N_9326,N_7747);
nand U12441 (N_12441,N_5415,N_9152);
and U12442 (N_12442,N_9397,N_7562);
or U12443 (N_12443,N_5922,N_8056);
and U12444 (N_12444,N_8657,N_6667);
nand U12445 (N_12445,N_6335,N_8007);
or U12446 (N_12446,N_5066,N_9711);
nand U12447 (N_12447,N_9795,N_9895);
nand U12448 (N_12448,N_8758,N_5588);
nand U12449 (N_12449,N_6111,N_7185);
and U12450 (N_12450,N_8915,N_5771);
nand U12451 (N_12451,N_6243,N_7049);
and U12452 (N_12452,N_9650,N_7629);
xor U12453 (N_12453,N_8639,N_5899);
or U12454 (N_12454,N_7021,N_9950);
nand U12455 (N_12455,N_8550,N_9075);
and U12456 (N_12456,N_7540,N_8979);
and U12457 (N_12457,N_6204,N_5844);
or U12458 (N_12458,N_5290,N_9198);
and U12459 (N_12459,N_8002,N_6515);
or U12460 (N_12460,N_7734,N_6123);
and U12461 (N_12461,N_8020,N_6124);
nand U12462 (N_12462,N_6979,N_9527);
or U12463 (N_12463,N_9017,N_9970);
nand U12464 (N_12464,N_6866,N_6920);
and U12465 (N_12465,N_6004,N_5381);
nand U12466 (N_12466,N_7018,N_5783);
and U12467 (N_12467,N_9735,N_9284);
nor U12468 (N_12468,N_7415,N_6303);
nor U12469 (N_12469,N_8932,N_7431);
nor U12470 (N_12470,N_5615,N_8246);
nor U12471 (N_12471,N_7459,N_6307);
nand U12472 (N_12472,N_6441,N_8353);
nor U12473 (N_12473,N_8404,N_9797);
and U12474 (N_12474,N_8673,N_5516);
nor U12475 (N_12475,N_6259,N_7245);
nor U12476 (N_12476,N_8552,N_7843);
nor U12477 (N_12477,N_8502,N_8869);
and U12478 (N_12478,N_7050,N_9288);
and U12479 (N_12479,N_7739,N_5965);
xor U12480 (N_12480,N_8711,N_9307);
or U12481 (N_12481,N_6162,N_8858);
xor U12482 (N_12482,N_8209,N_9232);
nor U12483 (N_12483,N_6238,N_7507);
and U12484 (N_12484,N_5033,N_7837);
nand U12485 (N_12485,N_7566,N_7466);
nand U12486 (N_12486,N_5408,N_6980);
and U12487 (N_12487,N_6630,N_6010);
or U12488 (N_12488,N_5496,N_9221);
nand U12489 (N_12489,N_5598,N_5685);
or U12490 (N_12490,N_6914,N_9636);
nor U12491 (N_12491,N_9991,N_6940);
nor U12492 (N_12492,N_8098,N_6757);
and U12493 (N_12493,N_9781,N_9700);
and U12494 (N_12494,N_9045,N_8291);
nand U12495 (N_12495,N_6827,N_7616);
or U12496 (N_12496,N_8723,N_5819);
nand U12497 (N_12497,N_9354,N_6359);
and U12498 (N_12498,N_5063,N_6578);
nor U12499 (N_12499,N_8413,N_5992);
nor U12500 (N_12500,N_8270,N_8580);
and U12501 (N_12501,N_6056,N_6818);
and U12502 (N_12502,N_5121,N_8916);
xor U12503 (N_12503,N_5439,N_5356);
or U12504 (N_12504,N_6774,N_5392);
nand U12505 (N_12505,N_7885,N_6066);
nand U12506 (N_12506,N_9906,N_5760);
xnor U12507 (N_12507,N_7250,N_8717);
nor U12508 (N_12508,N_7995,N_6432);
or U12509 (N_12509,N_9085,N_6133);
or U12510 (N_12510,N_6338,N_7813);
xor U12511 (N_12511,N_8013,N_7093);
and U12512 (N_12512,N_7572,N_9401);
or U12513 (N_12513,N_7758,N_7398);
xnor U12514 (N_12514,N_6709,N_9138);
nand U12515 (N_12515,N_8338,N_6955);
xor U12516 (N_12516,N_8929,N_9263);
or U12517 (N_12517,N_8490,N_5335);
or U12518 (N_12518,N_9721,N_6529);
xor U12519 (N_12519,N_7053,N_7359);
and U12520 (N_12520,N_5392,N_7406);
nor U12521 (N_12521,N_5637,N_5921);
and U12522 (N_12522,N_8459,N_9935);
xor U12523 (N_12523,N_6942,N_8718);
and U12524 (N_12524,N_7989,N_5378);
nand U12525 (N_12525,N_7628,N_8329);
nor U12526 (N_12526,N_9646,N_5077);
nor U12527 (N_12527,N_7300,N_7258);
nor U12528 (N_12528,N_5304,N_6631);
nand U12529 (N_12529,N_7093,N_8425);
and U12530 (N_12530,N_8656,N_5727);
or U12531 (N_12531,N_7826,N_9074);
nor U12532 (N_12532,N_5117,N_5663);
nor U12533 (N_12533,N_8115,N_7857);
or U12534 (N_12534,N_9523,N_7598);
xor U12535 (N_12535,N_5156,N_5273);
nand U12536 (N_12536,N_8257,N_9649);
nand U12537 (N_12537,N_8144,N_5983);
or U12538 (N_12538,N_9844,N_8349);
nand U12539 (N_12539,N_7091,N_5589);
nor U12540 (N_12540,N_5886,N_6167);
nand U12541 (N_12541,N_5064,N_7446);
and U12542 (N_12542,N_8393,N_5388);
nor U12543 (N_12543,N_7336,N_8093);
or U12544 (N_12544,N_9936,N_6777);
and U12545 (N_12545,N_6555,N_5527);
or U12546 (N_12546,N_7779,N_9259);
nand U12547 (N_12547,N_9816,N_6949);
nand U12548 (N_12548,N_5874,N_5206);
nand U12549 (N_12549,N_5372,N_6378);
nor U12550 (N_12550,N_6215,N_6863);
nor U12551 (N_12551,N_6179,N_9793);
or U12552 (N_12552,N_8952,N_9617);
nand U12553 (N_12553,N_6583,N_7836);
or U12554 (N_12554,N_5081,N_9271);
nand U12555 (N_12555,N_8888,N_9249);
nand U12556 (N_12556,N_6313,N_8788);
or U12557 (N_12557,N_8385,N_6895);
and U12558 (N_12558,N_9101,N_9138);
and U12559 (N_12559,N_7206,N_8280);
and U12560 (N_12560,N_5659,N_7926);
or U12561 (N_12561,N_9494,N_7601);
xnor U12562 (N_12562,N_6732,N_8435);
and U12563 (N_12563,N_8809,N_9667);
nand U12564 (N_12564,N_8810,N_9113);
and U12565 (N_12565,N_8067,N_6432);
nand U12566 (N_12566,N_9518,N_7160);
or U12567 (N_12567,N_5385,N_7860);
and U12568 (N_12568,N_9433,N_6011);
and U12569 (N_12569,N_5733,N_9619);
and U12570 (N_12570,N_5293,N_6430);
xnor U12571 (N_12571,N_7973,N_7055);
nor U12572 (N_12572,N_6768,N_8127);
nor U12573 (N_12573,N_7362,N_7706);
nand U12574 (N_12574,N_6706,N_5181);
xnor U12575 (N_12575,N_6119,N_7623);
xor U12576 (N_12576,N_6993,N_5825);
nor U12577 (N_12577,N_7218,N_8410);
and U12578 (N_12578,N_6361,N_8921);
nor U12579 (N_12579,N_6396,N_8224);
and U12580 (N_12580,N_5081,N_7669);
nand U12581 (N_12581,N_5286,N_8160);
and U12582 (N_12582,N_7467,N_6775);
or U12583 (N_12583,N_5773,N_6794);
or U12584 (N_12584,N_7731,N_6884);
or U12585 (N_12585,N_7597,N_9441);
nor U12586 (N_12586,N_8180,N_7854);
xor U12587 (N_12587,N_7492,N_9247);
nor U12588 (N_12588,N_6009,N_5237);
nor U12589 (N_12589,N_6990,N_7181);
nor U12590 (N_12590,N_8162,N_8340);
nor U12591 (N_12591,N_5863,N_7483);
and U12592 (N_12592,N_9372,N_6454);
or U12593 (N_12593,N_8139,N_9701);
or U12594 (N_12594,N_6864,N_7536);
or U12595 (N_12595,N_5966,N_7679);
nor U12596 (N_12596,N_8151,N_6991);
nor U12597 (N_12597,N_7990,N_8755);
nand U12598 (N_12598,N_6645,N_5659);
nand U12599 (N_12599,N_5654,N_7318);
or U12600 (N_12600,N_5585,N_7952);
xnor U12601 (N_12601,N_7998,N_5642);
or U12602 (N_12602,N_9344,N_5984);
and U12603 (N_12603,N_5984,N_7165);
nor U12604 (N_12604,N_8773,N_9506);
or U12605 (N_12605,N_5408,N_5595);
and U12606 (N_12606,N_5526,N_6521);
xnor U12607 (N_12607,N_5359,N_7262);
nor U12608 (N_12608,N_7304,N_9656);
nand U12609 (N_12609,N_5291,N_7784);
or U12610 (N_12610,N_8318,N_8978);
nand U12611 (N_12611,N_8728,N_8162);
or U12612 (N_12612,N_5479,N_8039);
xor U12613 (N_12613,N_8415,N_5445);
xnor U12614 (N_12614,N_7235,N_9628);
and U12615 (N_12615,N_7782,N_8115);
xor U12616 (N_12616,N_9302,N_6027);
and U12617 (N_12617,N_9283,N_9938);
nor U12618 (N_12618,N_8691,N_5925);
nor U12619 (N_12619,N_8413,N_7573);
nand U12620 (N_12620,N_7976,N_7142);
and U12621 (N_12621,N_6025,N_8517);
nor U12622 (N_12622,N_8521,N_8833);
nand U12623 (N_12623,N_5454,N_9350);
nor U12624 (N_12624,N_9714,N_7461);
nor U12625 (N_12625,N_8134,N_7611);
or U12626 (N_12626,N_5127,N_7270);
and U12627 (N_12627,N_6401,N_9896);
and U12628 (N_12628,N_6301,N_9833);
xor U12629 (N_12629,N_8065,N_7439);
or U12630 (N_12630,N_7194,N_7789);
nand U12631 (N_12631,N_8436,N_6630);
and U12632 (N_12632,N_6928,N_9001);
and U12633 (N_12633,N_9009,N_6013);
nand U12634 (N_12634,N_8532,N_6327);
or U12635 (N_12635,N_9623,N_7001);
and U12636 (N_12636,N_9050,N_7252);
and U12637 (N_12637,N_9057,N_8297);
or U12638 (N_12638,N_8248,N_7471);
and U12639 (N_12639,N_9949,N_8912);
or U12640 (N_12640,N_7071,N_9073);
nor U12641 (N_12641,N_7280,N_5996);
or U12642 (N_12642,N_9334,N_9719);
nand U12643 (N_12643,N_7376,N_8824);
and U12644 (N_12644,N_7932,N_8893);
nand U12645 (N_12645,N_5381,N_9158);
nor U12646 (N_12646,N_7467,N_9868);
nor U12647 (N_12647,N_6676,N_6733);
or U12648 (N_12648,N_6592,N_8004);
and U12649 (N_12649,N_6352,N_9061);
or U12650 (N_12650,N_9350,N_6207);
or U12651 (N_12651,N_9589,N_6004);
and U12652 (N_12652,N_8903,N_7232);
or U12653 (N_12653,N_6042,N_6045);
nand U12654 (N_12654,N_9458,N_8134);
nor U12655 (N_12655,N_8813,N_8245);
nand U12656 (N_12656,N_6131,N_5861);
or U12657 (N_12657,N_6723,N_5844);
nand U12658 (N_12658,N_9546,N_6674);
and U12659 (N_12659,N_9465,N_9921);
and U12660 (N_12660,N_6815,N_6481);
nor U12661 (N_12661,N_5417,N_5785);
or U12662 (N_12662,N_6162,N_8141);
nor U12663 (N_12663,N_9322,N_5334);
nor U12664 (N_12664,N_5078,N_7020);
or U12665 (N_12665,N_5113,N_6746);
or U12666 (N_12666,N_6329,N_6418);
xor U12667 (N_12667,N_5001,N_7557);
nor U12668 (N_12668,N_6844,N_6770);
or U12669 (N_12669,N_6890,N_9336);
nand U12670 (N_12670,N_7142,N_5826);
or U12671 (N_12671,N_5104,N_9304);
and U12672 (N_12672,N_6224,N_6236);
nor U12673 (N_12673,N_7088,N_9383);
nor U12674 (N_12674,N_5363,N_6369);
nor U12675 (N_12675,N_9379,N_8646);
and U12676 (N_12676,N_5261,N_7239);
and U12677 (N_12677,N_8147,N_5416);
and U12678 (N_12678,N_7720,N_6011);
nand U12679 (N_12679,N_9683,N_7484);
or U12680 (N_12680,N_7331,N_5952);
and U12681 (N_12681,N_9409,N_6636);
nand U12682 (N_12682,N_6537,N_6357);
or U12683 (N_12683,N_8618,N_7863);
and U12684 (N_12684,N_9678,N_7754);
or U12685 (N_12685,N_6757,N_9071);
nand U12686 (N_12686,N_5560,N_9119);
nand U12687 (N_12687,N_5325,N_6819);
and U12688 (N_12688,N_7466,N_7478);
xor U12689 (N_12689,N_7756,N_5074);
nand U12690 (N_12690,N_8158,N_5526);
or U12691 (N_12691,N_7320,N_8718);
nor U12692 (N_12692,N_5770,N_8193);
nor U12693 (N_12693,N_8801,N_9556);
nor U12694 (N_12694,N_5372,N_5674);
nor U12695 (N_12695,N_6986,N_5643);
nand U12696 (N_12696,N_9230,N_5862);
and U12697 (N_12697,N_8240,N_6411);
nand U12698 (N_12698,N_6432,N_5227);
nor U12699 (N_12699,N_7814,N_6205);
nand U12700 (N_12700,N_5231,N_9224);
and U12701 (N_12701,N_8867,N_8939);
and U12702 (N_12702,N_9831,N_8560);
xnor U12703 (N_12703,N_8319,N_5441);
and U12704 (N_12704,N_5625,N_6528);
or U12705 (N_12705,N_6162,N_5462);
nand U12706 (N_12706,N_8823,N_8508);
nand U12707 (N_12707,N_7510,N_8140);
or U12708 (N_12708,N_8892,N_9554);
and U12709 (N_12709,N_8569,N_7276);
nand U12710 (N_12710,N_6917,N_8205);
nor U12711 (N_12711,N_7354,N_7544);
and U12712 (N_12712,N_7906,N_8383);
nor U12713 (N_12713,N_7936,N_7260);
or U12714 (N_12714,N_8979,N_9225);
or U12715 (N_12715,N_7299,N_5621);
or U12716 (N_12716,N_7032,N_6224);
nor U12717 (N_12717,N_8113,N_6025);
and U12718 (N_12718,N_6299,N_5316);
or U12719 (N_12719,N_8475,N_6123);
nor U12720 (N_12720,N_9824,N_9573);
and U12721 (N_12721,N_6910,N_5345);
and U12722 (N_12722,N_5415,N_7730);
nor U12723 (N_12723,N_7303,N_9849);
xor U12724 (N_12724,N_6946,N_9519);
and U12725 (N_12725,N_5314,N_9236);
or U12726 (N_12726,N_9738,N_8000);
or U12727 (N_12727,N_6475,N_6989);
nand U12728 (N_12728,N_7336,N_5876);
nor U12729 (N_12729,N_7057,N_5032);
or U12730 (N_12730,N_6649,N_5602);
and U12731 (N_12731,N_7928,N_7550);
or U12732 (N_12732,N_6896,N_7427);
nand U12733 (N_12733,N_6902,N_6689);
xor U12734 (N_12734,N_6529,N_5212);
and U12735 (N_12735,N_5845,N_5479);
nand U12736 (N_12736,N_8324,N_9776);
nor U12737 (N_12737,N_6803,N_8748);
and U12738 (N_12738,N_5059,N_5533);
or U12739 (N_12739,N_7038,N_7644);
nand U12740 (N_12740,N_8325,N_6300);
nor U12741 (N_12741,N_6630,N_8557);
nor U12742 (N_12742,N_9938,N_8978);
and U12743 (N_12743,N_5997,N_9121);
nand U12744 (N_12744,N_8161,N_7353);
nor U12745 (N_12745,N_6508,N_8854);
and U12746 (N_12746,N_9430,N_8566);
or U12747 (N_12747,N_7365,N_7755);
and U12748 (N_12748,N_5481,N_7055);
nor U12749 (N_12749,N_5821,N_5981);
and U12750 (N_12750,N_9378,N_9259);
or U12751 (N_12751,N_6454,N_5622);
and U12752 (N_12752,N_9186,N_7155);
xnor U12753 (N_12753,N_5938,N_8027);
nor U12754 (N_12754,N_6251,N_7986);
nand U12755 (N_12755,N_6368,N_5356);
nand U12756 (N_12756,N_8116,N_7071);
nand U12757 (N_12757,N_9450,N_7763);
nor U12758 (N_12758,N_9669,N_8904);
nor U12759 (N_12759,N_6537,N_7396);
nand U12760 (N_12760,N_5575,N_7181);
nor U12761 (N_12761,N_6789,N_6387);
xor U12762 (N_12762,N_7526,N_7108);
and U12763 (N_12763,N_7308,N_7631);
and U12764 (N_12764,N_5667,N_5519);
and U12765 (N_12765,N_8352,N_5440);
or U12766 (N_12766,N_5924,N_6336);
and U12767 (N_12767,N_5844,N_9075);
and U12768 (N_12768,N_6123,N_8256);
nand U12769 (N_12769,N_5392,N_7252);
nand U12770 (N_12770,N_9381,N_5963);
xnor U12771 (N_12771,N_7537,N_6873);
nand U12772 (N_12772,N_7651,N_9657);
and U12773 (N_12773,N_6147,N_5515);
and U12774 (N_12774,N_7530,N_6264);
nand U12775 (N_12775,N_7981,N_8552);
nor U12776 (N_12776,N_8236,N_7244);
or U12777 (N_12777,N_8314,N_7810);
and U12778 (N_12778,N_5103,N_5638);
nor U12779 (N_12779,N_6686,N_5110);
nand U12780 (N_12780,N_8621,N_6289);
nor U12781 (N_12781,N_8785,N_9039);
nor U12782 (N_12782,N_7011,N_5175);
nand U12783 (N_12783,N_8644,N_7475);
nor U12784 (N_12784,N_8442,N_7883);
nand U12785 (N_12785,N_5167,N_7591);
or U12786 (N_12786,N_9676,N_5912);
or U12787 (N_12787,N_6983,N_5921);
or U12788 (N_12788,N_5404,N_6038);
nand U12789 (N_12789,N_9589,N_6258);
or U12790 (N_12790,N_8628,N_6657);
nand U12791 (N_12791,N_7076,N_5146);
or U12792 (N_12792,N_9759,N_6525);
nor U12793 (N_12793,N_8092,N_5375);
xnor U12794 (N_12794,N_9359,N_7774);
and U12795 (N_12795,N_5349,N_5723);
nor U12796 (N_12796,N_9623,N_5137);
xor U12797 (N_12797,N_9742,N_6569);
nand U12798 (N_12798,N_6982,N_7099);
or U12799 (N_12799,N_6068,N_6077);
nand U12800 (N_12800,N_9425,N_8163);
nor U12801 (N_12801,N_9449,N_5672);
nand U12802 (N_12802,N_5666,N_9086);
nor U12803 (N_12803,N_6317,N_6841);
nor U12804 (N_12804,N_7442,N_8005);
nor U12805 (N_12805,N_5428,N_7556);
and U12806 (N_12806,N_8701,N_9811);
nor U12807 (N_12807,N_7887,N_5742);
nor U12808 (N_12808,N_6681,N_7626);
and U12809 (N_12809,N_7001,N_6987);
xnor U12810 (N_12810,N_9788,N_8047);
nor U12811 (N_12811,N_9364,N_7318);
or U12812 (N_12812,N_8407,N_8746);
and U12813 (N_12813,N_5115,N_9958);
or U12814 (N_12814,N_9370,N_5779);
nand U12815 (N_12815,N_8511,N_8987);
xnor U12816 (N_12816,N_9158,N_8587);
and U12817 (N_12817,N_8993,N_9422);
nand U12818 (N_12818,N_9345,N_7130);
and U12819 (N_12819,N_8059,N_8026);
nor U12820 (N_12820,N_9967,N_5309);
nand U12821 (N_12821,N_7846,N_9722);
nand U12822 (N_12822,N_6304,N_8605);
nor U12823 (N_12823,N_6909,N_9897);
xor U12824 (N_12824,N_7288,N_9944);
or U12825 (N_12825,N_7744,N_6797);
nor U12826 (N_12826,N_8148,N_9535);
nand U12827 (N_12827,N_7844,N_7050);
nor U12828 (N_12828,N_7726,N_9371);
and U12829 (N_12829,N_5312,N_5022);
and U12830 (N_12830,N_8177,N_6518);
nand U12831 (N_12831,N_6860,N_6597);
nand U12832 (N_12832,N_6081,N_6221);
nor U12833 (N_12833,N_9986,N_5123);
nand U12834 (N_12834,N_9567,N_7097);
nand U12835 (N_12835,N_6695,N_5779);
nor U12836 (N_12836,N_9460,N_9086);
nor U12837 (N_12837,N_7496,N_6174);
xnor U12838 (N_12838,N_9332,N_8227);
nor U12839 (N_12839,N_5777,N_8057);
and U12840 (N_12840,N_8015,N_5566);
nand U12841 (N_12841,N_8490,N_6052);
or U12842 (N_12842,N_5350,N_5150);
nand U12843 (N_12843,N_8486,N_6034);
nand U12844 (N_12844,N_8791,N_7914);
and U12845 (N_12845,N_8975,N_5800);
nor U12846 (N_12846,N_5611,N_6527);
or U12847 (N_12847,N_8142,N_8751);
xnor U12848 (N_12848,N_5203,N_9279);
or U12849 (N_12849,N_9267,N_9814);
nor U12850 (N_12850,N_6378,N_9857);
nor U12851 (N_12851,N_9378,N_5949);
or U12852 (N_12852,N_9576,N_5910);
or U12853 (N_12853,N_7848,N_6929);
and U12854 (N_12854,N_6584,N_8855);
nor U12855 (N_12855,N_7231,N_6961);
nand U12856 (N_12856,N_7513,N_7982);
nand U12857 (N_12857,N_9466,N_8184);
or U12858 (N_12858,N_6632,N_7695);
or U12859 (N_12859,N_7812,N_9820);
nand U12860 (N_12860,N_8847,N_9391);
or U12861 (N_12861,N_8317,N_9904);
nand U12862 (N_12862,N_7707,N_5953);
nor U12863 (N_12863,N_5244,N_6185);
xor U12864 (N_12864,N_8916,N_8863);
nor U12865 (N_12865,N_6803,N_7284);
or U12866 (N_12866,N_7923,N_5377);
xnor U12867 (N_12867,N_8490,N_8062);
nor U12868 (N_12868,N_7366,N_8864);
nand U12869 (N_12869,N_5123,N_8791);
nor U12870 (N_12870,N_9160,N_6928);
nand U12871 (N_12871,N_6505,N_8630);
nand U12872 (N_12872,N_5209,N_9683);
or U12873 (N_12873,N_5434,N_9289);
nor U12874 (N_12874,N_9675,N_8834);
nand U12875 (N_12875,N_7311,N_8486);
nand U12876 (N_12876,N_6362,N_8961);
nand U12877 (N_12877,N_9294,N_9807);
and U12878 (N_12878,N_8706,N_9272);
nor U12879 (N_12879,N_9287,N_7511);
or U12880 (N_12880,N_7301,N_6244);
nand U12881 (N_12881,N_8982,N_7844);
nand U12882 (N_12882,N_5559,N_5121);
nor U12883 (N_12883,N_5667,N_5208);
nand U12884 (N_12884,N_7866,N_9743);
or U12885 (N_12885,N_9678,N_7962);
nor U12886 (N_12886,N_8397,N_8648);
nor U12887 (N_12887,N_7929,N_6507);
and U12888 (N_12888,N_8301,N_5667);
nand U12889 (N_12889,N_7488,N_7635);
nor U12890 (N_12890,N_9245,N_9251);
and U12891 (N_12891,N_8757,N_7222);
nand U12892 (N_12892,N_8625,N_5496);
or U12893 (N_12893,N_6945,N_8533);
nor U12894 (N_12894,N_7167,N_8339);
nand U12895 (N_12895,N_8811,N_9276);
and U12896 (N_12896,N_8905,N_6508);
and U12897 (N_12897,N_6788,N_6627);
nor U12898 (N_12898,N_7532,N_9843);
xor U12899 (N_12899,N_8768,N_8933);
nor U12900 (N_12900,N_9591,N_5803);
or U12901 (N_12901,N_7317,N_6897);
or U12902 (N_12902,N_5516,N_6553);
nor U12903 (N_12903,N_7085,N_6514);
or U12904 (N_12904,N_7012,N_8113);
and U12905 (N_12905,N_5838,N_8646);
nand U12906 (N_12906,N_8995,N_9098);
nor U12907 (N_12907,N_6225,N_8728);
nand U12908 (N_12908,N_9488,N_7071);
nor U12909 (N_12909,N_5292,N_8540);
nor U12910 (N_12910,N_7344,N_6890);
nand U12911 (N_12911,N_5883,N_7827);
nor U12912 (N_12912,N_5311,N_9726);
nand U12913 (N_12913,N_8428,N_8497);
nor U12914 (N_12914,N_9630,N_6679);
nand U12915 (N_12915,N_6748,N_7970);
or U12916 (N_12916,N_9805,N_7301);
xnor U12917 (N_12917,N_8425,N_5907);
nor U12918 (N_12918,N_5638,N_9501);
and U12919 (N_12919,N_7110,N_5359);
nand U12920 (N_12920,N_6931,N_7911);
and U12921 (N_12921,N_8035,N_8257);
nand U12922 (N_12922,N_6152,N_7422);
and U12923 (N_12923,N_5628,N_9114);
and U12924 (N_12924,N_7105,N_8623);
or U12925 (N_12925,N_9696,N_5259);
and U12926 (N_12926,N_6707,N_5817);
nand U12927 (N_12927,N_5442,N_5699);
or U12928 (N_12928,N_8362,N_9477);
or U12929 (N_12929,N_5324,N_5096);
nor U12930 (N_12930,N_6519,N_5678);
nor U12931 (N_12931,N_6618,N_6596);
nand U12932 (N_12932,N_7347,N_5975);
nand U12933 (N_12933,N_6581,N_5101);
nand U12934 (N_12934,N_7660,N_6123);
xor U12935 (N_12935,N_7295,N_6794);
xnor U12936 (N_12936,N_5479,N_5769);
or U12937 (N_12937,N_8930,N_6528);
nor U12938 (N_12938,N_7878,N_7485);
nand U12939 (N_12939,N_7685,N_6454);
or U12940 (N_12940,N_9195,N_9251);
or U12941 (N_12941,N_7860,N_5702);
or U12942 (N_12942,N_9901,N_6753);
nor U12943 (N_12943,N_8481,N_8893);
and U12944 (N_12944,N_8904,N_5816);
nor U12945 (N_12945,N_8381,N_8801);
nand U12946 (N_12946,N_6088,N_5043);
nand U12947 (N_12947,N_9621,N_8274);
and U12948 (N_12948,N_6105,N_8191);
nand U12949 (N_12949,N_7383,N_6484);
nand U12950 (N_12950,N_8355,N_9873);
nor U12951 (N_12951,N_9016,N_8641);
and U12952 (N_12952,N_6967,N_5775);
or U12953 (N_12953,N_5991,N_8525);
or U12954 (N_12954,N_8755,N_7610);
nand U12955 (N_12955,N_7964,N_6131);
or U12956 (N_12956,N_7743,N_8403);
or U12957 (N_12957,N_9784,N_7668);
or U12958 (N_12958,N_7370,N_6038);
nor U12959 (N_12959,N_9908,N_9174);
xnor U12960 (N_12960,N_5145,N_8862);
or U12961 (N_12961,N_7562,N_8909);
nor U12962 (N_12962,N_9098,N_9464);
xnor U12963 (N_12963,N_6095,N_8313);
nor U12964 (N_12964,N_8892,N_9238);
nand U12965 (N_12965,N_5667,N_9009);
nor U12966 (N_12966,N_5007,N_5281);
nand U12967 (N_12967,N_8861,N_9063);
nand U12968 (N_12968,N_9976,N_5753);
and U12969 (N_12969,N_9374,N_5701);
or U12970 (N_12970,N_9859,N_9985);
or U12971 (N_12971,N_9240,N_5196);
nand U12972 (N_12972,N_8188,N_5444);
or U12973 (N_12973,N_7645,N_5420);
and U12974 (N_12974,N_7113,N_6844);
nor U12975 (N_12975,N_5856,N_8738);
and U12976 (N_12976,N_5446,N_9980);
nor U12977 (N_12977,N_5249,N_7374);
nand U12978 (N_12978,N_9945,N_5696);
nand U12979 (N_12979,N_9723,N_6026);
and U12980 (N_12980,N_5026,N_9724);
xor U12981 (N_12981,N_7540,N_7923);
nand U12982 (N_12982,N_9589,N_6529);
nor U12983 (N_12983,N_7444,N_9481);
and U12984 (N_12984,N_9027,N_9297);
or U12985 (N_12985,N_7355,N_6759);
or U12986 (N_12986,N_7880,N_7575);
and U12987 (N_12987,N_5158,N_5857);
and U12988 (N_12988,N_6874,N_6544);
nor U12989 (N_12989,N_5874,N_9657);
nor U12990 (N_12990,N_8713,N_7520);
and U12991 (N_12991,N_5735,N_7952);
nor U12992 (N_12992,N_9371,N_9527);
and U12993 (N_12993,N_7998,N_7737);
nand U12994 (N_12994,N_7017,N_9062);
nand U12995 (N_12995,N_7280,N_8610);
nor U12996 (N_12996,N_8754,N_9202);
nand U12997 (N_12997,N_6189,N_5761);
and U12998 (N_12998,N_6155,N_6487);
nor U12999 (N_12999,N_5541,N_8406);
nor U13000 (N_13000,N_8897,N_9368);
or U13001 (N_13001,N_7953,N_7932);
nand U13002 (N_13002,N_6036,N_7789);
nor U13003 (N_13003,N_9967,N_7951);
or U13004 (N_13004,N_5718,N_9676);
nand U13005 (N_13005,N_8877,N_7521);
nor U13006 (N_13006,N_8846,N_9921);
and U13007 (N_13007,N_9408,N_7177);
xor U13008 (N_13008,N_8447,N_8485);
or U13009 (N_13009,N_5558,N_7983);
or U13010 (N_13010,N_9737,N_5218);
nor U13011 (N_13011,N_7657,N_7370);
and U13012 (N_13012,N_8350,N_6762);
and U13013 (N_13013,N_8945,N_6347);
nor U13014 (N_13014,N_7096,N_8884);
nand U13015 (N_13015,N_7746,N_7425);
or U13016 (N_13016,N_7021,N_5627);
or U13017 (N_13017,N_9696,N_5425);
or U13018 (N_13018,N_8605,N_5892);
nand U13019 (N_13019,N_8580,N_6486);
nand U13020 (N_13020,N_8386,N_6217);
or U13021 (N_13021,N_5125,N_8548);
and U13022 (N_13022,N_8829,N_7347);
xnor U13023 (N_13023,N_8007,N_5461);
nor U13024 (N_13024,N_6390,N_8513);
and U13025 (N_13025,N_8852,N_8298);
or U13026 (N_13026,N_9518,N_5450);
nand U13027 (N_13027,N_6056,N_5546);
nor U13028 (N_13028,N_9967,N_9210);
or U13029 (N_13029,N_6833,N_7830);
nor U13030 (N_13030,N_5559,N_8879);
and U13031 (N_13031,N_9241,N_5369);
nand U13032 (N_13032,N_8595,N_5525);
nand U13033 (N_13033,N_6746,N_9207);
and U13034 (N_13034,N_8369,N_7794);
or U13035 (N_13035,N_6296,N_6956);
nand U13036 (N_13036,N_6828,N_9319);
nand U13037 (N_13037,N_8922,N_5622);
and U13038 (N_13038,N_8088,N_8134);
or U13039 (N_13039,N_7891,N_6064);
and U13040 (N_13040,N_9023,N_6390);
xor U13041 (N_13041,N_6124,N_9896);
and U13042 (N_13042,N_8215,N_7295);
or U13043 (N_13043,N_9373,N_8642);
or U13044 (N_13044,N_9853,N_8688);
and U13045 (N_13045,N_7616,N_9976);
nor U13046 (N_13046,N_6977,N_8794);
xor U13047 (N_13047,N_7555,N_6365);
or U13048 (N_13048,N_8465,N_9017);
nor U13049 (N_13049,N_5844,N_7681);
and U13050 (N_13050,N_7634,N_6106);
nor U13051 (N_13051,N_7905,N_6344);
nor U13052 (N_13052,N_5272,N_6985);
xor U13053 (N_13053,N_8952,N_7702);
nand U13054 (N_13054,N_8480,N_5152);
nand U13055 (N_13055,N_5290,N_9533);
nor U13056 (N_13056,N_7385,N_9296);
and U13057 (N_13057,N_5508,N_5942);
nor U13058 (N_13058,N_8502,N_5998);
nor U13059 (N_13059,N_5877,N_9840);
nor U13060 (N_13060,N_7326,N_5014);
nor U13061 (N_13061,N_6591,N_8054);
nand U13062 (N_13062,N_9836,N_5675);
nor U13063 (N_13063,N_6498,N_9502);
and U13064 (N_13064,N_7561,N_6905);
nand U13065 (N_13065,N_9735,N_6707);
or U13066 (N_13066,N_5469,N_9345);
nand U13067 (N_13067,N_8788,N_6401);
nand U13068 (N_13068,N_6723,N_7461);
or U13069 (N_13069,N_7282,N_7346);
and U13070 (N_13070,N_5626,N_5200);
or U13071 (N_13071,N_8137,N_7054);
xnor U13072 (N_13072,N_9677,N_7433);
nand U13073 (N_13073,N_7836,N_9114);
or U13074 (N_13074,N_5579,N_8705);
nand U13075 (N_13075,N_7284,N_6279);
xor U13076 (N_13076,N_9221,N_8699);
or U13077 (N_13077,N_8822,N_6601);
nand U13078 (N_13078,N_7657,N_5734);
nand U13079 (N_13079,N_8599,N_9773);
nand U13080 (N_13080,N_5743,N_6211);
and U13081 (N_13081,N_6876,N_9313);
and U13082 (N_13082,N_8921,N_5787);
and U13083 (N_13083,N_8581,N_8297);
nand U13084 (N_13084,N_9691,N_7306);
or U13085 (N_13085,N_6155,N_6966);
nand U13086 (N_13086,N_5270,N_7122);
nand U13087 (N_13087,N_5869,N_8463);
or U13088 (N_13088,N_9913,N_5761);
nor U13089 (N_13089,N_9132,N_9735);
or U13090 (N_13090,N_8440,N_6331);
or U13091 (N_13091,N_6497,N_8699);
nor U13092 (N_13092,N_9200,N_5116);
and U13093 (N_13093,N_7576,N_8993);
or U13094 (N_13094,N_7116,N_5506);
and U13095 (N_13095,N_6032,N_7641);
or U13096 (N_13096,N_9358,N_7550);
and U13097 (N_13097,N_8926,N_9639);
nor U13098 (N_13098,N_6585,N_6138);
nand U13099 (N_13099,N_7398,N_9710);
and U13100 (N_13100,N_8716,N_7740);
or U13101 (N_13101,N_6007,N_5244);
nor U13102 (N_13102,N_8520,N_6998);
nand U13103 (N_13103,N_8811,N_8763);
nand U13104 (N_13104,N_7817,N_5979);
or U13105 (N_13105,N_8021,N_5234);
nor U13106 (N_13106,N_8054,N_8679);
nor U13107 (N_13107,N_6791,N_7715);
and U13108 (N_13108,N_8484,N_6587);
or U13109 (N_13109,N_5438,N_8230);
and U13110 (N_13110,N_6770,N_6951);
or U13111 (N_13111,N_6162,N_6124);
and U13112 (N_13112,N_5545,N_6361);
or U13113 (N_13113,N_8014,N_7881);
and U13114 (N_13114,N_8016,N_7968);
or U13115 (N_13115,N_8339,N_7829);
nand U13116 (N_13116,N_9156,N_6527);
or U13117 (N_13117,N_8200,N_8115);
nand U13118 (N_13118,N_7166,N_7896);
nor U13119 (N_13119,N_7787,N_5936);
nor U13120 (N_13120,N_5716,N_7711);
nand U13121 (N_13121,N_8963,N_7644);
and U13122 (N_13122,N_9978,N_9422);
or U13123 (N_13123,N_8944,N_7340);
nor U13124 (N_13124,N_7237,N_5826);
and U13125 (N_13125,N_6495,N_5864);
or U13126 (N_13126,N_7366,N_8378);
xor U13127 (N_13127,N_9125,N_8309);
or U13128 (N_13128,N_9436,N_9850);
nand U13129 (N_13129,N_7121,N_8091);
and U13130 (N_13130,N_6666,N_7841);
or U13131 (N_13131,N_9385,N_9801);
and U13132 (N_13132,N_5857,N_9757);
and U13133 (N_13133,N_6959,N_6358);
nand U13134 (N_13134,N_5373,N_6261);
nand U13135 (N_13135,N_6247,N_6766);
and U13136 (N_13136,N_8277,N_6544);
nor U13137 (N_13137,N_6039,N_9267);
and U13138 (N_13138,N_8416,N_9202);
xor U13139 (N_13139,N_6391,N_7030);
or U13140 (N_13140,N_6752,N_7601);
nor U13141 (N_13141,N_9058,N_8520);
and U13142 (N_13142,N_5857,N_6287);
nand U13143 (N_13143,N_9389,N_7494);
and U13144 (N_13144,N_8795,N_7281);
and U13145 (N_13145,N_8169,N_5828);
nand U13146 (N_13146,N_9080,N_8187);
and U13147 (N_13147,N_8818,N_7881);
or U13148 (N_13148,N_6512,N_6948);
or U13149 (N_13149,N_7821,N_7394);
and U13150 (N_13150,N_8632,N_8646);
and U13151 (N_13151,N_8232,N_8439);
nand U13152 (N_13152,N_8896,N_9694);
nand U13153 (N_13153,N_9949,N_7936);
nor U13154 (N_13154,N_5242,N_7699);
xor U13155 (N_13155,N_7227,N_6188);
nand U13156 (N_13156,N_9372,N_6066);
nand U13157 (N_13157,N_7938,N_8151);
nand U13158 (N_13158,N_9146,N_6336);
and U13159 (N_13159,N_9215,N_8230);
and U13160 (N_13160,N_5943,N_8454);
and U13161 (N_13161,N_9950,N_5012);
xnor U13162 (N_13162,N_5815,N_8737);
and U13163 (N_13163,N_9085,N_8367);
nor U13164 (N_13164,N_7487,N_8923);
and U13165 (N_13165,N_8471,N_8638);
and U13166 (N_13166,N_6250,N_6513);
or U13167 (N_13167,N_8205,N_8420);
nand U13168 (N_13168,N_6897,N_8715);
and U13169 (N_13169,N_7400,N_9535);
and U13170 (N_13170,N_9480,N_8120);
or U13171 (N_13171,N_6365,N_9351);
nor U13172 (N_13172,N_5878,N_7870);
nor U13173 (N_13173,N_7182,N_9751);
or U13174 (N_13174,N_6515,N_7584);
or U13175 (N_13175,N_6924,N_5262);
nand U13176 (N_13176,N_9725,N_9212);
or U13177 (N_13177,N_9813,N_9416);
and U13178 (N_13178,N_7797,N_7047);
or U13179 (N_13179,N_8221,N_5772);
nor U13180 (N_13180,N_8307,N_9019);
and U13181 (N_13181,N_6631,N_9191);
xor U13182 (N_13182,N_6621,N_6216);
xor U13183 (N_13183,N_6183,N_6405);
nand U13184 (N_13184,N_7842,N_8851);
and U13185 (N_13185,N_8048,N_5606);
nor U13186 (N_13186,N_7682,N_8181);
or U13187 (N_13187,N_7333,N_6997);
and U13188 (N_13188,N_8336,N_5048);
nand U13189 (N_13189,N_5588,N_9815);
or U13190 (N_13190,N_5879,N_5498);
xnor U13191 (N_13191,N_5033,N_7328);
and U13192 (N_13192,N_8058,N_9696);
and U13193 (N_13193,N_7627,N_7208);
and U13194 (N_13194,N_5232,N_9200);
nor U13195 (N_13195,N_9371,N_8359);
or U13196 (N_13196,N_6393,N_6320);
nor U13197 (N_13197,N_9229,N_9251);
or U13198 (N_13198,N_6613,N_6896);
xor U13199 (N_13199,N_7993,N_5944);
and U13200 (N_13200,N_5255,N_6740);
nand U13201 (N_13201,N_9207,N_5438);
or U13202 (N_13202,N_9360,N_8763);
and U13203 (N_13203,N_7074,N_9878);
xor U13204 (N_13204,N_5290,N_9724);
or U13205 (N_13205,N_6847,N_7759);
or U13206 (N_13206,N_6902,N_8293);
xnor U13207 (N_13207,N_9690,N_7719);
and U13208 (N_13208,N_7709,N_6306);
nand U13209 (N_13209,N_7681,N_7796);
and U13210 (N_13210,N_6563,N_9757);
xor U13211 (N_13211,N_9944,N_9060);
xor U13212 (N_13212,N_7292,N_8245);
and U13213 (N_13213,N_7069,N_9189);
or U13214 (N_13214,N_5401,N_5482);
and U13215 (N_13215,N_7490,N_8726);
and U13216 (N_13216,N_6831,N_5973);
nor U13217 (N_13217,N_9558,N_7799);
nor U13218 (N_13218,N_7040,N_9848);
or U13219 (N_13219,N_5959,N_9522);
nor U13220 (N_13220,N_7425,N_8339);
nand U13221 (N_13221,N_5230,N_5305);
nor U13222 (N_13222,N_6972,N_6938);
xor U13223 (N_13223,N_8959,N_5348);
and U13224 (N_13224,N_8158,N_7057);
or U13225 (N_13225,N_7808,N_7681);
xnor U13226 (N_13226,N_8726,N_7165);
xor U13227 (N_13227,N_5361,N_6735);
and U13228 (N_13228,N_8597,N_6069);
nand U13229 (N_13229,N_9374,N_7100);
or U13230 (N_13230,N_6929,N_9973);
nor U13231 (N_13231,N_8188,N_8387);
nand U13232 (N_13232,N_6534,N_6714);
and U13233 (N_13233,N_9765,N_9566);
or U13234 (N_13234,N_6073,N_5442);
nor U13235 (N_13235,N_5648,N_5454);
nand U13236 (N_13236,N_9389,N_8626);
or U13237 (N_13237,N_5448,N_9473);
nand U13238 (N_13238,N_7673,N_8594);
nor U13239 (N_13239,N_7885,N_5306);
or U13240 (N_13240,N_7532,N_8926);
nor U13241 (N_13241,N_6628,N_5137);
and U13242 (N_13242,N_6312,N_5888);
and U13243 (N_13243,N_6233,N_6336);
or U13244 (N_13244,N_8782,N_7154);
nand U13245 (N_13245,N_7953,N_6081);
nand U13246 (N_13246,N_7992,N_6437);
and U13247 (N_13247,N_5861,N_8081);
nor U13248 (N_13248,N_9741,N_7645);
nor U13249 (N_13249,N_7925,N_9973);
nor U13250 (N_13250,N_7633,N_7240);
xnor U13251 (N_13251,N_8860,N_8945);
nor U13252 (N_13252,N_9608,N_8328);
xor U13253 (N_13253,N_9622,N_7688);
nor U13254 (N_13254,N_9067,N_6424);
xor U13255 (N_13255,N_8416,N_6753);
or U13256 (N_13256,N_8582,N_9113);
xnor U13257 (N_13257,N_8649,N_7007);
xor U13258 (N_13258,N_5589,N_7427);
or U13259 (N_13259,N_9965,N_9541);
and U13260 (N_13260,N_7860,N_9320);
nand U13261 (N_13261,N_7250,N_8352);
nor U13262 (N_13262,N_6905,N_7417);
xor U13263 (N_13263,N_8262,N_8457);
nand U13264 (N_13264,N_9952,N_6910);
nand U13265 (N_13265,N_8479,N_9267);
or U13266 (N_13266,N_8100,N_7793);
nand U13267 (N_13267,N_6968,N_7346);
or U13268 (N_13268,N_5913,N_7661);
or U13269 (N_13269,N_8235,N_9294);
or U13270 (N_13270,N_8935,N_7661);
nand U13271 (N_13271,N_9243,N_9434);
or U13272 (N_13272,N_6318,N_7900);
nor U13273 (N_13273,N_9754,N_5698);
and U13274 (N_13274,N_9901,N_8485);
and U13275 (N_13275,N_7528,N_8599);
and U13276 (N_13276,N_6713,N_6866);
nand U13277 (N_13277,N_5978,N_7290);
nand U13278 (N_13278,N_8939,N_7625);
nor U13279 (N_13279,N_9481,N_5954);
or U13280 (N_13280,N_5993,N_6538);
nand U13281 (N_13281,N_9556,N_8192);
and U13282 (N_13282,N_9701,N_5466);
xnor U13283 (N_13283,N_5359,N_6877);
nor U13284 (N_13284,N_9090,N_5366);
nand U13285 (N_13285,N_9184,N_9482);
or U13286 (N_13286,N_7979,N_9864);
xnor U13287 (N_13287,N_5031,N_7669);
xor U13288 (N_13288,N_7881,N_6990);
or U13289 (N_13289,N_5498,N_8998);
and U13290 (N_13290,N_9537,N_8922);
or U13291 (N_13291,N_8818,N_5991);
nand U13292 (N_13292,N_9526,N_7505);
and U13293 (N_13293,N_7952,N_9774);
and U13294 (N_13294,N_6741,N_6519);
nor U13295 (N_13295,N_9359,N_5149);
xnor U13296 (N_13296,N_6823,N_6359);
and U13297 (N_13297,N_6676,N_7312);
or U13298 (N_13298,N_7478,N_7416);
nor U13299 (N_13299,N_8134,N_6877);
nor U13300 (N_13300,N_5934,N_5437);
nor U13301 (N_13301,N_7155,N_5266);
nor U13302 (N_13302,N_6558,N_5996);
and U13303 (N_13303,N_6646,N_5210);
nor U13304 (N_13304,N_6865,N_5901);
or U13305 (N_13305,N_8926,N_7638);
xor U13306 (N_13306,N_8905,N_5973);
nand U13307 (N_13307,N_5744,N_9226);
nor U13308 (N_13308,N_8739,N_7330);
or U13309 (N_13309,N_6764,N_6932);
nand U13310 (N_13310,N_8711,N_9330);
nor U13311 (N_13311,N_5883,N_5010);
and U13312 (N_13312,N_6933,N_7313);
and U13313 (N_13313,N_5973,N_7255);
xor U13314 (N_13314,N_6734,N_7380);
nor U13315 (N_13315,N_8588,N_7391);
nand U13316 (N_13316,N_9667,N_5144);
and U13317 (N_13317,N_7604,N_7568);
or U13318 (N_13318,N_8870,N_7727);
nor U13319 (N_13319,N_9807,N_8485);
nor U13320 (N_13320,N_9432,N_8358);
or U13321 (N_13321,N_8891,N_5146);
xor U13322 (N_13322,N_5128,N_8556);
or U13323 (N_13323,N_8980,N_8260);
nand U13324 (N_13324,N_5397,N_7678);
xor U13325 (N_13325,N_8328,N_8672);
nor U13326 (N_13326,N_5647,N_6611);
and U13327 (N_13327,N_5306,N_7536);
nand U13328 (N_13328,N_5128,N_9566);
and U13329 (N_13329,N_7344,N_7472);
or U13330 (N_13330,N_6446,N_9914);
and U13331 (N_13331,N_7817,N_9067);
xor U13332 (N_13332,N_8060,N_6857);
or U13333 (N_13333,N_6398,N_6045);
and U13334 (N_13334,N_5163,N_5977);
nand U13335 (N_13335,N_7988,N_8118);
nor U13336 (N_13336,N_6045,N_9087);
nand U13337 (N_13337,N_7438,N_9963);
and U13338 (N_13338,N_5832,N_8865);
xor U13339 (N_13339,N_9008,N_8731);
nor U13340 (N_13340,N_8614,N_8591);
xnor U13341 (N_13341,N_5507,N_9892);
or U13342 (N_13342,N_9835,N_6805);
or U13343 (N_13343,N_9406,N_7108);
nand U13344 (N_13344,N_9602,N_5853);
nor U13345 (N_13345,N_9039,N_5978);
nand U13346 (N_13346,N_6612,N_7323);
or U13347 (N_13347,N_5797,N_5736);
nor U13348 (N_13348,N_5996,N_5389);
and U13349 (N_13349,N_7617,N_6022);
xor U13350 (N_13350,N_7199,N_9833);
or U13351 (N_13351,N_6305,N_8854);
nor U13352 (N_13352,N_7981,N_7769);
nand U13353 (N_13353,N_6870,N_6277);
nor U13354 (N_13354,N_5076,N_8924);
or U13355 (N_13355,N_6691,N_8353);
and U13356 (N_13356,N_5134,N_7737);
or U13357 (N_13357,N_6487,N_8160);
or U13358 (N_13358,N_6309,N_6027);
or U13359 (N_13359,N_8015,N_9871);
nand U13360 (N_13360,N_6202,N_8374);
or U13361 (N_13361,N_9012,N_5920);
or U13362 (N_13362,N_7027,N_8725);
nand U13363 (N_13363,N_5926,N_6763);
nand U13364 (N_13364,N_6864,N_5373);
and U13365 (N_13365,N_7816,N_5674);
nand U13366 (N_13366,N_8815,N_7832);
nand U13367 (N_13367,N_8154,N_9320);
nor U13368 (N_13368,N_8247,N_6199);
or U13369 (N_13369,N_8791,N_8295);
or U13370 (N_13370,N_5398,N_5712);
or U13371 (N_13371,N_9885,N_6834);
nor U13372 (N_13372,N_5608,N_8348);
nand U13373 (N_13373,N_5276,N_6122);
and U13374 (N_13374,N_7422,N_7669);
nor U13375 (N_13375,N_9713,N_9531);
nand U13376 (N_13376,N_9308,N_7120);
xor U13377 (N_13377,N_7388,N_7036);
nor U13378 (N_13378,N_6738,N_9308);
nand U13379 (N_13379,N_8219,N_8931);
nand U13380 (N_13380,N_5142,N_5390);
nor U13381 (N_13381,N_8830,N_9045);
nor U13382 (N_13382,N_8219,N_8354);
nand U13383 (N_13383,N_9979,N_6354);
or U13384 (N_13384,N_9479,N_9795);
nor U13385 (N_13385,N_7128,N_9608);
nand U13386 (N_13386,N_8245,N_5806);
nand U13387 (N_13387,N_5511,N_8058);
or U13388 (N_13388,N_5747,N_9135);
or U13389 (N_13389,N_9896,N_8282);
nor U13390 (N_13390,N_9180,N_5039);
nor U13391 (N_13391,N_5348,N_6659);
nor U13392 (N_13392,N_5173,N_7955);
and U13393 (N_13393,N_8168,N_7124);
xor U13394 (N_13394,N_6634,N_9449);
and U13395 (N_13395,N_8675,N_5645);
nand U13396 (N_13396,N_7115,N_9244);
nand U13397 (N_13397,N_9899,N_7983);
nor U13398 (N_13398,N_8195,N_7181);
and U13399 (N_13399,N_8702,N_9143);
and U13400 (N_13400,N_5602,N_5923);
or U13401 (N_13401,N_5379,N_6004);
or U13402 (N_13402,N_7881,N_5603);
or U13403 (N_13403,N_8094,N_9774);
nor U13404 (N_13404,N_5054,N_7790);
or U13405 (N_13405,N_8046,N_8779);
nor U13406 (N_13406,N_9916,N_9193);
nor U13407 (N_13407,N_5970,N_7831);
nand U13408 (N_13408,N_8898,N_9756);
and U13409 (N_13409,N_6863,N_6955);
nor U13410 (N_13410,N_9307,N_7097);
nor U13411 (N_13411,N_9292,N_5922);
and U13412 (N_13412,N_7954,N_8432);
nor U13413 (N_13413,N_9640,N_8575);
and U13414 (N_13414,N_7277,N_6114);
and U13415 (N_13415,N_6667,N_9336);
nand U13416 (N_13416,N_7635,N_6573);
nand U13417 (N_13417,N_7884,N_5213);
or U13418 (N_13418,N_6316,N_7793);
nor U13419 (N_13419,N_8411,N_6387);
and U13420 (N_13420,N_5969,N_7304);
and U13421 (N_13421,N_9085,N_8388);
nor U13422 (N_13422,N_8846,N_7387);
nand U13423 (N_13423,N_7340,N_9058);
nand U13424 (N_13424,N_9318,N_5049);
nor U13425 (N_13425,N_5342,N_6790);
or U13426 (N_13426,N_5983,N_5487);
and U13427 (N_13427,N_6211,N_6279);
nor U13428 (N_13428,N_5144,N_8851);
and U13429 (N_13429,N_7861,N_5486);
and U13430 (N_13430,N_9865,N_5946);
and U13431 (N_13431,N_7648,N_6205);
and U13432 (N_13432,N_5823,N_6067);
nor U13433 (N_13433,N_6901,N_8530);
and U13434 (N_13434,N_6828,N_6806);
or U13435 (N_13435,N_9084,N_9279);
nor U13436 (N_13436,N_5529,N_8569);
nor U13437 (N_13437,N_8809,N_7184);
and U13438 (N_13438,N_6353,N_7958);
and U13439 (N_13439,N_5682,N_6416);
and U13440 (N_13440,N_5055,N_9440);
or U13441 (N_13441,N_8064,N_5936);
and U13442 (N_13442,N_5544,N_7467);
nor U13443 (N_13443,N_5695,N_5916);
nand U13444 (N_13444,N_5171,N_7829);
and U13445 (N_13445,N_6304,N_5046);
and U13446 (N_13446,N_5927,N_9906);
and U13447 (N_13447,N_9898,N_7065);
nand U13448 (N_13448,N_6862,N_5588);
xnor U13449 (N_13449,N_5971,N_7432);
and U13450 (N_13450,N_6277,N_6468);
and U13451 (N_13451,N_5685,N_5652);
xor U13452 (N_13452,N_6575,N_9874);
nand U13453 (N_13453,N_9472,N_7262);
nor U13454 (N_13454,N_9584,N_7533);
xnor U13455 (N_13455,N_7030,N_5638);
nand U13456 (N_13456,N_6967,N_5053);
and U13457 (N_13457,N_6145,N_5489);
or U13458 (N_13458,N_8215,N_9141);
nand U13459 (N_13459,N_6801,N_7243);
or U13460 (N_13460,N_9426,N_7937);
and U13461 (N_13461,N_5790,N_9231);
nor U13462 (N_13462,N_8769,N_5087);
or U13463 (N_13463,N_5034,N_6490);
xor U13464 (N_13464,N_7915,N_9080);
and U13465 (N_13465,N_7440,N_5488);
or U13466 (N_13466,N_6093,N_7690);
xnor U13467 (N_13467,N_9093,N_6175);
or U13468 (N_13468,N_8972,N_6531);
nand U13469 (N_13469,N_7213,N_9744);
nand U13470 (N_13470,N_5576,N_7793);
or U13471 (N_13471,N_8796,N_5815);
or U13472 (N_13472,N_7644,N_8378);
nor U13473 (N_13473,N_5350,N_8423);
nand U13474 (N_13474,N_8614,N_6158);
nor U13475 (N_13475,N_9076,N_6585);
nand U13476 (N_13476,N_6997,N_6359);
nand U13477 (N_13477,N_8419,N_5144);
nand U13478 (N_13478,N_5674,N_7932);
nor U13479 (N_13479,N_6662,N_8581);
nor U13480 (N_13480,N_6652,N_7215);
or U13481 (N_13481,N_9305,N_7629);
nor U13482 (N_13482,N_5496,N_5900);
xnor U13483 (N_13483,N_7784,N_5217);
and U13484 (N_13484,N_6853,N_5344);
and U13485 (N_13485,N_9726,N_7868);
nor U13486 (N_13486,N_8324,N_9178);
nor U13487 (N_13487,N_7426,N_8424);
and U13488 (N_13488,N_6549,N_5687);
and U13489 (N_13489,N_6596,N_5294);
or U13490 (N_13490,N_9816,N_8402);
or U13491 (N_13491,N_6664,N_7074);
nor U13492 (N_13492,N_5539,N_8365);
nand U13493 (N_13493,N_9071,N_6727);
or U13494 (N_13494,N_8715,N_9865);
and U13495 (N_13495,N_5769,N_7606);
or U13496 (N_13496,N_8999,N_5622);
and U13497 (N_13497,N_8207,N_5736);
nand U13498 (N_13498,N_9134,N_5629);
nor U13499 (N_13499,N_5303,N_8155);
or U13500 (N_13500,N_9636,N_5054);
or U13501 (N_13501,N_8893,N_6039);
nand U13502 (N_13502,N_9177,N_8825);
nor U13503 (N_13503,N_9955,N_8387);
nand U13504 (N_13504,N_8435,N_7374);
nor U13505 (N_13505,N_9313,N_6275);
nand U13506 (N_13506,N_7842,N_5060);
nand U13507 (N_13507,N_7585,N_6854);
and U13508 (N_13508,N_7109,N_9649);
nor U13509 (N_13509,N_9242,N_8758);
xor U13510 (N_13510,N_6125,N_8247);
or U13511 (N_13511,N_9738,N_7257);
or U13512 (N_13512,N_5373,N_6317);
nand U13513 (N_13513,N_6861,N_5967);
and U13514 (N_13514,N_9750,N_6921);
and U13515 (N_13515,N_7700,N_7128);
xnor U13516 (N_13516,N_5405,N_6300);
or U13517 (N_13517,N_9996,N_9696);
xnor U13518 (N_13518,N_8525,N_9447);
nor U13519 (N_13519,N_6214,N_7641);
nand U13520 (N_13520,N_7090,N_7887);
and U13521 (N_13521,N_8309,N_8389);
nor U13522 (N_13522,N_9680,N_5052);
nand U13523 (N_13523,N_9129,N_7063);
nand U13524 (N_13524,N_8568,N_7664);
nand U13525 (N_13525,N_9419,N_5334);
or U13526 (N_13526,N_8616,N_6564);
or U13527 (N_13527,N_9296,N_9931);
nor U13528 (N_13528,N_6999,N_6006);
and U13529 (N_13529,N_9103,N_8295);
and U13530 (N_13530,N_6409,N_5290);
nor U13531 (N_13531,N_5217,N_7478);
and U13532 (N_13532,N_8028,N_5500);
nand U13533 (N_13533,N_5527,N_7709);
or U13534 (N_13534,N_5203,N_8815);
nor U13535 (N_13535,N_8671,N_8819);
nand U13536 (N_13536,N_5745,N_6344);
nor U13537 (N_13537,N_8802,N_8990);
nand U13538 (N_13538,N_5178,N_8457);
nand U13539 (N_13539,N_9602,N_9697);
nand U13540 (N_13540,N_5370,N_9329);
nor U13541 (N_13541,N_7501,N_8047);
and U13542 (N_13542,N_5990,N_6135);
nor U13543 (N_13543,N_9663,N_7847);
xor U13544 (N_13544,N_6492,N_8672);
nand U13545 (N_13545,N_8475,N_6181);
nand U13546 (N_13546,N_9819,N_6028);
and U13547 (N_13547,N_7630,N_9775);
nor U13548 (N_13548,N_7203,N_7118);
xor U13549 (N_13549,N_6933,N_9537);
and U13550 (N_13550,N_9849,N_7862);
nand U13551 (N_13551,N_9075,N_8664);
nand U13552 (N_13552,N_5348,N_5049);
or U13553 (N_13553,N_5727,N_6590);
or U13554 (N_13554,N_9222,N_7273);
or U13555 (N_13555,N_7875,N_7232);
or U13556 (N_13556,N_5249,N_9953);
nand U13557 (N_13557,N_5639,N_5736);
or U13558 (N_13558,N_6671,N_6372);
or U13559 (N_13559,N_6396,N_5909);
or U13560 (N_13560,N_7227,N_5093);
nand U13561 (N_13561,N_9232,N_7556);
nor U13562 (N_13562,N_9882,N_6942);
nor U13563 (N_13563,N_9736,N_7619);
nor U13564 (N_13564,N_7281,N_8770);
and U13565 (N_13565,N_5686,N_5585);
xnor U13566 (N_13566,N_5904,N_6001);
nand U13567 (N_13567,N_6677,N_8035);
nor U13568 (N_13568,N_6901,N_8300);
or U13569 (N_13569,N_6520,N_5249);
nand U13570 (N_13570,N_5465,N_9540);
and U13571 (N_13571,N_9234,N_9054);
nand U13572 (N_13572,N_8366,N_8017);
and U13573 (N_13573,N_9728,N_7011);
or U13574 (N_13574,N_5978,N_7608);
and U13575 (N_13575,N_5720,N_6367);
and U13576 (N_13576,N_9458,N_7608);
nand U13577 (N_13577,N_9087,N_5814);
and U13578 (N_13578,N_7389,N_5632);
or U13579 (N_13579,N_7980,N_5553);
and U13580 (N_13580,N_5287,N_6572);
nand U13581 (N_13581,N_8570,N_7107);
and U13582 (N_13582,N_5198,N_7950);
or U13583 (N_13583,N_7661,N_6331);
nor U13584 (N_13584,N_8888,N_6936);
nor U13585 (N_13585,N_7667,N_8077);
nor U13586 (N_13586,N_8000,N_5253);
nand U13587 (N_13587,N_6517,N_7947);
and U13588 (N_13588,N_8601,N_6505);
and U13589 (N_13589,N_6679,N_8344);
xor U13590 (N_13590,N_8615,N_8940);
or U13591 (N_13591,N_6598,N_6439);
and U13592 (N_13592,N_5059,N_9362);
or U13593 (N_13593,N_8604,N_9315);
nor U13594 (N_13594,N_5397,N_6044);
or U13595 (N_13595,N_6837,N_7816);
nand U13596 (N_13596,N_9339,N_5891);
or U13597 (N_13597,N_6436,N_8894);
xnor U13598 (N_13598,N_6605,N_6702);
xor U13599 (N_13599,N_6703,N_7197);
and U13600 (N_13600,N_9217,N_8136);
and U13601 (N_13601,N_5510,N_8024);
nand U13602 (N_13602,N_5641,N_8262);
or U13603 (N_13603,N_5952,N_9922);
and U13604 (N_13604,N_5861,N_9094);
nor U13605 (N_13605,N_9061,N_9892);
and U13606 (N_13606,N_7252,N_9251);
xor U13607 (N_13607,N_6550,N_9749);
and U13608 (N_13608,N_9500,N_5184);
nor U13609 (N_13609,N_6705,N_8431);
nor U13610 (N_13610,N_8038,N_9461);
nand U13611 (N_13611,N_7839,N_9572);
nand U13612 (N_13612,N_6682,N_6797);
or U13613 (N_13613,N_6204,N_5904);
or U13614 (N_13614,N_7988,N_8811);
nand U13615 (N_13615,N_5027,N_7642);
nor U13616 (N_13616,N_8065,N_6397);
nor U13617 (N_13617,N_7809,N_6661);
nor U13618 (N_13618,N_8394,N_7900);
or U13619 (N_13619,N_7302,N_8247);
nand U13620 (N_13620,N_5884,N_7131);
nor U13621 (N_13621,N_5134,N_6155);
and U13622 (N_13622,N_9360,N_7328);
nand U13623 (N_13623,N_9430,N_8403);
xor U13624 (N_13624,N_5607,N_8196);
and U13625 (N_13625,N_7044,N_8999);
or U13626 (N_13626,N_7858,N_6274);
or U13627 (N_13627,N_6131,N_5035);
xor U13628 (N_13628,N_6001,N_6122);
and U13629 (N_13629,N_5218,N_8037);
and U13630 (N_13630,N_8133,N_9779);
nand U13631 (N_13631,N_7164,N_7320);
or U13632 (N_13632,N_9369,N_8524);
or U13633 (N_13633,N_8712,N_8251);
nand U13634 (N_13634,N_5948,N_5387);
nand U13635 (N_13635,N_7167,N_8752);
and U13636 (N_13636,N_5442,N_8816);
xor U13637 (N_13637,N_9475,N_6966);
nand U13638 (N_13638,N_7767,N_6411);
or U13639 (N_13639,N_7416,N_5291);
nand U13640 (N_13640,N_5529,N_8247);
nand U13641 (N_13641,N_5495,N_7673);
nand U13642 (N_13642,N_9979,N_5441);
and U13643 (N_13643,N_5334,N_7018);
and U13644 (N_13644,N_5063,N_6852);
or U13645 (N_13645,N_9473,N_9230);
and U13646 (N_13646,N_6107,N_5707);
or U13647 (N_13647,N_5295,N_5737);
or U13648 (N_13648,N_8240,N_6308);
nor U13649 (N_13649,N_7768,N_5825);
nand U13650 (N_13650,N_5688,N_7893);
nand U13651 (N_13651,N_8249,N_9740);
nand U13652 (N_13652,N_6753,N_8705);
nor U13653 (N_13653,N_9758,N_5010);
xnor U13654 (N_13654,N_6479,N_9035);
nand U13655 (N_13655,N_5645,N_7722);
or U13656 (N_13656,N_9919,N_6462);
and U13657 (N_13657,N_6331,N_9057);
and U13658 (N_13658,N_6506,N_6676);
nand U13659 (N_13659,N_6190,N_7840);
or U13660 (N_13660,N_6576,N_8399);
nor U13661 (N_13661,N_9917,N_9326);
and U13662 (N_13662,N_9761,N_6762);
nor U13663 (N_13663,N_9056,N_8111);
or U13664 (N_13664,N_6382,N_7880);
nor U13665 (N_13665,N_6308,N_9229);
or U13666 (N_13666,N_9792,N_8604);
and U13667 (N_13667,N_8988,N_7756);
or U13668 (N_13668,N_6196,N_8798);
and U13669 (N_13669,N_6828,N_7879);
and U13670 (N_13670,N_9890,N_9277);
nand U13671 (N_13671,N_8405,N_5139);
or U13672 (N_13672,N_5486,N_9491);
nand U13673 (N_13673,N_7026,N_5430);
xor U13674 (N_13674,N_8954,N_6716);
nand U13675 (N_13675,N_8158,N_6598);
and U13676 (N_13676,N_7234,N_8590);
xor U13677 (N_13677,N_7249,N_6640);
and U13678 (N_13678,N_9631,N_8240);
or U13679 (N_13679,N_8691,N_9554);
or U13680 (N_13680,N_9657,N_5109);
and U13681 (N_13681,N_5733,N_7919);
nor U13682 (N_13682,N_5225,N_9031);
nand U13683 (N_13683,N_7857,N_5425);
and U13684 (N_13684,N_8391,N_5650);
xnor U13685 (N_13685,N_9313,N_6981);
nand U13686 (N_13686,N_7736,N_9068);
xnor U13687 (N_13687,N_8054,N_6485);
nor U13688 (N_13688,N_6571,N_8511);
xor U13689 (N_13689,N_8488,N_6480);
or U13690 (N_13690,N_7106,N_8940);
xnor U13691 (N_13691,N_5996,N_6754);
and U13692 (N_13692,N_9817,N_8209);
and U13693 (N_13693,N_5798,N_6566);
or U13694 (N_13694,N_7516,N_7332);
or U13695 (N_13695,N_6733,N_6314);
xnor U13696 (N_13696,N_6532,N_6754);
or U13697 (N_13697,N_5228,N_8686);
and U13698 (N_13698,N_9696,N_7133);
nand U13699 (N_13699,N_7558,N_7701);
and U13700 (N_13700,N_8163,N_6606);
and U13701 (N_13701,N_6134,N_8823);
nor U13702 (N_13702,N_7543,N_5275);
and U13703 (N_13703,N_8598,N_9315);
and U13704 (N_13704,N_6625,N_6707);
nand U13705 (N_13705,N_9149,N_5679);
or U13706 (N_13706,N_8100,N_6013);
nor U13707 (N_13707,N_6099,N_9354);
nand U13708 (N_13708,N_9345,N_7813);
or U13709 (N_13709,N_6836,N_8219);
and U13710 (N_13710,N_5296,N_5840);
and U13711 (N_13711,N_5319,N_6153);
and U13712 (N_13712,N_5715,N_5662);
xor U13713 (N_13713,N_7500,N_6160);
or U13714 (N_13714,N_7308,N_8314);
or U13715 (N_13715,N_8324,N_6954);
xor U13716 (N_13716,N_8708,N_9306);
nand U13717 (N_13717,N_9707,N_9314);
and U13718 (N_13718,N_6668,N_9837);
or U13719 (N_13719,N_8112,N_5213);
nand U13720 (N_13720,N_7956,N_5012);
and U13721 (N_13721,N_9211,N_7563);
or U13722 (N_13722,N_7976,N_9118);
or U13723 (N_13723,N_7269,N_7877);
xor U13724 (N_13724,N_9536,N_5321);
and U13725 (N_13725,N_8301,N_9934);
and U13726 (N_13726,N_5697,N_8335);
nor U13727 (N_13727,N_8930,N_7224);
nand U13728 (N_13728,N_6003,N_6486);
or U13729 (N_13729,N_8023,N_6285);
nand U13730 (N_13730,N_5009,N_5001);
nor U13731 (N_13731,N_8681,N_8206);
nor U13732 (N_13732,N_9602,N_8742);
or U13733 (N_13733,N_5259,N_8980);
nor U13734 (N_13734,N_6323,N_6820);
or U13735 (N_13735,N_7521,N_6643);
nor U13736 (N_13736,N_6051,N_6727);
or U13737 (N_13737,N_6107,N_9109);
nor U13738 (N_13738,N_5655,N_8094);
or U13739 (N_13739,N_7900,N_9088);
or U13740 (N_13740,N_9365,N_6614);
nor U13741 (N_13741,N_7899,N_7472);
and U13742 (N_13742,N_7048,N_6103);
nor U13743 (N_13743,N_5819,N_7209);
or U13744 (N_13744,N_7780,N_9202);
and U13745 (N_13745,N_9285,N_8010);
nor U13746 (N_13746,N_7583,N_7876);
or U13747 (N_13747,N_9615,N_7529);
nor U13748 (N_13748,N_9686,N_5993);
and U13749 (N_13749,N_7280,N_8004);
xor U13750 (N_13750,N_8827,N_6651);
nor U13751 (N_13751,N_9308,N_8265);
nor U13752 (N_13752,N_9768,N_7131);
nor U13753 (N_13753,N_7850,N_6054);
nor U13754 (N_13754,N_6315,N_5134);
nor U13755 (N_13755,N_9095,N_8362);
nor U13756 (N_13756,N_8244,N_7621);
or U13757 (N_13757,N_8925,N_7167);
nor U13758 (N_13758,N_9882,N_6479);
nor U13759 (N_13759,N_5650,N_7573);
and U13760 (N_13760,N_6012,N_8012);
and U13761 (N_13761,N_9211,N_9399);
nor U13762 (N_13762,N_8133,N_7357);
nor U13763 (N_13763,N_7535,N_5086);
nor U13764 (N_13764,N_5314,N_6394);
nand U13765 (N_13765,N_6865,N_6774);
or U13766 (N_13766,N_9240,N_8614);
xnor U13767 (N_13767,N_6146,N_9321);
and U13768 (N_13768,N_6844,N_7496);
nor U13769 (N_13769,N_6704,N_9624);
nor U13770 (N_13770,N_5216,N_7055);
and U13771 (N_13771,N_7710,N_8024);
nor U13772 (N_13772,N_9446,N_5731);
nor U13773 (N_13773,N_7734,N_7320);
nand U13774 (N_13774,N_8250,N_9023);
nor U13775 (N_13775,N_7657,N_9583);
nand U13776 (N_13776,N_8639,N_9615);
or U13777 (N_13777,N_8353,N_8656);
and U13778 (N_13778,N_8320,N_6353);
and U13779 (N_13779,N_8336,N_8958);
nor U13780 (N_13780,N_8945,N_5888);
nand U13781 (N_13781,N_6616,N_7751);
and U13782 (N_13782,N_7429,N_5868);
nand U13783 (N_13783,N_6322,N_8026);
or U13784 (N_13784,N_5479,N_7788);
nor U13785 (N_13785,N_8994,N_8720);
nand U13786 (N_13786,N_8908,N_9413);
nand U13787 (N_13787,N_6106,N_7475);
nand U13788 (N_13788,N_6453,N_8288);
nor U13789 (N_13789,N_8876,N_6900);
or U13790 (N_13790,N_7079,N_9611);
or U13791 (N_13791,N_6926,N_5999);
nand U13792 (N_13792,N_8225,N_9044);
nand U13793 (N_13793,N_8682,N_9673);
nor U13794 (N_13794,N_8834,N_9918);
nand U13795 (N_13795,N_6021,N_6026);
or U13796 (N_13796,N_7930,N_6186);
xor U13797 (N_13797,N_5797,N_5599);
or U13798 (N_13798,N_7718,N_9999);
nor U13799 (N_13799,N_6196,N_8500);
nor U13800 (N_13800,N_9712,N_7700);
nor U13801 (N_13801,N_6288,N_5346);
nor U13802 (N_13802,N_7288,N_8753);
or U13803 (N_13803,N_9761,N_9150);
and U13804 (N_13804,N_8059,N_7415);
nand U13805 (N_13805,N_6940,N_8974);
and U13806 (N_13806,N_6905,N_8169);
xor U13807 (N_13807,N_7555,N_7694);
nand U13808 (N_13808,N_6731,N_6505);
nand U13809 (N_13809,N_6435,N_9105);
nor U13810 (N_13810,N_7987,N_6359);
and U13811 (N_13811,N_6167,N_7306);
and U13812 (N_13812,N_6698,N_7741);
nand U13813 (N_13813,N_7591,N_6194);
and U13814 (N_13814,N_5370,N_5322);
and U13815 (N_13815,N_9058,N_5928);
xor U13816 (N_13816,N_7248,N_8808);
xor U13817 (N_13817,N_8693,N_9564);
xor U13818 (N_13818,N_8113,N_5281);
nand U13819 (N_13819,N_5589,N_9544);
or U13820 (N_13820,N_6716,N_5357);
or U13821 (N_13821,N_5743,N_8348);
nor U13822 (N_13822,N_8459,N_7335);
nor U13823 (N_13823,N_6658,N_5880);
and U13824 (N_13824,N_6404,N_5280);
nand U13825 (N_13825,N_8523,N_8125);
and U13826 (N_13826,N_9264,N_6738);
xnor U13827 (N_13827,N_9412,N_8091);
nor U13828 (N_13828,N_6362,N_5099);
nand U13829 (N_13829,N_7587,N_7408);
and U13830 (N_13830,N_9266,N_7279);
or U13831 (N_13831,N_8673,N_8425);
and U13832 (N_13832,N_6958,N_5928);
nor U13833 (N_13833,N_7202,N_6720);
xnor U13834 (N_13834,N_5940,N_7728);
and U13835 (N_13835,N_6315,N_5140);
or U13836 (N_13836,N_8286,N_9350);
nor U13837 (N_13837,N_6594,N_6244);
xnor U13838 (N_13838,N_6168,N_7142);
or U13839 (N_13839,N_9150,N_8711);
and U13840 (N_13840,N_9865,N_7030);
and U13841 (N_13841,N_7581,N_5745);
nor U13842 (N_13842,N_8512,N_7061);
nand U13843 (N_13843,N_8684,N_6250);
xnor U13844 (N_13844,N_8706,N_5339);
xnor U13845 (N_13845,N_7477,N_9630);
xnor U13846 (N_13846,N_5071,N_8793);
nand U13847 (N_13847,N_9337,N_6642);
nor U13848 (N_13848,N_6245,N_6200);
nand U13849 (N_13849,N_6629,N_9720);
xor U13850 (N_13850,N_7311,N_5335);
nand U13851 (N_13851,N_7123,N_8746);
xor U13852 (N_13852,N_9434,N_5545);
nand U13853 (N_13853,N_9575,N_7496);
nor U13854 (N_13854,N_9691,N_8499);
or U13855 (N_13855,N_7771,N_5141);
and U13856 (N_13856,N_7119,N_7881);
xnor U13857 (N_13857,N_8938,N_5343);
or U13858 (N_13858,N_5578,N_8469);
and U13859 (N_13859,N_7880,N_9774);
nor U13860 (N_13860,N_5260,N_7260);
nor U13861 (N_13861,N_9732,N_5015);
and U13862 (N_13862,N_6431,N_5811);
nor U13863 (N_13863,N_9512,N_8372);
nand U13864 (N_13864,N_5308,N_6067);
nor U13865 (N_13865,N_7116,N_9599);
nand U13866 (N_13866,N_9868,N_8099);
xnor U13867 (N_13867,N_7901,N_5844);
nor U13868 (N_13868,N_7677,N_8425);
or U13869 (N_13869,N_5384,N_6511);
or U13870 (N_13870,N_7513,N_7125);
or U13871 (N_13871,N_7950,N_9551);
nand U13872 (N_13872,N_5440,N_8594);
xnor U13873 (N_13873,N_6938,N_7893);
nand U13874 (N_13874,N_5554,N_7437);
nand U13875 (N_13875,N_6768,N_6623);
nand U13876 (N_13876,N_8659,N_7196);
or U13877 (N_13877,N_9412,N_7704);
nand U13878 (N_13878,N_6881,N_8556);
nor U13879 (N_13879,N_7608,N_5277);
and U13880 (N_13880,N_9792,N_6887);
and U13881 (N_13881,N_8638,N_8660);
or U13882 (N_13882,N_6216,N_9185);
and U13883 (N_13883,N_8639,N_7250);
and U13884 (N_13884,N_9077,N_7470);
nor U13885 (N_13885,N_8782,N_6986);
nand U13886 (N_13886,N_6550,N_7069);
nor U13887 (N_13887,N_5945,N_6609);
nor U13888 (N_13888,N_6537,N_5808);
nor U13889 (N_13889,N_6039,N_9877);
nor U13890 (N_13890,N_7891,N_5836);
and U13891 (N_13891,N_9091,N_9588);
or U13892 (N_13892,N_9546,N_7609);
or U13893 (N_13893,N_8947,N_8544);
or U13894 (N_13894,N_6028,N_5167);
nand U13895 (N_13895,N_9957,N_6273);
nor U13896 (N_13896,N_9387,N_8006);
nor U13897 (N_13897,N_7928,N_6435);
or U13898 (N_13898,N_6496,N_6774);
or U13899 (N_13899,N_5498,N_6005);
nand U13900 (N_13900,N_8551,N_7666);
or U13901 (N_13901,N_8841,N_9864);
xnor U13902 (N_13902,N_5037,N_9527);
nor U13903 (N_13903,N_8569,N_7198);
nor U13904 (N_13904,N_9865,N_9105);
xnor U13905 (N_13905,N_7767,N_7158);
or U13906 (N_13906,N_6055,N_6745);
nor U13907 (N_13907,N_6616,N_6977);
nor U13908 (N_13908,N_8317,N_9541);
nand U13909 (N_13909,N_6584,N_5518);
nand U13910 (N_13910,N_8776,N_7900);
nand U13911 (N_13911,N_5638,N_9465);
xor U13912 (N_13912,N_7188,N_8083);
nor U13913 (N_13913,N_5836,N_7628);
xnor U13914 (N_13914,N_6551,N_6848);
nor U13915 (N_13915,N_5217,N_8235);
or U13916 (N_13916,N_9602,N_8766);
or U13917 (N_13917,N_7149,N_9464);
xnor U13918 (N_13918,N_7476,N_8834);
xnor U13919 (N_13919,N_5981,N_6623);
and U13920 (N_13920,N_6478,N_8669);
and U13921 (N_13921,N_6008,N_6025);
and U13922 (N_13922,N_6635,N_7083);
nand U13923 (N_13923,N_5673,N_7716);
or U13924 (N_13924,N_5652,N_7036);
nand U13925 (N_13925,N_6039,N_6221);
nor U13926 (N_13926,N_8240,N_6621);
nor U13927 (N_13927,N_5616,N_7993);
or U13928 (N_13928,N_6685,N_7109);
nand U13929 (N_13929,N_6330,N_7683);
or U13930 (N_13930,N_5525,N_5201);
xnor U13931 (N_13931,N_6848,N_7405);
or U13932 (N_13932,N_7571,N_5277);
and U13933 (N_13933,N_6646,N_9973);
nand U13934 (N_13934,N_8263,N_8378);
or U13935 (N_13935,N_6119,N_7071);
and U13936 (N_13936,N_8614,N_7232);
or U13937 (N_13937,N_5273,N_7879);
nand U13938 (N_13938,N_9129,N_6931);
and U13939 (N_13939,N_9851,N_5635);
nand U13940 (N_13940,N_9510,N_6109);
nand U13941 (N_13941,N_6501,N_9355);
nand U13942 (N_13942,N_8378,N_8251);
and U13943 (N_13943,N_9741,N_7647);
nor U13944 (N_13944,N_8090,N_7321);
or U13945 (N_13945,N_6571,N_7852);
or U13946 (N_13946,N_8224,N_6258);
and U13947 (N_13947,N_7370,N_9549);
nor U13948 (N_13948,N_8621,N_6076);
nand U13949 (N_13949,N_5224,N_8046);
nor U13950 (N_13950,N_9653,N_8320);
xnor U13951 (N_13951,N_6744,N_9340);
and U13952 (N_13952,N_9053,N_5840);
nor U13953 (N_13953,N_5097,N_5453);
nor U13954 (N_13954,N_8488,N_7793);
nor U13955 (N_13955,N_8582,N_8550);
or U13956 (N_13956,N_7343,N_7409);
or U13957 (N_13957,N_7599,N_8713);
nor U13958 (N_13958,N_5047,N_9437);
nand U13959 (N_13959,N_5964,N_6117);
and U13960 (N_13960,N_6601,N_8258);
nor U13961 (N_13961,N_7956,N_8622);
nand U13962 (N_13962,N_9571,N_6516);
nor U13963 (N_13963,N_6387,N_6994);
nor U13964 (N_13964,N_9705,N_8051);
xor U13965 (N_13965,N_5255,N_5171);
nor U13966 (N_13966,N_9565,N_5664);
or U13967 (N_13967,N_6539,N_6046);
xor U13968 (N_13968,N_5959,N_6578);
nor U13969 (N_13969,N_8292,N_8759);
and U13970 (N_13970,N_9850,N_9826);
and U13971 (N_13971,N_5809,N_7797);
xnor U13972 (N_13972,N_6117,N_6109);
nor U13973 (N_13973,N_7344,N_8729);
nand U13974 (N_13974,N_6723,N_6832);
or U13975 (N_13975,N_5957,N_8827);
and U13976 (N_13976,N_6197,N_5663);
xnor U13977 (N_13977,N_6551,N_7063);
nor U13978 (N_13978,N_5954,N_7563);
nand U13979 (N_13979,N_8424,N_9170);
and U13980 (N_13980,N_9663,N_7363);
or U13981 (N_13981,N_7220,N_6981);
nand U13982 (N_13982,N_7641,N_7455);
xor U13983 (N_13983,N_8057,N_7452);
nor U13984 (N_13984,N_5872,N_8283);
nand U13985 (N_13985,N_9966,N_7279);
nand U13986 (N_13986,N_5584,N_8512);
nand U13987 (N_13987,N_7529,N_6046);
xor U13988 (N_13988,N_6145,N_9150);
or U13989 (N_13989,N_9502,N_8822);
nor U13990 (N_13990,N_7021,N_9196);
nor U13991 (N_13991,N_5632,N_8073);
nand U13992 (N_13992,N_9341,N_5769);
or U13993 (N_13993,N_9792,N_9719);
or U13994 (N_13994,N_7052,N_5507);
xnor U13995 (N_13995,N_7854,N_5321);
nor U13996 (N_13996,N_8312,N_7187);
nand U13997 (N_13997,N_7461,N_7159);
or U13998 (N_13998,N_9764,N_6588);
nand U13999 (N_13999,N_7977,N_8939);
xor U14000 (N_14000,N_9330,N_6719);
nand U14001 (N_14001,N_6219,N_9692);
nand U14002 (N_14002,N_9033,N_7200);
xor U14003 (N_14003,N_8460,N_6630);
and U14004 (N_14004,N_9675,N_7878);
or U14005 (N_14005,N_8804,N_9324);
nor U14006 (N_14006,N_5215,N_9303);
nand U14007 (N_14007,N_6618,N_5920);
nor U14008 (N_14008,N_5782,N_8997);
xnor U14009 (N_14009,N_6020,N_5544);
and U14010 (N_14010,N_8502,N_7488);
and U14011 (N_14011,N_8279,N_6995);
and U14012 (N_14012,N_5793,N_6832);
nor U14013 (N_14013,N_5466,N_8309);
and U14014 (N_14014,N_9210,N_5190);
nand U14015 (N_14015,N_6358,N_7152);
or U14016 (N_14016,N_6405,N_8808);
and U14017 (N_14017,N_6908,N_7075);
xor U14018 (N_14018,N_5526,N_7161);
nand U14019 (N_14019,N_6527,N_8552);
or U14020 (N_14020,N_5439,N_5868);
nor U14021 (N_14021,N_6095,N_7479);
xor U14022 (N_14022,N_6183,N_5100);
or U14023 (N_14023,N_7431,N_6164);
nor U14024 (N_14024,N_6801,N_8748);
nor U14025 (N_14025,N_5064,N_6085);
nand U14026 (N_14026,N_5239,N_7173);
or U14027 (N_14027,N_5160,N_5047);
or U14028 (N_14028,N_8274,N_7019);
nand U14029 (N_14029,N_5946,N_6120);
nor U14030 (N_14030,N_5900,N_9723);
and U14031 (N_14031,N_9211,N_9361);
nand U14032 (N_14032,N_7195,N_5416);
or U14033 (N_14033,N_6201,N_6974);
nor U14034 (N_14034,N_7533,N_5049);
nor U14035 (N_14035,N_5667,N_8174);
nand U14036 (N_14036,N_7691,N_6281);
and U14037 (N_14037,N_6454,N_5668);
and U14038 (N_14038,N_6933,N_9878);
nor U14039 (N_14039,N_9891,N_9782);
or U14040 (N_14040,N_6350,N_9472);
or U14041 (N_14041,N_9472,N_5922);
and U14042 (N_14042,N_5805,N_7690);
and U14043 (N_14043,N_7881,N_5204);
nor U14044 (N_14044,N_8243,N_6836);
nor U14045 (N_14045,N_6302,N_8189);
nor U14046 (N_14046,N_5821,N_5038);
or U14047 (N_14047,N_7245,N_8877);
and U14048 (N_14048,N_9204,N_8152);
nor U14049 (N_14049,N_7670,N_5691);
and U14050 (N_14050,N_5213,N_8048);
or U14051 (N_14051,N_6460,N_7383);
and U14052 (N_14052,N_5460,N_9193);
nand U14053 (N_14053,N_6514,N_5401);
nor U14054 (N_14054,N_6650,N_5995);
nand U14055 (N_14055,N_8605,N_6546);
and U14056 (N_14056,N_6039,N_7417);
and U14057 (N_14057,N_8446,N_7266);
nand U14058 (N_14058,N_9452,N_7701);
and U14059 (N_14059,N_6182,N_5175);
nor U14060 (N_14060,N_5407,N_9726);
or U14061 (N_14061,N_8647,N_7016);
and U14062 (N_14062,N_6823,N_5349);
or U14063 (N_14063,N_8362,N_5735);
nor U14064 (N_14064,N_8571,N_8708);
xnor U14065 (N_14065,N_9403,N_6558);
or U14066 (N_14066,N_9011,N_6915);
nor U14067 (N_14067,N_7501,N_7863);
and U14068 (N_14068,N_8702,N_6877);
and U14069 (N_14069,N_7341,N_9114);
or U14070 (N_14070,N_8310,N_8302);
nor U14071 (N_14071,N_9459,N_5291);
nor U14072 (N_14072,N_8547,N_7837);
and U14073 (N_14073,N_8421,N_5535);
nand U14074 (N_14074,N_9538,N_5183);
or U14075 (N_14075,N_6636,N_5062);
nand U14076 (N_14076,N_9947,N_9918);
or U14077 (N_14077,N_6832,N_7944);
or U14078 (N_14078,N_6330,N_9678);
nand U14079 (N_14079,N_9387,N_9528);
nand U14080 (N_14080,N_8444,N_5479);
nor U14081 (N_14081,N_7472,N_9092);
and U14082 (N_14082,N_9104,N_7910);
xnor U14083 (N_14083,N_7018,N_7921);
xor U14084 (N_14084,N_5630,N_9881);
and U14085 (N_14085,N_5753,N_5879);
nand U14086 (N_14086,N_9857,N_7769);
or U14087 (N_14087,N_7479,N_8323);
and U14088 (N_14088,N_6255,N_8645);
xor U14089 (N_14089,N_7517,N_6348);
xor U14090 (N_14090,N_6226,N_7858);
or U14091 (N_14091,N_9171,N_8060);
nand U14092 (N_14092,N_9912,N_9003);
xor U14093 (N_14093,N_8899,N_9679);
nor U14094 (N_14094,N_8809,N_9747);
nor U14095 (N_14095,N_6595,N_8807);
nor U14096 (N_14096,N_5827,N_7619);
or U14097 (N_14097,N_6612,N_5836);
and U14098 (N_14098,N_7072,N_6966);
nor U14099 (N_14099,N_9817,N_5043);
or U14100 (N_14100,N_6248,N_5796);
nand U14101 (N_14101,N_5427,N_6932);
and U14102 (N_14102,N_5046,N_5528);
or U14103 (N_14103,N_6695,N_7366);
or U14104 (N_14104,N_6347,N_9513);
or U14105 (N_14105,N_7875,N_5547);
or U14106 (N_14106,N_9449,N_9483);
nor U14107 (N_14107,N_5693,N_8386);
or U14108 (N_14108,N_7580,N_7095);
and U14109 (N_14109,N_8701,N_6067);
nor U14110 (N_14110,N_7999,N_8156);
and U14111 (N_14111,N_9334,N_8968);
nand U14112 (N_14112,N_8361,N_7962);
nand U14113 (N_14113,N_6808,N_6891);
and U14114 (N_14114,N_6027,N_5276);
nor U14115 (N_14115,N_6693,N_9064);
nor U14116 (N_14116,N_9791,N_8981);
nand U14117 (N_14117,N_7729,N_9502);
or U14118 (N_14118,N_9335,N_8775);
nand U14119 (N_14119,N_8449,N_6534);
nor U14120 (N_14120,N_7266,N_5794);
nor U14121 (N_14121,N_8666,N_9086);
nand U14122 (N_14122,N_7790,N_5814);
and U14123 (N_14123,N_6473,N_5646);
and U14124 (N_14124,N_9698,N_9020);
and U14125 (N_14125,N_7323,N_5736);
nor U14126 (N_14126,N_9540,N_7630);
nor U14127 (N_14127,N_8449,N_7581);
or U14128 (N_14128,N_7551,N_5443);
and U14129 (N_14129,N_9287,N_9443);
nor U14130 (N_14130,N_8710,N_7046);
xnor U14131 (N_14131,N_7193,N_6255);
nor U14132 (N_14132,N_8588,N_6352);
nor U14133 (N_14133,N_7243,N_5989);
nand U14134 (N_14134,N_9156,N_6170);
nor U14135 (N_14135,N_9586,N_6325);
nor U14136 (N_14136,N_6351,N_6565);
xor U14137 (N_14137,N_6785,N_8116);
or U14138 (N_14138,N_6275,N_5058);
nand U14139 (N_14139,N_6445,N_6526);
or U14140 (N_14140,N_6257,N_8685);
nor U14141 (N_14141,N_6292,N_6973);
nand U14142 (N_14142,N_5508,N_6457);
and U14143 (N_14143,N_6141,N_5916);
and U14144 (N_14144,N_7169,N_9765);
or U14145 (N_14145,N_6427,N_9799);
and U14146 (N_14146,N_6789,N_7370);
and U14147 (N_14147,N_6506,N_9933);
xor U14148 (N_14148,N_5853,N_7976);
or U14149 (N_14149,N_8057,N_9087);
nand U14150 (N_14150,N_7788,N_7179);
or U14151 (N_14151,N_6562,N_9238);
nor U14152 (N_14152,N_9217,N_6864);
and U14153 (N_14153,N_5069,N_5861);
nor U14154 (N_14154,N_7360,N_5027);
and U14155 (N_14155,N_5140,N_7686);
and U14156 (N_14156,N_6772,N_9560);
nand U14157 (N_14157,N_7655,N_8829);
and U14158 (N_14158,N_6877,N_9371);
nor U14159 (N_14159,N_6158,N_9127);
or U14160 (N_14160,N_7544,N_9794);
xor U14161 (N_14161,N_8187,N_7404);
xor U14162 (N_14162,N_7718,N_8055);
xor U14163 (N_14163,N_7344,N_8284);
nor U14164 (N_14164,N_7058,N_6612);
nand U14165 (N_14165,N_5890,N_8904);
nand U14166 (N_14166,N_9896,N_8813);
nor U14167 (N_14167,N_5211,N_5825);
or U14168 (N_14168,N_7245,N_8319);
xor U14169 (N_14169,N_5802,N_8793);
nor U14170 (N_14170,N_6050,N_6881);
nor U14171 (N_14171,N_6950,N_5074);
nor U14172 (N_14172,N_9164,N_7984);
nand U14173 (N_14173,N_8102,N_5356);
and U14174 (N_14174,N_5824,N_6166);
nand U14175 (N_14175,N_7200,N_6042);
or U14176 (N_14176,N_8482,N_8176);
and U14177 (N_14177,N_5220,N_5269);
nor U14178 (N_14178,N_7973,N_5004);
and U14179 (N_14179,N_5654,N_8389);
nand U14180 (N_14180,N_6905,N_5553);
nand U14181 (N_14181,N_7468,N_8439);
nand U14182 (N_14182,N_6715,N_5261);
nor U14183 (N_14183,N_9661,N_6815);
or U14184 (N_14184,N_9044,N_7475);
nand U14185 (N_14185,N_5559,N_7596);
nand U14186 (N_14186,N_8466,N_7488);
nand U14187 (N_14187,N_5690,N_7412);
nand U14188 (N_14188,N_9935,N_9934);
and U14189 (N_14189,N_6775,N_6412);
xnor U14190 (N_14190,N_6981,N_6626);
or U14191 (N_14191,N_6224,N_6589);
or U14192 (N_14192,N_9414,N_8233);
nand U14193 (N_14193,N_7720,N_6127);
nand U14194 (N_14194,N_8963,N_6743);
nand U14195 (N_14195,N_8681,N_9034);
nor U14196 (N_14196,N_6096,N_9206);
and U14197 (N_14197,N_9702,N_8652);
nor U14198 (N_14198,N_5644,N_8066);
nor U14199 (N_14199,N_6960,N_9272);
and U14200 (N_14200,N_6333,N_6702);
nor U14201 (N_14201,N_8181,N_5827);
and U14202 (N_14202,N_8904,N_8363);
or U14203 (N_14203,N_6792,N_6432);
or U14204 (N_14204,N_6354,N_9694);
nor U14205 (N_14205,N_9075,N_9923);
nor U14206 (N_14206,N_9065,N_5891);
nand U14207 (N_14207,N_8853,N_5424);
nor U14208 (N_14208,N_5138,N_8366);
nor U14209 (N_14209,N_6113,N_7647);
and U14210 (N_14210,N_7448,N_8829);
or U14211 (N_14211,N_7336,N_5372);
nor U14212 (N_14212,N_5967,N_7503);
or U14213 (N_14213,N_5609,N_6402);
nor U14214 (N_14214,N_7896,N_9814);
and U14215 (N_14215,N_8953,N_9603);
nor U14216 (N_14216,N_7439,N_8941);
and U14217 (N_14217,N_8292,N_8516);
nor U14218 (N_14218,N_5784,N_5641);
and U14219 (N_14219,N_8506,N_6880);
and U14220 (N_14220,N_5165,N_7403);
nand U14221 (N_14221,N_5959,N_5786);
nor U14222 (N_14222,N_5254,N_5029);
nor U14223 (N_14223,N_9865,N_9400);
nor U14224 (N_14224,N_5490,N_7040);
xor U14225 (N_14225,N_6845,N_5245);
or U14226 (N_14226,N_9930,N_5507);
nor U14227 (N_14227,N_5870,N_5519);
nor U14228 (N_14228,N_9171,N_5300);
and U14229 (N_14229,N_5252,N_6830);
nor U14230 (N_14230,N_5113,N_8729);
or U14231 (N_14231,N_8589,N_9017);
nand U14232 (N_14232,N_9531,N_9774);
xor U14233 (N_14233,N_6608,N_8608);
and U14234 (N_14234,N_6968,N_6414);
nor U14235 (N_14235,N_9223,N_6493);
nor U14236 (N_14236,N_9480,N_7665);
and U14237 (N_14237,N_8080,N_7350);
nor U14238 (N_14238,N_5783,N_8476);
nor U14239 (N_14239,N_9641,N_5491);
xnor U14240 (N_14240,N_8554,N_7517);
and U14241 (N_14241,N_8210,N_8423);
xnor U14242 (N_14242,N_7370,N_9668);
and U14243 (N_14243,N_6650,N_9242);
nor U14244 (N_14244,N_7808,N_8048);
and U14245 (N_14245,N_9922,N_5670);
nor U14246 (N_14246,N_6304,N_6725);
xor U14247 (N_14247,N_5207,N_5701);
and U14248 (N_14248,N_8745,N_9910);
nor U14249 (N_14249,N_7797,N_6038);
or U14250 (N_14250,N_7235,N_8135);
and U14251 (N_14251,N_8804,N_9153);
nand U14252 (N_14252,N_8467,N_7829);
and U14253 (N_14253,N_7469,N_9160);
xor U14254 (N_14254,N_7090,N_5082);
nor U14255 (N_14255,N_7237,N_7916);
nand U14256 (N_14256,N_6390,N_9805);
and U14257 (N_14257,N_6758,N_6235);
or U14258 (N_14258,N_8259,N_8812);
xnor U14259 (N_14259,N_7111,N_7706);
nand U14260 (N_14260,N_6862,N_5633);
and U14261 (N_14261,N_8543,N_9568);
nand U14262 (N_14262,N_9151,N_7609);
or U14263 (N_14263,N_8243,N_6967);
nor U14264 (N_14264,N_7841,N_9054);
and U14265 (N_14265,N_7318,N_7083);
nor U14266 (N_14266,N_5158,N_7674);
nand U14267 (N_14267,N_6537,N_9892);
nor U14268 (N_14268,N_6014,N_8060);
xnor U14269 (N_14269,N_8535,N_8974);
or U14270 (N_14270,N_8016,N_5917);
nor U14271 (N_14271,N_8691,N_6165);
and U14272 (N_14272,N_9097,N_7898);
xor U14273 (N_14273,N_8935,N_8711);
xor U14274 (N_14274,N_8251,N_8122);
or U14275 (N_14275,N_5012,N_6480);
nor U14276 (N_14276,N_6012,N_9034);
or U14277 (N_14277,N_5589,N_6024);
nand U14278 (N_14278,N_5311,N_8400);
or U14279 (N_14279,N_9585,N_7110);
and U14280 (N_14280,N_8830,N_8044);
or U14281 (N_14281,N_6374,N_5940);
xnor U14282 (N_14282,N_8477,N_9176);
and U14283 (N_14283,N_6504,N_5658);
xnor U14284 (N_14284,N_5255,N_9608);
or U14285 (N_14285,N_6100,N_8980);
and U14286 (N_14286,N_6309,N_8761);
and U14287 (N_14287,N_9806,N_9430);
or U14288 (N_14288,N_7051,N_6680);
nor U14289 (N_14289,N_5464,N_9131);
and U14290 (N_14290,N_6907,N_7702);
and U14291 (N_14291,N_8471,N_9928);
or U14292 (N_14292,N_8073,N_9966);
and U14293 (N_14293,N_5243,N_5672);
nand U14294 (N_14294,N_5468,N_6502);
and U14295 (N_14295,N_9786,N_9085);
or U14296 (N_14296,N_6390,N_8966);
or U14297 (N_14297,N_6119,N_5465);
or U14298 (N_14298,N_6911,N_9910);
and U14299 (N_14299,N_8629,N_5261);
and U14300 (N_14300,N_5014,N_8746);
and U14301 (N_14301,N_7941,N_8406);
nor U14302 (N_14302,N_9561,N_8622);
and U14303 (N_14303,N_5112,N_7238);
or U14304 (N_14304,N_9019,N_8496);
nand U14305 (N_14305,N_6722,N_6824);
or U14306 (N_14306,N_5174,N_9699);
or U14307 (N_14307,N_7514,N_5797);
and U14308 (N_14308,N_7930,N_6577);
or U14309 (N_14309,N_6403,N_5991);
or U14310 (N_14310,N_6731,N_8988);
nand U14311 (N_14311,N_9269,N_6203);
nor U14312 (N_14312,N_8634,N_8989);
xor U14313 (N_14313,N_6443,N_8472);
nand U14314 (N_14314,N_6464,N_9584);
xnor U14315 (N_14315,N_6141,N_6354);
and U14316 (N_14316,N_7187,N_9188);
or U14317 (N_14317,N_7551,N_5679);
nand U14318 (N_14318,N_8418,N_9588);
or U14319 (N_14319,N_8435,N_8723);
xor U14320 (N_14320,N_9203,N_9384);
nand U14321 (N_14321,N_7619,N_8264);
and U14322 (N_14322,N_7083,N_9638);
nand U14323 (N_14323,N_7114,N_9983);
nor U14324 (N_14324,N_7880,N_5046);
nand U14325 (N_14325,N_9496,N_7259);
and U14326 (N_14326,N_5258,N_7045);
nand U14327 (N_14327,N_7178,N_9874);
and U14328 (N_14328,N_9650,N_5282);
nand U14329 (N_14329,N_6761,N_6964);
nor U14330 (N_14330,N_9389,N_9858);
and U14331 (N_14331,N_7043,N_8507);
and U14332 (N_14332,N_7536,N_6533);
xnor U14333 (N_14333,N_7434,N_5655);
and U14334 (N_14334,N_9179,N_6630);
nand U14335 (N_14335,N_8713,N_5638);
or U14336 (N_14336,N_6400,N_6221);
or U14337 (N_14337,N_5161,N_9524);
nor U14338 (N_14338,N_6771,N_5825);
nor U14339 (N_14339,N_7474,N_6753);
or U14340 (N_14340,N_7708,N_8263);
nor U14341 (N_14341,N_7340,N_7111);
and U14342 (N_14342,N_9305,N_6413);
nand U14343 (N_14343,N_5482,N_7948);
nand U14344 (N_14344,N_9700,N_6782);
nand U14345 (N_14345,N_7051,N_8543);
nand U14346 (N_14346,N_7234,N_6616);
nand U14347 (N_14347,N_6065,N_5255);
or U14348 (N_14348,N_5564,N_5460);
or U14349 (N_14349,N_6231,N_8478);
and U14350 (N_14350,N_8224,N_5683);
nand U14351 (N_14351,N_6529,N_9128);
nand U14352 (N_14352,N_8479,N_9618);
and U14353 (N_14353,N_9791,N_6087);
nor U14354 (N_14354,N_7682,N_5936);
nor U14355 (N_14355,N_9439,N_7713);
nor U14356 (N_14356,N_7424,N_9515);
xnor U14357 (N_14357,N_8684,N_9127);
xor U14358 (N_14358,N_5413,N_8150);
and U14359 (N_14359,N_6931,N_7404);
or U14360 (N_14360,N_7267,N_8289);
and U14361 (N_14361,N_5423,N_7094);
nor U14362 (N_14362,N_7894,N_9138);
nor U14363 (N_14363,N_9868,N_7279);
and U14364 (N_14364,N_5061,N_7952);
or U14365 (N_14365,N_5154,N_8875);
nand U14366 (N_14366,N_9521,N_9686);
nor U14367 (N_14367,N_5475,N_7959);
nor U14368 (N_14368,N_7052,N_9405);
nor U14369 (N_14369,N_6643,N_6224);
xnor U14370 (N_14370,N_9674,N_5364);
or U14371 (N_14371,N_8519,N_9042);
xnor U14372 (N_14372,N_7411,N_7461);
and U14373 (N_14373,N_9051,N_8634);
nor U14374 (N_14374,N_7508,N_6758);
or U14375 (N_14375,N_9431,N_5872);
nand U14376 (N_14376,N_8004,N_5758);
or U14377 (N_14377,N_9750,N_7741);
or U14378 (N_14378,N_6521,N_9548);
nor U14379 (N_14379,N_9555,N_6228);
or U14380 (N_14380,N_9471,N_7759);
xor U14381 (N_14381,N_8088,N_6732);
nand U14382 (N_14382,N_6922,N_9471);
nand U14383 (N_14383,N_5924,N_9668);
and U14384 (N_14384,N_9901,N_6706);
nand U14385 (N_14385,N_8197,N_8127);
nor U14386 (N_14386,N_7545,N_7701);
xor U14387 (N_14387,N_6241,N_7510);
nor U14388 (N_14388,N_9724,N_7053);
nor U14389 (N_14389,N_5240,N_6918);
xor U14390 (N_14390,N_7026,N_7520);
or U14391 (N_14391,N_5209,N_8169);
nand U14392 (N_14392,N_5010,N_7620);
nand U14393 (N_14393,N_7902,N_5293);
nand U14394 (N_14394,N_8228,N_9378);
or U14395 (N_14395,N_5967,N_7193);
or U14396 (N_14396,N_5868,N_9894);
and U14397 (N_14397,N_5120,N_6167);
and U14398 (N_14398,N_9070,N_8706);
or U14399 (N_14399,N_7761,N_8939);
and U14400 (N_14400,N_5812,N_8163);
nor U14401 (N_14401,N_6965,N_5805);
nand U14402 (N_14402,N_9547,N_9916);
nor U14403 (N_14403,N_6379,N_8844);
nand U14404 (N_14404,N_6577,N_7776);
and U14405 (N_14405,N_5453,N_5971);
or U14406 (N_14406,N_6275,N_7741);
and U14407 (N_14407,N_5632,N_5168);
nand U14408 (N_14408,N_9835,N_5459);
xor U14409 (N_14409,N_8433,N_8948);
or U14410 (N_14410,N_8241,N_9870);
nor U14411 (N_14411,N_5153,N_8834);
nor U14412 (N_14412,N_9015,N_9768);
or U14413 (N_14413,N_9708,N_6325);
nand U14414 (N_14414,N_6697,N_6295);
nand U14415 (N_14415,N_5960,N_6125);
and U14416 (N_14416,N_6179,N_7037);
nand U14417 (N_14417,N_9592,N_5256);
or U14418 (N_14418,N_5504,N_5155);
or U14419 (N_14419,N_5999,N_7079);
and U14420 (N_14420,N_9331,N_8591);
nor U14421 (N_14421,N_8361,N_5649);
and U14422 (N_14422,N_7936,N_8616);
nor U14423 (N_14423,N_5386,N_6168);
and U14424 (N_14424,N_8383,N_7590);
or U14425 (N_14425,N_9505,N_6903);
or U14426 (N_14426,N_8780,N_5150);
nor U14427 (N_14427,N_8673,N_7777);
nand U14428 (N_14428,N_7134,N_9487);
or U14429 (N_14429,N_7711,N_8329);
nand U14430 (N_14430,N_6106,N_7432);
or U14431 (N_14431,N_8173,N_9933);
or U14432 (N_14432,N_6318,N_6444);
and U14433 (N_14433,N_8852,N_9053);
nor U14434 (N_14434,N_8443,N_9937);
or U14435 (N_14435,N_6858,N_7846);
or U14436 (N_14436,N_8808,N_9510);
nor U14437 (N_14437,N_5614,N_5139);
nand U14438 (N_14438,N_5272,N_5910);
xnor U14439 (N_14439,N_6084,N_5199);
and U14440 (N_14440,N_7513,N_9337);
nor U14441 (N_14441,N_8313,N_5805);
or U14442 (N_14442,N_7236,N_5704);
and U14443 (N_14443,N_5419,N_9116);
xor U14444 (N_14444,N_8857,N_9511);
nand U14445 (N_14445,N_9615,N_5410);
nand U14446 (N_14446,N_6987,N_8981);
or U14447 (N_14447,N_6603,N_6918);
or U14448 (N_14448,N_6783,N_9734);
nand U14449 (N_14449,N_6797,N_6305);
nor U14450 (N_14450,N_5766,N_6214);
xnor U14451 (N_14451,N_8567,N_6908);
nand U14452 (N_14452,N_9434,N_6929);
and U14453 (N_14453,N_9259,N_9482);
and U14454 (N_14454,N_5636,N_5368);
nor U14455 (N_14455,N_5296,N_9913);
or U14456 (N_14456,N_7001,N_6451);
nor U14457 (N_14457,N_5674,N_6270);
nand U14458 (N_14458,N_8259,N_8912);
nand U14459 (N_14459,N_8605,N_8670);
nand U14460 (N_14460,N_6278,N_7383);
and U14461 (N_14461,N_9623,N_8200);
nand U14462 (N_14462,N_8559,N_5682);
nand U14463 (N_14463,N_8143,N_6802);
and U14464 (N_14464,N_7163,N_6710);
or U14465 (N_14465,N_8694,N_6551);
and U14466 (N_14466,N_5425,N_7529);
nor U14467 (N_14467,N_8426,N_5614);
nor U14468 (N_14468,N_8512,N_6057);
nor U14469 (N_14469,N_5368,N_8432);
nor U14470 (N_14470,N_8582,N_8589);
nand U14471 (N_14471,N_7467,N_8155);
or U14472 (N_14472,N_6433,N_8135);
nand U14473 (N_14473,N_9951,N_7206);
nor U14474 (N_14474,N_6002,N_6086);
or U14475 (N_14475,N_9317,N_5369);
xnor U14476 (N_14476,N_5628,N_8395);
and U14477 (N_14477,N_8435,N_6681);
nor U14478 (N_14478,N_9434,N_6456);
and U14479 (N_14479,N_8261,N_6322);
nor U14480 (N_14480,N_5532,N_6173);
or U14481 (N_14481,N_8997,N_9425);
nor U14482 (N_14482,N_6484,N_6012);
nor U14483 (N_14483,N_7911,N_9815);
nor U14484 (N_14484,N_7464,N_5106);
and U14485 (N_14485,N_7072,N_9759);
and U14486 (N_14486,N_5122,N_5304);
or U14487 (N_14487,N_5283,N_8732);
nand U14488 (N_14488,N_6925,N_7040);
nand U14489 (N_14489,N_7848,N_8039);
or U14490 (N_14490,N_7427,N_8673);
or U14491 (N_14491,N_6877,N_9330);
nand U14492 (N_14492,N_5246,N_7707);
or U14493 (N_14493,N_8729,N_7716);
or U14494 (N_14494,N_8650,N_6766);
nand U14495 (N_14495,N_6241,N_6462);
and U14496 (N_14496,N_6301,N_9877);
nand U14497 (N_14497,N_6085,N_5634);
nor U14498 (N_14498,N_9816,N_7592);
nand U14499 (N_14499,N_9889,N_7134);
nor U14500 (N_14500,N_6361,N_5833);
or U14501 (N_14501,N_5706,N_9602);
and U14502 (N_14502,N_5256,N_6656);
or U14503 (N_14503,N_5400,N_8091);
and U14504 (N_14504,N_7058,N_8376);
and U14505 (N_14505,N_8613,N_7487);
or U14506 (N_14506,N_7150,N_7369);
nand U14507 (N_14507,N_7141,N_6074);
or U14508 (N_14508,N_5235,N_6666);
and U14509 (N_14509,N_7517,N_9045);
or U14510 (N_14510,N_6197,N_7735);
nand U14511 (N_14511,N_9733,N_8857);
or U14512 (N_14512,N_9796,N_8847);
and U14513 (N_14513,N_7991,N_6450);
or U14514 (N_14514,N_6400,N_5300);
nor U14515 (N_14515,N_8319,N_8154);
nand U14516 (N_14516,N_6800,N_7956);
nor U14517 (N_14517,N_5499,N_9570);
nor U14518 (N_14518,N_8579,N_7284);
and U14519 (N_14519,N_7360,N_7684);
nand U14520 (N_14520,N_7478,N_6388);
or U14521 (N_14521,N_9392,N_8750);
and U14522 (N_14522,N_5492,N_6082);
or U14523 (N_14523,N_6157,N_7501);
nand U14524 (N_14524,N_7824,N_6531);
or U14525 (N_14525,N_8181,N_9820);
nand U14526 (N_14526,N_8170,N_9706);
nor U14527 (N_14527,N_6759,N_9811);
and U14528 (N_14528,N_7752,N_7973);
or U14529 (N_14529,N_7443,N_6481);
or U14530 (N_14530,N_5997,N_8078);
or U14531 (N_14531,N_8782,N_8152);
nand U14532 (N_14532,N_8030,N_9905);
nand U14533 (N_14533,N_9711,N_7272);
nand U14534 (N_14534,N_5700,N_9371);
and U14535 (N_14535,N_7981,N_8042);
nand U14536 (N_14536,N_6717,N_5110);
nand U14537 (N_14537,N_8627,N_5897);
nor U14538 (N_14538,N_6807,N_7846);
or U14539 (N_14539,N_6094,N_7535);
or U14540 (N_14540,N_9927,N_7837);
and U14541 (N_14541,N_9780,N_8228);
nor U14542 (N_14542,N_9802,N_7996);
or U14543 (N_14543,N_9586,N_8024);
or U14544 (N_14544,N_8431,N_5001);
nor U14545 (N_14545,N_7718,N_9876);
or U14546 (N_14546,N_9085,N_6027);
nand U14547 (N_14547,N_9691,N_6729);
or U14548 (N_14548,N_5655,N_5719);
and U14549 (N_14549,N_7394,N_9696);
and U14550 (N_14550,N_8177,N_8278);
and U14551 (N_14551,N_7288,N_8371);
nor U14552 (N_14552,N_5499,N_8740);
xnor U14553 (N_14553,N_6883,N_6586);
nor U14554 (N_14554,N_7756,N_9496);
xnor U14555 (N_14555,N_9031,N_7858);
and U14556 (N_14556,N_9841,N_9133);
and U14557 (N_14557,N_7732,N_9503);
or U14558 (N_14558,N_8632,N_6055);
nor U14559 (N_14559,N_7752,N_6440);
xnor U14560 (N_14560,N_9240,N_5827);
nor U14561 (N_14561,N_7662,N_9400);
nand U14562 (N_14562,N_9934,N_8942);
nor U14563 (N_14563,N_9329,N_6239);
nor U14564 (N_14564,N_5928,N_5465);
nor U14565 (N_14565,N_5583,N_5532);
and U14566 (N_14566,N_7544,N_6148);
or U14567 (N_14567,N_5533,N_8521);
and U14568 (N_14568,N_8321,N_5198);
nand U14569 (N_14569,N_7509,N_8577);
xnor U14570 (N_14570,N_9719,N_5766);
nor U14571 (N_14571,N_8218,N_8114);
nand U14572 (N_14572,N_8520,N_9262);
and U14573 (N_14573,N_7474,N_6785);
xnor U14574 (N_14574,N_9597,N_6967);
nand U14575 (N_14575,N_9588,N_6650);
or U14576 (N_14576,N_5118,N_9317);
nor U14577 (N_14577,N_5490,N_5143);
nor U14578 (N_14578,N_9372,N_9403);
or U14579 (N_14579,N_7414,N_5161);
or U14580 (N_14580,N_8742,N_8909);
nand U14581 (N_14581,N_6667,N_7824);
xor U14582 (N_14582,N_9084,N_9667);
or U14583 (N_14583,N_8345,N_7928);
or U14584 (N_14584,N_8850,N_9722);
xor U14585 (N_14585,N_9471,N_9225);
and U14586 (N_14586,N_5918,N_6868);
or U14587 (N_14587,N_8631,N_6087);
nand U14588 (N_14588,N_9254,N_9247);
and U14589 (N_14589,N_5336,N_8100);
nand U14590 (N_14590,N_8315,N_9096);
nand U14591 (N_14591,N_8722,N_9375);
and U14592 (N_14592,N_6042,N_9515);
and U14593 (N_14593,N_8760,N_9251);
nand U14594 (N_14594,N_5326,N_7955);
nand U14595 (N_14595,N_8193,N_5041);
and U14596 (N_14596,N_8734,N_9741);
xor U14597 (N_14597,N_8652,N_8434);
or U14598 (N_14598,N_8103,N_9155);
or U14599 (N_14599,N_5160,N_7061);
and U14600 (N_14600,N_7802,N_6703);
nand U14601 (N_14601,N_7281,N_5801);
or U14602 (N_14602,N_5179,N_9227);
or U14603 (N_14603,N_5283,N_9946);
nand U14604 (N_14604,N_8100,N_7468);
nor U14605 (N_14605,N_6770,N_9115);
nand U14606 (N_14606,N_5993,N_8439);
and U14607 (N_14607,N_8504,N_9216);
or U14608 (N_14608,N_5029,N_8515);
or U14609 (N_14609,N_5295,N_6849);
and U14610 (N_14610,N_9474,N_5967);
and U14611 (N_14611,N_5731,N_5038);
or U14612 (N_14612,N_9531,N_8314);
and U14613 (N_14613,N_8760,N_9335);
or U14614 (N_14614,N_6219,N_7789);
nand U14615 (N_14615,N_8327,N_9707);
or U14616 (N_14616,N_7181,N_6863);
xnor U14617 (N_14617,N_7030,N_7196);
nor U14618 (N_14618,N_9530,N_8454);
and U14619 (N_14619,N_7771,N_7489);
and U14620 (N_14620,N_9207,N_9758);
nand U14621 (N_14621,N_7267,N_8641);
and U14622 (N_14622,N_8202,N_5210);
nor U14623 (N_14623,N_7718,N_6187);
or U14624 (N_14624,N_6640,N_6081);
nand U14625 (N_14625,N_7541,N_7346);
or U14626 (N_14626,N_6737,N_6257);
nor U14627 (N_14627,N_8865,N_9069);
nand U14628 (N_14628,N_5357,N_8939);
xnor U14629 (N_14629,N_6475,N_6248);
and U14630 (N_14630,N_9546,N_9188);
nand U14631 (N_14631,N_7741,N_7142);
nand U14632 (N_14632,N_5583,N_7504);
nand U14633 (N_14633,N_5921,N_8237);
or U14634 (N_14634,N_6214,N_9510);
nand U14635 (N_14635,N_9471,N_7120);
or U14636 (N_14636,N_8629,N_8808);
nand U14637 (N_14637,N_8614,N_9144);
and U14638 (N_14638,N_5440,N_7166);
nor U14639 (N_14639,N_8342,N_8276);
nor U14640 (N_14640,N_7729,N_5932);
nor U14641 (N_14641,N_9417,N_9234);
nand U14642 (N_14642,N_8627,N_8609);
or U14643 (N_14643,N_5813,N_5973);
nor U14644 (N_14644,N_6733,N_6020);
or U14645 (N_14645,N_8362,N_5411);
and U14646 (N_14646,N_8037,N_9727);
nor U14647 (N_14647,N_8164,N_5483);
nand U14648 (N_14648,N_9147,N_5828);
or U14649 (N_14649,N_7280,N_8683);
or U14650 (N_14650,N_5801,N_7032);
nor U14651 (N_14651,N_5930,N_8149);
or U14652 (N_14652,N_6435,N_5499);
nor U14653 (N_14653,N_6109,N_6371);
xor U14654 (N_14654,N_7379,N_7108);
and U14655 (N_14655,N_9426,N_7158);
and U14656 (N_14656,N_7656,N_7661);
nand U14657 (N_14657,N_8377,N_8386);
and U14658 (N_14658,N_5053,N_7222);
and U14659 (N_14659,N_5301,N_6264);
nand U14660 (N_14660,N_7171,N_6927);
and U14661 (N_14661,N_9427,N_9022);
xnor U14662 (N_14662,N_9933,N_6505);
and U14663 (N_14663,N_7415,N_7785);
xor U14664 (N_14664,N_6045,N_8743);
xor U14665 (N_14665,N_5516,N_6458);
or U14666 (N_14666,N_6931,N_5010);
and U14667 (N_14667,N_6302,N_5155);
and U14668 (N_14668,N_8597,N_5354);
or U14669 (N_14669,N_5842,N_6670);
nand U14670 (N_14670,N_6402,N_8804);
nand U14671 (N_14671,N_5152,N_6007);
nand U14672 (N_14672,N_8570,N_6788);
nand U14673 (N_14673,N_9665,N_9691);
nor U14674 (N_14674,N_5857,N_7228);
or U14675 (N_14675,N_6558,N_5496);
nor U14676 (N_14676,N_8284,N_8192);
or U14677 (N_14677,N_9419,N_8395);
and U14678 (N_14678,N_9926,N_5387);
nand U14679 (N_14679,N_7730,N_5702);
and U14680 (N_14680,N_9455,N_9166);
nor U14681 (N_14681,N_8142,N_7489);
and U14682 (N_14682,N_9457,N_5920);
or U14683 (N_14683,N_6527,N_6342);
nor U14684 (N_14684,N_8730,N_9858);
or U14685 (N_14685,N_8298,N_6076);
xnor U14686 (N_14686,N_6521,N_5166);
nand U14687 (N_14687,N_6394,N_6189);
or U14688 (N_14688,N_7062,N_5400);
and U14689 (N_14689,N_6883,N_9373);
xnor U14690 (N_14690,N_7821,N_8657);
nor U14691 (N_14691,N_8444,N_5681);
nor U14692 (N_14692,N_9821,N_6247);
and U14693 (N_14693,N_8428,N_9458);
xor U14694 (N_14694,N_9410,N_5916);
xnor U14695 (N_14695,N_8809,N_6056);
or U14696 (N_14696,N_6972,N_6767);
and U14697 (N_14697,N_8126,N_9598);
and U14698 (N_14698,N_5000,N_8110);
nand U14699 (N_14699,N_5224,N_5881);
nand U14700 (N_14700,N_9126,N_6734);
nand U14701 (N_14701,N_5252,N_6688);
or U14702 (N_14702,N_9494,N_9735);
and U14703 (N_14703,N_6136,N_5641);
nand U14704 (N_14704,N_6833,N_7108);
nor U14705 (N_14705,N_8589,N_7413);
xor U14706 (N_14706,N_5039,N_5453);
xnor U14707 (N_14707,N_8224,N_6951);
xor U14708 (N_14708,N_6748,N_6987);
and U14709 (N_14709,N_8518,N_5749);
or U14710 (N_14710,N_5540,N_6422);
or U14711 (N_14711,N_5502,N_9361);
and U14712 (N_14712,N_9741,N_7189);
or U14713 (N_14713,N_9545,N_8081);
or U14714 (N_14714,N_7093,N_8942);
xor U14715 (N_14715,N_9239,N_9123);
xor U14716 (N_14716,N_7753,N_8265);
nor U14717 (N_14717,N_9544,N_9865);
and U14718 (N_14718,N_7679,N_7995);
nand U14719 (N_14719,N_7085,N_7856);
and U14720 (N_14720,N_8534,N_8601);
and U14721 (N_14721,N_8258,N_9167);
xnor U14722 (N_14722,N_7499,N_7131);
nand U14723 (N_14723,N_6261,N_7831);
or U14724 (N_14724,N_9078,N_8315);
nor U14725 (N_14725,N_9447,N_9398);
and U14726 (N_14726,N_7167,N_8718);
nor U14727 (N_14727,N_8820,N_5478);
xnor U14728 (N_14728,N_8723,N_8919);
and U14729 (N_14729,N_9792,N_6453);
or U14730 (N_14730,N_9009,N_7840);
and U14731 (N_14731,N_9936,N_5788);
or U14732 (N_14732,N_6478,N_9276);
or U14733 (N_14733,N_9703,N_8564);
and U14734 (N_14734,N_5209,N_8868);
and U14735 (N_14735,N_7609,N_5979);
nor U14736 (N_14736,N_7877,N_8350);
nand U14737 (N_14737,N_6335,N_5222);
nor U14738 (N_14738,N_8694,N_5548);
or U14739 (N_14739,N_7658,N_6180);
nor U14740 (N_14740,N_9356,N_7418);
nor U14741 (N_14741,N_5103,N_7779);
nand U14742 (N_14742,N_9210,N_5942);
nor U14743 (N_14743,N_9270,N_8888);
or U14744 (N_14744,N_6522,N_8706);
nand U14745 (N_14745,N_8846,N_8069);
nor U14746 (N_14746,N_8038,N_5205);
nand U14747 (N_14747,N_6402,N_9097);
nor U14748 (N_14748,N_8692,N_6777);
nand U14749 (N_14749,N_7492,N_7283);
nand U14750 (N_14750,N_5259,N_9722);
xor U14751 (N_14751,N_5974,N_6786);
and U14752 (N_14752,N_5611,N_5762);
nor U14753 (N_14753,N_9513,N_5604);
or U14754 (N_14754,N_5353,N_8785);
or U14755 (N_14755,N_8654,N_8132);
nand U14756 (N_14756,N_7598,N_8380);
and U14757 (N_14757,N_8476,N_5396);
nand U14758 (N_14758,N_5950,N_5643);
or U14759 (N_14759,N_5886,N_7447);
nand U14760 (N_14760,N_6359,N_7780);
and U14761 (N_14761,N_7978,N_6833);
and U14762 (N_14762,N_5088,N_7461);
or U14763 (N_14763,N_9621,N_7403);
and U14764 (N_14764,N_8860,N_7324);
and U14765 (N_14765,N_9093,N_6903);
nand U14766 (N_14766,N_5423,N_6426);
or U14767 (N_14767,N_5146,N_5286);
nand U14768 (N_14768,N_5061,N_7234);
nor U14769 (N_14769,N_8053,N_7724);
and U14770 (N_14770,N_8950,N_8787);
nor U14771 (N_14771,N_6904,N_6253);
nor U14772 (N_14772,N_7095,N_6585);
nand U14773 (N_14773,N_7668,N_6786);
nand U14774 (N_14774,N_8706,N_6110);
or U14775 (N_14775,N_7561,N_5956);
nor U14776 (N_14776,N_9432,N_8397);
xnor U14777 (N_14777,N_9065,N_9884);
and U14778 (N_14778,N_5547,N_8774);
or U14779 (N_14779,N_8307,N_8318);
nor U14780 (N_14780,N_8296,N_5080);
nor U14781 (N_14781,N_5317,N_8830);
and U14782 (N_14782,N_6017,N_7005);
nand U14783 (N_14783,N_5939,N_8947);
or U14784 (N_14784,N_5140,N_8739);
or U14785 (N_14785,N_7510,N_8722);
or U14786 (N_14786,N_5612,N_8107);
xor U14787 (N_14787,N_7120,N_9942);
nor U14788 (N_14788,N_5294,N_8464);
xnor U14789 (N_14789,N_9686,N_5647);
nand U14790 (N_14790,N_8207,N_9379);
or U14791 (N_14791,N_8856,N_8750);
nor U14792 (N_14792,N_7133,N_6111);
or U14793 (N_14793,N_8415,N_5170);
nor U14794 (N_14794,N_9454,N_7052);
nor U14795 (N_14795,N_7485,N_6835);
nand U14796 (N_14796,N_8693,N_5153);
nor U14797 (N_14797,N_5878,N_9913);
nand U14798 (N_14798,N_9361,N_5734);
or U14799 (N_14799,N_8239,N_8484);
and U14800 (N_14800,N_6028,N_9390);
and U14801 (N_14801,N_9159,N_8556);
nor U14802 (N_14802,N_6828,N_6276);
nor U14803 (N_14803,N_5806,N_6633);
or U14804 (N_14804,N_5460,N_8148);
nor U14805 (N_14805,N_7172,N_9426);
or U14806 (N_14806,N_9340,N_9106);
or U14807 (N_14807,N_9005,N_7224);
nand U14808 (N_14808,N_8114,N_9813);
or U14809 (N_14809,N_6570,N_6518);
nand U14810 (N_14810,N_7087,N_9606);
xor U14811 (N_14811,N_9299,N_8727);
nor U14812 (N_14812,N_7407,N_7585);
nand U14813 (N_14813,N_9833,N_7300);
or U14814 (N_14814,N_9404,N_8790);
or U14815 (N_14815,N_6354,N_6383);
nor U14816 (N_14816,N_5454,N_8083);
xor U14817 (N_14817,N_8537,N_8585);
and U14818 (N_14818,N_6925,N_8234);
nor U14819 (N_14819,N_7037,N_8836);
nand U14820 (N_14820,N_5474,N_6918);
and U14821 (N_14821,N_6054,N_5253);
nand U14822 (N_14822,N_9921,N_7379);
or U14823 (N_14823,N_8540,N_5230);
xor U14824 (N_14824,N_7047,N_7304);
or U14825 (N_14825,N_8133,N_6902);
xnor U14826 (N_14826,N_8148,N_9660);
nor U14827 (N_14827,N_9953,N_8104);
nand U14828 (N_14828,N_9227,N_7897);
and U14829 (N_14829,N_6069,N_7628);
or U14830 (N_14830,N_7809,N_7647);
or U14831 (N_14831,N_6881,N_7176);
nand U14832 (N_14832,N_7234,N_5541);
nand U14833 (N_14833,N_8805,N_7479);
and U14834 (N_14834,N_5234,N_8067);
nor U14835 (N_14835,N_6458,N_8361);
nand U14836 (N_14836,N_9217,N_6689);
or U14837 (N_14837,N_5790,N_5410);
nor U14838 (N_14838,N_8357,N_8268);
and U14839 (N_14839,N_6951,N_6136);
or U14840 (N_14840,N_8549,N_7360);
nor U14841 (N_14841,N_9993,N_5652);
nor U14842 (N_14842,N_8641,N_7092);
xor U14843 (N_14843,N_7091,N_5860);
nor U14844 (N_14844,N_5340,N_9009);
and U14845 (N_14845,N_9547,N_8386);
nor U14846 (N_14846,N_5305,N_8403);
nor U14847 (N_14847,N_5240,N_8533);
and U14848 (N_14848,N_6352,N_7217);
xnor U14849 (N_14849,N_5184,N_8423);
xor U14850 (N_14850,N_5721,N_8251);
or U14851 (N_14851,N_7526,N_8452);
and U14852 (N_14852,N_7794,N_8531);
nand U14853 (N_14853,N_7886,N_7690);
and U14854 (N_14854,N_7834,N_6950);
or U14855 (N_14855,N_5141,N_5611);
xor U14856 (N_14856,N_7729,N_8948);
nor U14857 (N_14857,N_8230,N_8677);
xor U14858 (N_14858,N_9303,N_5106);
nand U14859 (N_14859,N_8505,N_8119);
and U14860 (N_14860,N_8592,N_8802);
nor U14861 (N_14861,N_9998,N_9248);
and U14862 (N_14862,N_6164,N_5055);
or U14863 (N_14863,N_6935,N_9442);
xnor U14864 (N_14864,N_5919,N_5298);
nor U14865 (N_14865,N_7441,N_6811);
and U14866 (N_14866,N_5948,N_5716);
nor U14867 (N_14867,N_5366,N_8235);
and U14868 (N_14868,N_6650,N_6296);
and U14869 (N_14869,N_7590,N_9113);
nand U14870 (N_14870,N_7107,N_6826);
nand U14871 (N_14871,N_5918,N_9426);
xnor U14872 (N_14872,N_5829,N_8538);
nor U14873 (N_14873,N_5936,N_8048);
nor U14874 (N_14874,N_7704,N_5493);
or U14875 (N_14875,N_7858,N_9571);
xnor U14876 (N_14876,N_9890,N_6226);
xor U14877 (N_14877,N_9964,N_8457);
nand U14878 (N_14878,N_5435,N_8219);
or U14879 (N_14879,N_8586,N_8190);
and U14880 (N_14880,N_7017,N_7334);
or U14881 (N_14881,N_8912,N_8507);
or U14882 (N_14882,N_6349,N_6625);
and U14883 (N_14883,N_7166,N_6087);
and U14884 (N_14884,N_6578,N_9654);
or U14885 (N_14885,N_6588,N_8173);
and U14886 (N_14886,N_8837,N_5779);
nor U14887 (N_14887,N_9512,N_9138);
or U14888 (N_14888,N_5796,N_6311);
or U14889 (N_14889,N_6022,N_7423);
xor U14890 (N_14890,N_9605,N_5618);
or U14891 (N_14891,N_6890,N_7975);
nand U14892 (N_14892,N_6218,N_6226);
and U14893 (N_14893,N_9190,N_8618);
or U14894 (N_14894,N_7780,N_8079);
nor U14895 (N_14895,N_7136,N_9302);
and U14896 (N_14896,N_8476,N_8429);
and U14897 (N_14897,N_9538,N_5403);
nand U14898 (N_14898,N_5589,N_8526);
or U14899 (N_14899,N_9831,N_6723);
nand U14900 (N_14900,N_6353,N_9939);
nor U14901 (N_14901,N_9734,N_8219);
nor U14902 (N_14902,N_5817,N_7801);
and U14903 (N_14903,N_5866,N_8110);
or U14904 (N_14904,N_5258,N_8445);
nor U14905 (N_14905,N_6248,N_5752);
xor U14906 (N_14906,N_8105,N_9035);
nor U14907 (N_14907,N_9736,N_6052);
nand U14908 (N_14908,N_9501,N_6144);
nand U14909 (N_14909,N_5212,N_9237);
nand U14910 (N_14910,N_8952,N_9764);
nor U14911 (N_14911,N_6761,N_6480);
nand U14912 (N_14912,N_9609,N_5516);
and U14913 (N_14913,N_9255,N_8568);
nor U14914 (N_14914,N_6670,N_6358);
and U14915 (N_14915,N_5817,N_5359);
and U14916 (N_14916,N_5989,N_9534);
nor U14917 (N_14917,N_7732,N_7229);
nand U14918 (N_14918,N_7883,N_5788);
or U14919 (N_14919,N_6926,N_9163);
nand U14920 (N_14920,N_7771,N_5309);
or U14921 (N_14921,N_9296,N_7943);
or U14922 (N_14922,N_5217,N_8773);
xor U14923 (N_14923,N_5973,N_9405);
or U14924 (N_14924,N_7671,N_6560);
and U14925 (N_14925,N_6844,N_8646);
and U14926 (N_14926,N_5436,N_8063);
nand U14927 (N_14927,N_7245,N_9807);
and U14928 (N_14928,N_6043,N_8236);
nor U14929 (N_14929,N_5762,N_6375);
and U14930 (N_14930,N_9359,N_7815);
nand U14931 (N_14931,N_5538,N_7486);
or U14932 (N_14932,N_5521,N_5179);
and U14933 (N_14933,N_7449,N_6084);
and U14934 (N_14934,N_8294,N_6488);
or U14935 (N_14935,N_8165,N_8784);
or U14936 (N_14936,N_8859,N_8845);
nor U14937 (N_14937,N_9100,N_6772);
nand U14938 (N_14938,N_6250,N_7393);
nor U14939 (N_14939,N_7651,N_8343);
or U14940 (N_14940,N_8940,N_6481);
or U14941 (N_14941,N_9208,N_8786);
and U14942 (N_14942,N_9228,N_8669);
or U14943 (N_14943,N_9879,N_5009);
nor U14944 (N_14944,N_6173,N_6655);
or U14945 (N_14945,N_9717,N_5956);
nor U14946 (N_14946,N_9418,N_5556);
or U14947 (N_14947,N_6794,N_7223);
nor U14948 (N_14948,N_9446,N_7743);
nand U14949 (N_14949,N_9621,N_7415);
xnor U14950 (N_14950,N_7236,N_8999);
nor U14951 (N_14951,N_6683,N_8551);
nand U14952 (N_14952,N_5255,N_6369);
nor U14953 (N_14953,N_8405,N_6413);
and U14954 (N_14954,N_9974,N_7352);
nor U14955 (N_14955,N_5988,N_8236);
and U14956 (N_14956,N_7169,N_7998);
nor U14957 (N_14957,N_6280,N_5613);
xnor U14958 (N_14958,N_9323,N_5089);
nand U14959 (N_14959,N_5552,N_6072);
nand U14960 (N_14960,N_8915,N_6506);
nand U14961 (N_14961,N_5528,N_8986);
nor U14962 (N_14962,N_6386,N_9220);
nand U14963 (N_14963,N_6820,N_8524);
nand U14964 (N_14964,N_5151,N_5635);
or U14965 (N_14965,N_6303,N_6541);
or U14966 (N_14966,N_7247,N_8096);
nor U14967 (N_14967,N_9530,N_8734);
nor U14968 (N_14968,N_8776,N_6748);
or U14969 (N_14969,N_9098,N_5759);
and U14970 (N_14970,N_8334,N_8545);
or U14971 (N_14971,N_5167,N_5131);
nor U14972 (N_14972,N_9480,N_6709);
nand U14973 (N_14973,N_6779,N_9558);
and U14974 (N_14974,N_9915,N_8408);
or U14975 (N_14975,N_9920,N_6206);
nor U14976 (N_14976,N_5553,N_7462);
nor U14977 (N_14977,N_7998,N_8087);
and U14978 (N_14978,N_7393,N_7460);
xor U14979 (N_14979,N_6942,N_9058);
or U14980 (N_14980,N_8037,N_8696);
nor U14981 (N_14981,N_6838,N_5676);
or U14982 (N_14982,N_6212,N_6179);
nor U14983 (N_14983,N_5405,N_9008);
and U14984 (N_14984,N_5734,N_9746);
nand U14985 (N_14985,N_5099,N_7154);
nand U14986 (N_14986,N_9823,N_9046);
and U14987 (N_14987,N_8462,N_9748);
xor U14988 (N_14988,N_6025,N_6609);
and U14989 (N_14989,N_7549,N_8232);
and U14990 (N_14990,N_9496,N_6519);
nor U14991 (N_14991,N_5874,N_5256);
and U14992 (N_14992,N_5970,N_7166);
and U14993 (N_14993,N_9212,N_5258);
or U14994 (N_14994,N_7463,N_9390);
or U14995 (N_14995,N_6017,N_5490);
nor U14996 (N_14996,N_8630,N_8909);
or U14997 (N_14997,N_5076,N_7062);
xnor U14998 (N_14998,N_8979,N_9208);
and U14999 (N_14999,N_8628,N_8718);
nand U15000 (N_15000,N_12242,N_10543);
nor U15001 (N_15001,N_12642,N_12864);
and U15002 (N_15002,N_14599,N_10713);
nor U15003 (N_15003,N_11966,N_11878);
or U15004 (N_15004,N_11594,N_13564);
and U15005 (N_15005,N_12883,N_13443);
and U15006 (N_15006,N_11865,N_12919);
nand U15007 (N_15007,N_14779,N_11434);
nor U15008 (N_15008,N_10773,N_11139);
and U15009 (N_15009,N_14640,N_10707);
nor U15010 (N_15010,N_12522,N_11922);
or U15011 (N_15011,N_12388,N_11032);
nor U15012 (N_15012,N_14787,N_12915);
or U15013 (N_15013,N_10509,N_11831);
or U15014 (N_15014,N_13297,N_10743);
nor U15015 (N_15015,N_14607,N_11274);
and U15016 (N_15016,N_12824,N_14688);
xor U15017 (N_15017,N_10994,N_14956);
nand U15018 (N_15018,N_11523,N_14212);
and U15019 (N_15019,N_11035,N_14389);
and U15020 (N_15020,N_13899,N_11088);
and U15021 (N_15021,N_10189,N_14782);
nor U15022 (N_15022,N_10558,N_14029);
or U15023 (N_15023,N_12782,N_13819);
or U15024 (N_15024,N_10031,N_11517);
nand U15025 (N_15025,N_13029,N_11826);
and U15026 (N_15026,N_13008,N_12934);
nor U15027 (N_15027,N_13292,N_10833);
and U15028 (N_15028,N_10961,N_10179);
xnor U15029 (N_15029,N_14143,N_12470);
xnor U15030 (N_15030,N_11267,N_14434);
nand U15031 (N_15031,N_14487,N_12145);
or U15032 (N_15032,N_11169,N_14246);
or U15033 (N_15033,N_11622,N_10537);
and U15034 (N_15034,N_14998,N_12385);
or U15035 (N_15035,N_11516,N_13694);
nor U15036 (N_15036,N_13365,N_12949);
nand U15037 (N_15037,N_11935,N_10075);
nand U15038 (N_15038,N_14197,N_14247);
and U15039 (N_15039,N_13605,N_10508);
or U15040 (N_15040,N_13797,N_10125);
nand U15041 (N_15041,N_10646,N_10751);
nor U15042 (N_15042,N_12423,N_13919);
or U15043 (N_15043,N_13254,N_10796);
and U15044 (N_15044,N_12087,N_11754);
and U15045 (N_15045,N_10856,N_13997);
nor U15046 (N_15046,N_10442,N_10182);
or U15047 (N_15047,N_14366,N_11583);
xnor U15048 (N_15048,N_14129,N_12384);
or U15049 (N_15049,N_10127,N_10056);
nor U15050 (N_15050,N_11307,N_14771);
nor U15051 (N_15051,N_11790,N_13743);
nand U15052 (N_15052,N_14381,N_14267);
nor U15053 (N_15053,N_14110,N_14077);
and U15054 (N_15054,N_10811,N_13717);
and U15055 (N_15055,N_13406,N_11546);
or U15056 (N_15056,N_13268,N_13712);
or U15057 (N_15057,N_12316,N_11219);
or U15058 (N_15058,N_12575,N_13649);
nand U15059 (N_15059,N_12537,N_14402);
or U15060 (N_15060,N_12201,N_10030);
and U15061 (N_15061,N_14822,N_13833);
nor U15062 (N_15062,N_13820,N_13534);
and U15063 (N_15063,N_12785,N_14061);
nor U15064 (N_15064,N_13862,N_14447);
or U15065 (N_15065,N_11627,N_10406);
xnor U15066 (N_15066,N_10494,N_14195);
nand U15067 (N_15067,N_12028,N_13053);
and U15068 (N_15068,N_14769,N_14756);
and U15069 (N_15069,N_14615,N_10403);
and U15070 (N_15070,N_10495,N_14325);
and U15071 (N_15071,N_11985,N_11052);
or U15072 (N_15072,N_14233,N_10821);
nor U15073 (N_15073,N_13135,N_12235);
nand U15074 (N_15074,N_14322,N_11655);
nor U15075 (N_15075,N_13229,N_12783);
nor U15076 (N_15076,N_11196,N_14758);
or U15077 (N_15077,N_12222,N_13674);
nand U15078 (N_15078,N_11941,N_12987);
and U15079 (N_15079,N_10648,N_14052);
xnor U15080 (N_15080,N_12539,N_12357);
and U15081 (N_15081,N_10855,N_13474);
and U15082 (N_15082,N_14650,N_11823);
or U15083 (N_15083,N_10105,N_13584);
and U15084 (N_15084,N_12136,N_11293);
nor U15085 (N_15085,N_10297,N_11575);
nor U15086 (N_15086,N_14789,N_11037);
nor U15087 (N_15087,N_11634,N_13464);
nor U15088 (N_15088,N_13956,N_10458);
nor U15089 (N_15089,N_14488,N_11156);
nand U15090 (N_15090,N_11202,N_11109);
nand U15091 (N_15091,N_14617,N_13173);
or U15092 (N_15092,N_10374,N_11694);
or U15093 (N_15093,N_12180,N_10376);
and U15094 (N_15094,N_12232,N_14836);
and U15095 (N_15095,N_11152,N_13682);
nand U15096 (N_15096,N_11953,N_11129);
nor U15097 (N_15097,N_12960,N_10151);
nor U15098 (N_15098,N_11449,N_11433);
nor U15099 (N_15099,N_10363,N_12627);
xnor U15100 (N_15100,N_11623,N_13115);
and U15101 (N_15101,N_11155,N_11715);
nand U15102 (N_15102,N_12431,N_11447);
and U15103 (N_15103,N_11319,N_10096);
nand U15104 (N_15104,N_12330,N_12464);
nand U15105 (N_15105,N_13739,N_10430);
nor U15106 (N_15106,N_12765,N_10906);
nor U15107 (N_15107,N_13400,N_12152);
and U15108 (N_15108,N_13015,N_11801);
nand U15109 (N_15109,N_10530,N_10121);
or U15110 (N_15110,N_11214,N_13526);
nand U15111 (N_15111,N_14042,N_14206);
nor U15112 (N_15112,N_11595,N_14625);
nand U15113 (N_15113,N_11301,N_14940);
nor U15114 (N_15114,N_11740,N_14275);
nand U15115 (N_15115,N_14271,N_10724);
or U15116 (N_15116,N_11412,N_11406);
xor U15117 (N_15117,N_11673,N_12014);
nor U15118 (N_15118,N_13275,N_11098);
nor U15119 (N_15119,N_12255,N_14657);
and U15120 (N_15120,N_12689,N_10378);
nor U15121 (N_15121,N_14123,N_13783);
and U15122 (N_15122,N_14482,N_13707);
and U15123 (N_15123,N_14125,N_12555);
nand U15124 (N_15124,N_14790,N_10071);
nor U15125 (N_15125,N_10557,N_11776);
nand U15126 (N_15126,N_13066,N_10476);
nor U15127 (N_15127,N_14065,N_14205);
nand U15128 (N_15128,N_13859,N_14258);
or U15129 (N_15129,N_14556,N_12270);
and U15130 (N_15130,N_11276,N_10827);
nand U15131 (N_15131,N_13886,N_14108);
nor U15132 (N_15132,N_12159,N_11228);
nand U15133 (N_15133,N_11311,N_14504);
and U15134 (N_15134,N_12612,N_13112);
or U15135 (N_15135,N_10319,N_11869);
xnor U15136 (N_15136,N_10969,N_11666);
nor U15137 (N_15137,N_11306,N_10489);
nor U15138 (N_15138,N_11289,N_12378);
or U15139 (N_15139,N_14598,N_10852);
and U15140 (N_15140,N_12490,N_13352);
xor U15141 (N_15141,N_12418,N_11193);
xnor U15142 (N_15142,N_11163,N_11074);
or U15143 (N_15143,N_14888,N_10902);
or U15144 (N_15144,N_11501,N_12216);
nand U15145 (N_15145,N_10138,N_12639);
or U15146 (N_15146,N_14418,N_10446);
and U15147 (N_15147,N_10365,N_10545);
or U15148 (N_15148,N_12476,N_12295);
nor U15149 (N_15149,N_14043,N_11678);
or U15150 (N_15150,N_13932,N_13439);
nand U15151 (N_15151,N_11668,N_13602);
and U15152 (N_15152,N_14364,N_10589);
and U15153 (N_15153,N_13647,N_13263);
and U15154 (N_15154,N_11153,N_12882);
xor U15155 (N_15155,N_13214,N_14412);
or U15156 (N_15156,N_12250,N_12991);
and U15157 (N_15157,N_14926,N_12404);
or U15158 (N_15158,N_11988,N_10695);
or U15159 (N_15159,N_14326,N_11252);
and U15160 (N_15160,N_14950,N_12358);
nor U15161 (N_15161,N_10418,N_14268);
nor U15162 (N_15162,N_13837,N_14965);
and U15163 (N_15163,N_10147,N_14387);
xnor U15164 (N_15164,N_13349,N_11427);
nor U15165 (N_15165,N_12871,N_13461);
and U15166 (N_15166,N_10413,N_10562);
or U15167 (N_15167,N_10130,N_14085);
nor U15168 (N_15168,N_11898,N_10627);
nor U15169 (N_15169,N_11134,N_11987);
xor U15170 (N_15170,N_14424,N_12684);
nor U15171 (N_15171,N_12995,N_13701);
or U15172 (N_15172,N_11648,N_12885);
nand U15173 (N_15173,N_14145,N_10060);
and U15174 (N_15174,N_10477,N_13855);
and U15175 (N_15175,N_11887,N_13508);
and U15176 (N_15176,N_12756,N_11933);
or U15177 (N_15177,N_10380,N_14928);
nor U15178 (N_15178,N_10612,N_10370);
or U15179 (N_15179,N_12015,N_14457);
and U15180 (N_15180,N_10128,N_12942);
and U15181 (N_15181,N_14055,N_14335);
nand U15182 (N_15182,N_14802,N_13442);
or U15183 (N_15183,N_14860,N_13742);
nand U15184 (N_15184,N_10340,N_11458);
xor U15185 (N_15185,N_13511,N_13721);
xnor U15186 (N_15186,N_12424,N_12382);
nor U15187 (N_15187,N_11533,N_12896);
and U15188 (N_15188,N_11361,N_13553);
and U15189 (N_15189,N_11264,N_13475);
nor U15190 (N_15190,N_10354,N_11029);
and U15191 (N_15191,N_14652,N_14338);
xor U15192 (N_15192,N_10131,N_11779);
or U15193 (N_15193,N_12862,N_11840);
nor U15194 (N_15194,N_14005,N_12692);
and U15195 (N_15195,N_14273,N_13497);
or U15196 (N_15196,N_12978,N_14603);
nor U15197 (N_15197,N_10234,N_14136);
and U15198 (N_15198,N_11797,N_10536);
xor U15199 (N_15199,N_14717,N_13054);
and U15200 (N_15200,N_14834,N_11907);
nand U15201 (N_15201,N_11856,N_14979);
or U15202 (N_15202,N_13928,N_13830);
nor U15203 (N_15203,N_10388,N_11625);
or U15204 (N_15204,N_10335,N_12694);
and U15205 (N_15205,N_14889,N_14220);
nand U15206 (N_15206,N_14721,N_10710);
and U15207 (N_15207,N_14153,N_13690);
and U15208 (N_15208,N_11934,N_13560);
and U15209 (N_15209,N_10146,N_10723);
and U15210 (N_15210,N_12870,N_10014);
and U15211 (N_15211,N_14303,N_12079);
nor U15212 (N_15212,N_11290,N_11036);
nor U15213 (N_15213,N_10824,N_13308);
xor U15214 (N_15214,N_11841,N_10565);
and U15215 (N_15215,N_10568,N_10775);
or U15216 (N_15216,N_11386,N_10638);
nand U15217 (N_15217,N_11184,N_14701);
nor U15218 (N_15218,N_11931,N_11068);
nand U15219 (N_15219,N_12195,N_11329);
nand U15220 (N_15220,N_13179,N_11158);
or U15221 (N_15221,N_11070,N_12602);
nand U15222 (N_15222,N_14353,N_14171);
or U15223 (N_15223,N_14528,N_12702);
or U15224 (N_15224,N_12772,N_12880);
and U15225 (N_15225,N_11631,N_13033);
xor U15226 (N_15226,N_12899,N_13389);
or U15227 (N_15227,N_11205,N_13834);
or U15228 (N_15228,N_11031,N_12593);
nand U15229 (N_15229,N_11705,N_14762);
nand U15230 (N_15230,N_12531,N_12737);
nand U15231 (N_15231,N_14886,N_13177);
and U15232 (N_15232,N_12840,N_10625);
and U15233 (N_15233,N_12711,N_11423);
and U15234 (N_15234,N_13084,N_11891);
and U15235 (N_15235,N_10745,N_12908);
nor U15236 (N_15236,N_10364,N_13273);
or U15237 (N_15237,N_14639,N_13800);
or U15238 (N_15238,N_13014,N_13515);
and U15239 (N_15239,N_10221,N_10350);
nand U15240 (N_15240,N_12691,N_11468);
or U15241 (N_15241,N_13217,N_11913);
nor U15242 (N_15242,N_11958,N_13462);
nand U15243 (N_15243,N_11519,N_11905);
nand U15244 (N_15244,N_14962,N_13999);
and U15245 (N_15245,N_12096,N_12874);
nor U15246 (N_15246,N_10945,N_14227);
nor U15247 (N_15247,N_12664,N_11954);
and U15248 (N_15248,N_14946,N_13924);
nor U15249 (N_15249,N_14374,N_10177);
nand U15250 (N_15250,N_11961,N_14058);
nand U15251 (N_15251,N_14677,N_13918);
nand U15252 (N_15252,N_11483,N_12320);
nand U15253 (N_15253,N_12116,N_12911);
or U15254 (N_15254,N_11246,N_12727);
nor U15255 (N_15255,N_10986,N_11313);
nor U15256 (N_15256,N_12563,N_13657);
or U15257 (N_15257,N_14296,N_12027);
nor U15258 (N_15258,N_10957,N_10581);
nand U15259 (N_15259,N_12724,N_11591);
nor U15260 (N_15260,N_13299,N_10661);
and U15261 (N_15261,N_11669,N_10339);
and U15262 (N_15262,N_12552,N_14653);
and U15263 (N_15263,N_10412,N_13518);
or U15264 (N_15264,N_10542,N_10830);
xnor U15265 (N_15265,N_12913,N_12178);
nand U15266 (N_15266,N_14416,N_11530);
and U15267 (N_15267,N_13608,N_13642);
or U15268 (N_15268,N_14551,N_10402);
and U15269 (N_15269,N_12102,N_11233);
or U15270 (N_15270,N_11885,N_10460);
nor U15271 (N_15271,N_12947,N_12381);
or U15272 (N_15272,N_10635,N_13887);
or U15273 (N_15273,N_10401,N_10260);
nand U15274 (N_15274,N_14839,N_13844);
nor U15275 (N_15275,N_14898,N_13525);
nand U15276 (N_15276,N_13946,N_14509);
nand U15277 (N_15277,N_13000,N_11771);
nand U15278 (N_15278,N_12472,N_13494);
or U15279 (N_15279,N_14942,N_10813);
xnor U15280 (N_15280,N_10432,N_11257);
nor U15281 (N_15281,N_14713,N_12266);
nand U15282 (N_15282,N_12721,N_10750);
nor U15283 (N_15283,N_10486,N_13197);
and U15284 (N_15284,N_14294,N_10787);
xnor U15285 (N_15285,N_10839,N_12997);
and U15286 (N_15286,N_13391,N_10324);
or U15287 (N_15287,N_10439,N_12802);
nor U15288 (N_15288,N_14433,N_13267);
and U15289 (N_15289,N_10577,N_11883);
nand U15290 (N_15290,N_10452,N_14229);
nand U15291 (N_15291,N_11963,N_13204);
and U15292 (N_15292,N_13902,N_10535);
nor U15293 (N_15293,N_12940,N_12543);
or U15294 (N_15294,N_12823,N_14327);
and U15295 (N_15295,N_14132,N_10045);
nand U15296 (N_15296,N_10689,N_10344);
or U15297 (N_15297,N_12615,N_10483);
nor U15298 (N_15298,N_13425,N_11662);
nand U15299 (N_15299,N_11154,N_11187);
or U15300 (N_15300,N_10999,N_10848);
nand U15301 (N_15301,N_13543,N_14156);
nand U15302 (N_15302,N_10355,N_14768);
nand U15303 (N_15303,N_11121,N_14534);
nand U15304 (N_15304,N_13333,N_12016);
xor U15305 (N_15305,N_12071,N_12925);
nor U15306 (N_15306,N_10600,N_14773);
xor U15307 (N_15307,N_11644,N_11316);
and U15308 (N_15308,N_14380,N_14211);
xor U15309 (N_15309,N_11309,N_14492);
nand U15310 (N_15310,N_14637,N_10893);
nor U15311 (N_15311,N_11380,N_10316);
and U15312 (N_15312,N_12077,N_12390);
or U15313 (N_15313,N_11957,N_11798);
nor U15314 (N_15314,N_11164,N_13858);
or U15315 (N_15315,N_10272,N_10454);
xnor U15316 (N_15316,N_12434,N_14936);
nand U15317 (N_15317,N_13710,N_14985);
nand U15318 (N_15318,N_12663,N_11294);
xnor U15319 (N_15319,N_12716,N_12117);
nand U15320 (N_15320,N_10399,N_10687);
and U15321 (N_15321,N_11632,N_10645);
nor U15322 (N_15322,N_10869,N_10069);
nand U15323 (N_15323,N_12483,N_10546);
and U15324 (N_15324,N_14250,N_11064);
or U15325 (N_15325,N_11189,N_14935);
nor U15326 (N_15326,N_11977,N_10939);
or U15327 (N_15327,N_12275,N_11227);
nor U15328 (N_15328,N_10907,N_11244);
and U15329 (N_15329,N_12749,N_11724);
and U15330 (N_15330,N_12514,N_13687);
and U15331 (N_15331,N_13253,N_12186);
nand U15332 (N_15332,N_12901,N_11166);
nor U15333 (N_15333,N_11105,N_12495);
nand U15334 (N_15334,N_13309,N_13099);
and U15335 (N_15335,N_11008,N_11752);
and U15336 (N_15336,N_14997,N_11171);
or U15337 (N_15337,N_12150,N_13424);
nor U15338 (N_15338,N_10461,N_13802);
and U15339 (N_15339,N_10634,N_13209);
or U15340 (N_15340,N_14214,N_14147);
or U15341 (N_15341,N_11493,N_13875);
nand U15342 (N_15342,N_10580,N_11221);
and U15343 (N_15343,N_11675,N_11401);
xnor U15344 (N_15344,N_12900,N_12393);
and U15345 (N_15345,N_14215,N_14170);
nor U15346 (N_15346,N_12905,N_12668);
and U15347 (N_15347,N_11521,N_13818);
nand U15348 (N_15348,N_12536,N_10865);
nand U15349 (N_15349,N_12304,N_14964);
nor U15350 (N_15350,N_13983,N_13157);
nor U15351 (N_15351,N_14245,N_10526);
nor U15352 (N_15352,N_12518,N_10041);
or U15353 (N_15353,N_12876,N_11364);
nand U15354 (N_15354,N_12392,N_14018);
nand U15355 (N_15355,N_12832,N_14319);
nand U15356 (N_15356,N_12810,N_10944);
nor U15357 (N_15357,N_12241,N_11653);
nand U15358 (N_15358,N_12355,N_10341);
nand U15359 (N_15359,N_10033,N_14328);
and U15360 (N_15360,N_13206,N_12482);
nand U15361 (N_15361,N_13122,N_13213);
and U15362 (N_15362,N_11371,N_11471);
and U15363 (N_15363,N_10591,N_11821);
xnor U15364 (N_15364,N_13676,N_11304);
nor U15365 (N_15365,N_12857,N_13043);
nor U15366 (N_15366,N_14814,N_12811);
or U15367 (N_15367,N_11002,N_14198);
and U15368 (N_15368,N_12115,N_14112);
nor U15369 (N_15369,N_12520,N_12594);
nor U15370 (N_15370,N_14696,N_10874);
nor U15371 (N_15371,N_10306,N_10931);
or U15372 (N_15372,N_12535,N_11038);
or U15373 (N_15373,N_12533,N_12521);
nor U15374 (N_15374,N_14765,N_14700);
nor U15375 (N_15375,N_13372,N_14672);
and U15376 (N_15376,N_12352,N_14954);
and U15377 (N_15377,N_14098,N_13144);
or U15378 (N_15378,N_13939,N_12155);
xnor U15379 (N_15379,N_10506,N_11286);
or U15380 (N_15380,N_14667,N_11281);
and U15381 (N_15381,N_10913,N_13361);
nand U15382 (N_15382,N_11350,N_14081);
and U15383 (N_15383,N_11700,N_13745);
and U15384 (N_15384,N_12970,N_13388);
nand U15385 (N_15385,N_10000,N_10064);
or U15386 (N_15386,N_10815,N_13554);
and U15387 (N_15387,N_11356,N_11084);
nand U15388 (N_15388,N_14941,N_13555);
or U15389 (N_15389,N_10076,N_11415);
or U15390 (N_15390,N_14261,N_12825);
nand U15391 (N_15391,N_14920,N_13387);
nand U15392 (N_15392,N_14025,N_12957);
nor U15393 (N_15393,N_11525,N_11866);
nor U15394 (N_15394,N_14394,N_14276);
or U15395 (N_15395,N_14122,N_10704);
nor U15396 (N_15396,N_13706,N_13485);
and U15397 (N_15397,N_13900,N_14991);
nor U15398 (N_15398,N_10866,N_14589);
nand U15399 (N_15399,N_10357,N_11515);
nor U15400 (N_15400,N_11201,N_11637);
or U15401 (N_15401,N_13139,N_14320);
xnor U15402 (N_15402,N_12127,N_12084);
nand U15403 (N_15403,N_10933,N_14225);
nor U15404 (N_15404,N_13644,N_11455);
nand U15405 (N_15405,N_14722,N_13082);
or U15406 (N_15406,N_13629,N_10150);
nand U15407 (N_15407,N_10731,N_10631);
xnor U15408 (N_15408,N_11145,N_12236);
or U15409 (N_15409,N_11762,N_13162);
or U15410 (N_15410,N_13930,N_10078);
and U15411 (N_15411,N_11333,N_14291);
and U15412 (N_15412,N_10711,N_10954);
or U15413 (N_15413,N_10622,N_14537);
or U15414 (N_15414,N_12524,N_12787);
nor U15415 (N_15415,N_12920,N_12784);
nor U15416 (N_15416,N_13113,N_12974);
xor U15417 (N_15417,N_14073,N_11976);
nor U15418 (N_15418,N_10681,N_11854);
and U15419 (N_15419,N_13416,N_12654);
and U15420 (N_15420,N_14629,N_13108);
nor U15421 (N_15421,N_14097,N_13149);
or U15422 (N_15422,N_10397,N_11643);
or U15423 (N_15423,N_13154,N_10888);
nor U15424 (N_15424,N_13619,N_11903);
xor U15425 (N_15425,N_14035,N_12829);
nand U15426 (N_15426,N_12414,N_14877);
nor U15427 (N_15427,N_10674,N_13342);
nor U15428 (N_15428,N_10936,N_10163);
nor U15429 (N_15429,N_13470,N_11410);
and U15430 (N_15430,N_13995,N_14500);
or U15431 (N_15431,N_12842,N_14620);
and U15432 (N_15432,N_12137,N_12188);
nand U15433 (N_15433,N_11279,N_12288);
xnor U15434 (N_15434,N_12487,N_11803);
nand U15435 (N_15435,N_11749,N_12826);
or U15436 (N_15436,N_10529,N_12872);
nand U15437 (N_15437,N_13377,N_10223);
nand U15438 (N_15438,N_13936,N_12572);
xor U15439 (N_15439,N_13714,N_12151);
or U15440 (N_15440,N_14350,N_11352);
and U15441 (N_15441,N_14907,N_14148);
and U15442 (N_15442,N_13131,N_13062);
or U15443 (N_15443,N_12119,N_11486);
xor U15444 (N_15444,N_11460,N_12626);
xor U15445 (N_15445,N_11747,N_11432);
nor U15446 (N_15446,N_14744,N_11871);
xor U15447 (N_15447,N_11900,N_10062);
and U15448 (N_15448,N_10336,N_10420);
nand U15449 (N_15449,N_12494,N_14601);
or U15450 (N_15450,N_10513,N_10479);
and U15451 (N_15451,N_11945,N_11204);
and U15452 (N_15452,N_10298,N_13246);
and U15453 (N_15453,N_13224,N_11241);
nor U15454 (N_15454,N_14689,N_13138);
or U15455 (N_15455,N_10794,N_12374);
nor U15456 (N_15456,N_10104,N_14235);
and U15457 (N_15457,N_12111,N_11843);
and U15458 (N_15458,N_13021,N_13677);
nand U15459 (N_15459,N_12379,N_10285);
xnor U15460 (N_15460,N_13295,N_13522);
nor U15461 (N_15461,N_12803,N_14107);
nor U15462 (N_15462,N_12794,N_10135);
nand U15463 (N_15463,N_10549,N_12364);
xnor U15464 (N_15464,N_13252,N_12394);
nor U15465 (N_15465,N_13659,N_13615);
nand U15466 (N_15466,N_13760,N_11972);
xnor U15467 (N_15467,N_12283,N_11978);
nand U15468 (N_15468,N_13272,N_11091);
and U15469 (N_15469,N_10482,N_12939);
nor U15470 (N_15470,N_10665,N_12109);
nand U15471 (N_15471,N_11962,N_13392);
nand U15472 (N_15472,N_14332,N_13166);
and U15473 (N_15473,N_11118,N_14003);
nand U15474 (N_15474,N_11490,N_12503);
and U15475 (N_15475,N_12979,N_11853);
or U15476 (N_15476,N_10682,N_14514);
and U15477 (N_15477,N_14764,N_12026);
nand U15478 (N_15478,N_11721,N_14925);
and U15479 (N_15479,N_10518,N_10466);
nor U15480 (N_15480,N_10253,N_14916);
or U15481 (N_15481,N_11407,N_14893);
or U15482 (N_15482,N_10192,N_12103);
nor U15483 (N_15483,N_10853,N_10292);
nor U15484 (N_15484,N_13093,N_13630);
nand U15485 (N_15485,N_11365,N_10585);
nor U15486 (N_15486,N_14086,N_12187);
or U15487 (N_15487,N_13842,N_14938);
and U15488 (N_15488,N_14159,N_12946);
xor U15489 (N_15489,N_10312,N_14630);
and U15490 (N_15490,N_14967,N_10161);
and U15491 (N_15491,N_14642,N_11811);
nor U15492 (N_15492,N_12886,N_10684);
xor U15493 (N_15493,N_14567,N_14352);
and U15494 (N_15494,N_14346,N_10919);
and U15495 (N_15495,N_11473,N_11599);
or U15496 (N_15496,N_14833,N_14955);
nand U15497 (N_15497,N_10735,N_14673);
or U15498 (N_15498,N_11082,N_14649);
and U15499 (N_15499,N_12921,N_10755);
or U15500 (N_15500,N_12750,N_10571);
xnor U15501 (N_15501,N_13289,N_10431);
and U15502 (N_15502,N_13190,N_10693);
xor U15503 (N_15503,N_14177,N_11693);
or U15504 (N_15504,N_10327,N_14062);
nand U15505 (N_15505,N_11278,N_12958);
and U15506 (N_15506,N_13145,N_14638);
or U15507 (N_15507,N_14518,N_12163);
nand U15508 (N_15508,N_12439,N_14697);
xor U15509 (N_15509,N_13410,N_12944);
or U15510 (N_15510,N_11175,N_10662);
and U15511 (N_15511,N_12133,N_13850);
or U15512 (N_15512,N_12945,N_11691);
nor U15513 (N_15513,N_10699,N_11973);
nor U15514 (N_15514,N_12313,N_13168);
xnor U15515 (N_15515,N_13772,N_10434);
xnor U15516 (N_15516,N_11734,N_10438);
or U15517 (N_15517,N_13814,N_11053);
nor U15518 (N_15518,N_13719,N_11711);
nand U15519 (N_15519,N_13925,N_12816);
nand U15520 (N_15520,N_10847,N_14747);
xnor U15521 (N_15521,N_10762,N_10663);
or U15522 (N_15522,N_12461,N_13734);
nor U15523 (N_15523,N_11565,N_14376);
or U15524 (N_15524,N_13729,N_13434);
nand U15525 (N_15525,N_13169,N_11641);
and U15526 (N_15526,N_10587,N_11127);
nor U15527 (N_15527,N_10108,N_11714);
or U15528 (N_15528,N_10770,N_14391);
and U15529 (N_15529,N_10023,N_10985);
nand U15530 (N_15530,N_14851,N_11851);
xnor U15531 (N_15531,N_14566,N_10720);
nand U15532 (N_15532,N_12298,N_10632);
xnor U15533 (N_15533,N_12637,N_12373);
or U15534 (N_15534,N_11026,N_14825);
nand U15535 (N_15535,N_14176,N_10098);
nor U15536 (N_15536,N_12805,N_14919);
xnor U15537 (N_15537,N_11272,N_11788);
or U15538 (N_15538,N_10791,N_11199);
or U15539 (N_15539,N_11028,N_11377);
nor U15540 (N_15540,N_12890,N_13907);
or U15541 (N_15541,N_11937,N_12184);
and U15542 (N_15542,N_11069,N_11019);
nand U15543 (N_15543,N_10763,N_13836);
and U15544 (N_15544,N_12516,N_10300);
or U15545 (N_15545,N_13781,N_11096);
nand U15546 (N_15546,N_13514,N_14435);
and U15547 (N_15547,N_11378,N_10222);
nand U15548 (N_15548,N_12259,N_13708);
nor U15549 (N_15549,N_14903,N_11079);
nor U15550 (N_15550,N_12203,N_11938);
or U15551 (N_15551,N_11424,N_10233);
nor U15552 (N_15552,N_12739,N_11782);
nand U15553 (N_15553,N_14983,N_13822);
or U15554 (N_15554,N_14659,N_12875);
nor U15555 (N_15555,N_13368,N_14579);
or U15556 (N_15556,N_10026,N_10923);
xnor U15557 (N_15557,N_10455,N_14587);
or U15558 (N_15558,N_12072,N_12812);
nor U15559 (N_15559,N_11908,N_13123);
and U15560 (N_15560,N_12475,N_14783);
xor U15561 (N_15561,N_13869,N_13612);
or U15562 (N_15562,N_14797,N_11054);
nand U15563 (N_15563,N_10754,N_13503);
or U15564 (N_15564,N_14723,N_14251);
or U15565 (N_15565,N_13792,N_12820);
nor U15566 (N_15566,N_11465,N_13579);
or U15567 (N_15567,N_14869,N_10828);
nand U15568 (N_15568,N_13556,N_11162);
nand U15569 (N_15569,N_13110,N_10840);
xor U15570 (N_15570,N_10410,N_14716);
nand U15571 (N_15571,N_11925,N_14614);
xnor U15572 (N_15572,N_13240,N_14707);
xor U15573 (N_15573,N_10169,N_13375);
nand U15574 (N_15574,N_13187,N_11536);
or U15575 (N_15575,N_10882,N_10911);
nor U15576 (N_15576,N_12768,N_13698);
xnor U15577 (N_15577,N_11131,N_13769);
or U15578 (N_15578,N_10946,N_11670);
and U15579 (N_15579,N_11774,N_12906);
nand U15580 (N_15580,N_12693,N_12606);
xor U15581 (N_15581,N_11690,N_11814);
nand U15582 (N_15582,N_12808,N_14952);
or U15583 (N_15583,N_11100,N_12931);
nand U15584 (N_15584,N_13271,N_11149);
nand U15585 (N_15585,N_10757,N_10216);
or U15586 (N_15586,N_12338,N_11126);
nor U15587 (N_15587,N_13089,N_10262);
and U15588 (N_15588,N_14980,N_12780);
or U15589 (N_15589,N_13358,N_10426);
and U15590 (N_15590,N_11360,N_11789);
or U15591 (N_15591,N_11807,N_10967);
nor U15592 (N_15592,N_13741,N_11943);
nor U15593 (N_15593,N_11766,N_11505);
and U15594 (N_15594,N_10917,N_12311);
nand U15595 (N_15595,N_14896,N_12511);
nor U15596 (N_15596,N_10774,N_13165);
and U15597 (N_15597,N_12179,N_13521);
and U15598 (N_15598,N_10926,N_12988);
nand U15599 (N_15599,N_13210,N_12881);
xnor U15600 (N_15600,N_13460,N_10552);
and U15601 (N_15601,N_14499,N_12923);
xnor U15602 (N_15602,N_10894,N_10955);
nor U15603 (N_15603,N_14815,N_13756);
and U15604 (N_15604,N_10531,N_10569);
and U15605 (N_15605,N_14648,N_12197);
and U15606 (N_15606,N_10052,N_13109);
nand U15607 (N_15607,N_10450,N_13095);
nand U15608 (N_15608,N_10572,N_10883);
and U15609 (N_15609,N_12359,N_11800);
xnor U15610 (N_15610,N_12713,N_14188);
xnor U15611 (N_15611,N_13408,N_14027);
or U15612 (N_15612,N_12795,N_12598);
nor U15613 (N_15613,N_12831,N_13990);
nand U15614 (N_15614,N_14423,N_14463);
and U15615 (N_15615,N_12801,N_11255);
or U15616 (N_15616,N_12181,N_12744);
nor U15617 (N_15617,N_10443,N_13988);
and U15618 (N_15618,N_10550,N_10705);
nor U15619 (N_15619,N_14008,N_10218);
nand U15620 (N_15620,N_13864,N_10798);
nand U15621 (N_15621,N_13637,N_11825);
or U15622 (N_15622,N_11722,N_13628);
nor U15623 (N_15623,N_11395,N_12300);
and U15624 (N_15624,N_13727,N_12858);
xnor U15625 (N_15625,N_13074,N_14585);
nand U15626 (N_15626,N_10671,N_14014);
xor U15627 (N_15627,N_12492,N_10633);
nor U15628 (N_15628,N_13293,N_12929);
nor U15629 (N_15629,N_10845,N_12786);
nor U15630 (N_15630,N_11579,N_13433);
nand U15631 (N_15631,N_12859,N_11075);
nor U15632 (N_15632,N_12686,N_12057);
xor U15633 (N_15633,N_12401,N_11042);
and U15634 (N_15634,N_12892,N_14185);
or U15635 (N_15635,N_10929,N_10072);
nand U15636 (N_15636,N_13790,N_10666);
nor U15637 (N_15637,N_13957,N_12760);
or U15638 (N_15638,N_10035,N_12608);
and U15639 (N_15639,N_12146,N_10502);
and U15640 (N_15640,N_11946,N_14977);
nor U15641 (N_15641,N_14680,N_13171);
nand U15642 (N_15642,N_11051,N_14420);
or U15643 (N_15643,N_10993,N_14984);
nor U15644 (N_15644,N_10748,N_14187);
or U15645 (N_15645,N_12326,N_11297);
nor U15646 (N_15646,N_11507,N_14887);
or U15647 (N_15647,N_11436,N_10602);
nand U15648 (N_15648,N_13558,N_13613);
and U15649 (N_15649,N_13037,N_11367);
nor U15650 (N_15650,N_11218,N_13551);
nand U15651 (N_15651,N_14236,N_11769);
and U15652 (N_15652,N_14610,N_10063);
or U15653 (N_15653,N_11004,N_12416);
or U15654 (N_15654,N_14910,N_13780);
and U15655 (N_15655,N_13696,N_13343);
or U15656 (N_15656,N_10347,N_10099);
nand U15657 (N_15657,N_12659,N_10293);
nor U15658 (N_15658,N_13380,N_14856);
nand U15659 (N_15659,N_11582,N_10892);
and U15660 (N_15660,N_14260,N_14189);
nand U15661 (N_15661,N_10042,N_13873);
or U15662 (N_15662,N_14994,N_14671);
or U15663 (N_15663,N_14921,N_12198);
nand U15664 (N_15664,N_13334,N_13467);
nor U15665 (N_15665,N_13689,N_14024);
or U15666 (N_15666,N_10889,N_12666);
nand U15667 (N_15667,N_11404,N_12771);
xor U15668 (N_15668,N_13473,N_12585);
and U15669 (N_15669,N_13782,N_11593);
nand U15670 (N_15670,N_13044,N_14777);
nand U15671 (N_15671,N_10353,N_12956);
and U15672 (N_15672,N_11614,N_12688);
nand U15673 (N_15673,N_10155,N_11451);
or U15674 (N_15674,N_14571,N_13282);
nor U15675 (N_15675,N_13175,N_11667);
nand U15676 (N_15676,N_13072,N_12441);
xor U15677 (N_15677,N_13301,N_10283);
or U15678 (N_15678,N_12459,N_13378);
xnor U15679 (N_15679,N_14811,N_14957);
or U15680 (N_15680,N_12284,N_12775);
or U15681 (N_15681,N_10564,N_12099);
xnor U15682 (N_15682,N_11431,N_13746);
xnor U15683 (N_15683,N_10044,N_10077);
nor U15684 (N_15684,N_13290,N_10448);
nand U15685 (N_15685,N_11442,N_11422);
nand U15686 (N_15686,N_13685,N_11093);
or U15687 (N_15687,N_12170,N_10212);
nor U15688 (N_15688,N_11538,N_10555);
xnor U15689 (N_15689,N_10520,N_12294);
or U15690 (N_15690,N_11229,N_13422);
nand U15691 (N_15691,N_13950,N_14682);
xor U15692 (N_15692,N_14874,N_13269);
or U15693 (N_15693,N_11366,N_12329);
nor U15694 (N_15694,N_13397,N_14109);
nand U15695 (N_15695,N_12809,N_13167);
nand U15696 (N_15696,N_11860,N_14739);
nand U15697 (N_15697,N_10084,N_13680);
nand U15698 (N_15698,N_13549,N_11062);
or U15699 (N_15699,N_14662,N_12336);
nor U15700 (N_15700,N_13603,N_14853);
nand U15701 (N_15701,N_14915,N_12806);
xor U15702 (N_15702,N_13303,N_14719);
nand U15703 (N_15703,N_14969,N_12963);
nand U15704 (N_15704,N_10820,N_10470);
nand U15705 (N_15705,N_10899,N_13453);
or U15706 (N_15706,N_11537,N_13901);
xor U15707 (N_15707,N_11503,N_13151);
nor U15708 (N_15708,N_10369,N_11877);
xnor U15709 (N_15709,N_13386,N_14026);
nor U15710 (N_15710,N_14686,N_13247);
nand U15711 (N_15711,N_13523,N_10029);
nand U15712 (N_15712,N_12599,N_14542);
nor U15713 (N_15713,N_13793,N_12292);
xnor U15714 (N_15714,N_10228,N_12339);
nor U15715 (N_15715,N_13330,N_13759);
and U15716 (N_15716,N_12916,N_13182);
xnor U15717 (N_15717,N_12411,N_12733);
nor U15718 (N_15718,N_14623,N_11191);
xor U15719 (N_15719,N_10090,N_12860);
and U15720 (N_15720,N_11999,N_11926);
or U15721 (N_15721,N_12354,N_14628);
nor U15722 (N_15722,N_11775,N_13816);
and U15723 (N_15723,N_12559,N_11894);
nand U15724 (N_15724,N_14793,N_10842);
nor U15725 (N_15725,N_12632,N_11334);
nor U15726 (N_15726,N_11485,N_13141);
and U15727 (N_15727,N_11209,N_13256);
or U15728 (N_15728,N_13218,N_14362);
xor U15729 (N_15729,N_10680,N_11492);
or U15730 (N_15730,N_12767,N_14039);
and U15731 (N_15731,N_14624,N_10895);
nand U15732 (N_15732,N_10139,N_10752);
nand U15733 (N_15733,N_11712,N_14805);
nand U15734 (N_15734,N_13005,N_13223);
and U15735 (N_15735,N_12030,N_13251);
nor U15736 (N_15736,N_14367,N_13038);
nand U15737 (N_15737,N_11245,N_11650);
nand U15738 (N_15738,N_10080,N_10213);
nor U15739 (N_15739,N_14681,N_13770);
or U15740 (N_15740,N_10019,N_12499);
nor U15741 (N_15741,N_14971,N_11370);
or U15742 (N_15742,N_13949,N_14495);
or U15743 (N_15743,N_10831,N_11013);
nand U15744 (N_15744,N_10254,N_12504);
nand U15745 (N_15745,N_10359,N_14612);
or U15746 (N_15746,N_12403,N_12985);
xnor U15747 (N_15747,N_12687,N_12898);
nor U15748 (N_15748,N_14754,N_14978);
or U15749 (N_15749,N_14804,N_13587);
nor U15750 (N_15750,N_14297,N_10259);
nor U15751 (N_15751,N_14490,N_12821);
nor U15752 (N_15752,N_10238,N_10055);
xor U15753 (N_15753,N_13180,N_14759);
and U15754 (N_15754,N_10349,N_12398);
nand U15755 (N_15755,N_10047,N_10230);
nand U15756 (N_15756,N_12081,N_11951);
nand U15757 (N_15757,N_13183,N_10965);
and U15758 (N_15758,N_11578,N_13673);
xnor U15759 (N_15759,N_14219,N_12722);
or U15760 (N_15760,N_14613,N_14767);
nor U15761 (N_15761,N_14485,N_12479);
and U15762 (N_15762,N_12777,N_10626);
xnor U15763 (N_15763,N_11960,N_10657);
and U15764 (N_15764,N_13843,N_11968);
or U15765 (N_15765,N_10497,N_13048);
nor U15766 (N_15766,N_12032,N_14507);
nand U15767 (N_15767,N_12493,N_12369);
xnor U15768 (N_15768,N_10858,N_11750);
and U15769 (N_15769,N_13028,N_11466);
or U15770 (N_15770,N_11628,N_14728);
nor U15771 (N_15771,N_10930,N_13607);
nor U15772 (N_15772,N_10516,N_12169);
nand U15773 (N_15773,N_13102,N_11238);
or U15774 (N_15774,N_13100,N_14895);
nand U15775 (N_15775,N_12271,N_14059);
and U15776 (N_15776,N_12258,N_11640);
or U15777 (N_15777,N_14807,N_14191);
xnor U15778 (N_15778,N_13845,N_13367);
and U15779 (N_15779,N_13402,N_12208);
or U15780 (N_15780,N_14788,N_12532);
nand U15781 (N_15781,N_11130,N_13625);
nor U15782 (N_15782,N_10901,N_12397);
nor U15783 (N_15783,N_13910,N_11833);
and U15784 (N_15784,N_11902,N_11018);
nand U15785 (N_15785,N_14604,N_12971);
and U15786 (N_15786,N_10709,N_14501);
nor U15787 (N_15787,N_13471,N_10039);
or U15788 (N_15788,N_10018,N_10091);
nor U15789 (N_15789,N_10166,N_12021);
nor U15790 (N_15790,N_10922,N_13969);
nand U15791 (N_15791,N_14780,N_11608);
nand U15792 (N_15792,N_13915,N_14987);
nand U15793 (N_15793,N_13888,N_10148);
nand U15794 (N_15794,N_13117,N_11930);
or U15795 (N_15795,N_10785,N_12229);
and U15796 (N_15796,N_14845,N_12661);
or U15797 (N_15797,N_14203,N_12725);
nand U15798 (N_15798,N_10079,N_13982);
and U15799 (N_15799,N_11730,N_13385);
or U15800 (N_15800,N_14150,N_10143);
and U15801 (N_15801,N_12773,N_13944);
xor U15802 (N_15802,N_13040,N_12590);
nand U15803 (N_15803,N_11760,N_13896);
or U15804 (N_15804,N_13895,N_14524);
or U15805 (N_15805,N_11413,N_13789);
or U15806 (N_15806,N_14806,N_13500);
nand U15807 (N_15807,N_13948,N_12243);
nand U15808 (N_15808,N_11190,N_10346);
nand U15809 (N_15809,N_12730,N_12205);
or U15810 (N_15810,N_10377,N_12177);
and U15811 (N_15811,N_10067,N_10366);
or U15812 (N_15812,N_12544,N_14208);
nor U15813 (N_15813,N_14302,N_14255);
and U15814 (N_15814,N_12796,N_11007);
nand U15815 (N_15815,N_13627,N_10241);
xnor U15816 (N_15816,N_14193,N_14175);
and U15817 (N_15817,N_14298,N_12123);
or U15818 (N_15818,N_10948,N_13221);
xor U15819 (N_15819,N_13921,N_13614);
nand U15820 (N_15820,N_10025,N_12707);
and U15821 (N_15821,N_11123,N_10226);
nor U15822 (N_15822,N_14264,N_11464);
xor U15823 (N_15823,N_13513,N_11729);
and U15824 (N_15824,N_12049,N_12869);
nor U15825 (N_15825,N_13512,N_11893);
and U15826 (N_15826,N_12981,N_11733);
or U15827 (N_15827,N_11499,N_14196);
nor U15828 (N_15828,N_11997,N_10621);
and U15829 (N_15829,N_14540,N_14473);
and U15830 (N_15830,N_13401,N_12219);
nor U15831 (N_15831,N_13787,N_11200);
xor U15832 (N_15832,N_12943,N_11924);
nand U15833 (N_15833,N_10333,N_13312);
nand U15834 (N_15834,N_10053,N_13310);
and U15835 (N_15835,N_11083,N_10123);
or U15836 (N_15836,N_14040,N_10912);
nor U15837 (N_15837,N_12849,N_11596);
nand U15838 (N_15838,N_13242,N_13283);
and U15839 (N_15839,N_11959,N_11261);
nand U15840 (N_15840,N_12589,N_12568);
xor U15841 (N_15841,N_14092,N_12176);
and U15842 (N_15842,N_10252,N_14437);
or U15843 (N_15843,N_10616,N_10057);
and U15844 (N_15844,N_10291,N_13863);
xnor U15845 (N_15845,N_13912,N_11243);
nor U15846 (N_15846,N_10741,N_10953);
or U15847 (N_15847,N_12630,N_13118);
nand U15848 (N_15848,N_10758,N_12566);
nor U15849 (N_15849,N_14301,N_12223);
and U15850 (N_15850,N_11225,N_10844);
and U15851 (N_15851,N_12887,N_14742);
or U15852 (N_15852,N_10204,N_12315);
nor U15853 (N_15853,N_14323,N_12105);
nor U15854 (N_15854,N_10599,N_12265);
nor U15855 (N_15855,N_11102,N_14036);
or U15856 (N_15856,N_14349,N_13370);
or U15857 (N_15857,N_10541,N_14285);
nand U15858 (N_15858,N_11699,N_13848);
nand U15859 (N_15859,N_13019,N_12868);
xnor U15860 (N_15860,N_10698,N_11258);
and U15861 (N_15861,N_12800,N_10387);
and U15862 (N_15862,N_13496,N_12634);
nand U15863 (N_15863,N_12529,N_13345);
or U15864 (N_15864,N_11986,N_11741);
nand U15865 (N_15865,N_12221,N_13753);
or U15866 (N_15866,N_10609,N_10049);
and U15867 (N_15867,N_14685,N_10769);
and U15868 (N_15868,N_14242,N_11580);
nand U15869 (N_15869,N_14114,N_13632);
nand U15870 (N_15870,N_10214,N_11382);
or U15871 (N_15871,N_13011,N_14737);
or U15872 (N_15872,N_12955,N_11115);
and U15873 (N_15873,N_11544,N_12556);
or U15874 (N_15874,N_10517,N_12878);
and U15875 (N_15875,N_10037,N_14377);
nand U15876 (N_15876,N_14119,N_13531);
and U15877 (N_15877,N_11146,N_10947);
nor U15878 (N_15878,N_13479,N_14861);
and U15879 (N_15879,N_10396,N_14115);
or U15880 (N_15880,N_12211,N_13052);
or U15881 (N_15881,N_13591,N_14130);
nand U15882 (N_15882,N_14001,N_12833);
nand U15883 (N_15883,N_14970,N_13758);
and U15884 (N_15884,N_10659,N_12282);
and U15885 (N_15885,N_11868,N_10407);
and U15886 (N_15886,N_13762,N_12484);
or U15887 (N_15887,N_13056,N_11336);
nor U15888 (N_15888,N_10287,N_14778);
or U15889 (N_15889,N_10284,N_10582);
xnor U15890 (N_15890,N_14329,N_14660);
or U15891 (N_15891,N_11511,N_14382);
or U15892 (N_15892,N_12427,N_12445);
or U15893 (N_15893,N_12620,N_11810);
nand U15894 (N_15894,N_10304,N_11607);
nor U15895 (N_15895,N_11658,N_11692);
nand U15896 (N_15896,N_12469,N_14467);
nand U15897 (N_15897,N_13764,N_11630);
nor U15898 (N_15898,N_11381,N_12052);
and U15899 (N_15899,N_11557,N_11828);
and U15900 (N_15900,N_10173,N_14045);
xnor U15901 (N_15901,N_13853,N_14626);
nor U15902 (N_15902,N_12025,N_10381);
nor U15903 (N_15903,N_11504,N_11500);
nor U15904 (N_15904,N_14358,N_14491);
xnor U15905 (N_15905,N_11363,N_11253);
nand U15906 (N_15906,N_12192,N_11239);
xor U15907 (N_15907,N_12370,N_14262);
and U15908 (N_15908,N_11842,N_12098);
and U15909 (N_15909,N_12933,N_12660);
nand U15910 (N_15910,N_13773,N_14417);
nand U15911 (N_15911,N_14438,N_10641);
and U15912 (N_15912,N_11005,N_10675);
nor U15913 (N_15913,N_11183,N_13672);
nor U15914 (N_15914,N_14128,N_14812);
nor U15915 (N_15915,N_14558,N_11964);
or U15916 (N_15916,N_14078,N_11615);
or U15917 (N_15917,N_13973,N_13810);
nor U15918 (N_15918,N_13767,N_10332);
or U15919 (N_15919,N_11170,N_13502);
nor U15920 (N_15920,N_10668,N_11402);
and U15921 (N_15921,N_14127,N_11049);
nor U15922 (N_15922,N_10282,N_11689);
and U15923 (N_15923,N_10258,N_12287);
nand U15924 (N_15924,N_14184,N_11179);
and U15925 (N_15925,N_13538,N_13572);
and U15926 (N_15926,N_11996,N_13390);
nand U15927 (N_15927,N_10474,N_12185);
and U15928 (N_15928,N_13586,N_13828);
or U15929 (N_15929,N_11649,N_14067);
nor U15930 (N_15930,N_10719,N_13329);
or U15931 (N_15931,N_10722,N_12752);
and U15932 (N_15932,N_13877,N_11144);
nor U15933 (N_15933,N_14801,N_14959);
nor U15934 (N_15934,N_10484,N_12249);
or U15935 (N_15935,N_14691,N_12853);
or U15936 (N_15936,N_10759,N_12835);
nor U15937 (N_15937,N_10623,N_10225);
and U15938 (N_15938,N_11748,N_12093);
nand U15939 (N_15939,N_12432,N_12363);
nand U15940 (N_15940,N_13255,N_12545);
nand U15941 (N_15941,N_11024,N_10511);
or U15942 (N_15942,N_14408,N_11916);
and U15943 (N_15943,N_14063,N_11681);
xor U15944 (N_15944,N_12017,N_14337);
or U15945 (N_15945,N_11488,N_11119);
nand U15946 (N_15946,N_12967,N_12621);
or U15947 (N_15947,N_14796,N_13232);
or U15948 (N_15948,N_14633,N_14711);
or U15949 (N_15949,N_12426,N_11172);
xnor U15950 (N_15950,N_12387,N_12091);
nor U15951 (N_15951,N_11513,N_10095);
and U15952 (N_15952,N_14512,N_10290);
nand U15953 (N_15953,N_10679,N_12735);
xor U15954 (N_15954,N_12798,N_14654);
nor U15955 (N_15955,N_10022,N_10456);
or U15956 (N_15956,N_11777,N_12366);
nand U15957 (N_15957,N_11528,N_12891);
or U15958 (N_15958,N_14373,N_12895);
nor U15959 (N_15959,N_13120,N_10136);
and U15960 (N_15960,N_13194,N_11186);
or U15961 (N_15961,N_11339,N_10274);
or U15962 (N_15962,N_11160,N_12332);
nor U15963 (N_15963,N_10978,N_13594);
or U15964 (N_15964,N_12449,N_12581);
or U15965 (N_15965,N_11292,N_11560);
xor U15966 (N_15966,N_13519,N_14121);
and U15967 (N_15967,N_14670,N_11323);
or U15968 (N_15968,N_14486,N_10656);
or U15969 (N_15969,N_13544,N_10620);
or U15970 (N_15970,N_11262,N_13073);
and U15971 (N_15971,N_13601,N_11463);
nor U15972 (N_15972,N_13280,N_11892);
nor U15973 (N_15973,N_11110,N_10975);
or U15974 (N_15974,N_13478,N_12008);
nor U15975 (N_15975,N_13452,N_11895);
and U15976 (N_15976,N_11563,N_13286);
xor U15977 (N_15977,N_13640,N_10188);
and U15978 (N_15978,N_14878,N_12172);
nand U15979 (N_15979,N_12331,N_10624);
and U15980 (N_15980,N_14675,N_10323);
and U15981 (N_15981,N_11320,N_12281);
xnor U15982 (N_15982,N_11547,N_11755);
nand U15983 (N_15983,N_12097,N_11532);
nand U15984 (N_15984,N_11592,N_13225);
and U15985 (N_15985,N_14810,N_14849);
or U15986 (N_15986,N_11695,N_11848);
nor U15987 (N_15987,N_12070,N_13911);
or U15988 (N_15988,N_12220,N_11646);
nor U15989 (N_15989,N_10561,N_13976);
and U15990 (N_15990,N_13230,N_14531);
nand U15991 (N_15991,N_14658,N_10881);
or U15992 (N_15992,N_10120,N_10314);
or U15993 (N_15993,N_11045,N_13909);
and U15994 (N_15994,N_14053,N_10414);
and U15995 (N_15995,N_10925,N_10066);
nor U15996 (N_15996,N_12819,N_14311);
nand U15997 (N_15997,N_14484,N_14729);
nand U15998 (N_15998,N_10036,N_11321);
or U15999 (N_15999,N_10527,N_12546);
or U16000 (N_16000,N_12910,N_14396);
nand U16001 (N_16001,N_14428,N_10183);
or U16002 (N_16002,N_14733,N_11266);
nand U16003 (N_16003,N_14210,N_10167);
or U16004 (N_16004,N_14761,N_13631);
nor U16005 (N_16005,N_14816,N_12082);
nor U16006 (N_16006,N_13667,N_10573);
xnor U16007 (N_16007,N_10394,N_10352);
nand U16008 (N_16008,N_14033,N_11548);
nand U16009 (N_16009,N_14347,N_11876);
nand U16010 (N_16010,N_10736,N_14891);
nand U16011 (N_16011,N_13679,N_10615);
or U16012 (N_16012,N_13111,N_14162);
or U16013 (N_16013,N_11388,N_10313);
or U16014 (N_16014,N_12657,N_13128);
nand U16015 (N_16015,N_14458,N_13985);
nor U16016 (N_16016,N_10647,N_14464);
or U16017 (N_16017,N_14202,N_10559);
nor U16018 (N_16018,N_12010,N_12204);
nor U16019 (N_16019,N_13004,N_13980);
and U16020 (N_16020,N_13732,N_13327);
nor U16021 (N_16021,N_14541,N_11099);
and U16022 (N_16022,N_13382,N_12914);
or U16023 (N_16023,N_11300,N_12322);
nand U16024 (N_16024,N_14600,N_14792);
xnor U16025 (N_16025,N_10061,N_12625);
nor U16026 (N_16026,N_13784,N_12611);
or U16027 (N_16027,N_14331,N_10021);
and U16028 (N_16028,N_13691,N_13486);
nor U16029 (N_16029,N_12306,N_13350);
nand U16030 (N_16030,N_13163,N_14702);
and U16031 (N_16031,N_10275,N_10920);
or U16032 (N_16032,N_13589,N_12291);
nor U16033 (N_16033,N_13346,N_13879);
nand U16034 (N_16034,N_11358,N_12903);
and U16035 (N_16035,N_14703,N_11269);
nor U16036 (N_16036,N_13639,N_13581);
xnor U16037 (N_16037,N_13060,N_10174);
and U16038 (N_16038,N_10678,N_10799);
nand U16039 (N_16039,N_14183,N_13516);
nand U16040 (N_16040,N_12534,N_12700);
and U16041 (N_16041,N_14829,N_13105);
nor U16042 (N_16042,N_12158,N_13927);
or U16043 (N_16043,N_12527,N_11452);
nor U16044 (N_16044,N_14270,N_10249);
nand U16045 (N_16045,N_13520,N_11795);
and U16046 (N_16046,N_12227,N_14154);
nand U16047 (N_16047,N_11192,N_10595);
and U16048 (N_16048,N_13306,N_14074);
nand U16049 (N_16049,N_10880,N_10303);
nand U16050 (N_16050,N_13646,N_14532);
nand U16051 (N_16051,N_14618,N_11727);
and U16052 (N_16052,N_13039,N_12108);
and U16053 (N_16053,N_12743,N_12444);
and U16054 (N_16054,N_11708,N_11114);
nand U16055 (N_16055,N_13136,N_14862);
and U16056 (N_16056,N_11794,N_13655);
or U16057 (N_16057,N_14456,N_10744);
nand U16058 (N_16058,N_10503,N_14315);
or U16059 (N_16059,N_14300,N_13527);
and U16060 (N_16060,N_14646,N_12501);
nor U16061 (N_16061,N_14037,N_13542);
or U16062 (N_16062,N_13491,N_10747);
nand U16063 (N_16063,N_10868,N_10891);
nor U16064 (N_16064,N_14359,N_13536);
and U16065 (N_16065,N_12618,N_10043);
or U16066 (N_16066,N_12245,N_14602);
and U16067 (N_16067,N_13031,N_11549);
nor U16068 (N_16068,N_12841,N_14089);
and U16069 (N_16069,N_12924,N_14554);
or U16070 (N_16070,N_13970,N_11012);
or U16071 (N_16071,N_10950,N_11703);
xnor U16072 (N_16072,N_12035,N_14266);
nand U16073 (N_16073,N_14209,N_12312);
xnor U16074 (N_16074,N_14489,N_14124);
nor U16075 (N_16075,N_10667,N_10311);
nor U16076 (N_16076,N_12064,N_11324);
and U16077 (N_16077,N_14511,N_14278);
or U16078 (N_16078,N_12542,N_14330);
and U16079 (N_16079,N_11685,N_14048);
nand U16080 (N_16080,N_13592,N_12701);
xnor U16081 (N_16081,N_14683,N_13369);
nor U16082 (N_16082,N_10235,N_12751);
and U16083 (N_16083,N_11884,N_14982);
nor U16084 (N_16084,N_14866,N_14075);
or U16085 (N_16085,N_10384,N_11906);
xor U16086 (N_16086,N_12248,N_10152);
or U16087 (N_16087,N_11518,N_12989);
and U16088 (N_16088,N_14137,N_12024);
nor U16089 (N_16089,N_13143,N_13124);
nand U16090 (N_16090,N_13156,N_10164);
nand U16091 (N_16091,N_10199,N_12617);
nor U16092 (N_16092,N_11830,N_10829);
and U16093 (N_16093,N_10032,N_13761);
nor U16094 (N_16094,N_12966,N_13265);
and U16095 (N_16095,N_11450,N_10918);
or U16096 (N_16096,N_12778,N_10760);
and U16097 (N_16097,N_10694,N_14875);
nor U16098 (N_16098,N_10471,N_13107);
and U16099 (N_16099,N_14766,N_12624);
and U16100 (N_16100,N_12571,N_14911);
or U16101 (N_16101,N_13086,N_12623);
and U16102 (N_16102,N_10809,N_14351);
nand U16103 (N_16103,N_14113,N_14355);
nand U16104 (N_16104,N_10935,N_12060);
and U16105 (N_16105,N_12973,N_10268);
xnor U16106 (N_16106,N_13846,N_14989);
or U16107 (N_16107,N_12196,N_14388);
or U16108 (N_16108,N_13034,N_10140);
nor U16109 (N_16109,N_12474,N_10879);
and U16110 (N_16110,N_10943,N_14993);
and U16111 (N_16111,N_11975,N_11435);
nor U16112 (N_16112,N_13775,N_13222);
and U16113 (N_16113,N_13080,N_14234);
nor U16114 (N_16114,N_10206,N_12558);
nand U16115 (N_16115,N_11185,N_11805);
nor U16116 (N_16116,N_11181,N_11399);
xor U16117 (N_16117,N_12126,N_10566);
or U16118 (N_16118,N_11359,N_11832);
nand U16119 (N_16119,N_13645,N_11215);
and U16120 (N_16120,N_13824,N_13411);
nand U16121 (N_16121,N_13904,N_14370);
or U16122 (N_16122,N_14569,N_10210);
nor U16123 (N_16123,N_13811,N_14799);
or U16124 (N_16124,N_14647,N_12310);
and U16125 (N_16125,N_14539,N_12828);
xor U16126 (N_16126,N_12047,N_14868);
and U16127 (N_16127,N_14975,N_13499);
nor U16128 (N_16128,N_12561,N_13723);
or U16129 (N_16129,N_10576,N_11645);
nand U16130 (N_16130,N_14945,N_14584);
nor U16131 (N_16131,N_11919,N_10778);
or U16132 (N_16132,N_11998,N_12375);
and U16133 (N_16133,N_13813,N_12652);
and U16134 (N_16134,N_14953,N_14870);
nor U16135 (N_16135,N_12400,N_11656);
and U16136 (N_16136,N_14641,N_14864);
nor U16137 (N_16137,N_12996,N_14712);
xnor U16138 (N_16138,N_10040,N_11562);
nor U16139 (N_16139,N_13148,N_10276);
nand U16140 (N_16140,N_10504,N_10081);
nand U16141 (N_16141,N_11652,N_11213);
nor U16142 (N_16142,N_11176,N_11929);
and U16143 (N_16143,N_13300,N_11654);
nand U16144 (N_16144,N_14720,N_11918);
or U16145 (N_16145,N_12644,N_13200);
and U16146 (N_16146,N_12230,N_10278);
nand U16147 (N_16147,N_14199,N_13371);
nand U16148 (N_16148,N_10372,N_13882);
or U16149 (N_16149,N_12641,N_13940);
and U16150 (N_16150,N_12628,N_12455);
nand U16151 (N_16151,N_11288,N_13713);
or U16152 (N_16152,N_12042,N_11445);
xnor U16153 (N_16153,N_14368,N_14348);
or U16154 (N_16154,N_10185,N_14111);
or U16155 (N_16155,N_14844,N_13765);
xnor U16156 (N_16156,N_13212,N_14000);
and U16157 (N_16157,N_10317,N_12646);
or U16158 (N_16158,N_10823,N_10708);
or U16159 (N_16159,N_11453,N_13506);
and U16160 (N_16160,N_14313,N_12746);
nand U16161 (N_16161,N_14831,N_10112);
nor U16162 (N_16162,N_10941,N_11237);
and U16163 (N_16163,N_13847,N_14047);
nor U16164 (N_16164,N_10261,N_12106);
and U16165 (N_16165,N_13951,N_10924);
nor U16166 (N_16166,N_11440,N_10547);
or U16167 (N_16167,N_11372,N_13236);
nor U16168 (N_16168,N_12675,N_10500);
nor U16169 (N_16169,N_12465,N_14502);
nor U16170 (N_16170,N_14240,N_10949);
nand U16171 (N_16171,N_10619,N_14755);
nor U16172 (N_16172,N_10048,N_11763);
and U16173 (N_16173,N_14411,N_13849);
nand U16174 (N_16174,N_14854,N_10086);
xor U16175 (N_16175,N_14104,N_14336);
nand U16176 (N_16176,N_13396,N_12792);
or U16177 (N_16177,N_14974,N_10237);
nand U16178 (N_16178,N_13922,N_12349);
and U16179 (N_16179,N_14099,N_14931);
or U16180 (N_16180,N_12438,N_12553);
or U16181 (N_16181,N_11799,N_11683);
and U16182 (N_16182,N_12078,N_10440);
nand U16183 (N_16183,N_11702,N_10887);
nor U16184 (N_16184,N_11687,N_10271);
xnor U16185 (N_16185,N_13198,N_11178);
nand U16186 (N_16186,N_10672,N_12273);
and U16187 (N_16187,N_12446,N_13718);
nor U16188 (N_16188,N_10195,N_10697);
nand U16189 (N_16189,N_11055,N_13359);
and U16190 (N_16190,N_13656,N_12975);
nor U16191 (N_16191,N_11151,N_13711);
nor U16192 (N_16192,N_12846,N_14521);
and U16193 (N_16193,N_10964,N_13181);
nor U16194 (N_16194,N_11584,N_14846);
xor U16195 (N_16195,N_11389,N_13270);
or U16196 (N_16196,N_14400,N_13751);
nand U16197 (N_16197,N_10610,N_14763);
nor U16198 (N_16198,N_12976,N_11439);
nand U16199 (N_16199,N_11496,N_10800);
nand U16200 (N_16200,N_11376,N_10642);
nor U16201 (N_16201,N_11067,N_11347);
nand U16202 (N_16202,N_12759,N_13565);
nor U16203 (N_16203,N_14179,N_13653);
or U16204 (N_16204,N_12001,N_13641);
and U16205 (N_16205,N_14823,N_14995);
and U16206 (N_16206,N_13114,N_12670);
xnor U16207 (N_16207,N_11226,N_13867);
or U16208 (N_16208,N_13261,N_11904);
nand U16209 (N_16209,N_10505,N_12264);
or U16210 (N_16210,N_14103,N_13684);
nand U16211 (N_16211,N_14357,N_14574);
xor U16212 (N_16212,N_13533,N_14019);
nor U16213 (N_16213,N_13484,N_10248);
or U16214 (N_16214,N_14249,N_11487);
and U16215 (N_16215,N_13777,N_11743);
and U16216 (N_16216,N_13215,N_11420);
nand U16217 (N_16217,N_12927,N_14265);
nand U16218 (N_16218,N_12085,N_14519);
or U16219 (N_16219,N_10974,N_11430);
nor U16220 (N_16220,N_11497,N_10532);
and U16221 (N_16221,N_10217,N_13968);
nor U16222 (N_16222,N_13929,N_11617);
or U16223 (N_16223,N_13315,N_11419);
xnor U16224 (N_16224,N_12683,N_11409);
nand U16225 (N_16225,N_13020,N_14842);
and U16226 (N_16226,N_12718,N_11940);
nor U16227 (N_16227,N_10453,N_12043);
or U16228 (N_16228,N_13894,N_14071);
nor U16229 (N_16229,N_14809,N_11256);
or U16230 (N_16230,N_11344,N_14004);
or U16231 (N_16231,N_13495,N_10725);
or U16232 (N_16232,N_11888,N_13153);
nand U16233 (N_16233,N_11742,N_14960);
nand U16234 (N_16234,N_13501,N_11438);
and U16235 (N_16235,N_14913,N_13636);
nor U16236 (N_16236,N_10165,N_10244);
nand U16237 (N_16237,N_14565,N_12486);
xnor U16238 (N_16238,N_14390,N_13488);
nor U16239 (N_16239,N_11161,N_13338);
and U16240 (N_16240,N_14505,N_13815);
and U16241 (N_16241,N_10938,N_10348);
xnor U16242 (N_16242,N_13883,N_14847);
or U16243 (N_16243,N_13085,N_10789);
and U16244 (N_16244,N_10996,N_10721);
nor U16245 (N_16245,N_13278,N_11022);
and U16246 (N_16246,N_13318,N_10768);
or U16247 (N_16247,N_13429,N_10024);
nand U16248 (N_16248,N_12847,N_10959);
or U16249 (N_16249,N_12372,N_11679);
and U16250 (N_16250,N_14079,N_11223);
or U16251 (N_16251,N_12065,N_11397);
nand U16252 (N_16252,N_11136,N_10544);
nor U16253 (N_16253,N_13027,N_13150);
nand U16254 (N_16254,N_11414,N_13971);
or U16255 (N_16255,N_13458,N_13938);
nor U16256 (N_16256,N_12498,N_14666);
nor U16257 (N_16257,N_13091,N_13541);
and U16258 (N_16258,N_13635,N_13574);
or U16259 (N_16259,N_12362,N_12580);
or U16260 (N_16260,N_13795,N_12343);
and U16261 (N_16261,N_11141,N_12523);
nor U16262 (N_16262,N_11915,N_14695);
or U16263 (N_16263,N_12226,N_14280);
or U16264 (N_16264,N_11482,N_13419);
xor U16265 (N_16265,N_12982,N_12005);
nor U16266 (N_16266,N_10570,N_10117);
nand U16267 (N_16267,N_14431,N_12462);
or U16268 (N_16268,N_14469,N_12609);
or U16269 (N_16269,N_13432,N_10514);
and U16270 (N_16270,N_13158,N_12822);
and U16271 (N_16271,N_11220,N_12936);
xor U16272 (N_16272,N_10592,N_14100);
nand U16273 (N_16273,N_14879,N_12067);
and U16274 (N_16274,N_13276,N_11326);
nor U16275 (N_16275,N_11287,N_12253);
xor U16276 (N_16276,N_11677,N_13469);
xnor U16277 (N_16277,N_10764,N_14105);
nor U16278 (N_16278,N_14427,N_14546);
or U16279 (N_16279,N_13493,N_11056);
or U16280 (N_16280,N_10263,N_13611);
nor U16281 (N_16281,N_12409,N_10835);
nor U16282 (N_16282,N_10849,N_12428);
or U16283 (N_16283,N_11222,N_14674);
nand U16284 (N_16284,N_12838,N_12433);
and U16285 (N_16285,N_12327,N_11242);
or U16286 (N_16286,N_11786,N_14506);
and U16287 (N_16287,N_10094,N_13101);
or U16288 (N_16288,N_14474,N_14684);
nor U16289 (N_16289,N_13125,N_13835);
or U16290 (N_16290,N_12165,N_10405);
nor U16291 (N_16291,N_10015,N_14483);
and U16292 (N_16292,N_14462,N_10510);
and U16293 (N_16293,N_12419,N_14361);
nand U16294 (N_16294,N_14470,N_13069);
and U16295 (N_16295,N_11819,N_14312);
nand U16296 (N_16296,N_12144,N_12351);
or U16297 (N_16297,N_12277,N_11955);
or U16298 (N_16298,N_14867,N_10428);
and U16299 (N_16299,N_11772,N_10101);
xor U16300 (N_16300,N_14192,N_12377);
or U16301 (N_16301,N_11849,N_12510);
nor U16302 (N_16302,N_12505,N_14222);
nand U16303 (N_16303,N_10157,N_10269);
and U16304 (N_16304,N_14363,N_14550);
or U16305 (N_16305,N_10351,N_11527);
or U16306 (N_16306,N_10900,N_11816);
nor U16307 (N_16307,N_11400,N_14068);
xor U16308 (N_16308,N_11212,N_13955);
and U16309 (N_16309,N_11857,N_12139);
nand U16310 (N_16310,N_10279,N_14354);
nand U16311 (N_16311,N_10655,N_12696);
and U16312 (N_16312,N_12061,N_13595);
xor U16313 (N_16313,N_10144,N_14837);
and U16314 (N_16314,N_14436,N_14282);
nand U16315 (N_16315,N_11616,N_10819);
or U16316 (N_16316,N_11731,N_11330);
or U16317 (N_16317,N_11006,N_14619);
nand U16318 (N_16318,N_12305,N_11806);
and U16319 (N_16319,N_11000,N_12478);
nand U16320 (N_16320,N_10522,N_13752);
or U16321 (N_16321,N_10927,N_12162);
xor U16322 (N_16322,N_12672,N_13665);
and U16323 (N_16323,N_10342,N_10436);
and U16324 (N_16324,N_11041,N_13778);
nand U16325 (N_16325,N_14961,N_12347);
xnor U16326 (N_16326,N_12443,N_13963);
nor U16327 (N_16327,N_12889,N_14010);
nor U16328 (N_16328,N_14015,N_13321);
nand U16329 (N_16329,N_10153,N_12054);
and U16330 (N_16330,N_11348,N_11539);
xor U16331 (N_16331,N_11140,N_10498);
nor U16332 (N_16332,N_11920,N_12101);
nor U16333 (N_16333,N_11437,N_14006);
nand U16334 (N_16334,N_12452,N_12405);
nand U16335 (N_16335,N_10896,N_13063);
or U16336 (N_16336,N_11651,N_12538);
xor U16337 (N_16337,N_12214,N_11128);
xnor U16338 (N_16338,N_11822,N_10395);
nand U16339 (N_16339,N_12551,N_13740);
nor U16340 (N_16340,N_10877,N_14552);
nor U16341 (N_16341,N_13185,N_13668);
nor U16342 (N_16342,N_13420,N_13776);
and U16343 (N_16343,N_10286,N_13248);
and U16344 (N_16344,N_12658,N_13174);
nor U16345 (N_16345,N_12793,N_11707);
nand U16346 (N_16346,N_13570,N_11590);
nor U16347 (N_16347,N_13914,N_10016);
and U16348 (N_16348,N_13700,N_12193);
nand U16349 (N_16349,N_12038,N_13126);
nor U16350 (N_16350,N_11143,N_14308);
and U16351 (N_16351,N_10463,N_11717);
nor U16352 (N_16352,N_10360,N_10733);
or U16353 (N_16353,N_13774,N_13546);
nand U16354 (N_16354,N_10065,N_14310);
and U16355 (N_16355,N_12512,N_12134);
nand U16356 (N_16356,N_14529,N_13235);
nor U16357 (N_16357,N_13733,N_12954);
or U16358 (N_16358,N_10998,N_14087);
and U16359 (N_16359,N_11394,N_10408);
and U16360 (N_16360,N_14166,N_14698);
nand U16361 (N_16361,N_12396,N_10424);
or U16362 (N_16362,N_10429,N_13618);
nor U16363 (N_16363,N_13906,N_14158);
or U16364 (N_16364,N_13250,N_11077);
nor U16365 (N_16365,N_10160,N_13633);
or U16366 (N_16366,N_12122,N_11273);
or U16367 (N_16367,N_12006,N_11812);
xor U16368 (N_16368,N_10318,N_14776);
xor U16369 (N_16369,N_10330,N_13539);
xnor U16370 (N_16370,N_14446,N_14453);
or U16371 (N_16371,N_12804,N_14795);
nand U16372 (N_16372,N_11604,N_14066);
or U16373 (N_16373,N_14080,N_13356);
nand U16374 (N_16374,N_13737,N_12420);
and U16375 (N_16375,N_13050,N_13258);
and U16376 (N_16376,N_14263,N_12904);
nand U16377 (N_16377,N_13159,N_11991);
nand U16378 (N_16378,N_13889,N_13731);
nor U16379 (N_16379,N_11873,N_14237);
nor U16380 (N_16380,N_13347,N_13590);
and U16381 (N_16381,N_10932,N_14410);
and U16382 (N_16382,N_11299,N_11081);
and U16383 (N_16383,N_10756,N_13935);
nand U16384 (N_16384,N_14477,N_12224);
xnor U16385 (N_16385,N_14561,N_11457);
nor U16386 (N_16386,N_11824,N_13872);
and U16387 (N_16387,N_10097,N_12194);
or U16388 (N_16388,N_13030,N_12530);
nand U16389 (N_16389,N_12413,N_12040);
or U16390 (N_16390,N_13583,N_12050);
or U16391 (N_16391,N_14383,N_11232);
nand U16392 (N_16392,N_11889,N_12648);
xnor U16393 (N_16393,N_14223,N_14218);
or U16394 (N_16394,N_10990,N_14386);
nand U16395 (N_16395,N_11097,N_10496);
or U16396 (N_16396,N_10159,N_14665);
or U16397 (N_16397,N_12261,N_12272);
nand U16398 (N_16398,N_14238,N_11203);
and U16399 (N_16399,N_13622,N_11159);
and U16400 (N_16400,N_14095,N_12592);
nor U16401 (N_16401,N_14892,N_12500);
or U16402 (N_16402,N_10034,N_11351);
nand U16403 (N_16403,N_13807,N_11974);
xor U16404 (N_16404,N_13418,N_11709);
and U16405 (N_16405,N_12406,N_11555);
xor U16406 (N_16406,N_12348,N_12845);
nor U16407 (N_16407,N_11572,N_11443);
nand U16408 (N_16408,N_12286,N_14527);
or U16409 (N_16409,N_13234,N_13064);
or U16410 (N_16410,N_11211,N_13357);
and U16411 (N_16411,N_12189,N_11665);
nor U16412 (N_16412,N_10810,N_13898);
and U16413 (N_16413,N_11739,N_11194);
nor U16414 (N_16414,N_13596,N_11475);
xor U16415 (N_16415,N_10534,N_14461);
and U16416 (N_16416,N_11657,N_12262);
nor U16417 (N_16417,N_11182,N_13724);
xnor U16418 (N_16418,N_10423,N_11636);
or U16419 (N_16419,N_14570,N_11573);
or U16420 (N_16420,N_14622,N_13961);
and U16421 (N_16421,N_14990,N_12762);
xnor U16422 (N_16422,N_14316,N_11956);
or U16423 (N_16423,N_11897,N_13127);
or U16424 (N_16424,N_14479,N_14855);
and U16425 (N_16425,N_14342,N_12456);
nand U16426 (N_16426,N_12022,N_13016);
xor U16427 (N_16427,N_14840,N_12645);
nand U16428 (N_16428,N_12477,N_14070);
and U16429 (N_16429,N_14448,N_10981);
nor U16430 (N_16430,N_10251,N_14375);
xor U16431 (N_16431,N_11781,N_13448);
nand U16432 (N_16432,N_13692,N_10264);
nand U16433 (N_16433,N_12964,N_13597);
nand U16434 (N_16434,N_11612,N_14401);
and U16435 (N_16435,N_13540,N_13035);
and U16436 (N_16436,N_14429,N_10822);
and U16437 (N_16437,N_12852,N_13576);
nor U16438 (N_16438,N_13977,N_13070);
xor U16439 (N_16439,N_13284,N_10398);
or U16440 (N_16440,N_14011,N_13662);
nor U16441 (N_16441,N_13623,N_14378);
nor U16442 (N_16442,N_14091,N_14157);
xor U16443 (N_16443,N_11661,N_14466);
and U16444 (N_16444,N_12613,N_12507);
and U16445 (N_16445,N_13106,N_12865);
xor U16446 (N_16446,N_14865,N_13557);
and U16447 (N_16447,N_14333,N_13986);
nor U16448 (N_16448,N_10007,N_11936);
nor U16449 (N_16449,N_12089,N_12741);
or U16450 (N_16450,N_14146,N_13962);
or U16451 (N_16451,N_12576,N_13220);
or U16452 (N_16452,N_10908,N_14134);
xnor U16453 (N_16453,N_11459,N_14901);
and U16454 (N_16454,N_12303,N_13336);
or U16455 (N_16455,N_10928,N_13147);
xor U16456 (N_16456,N_10107,N_13322);
xor U16457 (N_16457,N_14517,N_10614);
nand U16458 (N_16458,N_14929,N_11626);
nand U16459 (N_16459,N_14576,N_13354);
and U16460 (N_16460,N_12073,N_14049);
xor U16461 (N_16461,N_11713,N_11598);
xnor U16462 (N_16462,N_13823,N_12231);
and U16463 (N_16463,N_13825,N_10843);
and U16464 (N_16464,N_13412,N_14284);
xnor U16465 (N_16465,N_13009,N_12345);
or U16466 (N_16466,N_13373,N_10404);
xnor U16467 (N_16467,N_11647,N_11529);
nor U16468 (N_16468,N_13703,N_14668);
or U16469 (N_16469,N_13663,N_11864);
nor U16470 (N_16470,N_11886,N_13097);
nor U16471 (N_16471,N_11362,N_13559);
and U16472 (N_16472,N_11249,N_14281);
and U16473 (N_16473,N_14072,N_11597);
and U16474 (N_16474,N_12206,N_10761);
or U16475 (N_16475,N_10113,N_13996);
nor U16476 (N_16476,N_12629,N_10859);
or U16477 (N_16477,N_11050,N_12149);
or U16478 (N_16478,N_10838,N_11120);
or U16479 (N_16479,N_10734,N_11845);
and U16480 (N_16480,N_13715,N_11556);
nand U16481 (N_16481,N_12519,N_12285);
nor U16482 (N_16482,N_12610,N_10669);
nor U16483 (N_16483,N_13861,N_10867);
nand U16484 (N_16484,N_12834,N_11844);
and U16485 (N_16485,N_14819,N_11701);
and U16486 (N_16486,N_10574,N_12059);
and U16487 (N_16487,N_12948,N_13307);
or U16488 (N_16488,N_12619,N_14678);
or U16489 (N_16489,N_12485,N_13407);
nand U16490 (N_16490,N_10551,N_13078);
nor U16491 (N_16491,N_13046,N_11558);
and U16492 (N_16492,N_13960,N_10400);
or U16493 (N_16493,N_13620,N_13884);
and U16494 (N_16494,N_11704,N_12567);
or U16495 (N_16495,N_14572,N_14621);
and U16496 (N_16496,N_11498,N_13003);
nand U16497 (N_16497,N_11085,N_10119);
xnor U16498 (N_16498,N_14578,N_11710);
nand U16499 (N_16499,N_14178,N_14194);
or U16500 (N_16500,N_10915,N_13798);
xnor U16501 (N_16501,N_13992,N_12376);
and U16502 (N_16502,N_14748,N_11698);
and U16503 (N_16503,N_11838,N_12560);
and U16504 (N_16504,N_11216,N_13231);
nor U16505 (N_16505,N_10126,N_13160);
or U16506 (N_16506,N_10792,N_13287);
nand U16507 (N_16507,N_13476,N_12153);
nor U16508 (N_16508,N_10328,N_14597);
or U16509 (N_16509,N_11392,N_13413);
nand U16510 (N_16510,N_11346,N_14568);
nor U16511 (N_16511,N_11305,N_11312);
nand U16512 (N_16512,N_11984,N_12926);
xnor U16513 (N_16513,N_11011,N_10654);
or U16514 (N_16514,N_10011,N_13991);
and U16515 (N_16515,N_11982,N_12999);
xor U16516 (N_16516,N_13903,N_10685);
nand U16517 (N_16517,N_12239,N_10553);
nor U16518 (N_16518,N_10170,N_14732);
nor U16519 (N_16519,N_13805,N_12147);
and U16520 (N_16520,N_13865,N_13702);
nand U16521 (N_16521,N_12120,N_11568);
nor U16522 (N_16522,N_10280,N_11429);
nor U16523 (N_16523,N_14449,N_11009);
and U16524 (N_16524,N_14472,N_13405);
or U16525 (N_16525,N_11552,N_10909);
and U16526 (N_16526,N_14254,N_10578);
nor U16527 (N_16527,N_10427,N_10876);
and U16528 (N_16528,N_14480,N_13304);
and U16529 (N_16529,N_11448,N_12256);
or U16530 (N_16530,N_11663,N_11165);
xnor U16531 (N_16531,N_13042,N_10802);
or U16532 (N_16532,N_13294,N_12697);
nand U16533 (N_16533,N_10132,N_10273);
or U16534 (N_16534,N_12799,N_12565);
nand U16535 (N_16535,N_11508,N_12582);
xnor U16536 (N_16536,N_11506,N_14526);
or U16537 (N_16537,N_13317,N_11396);
nor U16538 (N_16538,N_12729,N_11720);
and U16539 (N_16539,N_10320,N_14586);
nand U16540 (N_16540,N_11928,N_14876);
nand U16541 (N_16541,N_12506,N_12094);
nor U16542 (N_16542,N_14174,N_10239);
nand U16543 (N_16543,N_13341,N_12069);
nor U16544 (N_16544,N_10686,N_13989);
nor U16545 (N_16545,N_13079,N_12131);
nor U16546 (N_16546,N_13426,N_13428);
and U16547 (N_16547,N_14243,N_12466);
xnor U16548 (N_16548,N_14515,N_11784);
and U16549 (N_16549,N_10611,N_13978);
nor U16550 (N_16550,N_13664,N_13032);
or U16551 (N_16551,N_14976,N_13302);
or U16552 (N_16552,N_12086,N_10776);
nand U16553 (N_16553,N_10637,N_14277);
or U16554 (N_16554,N_11379,N_13933);
nand U16555 (N_16555,N_14016,N_10940);
or U16556 (N_16556,N_12766,N_13238);
or U16557 (N_16557,N_10051,N_13947);
or U16558 (N_16558,N_10417,N_11113);
or U16559 (N_16559,N_14743,N_10753);
nor U16560 (N_16560,N_12045,N_14881);
nand U16561 (N_16561,N_11195,N_12386);
nand U16562 (N_16562,N_13838,N_11697);
nor U16563 (N_16563,N_13017,N_10073);
or U16564 (N_16564,N_13517,N_11325);
and U16565 (N_16565,N_11726,N_14687);
and U16566 (N_16566,N_10652,N_10368);
xnor U16567 (N_16567,N_10288,N_10373);
and U16568 (N_16568,N_12977,N_13445);
or U16569 (N_16569,N_10870,N_10688);
nand U16570 (N_16570,N_11023,N_14404);
nor U16571 (N_16571,N_13874,N_11541);
nand U16572 (N_16572,N_10343,N_12171);
and U16573 (N_16573,N_10715,N_12922);
and U16574 (N_16574,N_13736,N_13532);
nand U16575 (N_16575,N_14520,N_14443);
or U16576 (N_16576,N_11502,N_14139);
or U16577 (N_16577,N_10194,N_11280);
or U16578 (N_16578,N_12791,N_10133);
or U16579 (N_16579,N_13893,N_10914);
or U16580 (N_16580,N_13683,N_13313);
nand U16581 (N_16581,N_10739,N_13966);
nor U16582 (N_16582,N_13785,N_12212);
and U16583 (N_16583,N_12412,N_12649);
and U16584 (N_16584,N_14207,N_12307);
nand U16585 (N_16585,N_10729,N_11585);
nand U16586 (N_16586,N_14699,N_11478);
nand U16587 (N_16587,N_10898,N_13832);
nor U16588 (N_16588,N_14906,N_11574);
and U16589 (N_16589,N_11862,N_11567);
or U16590 (N_16590,N_11639,N_13067);
nand U16591 (N_16591,N_12274,N_10951);
xnor U16592 (N_16592,N_10299,N_13456);
or U16593 (N_16593,N_13103,N_13803);
and U16594 (N_16594,N_14221,N_14972);
xor U16595 (N_16595,N_14692,N_13417);
nand U16596 (N_16596,N_12435,N_11112);
and U16597 (N_16597,N_13196,N_12909);
or U16598 (N_16598,N_10963,N_11688);
xnor U16599 (N_16599,N_13132,N_13498);
and U16600 (N_16600,N_13013,N_10596);
and U16601 (N_16601,N_13170,N_12677);
xnor U16602 (N_16602,N_13720,N_12515);
nand U16603 (N_16603,N_11108,N_11660);
or U16604 (N_16604,N_10129,N_13444);
or U16605 (N_16605,N_12217,N_11147);
and U16606 (N_16606,N_14425,N_10141);
nand U16607 (N_16607,N_13055,N_10548);
nand U16608 (N_16608,N_10010,N_13116);
or U16609 (N_16609,N_10003,N_11357);
nor U16610 (N_16610,N_10814,N_12848);
and U16611 (N_16611,N_13449,N_11047);
nand U16612 (N_16612,N_10540,N_14523);
xnor U16613 (N_16613,N_12410,N_11944);
and U16614 (N_16614,N_11980,N_14645);
xnor U16615 (N_16615,N_14385,N_11322);
or U16616 (N_16616,N_12437,N_13885);
or U16617 (N_16617,N_13763,N_10002);
and U16618 (N_16618,N_13025,N_10267);
nor U16619 (N_16619,N_10301,N_13757);
nor U16620 (N_16620,N_10180,N_13730);
nor U16621 (N_16621,N_11927,N_14287);
or U16622 (N_16622,N_14496,N_12234);
nand U16623 (N_16623,N_13096,N_11576);
xnor U16624 (N_16624,N_13454,N_10702);
or U16625 (N_16625,N_13801,N_10873);
and U16626 (N_16626,N_13926,N_10860);
and U16627 (N_16627,N_13610,N_11796);
nor U16628 (N_16628,N_11177,N_14041);
or U16629 (N_16629,N_14430,N_10490);
nand U16630 (N_16630,N_14930,N_10302);
nand U16631 (N_16631,N_10422,N_10187);
and U16632 (N_16632,N_11768,N_14399);
or U16633 (N_16633,N_12280,N_13705);
nor U16634 (N_16634,N_12460,N_13340);
or U16635 (N_16635,N_13483,N_14293);
or U16636 (N_16636,N_14547,N_10608);
nand U16637 (N_16637,N_10154,N_13477);
xor U16638 (N_16638,N_13722,N_10106);
nand U16639 (N_16639,N_13529,N_10738);
and U16640 (N_16640,N_13666,N_11758);
nand U16641 (N_16641,N_14912,N_12650);
or U16642 (N_16642,N_10115,N_13438);
and U16643 (N_16643,N_14031,N_14356);
nand U16644 (N_16644,N_10393,N_14873);
nor U16645 (N_16645,N_13090,N_11174);
and U16646 (N_16646,N_11952,N_13547);
and U16647 (N_16647,N_14050,N_13771);
nor U16648 (N_16648,N_12807,N_11759);
nand U16649 (N_16649,N_10326,N_14432);
and U16650 (N_16650,N_10172,N_14167);
nor U16651 (N_16651,N_13964,N_12013);
nor U16652 (N_16652,N_11495,N_11965);
xnor U16653 (N_16653,N_13604,N_11087);
or U16654 (N_16654,N_11514,N_13259);
or U16655 (N_16655,N_12046,N_13799);
and U16656 (N_16656,N_10991,N_12699);
nor U16657 (N_16657,N_10337,N_14083);
or U16658 (N_16658,N_11706,N_12671);
or U16659 (N_16659,N_11494,N_12814);
nor U16660 (N_16660,N_10934,N_13528);
nor U16661 (N_16661,N_14451,N_13296);
and U16662 (N_16662,N_10468,N_12564);
nand U16663 (N_16663,N_14902,N_12051);
nand U16664 (N_16664,N_14244,N_10231);
and U16665 (N_16665,N_13395,N_14064);
nor U16666 (N_16666,N_12278,N_11368);
and U16667 (N_16667,N_13075,N_14850);
or U16668 (N_16668,N_13065,N_14038);
nor U16669 (N_16669,N_10872,N_13725);
xor U16670 (N_16670,N_12199,N_13796);
or U16671 (N_16671,N_10977,N_10980);
or U16672 (N_16672,N_12314,N_12260);
nor U16673 (N_16673,N_11813,N_13233);
nor U16674 (N_16674,N_14718,N_12247);
or U16675 (N_16675,N_11682,N_12574);
nand U16676 (N_16676,N_10617,N_12041);
or U16677 (N_16677,N_14407,N_11342);
and U16678 (N_16678,N_10197,N_14714);
nor U16679 (N_16679,N_13435,N_13786);
and U16680 (N_16680,N_13351,N_12125);
nor U16681 (N_16681,N_14164,N_10001);
nor U16682 (N_16682,N_13393,N_14923);
and U16683 (N_16683,N_11899,N_12297);
nand U16684 (N_16684,N_14118,N_14852);
or U16685 (N_16685,N_10229,N_13578);
nor U16686 (N_16686,N_12000,N_14857);
or U16687 (N_16687,N_12402,N_14239);
nor U16688 (N_16688,N_12757,N_14944);
or U16689 (N_16689,N_14830,N_10092);
nand U16690 (N_16690,N_12124,N_13600);
and U16691 (N_16691,N_13923,N_12167);
nand U16692 (N_16692,N_14843,N_12747);
nor U16693 (N_16693,N_14557,N_12643);
nor U16694 (N_16694,N_13459,N_11282);
xnor U16695 (N_16695,N_10491,N_12293);
nand U16696 (N_16696,N_14800,N_13716);
or U16697 (N_16697,N_11737,N_13323);
or U16698 (N_16698,N_10676,N_10519);
or U16699 (N_16699,N_11043,N_13355);
nor U16700 (N_16700,N_10236,N_14082);
nand U16701 (N_16701,N_10289,N_14279);
nor U16702 (N_16702,N_13326,N_14937);
xnor U16703 (N_16703,N_10850,N_14730);
nand U16704 (N_16704,N_10134,N_14309);
nand U16705 (N_16705,N_13954,N_14306);
nand U16706 (N_16706,N_13892,N_14180);
nand U16707 (N_16707,N_12635,N_12588);
or U16708 (N_16708,N_10700,N_14290);
nand U16709 (N_16709,N_11101,N_13617);
nor U16710 (N_16710,N_11059,N_10202);
or U16711 (N_16711,N_10782,N_14909);
and U16712 (N_16712,N_14295,N_10070);
or U16713 (N_16713,N_14009,N_11736);
or U16714 (N_16714,N_14259,N_13697);
nand U16715 (N_16715,N_14943,N_10307);
nor U16716 (N_16716,N_14256,N_12980);
nor U16717 (N_16717,N_11767,N_10658);
or U16718 (N_16718,N_11659,N_10834);
xor U16719 (N_16719,N_14379,N_10059);
and U16720 (N_16720,N_13257,N_14226);
and U16721 (N_16721,N_11863,N_11586);
nand U16722 (N_16722,N_10006,N_14522);
and U16723 (N_16723,N_11872,N_14093);
nand U16724 (N_16724,N_14549,N_14841);
or U16725 (N_16725,N_12034,N_11393);
nand U16726 (N_16726,N_12965,N_12631);
nand U16727 (N_16727,N_14736,N_13176);
and U16728 (N_16728,N_13535,N_11408);
xnor U16729 (N_16729,N_13192,N_12399);
xor U16730 (N_16730,N_12540,N_11444);
and U16731 (N_16731,N_12251,N_14595);
nand U16732 (N_16732,N_10971,N_11353);
nor U16733 (N_16733,N_10441,N_10362);
nor U16734 (N_16734,N_14575,N_10485);
or U16735 (N_16735,N_10683,N_11875);
nor U16736 (N_16736,N_12140,N_11820);
or U16737 (N_16737,N_12436,N_10651);
xnor U16738 (N_16738,N_12092,N_12781);
or U16739 (N_16739,N_13071,N_12011);
nor U16740 (N_16740,N_14559,N_10116);
nand U16741 (N_16741,N_11033,N_12992);
nand U16742 (N_16742,N_10772,N_10247);
nor U16743 (N_16743,N_13616,N_13967);
or U16744 (N_16744,N_12246,N_13146);
nand U16745 (N_16745,N_14715,N_11850);
or U16746 (N_16746,N_14828,N_10200);
xnor U16747 (N_16747,N_12941,N_12244);
xor U16748 (N_16748,N_13362,N_12457);
nand U16749 (N_16749,N_10038,N_14905);
nor U16750 (N_16750,N_14746,N_11990);
or U16751 (N_16751,N_11791,N_12554);
nand U16752 (N_16752,N_11421,N_11039);
nand U16753 (N_16753,N_10122,N_11476);
and U16754 (N_16754,N_11071,N_13804);
xor U16755 (N_16755,N_10817,N_13750);
nor U16756 (N_16756,N_11398,N_12930);
or U16757 (N_16757,N_12638,N_10028);
or U16758 (N_16758,N_12324,N_14023);
nor U16759 (N_16759,N_14538,N_13202);
or U16760 (N_16760,N_10383,N_11263);
or U16761 (N_16761,N_13826,N_10864);
nand U16762 (N_16762,N_12174,N_14439);
and U16763 (N_16763,N_10118,N_11061);
nand U16764 (N_16764,N_12491,N_10937);
or U16765 (N_16765,N_10837,N_10190);
xnor U16766 (N_16766,N_13155,N_14751);
and U16767 (N_16767,N_10584,N_10379);
and U16768 (N_16768,N_11910,N_12508);
nand U16769 (N_16769,N_12705,N_12207);
nand U16770 (N_16770,N_12728,N_14560);
nor U16771 (N_16771,N_10538,N_13451);
and U16772 (N_16772,N_12019,N_14582);
and U16773 (N_16773,N_12012,N_12938);
and U16774 (N_16774,N_13566,N_12451);
nor U16775 (N_16775,N_14144,N_13569);
and U16776 (N_16776,N_14201,N_14706);
nand U16777 (N_16777,N_14738,N_10629);
nor U16778 (N_16778,N_14450,N_13305);
or U16779 (N_16779,N_12238,N_14933);
nor U16780 (N_16780,N_11428,N_12731);
and U16781 (N_16781,N_13199,N_10613);
nand U16782 (N_16782,N_11948,N_12827);
or U16783 (N_16783,N_12937,N_11581);
xnor U16784 (N_16784,N_10009,N_13987);
nand U16785 (N_16785,N_10409,N_14999);
nand U16786 (N_16786,N_10445,N_11462);
xnor U16787 (N_16787,N_12425,N_14750);
nor U16788 (N_16788,N_11198,N_13087);
and U16789 (N_16789,N_12837,N_10186);
xnor U16790 (N_16790,N_11385,N_14460);
and U16791 (N_16791,N_11674,N_12448);
nor U16792 (N_16792,N_10594,N_12076);
nor U16793 (N_16793,N_14690,N_10528);
nor U16794 (N_16794,N_14922,N_10345);
nand U16795 (N_16795,N_13057,N_10158);
and U16796 (N_16796,N_11441,N_10459);
and U16797 (N_16797,N_13415,N_12044);
nor U16798 (N_16798,N_14272,N_14904);
or U16799 (N_16799,N_13374,N_11738);
and U16800 (N_16800,N_14770,N_11969);
nor U16801 (N_16801,N_13744,N_12023);
nor U16802 (N_16802,N_13548,N_12647);
nor U16803 (N_16803,N_12090,N_10973);
and U16804 (N_16804,N_13226,N_10890);
or U16805 (N_16805,N_11993,N_12215);
xor U16806 (N_16806,N_12328,N_13754);
nor U16807 (N_16807,N_11846,N_14002);
or U16808 (N_16808,N_12665,N_13965);
nor U16809 (N_16809,N_14932,N_12473);
xor U16810 (N_16810,N_11602,N_14117);
or U16811 (N_16811,N_13958,N_12843);
and U16812 (N_16812,N_14345,N_10058);
nor U16813 (N_16813,N_12335,N_14181);
and U16814 (N_16814,N_13738,N_11725);
nor U16815 (N_16815,N_11328,N_14581);
nor U16816 (N_16816,N_11089,N_12952);
and U16817 (N_16817,N_14253,N_14138);
and U16818 (N_16818,N_14821,N_11295);
and U16819 (N_16819,N_10416,N_14413);
nor U16820 (N_16820,N_10325,N_10921);
or U16821 (N_16821,N_14634,N_10196);
or U16822 (N_16822,N_11416,N_11470);
and U16823 (N_16823,N_13134,N_11912);
nand U16824 (N_16824,N_11874,N_12549);
or U16825 (N_16825,N_13937,N_12587);
xnor U16826 (N_16826,N_12068,N_14151);
and U16827 (N_16827,N_11611,N_14228);
nand U16828 (N_16828,N_10469,N_10960);
and U16829 (N_16829,N_11298,N_10281);
and U16830 (N_16830,N_13567,N_11751);
nor U16831 (N_16831,N_10507,N_12309);
or U16832 (N_16832,N_10597,N_14409);
and U16833 (N_16833,N_12325,N_12573);
or U16834 (N_16834,N_12622,N_14341);
nor U16835 (N_16835,N_11133,N_12667);
xnor U16836 (N_16836,N_14165,N_13860);
nor U16837 (N_16837,N_10885,N_14149);
or U16838 (N_16838,N_12353,N_12302);
or U16839 (N_16839,N_14017,N_12673);
nand U16840 (N_16840,N_11073,N_14106);
nor U16841 (N_16841,N_10462,N_13203);
nand U16842 (N_16842,N_11020,N_11284);
or U16843 (N_16843,N_12157,N_13191);
or U16844 (N_16844,N_10331,N_11446);
nor U16845 (N_16845,N_13671,N_14419);
nand U16846 (N_16846,N_11124,N_11881);
or U16847 (N_16847,N_11793,N_11355);
and U16848 (N_16848,N_10781,N_11570);
or U16849 (N_16849,N_10989,N_11569);
or U16850 (N_16850,N_13208,N_11260);
or U16851 (N_16851,N_14028,N_12356);
and U16852 (N_16852,N_10712,N_11829);
or U16853 (N_16853,N_11285,N_11341);
or U16854 (N_16854,N_11577,N_11808);
nor U16855 (N_16855,N_13227,N_14608);
or U16856 (N_16856,N_12866,N_13748);
xnor U16857 (N_16857,N_12753,N_11600);
nand U16858 (N_16858,N_13094,N_11858);
nand U16859 (N_16859,N_11542,N_10270);
nand U16860 (N_16860,N_12334,N_11921);
or U16861 (N_16861,N_10997,N_12408);
nand U16862 (N_16862,N_13364,N_10451);
and U16863 (N_16863,N_10740,N_11116);
or U16864 (N_16864,N_10703,N_10114);
and U16865 (N_16865,N_12935,N_10563);
or U16866 (N_16866,N_10020,N_12080);
or U16867 (N_16867,N_13404,N_13598);
or U16868 (N_16868,N_14899,N_14020);
or U16869 (N_16869,N_11967,N_14631);
nor U16870 (N_16870,N_10142,N_12317);
nand U16871 (N_16871,N_12056,N_11086);
and U16872 (N_16872,N_14871,N_10803);
nand U16873 (N_16873,N_11080,N_13972);
nand U16874 (N_16874,N_12703,N_11230);
or U16875 (N_16875,N_10464,N_10604);
and U16876 (N_16876,N_12202,N_14471);
and U16877 (N_16877,N_14591,N_13376);
nor U16878 (N_16878,N_11331,N_14497);
xor U16879 (N_16879,N_14914,N_13481);
and U16880 (N_16880,N_12020,N_13669);
nor U16881 (N_16881,N_14533,N_10305);
or U16882 (N_16882,N_14724,N_13023);
and U16883 (N_16883,N_13140,N_10310);
nand U16884 (N_16884,N_14163,N_13081);
xor U16885 (N_16885,N_11785,N_10111);
nand U16886 (N_16886,N_13913,N_13908);
or U16887 (N_16887,N_12321,N_13856);
nor U16888 (N_16888,N_10727,N_12704);
nand U16889 (N_16889,N_13001,N_10749);
xor U16890 (N_16890,N_14704,N_12129);
nor U16891 (N_16891,N_12698,N_12344);
or U16892 (N_16892,N_10083,N_13952);
or U16893 (N_16893,N_14564,N_14094);
nor U16894 (N_16894,N_13582,N_12279);
nor U16895 (N_16895,N_10137,N_11106);
nor U16896 (N_16896,N_13414,N_10603);
nand U16897 (N_16897,N_12774,N_13699);
and U16898 (N_16898,N_12951,N_12257);
nor U16899 (N_16899,N_10329,N_10361);
nor U16900 (N_16900,N_14543,N_12562);
or U16901 (N_16901,N_13381,N_14384);
and U16902 (N_16902,N_10664,N_12062);
nand U16903 (N_16903,N_10886,N_13195);
and U16904 (N_16904,N_13431,N_11638);
nor U16905 (N_16905,N_14034,N_12674);
or U16906 (N_16906,N_11618,N_14044);
nand U16907 (N_16907,N_11855,N_11308);
nor U16908 (N_16908,N_14669,N_11870);
or U16909 (N_16909,N_11343,N_11836);
or U16910 (N_16910,N_10805,N_11117);
xor U16911 (N_16911,N_13288,N_14304);
nor U16912 (N_16912,N_11773,N_14516);
xor U16913 (N_16913,N_13530,N_11072);
and U16914 (N_16914,N_14468,N_14596);
nand U16915 (N_16915,N_13383,N_13164);
nor U16916 (N_16916,N_14791,N_13427);
and U16917 (N_16917,N_12148,N_10801);
nor U16918 (N_16918,N_13870,N_11484);
or U16919 (N_16919,N_10618,N_10391);
nor U16920 (N_16920,N_10294,N_12984);
xor U16921 (N_16921,N_10478,N_12962);
xor U16922 (N_16922,N_12712,N_10586);
and U16923 (N_16923,N_10818,N_10588);
and U16924 (N_16924,N_13599,N_14588);
or U16925 (N_16925,N_11390,N_12888);
nand U16926 (N_16926,N_10246,N_13068);
and U16927 (N_16927,N_13245,N_12033);
or U16928 (N_16928,N_12083,N_10628);
nor U16929 (N_16929,N_10201,N_11259);
nand U16930 (N_16930,N_12200,N_13077);
nor U16931 (N_16931,N_13808,N_11942);
and U16932 (N_16932,N_10027,N_10970);
and U16933 (N_16933,N_10701,N_13634);
nor U16934 (N_16934,N_12104,N_10716);
nor U16935 (N_16935,N_13505,N_11224);
nand U16936 (N_16936,N_11559,N_11461);
xnor U16937 (N_16937,N_12710,N_14752);
and U16938 (N_16938,N_10575,N_10692);
nand U16939 (N_16939,N_12726,N_14609);
or U16940 (N_16940,N_11277,N_13216);
or U16941 (N_16941,N_12480,N_14592);
and U16942 (N_16942,N_12616,N_14142);
nand U16943 (N_16943,N_11566,N_11337);
or U16944 (N_16944,N_12884,N_14775);
or U16945 (N_16945,N_14820,N_11787);
and U16946 (N_16946,N_14455,N_13161);
nor U16947 (N_16947,N_10250,N_10524);
nor U16948 (N_16948,N_14204,N_11564);
or U16949 (N_16949,N_10952,N_12680);
and U16950 (N_16950,N_11283,N_10175);
or U16951 (N_16951,N_14835,N_13466);
or U16952 (N_16952,N_12817,N_13959);
nand U16953 (N_16953,N_13568,N_10176);
nor U16954 (N_16954,N_14949,N_13755);
nand U16955 (N_16955,N_13588,N_14252);
nand U16956 (N_16956,N_10255,N_12318);
and U16957 (N_16957,N_12468,N_11338);
or U16958 (N_16958,N_10449,N_11040);
and U16959 (N_16959,N_10905,N_10560);
or U16960 (N_16960,N_14749,N_10447);
nor U16961 (N_16961,N_12053,N_14395);
and U16962 (N_16962,N_13088,N_14007);
or U16963 (N_16963,N_11207,N_12769);
or U16964 (N_16964,N_12467,N_12776);
and U16965 (N_16965,N_11620,N_13205);
or U16966 (N_16966,N_11723,N_11757);
nand U16967 (N_16967,N_10046,N_12601);
nor U16968 (N_16968,N_14365,N_13324);
or U16969 (N_16969,N_14116,N_12276);
xnor U16970 (N_16970,N_12160,N_13681);
nor U16971 (N_16971,N_12917,N_12603);
nand U16972 (N_16972,N_13890,N_12968);
or U16973 (N_16973,N_12969,N_13561);
or U16974 (N_16974,N_14798,N_12912);
nand U16975 (N_16975,N_11015,N_13998);
nor U16976 (N_16976,N_13979,N_13489);
or U16977 (N_16977,N_11992,N_12450);
nor U16978 (N_16978,N_14740,N_10639);
or U16979 (N_16979,N_14269,N_10004);
nand U16980 (N_16980,N_14827,N_14884);
or U16981 (N_16981,N_13688,N_11684);
nand U16982 (N_16982,N_10984,N_10492);
nor U16983 (N_16983,N_10630,N_10232);
xor U16984 (N_16984,N_12651,N_12740);
nand U16985 (N_16985,N_12873,N_12855);
and U16986 (N_16986,N_11250,N_11315);
nor U16987 (N_16987,N_11349,N_13010);
nand U16988 (N_16988,N_12290,N_11606);
and U16989 (N_16989,N_11254,N_10606);
and U16990 (N_16990,N_13626,N_11302);
and U16991 (N_16991,N_11561,N_14084);
nor U16992 (N_16992,N_10168,N_14054);
or U16993 (N_16993,N_12541,N_12894);
nand U16994 (N_16994,N_12268,N_14257);
and U16995 (N_16995,N_11168,N_11030);
and U16996 (N_16996,N_12605,N_14644);
nor U16997 (N_16997,N_10512,N_13747);
and U16998 (N_16998,N_10392,N_12453);
nand U16999 (N_16999,N_12039,N_13524);
and U17000 (N_17000,N_12267,N_14605);
or U17001 (N_17001,N_14745,N_13537);
or U17002 (N_17002,N_11671,N_14663);
nor U17003 (N_17003,N_14046,N_11917);
and U17004 (N_17004,N_13916,N_14664);
xor U17005 (N_17005,N_10673,N_10841);
and U17006 (N_17006,N_13239,N_13652);
or U17007 (N_17007,N_10742,N_12738);
and U17008 (N_17008,N_11234,N_10650);
and U17009 (N_17009,N_14594,N_14340);
or U17010 (N_17010,N_14838,N_13917);
xor U17011 (N_17011,N_11048,N_10995);
nand U17012 (N_17012,N_13726,N_12596);
and U17013 (N_17013,N_10171,N_12003);
and U17014 (N_17014,N_11248,N_12209);
nand U17015 (N_17015,N_12361,N_12154);
nand U17016 (N_17016,N_10227,N_11554);
and U17017 (N_17017,N_10103,N_13545);
nor U17018 (N_17018,N_11340,N_13809);
nor U17019 (N_17019,N_12263,N_10539);
or U17020 (N_17020,N_12168,N_11240);
nor U17021 (N_17021,N_13891,N_11210);
nor U17022 (N_17022,N_12121,N_12547);
nand U17023 (N_17023,N_10795,N_10983);
and U17024 (N_17024,N_12986,N_14200);
or U17025 (N_17025,N_12031,N_11418);
nor U17026 (N_17026,N_13083,N_12714);
nand U17027 (N_17027,N_12591,N_11534);
or U17028 (N_17028,N_11551,N_13465);
nand U17029 (N_17029,N_11818,N_13794);
nand U17030 (N_17030,N_10790,N_10321);
and U17031 (N_17031,N_11676,N_10088);
nor U17032 (N_17032,N_12569,N_12758);
nor U17033 (N_17033,N_12998,N_12706);
and U17034 (N_17034,N_14734,N_14169);
nor U17035 (N_17035,N_14709,N_10875);
nor U17036 (N_17036,N_14452,N_10013);
nor U17037 (N_17037,N_12009,N_10903);
and U17038 (N_17038,N_13188,N_12690);
or U17039 (N_17039,N_14305,N_14493);
nor U17040 (N_17040,N_13941,N_14172);
nand U17041 (N_17041,N_11613,N_11265);
nor U17042 (N_17042,N_13193,N_14056);
and U17043 (N_17043,N_10178,N_10521);
nand U17044 (N_17044,N_10968,N_12993);
nand U17045 (N_17045,N_13839,N_14397);
or U17046 (N_17046,N_14635,N_14676);
nand U17047 (N_17047,N_11950,N_11778);
nor U17048 (N_17048,N_11764,N_11481);
xnor U17049 (N_17049,N_14231,N_14661);
nor U17050 (N_17050,N_11474,N_13492);
nand U17051 (N_17051,N_14510,N_12138);
nor U17052 (N_17052,N_12346,N_14725);
and U17053 (N_17053,N_10093,N_13482);
xnor U17054 (N_17054,N_14727,N_14141);
nor U17055 (N_17055,N_13686,N_12407);
or U17056 (N_17056,N_12075,N_12815);
nand U17057 (N_17057,N_14096,N_11587);
nor U17058 (N_17058,N_10074,N_11291);
and U17059 (N_17059,N_14553,N_13045);
nand U17060 (N_17060,N_11310,N_10766);
nand U17061 (N_17061,N_11753,N_13316);
nor U17062 (N_17062,N_13550,N_13670);
nor U17063 (N_17063,N_12607,N_11815);
nand U17064 (N_17064,N_12836,N_11135);
nor U17065 (N_17065,N_13184,N_10334);
and U17066 (N_17066,N_10110,N_11994);
and U17067 (N_17067,N_13480,N_12509);
nand U17068 (N_17068,N_14190,N_14934);
nor U17069 (N_17069,N_10832,N_11066);
nor U17070 (N_17070,N_13766,N_10481);
and U17071 (N_17071,N_12240,N_13279);
nand U17072 (N_17072,N_11314,N_10966);
nand U17073 (N_17073,N_14786,N_11111);
nand U17074 (N_17074,N_12734,N_10265);
nand U17075 (N_17075,N_12597,N_14299);
and U17076 (N_17076,N_11847,N_13059);
or U17077 (N_17077,N_13447,N_12301);
nor U17078 (N_17078,N_12994,N_13119);
nand U17079 (N_17079,N_14283,N_14186);
nor U17080 (N_17080,N_11512,N_10904);
or U17081 (N_17081,N_10205,N_14958);
nand U17082 (N_17082,N_13821,N_14694);
or U17083 (N_17083,N_14334,N_10515);
xor U17084 (N_17084,N_10767,N_12454);
and U17085 (N_17085,N_14030,N_12656);
nand U17086 (N_17086,N_10219,N_14216);
nor U17087 (N_17087,N_12604,N_11911);
or U17088 (N_17088,N_12074,N_10256);
or U17089 (N_17089,N_10854,N_12844);
or U17090 (N_17090,N_11971,N_11896);
and U17091 (N_17091,N_11545,N_12669);
and U17092 (N_17092,N_12856,N_13421);
and U17093 (N_17093,N_13129,N_12789);
nor U17094 (N_17094,N_14135,N_13827);
and U17095 (N_17095,N_12720,N_12502);
or U17096 (N_17096,N_13562,N_14476);
nor U17097 (N_17097,N_10826,N_13791);
and U17098 (N_17098,N_11025,N_10054);
and U17099 (N_17099,N_10087,N_12790);
or U17100 (N_17100,N_13678,N_12389);
nor U17101 (N_17101,N_14616,N_11354);
nor U17102 (N_17102,N_12959,N_11509);
nand U17103 (N_17103,N_12640,N_12779);
xor U17104 (N_17104,N_11065,N_12114);
nand U17105 (N_17105,N_12066,N_11520);
nor U17106 (N_17106,N_10714,N_11270);
or U17107 (N_17107,N_12897,N_13337);
or U17108 (N_17108,N_12463,N_13241);
or U17109 (N_17109,N_12380,N_11909);
nand U17110 (N_17110,N_11629,N_10717);
nand U17111 (N_17111,N_10390,N_10475);
nand U17112 (N_17112,N_12036,N_12557);
nand U17113 (N_17113,N_10804,N_10779);
nand U17114 (N_17114,N_12813,N_14426);
nor U17115 (N_17115,N_12183,N_10419);
nor U17116 (N_17116,N_10640,N_13403);
nand U17117 (N_17117,N_11454,N_13880);
nand U17118 (N_17118,N_12600,N_12383);
nand U17119 (N_17119,N_11173,N_12191);
nor U17120 (N_17120,N_12161,N_13348);
or U17121 (N_17121,N_14794,N_12341);
or U17122 (N_17122,N_10979,N_13430);
nand U17123 (N_17123,N_14415,N_11425);
or U17124 (N_17124,N_10124,N_11901);
nor U17125 (N_17125,N_13552,N_10765);
nand U17126 (N_17126,N_13953,N_13577);
nor U17127 (N_17127,N_11809,N_12156);
and U17128 (N_17128,N_11275,N_10988);
nand U17129 (N_17129,N_10315,N_13510);
or U17130 (N_17130,N_13379,N_11016);
and U17131 (N_17131,N_14369,N_14140);
nand U17132 (N_17132,N_11672,N_12037);
and U17133 (N_17133,N_13942,N_13871);
or U17134 (N_17134,N_10806,N_13661);
nand U17135 (N_17135,N_13384,N_10636);
and U17136 (N_17136,N_10884,N_12754);
or U17137 (N_17137,N_14032,N_13277);
xnor U17138 (N_17138,N_14481,N_14475);
nor U17139 (N_17139,N_11391,N_14863);
and U17140 (N_17140,N_14445,N_12299);
nor U17141 (N_17141,N_14133,N_14818);
nor U17142 (N_17142,N_12614,N_12717);
or U17143 (N_17143,N_10718,N_12839);
nand U17144 (N_17144,N_10653,N_12770);
nand U17145 (N_17145,N_13993,N_10784);
nand U17146 (N_17146,N_11553,N_14403);
and U17147 (N_17147,N_11383,N_12961);
and U17148 (N_17148,N_10846,N_10956);
nor U17149 (N_17149,N_13441,N_10487);
and U17150 (N_17150,N_12861,N_11680);
nand U17151 (N_17151,N_11624,N_11664);
nand U17152 (N_17152,N_14131,N_10863);
and U17153 (N_17153,N_14813,N_13817);
nand U17154 (N_17154,N_12391,N_10812);
xnor U17155 (N_17155,N_13606,N_12854);
nand U17156 (N_17156,N_11417,N_14535);
and U17157 (N_17157,N_12584,N_10411);
or U17158 (N_17158,N_14966,N_14883);
nor U17159 (N_17159,N_13455,N_12548);
or U17160 (N_17160,N_14753,N_13130);
xor U17161 (N_17161,N_10102,N_14513);
or U17162 (N_17162,N_11403,N_11601);
and U17163 (N_17163,N_11867,N_11882);
or U17164 (N_17164,N_13092,N_12990);
xor U17165 (N_17165,N_14441,N_12742);
and U17166 (N_17166,N_11696,N_14544);
nor U17167 (N_17167,N_12095,N_10691);
and U17168 (N_17168,N_11477,N_11526);
and U17169 (N_17169,N_13446,N_10389);
and U17170 (N_17170,N_14897,N_12018);
xor U17171 (N_17171,N_11001,N_12063);
or U17172 (N_17172,N_11923,N_12088);
nand U17173 (N_17173,N_13325,N_13509);
or U17174 (N_17174,N_10005,N_14636);
nand U17175 (N_17175,N_14152,N_13457);
or U17176 (N_17176,N_11247,N_11231);
nand U17177 (N_17177,N_13931,N_10050);
xor U17178 (N_17178,N_14848,N_10488);
or U17179 (N_17179,N_12367,N_12489);
nor U17180 (N_17180,N_13490,N_12497);
nand U17181 (N_17181,N_11148,N_10309);
nand U17182 (N_17182,N_11718,N_11852);
nor U17183 (N_17183,N_12719,N_12395);
and U17184 (N_17184,N_11686,N_12577);
nand U17185 (N_17185,N_14859,N_13363);
and U17186 (N_17186,N_10987,N_11770);
and U17187 (N_17187,N_12319,N_11880);
nand U17188 (N_17188,N_10203,N_11804);
nand U17189 (N_17189,N_12141,N_10435);
and U17190 (N_17190,N_14939,N_14414);
or U17191 (N_17191,N_11188,N_14992);
nor U17192 (N_17192,N_13878,N_10732);
and U17193 (N_17193,N_10008,N_14726);
nor U17194 (N_17194,N_14593,N_11995);
nand U17195 (N_17195,N_10972,N_11524);
nor U17196 (N_17196,N_10240,N_13423);
nor U17197 (N_17197,N_12928,N_11150);
nand U17198 (N_17198,N_14224,N_10690);
or U17199 (N_17199,N_10649,N_10444);
or U17200 (N_17200,N_14927,N_11122);
and U17201 (N_17201,N_13243,N_13178);
nor U17202 (N_17202,N_11835,N_12851);
or U17203 (N_17203,N_14274,N_14508);
and U17204 (N_17204,N_10533,N_12417);
xnor U17205 (N_17205,N_11914,N_10385);
xnor U17206 (N_17206,N_12142,N_11605);
nor U17207 (N_17207,N_14344,N_11167);
and U17208 (N_17208,N_14405,N_14182);
nor U17209 (N_17209,N_12653,N_13975);
nor U17210 (N_17210,N_14360,N_13851);
and U17211 (N_17211,N_10797,N_12570);
nand U17212 (N_17212,N_14924,N_13866);
or U17213 (N_17213,N_10382,N_13857);
or U17214 (N_17214,N_12877,N_11719);
and U17215 (N_17215,N_10525,N_10816);
and U17216 (N_17216,N_14882,N_11076);
xor U17217 (N_17217,N_10910,N_11522);
nand U17218 (N_17218,N_12421,N_13319);
and U17219 (N_17219,N_11744,N_14022);
nor U17220 (N_17220,N_13133,N_13436);
nand U17221 (N_17221,N_11369,N_13142);
and U17222 (N_17222,N_11014,N_10499);
nor U17223 (N_17223,N_12695,N_14444);
nor U17224 (N_17224,N_10861,N_10982);
nor U17225 (N_17225,N_14963,N_11837);
nor U17226 (N_17226,N_11989,N_12110);
and U17227 (N_17227,N_10211,N_12662);
nand U17228 (N_17228,N_12682,N_11479);
xor U17229 (N_17229,N_14996,N_12893);
nor U17230 (N_17230,N_10386,N_12228);
nand U17231 (N_17231,N_13945,N_10473);
and U17232 (N_17232,N_13207,N_14421);
nand U17233 (N_17233,N_10181,N_11480);
or U17234 (N_17234,N_14988,N_10012);
or U17235 (N_17235,N_11543,N_12458);
nand U17236 (N_17236,N_11588,N_14060);
or U17237 (N_17237,N_14632,N_14562);
or U17238 (N_17238,N_14611,N_12709);
or U17239 (N_17239,N_14406,N_10156);
and U17240 (N_17240,N_12708,N_14880);
or U17241 (N_17241,N_14973,N_13281);
nor U17242 (N_17242,N_12655,N_11932);
and U17243 (N_17243,N_10836,N_14918);
or U17244 (N_17244,N_10696,N_14217);
nand U17245 (N_17245,N_10857,N_13463);
and U17246 (N_17246,N_11642,N_14710);
and U17247 (N_17247,N_11609,N_12579);
xor U17248 (N_17248,N_11318,N_14656);
nand U17249 (N_17249,N_12113,N_13658);
xor U17250 (N_17250,N_10245,N_12972);
nand U17251 (N_17251,N_11839,N_12365);
nor U17252 (N_17252,N_11375,N_14120);
or U17253 (N_17253,N_14741,N_13022);
nand U17254 (N_17254,N_14708,N_14781);
xor U17255 (N_17255,N_12135,N_10916);
and U17256 (N_17256,N_14021,N_13575);
and U17257 (N_17257,N_13344,N_11879);
xor U17258 (N_17258,N_12107,N_14232);
or U17259 (N_17259,N_13487,N_10089);
nand U17260 (N_17260,N_14894,N_14372);
and U17261 (N_17261,N_13007,N_14013);
or U17262 (N_17262,N_11610,N_13695);
nor U17263 (N_17263,N_12748,N_14606);
nor U17264 (N_17264,N_13394,N_13026);
and U17265 (N_17265,N_14580,N_13264);
and U17266 (N_17266,N_11303,N_14393);
nor U17267 (N_17267,N_13353,N_13749);
and U17268 (N_17268,N_10601,N_11621);
nor U17269 (N_17269,N_10862,N_11949);
and U17270 (N_17270,N_12128,N_13311);
nor U17271 (N_17271,N_10746,N_14012);
nor U17272 (N_17272,N_12528,N_13437);
nor U17273 (N_17273,N_10437,N_10607);
nor U17274 (N_17274,N_14398,N_11345);
xnor U17275 (N_17275,N_13654,N_13841);
and U17276 (N_17276,N_10593,N_11217);
nor U17277 (N_17277,N_11939,N_14339);
or U17278 (N_17278,N_12342,N_14248);
nand U17279 (N_17279,N_13047,N_13137);
or U17280 (N_17280,N_12907,N_11947);
nor U17281 (N_17281,N_11021,N_13049);
or U17282 (N_17282,N_12481,N_14454);
or U17283 (N_17283,N_13298,N_12863);
nor U17284 (N_17284,N_12004,N_12112);
and U17285 (N_17285,N_10962,N_12252);
nor U17286 (N_17286,N_13104,N_13152);
xor U17287 (N_17287,N_11472,N_14908);
or U17288 (N_17288,N_10296,N_11335);
nor U17289 (N_17289,N_14102,N_12130);
nand U17290 (N_17290,N_14826,N_10068);
nand U17291 (N_17291,N_10583,N_10807);
or U17292 (N_17292,N_13624,N_10598);
xnor U17293 (N_17293,N_14890,N_13994);
nor U17294 (N_17294,N_14314,N_12550);
and U17295 (N_17295,N_13320,N_12308);
nor U17296 (N_17296,N_13934,N_14155);
and U17297 (N_17297,N_12867,N_10082);
nand U17298 (N_17298,N_10605,N_12132);
nand U17299 (N_17299,N_10100,N_12269);
nand U17300 (N_17300,N_12676,N_12932);
xor U17301 (N_17301,N_12850,N_10224);
or U17302 (N_17302,N_10567,N_10730);
or U17303 (N_17303,N_11327,N_10338);
nor U17304 (N_17304,N_11489,N_14968);
nand U17305 (N_17305,N_12633,N_11125);
nand U17306 (N_17306,N_11063,N_11268);
nand U17307 (N_17307,N_11387,N_10777);
or U17308 (N_17308,N_13650,N_10788);
and U17309 (N_17309,N_13328,N_13905);
or U17310 (N_17310,N_13440,N_12323);
and U17311 (N_17311,N_14168,N_14590);
or U17312 (N_17312,N_13291,N_12526);
and U17313 (N_17313,N_14161,N_11090);
nand U17314 (N_17314,N_11317,N_13041);
and U17315 (N_17315,N_13260,N_14307);
or U17316 (N_17316,N_10277,N_12337);
xor U17317 (N_17317,N_12100,N_14885);
nand U17318 (N_17318,N_11094,N_13660);
and U17319 (N_17319,N_10207,N_10825);
nor U17320 (N_17320,N_14088,N_10493);
nor U17321 (N_17321,N_12055,N_10579);
or U17322 (N_17322,N_11208,N_11745);
nor U17323 (N_17323,N_10706,N_10375);
or U17324 (N_17324,N_10162,N_11550);
and U17325 (N_17325,N_11802,N_13244);
nor U17326 (N_17326,N_11104,N_11057);
and U17327 (N_17327,N_12440,N_10878);
or U17328 (N_17328,N_10590,N_13249);
nand U17329 (N_17329,N_11716,N_11374);
or U17330 (N_17330,N_11756,N_13735);
or U17331 (N_17331,N_14757,N_14986);
and U17332 (N_17332,N_10465,N_14573);
or U17333 (N_17333,N_14808,N_10771);
nor U17334 (N_17334,N_10942,N_12371);
nand U17335 (N_17335,N_11236,N_13366);
nand U17336 (N_17336,N_11332,N_13266);
nor U17337 (N_17337,N_13704,N_14545);
and U17338 (N_17338,N_14160,N_13228);
nor U17339 (N_17339,N_11970,N_10191);
nor U17340 (N_17340,N_13036,N_12048);
nor U17341 (N_17341,N_14760,N_13876);
xnor U17342 (N_17342,N_11732,N_12525);
xor U17343 (N_17343,N_12879,N_14459);
nor U17344 (N_17344,N_12173,N_10356);
xor U17345 (N_17345,N_11296,N_14536);
nand U17346 (N_17346,N_14478,N_12422);
nand U17347 (N_17347,N_11060,N_11027);
nand U17348 (N_17348,N_12953,N_12296);
and U17349 (N_17349,N_13335,N_14858);
nor U17350 (N_17350,N_14530,N_10644);
or U17351 (N_17351,N_12340,N_13768);
and U17352 (N_17352,N_13211,N_10145);
nor U17353 (N_17353,N_14555,N_14230);
nand U17354 (N_17354,N_13648,N_12586);
and U17355 (N_17355,N_11034,N_10780);
nand U17356 (N_17356,N_13189,N_12360);
and U17357 (N_17357,N_10472,N_11510);
nand U17358 (N_17358,N_10209,N_12218);
nand U17359 (N_17359,N_12715,N_11827);
or U17360 (N_17360,N_12755,N_12213);
xor U17361 (N_17361,N_12143,N_10243);
or U17362 (N_17362,N_12513,N_13920);
xor U17363 (N_17363,N_12002,N_12636);
nand U17364 (N_17364,N_14583,N_14655);
and U17365 (N_17365,N_12007,N_11411);
and U17366 (N_17366,N_10109,N_11728);
or U17367 (N_17367,N_10793,N_11633);
xor U17368 (N_17368,N_14498,N_13058);
nand U17369 (N_17369,N_11783,N_11046);
nand U17370 (N_17370,N_10208,N_12225);
or U17371 (N_17371,N_12736,N_13693);
nor U17372 (N_17372,N_13854,N_14784);
xor U17373 (N_17373,N_11235,N_11010);
and U17374 (N_17374,N_14317,N_14824);
nor U17375 (N_17375,N_10257,N_12442);
xnor U17376 (N_17376,N_11834,N_14051);
nand U17377 (N_17377,N_13580,N_13285);
xor U17378 (N_17378,N_14525,N_12830);
and U17379 (N_17379,N_12764,N_13984);
or U17380 (N_17380,N_10184,N_12182);
nor U17381 (N_17381,N_14392,N_10367);
nand U17382 (N_17382,N_13262,N_11746);
nor U17383 (N_17383,N_13621,N_12254);
nand U17384 (N_17384,N_14286,N_11859);
and U17385 (N_17385,N_10556,N_14774);
nor U17386 (N_17386,N_13002,N_12681);
and U17387 (N_17387,N_13812,N_13006);
nand U17388 (N_17388,N_14503,N_12368);
and U17389 (N_17389,N_10467,N_12233);
and U17390 (N_17390,N_13201,N_11142);
nand U17391 (N_17391,N_10085,N_12429);
nor U17392 (N_17392,N_11735,N_14679);
nand U17393 (N_17393,N_12763,N_11619);
nand U17394 (N_17394,N_11251,N_12029);
and U17395 (N_17395,N_10808,N_13638);
nand U17396 (N_17396,N_13274,N_13840);
nor U17397 (N_17397,N_10371,N_14440);
nand U17398 (N_17398,N_13609,N_14213);
and U17399 (N_17399,N_13868,N_14832);
nand U17400 (N_17400,N_13675,N_12333);
nor U17401 (N_17401,N_12797,N_14076);
and U17402 (N_17402,N_11531,N_10425);
and U17403 (N_17403,N_12175,N_13339);
and U17404 (N_17404,N_13651,N_11384);
nand U17405 (N_17405,N_11017,N_13121);
xor U17406 (N_17406,N_13709,N_13943);
nor U17407 (N_17407,N_11405,N_14693);
and U17408 (N_17408,N_10958,N_12723);
or U17409 (N_17409,N_11137,N_13728);
nor U17410 (N_17410,N_10295,N_14981);
or U17411 (N_17411,N_11981,N_13643);
and U17412 (N_17412,N_10976,N_13468);
nand U17413 (N_17413,N_10308,N_14872);
nand U17414 (N_17414,N_11092,N_11571);
or U17415 (N_17415,N_12166,N_12350);
nand U17416 (N_17416,N_14772,N_14422);
nor U17417 (N_17417,N_12578,N_10670);
or U17418 (N_17418,N_14371,N_12430);
nor U17419 (N_17419,N_11103,N_13852);
and U17420 (N_17420,N_10433,N_11491);
xnor U17421 (N_17421,N_11373,N_14917);
or U17422 (N_17422,N_13573,N_13076);
xor U17423 (N_17423,N_12488,N_13219);
or U17424 (N_17424,N_12164,N_14126);
nand U17425 (N_17425,N_12190,N_12583);
nor U17426 (N_17426,N_14465,N_11180);
or U17427 (N_17427,N_11206,N_12761);
or U17428 (N_17428,N_13829,N_12902);
nand U17429 (N_17429,N_14090,N_13332);
nor U17430 (N_17430,N_12471,N_12678);
and U17431 (N_17431,N_12679,N_12496);
nor U17432 (N_17432,N_13186,N_13398);
nor U17433 (N_17433,N_11603,N_10242);
nand U17434 (N_17434,N_11535,N_13024);
nand U17435 (N_17435,N_11780,N_12517);
or U17436 (N_17436,N_14563,N_10737);
xnor U17437 (N_17437,N_12210,N_11058);
or U17438 (N_17438,N_14803,N_13314);
nand U17439 (N_17439,N_11983,N_11044);
or U17440 (N_17440,N_11197,N_11861);
or U17441 (N_17441,N_10480,N_12237);
or U17442 (N_17442,N_12595,N_14343);
and U17443 (N_17443,N_10786,N_11132);
nor U17444 (N_17444,N_13472,N_13504);
xor U17445 (N_17445,N_12058,N_13507);
nand U17446 (N_17446,N_10677,N_13360);
nand U17447 (N_17447,N_11456,N_10783);
or U17448 (N_17448,N_14324,N_14577);
and U17449 (N_17449,N_14785,N_14731);
and U17450 (N_17450,N_11765,N_14292);
nor U17451 (N_17451,N_12118,N_13331);
and U17452 (N_17452,N_10322,N_14318);
xnor U17453 (N_17453,N_14643,N_11589);
nor U17454 (N_17454,N_10992,N_10220);
or U17455 (N_17455,N_14948,N_13237);
nand U17456 (N_17456,N_14651,N_13409);
nor U17457 (N_17457,N_14069,N_14442);
nand U17458 (N_17458,N_11078,N_13779);
nor U17459 (N_17459,N_14494,N_11271);
nor U17460 (N_17460,N_11979,N_13571);
and U17461 (N_17461,N_12788,N_14951);
and U17462 (N_17462,N_10897,N_12415);
nand U17463 (N_17463,N_10871,N_10726);
nand U17464 (N_17464,N_14057,N_12732);
nor U17465 (N_17465,N_14289,N_13051);
nor U17466 (N_17466,N_11469,N_13806);
or U17467 (N_17467,N_11792,N_13563);
nor U17468 (N_17468,N_11107,N_13897);
nand U17469 (N_17469,N_11761,N_12447);
xor U17470 (N_17470,N_14947,N_13788);
nor U17471 (N_17471,N_10017,N_10421);
or U17472 (N_17472,N_14101,N_14548);
or U17473 (N_17473,N_11817,N_12289);
nand U17474 (N_17474,N_10215,N_12950);
nor U17475 (N_17475,N_13981,N_10523);
and U17476 (N_17476,N_10358,N_11426);
and U17477 (N_17477,N_12983,N_12685);
and U17478 (N_17478,N_14735,N_13881);
and U17479 (N_17479,N_14705,N_14321);
and U17480 (N_17480,N_10457,N_13974);
nor U17481 (N_17481,N_13098,N_13061);
nor U17482 (N_17482,N_14817,N_11467);
xor U17483 (N_17483,N_11095,N_13012);
nor U17484 (N_17484,N_14900,N_14288);
and U17485 (N_17485,N_10415,N_14241);
or U17486 (N_17486,N_13831,N_13450);
and U17487 (N_17487,N_10643,N_10851);
nor U17488 (N_17488,N_13593,N_13585);
nand U17489 (N_17489,N_13399,N_10501);
nor U17490 (N_17490,N_13018,N_12818);
or U17491 (N_17491,N_11890,N_10266);
nor U17492 (N_17492,N_11540,N_10149);
or U17493 (N_17493,N_12918,N_10728);
nor U17494 (N_17494,N_10198,N_10193);
nand U17495 (N_17495,N_11635,N_11138);
nand U17496 (N_17496,N_14173,N_12745);
and U17497 (N_17497,N_14627,N_13172);
or U17498 (N_17498,N_10660,N_10554);
or U17499 (N_17499,N_11157,N_11003);
nand U17500 (N_17500,N_10785,N_14543);
or U17501 (N_17501,N_10997,N_12897);
nand U17502 (N_17502,N_14904,N_14216);
and U17503 (N_17503,N_12564,N_12945);
nor U17504 (N_17504,N_10401,N_12993);
and U17505 (N_17505,N_14885,N_11887);
nand U17506 (N_17506,N_10809,N_11422);
xnor U17507 (N_17507,N_10761,N_12688);
xor U17508 (N_17508,N_10438,N_13856);
or U17509 (N_17509,N_11357,N_13395);
nand U17510 (N_17510,N_12512,N_14959);
nand U17511 (N_17511,N_12143,N_14973);
nand U17512 (N_17512,N_12037,N_12906);
nor U17513 (N_17513,N_13439,N_12960);
nand U17514 (N_17514,N_12567,N_14878);
nor U17515 (N_17515,N_13913,N_10605);
nand U17516 (N_17516,N_11549,N_10937);
and U17517 (N_17517,N_10323,N_13086);
nand U17518 (N_17518,N_11608,N_14684);
nor U17519 (N_17519,N_10395,N_11419);
nand U17520 (N_17520,N_14183,N_11960);
xnor U17521 (N_17521,N_14056,N_13637);
and U17522 (N_17522,N_12290,N_12017);
nor U17523 (N_17523,N_11483,N_10332);
and U17524 (N_17524,N_13197,N_12695);
and U17525 (N_17525,N_10452,N_10816);
nor U17526 (N_17526,N_12721,N_11848);
or U17527 (N_17527,N_14479,N_11414);
nand U17528 (N_17528,N_13120,N_11715);
nand U17529 (N_17529,N_13825,N_13161);
and U17530 (N_17530,N_10170,N_12194);
nor U17531 (N_17531,N_11683,N_12521);
nand U17532 (N_17532,N_11005,N_10794);
nand U17533 (N_17533,N_10872,N_12069);
nand U17534 (N_17534,N_11050,N_11905);
xor U17535 (N_17535,N_12293,N_14253);
nor U17536 (N_17536,N_11528,N_10312);
nand U17537 (N_17537,N_10851,N_10860);
or U17538 (N_17538,N_12736,N_10016);
and U17539 (N_17539,N_14354,N_10985);
nor U17540 (N_17540,N_13918,N_13163);
nor U17541 (N_17541,N_13149,N_14297);
nand U17542 (N_17542,N_10439,N_12337);
and U17543 (N_17543,N_12298,N_13338);
and U17544 (N_17544,N_11664,N_13780);
nor U17545 (N_17545,N_10400,N_12671);
or U17546 (N_17546,N_12925,N_10951);
and U17547 (N_17547,N_13308,N_14672);
and U17548 (N_17548,N_11881,N_11467);
nor U17549 (N_17549,N_13962,N_13519);
nand U17550 (N_17550,N_12030,N_10157);
nand U17551 (N_17551,N_10800,N_11137);
nor U17552 (N_17552,N_14521,N_12537);
or U17553 (N_17553,N_11663,N_14439);
nor U17554 (N_17554,N_12653,N_13707);
nor U17555 (N_17555,N_14986,N_12919);
nand U17556 (N_17556,N_10666,N_12054);
nor U17557 (N_17557,N_14821,N_11058);
and U17558 (N_17558,N_11552,N_11342);
nand U17559 (N_17559,N_11356,N_14898);
and U17560 (N_17560,N_10488,N_13807);
or U17561 (N_17561,N_11429,N_12974);
nor U17562 (N_17562,N_10998,N_13328);
nor U17563 (N_17563,N_13546,N_10745);
nor U17564 (N_17564,N_13294,N_14253);
xor U17565 (N_17565,N_12267,N_13459);
or U17566 (N_17566,N_13105,N_13891);
and U17567 (N_17567,N_11068,N_11495);
nor U17568 (N_17568,N_14665,N_12165);
xor U17569 (N_17569,N_10984,N_14800);
or U17570 (N_17570,N_13554,N_12033);
and U17571 (N_17571,N_12707,N_12049);
nor U17572 (N_17572,N_12498,N_11701);
and U17573 (N_17573,N_14798,N_12422);
nand U17574 (N_17574,N_10007,N_10888);
and U17575 (N_17575,N_11589,N_11308);
xnor U17576 (N_17576,N_11746,N_10218);
and U17577 (N_17577,N_14909,N_12935);
nor U17578 (N_17578,N_14833,N_14987);
or U17579 (N_17579,N_11977,N_14061);
nand U17580 (N_17580,N_14916,N_14320);
and U17581 (N_17581,N_12516,N_10666);
or U17582 (N_17582,N_14421,N_12077);
and U17583 (N_17583,N_11959,N_14928);
nor U17584 (N_17584,N_11790,N_13579);
xnor U17585 (N_17585,N_10959,N_12675);
nor U17586 (N_17586,N_12598,N_11662);
nand U17587 (N_17587,N_10392,N_14822);
nor U17588 (N_17588,N_10045,N_14976);
nand U17589 (N_17589,N_14387,N_12319);
nand U17590 (N_17590,N_11425,N_14093);
and U17591 (N_17591,N_10865,N_12619);
nand U17592 (N_17592,N_13066,N_10152);
nand U17593 (N_17593,N_14843,N_14970);
nor U17594 (N_17594,N_13321,N_12509);
and U17595 (N_17595,N_14929,N_14507);
nor U17596 (N_17596,N_12963,N_11781);
nor U17597 (N_17597,N_10532,N_13265);
or U17598 (N_17598,N_13121,N_13356);
or U17599 (N_17599,N_11750,N_12401);
nor U17600 (N_17600,N_10332,N_10929);
nor U17601 (N_17601,N_11238,N_13998);
or U17602 (N_17602,N_13220,N_11877);
nand U17603 (N_17603,N_11506,N_12210);
nor U17604 (N_17604,N_11291,N_13923);
and U17605 (N_17605,N_11124,N_13312);
or U17606 (N_17606,N_13480,N_14603);
nor U17607 (N_17607,N_11345,N_13328);
xnor U17608 (N_17608,N_10631,N_11731);
or U17609 (N_17609,N_10606,N_12581);
xnor U17610 (N_17610,N_14272,N_14473);
nand U17611 (N_17611,N_14592,N_10539);
nor U17612 (N_17612,N_11855,N_10763);
and U17613 (N_17613,N_11351,N_10509);
nor U17614 (N_17614,N_14974,N_10860);
nand U17615 (N_17615,N_11340,N_12003);
nand U17616 (N_17616,N_12594,N_10713);
or U17617 (N_17617,N_11432,N_13381);
nor U17618 (N_17618,N_14098,N_13998);
and U17619 (N_17619,N_14777,N_14631);
nand U17620 (N_17620,N_10314,N_11623);
xnor U17621 (N_17621,N_12211,N_13530);
nand U17622 (N_17622,N_14936,N_10266);
nand U17623 (N_17623,N_14921,N_14555);
and U17624 (N_17624,N_11860,N_12463);
nor U17625 (N_17625,N_11721,N_14715);
nand U17626 (N_17626,N_14272,N_11364);
nand U17627 (N_17627,N_12646,N_10917);
xnor U17628 (N_17628,N_14157,N_12319);
nor U17629 (N_17629,N_11578,N_10887);
or U17630 (N_17630,N_10991,N_12063);
and U17631 (N_17631,N_14716,N_11749);
or U17632 (N_17632,N_11693,N_13619);
or U17633 (N_17633,N_10493,N_12079);
xor U17634 (N_17634,N_12925,N_11110);
or U17635 (N_17635,N_10772,N_14817);
and U17636 (N_17636,N_12363,N_11237);
nand U17637 (N_17637,N_14980,N_12062);
nand U17638 (N_17638,N_10553,N_12184);
or U17639 (N_17639,N_13970,N_10903);
nand U17640 (N_17640,N_12479,N_14900);
nand U17641 (N_17641,N_12043,N_13624);
and U17642 (N_17642,N_10027,N_10649);
or U17643 (N_17643,N_12647,N_13871);
or U17644 (N_17644,N_13362,N_13673);
or U17645 (N_17645,N_14341,N_10435);
nand U17646 (N_17646,N_14947,N_14721);
and U17647 (N_17647,N_12937,N_14522);
nor U17648 (N_17648,N_10676,N_14256);
nand U17649 (N_17649,N_14016,N_11269);
and U17650 (N_17650,N_10951,N_10234);
and U17651 (N_17651,N_10912,N_11012);
or U17652 (N_17652,N_10538,N_13047);
nor U17653 (N_17653,N_10535,N_11788);
or U17654 (N_17654,N_13378,N_11855);
nand U17655 (N_17655,N_10633,N_12704);
and U17656 (N_17656,N_13570,N_13657);
and U17657 (N_17657,N_11248,N_13739);
or U17658 (N_17658,N_12189,N_11959);
or U17659 (N_17659,N_14151,N_10314);
nand U17660 (N_17660,N_14937,N_12692);
and U17661 (N_17661,N_14730,N_12180);
nor U17662 (N_17662,N_10226,N_14960);
and U17663 (N_17663,N_10484,N_11788);
xnor U17664 (N_17664,N_14064,N_13103);
or U17665 (N_17665,N_12426,N_13854);
nor U17666 (N_17666,N_14084,N_14948);
nor U17667 (N_17667,N_13164,N_11848);
and U17668 (N_17668,N_14049,N_11727);
and U17669 (N_17669,N_14075,N_13384);
or U17670 (N_17670,N_10759,N_14743);
or U17671 (N_17671,N_13527,N_12608);
nand U17672 (N_17672,N_14696,N_10153);
nand U17673 (N_17673,N_11558,N_12490);
nand U17674 (N_17674,N_10563,N_11160);
and U17675 (N_17675,N_14736,N_11786);
nand U17676 (N_17676,N_14028,N_14481);
or U17677 (N_17677,N_10243,N_14337);
xnor U17678 (N_17678,N_12952,N_14497);
or U17679 (N_17679,N_14466,N_14662);
or U17680 (N_17680,N_13440,N_11178);
nor U17681 (N_17681,N_10141,N_10301);
and U17682 (N_17682,N_10561,N_10678);
and U17683 (N_17683,N_11740,N_11803);
and U17684 (N_17684,N_10394,N_14341);
nand U17685 (N_17685,N_14002,N_11624);
nand U17686 (N_17686,N_13926,N_10415);
nor U17687 (N_17687,N_13806,N_12100);
or U17688 (N_17688,N_14479,N_14686);
nor U17689 (N_17689,N_12573,N_10330);
nand U17690 (N_17690,N_10742,N_12289);
nand U17691 (N_17691,N_10467,N_11972);
or U17692 (N_17692,N_13180,N_11725);
and U17693 (N_17693,N_11184,N_11888);
or U17694 (N_17694,N_11303,N_12711);
or U17695 (N_17695,N_13055,N_14107);
and U17696 (N_17696,N_11970,N_12265);
or U17697 (N_17697,N_12229,N_10830);
or U17698 (N_17698,N_11813,N_11500);
xnor U17699 (N_17699,N_13621,N_10332);
or U17700 (N_17700,N_14256,N_12143);
nand U17701 (N_17701,N_12480,N_14084);
and U17702 (N_17702,N_10215,N_13243);
or U17703 (N_17703,N_14479,N_12455);
and U17704 (N_17704,N_14235,N_10561);
or U17705 (N_17705,N_14683,N_14643);
nor U17706 (N_17706,N_10725,N_10586);
nand U17707 (N_17707,N_11938,N_10094);
or U17708 (N_17708,N_12791,N_12733);
nand U17709 (N_17709,N_10899,N_10631);
and U17710 (N_17710,N_10365,N_13699);
or U17711 (N_17711,N_11594,N_10741);
nand U17712 (N_17712,N_13015,N_14225);
xor U17713 (N_17713,N_10070,N_10638);
nor U17714 (N_17714,N_12941,N_10965);
nand U17715 (N_17715,N_14347,N_12870);
and U17716 (N_17716,N_14411,N_10638);
and U17717 (N_17717,N_12729,N_14242);
xnor U17718 (N_17718,N_12051,N_14522);
nor U17719 (N_17719,N_12836,N_10246);
or U17720 (N_17720,N_11480,N_11864);
or U17721 (N_17721,N_14228,N_12990);
nand U17722 (N_17722,N_10659,N_11732);
and U17723 (N_17723,N_11765,N_10172);
xor U17724 (N_17724,N_12781,N_13123);
nor U17725 (N_17725,N_14186,N_10399);
and U17726 (N_17726,N_14319,N_10226);
or U17727 (N_17727,N_10597,N_13988);
and U17728 (N_17728,N_10911,N_12074);
or U17729 (N_17729,N_14805,N_12903);
and U17730 (N_17730,N_12170,N_12342);
xor U17731 (N_17731,N_10324,N_10417);
or U17732 (N_17732,N_13706,N_12307);
and U17733 (N_17733,N_12768,N_12533);
or U17734 (N_17734,N_12899,N_10261);
nor U17735 (N_17735,N_12009,N_10826);
nor U17736 (N_17736,N_12568,N_11538);
xnor U17737 (N_17737,N_14699,N_13823);
or U17738 (N_17738,N_14735,N_10524);
nor U17739 (N_17739,N_14491,N_12804);
or U17740 (N_17740,N_12693,N_11691);
nor U17741 (N_17741,N_13182,N_13508);
and U17742 (N_17742,N_11814,N_12700);
and U17743 (N_17743,N_14275,N_11880);
and U17744 (N_17744,N_14850,N_10586);
nor U17745 (N_17745,N_12502,N_10379);
or U17746 (N_17746,N_14962,N_11956);
nor U17747 (N_17747,N_13851,N_10051);
nand U17748 (N_17748,N_11020,N_10649);
and U17749 (N_17749,N_11397,N_12976);
nand U17750 (N_17750,N_14091,N_10919);
nand U17751 (N_17751,N_13645,N_12842);
nand U17752 (N_17752,N_14679,N_13993);
nor U17753 (N_17753,N_13883,N_11358);
nand U17754 (N_17754,N_11706,N_11348);
and U17755 (N_17755,N_10761,N_10012);
nor U17756 (N_17756,N_14376,N_11508);
or U17757 (N_17757,N_12455,N_14355);
nor U17758 (N_17758,N_10895,N_13111);
xnor U17759 (N_17759,N_11284,N_12638);
nor U17760 (N_17760,N_13329,N_12231);
or U17761 (N_17761,N_12511,N_10065);
xnor U17762 (N_17762,N_14799,N_13769);
or U17763 (N_17763,N_11383,N_10480);
nor U17764 (N_17764,N_14444,N_13921);
nand U17765 (N_17765,N_14579,N_10143);
and U17766 (N_17766,N_13057,N_11089);
nor U17767 (N_17767,N_12148,N_10757);
or U17768 (N_17768,N_11223,N_10156);
and U17769 (N_17769,N_14441,N_11428);
and U17770 (N_17770,N_13924,N_11498);
or U17771 (N_17771,N_10979,N_11435);
nor U17772 (N_17772,N_11276,N_10484);
nor U17773 (N_17773,N_10318,N_13700);
and U17774 (N_17774,N_14360,N_13372);
or U17775 (N_17775,N_10828,N_10520);
or U17776 (N_17776,N_11358,N_10291);
xor U17777 (N_17777,N_12724,N_10876);
nor U17778 (N_17778,N_12049,N_14645);
or U17779 (N_17779,N_10910,N_13700);
and U17780 (N_17780,N_14489,N_11393);
or U17781 (N_17781,N_10337,N_14989);
nor U17782 (N_17782,N_10227,N_13527);
or U17783 (N_17783,N_10982,N_14316);
nand U17784 (N_17784,N_11191,N_12957);
and U17785 (N_17785,N_11913,N_13014);
nor U17786 (N_17786,N_14361,N_11289);
and U17787 (N_17787,N_11554,N_10622);
nand U17788 (N_17788,N_13161,N_11119);
or U17789 (N_17789,N_10025,N_11385);
nand U17790 (N_17790,N_12326,N_13981);
and U17791 (N_17791,N_13008,N_11254);
xnor U17792 (N_17792,N_11004,N_12390);
nor U17793 (N_17793,N_14316,N_11594);
xnor U17794 (N_17794,N_10027,N_10933);
and U17795 (N_17795,N_11845,N_13262);
nor U17796 (N_17796,N_13182,N_10565);
and U17797 (N_17797,N_14496,N_10284);
or U17798 (N_17798,N_10745,N_13793);
nand U17799 (N_17799,N_11957,N_10865);
and U17800 (N_17800,N_11487,N_10654);
nor U17801 (N_17801,N_12661,N_11970);
nand U17802 (N_17802,N_11199,N_12533);
nor U17803 (N_17803,N_11248,N_14786);
nor U17804 (N_17804,N_12150,N_13541);
xnor U17805 (N_17805,N_12909,N_14027);
and U17806 (N_17806,N_13275,N_11884);
xor U17807 (N_17807,N_13149,N_14410);
and U17808 (N_17808,N_12082,N_10528);
and U17809 (N_17809,N_10612,N_14885);
xor U17810 (N_17810,N_14111,N_10196);
and U17811 (N_17811,N_13634,N_10956);
nor U17812 (N_17812,N_13689,N_11040);
xor U17813 (N_17813,N_13463,N_11257);
and U17814 (N_17814,N_14599,N_11859);
nor U17815 (N_17815,N_14275,N_11388);
nand U17816 (N_17816,N_11500,N_12288);
and U17817 (N_17817,N_13281,N_11463);
nor U17818 (N_17818,N_11676,N_13991);
and U17819 (N_17819,N_10158,N_12171);
or U17820 (N_17820,N_11381,N_12091);
nor U17821 (N_17821,N_13503,N_10657);
nand U17822 (N_17822,N_12318,N_13341);
xnor U17823 (N_17823,N_11605,N_14738);
nand U17824 (N_17824,N_14779,N_13062);
nand U17825 (N_17825,N_10809,N_11722);
nor U17826 (N_17826,N_12991,N_14795);
nand U17827 (N_17827,N_13462,N_14951);
or U17828 (N_17828,N_14931,N_13957);
and U17829 (N_17829,N_14370,N_12213);
nand U17830 (N_17830,N_14632,N_11335);
or U17831 (N_17831,N_10374,N_10082);
or U17832 (N_17832,N_12143,N_12410);
xor U17833 (N_17833,N_14402,N_11224);
or U17834 (N_17834,N_10218,N_11200);
nor U17835 (N_17835,N_11312,N_11480);
xnor U17836 (N_17836,N_13415,N_11695);
or U17837 (N_17837,N_11046,N_14028);
nor U17838 (N_17838,N_12267,N_14104);
and U17839 (N_17839,N_14846,N_11419);
or U17840 (N_17840,N_14850,N_12175);
nand U17841 (N_17841,N_14034,N_12090);
xnor U17842 (N_17842,N_13984,N_10759);
or U17843 (N_17843,N_14581,N_14856);
nor U17844 (N_17844,N_13331,N_13703);
nand U17845 (N_17845,N_13435,N_10255);
and U17846 (N_17846,N_12581,N_14818);
nor U17847 (N_17847,N_10537,N_11376);
nand U17848 (N_17848,N_10030,N_11302);
xor U17849 (N_17849,N_13069,N_13327);
nand U17850 (N_17850,N_10835,N_10983);
nand U17851 (N_17851,N_10045,N_14043);
nand U17852 (N_17852,N_13212,N_13927);
or U17853 (N_17853,N_11978,N_14714);
or U17854 (N_17854,N_12930,N_13330);
and U17855 (N_17855,N_13937,N_12466);
nand U17856 (N_17856,N_12521,N_13258);
and U17857 (N_17857,N_13395,N_11301);
and U17858 (N_17858,N_10733,N_11326);
nand U17859 (N_17859,N_12808,N_10376);
and U17860 (N_17860,N_14824,N_12653);
nor U17861 (N_17861,N_12673,N_14093);
or U17862 (N_17862,N_11721,N_14269);
or U17863 (N_17863,N_11091,N_11343);
or U17864 (N_17864,N_13809,N_10772);
and U17865 (N_17865,N_10629,N_10388);
nand U17866 (N_17866,N_10809,N_12920);
nor U17867 (N_17867,N_11491,N_10735);
and U17868 (N_17868,N_13784,N_11749);
xor U17869 (N_17869,N_14473,N_11557);
nor U17870 (N_17870,N_13321,N_14257);
nor U17871 (N_17871,N_11443,N_11495);
and U17872 (N_17872,N_13505,N_10940);
nor U17873 (N_17873,N_10598,N_10156);
and U17874 (N_17874,N_11239,N_12098);
nor U17875 (N_17875,N_14705,N_12401);
nand U17876 (N_17876,N_12749,N_13095);
nand U17877 (N_17877,N_12075,N_14532);
nor U17878 (N_17878,N_10766,N_12349);
or U17879 (N_17879,N_12245,N_13993);
nor U17880 (N_17880,N_10414,N_13812);
or U17881 (N_17881,N_10465,N_10445);
and U17882 (N_17882,N_11958,N_11268);
nor U17883 (N_17883,N_10248,N_13638);
nand U17884 (N_17884,N_14185,N_10331);
nand U17885 (N_17885,N_13987,N_13670);
or U17886 (N_17886,N_12181,N_10495);
and U17887 (N_17887,N_13310,N_11007);
and U17888 (N_17888,N_10266,N_14458);
and U17889 (N_17889,N_10879,N_10230);
or U17890 (N_17890,N_13962,N_13657);
nand U17891 (N_17891,N_10110,N_10654);
or U17892 (N_17892,N_13739,N_10429);
or U17893 (N_17893,N_12400,N_10412);
or U17894 (N_17894,N_14557,N_14106);
nand U17895 (N_17895,N_13926,N_10259);
nor U17896 (N_17896,N_11760,N_10775);
nand U17897 (N_17897,N_14048,N_12728);
or U17898 (N_17898,N_13251,N_13064);
nand U17899 (N_17899,N_11349,N_14866);
or U17900 (N_17900,N_14319,N_12616);
and U17901 (N_17901,N_12447,N_13458);
and U17902 (N_17902,N_10303,N_10944);
nand U17903 (N_17903,N_10155,N_11819);
xnor U17904 (N_17904,N_13806,N_14116);
xnor U17905 (N_17905,N_11275,N_13849);
or U17906 (N_17906,N_11436,N_14179);
nand U17907 (N_17907,N_14272,N_14648);
and U17908 (N_17908,N_10835,N_13954);
or U17909 (N_17909,N_14814,N_12205);
nand U17910 (N_17910,N_14287,N_14418);
nor U17911 (N_17911,N_13569,N_14099);
or U17912 (N_17912,N_13205,N_12871);
or U17913 (N_17913,N_12021,N_12130);
or U17914 (N_17914,N_11469,N_10427);
nor U17915 (N_17915,N_12954,N_14740);
or U17916 (N_17916,N_10876,N_14768);
and U17917 (N_17917,N_14284,N_10705);
nor U17918 (N_17918,N_10834,N_11783);
or U17919 (N_17919,N_12573,N_10466);
nor U17920 (N_17920,N_11703,N_10087);
nor U17921 (N_17921,N_10778,N_12808);
nor U17922 (N_17922,N_12152,N_13426);
nor U17923 (N_17923,N_14193,N_10369);
or U17924 (N_17924,N_13030,N_10816);
and U17925 (N_17925,N_14045,N_13804);
or U17926 (N_17926,N_10203,N_14958);
xnor U17927 (N_17927,N_13508,N_14727);
and U17928 (N_17928,N_11928,N_10677);
and U17929 (N_17929,N_14778,N_14577);
nand U17930 (N_17930,N_13919,N_11321);
and U17931 (N_17931,N_13464,N_11365);
xnor U17932 (N_17932,N_10546,N_11184);
or U17933 (N_17933,N_12819,N_11589);
nand U17934 (N_17934,N_12753,N_14801);
nand U17935 (N_17935,N_12102,N_12257);
nand U17936 (N_17936,N_14772,N_13409);
or U17937 (N_17937,N_14501,N_13093);
and U17938 (N_17938,N_14939,N_14528);
or U17939 (N_17939,N_10710,N_12129);
and U17940 (N_17940,N_11114,N_14470);
xor U17941 (N_17941,N_10836,N_12764);
nor U17942 (N_17942,N_12380,N_11599);
nand U17943 (N_17943,N_14503,N_12249);
and U17944 (N_17944,N_10818,N_11384);
nor U17945 (N_17945,N_14432,N_12969);
nor U17946 (N_17946,N_10664,N_14449);
or U17947 (N_17947,N_11564,N_11058);
and U17948 (N_17948,N_10527,N_14667);
and U17949 (N_17949,N_11108,N_12817);
nand U17950 (N_17950,N_11565,N_10133);
or U17951 (N_17951,N_10516,N_13121);
nor U17952 (N_17952,N_11514,N_14350);
or U17953 (N_17953,N_11185,N_14776);
and U17954 (N_17954,N_12151,N_11000);
nand U17955 (N_17955,N_14868,N_11578);
and U17956 (N_17956,N_10644,N_11653);
or U17957 (N_17957,N_11848,N_11948);
nand U17958 (N_17958,N_13277,N_14873);
nor U17959 (N_17959,N_10561,N_13349);
nand U17960 (N_17960,N_10375,N_14420);
and U17961 (N_17961,N_13585,N_13252);
nor U17962 (N_17962,N_10191,N_12057);
nand U17963 (N_17963,N_12429,N_11834);
nor U17964 (N_17964,N_14243,N_13625);
nand U17965 (N_17965,N_10651,N_12274);
or U17966 (N_17966,N_11833,N_13088);
nand U17967 (N_17967,N_12599,N_13272);
and U17968 (N_17968,N_14866,N_10551);
nor U17969 (N_17969,N_13067,N_13641);
or U17970 (N_17970,N_10258,N_11486);
or U17971 (N_17971,N_13619,N_14649);
nand U17972 (N_17972,N_11867,N_11057);
and U17973 (N_17973,N_14445,N_14488);
and U17974 (N_17974,N_12514,N_12493);
and U17975 (N_17975,N_11696,N_11158);
nand U17976 (N_17976,N_11677,N_10731);
nor U17977 (N_17977,N_11871,N_10520);
nand U17978 (N_17978,N_12450,N_13806);
or U17979 (N_17979,N_12738,N_14265);
nand U17980 (N_17980,N_13942,N_14346);
nor U17981 (N_17981,N_13675,N_14695);
xor U17982 (N_17982,N_12588,N_14721);
or U17983 (N_17983,N_11822,N_11430);
or U17984 (N_17984,N_11127,N_11908);
nor U17985 (N_17985,N_14501,N_13167);
nand U17986 (N_17986,N_14254,N_12403);
nor U17987 (N_17987,N_10883,N_14084);
nor U17988 (N_17988,N_12645,N_10543);
nor U17989 (N_17989,N_12709,N_10124);
nand U17990 (N_17990,N_14641,N_10824);
and U17991 (N_17991,N_11378,N_12164);
xor U17992 (N_17992,N_10622,N_14900);
and U17993 (N_17993,N_12158,N_10816);
nand U17994 (N_17994,N_14566,N_11922);
nand U17995 (N_17995,N_10342,N_10459);
nor U17996 (N_17996,N_14936,N_11842);
nand U17997 (N_17997,N_14510,N_13196);
nand U17998 (N_17998,N_10673,N_14418);
nand U17999 (N_17999,N_13525,N_13065);
nand U18000 (N_18000,N_11063,N_13460);
nor U18001 (N_18001,N_10579,N_13895);
or U18002 (N_18002,N_11135,N_10121);
nor U18003 (N_18003,N_11212,N_13221);
or U18004 (N_18004,N_11683,N_10405);
nand U18005 (N_18005,N_10912,N_12399);
and U18006 (N_18006,N_14331,N_10062);
or U18007 (N_18007,N_14020,N_14843);
or U18008 (N_18008,N_12706,N_10912);
nand U18009 (N_18009,N_10952,N_12134);
nand U18010 (N_18010,N_12146,N_11173);
nand U18011 (N_18011,N_11138,N_10716);
xnor U18012 (N_18012,N_10870,N_11534);
nand U18013 (N_18013,N_12262,N_12246);
xor U18014 (N_18014,N_12441,N_14567);
and U18015 (N_18015,N_10762,N_14765);
nor U18016 (N_18016,N_11942,N_12868);
nand U18017 (N_18017,N_13830,N_13837);
xor U18018 (N_18018,N_12288,N_12769);
or U18019 (N_18019,N_10540,N_11509);
xnor U18020 (N_18020,N_12681,N_12578);
nor U18021 (N_18021,N_11008,N_13933);
nand U18022 (N_18022,N_12346,N_14546);
nor U18023 (N_18023,N_13472,N_11268);
or U18024 (N_18024,N_14838,N_10454);
xor U18025 (N_18025,N_10623,N_11171);
nor U18026 (N_18026,N_12952,N_11552);
xnor U18027 (N_18027,N_12069,N_11037);
nor U18028 (N_18028,N_14542,N_11876);
or U18029 (N_18029,N_11143,N_10718);
or U18030 (N_18030,N_11787,N_13381);
or U18031 (N_18031,N_13558,N_11689);
xnor U18032 (N_18032,N_13909,N_10067);
nor U18033 (N_18033,N_13828,N_12204);
xnor U18034 (N_18034,N_14925,N_10851);
xnor U18035 (N_18035,N_13721,N_11304);
nand U18036 (N_18036,N_14161,N_13402);
nor U18037 (N_18037,N_14196,N_14263);
or U18038 (N_18038,N_12198,N_14210);
xor U18039 (N_18039,N_11237,N_13709);
nand U18040 (N_18040,N_13018,N_13738);
nand U18041 (N_18041,N_11892,N_10019);
xnor U18042 (N_18042,N_14380,N_12687);
nor U18043 (N_18043,N_14631,N_10520);
nand U18044 (N_18044,N_13570,N_11810);
nand U18045 (N_18045,N_13616,N_14471);
and U18046 (N_18046,N_12582,N_11027);
xor U18047 (N_18047,N_10404,N_13587);
nand U18048 (N_18048,N_14859,N_14002);
nor U18049 (N_18049,N_12214,N_10390);
or U18050 (N_18050,N_10982,N_14788);
nand U18051 (N_18051,N_10603,N_12478);
or U18052 (N_18052,N_14683,N_14175);
or U18053 (N_18053,N_10866,N_13626);
nand U18054 (N_18054,N_14419,N_13076);
or U18055 (N_18055,N_13353,N_13528);
nor U18056 (N_18056,N_10607,N_12648);
nand U18057 (N_18057,N_14327,N_12632);
nor U18058 (N_18058,N_12405,N_13787);
nand U18059 (N_18059,N_12867,N_10716);
nor U18060 (N_18060,N_11205,N_12538);
xnor U18061 (N_18061,N_12785,N_11219);
xnor U18062 (N_18062,N_12629,N_10382);
or U18063 (N_18063,N_10689,N_12456);
nor U18064 (N_18064,N_13295,N_14446);
and U18065 (N_18065,N_11171,N_12895);
nand U18066 (N_18066,N_14662,N_12419);
nand U18067 (N_18067,N_12231,N_12988);
nor U18068 (N_18068,N_13921,N_12019);
or U18069 (N_18069,N_14877,N_11532);
nand U18070 (N_18070,N_11513,N_13556);
or U18071 (N_18071,N_14004,N_10619);
and U18072 (N_18072,N_11704,N_10208);
or U18073 (N_18073,N_10247,N_10622);
and U18074 (N_18074,N_11486,N_10256);
nor U18075 (N_18075,N_12202,N_12255);
or U18076 (N_18076,N_13132,N_12200);
nand U18077 (N_18077,N_10978,N_13874);
nor U18078 (N_18078,N_11070,N_12012);
and U18079 (N_18079,N_12338,N_12342);
and U18080 (N_18080,N_13008,N_10301);
nor U18081 (N_18081,N_14680,N_11105);
and U18082 (N_18082,N_12083,N_11013);
nand U18083 (N_18083,N_11257,N_14387);
nor U18084 (N_18084,N_13862,N_12925);
nor U18085 (N_18085,N_13658,N_13220);
xor U18086 (N_18086,N_10569,N_11561);
nor U18087 (N_18087,N_10154,N_12239);
xnor U18088 (N_18088,N_11526,N_13657);
or U18089 (N_18089,N_13041,N_11598);
nor U18090 (N_18090,N_13789,N_12226);
and U18091 (N_18091,N_10811,N_12110);
nand U18092 (N_18092,N_14916,N_13939);
and U18093 (N_18093,N_10424,N_14420);
nor U18094 (N_18094,N_11657,N_10212);
nor U18095 (N_18095,N_14645,N_12485);
and U18096 (N_18096,N_14169,N_13375);
nor U18097 (N_18097,N_11554,N_12513);
or U18098 (N_18098,N_14736,N_11763);
xor U18099 (N_18099,N_11918,N_12012);
nor U18100 (N_18100,N_12567,N_14976);
xnor U18101 (N_18101,N_11212,N_13414);
nor U18102 (N_18102,N_12687,N_11744);
nor U18103 (N_18103,N_11575,N_13545);
xor U18104 (N_18104,N_14548,N_13338);
and U18105 (N_18105,N_13434,N_13102);
or U18106 (N_18106,N_12820,N_12382);
nor U18107 (N_18107,N_10129,N_14741);
and U18108 (N_18108,N_13431,N_12044);
and U18109 (N_18109,N_11599,N_14905);
and U18110 (N_18110,N_10624,N_12122);
xnor U18111 (N_18111,N_13671,N_10866);
xnor U18112 (N_18112,N_12487,N_11302);
nand U18113 (N_18113,N_10455,N_11872);
nor U18114 (N_18114,N_12177,N_12114);
and U18115 (N_18115,N_12041,N_14360);
nor U18116 (N_18116,N_13034,N_13409);
nor U18117 (N_18117,N_14561,N_12155);
or U18118 (N_18118,N_12809,N_13256);
nor U18119 (N_18119,N_14127,N_12696);
nand U18120 (N_18120,N_13111,N_11334);
or U18121 (N_18121,N_11348,N_14834);
nand U18122 (N_18122,N_11148,N_11411);
and U18123 (N_18123,N_13036,N_14969);
xnor U18124 (N_18124,N_10707,N_14042);
nand U18125 (N_18125,N_10842,N_14692);
nand U18126 (N_18126,N_11091,N_13335);
nand U18127 (N_18127,N_13989,N_11532);
or U18128 (N_18128,N_14804,N_12914);
or U18129 (N_18129,N_14865,N_14659);
nor U18130 (N_18130,N_12210,N_14451);
nor U18131 (N_18131,N_14422,N_13612);
or U18132 (N_18132,N_14874,N_11527);
or U18133 (N_18133,N_13767,N_11600);
xor U18134 (N_18134,N_12238,N_11901);
nand U18135 (N_18135,N_14313,N_13370);
nand U18136 (N_18136,N_14671,N_10764);
or U18137 (N_18137,N_14176,N_10726);
nand U18138 (N_18138,N_11769,N_11867);
or U18139 (N_18139,N_12751,N_12721);
and U18140 (N_18140,N_12743,N_14717);
xnor U18141 (N_18141,N_14885,N_10087);
and U18142 (N_18142,N_12026,N_14401);
or U18143 (N_18143,N_14657,N_14853);
nor U18144 (N_18144,N_11122,N_11026);
nor U18145 (N_18145,N_13713,N_11315);
or U18146 (N_18146,N_14672,N_13414);
xor U18147 (N_18147,N_13894,N_13304);
nand U18148 (N_18148,N_10725,N_13949);
nand U18149 (N_18149,N_11439,N_12871);
xor U18150 (N_18150,N_14796,N_11229);
or U18151 (N_18151,N_14147,N_12102);
nor U18152 (N_18152,N_14293,N_11910);
and U18153 (N_18153,N_13471,N_13766);
nand U18154 (N_18154,N_11474,N_12774);
nor U18155 (N_18155,N_10729,N_10055);
and U18156 (N_18156,N_10048,N_12703);
nand U18157 (N_18157,N_13743,N_12254);
nor U18158 (N_18158,N_12389,N_11821);
nor U18159 (N_18159,N_10231,N_12981);
xnor U18160 (N_18160,N_13490,N_14195);
nor U18161 (N_18161,N_10121,N_12339);
nor U18162 (N_18162,N_10368,N_14043);
and U18163 (N_18163,N_13111,N_13228);
nand U18164 (N_18164,N_13678,N_14313);
xor U18165 (N_18165,N_12138,N_11197);
nand U18166 (N_18166,N_11302,N_13640);
nand U18167 (N_18167,N_13097,N_11968);
or U18168 (N_18168,N_14056,N_12067);
nand U18169 (N_18169,N_12108,N_12744);
or U18170 (N_18170,N_10963,N_13900);
nand U18171 (N_18171,N_11365,N_10734);
nor U18172 (N_18172,N_14269,N_14595);
and U18173 (N_18173,N_11967,N_14658);
and U18174 (N_18174,N_13212,N_10266);
nand U18175 (N_18175,N_14241,N_13519);
and U18176 (N_18176,N_13195,N_12958);
xnor U18177 (N_18177,N_11920,N_10219);
and U18178 (N_18178,N_14052,N_14454);
nor U18179 (N_18179,N_14616,N_10194);
and U18180 (N_18180,N_13726,N_14774);
and U18181 (N_18181,N_12697,N_14714);
nor U18182 (N_18182,N_12839,N_11006);
and U18183 (N_18183,N_11309,N_11406);
xor U18184 (N_18184,N_10895,N_10840);
and U18185 (N_18185,N_12804,N_11856);
or U18186 (N_18186,N_14040,N_10049);
nand U18187 (N_18187,N_14821,N_12611);
nor U18188 (N_18188,N_12037,N_12043);
and U18189 (N_18189,N_11483,N_12361);
nor U18190 (N_18190,N_10796,N_11958);
nor U18191 (N_18191,N_10314,N_13765);
nor U18192 (N_18192,N_12570,N_11373);
and U18193 (N_18193,N_14849,N_10912);
nor U18194 (N_18194,N_11072,N_11608);
or U18195 (N_18195,N_14716,N_11615);
nand U18196 (N_18196,N_12875,N_12979);
and U18197 (N_18197,N_14954,N_12097);
or U18198 (N_18198,N_11682,N_13544);
or U18199 (N_18199,N_14420,N_10259);
or U18200 (N_18200,N_14546,N_10254);
xnor U18201 (N_18201,N_12854,N_13362);
nand U18202 (N_18202,N_13657,N_13722);
nor U18203 (N_18203,N_12452,N_11590);
and U18204 (N_18204,N_13679,N_11393);
or U18205 (N_18205,N_13866,N_10232);
nor U18206 (N_18206,N_11640,N_14238);
and U18207 (N_18207,N_11852,N_14599);
nand U18208 (N_18208,N_12471,N_10480);
nand U18209 (N_18209,N_10463,N_12806);
or U18210 (N_18210,N_12202,N_14810);
and U18211 (N_18211,N_14626,N_14801);
xnor U18212 (N_18212,N_14350,N_10526);
nor U18213 (N_18213,N_14931,N_13618);
nor U18214 (N_18214,N_13809,N_13001);
nor U18215 (N_18215,N_14925,N_12782);
nor U18216 (N_18216,N_11210,N_13123);
xor U18217 (N_18217,N_11122,N_13606);
xnor U18218 (N_18218,N_13842,N_10354);
and U18219 (N_18219,N_11124,N_12646);
or U18220 (N_18220,N_11471,N_14842);
or U18221 (N_18221,N_11905,N_13590);
or U18222 (N_18222,N_12256,N_11891);
nand U18223 (N_18223,N_13931,N_11390);
and U18224 (N_18224,N_13901,N_14354);
xor U18225 (N_18225,N_10757,N_11045);
nor U18226 (N_18226,N_10950,N_10936);
and U18227 (N_18227,N_14210,N_14711);
nand U18228 (N_18228,N_14830,N_13781);
or U18229 (N_18229,N_14730,N_14725);
nor U18230 (N_18230,N_14230,N_14040);
nor U18231 (N_18231,N_10831,N_12479);
and U18232 (N_18232,N_12504,N_10146);
nand U18233 (N_18233,N_11842,N_11699);
nor U18234 (N_18234,N_13960,N_11500);
and U18235 (N_18235,N_11924,N_12094);
or U18236 (N_18236,N_12772,N_13610);
nor U18237 (N_18237,N_11203,N_10942);
nand U18238 (N_18238,N_11743,N_11562);
xor U18239 (N_18239,N_11687,N_13454);
xor U18240 (N_18240,N_14298,N_12660);
or U18241 (N_18241,N_11637,N_10956);
or U18242 (N_18242,N_11865,N_14918);
nor U18243 (N_18243,N_10365,N_14946);
and U18244 (N_18244,N_10065,N_14847);
nor U18245 (N_18245,N_12167,N_11058);
nor U18246 (N_18246,N_12523,N_11113);
nand U18247 (N_18247,N_10190,N_11550);
or U18248 (N_18248,N_10081,N_13820);
and U18249 (N_18249,N_12702,N_13051);
nor U18250 (N_18250,N_11215,N_13739);
nor U18251 (N_18251,N_12208,N_12791);
or U18252 (N_18252,N_12490,N_11618);
nor U18253 (N_18253,N_10233,N_10113);
or U18254 (N_18254,N_13351,N_10379);
xnor U18255 (N_18255,N_14025,N_10197);
xor U18256 (N_18256,N_13404,N_13093);
and U18257 (N_18257,N_14340,N_13372);
nand U18258 (N_18258,N_10399,N_14297);
or U18259 (N_18259,N_12580,N_12581);
and U18260 (N_18260,N_10068,N_13313);
nor U18261 (N_18261,N_14811,N_11762);
and U18262 (N_18262,N_13851,N_11762);
or U18263 (N_18263,N_12273,N_14395);
or U18264 (N_18264,N_12045,N_14175);
and U18265 (N_18265,N_10802,N_11870);
nand U18266 (N_18266,N_11378,N_11871);
or U18267 (N_18267,N_12056,N_10685);
nand U18268 (N_18268,N_14160,N_13883);
or U18269 (N_18269,N_12983,N_13245);
xnor U18270 (N_18270,N_10445,N_11750);
and U18271 (N_18271,N_10849,N_13707);
nor U18272 (N_18272,N_11232,N_13463);
or U18273 (N_18273,N_10068,N_14803);
and U18274 (N_18274,N_11493,N_14571);
nand U18275 (N_18275,N_11757,N_11412);
xor U18276 (N_18276,N_13445,N_13596);
nand U18277 (N_18277,N_13383,N_14790);
or U18278 (N_18278,N_11577,N_10546);
or U18279 (N_18279,N_10753,N_14603);
xnor U18280 (N_18280,N_11859,N_10799);
nor U18281 (N_18281,N_10610,N_10993);
nand U18282 (N_18282,N_11763,N_10474);
nor U18283 (N_18283,N_13538,N_10941);
nand U18284 (N_18284,N_13863,N_11693);
or U18285 (N_18285,N_12075,N_13279);
and U18286 (N_18286,N_10309,N_10681);
nor U18287 (N_18287,N_11491,N_12257);
nand U18288 (N_18288,N_10228,N_13585);
or U18289 (N_18289,N_11539,N_13746);
and U18290 (N_18290,N_11774,N_14966);
or U18291 (N_18291,N_13930,N_10645);
and U18292 (N_18292,N_11435,N_12316);
nor U18293 (N_18293,N_10813,N_13924);
nand U18294 (N_18294,N_10543,N_10427);
xnor U18295 (N_18295,N_13402,N_11898);
nand U18296 (N_18296,N_12215,N_14738);
xor U18297 (N_18297,N_14798,N_10440);
xor U18298 (N_18298,N_14879,N_13025);
nand U18299 (N_18299,N_11094,N_13872);
or U18300 (N_18300,N_10017,N_13831);
nand U18301 (N_18301,N_10298,N_14389);
or U18302 (N_18302,N_13685,N_12279);
nor U18303 (N_18303,N_13811,N_13064);
and U18304 (N_18304,N_10911,N_10926);
nand U18305 (N_18305,N_13280,N_13650);
nor U18306 (N_18306,N_12973,N_13725);
or U18307 (N_18307,N_13038,N_10976);
and U18308 (N_18308,N_13111,N_12401);
and U18309 (N_18309,N_14714,N_13789);
and U18310 (N_18310,N_11457,N_13332);
and U18311 (N_18311,N_10161,N_12112);
and U18312 (N_18312,N_11619,N_14077);
and U18313 (N_18313,N_10781,N_10240);
and U18314 (N_18314,N_12817,N_12700);
nor U18315 (N_18315,N_14717,N_14608);
nor U18316 (N_18316,N_14170,N_13108);
nand U18317 (N_18317,N_12382,N_14045);
and U18318 (N_18318,N_10370,N_10857);
nand U18319 (N_18319,N_12990,N_13315);
nand U18320 (N_18320,N_10205,N_10107);
and U18321 (N_18321,N_13741,N_13880);
and U18322 (N_18322,N_10069,N_12557);
or U18323 (N_18323,N_12814,N_10547);
or U18324 (N_18324,N_11295,N_10472);
xnor U18325 (N_18325,N_11050,N_14778);
or U18326 (N_18326,N_12104,N_11263);
nand U18327 (N_18327,N_11054,N_12274);
nand U18328 (N_18328,N_14935,N_10464);
nor U18329 (N_18329,N_14089,N_13881);
or U18330 (N_18330,N_13522,N_12137);
or U18331 (N_18331,N_14570,N_10178);
nand U18332 (N_18332,N_10575,N_12113);
nor U18333 (N_18333,N_10623,N_12259);
nor U18334 (N_18334,N_12576,N_14463);
nor U18335 (N_18335,N_12150,N_11070);
nand U18336 (N_18336,N_13052,N_12557);
nand U18337 (N_18337,N_14593,N_11797);
or U18338 (N_18338,N_10787,N_10991);
xnor U18339 (N_18339,N_11627,N_11976);
and U18340 (N_18340,N_11648,N_10571);
nand U18341 (N_18341,N_11456,N_14261);
or U18342 (N_18342,N_13560,N_12409);
xor U18343 (N_18343,N_13422,N_14572);
nor U18344 (N_18344,N_13919,N_10497);
nor U18345 (N_18345,N_10850,N_11362);
nand U18346 (N_18346,N_12364,N_10530);
nor U18347 (N_18347,N_13314,N_11184);
and U18348 (N_18348,N_10741,N_13971);
nand U18349 (N_18349,N_10829,N_14376);
and U18350 (N_18350,N_13278,N_11594);
nor U18351 (N_18351,N_11401,N_12780);
and U18352 (N_18352,N_10271,N_11003);
nor U18353 (N_18353,N_10537,N_14340);
xnor U18354 (N_18354,N_12590,N_10287);
and U18355 (N_18355,N_10494,N_11277);
nor U18356 (N_18356,N_14955,N_12162);
nor U18357 (N_18357,N_14665,N_10388);
or U18358 (N_18358,N_12470,N_13558);
xor U18359 (N_18359,N_12343,N_11399);
nand U18360 (N_18360,N_13404,N_10027);
nor U18361 (N_18361,N_12615,N_11453);
and U18362 (N_18362,N_11535,N_11860);
nor U18363 (N_18363,N_14250,N_10562);
xor U18364 (N_18364,N_10584,N_13559);
nor U18365 (N_18365,N_10943,N_14846);
or U18366 (N_18366,N_14206,N_12996);
and U18367 (N_18367,N_10192,N_11607);
or U18368 (N_18368,N_10518,N_11796);
nand U18369 (N_18369,N_10989,N_12704);
nand U18370 (N_18370,N_10166,N_14228);
nand U18371 (N_18371,N_14554,N_10962);
nor U18372 (N_18372,N_11681,N_10059);
nor U18373 (N_18373,N_13081,N_12279);
nor U18374 (N_18374,N_13624,N_12113);
and U18375 (N_18375,N_12759,N_11984);
or U18376 (N_18376,N_12198,N_10494);
or U18377 (N_18377,N_13788,N_10133);
nor U18378 (N_18378,N_11163,N_12328);
and U18379 (N_18379,N_13800,N_12953);
and U18380 (N_18380,N_10803,N_14525);
or U18381 (N_18381,N_14193,N_14527);
and U18382 (N_18382,N_12687,N_13169);
nand U18383 (N_18383,N_11006,N_14033);
nand U18384 (N_18384,N_14069,N_11525);
or U18385 (N_18385,N_10287,N_11932);
nand U18386 (N_18386,N_14453,N_14767);
or U18387 (N_18387,N_14225,N_10687);
or U18388 (N_18388,N_14976,N_12219);
nand U18389 (N_18389,N_13126,N_13352);
or U18390 (N_18390,N_11732,N_11834);
xnor U18391 (N_18391,N_10591,N_13353);
nor U18392 (N_18392,N_14860,N_13773);
or U18393 (N_18393,N_12894,N_11507);
and U18394 (N_18394,N_11453,N_10601);
or U18395 (N_18395,N_14187,N_14411);
nand U18396 (N_18396,N_11553,N_13226);
nand U18397 (N_18397,N_14938,N_13265);
nor U18398 (N_18398,N_13926,N_10617);
and U18399 (N_18399,N_13283,N_13058);
or U18400 (N_18400,N_12016,N_12036);
or U18401 (N_18401,N_11388,N_14080);
nand U18402 (N_18402,N_14628,N_13737);
nor U18403 (N_18403,N_13708,N_13821);
xor U18404 (N_18404,N_14730,N_10496);
and U18405 (N_18405,N_14031,N_13310);
nor U18406 (N_18406,N_11884,N_13378);
nor U18407 (N_18407,N_14140,N_10327);
and U18408 (N_18408,N_11591,N_11747);
nor U18409 (N_18409,N_12380,N_11059);
nor U18410 (N_18410,N_14074,N_13859);
and U18411 (N_18411,N_14282,N_13450);
nand U18412 (N_18412,N_11997,N_11092);
nor U18413 (N_18413,N_11453,N_11559);
nand U18414 (N_18414,N_10087,N_12328);
nor U18415 (N_18415,N_11196,N_13697);
nor U18416 (N_18416,N_10635,N_12400);
and U18417 (N_18417,N_14287,N_10555);
nand U18418 (N_18418,N_10016,N_13305);
nor U18419 (N_18419,N_12341,N_13313);
or U18420 (N_18420,N_13491,N_14327);
and U18421 (N_18421,N_12558,N_14129);
nand U18422 (N_18422,N_11305,N_10428);
or U18423 (N_18423,N_13534,N_11028);
or U18424 (N_18424,N_13149,N_14753);
and U18425 (N_18425,N_12316,N_14138);
nor U18426 (N_18426,N_12185,N_10851);
and U18427 (N_18427,N_12157,N_12769);
nand U18428 (N_18428,N_14813,N_11361);
or U18429 (N_18429,N_14883,N_10454);
nand U18430 (N_18430,N_12540,N_14025);
or U18431 (N_18431,N_14910,N_13839);
or U18432 (N_18432,N_14248,N_13094);
and U18433 (N_18433,N_11125,N_10711);
or U18434 (N_18434,N_14903,N_13754);
nand U18435 (N_18435,N_13623,N_14133);
and U18436 (N_18436,N_11856,N_14179);
and U18437 (N_18437,N_11474,N_11450);
nand U18438 (N_18438,N_13515,N_14593);
nand U18439 (N_18439,N_14918,N_10398);
nand U18440 (N_18440,N_14037,N_10919);
nand U18441 (N_18441,N_10760,N_11123);
and U18442 (N_18442,N_11101,N_12768);
or U18443 (N_18443,N_14027,N_14168);
nand U18444 (N_18444,N_12809,N_13783);
or U18445 (N_18445,N_10915,N_13313);
and U18446 (N_18446,N_14550,N_13834);
xnor U18447 (N_18447,N_10059,N_13686);
xor U18448 (N_18448,N_11359,N_11177);
nor U18449 (N_18449,N_14008,N_14878);
xnor U18450 (N_18450,N_14428,N_13162);
nor U18451 (N_18451,N_14792,N_10920);
nor U18452 (N_18452,N_13147,N_14937);
xor U18453 (N_18453,N_11922,N_12267);
nand U18454 (N_18454,N_10641,N_14881);
or U18455 (N_18455,N_14296,N_12365);
and U18456 (N_18456,N_14295,N_11117);
or U18457 (N_18457,N_12677,N_13398);
and U18458 (N_18458,N_11763,N_13236);
nor U18459 (N_18459,N_11607,N_12755);
and U18460 (N_18460,N_13948,N_11663);
nand U18461 (N_18461,N_10801,N_11980);
nor U18462 (N_18462,N_14085,N_11903);
nor U18463 (N_18463,N_13262,N_11357);
nor U18464 (N_18464,N_10582,N_12180);
or U18465 (N_18465,N_10832,N_13930);
or U18466 (N_18466,N_14895,N_13781);
or U18467 (N_18467,N_10906,N_12214);
nor U18468 (N_18468,N_11885,N_11404);
or U18469 (N_18469,N_12492,N_10455);
or U18470 (N_18470,N_11306,N_13859);
nand U18471 (N_18471,N_11635,N_14312);
and U18472 (N_18472,N_13947,N_14310);
nor U18473 (N_18473,N_10806,N_12941);
and U18474 (N_18474,N_13942,N_13452);
nor U18475 (N_18475,N_11131,N_12420);
nor U18476 (N_18476,N_14220,N_10015);
nand U18477 (N_18477,N_13937,N_12006);
or U18478 (N_18478,N_14959,N_11031);
nand U18479 (N_18479,N_14031,N_12087);
and U18480 (N_18480,N_10841,N_14580);
and U18481 (N_18481,N_13686,N_11267);
xor U18482 (N_18482,N_13249,N_11009);
nand U18483 (N_18483,N_14551,N_11407);
xnor U18484 (N_18484,N_12048,N_10690);
or U18485 (N_18485,N_11996,N_14910);
and U18486 (N_18486,N_13796,N_13987);
nand U18487 (N_18487,N_11192,N_10086);
nand U18488 (N_18488,N_11447,N_14080);
nor U18489 (N_18489,N_14769,N_14057);
nand U18490 (N_18490,N_12949,N_12740);
nand U18491 (N_18491,N_12267,N_11786);
and U18492 (N_18492,N_12717,N_13611);
nand U18493 (N_18493,N_12288,N_11024);
xnor U18494 (N_18494,N_13303,N_12676);
nand U18495 (N_18495,N_10512,N_11618);
or U18496 (N_18496,N_11301,N_14550);
nor U18497 (N_18497,N_14685,N_13549);
or U18498 (N_18498,N_14707,N_14704);
nor U18499 (N_18499,N_10139,N_13834);
and U18500 (N_18500,N_12839,N_10470);
nor U18501 (N_18501,N_12455,N_12324);
and U18502 (N_18502,N_13545,N_14782);
nor U18503 (N_18503,N_11477,N_13586);
nand U18504 (N_18504,N_12988,N_14628);
or U18505 (N_18505,N_13548,N_11591);
nor U18506 (N_18506,N_11199,N_14266);
or U18507 (N_18507,N_12209,N_10891);
and U18508 (N_18508,N_14376,N_12981);
nand U18509 (N_18509,N_12782,N_14154);
nor U18510 (N_18510,N_11137,N_10213);
nor U18511 (N_18511,N_10588,N_13420);
and U18512 (N_18512,N_14966,N_12504);
nor U18513 (N_18513,N_14546,N_14846);
or U18514 (N_18514,N_10059,N_14400);
nand U18515 (N_18515,N_12150,N_12302);
nand U18516 (N_18516,N_13671,N_12337);
nor U18517 (N_18517,N_14916,N_10477);
or U18518 (N_18518,N_11837,N_10864);
nor U18519 (N_18519,N_13963,N_10235);
nand U18520 (N_18520,N_13545,N_13976);
nor U18521 (N_18521,N_10820,N_10289);
xor U18522 (N_18522,N_10026,N_10900);
or U18523 (N_18523,N_10639,N_12107);
or U18524 (N_18524,N_10060,N_11812);
and U18525 (N_18525,N_12686,N_11067);
nand U18526 (N_18526,N_11965,N_12248);
nand U18527 (N_18527,N_10652,N_12540);
and U18528 (N_18528,N_14952,N_14175);
nand U18529 (N_18529,N_11735,N_12514);
nand U18530 (N_18530,N_14767,N_14511);
nor U18531 (N_18531,N_13783,N_14735);
and U18532 (N_18532,N_10053,N_12182);
and U18533 (N_18533,N_11847,N_10627);
nand U18534 (N_18534,N_11283,N_10696);
or U18535 (N_18535,N_12991,N_10469);
xnor U18536 (N_18536,N_10615,N_14855);
and U18537 (N_18537,N_12036,N_14004);
nor U18538 (N_18538,N_10160,N_13420);
and U18539 (N_18539,N_13366,N_12719);
and U18540 (N_18540,N_11752,N_13685);
nor U18541 (N_18541,N_12052,N_13067);
nor U18542 (N_18542,N_12272,N_13137);
nor U18543 (N_18543,N_14440,N_10488);
nor U18544 (N_18544,N_10007,N_13291);
and U18545 (N_18545,N_14423,N_10477);
nor U18546 (N_18546,N_11033,N_10769);
nand U18547 (N_18547,N_11689,N_13258);
and U18548 (N_18548,N_11570,N_13825);
or U18549 (N_18549,N_14937,N_12704);
and U18550 (N_18550,N_13729,N_14778);
xnor U18551 (N_18551,N_14512,N_12274);
xor U18552 (N_18552,N_11640,N_14436);
xnor U18553 (N_18553,N_10786,N_11609);
or U18554 (N_18554,N_10821,N_13378);
and U18555 (N_18555,N_11956,N_14777);
nor U18556 (N_18556,N_12745,N_13606);
or U18557 (N_18557,N_11688,N_11103);
nor U18558 (N_18558,N_14051,N_13381);
and U18559 (N_18559,N_12550,N_12771);
and U18560 (N_18560,N_10240,N_12271);
or U18561 (N_18561,N_11749,N_14108);
nor U18562 (N_18562,N_10798,N_13640);
nand U18563 (N_18563,N_14108,N_14994);
nand U18564 (N_18564,N_11551,N_14517);
nand U18565 (N_18565,N_11768,N_11247);
or U18566 (N_18566,N_12691,N_12853);
or U18567 (N_18567,N_14098,N_11059);
nand U18568 (N_18568,N_14353,N_14655);
nand U18569 (N_18569,N_13186,N_13394);
nor U18570 (N_18570,N_14239,N_11629);
xor U18571 (N_18571,N_12162,N_13447);
or U18572 (N_18572,N_10265,N_14926);
and U18573 (N_18573,N_14873,N_13888);
xnor U18574 (N_18574,N_14925,N_10364);
and U18575 (N_18575,N_13752,N_14742);
nor U18576 (N_18576,N_11434,N_14384);
nor U18577 (N_18577,N_12325,N_11680);
or U18578 (N_18578,N_11524,N_12494);
nand U18579 (N_18579,N_14012,N_14455);
xnor U18580 (N_18580,N_10949,N_11762);
and U18581 (N_18581,N_14897,N_11885);
nor U18582 (N_18582,N_13562,N_14157);
nor U18583 (N_18583,N_12188,N_14469);
nand U18584 (N_18584,N_13565,N_10720);
nor U18585 (N_18585,N_11826,N_10873);
nand U18586 (N_18586,N_12210,N_13785);
or U18587 (N_18587,N_13430,N_11913);
nor U18588 (N_18588,N_13578,N_10884);
xor U18589 (N_18589,N_10529,N_14958);
nor U18590 (N_18590,N_10661,N_13756);
nor U18591 (N_18591,N_10247,N_12464);
nand U18592 (N_18592,N_10697,N_12259);
or U18593 (N_18593,N_11819,N_13535);
nor U18594 (N_18594,N_13439,N_13948);
or U18595 (N_18595,N_13357,N_14874);
nor U18596 (N_18596,N_11949,N_13017);
nor U18597 (N_18597,N_14092,N_12513);
or U18598 (N_18598,N_10749,N_11571);
and U18599 (N_18599,N_12636,N_13464);
nor U18600 (N_18600,N_13290,N_12901);
nand U18601 (N_18601,N_10605,N_14630);
xnor U18602 (N_18602,N_11996,N_13651);
nor U18603 (N_18603,N_12352,N_10782);
nor U18604 (N_18604,N_11586,N_11381);
or U18605 (N_18605,N_11587,N_10917);
or U18606 (N_18606,N_14018,N_11447);
and U18607 (N_18607,N_14766,N_11924);
nor U18608 (N_18608,N_13080,N_13949);
and U18609 (N_18609,N_13957,N_13420);
nand U18610 (N_18610,N_13897,N_10336);
nor U18611 (N_18611,N_13807,N_13518);
or U18612 (N_18612,N_11116,N_12940);
nand U18613 (N_18613,N_13512,N_11726);
and U18614 (N_18614,N_10931,N_11186);
xor U18615 (N_18615,N_14205,N_13446);
nand U18616 (N_18616,N_13097,N_12326);
or U18617 (N_18617,N_10283,N_10636);
or U18618 (N_18618,N_14672,N_14698);
or U18619 (N_18619,N_11867,N_13812);
nor U18620 (N_18620,N_14351,N_13240);
nand U18621 (N_18621,N_14172,N_11479);
nand U18622 (N_18622,N_11436,N_14104);
or U18623 (N_18623,N_14392,N_14240);
xor U18624 (N_18624,N_10794,N_13835);
nor U18625 (N_18625,N_10440,N_13326);
or U18626 (N_18626,N_14258,N_10567);
nor U18627 (N_18627,N_12849,N_11397);
and U18628 (N_18628,N_14127,N_13706);
nor U18629 (N_18629,N_12829,N_12035);
xnor U18630 (N_18630,N_10333,N_14712);
and U18631 (N_18631,N_10807,N_10224);
and U18632 (N_18632,N_14314,N_12989);
xnor U18633 (N_18633,N_10246,N_14146);
or U18634 (N_18634,N_14948,N_13078);
nor U18635 (N_18635,N_10900,N_10446);
nor U18636 (N_18636,N_11476,N_10346);
and U18637 (N_18637,N_12898,N_13574);
nand U18638 (N_18638,N_11549,N_10967);
or U18639 (N_18639,N_13296,N_14193);
and U18640 (N_18640,N_13014,N_11874);
nand U18641 (N_18641,N_10420,N_11381);
or U18642 (N_18642,N_12252,N_13726);
or U18643 (N_18643,N_12868,N_13781);
and U18644 (N_18644,N_12498,N_12314);
nand U18645 (N_18645,N_12045,N_12893);
nand U18646 (N_18646,N_10867,N_11688);
or U18647 (N_18647,N_12402,N_14115);
and U18648 (N_18648,N_10664,N_10103);
and U18649 (N_18649,N_13965,N_14487);
or U18650 (N_18650,N_11979,N_14386);
and U18651 (N_18651,N_13642,N_11481);
and U18652 (N_18652,N_12596,N_10349);
or U18653 (N_18653,N_12881,N_11024);
and U18654 (N_18654,N_12214,N_12909);
nor U18655 (N_18655,N_11288,N_11546);
nor U18656 (N_18656,N_14855,N_10268);
xnor U18657 (N_18657,N_11374,N_13446);
or U18658 (N_18658,N_11991,N_11095);
xor U18659 (N_18659,N_10042,N_13926);
nand U18660 (N_18660,N_14672,N_13535);
nor U18661 (N_18661,N_12828,N_10339);
and U18662 (N_18662,N_10701,N_11666);
nor U18663 (N_18663,N_11452,N_11574);
or U18664 (N_18664,N_14254,N_13053);
or U18665 (N_18665,N_12176,N_12057);
or U18666 (N_18666,N_10664,N_14607);
or U18667 (N_18667,N_12612,N_12724);
or U18668 (N_18668,N_11106,N_13330);
or U18669 (N_18669,N_11836,N_12063);
nand U18670 (N_18670,N_13272,N_13821);
or U18671 (N_18671,N_12651,N_14605);
nand U18672 (N_18672,N_13022,N_14190);
nor U18673 (N_18673,N_14791,N_11305);
or U18674 (N_18674,N_10902,N_13839);
or U18675 (N_18675,N_14584,N_13862);
or U18676 (N_18676,N_13719,N_13162);
and U18677 (N_18677,N_14360,N_10954);
nand U18678 (N_18678,N_12213,N_10234);
and U18679 (N_18679,N_14355,N_10759);
nand U18680 (N_18680,N_14619,N_12544);
nor U18681 (N_18681,N_12780,N_12913);
xnor U18682 (N_18682,N_12677,N_11017);
nand U18683 (N_18683,N_12524,N_11021);
or U18684 (N_18684,N_11399,N_14855);
and U18685 (N_18685,N_12159,N_10380);
and U18686 (N_18686,N_14619,N_13257);
nand U18687 (N_18687,N_14020,N_12980);
nor U18688 (N_18688,N_13639,N_13105);
nand U18689 (N_18689,N_11205,N_12173);
and U18690 (N_18690,N_14557,N_13753);
nor U18691 (N_18691,N_11776,N_12106);
nor U18692 (N_18692,N_11401,N_10807);
and U18693 (N_18693,N_11264,N_14882);
or U18694 (N_18694,N_10364,N_10934);
or U18695 (N_18695,N_12452,N_12532);
or U18696 (N_18696,N_11367,N_13274);
nor U18697 (N_18697,N_10190,N_14108);
nand U18698 (N_18698,N_10447,N_12104);
or U18699 (N_18699,N_13156,N_10439);
nor U18700 (N_18700,N_12210,N_13133);
nand U18701 (N_18701,N_14588,N_13386);
or U18702 (N_18702,N_10185,N_11237);
or U18703 (N_18703,N_12518,N_11782);
xnor U18704 (N_18704,N_11307,N_11494);
or U18705 (N_18705,N_10541,N_14716);
and U18706 (N_18706,N_13282,N_11383);
and U18707 (N_18707,N_14544,N_13748);
xnor U18708 (N_18708,N_11723,N_10406);
or U18709 (N_18709,N_10714,N_14109);
nor U18710 (N_18710,N_11198,N_13364);
xor U18711 (N_18711,N_14277,N_12504);
or U18712 (N_18712,N_14330,N_12018);
nand U18713 (N_18713,N_10878,N_11138);
xnor U18714 (N_18714,N_13476,N_13875);
nand U18715 (N_18715,N_13400,N_11882);
xor U18716 (N_18716,N_14457,N_14962);
or U18717 (N_18717,N_10064,N_14884);
and U18718 (N_18718,N_10530,N_10676);
or U18719 (N_18719,N_10704,N_12258);
nand U18720 (N_18720,N_14159,N_13736);
nand U18721 (N_18721,N_14726,N_14633);
nand U18722 (N_18722,N_10478,N_12929);
nor U18723 (N_18723,N_11849,N_11313);
and U18724 (N_18724,N_12232,N_12498);
or U18725 (N_18725,N_14807,N_13086);
and U18726 (N_18726,N_13911,N_12889);
or U18727 (N_18727,N_10792,N_13993);
or U18728 (N_18728,N_10636,N_14133);
or U18729 (N_18729,N_14939,N_14089);
nor U18730 (N_18730,N_13674,N_10132);
or U18731 (N_18731,N_10745,N_13223);
and U18732 (N_18732,N_12863,N_10659);
xnor U18733 (N_18733,N_11196,N_11538);
nor U18734 (N_18734,N_10689,N_13404);
nand U18735 (N_18735,N_13459,N_10098);
nand U18736 (N_18736,N_11499,N_14619);
nand U18737 (N_18737,N_14237,N_10433);
and U18738 (N_18738,N_10785,N_12621);
or U18739 (N_18739,N_12309,N_14045);
or U18740 (N_18740,N_10521,N_12314);
nor U18741 (N_18741,N_12241,N_13494);
nand U18742 (N_18742,N_13585,N_13901);
nor U18743 (N_18743,N_14464,N_13178);
nor U18744 (N_18744,N_14517,N_11603);
and U18745 (N_18745,N_12432,N_12248);
or U18746 (N_18746,N_14524,N_10983);
xor U18747 (N_18747,N_10313,N_13835);
or U18748 (N_18748,N_14196,N_14588);
and U18749 (N_18749,N_14210,N_11560);
or U18750 (N_18750,N_13392,N_10170);
or U18751 (N_18751,N_11821,N_11087);
and U18752 (N_18752,N_14710,N_14819);
nand U18753 (N_18753,N_11006,N_12531);
or U18754 (N_18754,N_11612,N_10421);
nand U18755 (N_18755,N_14847,N_13761);
or U18756 (N_18756,N_11708,N_10661);
nor U18757 (N_18757,N_13976,N_11046);
or U18758 (N_18758,N_13411,N_10827);
xnor U18759 (N_18759,N_14691,N_13954);
or U18760 (N_18760,N_14751,N_12544);
nor U18761 (N_18761,N_11045,N_11492);
and U18762 (N_18762,N_12385,N_13493);
nor U18763 (N_18763,N_13743,N_13680);
nand U18764 (N_18764,N_14201,N_11177);
or U18765 (N_18765,N_10956,N_14464);
nor U18766 (N_18766,N_10976,N_12618);
or U18767 (N_18767,N_10107,N_13329);
nor U18768 (N_18768,N_13651,N_10554);
and U18769 (N_18769,N_11306,N_12247);
and U18770 (N_18770,N_13766,N_12730);
and U18771 (N_18771,N_13138,N_14816);
or U18772 (N_18772,N_11500,N_13621);
and U18773 (N_18773,N_12581,N_11916);
nor U18774 (N_18774,N_12705,N_10257);
nor U18775 (N_18775,N_10794,N_12807);
nor U18776 (N_18776,N_11432,N_11867);
nand U18777 (N_18777,N_14877,N_12690);
nand U18778 (N_18778,N_11640,N_13120);
and U18779 (N_18779,N_11315,N_11492);
or U18780 (N_18780,N_13423,N_14980);
nor U18781 (N_18781,N_12255,N_12759);
and U18782 (N_18782,N_13743,N_11022);
or U18783 (N_18783,N_12216,N_10194);
and U18784 (N_18784,N_12692,N_14582);
and U18785 (N_18785,N_13045,N_14116);
or U18786 (N_18786,N_12957,N_10967);
nand U18787 (N_18787,N_12172,N_12767);
nand U18788 (N_18788,N_10586,N_14431);
xor U18789 (N_18789,N_11204,N_10319);
or U18790 (N_18790,N_11627,N_11519);
nand U18791 (N_18791,N_11436,N_11319);
and U18792 (N_18792,N_11710,N_10563);
nor U18793 (N_18793,N_10013,N_13445);
nor U18794 (N_18794,N_12993,N_12390);
nand U18795 (N_18795,N_11184,N_11203);
nand U18796 (N_18796,N_14184,N_10431);
and U18797 (N_18797,N_11433,N_11274);
or U18798 (N_18798,N_13651,N_11438);
nand U18799 (N_18799,N_13037,N_11920);
nor U18800 (N_18800,N_12270,N_14213);
nor U18801 (N_18801,N_11368,N_12961);
nand U18802 (N_18802,N_13404,N_11853);
nor U18803 (N_18803,N_12415,N_11064);
and U18804 (N_18804,N_12769,N_12134);
and U18805 (N_18805,N_14664,N_14997);
or U18806 (N_18806,N_14509,N_14162);
and U18807 (N_18807,N_12946,N_14092);
nor U18808 (N_18808,N_14218,N_11218);
and U18809 (N_18809,N_11231,N_10533);
nand U18810 (N_18810,N_12576,N_14773);
and U18811 (N_18811,N_14494,N_12089);
or U18812 (N_18812,N_12323,N_10177);
and U18813 (N_18813,N_11395,N_13160);
and U18814 (N_18814,N_11132,N_12682);
nor U18815 (N_18815,N_12251,N_10039);
and U18816 (N_18816,N_10631,N_11471);
nand U18817 (N_18817,N_11736,N_11079);
or U18818 (N_18818,N_10944,N_11293);
and U18819 (N_18819,N_13668,N_13867);
or U18820 (N_18820,N_14895,N_11359);
nand U18821 (N_18821,N_13982,N_12016);
and U18822 (N_18822,N_10745,N_11558);
nand U18823 (N_18823,N_14489,N_14708);
or U18824 (N_18824,N_12933,N_14397);
nor U18825 (N_18825,N_11026,N_13817);
nor U18826 (N_18826,N_13188,N_13919);
nand U18827 (N_18827,N_10187,N_11399);
nand U18828 (N_18828,N_11517,N_14408);
nor U18829 (N_18829,N_13780,N_10121);
nand U18830 (N_18830,N_10581,N_11169);
nor U18831 (N_18831,N_10031,N_10007);
or U18832 (N_18832,N_13092,N_14115);
nand U18833 (N_18833,N_14735,N_10610);
nor U18834 (N_18834,N_12642,N_11451);
xor U18835 (N_18835,N_10860,N_12682);
nand U18836 (N_18836,N_10813,N_10469);
or U18837 (N_18837,N_14467,N_10861);
and U18838 (N_18838,N_14182,N_12175);
or U18839 (N_18839,N_10918,N_14621);
and U18840 (N_18840,N_11156,N_11348);
and U18841 (N_18841,N_11822,N_14657);
nand U18842 (N_18842,N_12831,N_14401);
nand U18843 (N_18843,N_11961,N_10476);
nor U18844 (N_18844,N_13193,N_11486);
or U18845 (N_18845,N_10803,N_11189);
and U18846 (N_18846,N_13916,N_11618);
and U18847 (N_18847,N_14493,N_10839);
and U18848 (N_18848,N_14990,N_14098);
nand U18849 (N_18849,N_12370,N_11421);
xnor U18850 (N_18850,N_10514,N_12693);
or U18851 (N_18851,N_12264,N_14826);
nor U18852 (N_18852,N_13535,N_11161);
and U18853 (N_18853,N_12362,N_11430);
and U18854 (N_18854,N_10455,N_13025);
nand U18855 (N_18855,N_12103,N_14563);
and U18856 (N_18856,N_13316,N_13103);
or U18857 (N_18857,N_14949,N_10973);
or U18858 (N_18858,N_10605,N_11501);
or U18859 (N_18859,N_11806,N_13479);
and U18860 (N_18860,N_12771,N_14039);
nor U18861 (N_18861,N_13471,N_14883);
and U18862 (N_18862,N_11915,N_12492);
or U18863 (N_18863,N_10479,N_14696);
nand U18864 (N_18864,N_14866,N_11342);
or U18865 (N_18865,N_10500,N_11948);
nor U18866 (N_18866,N_14421,N_10867);
nor U18867 (N_18867,N_13144,N_10964);
or U18868 (N_18868,N_10130,N_14156);
and U18869 (N_18869,N_14906,N_12581);
nor U18870 (N_18870,N_11321,N_10844);
nand U18871 (N_18871,N_13952,N_14292);
nor U18872 (N_18872,N_10374,N_13757);
nor U18873 (N_18873,N_12133,N_13503);
nor U18874 (N_18874,N_12073,N_10957);
nor U18875 (N_18875,N_13920,N_14677);
and U18876 (N_18876,N_13544,N_13994);
xor U18877 (N_18877,N_10947,N_11331);
nor U18878 (N_18878,N_10256,N_10820);
and U18879 (N_18879,N_11718,N_13820);
nor U18880 (N_18880,N_14711,N_14563);
nand U18881 (N_18881,N_13271,N_10662);
or U18882 (N_18882,N_11538,N_11054);
and U18883 (N_18883,N_12818,N_13692);
nor U18884 (N_18884,N_14937,N_12188);
nor U18885 (N_18885,N_14678,N_14639);
nor U18886 (N_18886,N_14064,N_14947);
and U18887 (N_18887,N_11944,N_12732);
or U18888 (N_18888,N_10893,N_10338);
or U18889 (N_18889,N_13670,N_13422);
or U18890 (N_18890,N_11924,N_13186);
or U18891 (N_18891,N_11755,N_13275);
nand U18892 (N_18892,N_13504,N_11867);
nand U18893 (N_18893,N_11508,N_11313);
and U18894 (N_18894,N_10458,N_14586);
xnor U18895 (N_18895,N_10378,N_12200);
nand U18896 (N_18896,N_11018,N_14435);
nand U18897 (N_18897,N_12356,N_12816);
nor U18898 (N_18898,N_13517,N_14179);
or U18899 (N_18899,N_12036,N_10605);
xor U18900 (N_18900,N_11334,N_11260);
nand U18901 (N_18901,N_14101,N_10989);
and U18902 (N_18902,N_10720,N_13321);
or U18903 (N_18903,N_11953,N_12369);
nand U18904 (N_18904,N_12716,N_10191);
or U18905 (N_18905,N_13328,N_12832);
nand U18906 (N_18906,N_10595,N_12078);
nand U18907 (N_18907,N_10847,N_13269);
and U18908 (N_18908,N_12873,N_10833);
xor U18909 (N_18909,N_10389,N_13333);
and U18910 (N_18910,N_12141,N_11853);
and U18911 (N_18911,N_13310,N_14992);
nor U18912 (N_18912,N_13854,N_13594);
nand U18913 (N_18913,N_13818,N_11370);
and U18914 (N_18914,N_13150,N_13129);
xor U18915 (N_18915,N_14306,N_10903);
xnor U18916 (N_18916,N_12870,N_14205);
nand U18917 (N_18917,N_14307,N_10269);
nand U18918 (N_18918,N_10249,N_14342);
nand U18919 (N_18919,N_11736,N_10337);
nor U18920 (N_18920,N_12854,N_11100);
nand U18921 (N_18921,N_14527,N_13876);
and U18922 (N_18922,N_13200,N_14203);
xnor U18923 (N_18923,N_14211,N_12961);
xnor U18924 (N_18924,N_11609,N_12205);
xnor U18925 (N_18925,N_14360,N_14173);
and U18926 (N_18926,N_11019,N_10841);
or U18927 (N_18927,N_14975,N_11623);
nor U18928 (N_18928,N_10286,N_13843);
and U18929 (N_18929,N_14431,N_13484);
nor U18930 (N_18930,N_10618,N_13288);
nand U18931 (N_18931,N_14901,N_11635);
or U18932 (N_18932,N_12308,N_13325);
nor U18933 (N_18933,N_10130,N_11647);
or U18934 (N_18934,N_10835,N_14033);
and U18935 (N_18935,N_10370,N_14743);
and U18936 (N_18936,N_14465,N_12129);
or U18937 (N_18937,N_10340,N_13718);
nand U18938 (N_18938,N_14389,N_13257);
nand U18939 (N_18939,N_14377,N_13663);
and U18940 (N_18940,N_10545,N_10551);
xnor U18941 (N_18941,N_12715,N_10316);
nor U18942 (N_18942,N_14500,N_10662);
nand U18943 (N_18943,N_10067,N_13573);
nand U18944 (N_18944,N_14881,N_11358);
or U18945 (N_18945,N_14610,N_11667);
nand U18946 (N_18946,N_10796,N_12339);
nor U18947 (N_18947,N_11540,N_10866);
and U18948 (N_18948,N_11968,N_12225);
nand U18949 (N_18949,N_10203,N_10273);
or U18950 (N_18950,N_11050,N_12138);
nand U18951 (N_18951,N_11965,N_13196);
nand U18952 (N_18952,N_10173,N_12746);
nor U18953 (N_18953,N_13457,N_10636);
xnor U18954 (N_18954,N_12400,N_14933);
or U18955 (N_18955,N_13944,N_13077);
and U18956 (N_18956,N_12716,N_11683);
and U18957 (N_18957,N_14125,N_11280);
or U18958 (N_18958,N_13675,N_12639);
nor U18959 (N_18959,N_11569,N_14301);
xor U18960 (N_18960,N_10181,N_11104);
and U18961 (N_18961,N_13204,N_13814);
or U18962 (N_18962,N_10366,N_14994);
and U18963 (N_18963,N_14663,N_11297);
nor U18964 (N_18964,N_13428,N_12942);
nand U18965 (N_18965,N_11167,N_13095);
and U18966 (N_18966,N_14894,N_13109);
or U18967 (N_18967,N_14396,N_12066);
or U18968 (N_18968,N_12478,N_10882);
or U18969 (N_18969,N_10578,N_11580);
nand U18970 (N_18970,N_10772,N_10283);
or U18971 (N_18971,N_11291,N_10018);
nor U18972 (N_18972,N_14235,N_10874);
nand U18973 (N_18973,N_11457,N_10938);
or U18974 (N_18974,N_14038,N_13907);
nand U18975 (N_18975,N_11986,N_12629);
nand U18976 (N_18976,N_12140,N_13721);
nand U18977 (N_18977,N_10278,N_10675);
nand U18978 (N_18978,N_12799,N_12944);
or U18979 (N_18979,N_10132,N_13412);
or U18980 (N_18980,N_10916,N_11399);
nor U18981 (N_18981,N_14583,N_11794);
nor U18982 (N_18982,N_13520,N_13385);
nor U18983 (N_18983,N_14201,N_14422);
nor U18984 (N_18984,N_13782,N_11147);
nand U18985 (N_18985,N_12995,N_10107);
and U18986 (N_18986,N_11187,N_11906);
and U18987 (N_18987,N_13510,N_10527);
nand U18988 (N_18988,N_14990,N_12672);
xnor U18989 (N_18989,N_12718,N_14824);
nor U18990 (N_18990,N_12714,N_11356);
or U18991 (N_18991,N_10434,N_12216);
nand U18992 (N_18992,N_12245,N_13846);
or U18993 (N_18993,N_12584,N_11957);
and U18994 (N_18994,N_13394,N_10944);
nand U18995 (N_18995,N_10363,N_13001);
nor U18996 (N_18996,N_12956,N_14220);
nor U18997 (N_18997,N_10329,N_14460);
and U18998 (N_18998,N_11059,N_11157);
nand U18999 (N_18999,N_14265,N_14969);
and U19000 (N_19000,N_10299,N_10059);
nand U19001 (N_19001,N_12425,N_14310);
nor U19002 (N_19002,N_13250,N_13179);
or U19003 (N_19003,N_12156,N_14812);
or U19004 (N_19004,N_13439,N_10099);
nand U19005 (N_19005,N_14250,N_11544);
nor U19006 (N_19006,N_13832,N_14526);
or U19007 (N_19007,N_14276,N_14549);
or U19008 (N_19008,N_14422,N_13591);
xor U19009 (N_19009,N_12888,N_13949);
nand U19010 (N_19010,N_12135,N_12251);
nand U19011 (N_19011,N_13150,N_13098);
and U19012 (N_19012,N_12981,N_12036);
and U19013 (N_19013,N_14918,N_14336);
nor U19014 (N_19014,N_13184,N_10791);
nor U19015 (N_19015,N_13969,N_12118);
nand U19016 (N_19016,N_13345,N_10829);
nand U19017 (N_19017,N_14398,N_13779);
nor U19018 (N_19018,N_12848,N_13402);
xnor U19019 (N_19019,N_14285,N_12952);
xnor U19020 (N_19020,N_11844,N_13231);
nand U19021 (N_19021,N_11122,N_11234);
and U19022 (N_19022,N_10957,N_10101);
or U19023 (N_19023,N_12976,N_12757);
xor U19024 (N_19024,N_13019,N_13283);
xnor U19025 (N_19025,N_14989,N_10742);
nand U19026 (N_19026,N_12221,N_14428);
xor U19027 (N_19027,N_12462,N_12063);
or U19028 (N_19028,N_11502,N_10746);
nor U19029 (N_19029,N_14817,N_11325);
nor U19030 (N_19030,N_11966,N_11289);
and U19031 (N_19031,N_11941,N_13512);
nor U19032 (N_19032,N_11967,N_14870);
and U19033 (N_19033,N_10549,N_13779);
nor U19034 (N_19034,N_10123,N_14243);
nor U19035 (N_19035,N_10372,N_11666);
or U19036 (N_19036,N_14773,N_14013);
xnor U19037 (N_19037,N_11585,N_12753);
or U19038 (N_19038,N_12345,N_12843);
or U19039 (N_19039,N_14471,N_12438);
or U19040 (N_19040,N_12758,N_12376);
and U19041 (N_19041,N_14238,N_12074);
or U19042 (N_19042,N_12994,N_13916);
nand U19043 (N_19043,N_13859,N_14159);
nand U19044 (N_19044,N_11454,N_10855);
nor U19045 (N_19045,N_13439,N_13263);
and U19046 (N_19046,N_13812,N_12860);
or U19047 (N_19047,N_10235,N_14147);
nor U19048 (N_19048,N_11807,N_14748);
nand U19049 (N_19049,N_12413,N_14884);
and U19050 (N_19050,N_10501,N_10770);
or U19051 (N_19051,N_10894,N_10526);
nor U19052 (N_19052,N_11846,N_14382);
nand U19053 (N_19053,N_14633,N_14253);
nor U19054 (N_19054,N_14153,N_14122);
nor U19055 (N_19055,N_10265,N_14489);
nand U19056 (N_19056,N_10171,N_10096);
nand U19057 (N_19057,N_10081,N_11656);
or U19058 (N_19058,N_12353,N_11906);
nand U19059 (N_19059,N_10682,N_10205);
and U19060 (N_19060,N_13236,N_12988);
nand U19061 (N_19061,N_10335,N_13495);
or U19062 (N_19062,N_12717,N_14479);
nor U19063 (N_19063,N_10349,N_12713);
nand U19064 (N_19064,N_12530,N_10383);
nand U19065 (N_19065,N_12522,N_13769);
and U19066 (N_19066,N_10254,N_11245);
and U19067 (N_19067,N_12808,N_10555);
and U19068 (N_19068,N_12424,N_11026);
nand U19069 (N_19069,N_13349,N_11824);
or U19070 (N_19070,N_11279,N_10632);
or U19071 (N_19071,N_13017,N_10213);
nor U19072 (N_19072,N_11860,N_13875);
and U19073 (N_19073,N_12713,N_12061);
and U19074 (N_19074,N_10149,N_11214);
nand U19075 (N_19075,N_11949,N_10435);
nand U19076 (N_19076,N_12233,N_12305);
and U19077 (N_19077,N_12176,N_12277);
nor U19078 (N_19078,N_14143,N_14748);
nor U19079 (N_19079,N_10914,N_11046);
and U19080 (N_19080,N_13799,N_10803);
or U19081 (N_19081,N_12822,N_13822);
and U19082 (N_19082,N_10405,N_14696);
and U19083 (N_19083,N_10484,N_13031);
nor U19084 (N_19084,N_14606,N_10610);
nand U19085 (N_19085,N_12101,N_11219);
nand U19086 (N_19086,N_10847,N_10213);
and U19087 (N_19087,N_12199,N_12083);
nor U19088 (N_19088,N_14571,N_13385);
nand U19089 (N_19089,N_12289,N_10056);
or U19090 (N_19090,N_11772,N_11483);
xnor U19091 (N_19091,N_12063,N_11810);
and U19092 (N_19092,N_14043,N_11751);
nand U19093 (N_19093,N_12047,N_12767);
or U19094 (N_19094,N_14246,N_13250);
nor U19095 (N_19095,N_10807,N_14374);
nor U19096 (N_19096,N_12196,N_13089);
nand U19097 (N_19097,N_14097,N_11813);
and U19098 (N_19098,N_11207,N_11635);
nor U19099 (N_19099,N_12118,N_11782);
xor U19100 (N_19100,N_14957,N_10706);
nand U19101 (N_19101,N_11595,N_13340);
xnor U19102 (N_19102,N_10292,N_11026);
xnor U19103 (N_19103,N_14783,N_11273);
and U19104 (N_19104,N_11071,N_13349);
nand U19105 (N_19105,N_14172,N_11671);
and U19106 (N_19106,N_11253,N_11265);
or U19107 (N_19107,N_11489,N_12045);
nor U19108 (N_19108,N_10157,N_14376);
or U19109 (N_19109,N_10973,N_14299);
or U19110 (N_19110,N_10219,N_13419);
or U19111 (N_19111,N_10956,N_13876);
and U19112 (N_19112,N_11130,N_13588);
nand U19113 (N_19113,N_10645,N_10449);
xor U19114 (N_19114,N_12600,N_10323);
or U19115 (N_19115,N_14540,N_12182);
and U19116 (N_19116,N_13968,N_13292);
nand U19117 (N_19117,N_12013,N_10595);
or U19118 (N_19118,N_12511,N_11333);
or U19119 (N_19119,N_14369,N_11635);
nand U19120 (N_19120,N_12012,N_13393);
or U19121 (N_19121,N_10842,N_12199);
or U19122 (N_19122,N_10690,N_14755);
nand U19123 (N_19123,N_14452,N_10327);
or U19124 (N_19124,N_10212,N_12043);
xnor U19125 (N_19125,N_14219,N_14865);
nand U19126 (N_19126,N_14154,N_12757);
nand U19127 (N_19127,N_11120,N_10732);
nand U19128 (N_19128,N_14444,N_13053);
nor U19129 (N_19129,N_12231,N_10889);
or U19130 (N_19130,N_12285,N_12540);
or U19131 (N_19131,N_12548,N_11700);
and U19132 (N_19132,N_10304,N_11989);
or U19133 (N_19133,N_10743,N_12128);
nor U19134 (N_19134,N_10902,N_14310);
nand U19135 (N_19135,N_11657,N_12874);
or U19136 (N_19136,N_14712,N_13076);
xnor U19137 (N_19137,N_12255,N_12323);
nand U19138 (N_19138,N_12224,N_14742);
or U19139 (N_19139,N_13016,N_12441);
nor U19140 (N_19140,N_11389,N_14754);
nor U19141 (N_19141,N_12805,N_10156);
or U19142 (N_19142,N_13196,N_14291);
nor U19143 (N_19143,N_12156,N_12822);
or U19144 (N_19144,N_13424,N_13151);
nand U19145 (N_19145,N_10842,N_13895);
nor U19146 (N_19146,N_11309,N_10228);
nor U19147 (N_19147,N_11372,N_11113);
or U19148 (N_19148,N_11763,N_13584);
nand U19149 (N_19149,N_12912,N_12603);
and U19150 (N_19150,N_13521,N_12154);
nand U19151 (N_19151,N_14784,N_10961);
and U19152 (N_19152,N_13711,N_13016);
xnor U19153 (N_19153,N_14251,N_13087);
nor U19154 (N_19154,N_13462,N_14434);
or U19155 (N_19155,N_10223,N_11647);
nand U19156 (N_19156,N_12579,N_14397);
and U19157 (N_19157,N_12888,N_10546);
or U19158 (N_19158,N_10736,N_11289);
and U19159 (N_19159,N_13119,N_10524);
nand U19160 (N_19160,N_10947,N_11375);
nand U19161 (N_19161,N_13691,N_14401);
xor U19162 (N_19162,N_13126,N_12536);
nor U19163 (N_19163,N_13628,N_10725);
nor U19164 (N_19164,N_14490,N_12712);
nand U19165 (N_19165,N_11372,N_14745);
nand U19166 (N_19166,N_10181,N_10757);
and U19167 (N_19167,N_10206,N_14176);
and U19168 (N_19168,N_10699,N_12683);
or U19169 (N_19169,N_11178,N_10773);
nor U19170 (N_19170,N_13179,N_13382);
nand U19171 (N_19171,N_12454,N_10263);
and U19172 (N_19172,N_12195,N_14149);
nor U19173 (N_19173,N_11498,N_12743);
nand U19174 (N_19174,N_14392,N_14375);
and U19175 (N_19175,N_10226,N_14526);
and U19176 (N_19176,N_14744,N_10251);
and U19177 (N_19177,N_10378,N_12354);
nor U19178 (N_19178,N_10889,N_13810);
nand U19179 (N_19179,N_12406,N_14454);
and U19180 (N_19180,N_11206,N_13139);
nor U19181 (N_19181,N_14434,N_13926);
or U19182 (N_19182,N_10784,N_14823);
nor U19183 (N_19183,N_11007,N_12402);
or U19184 (N_19184,N_13610,N_13827);
or U19185 (N_19185,N_11435,N_11531);
nor U19186 (N_19186,N_14809,N_10115);
nor U19187 (N_19187,N_11184,N_11681);
nand U19188 (N_19188,N_12121,N_14425);
or U19189 (N_19189,N_14657,N_10109);
nand U19190 (N_19190,N_14749,N_13769);
nor U19191 (N_19191,N_12045,N_13189);
or U19192 (N_19192,N_12123,N_14927);
or U19193 (N_19193,N_14540,N_11845);
nor U19194 (N_19194,N_13656,N_13199);
nand U19195 (N_19195,N_11606,N_10336);
or U19196 (N_19196,N_14941,N_13702);
nor U19197 (N_19197,N_14699,N_12520);
or U19198 (N_19198,N_13747,N_11845);
xnor U19199 (N_19199,N_12591,N_10634);
and U19200 (N_19200,N_14270,N_12986);
and U19201 (N_19201,N_10246,N_12591);
or U19202 (N_19202,N_10772,N_11472);
or U19203 (N_19203,N_10153,N_13084);
xnor U19204 (N_19204,N_12237,N_11138);
xor U19205 (N_19205,N_11976,N_11901);
or U19206 (N_19206,N_11025,N_11331);
nand U19207 (N_19207,N_10560,N_10014);
nor U19208 (N_19208,N_11175,N_13161);
and U19209 (N_19209,N_10062,N_13618);
xnor U19210 (N_19210,N_14904,N_11571);
or U19211 (N_19211,N_14025,N_12925);
and U19212 (N_19212,N_12608,N_12627);
xnor U19213 (N_19213,N_10241,N_12995);
nor U19214 (N_19214,N_14779,N_10089);
nand U19215 (N_19215,N_14674,N_10936);
nand U19216 (N_19216,N_10228,N_12805);
and U19217 (N_19217,N_11371,N_10826);
or U19218 (N_19218,N_10847,N_13053);
nor U19219 (N_19219,N_13538,N_14034);
nor U19220 (N_19220,N_11164,N_12957);
or U19221 (N_19221,N_11809,N_12791);
nor U19222 (N_19222,N_14451,N_14630);
and U19223 (N_19223,N_13220,N_12453);
nor U19224 (N_19224,N_12833,N_11218);
nor U19225 (N_19225,N_14436,N_14710);
and U19226 (N_19226,N_10822,N_10313);
nand U19227 (N_19227,N_12384,N_12125);
xnor U19228 (N_19228,N_14696,N_13464);
or U19229 (N_19229,N_10609,N_10038);
or U19230 (N_19230,N_14376,N_10463);
nor U19231 (N_19231,N_11983,N_10326);
and U19232 (N_19232,N_11750,N_12616);
and U19233 (N_19233,N_11850,N_14609);
or U19234 (N_19234,N_10121,N_14776);
and U19235 (N_19235,N_13888,N_14858);
nor U19236 (N_19236,N_10560,N_13556);
or U19237 (N_19237,N_12124,N_14738);
nor U19238 (N_19238,N_13988,N_13857);
and U19239 (N_19239,N_12815,N_12347);
or U19240 (N_19240,N_10933,N_12975);
or U19241 (N_19241,N_14846,N_13738);
and U19242 (N_19242,N_12342,N_10920);
or U19243 (N_19243,N_14505,N_14336);
nand U19244 (N_19244,N_10516,N_10831);
or U19245 (N_19245,N_11943,N_10651);
nand U19246 (N_19246,N_12700,N_11337);
xor U19247 (N_19247,N_13852,N_12189);
and U19248 (N_19248,N_10304,N_12831);
and U19249 (N_19249,N_12081,N_14767);
or U19250 (N_19250,N_13659,N_13624);
or U19251 (N_19251,N_11377,N_14333);
or U19252 (N_19252,N_13779,N_14770);
xor U19253 (N_19253,N_12344,N_10476);
nor U19254 (N_19254,N_14497,N_13985);
and U19255 (N_19255,N_10635,N_11644);
and U19256 (N_19256,N_14803,N_12818);
xnor U19257 (N_19257,N_11657,N_10523);
or U19258 (N_19258,N_12239,N_10860);
and U19259 (N_19259,N_13540,N_14627);
nor U19260 (N_19260,N_11588,N_13370);
or U19261 (N_19261,N_11868,N_11892);
nand U19262 (N_19262,N_13357,N_13255);
xnor U19263 (N_19263,N_13594,N_12692);
or U19264 (N_19264,N_14942,N_11165);
nor U19265 (N_19265,N_14997,N_11820);
nor U19266 (N_19266,N_14403,N_14883);
or U19267 (N_19267,N_14446,N_10105);
nand U19268 (N_19268,N_13009,N_13142);
and U19269 (N_19269,N_11446,N_10005);
nand U19270 (N_19270,N_14092,N_13769);
xnor U19271 (N_19271,N_11987,N_14781);
xnor U19272 (N_19272,N_14614,N_13917);
and U19273 (N_19273,N_13071,N_13369);
nor U19274 (N_19274,N_14403,N_11028);
or U19275 (N_19275,N_11411,N_14962);
nor U19276 (N_19276,N_10028,N_10045);
and U19277 (N_19277,N_14911,N_10200);
and U19278 (N_19278,N_14461,N_13702);
nand U19279 (N_19279,N_10410,N_14682);
or U19280 (N_19280,N_14582,N_12995);
nor U19281 (N_19281,N_10377,N_10481);
nor U19282 (N_19282,N_10889,N_10096);
and U19283 (N_19283,N_14181,N_11821);
or U19284 (N_19284,N_10012,N_11271);
or U19285 (N_19285,N_14015,N_10014);
or U19286 (N_19286,N_10132,N_14021);
and U19287 (N_19287,N_12553,N_12095);
and U19288 (N_19288,N_12414,N_14439);
nor U19289 (N_19289,N_11561,N_12533);
and U19290 (N_19290,N_10681,N_10017);
nor U19291 (N_19291,N_10506,N_13412);
and U19292 (N_19292,N_13175,N_10564);
or U19293 (N_19293,N_14532,N_12239);
nor U19294 (N_19294,N_14983,N_13310);
and U19295 (N_19295,N_10713,N_12481);
nand U19296 (N_19296,N_10834,N_12119);
nor U19297 (N_19297,N_12175,N_12340);
or U19298 (N_19298,N_12190,N_10496);
nor U19299 (N_19299,N_14777,N_13055);
or U19300 (N_19300,N_13913,N_14312);
or U19301 (N_19301,N_14112,N_12187);
nand U19302 (N_19302,N_12792,N_13078);
or U19303 (N_19303,N_10125,N_10912);
nand U19304 (N_19304,N_13883,N_13380);
xor U19305 (N_19305,N_13774,N_11572);
nor U19306 (N_19306,N_11808,N_14778);
nor U19307 (N_19307,N_11098,N_13765);
nand U19308 (N_19308,N_11510,N_13949);
xnor U19309 (N_19309,N_11210,N_10217);
nor U19310 (N_19310,N_12619,N_14910);
xor U19311 (N_19311,N_14833,N_13382);
and U19312 (N_19312,N_13435,N_14801);
nor U19313 (N_19313,N_14884,N_14809);
and U19314 (N_19314,N_12927,N_12250);
nand U19315 (N_19315,N_14821,N_12468);
and U19316 (N_19316,N_12269,N_10301);
nor U19317 (N_19317,N_10536,N_10565);
xor U19318 (N_19318,N_10183,N_14914);
nand U19319 (N_19319,N_11115,N_11787);
nor U19320 (N_19320,N_13846,N_12248);
or U19321 (N_19321,N_12352,N_13610);
nor U19322 (N_19322,N_10164,N_10537);
nand U19323 (N_19323,N_14901,N_11285);
or U19324 (N_19324,N_11307,N_12897);
nand U19325 (N_19325,N_13545,N_11269);
and U19326 (N_19326,N_10091,N_13245);
nand U19327 (N_19327,N_13614,N_13060);
nor U19328 (N_19328,N_12050,N_10220);
or U19329 (N_19329,N_14938,N_13174);
and U19330 (N_19330,N_13058,N_12395);
or U19331 (N_19331,N_13027,N_14825);
nor U19332 (N_19332,N_14934,N_13618);
or U19333 (N_19333,N_13765,N_11161);
nor U19334 (N_19334,N_11963,N_10104);
and U19335 (N_19335,N_13004,N_10702);
nand U19336 (N_19336,N_14970,N_13432);
and U19337 (N_19337,N_13146,N_14017);
nor U19338 (N_19338,N_14077,N_10515);
nand U19339 (N_19339,N_12346,N_11415);
nor U19340 (N_19340,N_12132,N_10832);
and U19341 (N_19341,N_12029,N_10940);
xor U19342 (N_19342,N_14138,N_11039);
nand U19343 (N_19343,N_14519,N_11266);
nand U19344 (N_19344,N_11938,N_12089);
or U19345 (N_19345,N_14835,N_12359);
and U19346 (N_19346,N_10501,N_14093);
and U19347 (N_19347,N_11482,N_10599);
or U19348 (N_19348,N_12828,N_12706);
nand U19349 (N_19349,N_11259,N_11457);
or U19350 (N_19350,N_14156,N_13555);
or U19351 (N_19351,N_14121,N_13453);
nand U19352 (N_19352,N_11315,N_12692);
nand U19353 (N_19353,N_13762,N_12986);
or U19354 (N_19354,N_11869,N_10869);
nand U19355 (N_19355,N_14966,N_13365);
nand U19356 (N_19356,N_11413,N_13428);
nand U19357 (N_19357,N_11655,N_12998);
and U19358 (N_19358,N_13655,N_12130);
nor U19359 (N_19359,N_13419,N_11806);
or U19360 (N_19360,N_12929,N_11998);
nand U19361 (N_19361,N_14327,N_10974);
nor U19362 (N_19362,N_13100,N_12620);
and U19363 (N_19363,N_14309,N_11189);
and U19364 (N_19364,N_12669,N_12691);
and U19365 (N_19365,N_14976,N_11997);
and U19366 (N_19366,N_11833,N_14541);
and U19367 (N_19367,N_14997,N_13089);
nand U19368 (N_19368,N_11279,N_12554);
and U19369 (N_19369,N_14120,N_11025);
xnor U19370 (N_19370,N_14528,N_13529);
or U19371 (N_19371,N_11088,N_14255);
and U19372 (N_19372,N_14127,N_12148);
and U19373 (N_19373,N_10742,N_10700);
and U19374 (N_19374,N_14568,N_12068);
or U19375 (N_19375,N_12460,N_13470);
nand U19376 (N_19376,N_11122,N_11620);
nor U19377 (N_19377,N_14215,N_11618);
nor U19378 (N_19378,N_11106,N_12999);
nand U19379 (N_19379,N_10507,N_11743);
and U19380 (N_19380,N_13661,N_14759);
and U19381 (N_19381,N_11980,N_10635);
nor U19382 (N_19382,N_14811,N_13778);
nor U19383 (N_19383,N_12854,N_13066);
and U19384 (N_19384,N_14305,N_10744);
nand U19385 (N_19385,N_13953,N_13851);
or U19386 (N_19386,N_14194,N_14913);
nand U19387 (N_19387,N_11376,N_12920);
nor U19388 (N_19388,N_12656,N_12150);
nor U19389 (N_19389,N_10775,N_12239);
nor U19390 (N_19390,N_14723,N_10227);
nand U19391 (N_19391,N_14661,N_13981);
or U19392 (N_19392,N_12704,N_11617);
or U19393 (N_19393,N_10309,N_14406);
nand U19394 (N_19394,N_11012,N_13731);
nand U19395 (N_19395,N_13015,N_11764);
nor U19396 (N_19396,N_11227,N_13449);
nand U19397 (N_19397,N_11053,N_10647);
nor U19398 (N_19398,N_13733,N_12560);
nor U19399 (N_19399,N_11792,N_11381);
and U19400 (N_19400,N_12913,N_12604);
or U19401 (N_19401,N_14585,N_13001);
nor U19402 (N_19402,N_11512,N_11665);
nand U19403 (N_19403,N_14892,N_11987);
and U19404 (N_19404,N_13097,N_10543);
nor U19405 (N_19405,N_11372,N_14954);
nor U19406 (N_19406,N_10904,N_13782);
nor U19407 (N_19407,N_13026,N_14507);
nor U19408 (N_19408,N_13895,N_14941);
nand U19409 (N_19409,N_12326,N_11647);
and U19410 (N_19410,N_14346,N_12229);
nand U19411 (N_19411,N_12417,N_14051);
or U19412 (N_19412,N_12281,N_11899);
nor U19413 (N_19413,N_13200,N_13821);
or U19414 (N_19414,N_11738,N_10521);
nand U19415 (N_19415,N_13903,N_10663);
nand U19416 (N_19416,N_11583,N_14305);
and U19417 (N_19417,N_11190,N_14245);
nand U19418 (N_19418,N_13395,N_12937);
and U19419 (N_19419,N_12317,N_14051);
or U19420 (N_19420,N_13483,N_12359);
and U19421 (N_19421,N_13971,N_14995);
nor U19422 (N_19422,N_11795,N_14473);
nand U19423 (N_19423,N_10598,N_13629);
nand U19424 (N_19424,N_14986,N_11244);
xor U19425 (N_19425,N_10248,N_14668);
nor U19426 (N_19426,N_12604,N_10271);
and U19427 (N_19427,N_10418,N_12900);
or U19428 (N_19428,N_14213,N_13730);
nor U19429 (N_19429,N_13036,N_11578);
xor U19430 (N_19430,N_13645,N_13791);
or U19431 (N_19431,N_12757,N_13943);
nor U19432 (N_19432,N_13726,N_14198);
and U19433 (N_19433,N_12780,N_11387);
nand U19434 (N_19434,N_13813,N_13815);
and U19435 (N_19435,N_12603,N_12974);
nor U19436 (N_19436,N_12055,N_10062);
nor U19437 (N_19437,N_14255,N_11324);
and U19438 (N_19438,N_14922,N_10215);
nand U19439 (N_19439,N_10192,N_12220);
nor U19440 (N_19440,N_10539,N_10212);
nand U19441 (N_19441,N_12906,N_11836);
nor U19442 (N_19442,N_12986,N_10986);
nor U19443 (N_19443,N_14347,N_14295);
and U19444 (N_19444,N_10405,N_10892);
and U19445 (N_19445,N_11672,N_12313);
nand U19446 (N_19446,N_12727,N_12097);
or U19447 (N_19447,N_10917,N_11513);
or U19448 (N_19448,N_14451,N_12803);
nand U19449 (N_19449,N_12460,N_11003);
xor U19450 (N_19450,N_14868,N_13042);
nor U19451 (N_19451,N_14886,N_13058);
xor U19452 (N_19452,N_13054,N_12572);
and U19453 (N_19453,N_10000,N_11665);
or U19454 (N_19454,N_13726,N_10606);
or U19455 (N_19455,N_10284,N_12018);
or U19456 (N_19456,N_13753,N_10015);
and U19457 (N_19457,N_12868,N_12731);
or U19458 (N_19458,N_13862,N_12366);
or U19459 (N_19459,N_14910,N_13106);
xor U19460 (N_19460,N_11945,N_10753);
or U19461 (N_19461,N_11665,N_12568);
or U19462 (N_19462,N_12941,N_11237);
nor U19463 (N_19463,N_11749,N_10548);
nand U19464 (N_19464,N_14542,N_13472);
nor U19465 (N_19465,N_12578,N_11190);
nand U19466 (N_19466,N_12909,N_12363);
nor U19467 (N_19467,N_12575,N_13927);
nor U19468 (N_19468,N_11304,N_12421);
and U19469 (N_19469,N_12860,N_10064);
or U19470 (N_19470,N_10784,N_10779);
or U19471 (N_19471,N_14721,N_12195);
or U19472 (N_19472,N_14324,N_10015);
nand U19473 (N_19473,N_14156,N_13129);
nor U19474 (N_19474,N_10675,N_14366);
or U19475 (N_19475,N_12025,N_10143);
nand U19476 (N_19476,N_11146,N_12272);
or U19477 (N_19477,N_12709,N_14927);
nor U19478 (N_19478,N_12952,N_11427);
or U19479 (N_19479,N_13753,N_13951);
and U19480 (N_19480,N_12805,N_14639);
nand U19481 (N_19481,N_12893,N_11316);
xor U19482 (N_19482,N_10484,N_14537);
nand U19483 (N_19483,N_13756,N_11038);
xnor U19484 (N_19484,N_11707,N_12282);
and U19485 (N_19485,N_13866,N_11498);
nor U19486 (N_19486,N_14590,N_13181);
or U19487 (N_19487,N_13954,N_12854);
or U19488 (N_19488,N_13275,N_11771);
nand U19489 (N_19489,N_13457,N_12122);
xnor U19490 (N_19490,N_13118,N_10948);
nand U19491 (N_19491,N_13976,N_14717);
nor U19492 (N_19492,N_14310,N_14856);
or U19493 (N_19493,N_14151,N_14159);
and U19494 (N_19494,N_13794,N_14863);
nand U19495 (N_19495,N_13620,N_10350);
nand U19496 (N_19496,N_14577,N_12266);
nor U19497 (N_19497,N_10277,N_11545);
nand U19498 (N_19498,N_11864,N_14312);
and U19499 (N_19499,N_10835,N_12359);
and U19500 (N_19500,N_14357,N_13112);
nand U19501 (N_19501,N_11833,N_14589);
xor U19502 (N_19502,N_14318,N_12563);
nand U19503 (N_19503,N_11097,N_14726);
and U19504 (N_19504,N_14155,N_11550);
and U19505 (N_19505,N_11575,N_10212);
nand U19506 (N_19506,N_11734,N_10836);
nor U19507 (N_19507,N_11610,N_13155);
or U19508 (N_19508,N_13889,N_14958);
xor U19509 (N_19509,N_10207,N_10627);
nor U19510 (N_19510,N_12382,N_10013);
nand U19511 (N_19511,N_12006,N_11988);
or U19512 (N_19512,N_13084,N_13364);
nor U19513 (N_19513,N_10353,N_13458);
and U19514 (N_19514,N_12391,N_10377);
nand U19515 (N_19515,N_12713,N_11733);
nor U19516 (N_19516,N_14178,N_12984);
nand U19517 (N_19517,N_13999,N_12149);
nor U19518 (N_19518,N_12478,N_11946);
nand U19519 (N_19519,N_10864,N_10564);
or U19520 (N_19520,N_11116,N_10844);
and U19521 (N_19521,N_13871,N_13811);
xor U19522 (N_19522,N_10992,N_14851);
and U19523 (N_19523,N_14848,N_10724);
nor U19524 (N_19524,N_11117,N_10591);
xnor U19525 (N_19525,N_14047,N_10543);
xnor U19526 (N_19526,N_14403,N_13463);
or U19527 (N_19527,N_14546,N_13421);
or U19528 (N_19528,N_12570,N_11205);
or U19529 (N_19529,N_14303,N_12849);
or U19530 (N_19530,N_14535,N_10319);
xnor U19531 (N_19531,N_10582,N_12801);
or U19532 (N_19532,N_13157,N_11308);
xnor U19533 (N_19533,N_12137,N_11100);
nor U19534 (N_19534,N_14296,N_11566);
and U19535 (N_19535,N_13093,N_13620);
nor U19536 (N_19536,N_10606,N_12786);
nand U19537 (N_19537,N_10804,N_11271);
xor U19538 (N_19538,N_11864,N_11470);
nand U19539 (N_19539,N_11159,N_12908);
nor U19540 (N_19540,N_11684,N_12039);
or U19541 (N_19541,N_12792,N_10838);
nor U19542 (N_19542,N_12373,N_13876);
or U19543 (N_19543,N_12344,N_10465);
nor U19544 (N_19544,N_12859,N_12482);
nor U19545 (N_19545,N_14095,N_11855);
nand U19546 (N_19546,N_14023,N_13983);
and U19547 (N_19547,N_10211,N_12909);
nor U19548 (N_19548,N_10260,N_10663);
nand U19549 (N_19549,N_12417,N_13787);
xor U19550 (N_19550,N_12806,N_10502);
nand U19551 (N_19551,N_13818,N_11014);
or U19552 (N_19552,N_14041,N_12385);
xor U19553 (N_19553,N_12156,N_14866);
or U19554 (N_19554,N_11391,N_14240);
and U19555 (N_19555,N_13599,N_14253);
and U19556 (N_19556,N_12816,N_11450);
and U19557 (N_19557,N_11005,N_14698);
and U19558 (N_19558,N_12214,N_12198);
nor U19559 (N_19559,N_11608,N_11378);
or U19560 (N_19560,N_13958,N_12208);
nand U19561 (N_19561,N_13717,N_13646);
or U19562 (N_19562,N_13102,N_14648);
xnor U19563 (N_19563,N_13904,N_12367);
and U19564 (N_19564,N_13796,N_12882);
or U19565 (N_19565,N_13937,N_12996);
xor U19566 (N_19566,N_13485,N_11932);
nor U19567 (N_19567,N_12039,N_12492);
or U19568 (N_19568,N_13460,N_14679);
and U19569 (N_19569,N_11663,N_10909);
nor U19570 (N_19570,N_13196,N_14692);
nor U19571 (N_19571,N_10938,N_12019);
nor U19572 (N_19572,N_11246,N_10560);
and U19573 (N_19573,N_14313,N_11782);
xnor U19574 (N_19574,N_13128,N_14022);
nand U19575 (N_19575,N_13005,N_13992);
xor U19576 (N_19576,N_10741,N_10219);
nor U19577 (N_19577,N_12372,N_13844);
nand U19578 (N_19578,N_11482,N_10057);
nor U19579 (N_19579,N_13092,N_14767);
or U19580 (N_19580,N_12853,N_14045);
nand U19581 (N_19581,N_14691,N_14244);
and U19582 (N_19582,N_12587,N_10679);
nor U19583 (N_19583,N_11022,N_10327);
nand U19584 (N_19584,N_11171,N_14043);
xor U19585 (N_19585,N_14688,N_12125);
nor U19586 (N_19586,N_14593,N_12571);
nor U19587 (N_19587,N_10472,N_10812);
or U19588 (N_19588,N_10923,N_11638);
or U19589 (N_19589,N_11519,N_14435);
and U19590 (N_19590,N_13693,N_13205);
and U19591 (N_19591,N_14989,N_11630);
nand U19592 (N_19592,N_14027,N_14234);
nand U19593 (N_19593,N_14108,N_12476);
nor U19594 (N_19594,N_11605,N_12052);
nor U19595 (N_19595,N_12354,N_12340);
xor U19596 (N_19596,N_13230,N_12100);
nor U19597 (N_19597,N_14695,N_14381);
nand U19598 (N_19598,N_14532,N_14688);
nand U19599 (N_19599,N_11243,N_14688);
nor U19600 (N_19600,N_12788,N_13550);
and U19601 (N_19601,N_10423,N_11931);
nor U19602 (N_19602,N_11767,N_12222);
nand U19603 (N_19603,N_10000,N_12315);
and U19604 (N_19604,N_11741,N_10070);
nor U19605 (N_19605,N_10506,N_11706);
and U19606 (N_19606,N_13750,N_13248);
nor U19607 (N_19607,N_14918,N_12912);
nor U19608 (N_19608,N_10656,N_12221);
nor U19609 (N_19609,N_14925,N_11404);
or U19610 (N_19610,N_14628,N_12875);
nand U19611 (N_19611,N_13286,N_14383);
nand U19612 (N_19612,N_12420,N_11673);
nor U19613 (N_19613,N_13324,N_13742);
or U19614 (N_19614,N_11796,N_13174);
and U19615 (N_19615,N_11982,N_14369);
nor U19616 (N_19616,N_14089,N_11445);
and U19617 (N_19617,N_12649,N_12908);
xor U19618 (N_19618,N_12675,N_14951);
xnor U19619 (N_19619,N_10441,N_13222);
nor U19620 (N_19620,N_10587,N_14465);
nand U19621 (N_19621,N_14535,N_14000);
and U19622 (N_19622,N_14673,N_10124);
and U19623 (N_19623,N_10868,N_11851);
and U19624 (N_19624,N_13956,N_14687);
xor U19625 (N_19625,N_13845,N_13958);
and U19626 (N_19626,N_10356,N_13998);
and U19627 (N_19627,N_11956,N_11845);
xnor U19628 (N_19628,N_10242,N_14838);
and U19629 (N_19629,N_11721,N_14644);
and U19630 (N_19630,N_12086,N_11980);
nand U19631 (N_19631,N_10815,N_12236);
xor U19632 (N_19632,N_11005,N_12502);
or U19633 (N_19633,N_11430,N_10463);
nor U19634 (N_19634,N_12096,N_10078);
or U19635 (N_19635,N_14904,N_11976);
nor U19636 (N_19636,N_10661,N_14572);
and U19637 (N_19637,N_10714,N_11062);
or U19638 (N_19638,N_11500,N_12779);
and U19639 (N_19639,N_13748,N_12956);
nor U19640 (N_19640,N_12995,N_10247);
nand U19641 (N_19641,N_11123,N_11158);
nand U19642 (N_19642,N_12518,N_14933);
and U19643 (N_19643,N_14513,N_13810);
nand U19644 (N_19644,N_14517,N_14934);
nand U19645 (N_19645,N_11594,N_14336);
xor U19646 (N_19646,N_12617,N_11450);
xor U19647 (N_19647,N_13081,N_14863);
nand U19648 (N_19648,N_14937,N_11733);
nor U19649 (N_19649,N_12203,N_13059);
nor U19650 (N_19650,N_11014,N_11309);
or U19651 (N_19651,N_14381,N_13248);
nand U19652 (N_19652,N_10888,N_13975);
nor U19653 (N_19653,N_11676,N_12536);
and U19654 (N_19654,N_12960,N_12284);
or U19655 (N_19655,N_10109,N_11722);
xor U19656 (N_19656,N_12472,N_14597);
and U19657 (N_19657,N_11600,N_10475);
and U19658 (N_19658,N_12854,N_10527);
nand U19659 (N_19659,N_13387,N_14470);
and U19660 (N_19660,N_10686,N_10857);
nor U19661 (N_19661,N_10001,N_13058);
nand U19662 (N_19662,N_12339,N_14016);
and U19663 (N_19663,N_14726,N_12806);
xor U19664 (N_19664,N_14546,N_13858);
nor U19665 (N_19665,N_14446,N_13413);
nand U19666 (N_19666,N_14606,N_12999);
nand U19667 (N_19667,N_11835,N_12920);
and U19668 (N_19668,N_10488,N_13171);
nand U19669 (N_19669,N_11136,N_10632);
and U19670 (N_19670,N_13085,N_12435);
or U19671 (N_19671,N_11602,N_10192);
or U19672 (N_19672,N_13580,N_14457);
nand U19673 (N_19673,N_12685,N_14169);
and U19674 (N_19674,N_11480,N_10832);
xnor U19675 (N_19675,N_11915,N_13535);
nand U19676 (N_19676,N_12385,N_13268);
and U19677 (N_19677,N_10780,N_12069);
or U19678 (N_19678,N_12779,N_13237);
or U19679 (N_19679,N_10581,N_10041);
nand U19680 (N_19680,N_13086,N_14201);
and U19681 (N_19681,N_14336,N_14615);
or U19682 (N_19682,N_14098,N_10427);
nor U19683 (N_19683,N_14961,N_11730);
and U19684 (N_19684,N_13441,N_12339);
nand U19685 (N_19685,N_13141,N_11772);
or U19686 (N_19686,N_10338,N_14838);
and U19687 (N_19687,N_11956,N_11121);
xor U19688 (N_19688,N_14151,N_11102);
xnor U19689 (N_19689,N_14555,N_10290);
nand U19690 (N_19690,N_13020,N_13237);
and U19691 (N_19691,N_13987,N_12465);
or U19692 (N_19692,N_10976,N_13543);
and U19693 (N_19693,N_13000,N_14660);
or U19694 (N_19694,N_13490,N_11965);
and U19695 (N_19695,N_13917,N_11208);
and U19696 (N_19696,N_12392,N_12514);
xor U19697 (N_19697,N_11673,N_11860);
or U19698 (N_19698,N_13681,N_12681);
and U19699 (N_19699,N_10298,N_14767);
nor U19700 (N_19700,N_11177,N_14057);
and U19701 (N_19701,N_13177,N_13248);
nor U19702 (N_19702,N_10362,N_10354);
and U19703 (N_19703,N_14838,N_10207);
nand U19704 (N_19704,N_11084,N_11304);
and U19705 (N_19705,N_14131,N_11578);
or U19706 (N_19706,N_10057,N_12841);
nand U19707 (N_19707,N_12215,N_13452);
xor U19708 (N_19708,N_11622,N_11624);
nand U19709 (N_19709,N_12253,N_10072);
nor U19710 (N_19710,N_13960,N_10735);
and U19711 (N_19711,N_14993,N_11634);
nor U19712 (N_19712,N_10985,N_14051);
or U19713 (N_19713,N_10787,N_13023);
nand U19714 (N_19714,N_11546,N_10341);
nor U19715 (N_19715,N_10058,N_12580);
nand U19716 (N_19716,N_14989,N_14106);
and U19717 (N_19717,N_11719,N_13518);
nor U19718 (N_19718,N_11865,N_11475);
or U19719 (N_19719,N_13461,N_14499);
or U19720 (N_19720,N_11825,N_13900);
nand U19721 (N_19721,N_14752,N_13261);
nor U19722 (N_19722,N_13487,N_10163);
nand U19723 (N_19723,N_13505,N_12563);
nand U19724 (N_19724,N_13937,N_13394);
and U19725 (N_19725,N_10856,N_13468);
or U19726 (N_19726,N_11661,N_13609);
and U19727 (N_19727,N_11674,N_10713);
nand U19728 (N_19728,N_11965,N_12763);
xor U19729 (N_19729,N_14815,N_11939);
nand U19730 (N_19730,N_14411,N_13534);
and U19731 (N_19731,N_14175,N_10581);
or U19732 (N_19732,N_14111,N_13195);
and U19733 (N_19733,N_11462,N_12033);
or U19734 (N_19734,N_12201,N_13174);
nor U19735 (N_19735,N_11558,N_13634);
and U19736 (N_19736,N_11413,N_10100);
or U19737 (N_19737,N_12355,N_10512);
or U19738 (N_19738,N_13969,N_12940);
nor U19739 (N_19739,N_13729,N_12503);
nand U19740 (N_19740,N_12425,N_11031);
or U19741 (N_19741,N_13260,N_11313);
nand U19742 (N_19742,N_14668,N_13901);
or U19743 (N_19743,N_10062,N_14443);
nand U19744 (N_19744,N_12082,N_10983);
nand U19745 (N_19745,N_13224,N_10849);
and U19746 (N_19746,N_11249,N_12736);
and U19747 (N_19747,N_12183,N_13133);
nor U19748 (N_19748,N_13787,N_12111);
xor U19749 (N_19749,N_14653,N_12574);
and U19750 (N_19750,N_10649,N_10811);
or U19751 (N_19751,N_12638,N_10595);
nor U19752 (N_19752,N_11771,N_11935);
nor U19753 (N_19753,N_14857,N_12210);
and U19754 (N_19754,N_12601,N_13185);
xnor U19755 (N_19755,N_12097,N_13547);
xor U19756 (N_19756,N_10486,N_11806);
nand U19757 (N_19757,N_14967,N_13707);
nor U19758 (N_19758,N_12900,N_13714);
nand U19759 (N_19759,N_12703,N_12543);
and U19760 (N_19760,N_11141,N_13769);
and U19761 (N_19761,N_13302,N_12693);
and U19762 (N_19762,N_12438,N_14237);
nand U19763 (N_19763,N_10531,N_10231);
and U19764 (N_19764,N_13610,N_10119);
or U19765 (N_19765,N_11458,N_13849);
nand U19766 (N_19766,N_14098,N_11975);
and U19767 (N_19767,N_14534,N_10931);
or U19768 (N_19768,N_12990,N_13751);
nor U19769 (N_19769,N_10244,N_11008);
or U19770 (N_19770,N_13234,N_11208);
and U19771 (N_19771,N_12181,N_10953);
or U19772 (N_19772,N_13880,N_12155);
or U19773 (N_19773,N_12253,N_11089);
or U19774 (N_19774,N_14527,N_12333);
xnor U19775 (N_19775,N_13213,N_10510);
nand U19776 (N_19776,N_10285,N_12602);
nor U19777 (N_19777,N_11676,N_12860);
and U19778 (N_19778,N_13322,N_13794);
nand U19779 (N_19779,N_11615,N_12505);
and U19780 (N_19780,N_10173,N_10664);
nand U19781 (N_19781,N_12898,N_12164);
nor U19782 (N_19782,N_14765,N_13843);
and U19783 (N_19783,N_13044,N_11215);
nor U19784 (N_19784,N_10657,N_10225);
nand U19785 (N_19785,N_12356,N_11576);
xnor U19786 (N_19786,N_11284,N_11369);
nor U19787 (N_19787,N_10572,N_12711);
or U19788 (N_19788,N_12197,N_14560);
nor U19789 (N_19789,N_11514,N_10873);
or U19790 (N_19790,N_11999,N_11533);
nor U19791 (N_19791,N_12982,N_10208);
or U19792 (N_19792,N_12662,N_11462);
and U19793 (N_19793,N_11199,N_13216);
nand U19794 (N_19794,N_11191,N_10419);
or U19795 (N_19795,N_12143,N_11106);
xnor U19796 (N_19796,N_11055,N_14825);
and U19797 (N_19797,N_11413,N_13896);
nor U19798 (N_19798,N_11762,N_12153);
and U19799 (N_19799,N_12740,N_10010);
nor U19800 (N_19800,N_14536,N_12943);
nand U19801 (N_19801,N_12772,N_12099);
nor U19802 (N_19802,N_10799,N_10778);
and U19803 (N_19803,N_13076,N_14418);
or U19804 (N_19804,N_13530,N_13907);
and U19805 (N_19805,N_14620,N_11042);
nor U19806 (N_19806,N_10236,N_11078);
xor U19807 (N_19807,N_12736,N_14954);
xnor U19808 (N_19808,N_12095,N_11410);
and U19809 (N_19809,N_11683,N_10141);
or U19810 (N_19810,N_14864,N_12895);
nand U19811 (N_19811,N_12810,N_13651);
nand U19812 (N_19812,N_12141,N_13286);
and U19813 (N_19813,N_11796,N_12826);
and U19814 (N_19814,N_10089,N_10555);
nand U19815 (N_19815,N_11858,N_10987);
or U19816 (N_19816,N_13646,N_12315);
nand U19817 (N_19817,N_14223,N_10381);
and U19818 (N_19818,N_14236,N_13023);
or U19819 (N_19819,N_12423,N_13310);
nor U19820 (N_19820,N_12210,N_13155);
nand U19821 (N_19821,N_11457,N_13039);
and U19822 (N_19822,N_13129,N_13358);
nand U19823 (N_19823,N_13135,N_13011);
nor U19824 (N_19824,N_10877,N_11283);
xnor U19825 (N_19825,N_10201,N_11692);
nor U19826 (N_19826,N_13927,N_11252);
or U19827 (N_19827,N_12490,N_10757);
or U19828 (N_19828,N_13047,N_12595);
nor U19829 (N_19829,N_12846,N_14014);
nor U19830 (N_19830,N_12868,N_13147);
and U19831 (N_19831,N_12660,N_14891);
or U19832 (N_19832,N_14979,N_10898);
and U19833 (N_19833,N_12505,N_12645);
or U19834 (N_19834,N_10674,N_13309);
nand U19835 (N_19835,N_14634,N_13880);
nand U19836 (N_19836,N_12350,N_10296);
or U19837 (N_19837,N_12990,N_14526);
nor U19838 (N_19838,N_11463,N_13576);
and U19839 (N_19839,N_13434,N_13148);
nor U19840 (N_19840,N_13591,N_13439);
nor U19841 (N_19841,N_14291,N_12668);
nand U19842 (N_19842,N_13179,N_14197);
nor U19843 (N_19843,N_11247,N_11011);
xor U19844 (N_19844,N_10717,N_10215);
nand U19845 (N_19845,N_11054,N_13012);
and U19846 (N_19846,N_13779,N_13715);
nand U19847 (N_19847,N_14853,N_11147);
xor U19848 (N_19848,N_13979,N_13169);
nor U19849 (N_19849,N_13316,N_12977);
and U19850 (N_19850,N_10829,N_13928);
xor U19851 (N_19851,N_12331,N_11401);
nand U19852 (N_19852,N_14486,N_13737);
nor U19853 (N_19853,N_12330,N_13092);
nand U19854 (N_19854,N_13154,N_14616);
nand U19855 (N_19855,N_14436,N_12781);
nor U19856 (N_19856,N_13186,N_13828);
nand U19857 (N_19857,N_12714,N_10425);
or U19858 (N_19858,N_12648,N_11686);
nor U19859 (N_19859,N_13873,N_14662);
and U19860 (N_19860,N_11390,N_13302);
or U19861 (N_19861,N_12764,N_13910);
and U19862 (N_19862,N_12950,N_12345);
nor U19863 (N_19863,N_10065,N_12990);
nor U19864 (N_19864,N_10548,N_12844);
nor U19865 (N_19865,N_10975,N_11874);
nor U19866 (N_19866,N_14680,N_10819);
and U19867 (N_19867,N_14335,N_11417);
nor U19868 (N_19868,N_11125,N_14012);
nor U19869 (N_19869,N_12935,N_14220);
and U19870 (N_19870,N_11880,N_10588);
and U19871 (N_19871,N_12487,N_11599);
or U19872 (N_19872,N_14433,N_11572);
nor U19873 (N_19873,N_11750,N_13055);
xor U19874 (N_19874,N_10205,N_11818);
or U19875 (N_19875,N_13354,N_10777);
nor U19876 (N_19876,N_14528,N_14453);
or U19877 (N_19877,N_11192,N_10029);
and U19878 (N_19878,N_12978,N_13870);
nor U19879 (N_19879,N_13908,N_11966);
and U19880 (N_19880,N_14682,N_11817);
or U19881 (N_19881,N_14115,N_10640);
xor U19882 (N_19882,N_14242,N_12572);
and U19883 (N_19883,N_11795,N_10507);
xnor U19884 (N_19884,N_11965,N_10567);
nand U19885 (N_19885,N_11858,N_10964);
nor U19886 (N_19886,N_11798,N_11474);
nand U19887 (N_19887,N_10074,N_13556);
or U19888 (N_19888,N_10826,N_10180);
nor U19889 (N_19889,N_10324,N_10868);
or U19890 (N_19890,N_13338,N_12926);
nand U19891 (N_19891,N_11870,N_10924);
nor U19892 (N_19892,N_14645,N_12743);
or U19893 (N_19893,N_14433,N_12562);
xnor U19894 (N_19894,N_10946,N_14597);
or U19895 (N_19895,N_14049,N_10855);
nor U19896 (N_19896,N_14082,N_14505);
nand U19897 (N_19897,N_10906,N_13633);
or U19898 (N_19898,N_10290,N_13733);
nor U19899 (N_19899,N_14739,N_10238);
nand U19900 (N_19900,N_11617,N_11353);
nand U19901 (N_19901,N_10918,N_14700);
and U19902 (N_19902,N_12692,N_10644);
nand U19903 (N_19903,N_11157,N_13571);
and U19904 (N_19904,N_14833,N_12634);
nand U19905 (N_19905,N_12575,N_14187);
or U19906 (N_19906,N_10332,N_10495);
nand U19907 (N_19907,N_12607,N_11100);
or U19908 (N_19908,N_11973,N_14323);
and U19909 (N_19909,N_14547,N_11663);
xnor U19910 (N_19910,N_14367,N_11429);
or U19911 (N_19911,N_14081,N_14273);
xnor U19912 (N_19912,N_14867,N_10155);
xnor U19913 (N_19913,N_10925,N_10943);
nor U19914 (N_19914,N_12728,N_14548);
and U19915 (N_19915,N_12000,N_10308);
xnor U19916 (N_19916,N_14476,N_12606);
and U19917 (N_19917,N_12783,N_10486);
nand U19918 (N_19918,N_11052,N_13633);
nand U19919 (N_19919,N_11381,N_11954);
and U19920 (N_19920,N_10079,N_13493);
nand U19921 (N_19921,N_14962,N_11227);
or U19922 (N_19922,N_13904,N_10827);
nand U19923 (N_19923,N_12994,N_14996);
or U19924 (N_19924,N_11881,N_12522);
and U19925 (N_19925,N_11235,N_14343);
or U19926 (N_19926,N_13891,N_10488);
and U19927 (N_19927,N_12245,N_14348);
or U19928 (N_19928,N_14114,N_12722);
nand U19929 (N_19929,N_14920,N_10772);
nand U19930 (N_19930,N_14161,N_13687);
or U19931 (N_19931,N_14384,N_14373);
nand U19932 (N_19932,N_13416,N_13076);
and U19933 (N_19933,N_11162,N_14277);
or U19934 (N_19934,N_12109,N_12387);
xor U19935 (N_19935,N_12935,N_12082);
or U19936 (N_19936,N_10948,N_14470);
xor U19937 (N_19937,N_12813,N_12432);
or U19938 (N_19938,N_12671,N_13720);
and U19939 (N_19939,N_10447,N_11415);
nand U19940 (N_19940,N_14386,N_13432);
or U19941 (N_19941,N_13716,N_12128);
xor U19942 (N_19942,N_13575,N_12617);
or U19943 (N_19943,N_11940,N_14010);
and U19944 (N_19944,N_10340,N_12236);
nor U19945 (N_19945,N_12047,N_12894);
nand U19946 (N_19946,N_12798,N_10707);
and U19947 (N_19947,N_11944,N_12998);
or U19948 (N_19948,N_12582,N_12779);
nor U19949 (N_19949,N_12511,N_13997);
nor U19950 (N_19950,N_14247,N_11040);
or U19951 (N_19951,N_11758,N_12624);
and U19952 (N_19952,N_10527,N_14248);
nand U19953 (N_19953,N_11984,N_10939);
or U19954 (N_19954,N_12889,N_13244);
or U19955 (N_19955,N_10225,N_11155);
and U19956 (N_19956,N_14988,N_11074);
nor U19957 (N_19957,N_10694,N_14866);
nor U19958 (N_19958,N_10319,N_14260);
nand U19959 (N_19959,N_14058,N_14220);
or U19960 (N_19960,N_13496,N_11641);
nand U19961 (N_19961,N_13747,N_14924);
nor U19962 (N_19962,N_10371,N_10798);
nor U19963 (N_19963,N_14069,N_11824);
nand U19964 (N_19964,N_10697,N_13634);
xnor U19965 (N_19965,N_11387,N_13707);
nor U19966 (N_19966,N_14087,N_11344);
and U19967 (N_19967,N_12345,N_14410);
and U19968 (N_19968,N_12086,N_12469);
nand U19969 (N_19969,N_14292,N_14149);
nor U19970 (N_19970,N_11064,N_11858);
nor U19971 (N_19971,N_12938,N_14771);
and U19972 (N_19972,N_13002,N_13136);
or U19973 (N_19973,N_12861,N_14544);
and U19974 (N_19974,N_14623,N_13668);
and U19975 (N_19975,N_11328,N_13803);
nor U19976 (N_19976,N_14858,N_13511);
nor U19977 (N_19977,N_12938,N_14413);
xnor U19978 (N_19978,N_11619,N_10276);
nor U19979 (N_19979,N_13351,N_11076);
or U19980 (N_19980,N_10108,N_11518);
or U19981 (N_19981,N_13116,N_11140);
or U19982 (N_19982,N_14568,N_11988);
and U19983 (N_19983,N_14383,N_12286);
nor U19984 (N_19984,N_14837,N_11709);
nand U19985 (N_19985,N_13259,N_12559);
or U19986 (N_19986,N_10550,N_14353);
and U19987 (N_19987,N_11736,N_13530);
and U19988 (N_19988,N_11879,N_11659);
xor U19989 (N_19989,N_14526,N_14178);
nor U19990 (N_19990,N_14494,N_13705);
nand U19991 (N_19991,N_10443,N_11149);
or U19992 (N_19992,N_12033,N_12861);
nor U19993 (N_19993,N_13266,N_12028);
nand U19994 (N_19994,N_11027,N_11636);
or U19995 (N_19995,N_13750,N_11940);
and U19996 (N_19996,N_13348,N_13283);
nor U19997 (N_19997,N_10415,N_11322);
nor U19998 (N_19998,N_14774,N_11980);
and U19999 (N_19999,N_12729,N_10320);
and U20000 (N_20000,N_19525,N_16795);
and U20001 (N_20001,N_17758,N_16553);
and U20002 (N_20002,N_18457,N_18585);
and U20003 (N_20003,N_16572,N_16903);
nor U20004 (N_20004,N_18070,N_19671);
and U20005 (N_20005,N_16707,N_18150);
and U20006 (N_20006,N_16416,N_16494);
or U20007 (N_20007,N_18277,N_16090);
nand U20008 (N_20008,N_18290,N_15973);
xnor U20009 (N_20009,N_19890,N_16874);
nand U20010 (N_20010,N_17721,N_18535);
nor U20011 (N_20011,N_17619,N_17208);
and U20012 (N_20012,N_17897,N_16060);
nor U20013 (N_20013,N_16922,N_19881);
or U20014 (N_20014,N_17079,N_16630);
nor U20015 (N_20015,N_18245,N_18677);
or U20016 (N_20016,N_19505,N_16597);
nand U20017 (N_20017,N_17724,N_19927);
xnor U20018 (N_20018,N_16515,N_15779);
nor U20019 (N_20019,N_18176,N_18092);
nor U20020 (N_20020,N_19483,N_17108);
nand U20021 (N_20021,N_19828,N_19771);
or U20022 (N_20022,N_17520,N_16972);
and U20023 (N_20023,N_17007,N_17463);
nand U20024 (N_20024,N_16743,N_18663);
nor U20025 (N_20025,N_18059,N_16947);
and U20026 (N_20026,N_18167,N_15769);
nor U20027 (N_20027,N_18917,N_16289);
or U20028 (N_20028,N_15496,N_17708);
nand U20029 (N_20029,N_19552,N_17992);
nor U20030 (N_20030,N_19443,N_16190);
nand U20031 (N_20031,N_18750,N_15088);
nand U20032 (N_20032,N_19855,N_18863);
nor U20033 (N_20033,N_15199,N_16722);
nand U20034 (N_20034,N_19725,N_18537);
nand U20035 (N_20035,N_16902,N_16253);
and U20036 (N_20036,N_16221,N_18922);
or U20037 (N_20037,N_18182,N_19328);
and U20038 (N_20038,N_18437,N_17266);
and U20039 (N_20039,N_17197,N_19979);
nand U20040 (N_20040,N_19698,N_18301);
or U20041 (N_20041,N_18713,N_18539);
xor U20042 (N_20042,N_19223,N_16774);
nand U20043 (N_20043,N_18055,N_16917);
nor U20044 (N_20044,N_15747,N_15342);
nor U20045 (N_20045,N_16987,N_18840);
nor U20046 (N_20046,N_19187,N_19666);
and U20047 (N_20047,N_16831,N_16561);
nor U20048 (N_20048,N_15123,N_16834);
and U20049 (N_20049,N_18430,N_19951);
nand U20050 (N_20050,N_16143,N_17174);
nand U20051 (N_20051,N_16620,N_15096);
nor U20052 (N_20052,N_18013,N_16661);
nor U20053 (N_20053,N_19083,N_18734);
and U20054 (N_20054,N_15378,N_16042);
nor U20055 (N_20055,N_18199,N_15809);
nor U20056 (N_20056,N_19165,N_16039);
nor U20057 (N_20057,N_18074,N_17468);
or U20058 (N_20058,N_15466,N_18387);
or U20059 (N_20059,N_17765,N_19735);
and U20060 (N_20060,N_19542,N_19240);
nor U20061 (N_20061,N_18031,N_16918);
and U20062 (N_20062,N_17451,N_19945);
nand U20063 (N_20063,N_15283,N_17435);
and U20064 (N_20064,N_16666,N_19730);
or U20065 (N_20065,N_15002,N_18755);
nand U20066 (N_20066,N_18044,N_17403);
nor U20067 (N_20067,N_19239,N_15299);
or U20068 (N_20068,N_19308,N_17027);
nand U20069 (N_20069,N_15167,N_18994);
nand U20070 (N_20070,N_19019,N_15840);
and U20071 (N_20071,N_18156,N_15945);
nand U20072 (N_20072,N_19999,N_17582);
nand U20073 (N_20073,N_19392,N_15879);
nor U20074 (N_20074,N_15639,N_17168);
nand U20075 (N_20075,N_18588,N_15946);
and U20076 (N_20076,N_15994,N_18964);
or U20077 (N_20077,N_17531,N_15422);
nor U20078 (N_20078,N_15417,N_19621);
xor U20079 (N_20079,N_17204,N_15230);
and U20080 (N_20080,N_19491,N_19895);
nor U20081 (N_20081,N_16593,N_18073);
or U20082 (N_20082,N_17034,N_16485);
nor U20083 (N_20083,N_15381,N_17206);
nand U20084 (N_20084,N_15741,N_17839);
or U20085 (N_20085,N_17049,N_15428);
nand U20086 (N_20086,N_15780,N_15653);
nand U20087 (N_20087,N_15412,N_18339);
nand U20088 (N_20088,N_18586,N_15312);
xnor U20089 (N_20089,N_16808,N_18417);
and U20090 (N_20090,N_15166,N_18705);
nand U20091 (N_20091,N_17710,N_17396);
nor U20092 (N_20092,N_16235,N_16077);
or U20093 (N_20093,N_19184,N_19042);
nand U20094 (N_20094,N_19113,N_18855);
xor U20095 (N_20095,N_19602,N_18421);
nand U20096 (N_20096,N_17474,N_16968);
and U20097 (N_20097,N_17021,N_15313);
nor U20098 (N_20098,N_15213,N_16985);
nor U20099 (N_20099,N_15992,N_17249);
nand U20100 (N_20100,N_16714,N_16479);
nand U20101 (N_20101,N_17057,N_19422);
nand U20102 (N_20102,N_17660,N_16365);
nor U20103 (N_20103,N_19195,N_18386);
nand U20104 (N_20104,N_17088,N_19252);
and U20105 (N_20105,N_15191,N_16841);
or U20106 (N_20106,N_16934,N_17472);
nand U20107 (N_20107,N_19623,N_19038);
and U20108 (N_20108,N_19901,N_18095);
nor U20109 (N_20109,N_17343,N_16640);
and U20110 (N_20110,N_15884,N_18498);
and U20111 (N_20111,N_18419,N_18121);
xor U20112 (N_20112,N_17106,N_19864);
nand U20113 (N_20113,N_15696,N_17551);
nand U20114 (N_20114,N_18340,N_19333);
or U20115 (N_20115,N_15642,N_18448);
xnor U20116 (N_20116,N_18595,N_17571);
nand U20117 (N_20117,N_19986,N_18489);
and U20118 (N_20118,N_15515,N_16877);
nor U20119 (N_20119,N_18774,N_18392);
nor U20120 (N_20120,N_17385,N_19589);
nand U20121 (N_20121,N_16789,N_19772);
nand U20122 (N_20122,N_17828,N_17956);
and U20123 (N_20123,N_19037,N_17037);
or U20124 (N_20124,N_16034,N_17688);
and U20125 (N_20125,N_19952,N_17332);
nor U20126 (N_20126,N_19587,N_17600);
and U20127 (N_20127,N_17980,N_19801);
nor U20128 (N_20128,N_17450,N_19792);
xor U20129 (N_20129,N_18507,N_18493);
nor U20130 (N_20130,N_16772,N_19391);
nor U20131 (N_20131,N_18341,N_18980);
and U20132 (N_20132,N_18376,N_16786);
nor U20133 (N_20133,N_17193,N_15162);
or U20134 (N_20134,N_17547,N_19992);
and U20135 (N_20135,N_16096,N_15113);
nand U20136 (N_20136,N_16465,N_19168);
and U20137 (N_20137,N_16558,N_17277);
xnor U20138 (N_20138,N_15277,N_15452);
nand U20139 (N_20139,N_19747,N_19169);
nor U20140 (N_20140,N_16638,N_15483);
nor U20141 (N_20141,N_16125,N_18008);
nor U20142 (N_20142,N_15661,N_18096);
and U20143 (N_20143,N_17466,N_18864);
or U20144 (N_20144,N_17996,N_18977);
nor U20145 (N_20145,N_15393,N_17667);
and U20146 (N_20146,N_16989,N_18307);
xor U20147 (N_20147,N_18600,N_16738);
or U20148 (N_20148,N_18924,N_17824);
nand U20149 (N_20149,N_19371,N_17043);
or U20150 (N_20150,N_17275,N_17261);
nand U20151 (N_20151,N_16621,N_15603);
nor U20152 (N_20152,N_15938,N_16905);
nand U20153 (N_20153,N_19406,N_16976);
or U20154 (N_20154,N_16956,N_17822);
nand U20155 (N_20155,N_15771,N_17560);
nand U20156 (N_20156,N_18270,N_17963);
or U20157 (N_20157,N_16375,N_19858);
or U20158 (N_20158,N_15812,N_16059);
and U20159 (N_20159,N_17669,N_17642);
nor U20160 (N_20160,N_16313,N_18715);
nand U20161 (N_20161,N_18434,N_16281);
and U20162 (N_20162,N_19216,N_15392);
or U20163 (N_20163,N_19290,N_15244);
nand U20164 (N_20164,N_18674,N_19840);
nor U20165 (N_20165,N_15154,N_16857);
and U20166 (N_20166,N_17484,N_17630);
nor U20167 (N_20167,N_17480,N_18813);
xnor U20168 (N_20168,N_18184,N_18284);
or U20169 (N_20169,N_15280,N_15703);
or U20170 (N_20170,N_17747,N_15666);
nand U20171 (N_20171,N_15681,N_17664);
xnor U20172 (N_20172,N_16236,N_18825);
or U20173 (N_20173,N_16290,N_15424);
or U20174 (N_20174,N_19578,N_19056);
nand U20175 (N_20175,N_17938,N_15649);
or U20176 (N_20176,N_16346,N_19141);
xnor U20177 (N_20177,N_18278,N_17243);
xnor U20178 (N_20178,N_16624,N_15332);
nor U20179 (N_20179,N_16560,N_17247);
xnor U20180 (N_20180,N_15896,N_16896);
and U20181 (N_20181,N_16071,N_18928);
or U20182 (N_20182,N_19315,N_15009);
nor U20183 (N_20183,N_15804,N_15545);
nor U20184 (N_20184,N_18797,N_18068);
xnor U20185 (N_20185,N_18984,N_17175);
xor U20186 (N_20186,N_15608,N_19346);
or U20187 (N_20187,N_15212,N_16673);
nor U20188 (N_20188,N_15658,N_15498);
nand U20189 (N_20189,N_19605,N_16439);
xor U20190 (N_20190,N_17904,N_15012);
nand U20191 (N_20191,N_15526,N_15011);
nand U20192 (N_20192,N_18685,N_15750);
or U20193 (N_20193,N_15908,N_15484);
and U20194 (N_20194,N_16982,N_17264);
nand U20195 (N_20195,N_19917,N_16833);
and U20196 (N_20196,N_16403,N_15617);
and U20197 (N_20197,N_15411,N_16813);
xnor U20198 (N_20198,N_18959,N_19975);
nor U20199 (N_20199,N_17920,N_16233);
or U20200 (N_20200,N_15019,N_16156);
or U20201 (N_20201,N_15182,N_15200);
nand U20202 (N_20202,N_15263,N_15523);
nor U20203 (N_20203,N_16599,N_17580);
and U20204 (N_20204,N_17890,N_15298);
nand U20205 (N_20205,N_16598,N_17025);
and U20206 (N_20206,N_19852,N_17993);
and U20207 (N_20207,N_19379,N_19762);
or U20208 (N_20208,N_19726,N_17879);
nor U20209 (N_20209,N_16908,N_17382);
nor U20210 (N_20210,N_17769,N_16242);
or U20211 (N_20211,N_17540,N_18873);
xnor U20212 (N_20212,N_18117,N_16514);
or U20213 (N_20213,N_16304,N_16248);
or U20214 (N_20214,N_19384,N_16733);
and U20215 (N_20215,N_19791,N_15098);
and U20216 (N_20216,N_17233,N_19980);
and U20217 (N_20217,N_15099,N_17255);
nor U20218 (N_20218,N_19495,N_19508);
nor U20219 (N_20219,N_16647,N_19631);
nand U20220 (N_20220,N_17722,N_16822);
xor U20221 (N_20221,N_18583,N_17810);
and U20222 (N_20222,N_19268,N_15258);
nand U20223 (N_20223,N_19287,N_17651);
and U20224 (N_20224,N_19850,N_16108);
or U20225 (N_20225,N_17803,N_19301);
nor U20226 (N_20226,N_18312,N_17320);
or U20227 (N_20227,N_19954,N_18528);
or U20228 (N_20228,N_18453,N_19147);
nor U20229 (N_20229,N_18272,N_19217);
nand U20230 (N_20230,N_18519,N_19142);
or U20231 (N_20231,N_19106,N_15729);
and U20232 (N_20232,N_17067,N_18433);
nand U20233 (N_20233,N_17786,N_19736);
or U20234 (N_20234,N_15748,N_19242);
and U20235 (N_20235,N_17072,N_19245);
xor U20236 (N_20236,N_17137,N_19423);
nor U20237 (N_20237,N_15815,N_19732);
nand U20238 (N_20238,N_16137,N_17607);
and U20239 (N_20239,N_19398,N_15756);
nand U20240 (N_20240,N_15989,N_16352);
nand U20241 (N_20241,N_15219,N_16488);
nand U20242 (N_20242,N_18206,N_19533);
nor U20243 (N_20243,N_18534,N_16435);
xor U20244 (N_20244,N_15129,N_19462);
xor U20245 (N_20245,N_15024,N_16818);
or U20246 (N_20246,N_15594,N_18940);
nor U20247 (N_20247,N_15544,N_19058);
nand U20248 (N_20248,N_15928,N_19469);
nand U20249 (N_20249,N_19138,N_16040);
xnor U20250 (N_20250,N_15881,N_18274);
or U20251 (N_20251,N_15082,N_18574);
nor U20252 (N_20252,N_15487,N_19304);
nand U20253 (N_20253,N_19126,N_16981);
or U20254 (N_20254,N_16093,N_19063);
nor U20255 (N_20255,N_18052,N_18202);
or U20256 (N_20256,N_18110,N_16663);
and U20257 (N_20257,N_18644,N_17260);
and U20258 (N_20258,N_15648,N_18905);
nand U20259 (N_20259,N_16153,N_15157);
nand U20260 (N_20260,N_16091,N_17876);
and U20261 (N_20261,N_15349,N_15541);
nand U20262 (N_20262,N_18622,N_16207);
or U20263 (N_20263,N_15251,N_17154);
or U20264 (N_20264,N_16247,N_19718);
nand U20265 (N_20265,N_16219,N_15659);
or U20266 (N_20266,N_16878,N_16056);
nor U20267 (N_20267,N_16186,N_18298);
and U20268 (N_20268,N_16030,N_15664);
and U20269 (N_20269,N_19351,N_17603);
and U20270 (N_20270,N_16573,N_15930);
and U20271 (N_20271,N_16139,N_16317);
nand U20272 (N_20272,N_19254,N_17389);
or U20273 (N_20273,N_17358,N_15805);
or U20274 (N_20274,N_19200,N_17360);
or U20275 (N_20275,N_18309,N_15493);
or U20276 (N_20276,N_16316,N_16541);
nor U20277 (N_20277,N_17408,N_17035);
nand U20278 (N_20278,N_15404,N_19887);
or U20279 (N_20279,N_17924,N_19054);
nor U20280 (N_20280,N_15607,N_17189);
and U20281 (N_20281,N_15622,N_18660);
and U20282 (N_20282,N_16850,N_16428);
nand U20283 (N_20283,N_17728,N_18529);
and U20284 (N_20284,N_15232,N_15909);
nand U20285 (N_20285,N_19053,N_15846);
or U20286 (N_20286,N_18353,N_17988);
nor U20287 (N_20287,N_19360,N_15857);
and U20288 (N_20288,N_15387,N_19303);
and U20289 (N_20289,N_18992,N_16361);
nand U20290 (N_20290,N_18459,N_17680);
and U20291 (N_20291,N_16273,N_19585);
xnor U20292 (N_20292,N_16754,N_19550);
xor U20293 (N_20293,N_16283,N_19463);
or U20294 (N_20294,N_16583,N_15680);
or U20295 (N_20295,N_17666,N_17418);
nand U20296 (N_20296,N_16906,N_16759);
nand U20297 (N_20297,N_19484,N_19476);
and U20298 (N_20298,N_16064,N_15847);
and U20299 (N_20299,N_18690,N_17045);
and U20300 (N_20300,N_15851,N_15783);
nor U20301 (N_20301,N_16414,N_19586);
nand U20302 (N_20302,N_17796,N_17987);
or U20303 (N_20303,N_19410,N_16508);
or U20304 (N_20304,N_19665,N_18962);
nand U20305 (N_20305,N_16683,N_19436);
nand U20306 (N_20306,N_16832,N_17119);
and U20307 (N_20307,N_16250,N_17304);
or U20308 (N_20308,N_15524,N_16307);
and U20309 (N_20309,N_16282,N_18982);
nor U20310 (N_20310,N_18296,N_16036);
nor U20311 (N_20311,N_17729,N_17417);
and U20312 (N_20312,N_16204,N_15621);
or U20313 (N_20313,N_19784,N_19329);
and U20314 (N_20314,N_17731,N_16710);
nand U20315 (N_20315,N_19716,N_15873);
or U20316 (N_20316,N_15245,N_15132);
nor U20317 (N_20317,N_18165,N_17486);
nor U20318 (N_20318,N_17752,N_16345);
and U20319 (N_20319,N_15688,N_16404);
and U20320 (N_20320,N_16134,N_17345);
and U20321 (N_20321,N_15272,N_16766);
or U20322 (N_20322,N_17618,N_15409);
nand U20323 (N_20323,N_18602,N_18698);
and U20324 (N_20324,N_17354,N_18496);
and U20325 (N_20325,N_18803,N_18716);
nand U20326 (N_20326,N_18689,N_17171);
nor U20327 (N_20327,N_19556,N_15773);
or U20328 (N_20328,N_15331,N_19688);
or U20329 (N_20329,N_18142,N_18293);
or U20330 (N_20330,N_16923,N_17842);
nor U20331 (N_20331,N_19259,N_18868);
and U20332 (N_20332,N_17089,N_15148);
or U20333 (N_20333,N_19338,N_17179);
nand U20334 (N_20334,N_19651,N_16480);
and U20335 (N_20335,N_19934,N_17195);
nor U20336 (N_20336,N_15448,N_15604);
xor U20337 (N_20337,N_19886,N_17511);
or U20338 (N_20338,N_18799,N_19021);
nor U20339 (N_20339,N_16453,N_16379);
or U20340 (N_20340,N_18408,N_16546);
and U20341 (N_20341,N_17129,N_18083);
nand U20342 (N_20342,N_15538,N_15497);
and U20343 (N_20343,N_19930,N_15813);
xnor U20344 (N_20344,N_15619,N_19797);
nand U20345 (N_20345,N_18462,N_16065);
nor U20346 (N_20346,N_19776,N_19611);
nor U20347 (N_20347,N_16566,N_19669);
xnor U20348 (N_20348,N_18630,N_15318);
nand U20349 (N_20349,N_18933,N_18850);
nand U20350 (N_20350,N_18633,N_18703);
nor U20351 (N_20351,N_19158,N_19612);
nand U20352 (N_20352,N_16464,N_17479);
and U20353 (N_20353,N_15855,N_19906);
or U20354 (N_20354,N_18471,N_17392);
or U20355 (N_20355,N_16871,N_19117);
and U20356 (N_20356,N_17163,N_19427);
nor U20357 (N_20357,N_17982,N_17267);
nor U20358 (N_20358,N_17424,N_18772);
and U20359 (N_20359,N_16967,N_18533);
xnor U20360 (N_20360,N_18654,N_17279);
nand U20361 (N_20361,N_15955,N_19798);
nor U20362 (N_20362,N_16000,N_17973);
or U20363 (N_20363,N_18966,N_17159);
and U20364 (N_20364,N_16962,N_19615);
nor U20365 (N_20365,N_17807,N_15797);
nand U20366 (N_20366,N_16184,N_17614);
and U20367 (N_20367,N_15853,N_18047);
or U20368 (N_20368,N_15499,N_17525);
or U20369 (N_20369,N_17335,N_17010);
or U20370 (N_20370,N_16388,N_16697);
and U20371 (N_20371,N_16879,N_17570);
nor U20372 (N_20372,N_17646,N_19580);
and U20373 (N_20373,N_17581,N_16897);
or U20374 (N_20374,N_15517,N_16914);
nand U20375 (N_20375,N_18579,N_17470);
nand U20376 (N_20376,N_16536,N_15375);
nor U20377 (N_20377,N_18126,N_16021);
xor U20378 (N_20378,N_16168,N_15527);
and U20379 (N_20379,N_18919,N_19970);
nor U20380 (N_20380,N_15660,N_19847);
nor U20381 (N_20381,N_19105,N_18196);
nand U20382 (N_20382,N_15522,N_17832);
and U20383 (N_20383,N_19255,N_16991);
nand U20384 (N_20384,N_19595,N_15432);
nor U20385 (N_20385,N_18357,N_18480);
nand U20386 (N_20386,N_19222,N_18474);
or U20387 (N_20387,N_17659,N_17200);
nor U20388 (N_20388,N_16522,N_19551);
xor U20389 (N_20389,N_15044,N_19861);
nand U20390 (N_20390,N_17221,N_19738);
nand U20391 (N_20391,N_18168,N_15350);
nand U20392 (N_20392,N_18279,N_17593);
nand U20393 (N_20393,N_19134,N_18805);
nand U20394 (N_20394,N_15489,N_17544);
nand U20395 (N_20395,N_18643,N_17114);
or U20396 (N_20396,N_19029,N_16826);
xnor U20397 (N_20397,N_15788,N_19176);
and U20398 (N_20398,N_19543,N_17094);
nor U20399 (N_20399,N_16173,N_19645);
or U20400 (N_20400,N_17960,N_19081);
and U20401 (N_20401,N_16594,N_16852);
and U20402 (N_20402,N_18765,N_19994);
nand U20403 (N_20403,N_19089,N_17704);
nand U20404 (N_20404,N_15725,N_15511);
nand U20405 (N_20405,N_15941,N_16013);
nand U20406 (N_20406,N_19357,N_15704);
or U20407 (N_20407,N_17429,N_18219);
nor U20408 (N_20408,N_19995,N_17504);
xnor U20409 (N_20409,N_17113,N_19708);
xnor U20410 (N_20410,N_17060,N_15611);
and U20411 (N_20411,N_16605,N_15711);
nor U20412 (N_20412,N_15279,N_17866);
nand U20413 (N_20413,N_19232,N_17222);
or U20414 (N_20414,N_19783,N_16853);
nand U20415 (N_20415,N_19935,N_17181);
and U20416 (N_20416,N_15475,N_18870);
nand U20417 (N_20417,N_15792,N_16665);
and U20418 (N_20418,N_18422,N_18225);
nor U20419 (N_20419,N_15719,N_18443);
and U20420 (N_20420,N_16775,N_17742);
and U20421 (N_20421,N_15028,N_16158);
nand U20422 (N_20422,N_15801,N_16909);
and U20423 (N_20423,N_15051,N_15402);
nor U20424 (N_20424,N_18608,N_15702);
or U20425 (N_20425,N_18952,N_19929);
or U20426 (N_20426,N_17878,N_16147);
nor U20427 (N_20427,N_17042,N_17503);
nor U20428 (N_20428,N_16604,N_15975);
nand U20429 (N_20429,N_18758,N_15477);
nor U20430 (N_20430,N_18188,N_17490);
xnor U20431 (N_20431,N_19985,N_17228);
nor U20432 (N_20432,N_19793,N_16992);
nand U20433 (N_20433,N_18718,N_16112);
nand U20434 (N_20434,N_19757,N_18189);
and U20435 (N_20435,N_15900,N_16310);
and U20436 (N_20436,N_19100,N_15520);
nand U20437 (N_20437,N_18139,N_17574);
or U20438 (N_20438,N_16187,N_18696);
nand U20439 (N_20439,N_18505,N_18249);
nor U20440 (N_20440,N_16619,N_18368);
nand U20441 (N_20441,N_15363,N_15963);
nor U20442 (N_20442,N_19414,N_19274);
nor U20443 (N_20443,N_17427,N_15706);
nor U20444 (N_20444,N_17984,N_18769);
nand U20445 (N_20445,N_19354,N_16622);
nor U20446 (N_20446,N_18653,N_17976);
or U20447 (N_20447,N_15271,N_15737);
nand U20448 (N_20448,N_18846,N_19843);
and U20449 (N_20449,N_15882,N_16434);
nor U20450 (N_20450,N_16735,N_15636);
and U20451 (N_20451,N_16324,N_19109);
xor U20452 (N_20452,N_19872,N_17889);
nor U20453 (N_20453,N_19990,N_17147);
and U20454 (N_20454,N_15829,N_17573);
and U20455 (N_20455,N_16202,N_16681);
nor U20456 (N_20456,N_15228,N_19570);
nor U20457 (N_20457,N_19981,N_18647);
nor U20458 (N_20458,N_17990,N_17978);
nand U20459 (N_20459,N_18238,N_18406);
and U20460 (N_20460,N_15774,N_17860);
or U20461 (N_20461,N_18790,N_18134);
nand U20462 (N_20462,N_17109,N_17575);
or U20463 (N_20463,N_16883,N_18288);
nor U20464 (N_20464,N_15292,N_17937);
and U20465 (N_20465,N_16181,N_17843);
or U20466 (N_20466,N_19529,N_19010);
nand U20467 (N_20467,N_19524,N_17483);
nand U20468 (N_20468,N_17052,N_16255);
or U20469 (N_20469,N_16083,N_17846);
or U20470 (N_20470,N_18874,N_19916);
or U20471 (N_20471,N_17172,N_19711);
and U20472 (N_20472,N_18205,N_18043);
xnor U20473 (N_20473,N_16899,N_15290);
nand U20474 (N_20474,N_18458,N_17187);
nand U20475 (N_20475,N_17062,N_17734);
or U20476 (N_20476,N_15565,N_15159);
and U20477 (N_20477,N_16475,N_17955);
or U20478 (N_20478,N_15883,N_16405);
nor U20479 (N_20479,N_18263,N_19403);
and U20480 (N_20480,N_15924,N_18764);
and U20481 (N_20481,N_16623,N_19103);
or U20482 (N_20482,N_17442,N_16124);
nor U20483 (N_20483,N_17134,N_16753);
nand U20484 (N_20484,N_19225,N_18257);
nor U20485 (N_20485,N_19553,N_15395);
nor U20486 (N_20486,N_17554,N_16020);
nor U20487 (N_20487,N_19745,N_17962);
and U20488 (N_20488,N_16644,N_16109);
nand U20489 (N_20489,N_16506,N_16195);
nor U20490 (N_20490,N_15754,N_16526);
or U20491 (N_20491,N_18843,N_16466);
and U20492 (N_20492,N_19453,N_19499);
nor U20493 (N_20493,N_19073,N_19831);
nor U20494 (N_20494,N_16420,N_15764);
and U20495 (N_20495,N_15216,N_16120);
nand U20496 (N_20496,N_19183,N_17509);
nand U20497 (N_20497,N_19987,N_18720);
or U20498 (N_20498,N_16127,N_16130);
and U20499 (N_20499,N_15961,N_19057);
nor U20500 (N_20500,N_16286,N_16025);
nand U20501 (N_20501,N_15988,N_15856);
nand U20502 (N_20502,N_15786,N_17111);
nor U20503 (N_20503,N_15584,N_15715);
or U20504 (N_20504,N_15302,N_19236);
and U20505 (N_20505,N_17439,N_18435);
xor U20506 (N_20506,N_15508,N_18669);
or U20507 (N_20507,N_17199,N_17460);
or U20508 (N_20508,N_16476,N_17394);
or U20509 (N_20509,N_17006,N_15080);
nor U20510 (N_20510,N_19859,N_19402);
and U20511 (N_20511,N_17031,N_15482);
nor U20512 (N_20512,N_16835,N_15739);
and U20513 (N_20513,N_15506,N_17491);
nor U20514 (N_20514,N_15962,N_16861);
and U20515 (N_20515,N_19622,N_16949);
or U20516 (N_20516,N_18763,N_19721);
and U20517 (N_20517,N_17857,N_19870);
nor U20518 (N_20518,N_17847,N_16165);
xor U20519 (N_20519,N_18885,N_19956);
and U20520 (N_20520,N_17327,N_16384);
nor U20521 (N_20521,N_19786,N_16357);
and U20522 (N_20522,N_18082,N_19821);
nand U20523 (N_20523,N_15020,N_16237);
or U20524 (N_20524,N_18364,N_17709);
nand U20525 (N_20525,N_19297,N_17777);
nand U20526 (N_20526,N_15052,N_18968);
and U20527 (N_20527,N_15049,N_17023);
nor U20528 (N_20528,N_18818,N_15561);
xnor U20529 (N_20529,N_15807,N_17715);
and U20530 (N_20530,N_15481,N_19133);
nor U20531 (N_20531,N_15346,N_17967);
or U20532 (N_20532,N_15919,N_19210);
nand U20533 (N_20533,N_17622,N_19415);
nor U20534 (N_20534,N_17183,N_15556);
and U20535 (N_20535,N_19366,N_15059);
xnor U20536 (N_20536,N_16578,N_16596);
nor U20537 (N_20537,N_18502,N_17388);
or U20538 (N_20538,N_15674,N_15239);
nor U20539 (N_20539,N_19179,N_18640);
nor U20540 (N_20540,N_18484,N_18884);
nand U20541 (N_20541,N_18656,N_19382);
xor U20542 (N_20542,N_17446,N_17650);
and U20543 (N_20543,N_16145,N_17861);
nor U20544 (N_20544,N_19880,N_17003);
and U20545 (N_20545,N_18042,N_19982);
nand U20546 (N_20546,N_19490,N_15570);
or U20547 (N_20547,N_16979,N_18122);
nor U20548 (N_20548,N_17012,N_15104);
nor U20549 (N_20549,N_16746,N_18067);
nor U20550 (N_20550,N_18173,N_18547);
or U20551 (N_20551,N_19875,N_18651);
nand U20552 (N_20552,N_16499,N_17501);
xnor U20553 (N_20553,N_15000,N_15926);
nor U20554 (N_20554,N_18620,N_17105);
or U20555 (N_20555,N_15914,N_17453);
and U20556 (N_20556,N_18391,N_17311);
nor U20557 (N_20557,N_16073,N_17814);
nor U20558 (N_20558,N_17220,N_16162);
nand U20559 (N_20559,N_17300,N_18439);
nor U20560 (N_20560,N_17271,N_16511);
nand U20561 (N_20561,N_16787,N_19313);
nand U20562 (N_20562,N_17730,N_18405);
nand U20563 (N_20563,N_18518,N_18544);
nor U20564 (N_20564,N_15531,N_19310);
nand U20565 (N_20565,N_16924,N_16244);
and U20566 (N_20566,N_16291,N_16243);
and U20567 (N_20567,N_15360,N_17944);
nand U20568 (N_20568,N_19672,N_16827);
or U20569 (N_20569,N_19397,N_15361);
and U20570 (N_20570,N_15061,N_17321);
nand U20571 (N_20571,N_16193,N_15530);
or U20572 (N_20572,N_18495,N_16051);
nor U20573 (N_20573,N_15057,N_16362);
xor U20574 (N_20574,N_19347,N_18673);
nor U20575 (N_20575,N_16679,N_17557);
nor U20576 (N_20576,N_17083,N_15415);
and U20577 (N_20577,N_15705,N_17071);
xnor U20578 (N_20578,N_18226,N_18180);
or U20579 (N_20579,N_17077,N_18028);
and U20580 (N_20580,N_16702,N_16076);
or U20581 (N_20581,N_17258,N_16159);
xor U20582 (N_20582,N_19966,N_15922);
nor U20583 (N_20583,N_16582,N_18115);
nor U20584 (N_20584,N_17661,N_16969);
and U20585 (N_20585,N_18444,N_19794);
nor U20586 (N_20586,N_18823,N_19787);
and U20587 (N_20587,N_16095,N_16426);
and U20588 (N_20588,N_15032,N_16114);
or U20589 (N_20589,N_17329,N_15235);
or U20590 (N_20590,N_19075,N_18000);
nor U20591 (N_20591,N_17652,N_15753);
xnor U20592 (N_20592,N_15208,N_15321);
nand U20593 (N_20593,N_16067,N_19396);
and U20594 (N_20594,N_17288,N_15762);
or U20595 (N_20595,N_16033,N_17211);
xnor U20596 (N_20596,N_15981,N_17148);
or U20597 (N_20597,N_16574,N_19475);
nor U20598 (N_20598,N_19478,N_16579);
xor U20599 (N_20599,N_18066,N_18511);
or U20600 (N_20600,N_19824,N_16912);
and U20601 (N_20601,N_15274,N_18449);
nor U20602 (N_20602,N_15871,N_17009);
or U20603 (N_20603,N_15352,N_18411);
nand U20604 (N_20604,N_19321,N_19532);
nor U20605 (N_20605,N_16146,N_19269);
nand U20606 (N_20606,N_16699,N_17150);
xor U20607 (N_20607,N_17875,N_15550);
and U20608 (N_20608,N_17140,N_19016);
and U20609 (N_20609,N_19849,N_18963);
xnor U20610 (N_20610,N_19395,N_19362);
and U20611 (N_20611,N_16678,N_18076);
nor U20612 (N_20612,N_16645,N_19905);
or U20613 (N_20613,N_18235,N_16814);
nand U20614 (N_20614,N_18523,N_19068);
nand U20615 (N_20615,N_17589,N_15436);
nand U20616 (N_20616,N_18104,N_19441);
and U20617 (N_20617,N_18955,N_18568);
xnor U20618 (N_20618,N_18399,N_16577);
nor U20619 (N_20619,N_16552,N_17324);
and U20620 (N_20620,N_19795,N_17612);
and U20621 (N_20621,N_18308,N_18310);
nand U20622 (N_20622,N_15905,N_19640);
nand U20623 (N_20623,N_17475,N_17678);
and U20624 (N_20624,N_19618,N_16737);
nand U20625 (N_20625,N_16191,N_17706);
nand U20626 (N_20626,N_17346,N_19005);
or U20627 (N_20627,N_18046,N_17601);
and U20628 (N_20628,N_18702,N_17380);
and U20629 (N_20629,N_16950,N_17656);
nor U20630 (N_20630,N_18229,N_15918);
or U20631 (N_20631,N_18524,N_19048);
and U20632 (N_20632,N_16668,N_19860);
nor U20633 (N_20633,N_19502,N_19178);
nor U20634 (N_20634,N_19632,N_17645);
nand U20635 (N_20635,N_18007,N_15519);
nor U20636 (N_20636,N_19271,N_17124);
nor U20637 (N_20637,N_17838,N_19182);
nand U20638 (N_20638,N_19978,N_19627);
and U20639 (N_20639,N_17534,N_16309);
nor U20640 (N_20640,N_16695,N_17160);
xor U20641 (N_20641,N_16052,N_16262);
or U20642 (N_20642,N_17681,N_17892);
or U20643 (N_20643,N_17949,N_19567);
or U20644 (N_20644,N_16762,N_16133);
or U20645 (N_20645,N_17748,N_16224);
and U20646 (N_20646,N_15625,N_18596);
and U20647 (N_20647,N_17623,N_17438);
nor U20648 (N_20648,N_15430,N_16081);
xnor U20649 (N_20649,N_18889,N_16259);
and U20650 (N_20650,N_18351,N_15912);
and U20651 (N_20651,N_18314,N_19305);
or U20652 (N_20652,N_18324,N_15303);
and U20653 (N_20653,N_18925,N_15849);
nor U20654 (N_20654,N_18097,N_18701);
nor U20655 (N_20655,N_15369,N_16671);
or U20656 (N_20656,N_19868,N_16892);
or U20657 (N_20657,N_19957,N_15323);
or U20658 (N_20658,N_19394,N_18019);
or U20659 (N_20659,N_18866,N_17312);
nor U20660 (N_20660,N_18499,N_16171);
nor U20661 (N_20661,N_16728,N_16490);
and U20662 (N_20662,N_17947,N_16047);
nand U20663 (N_20663,N_15265,N_19235);
nand U20664 (N_20664,N_19959,N_18542);
nor U20665 (N_20665,N_16189,N_17338);
nor U20666 (N_20666,N_15789,N_18871);
or U20667 (N_20667,N_17720,N_19231);
or U20668 (N_20668,N_15215,N_15694);
nor U20669 (N_20669,N_17834,N_18809);
or U20670 (N_20670,N_18215,N_16182);
nand U20671 (N_20671,N_19292,N_15109);
or U20672 (N_20672,N_15599,N_18900);
and U20673 (N_20673,N_16400,N_16828);
nor U20674 (N_20674,N_17610,N_15003);
nand U20675 (N_20675,N_17120,N_15578);
or U20676 (N_20676,N_16531,N_19348);
or U20677 (N_20677,N_18363,N_18751);
and U20678 (N_20678,N_19922,N_19112);
xnor U20679 (N_20679,N_16393,N_15501);
nor U20680 (N_20680,N_18915,N_19326);
nand U20681 (N_20681,N_18881,N_18409);
or U20682 (N_20682,N_18562,N_17792);
or U20683 (N_20683,N_17158,N_16755);
and U20684 (N_20684,N_19001,N_16367);
xnor U20685 (N_20685,N_16926,N_16394);
or U20686 (N_20686,N_18795,N_19825);
nand U20687 (N_20687,N_18098,N_15429);
or U20688 (N_20688,N_18561,N_19941);
xnor U20689 (N_20689,N_16467,N_16113);
xor U20690 (N_20690,N_15934,N_15240);
xor U20691 (N_20691,N_19693,N_16217);
nor U20692 (N_20692,N_15455,N_16211);
or U20693 (N_20693,N_15631,N_18678);
nor U20694 (N_20694,N_18909,N_16089);
nor U20695 (N_20695,N_16614,N_18890);
nand U20696 (N_20696,N_19458,N_18628);
nand U20697 (N_20697,N_19020,N_17663);
or U20698 (N_20698,N_19108,N_19241);
nor U20699 (N_20699,N_19710,N_16829);
nor U20700 (N_20700,N_15670,N_16206);
nor U20701 (N_20701,N_18362,N_17611);
nor U20702 (N_20702,N_17217,N_15102);
nor U20703 (N_20703,N_19677,N_16625);
nand U20704 (N_20704,N_17085,N_15067);
and U20705 (N_20705,N_18243,N_19845);
xnor U20706 (N_20706,N_16586,N_15300);
nor U20707 (N_20707,N_17241,N_16978);
nand U20708 (N_20708,N_16650,N_19583);
and U20709 (N_20709,N_15645,N_18036);
nand U20710 (N_20710,N_15419,N_17232);
xor U20711 (N_20711,N_15824,N_19472);
nor U20712 (N_20712,N_19171,N_16246);
nand U20713 (N_20713,N_19185,N_16174);
nor U20714 (N_20714,N_18625,N_19092);
and U20715 (N_20715,N_18468,N_17858);
and U20716 (N_20716,N_19661,N_15327);
or U20717 (N_20717,N_15178,N_18517);
nand U20718 (N_20718,N_18381,N_15056);
nand U20719 (N_20719,N_19342,N_15586);
xnor U20720 (N_20720,N_19181,N_15876);
and U20721 (N_20721,N_19522,N_15572);
or U20722 (N_20722,N_15267,N_17771);
and U20723 (N_20723,N_18532,N_16704);
nor U20724 (N_20724,N_17772,N_18365);
and U20725 (N_20725,N_19755,N_18374);
nand U20726 (N_20726,N_18508,N_17038);
nand U20727 (N_20727,N_18491,N_16615);
nor U20728 (N_20728,N_18831,N_18892);
nor U20729 (N_20729,N_17118,N_18609);
or U20730 (N_20730,N_18125,N_18906);
xnor U20731 (N_20731,N_19358,N_19211);
nand U20732 (N_20732,N_17367,N_16919);
and U20733 (N_20733,N_19913,N_18255);
nand U20734 (N_20734,N_18637,N_16274);
and U20735 (N_20735,N_16631,N_17998);
nand U20736 (N_20736,N_17999,N_18961);
nor U20737 (N_20737,N_16649,N_15140);
and U20738 (N_20738,N_15859,N_19903);
or U20739 (N_20739,N_16203,N_19203);
and U20740 (N_20740,N_15054,N_17854);
nor U20741 (N_20741,N_19882,N_15246);
or U20742 (N_20742,N_16955,N_19538);
nand U20743 (N_20743,N_19102,N_18590);
xnor U20744 (N_20744,N_18942,N_18001);
or U20745 (N_20745,N_15194,N_19162);
and U20746 (N_20746,N_17449,N_16331);
nor U20747 (N_20747,N_17867,N_15401);
and U20748 (N_20748,N_16889,N_19614);
or U20749 (N_20749,N_18717,N_19867);
nand U20750 (N_20750,N_19153,N_17906);
and U20751 (N_20751,N_18744,N_18995);
nor U20752 (N_20752,N_16609,N_16997);
or U20753 (N_20753,N_15030,N_18655);
nor U20754 (N_20754,N_19026,N_15440);
nor U20755 (N_20755,N_18615,N_16401);
nor U20756 (N_20756,N_19331,N_19457);
nor U20757 (N_20757,N_17675,N_17820);
or U20758 (N_20758,N_16132,N_16780);
and U20759 (N_20759,N_18724,N_16385);
nand U20760 (N_20760,N_17384,N_19856);
or U20761 (N_20761,N_16752,N_19604);
and U20762 (N_20762,N_19997,N_15833);
nor U20763 (N_20763,N_15071,N_15207);
and U20764 (N_20764,N_17143,N_17326);
and U20765 (N_20765,N_16726,N_15287);
and U20766 (N_20766,N_17084,N_15142);
nor U20767 (N_20767,N_19526,N_15115);
and U20768 (N_20768,N_19208,N_15330);
and U20769 (N_20769,N_19359,N_17827);
and U20770 (N_20770,N_17428,N_16321);
nor U20771 (N_20771,N_17514,N_16970);
nor U20772 (N_20772,N_16024,N_16504);
nor U20773 (N_20773,N_16141,N_15770);
nor U20774 (N_20774,N_17821,N_19468);
nor U20775 (N_20775,N_18838,N_15177);
nand U20776 (N_20776,N_15820,N_16449);
nand U20777 (N_20777,N_17558,N_15260);
and U20778 (N_20778,N_17323,N_18573);
and U20779 (N_20779,N_16646,N_18947);
nand U20780 (N_20780,N_17936,N_16409);
nand U20781 (N_20781,N_16129,N_19961);
nor U20782 (N_20782,N_16974,N_18883);
nor U20783 (N_20783,N_16212,N_19413);
xor U20784 (N_20784,N_18627,N_15800);
or U20785 (N_20785,N_19660,N_15875);
nand U20786 (N_20786,N_17787,N_18345);
nand U20787 (N_20787,N_16535,N_16751);
nand U20788 (N_20788,N_16399,N_17727);
or U20789 (N_20789,N_18081,N_19844);
nor U20790 (N_20790,N_17457,N_17272);
and U20791 (N_20791,N_16482,N_15491);
and U20792 (N_20792,N_15993,N_17567);
nor U20793 (N_20793,N_17994,N_15062);
or U20794 (N_20794,N_16017,N_19352);
nor U20795 (N_20795,N_16525,N_15066);
nand U20796 (N_20796,N_17069,N_19657);
or U20797 (N_20797,N_19931,N_17918);
nor U20798 (N_20798,N_16980,N_18935);
or U20799 (N_20799,N_18631,N_18476);
nand U20800 (N_20800,N_17316,N_18852);
nand U20801 (N_20801,N_19851,N_18040);
or U20802 (N_20802,N_15420,N_17125);
nand U20803 (N_20803,N_18965,N_18956);
xnor U20804 (N_20804,N_15828,N_17494);
nor U20805 (N_20805,N_16094,N_18079);
nand U20806 (N_20806,N_15095,N_17224);
nand U20807 (N_20807,N_18867,N_18137);
or U20808 (N_20808,N_17308,N_18352);
and U20809 (N_20809,N_19251,N_16268);
nor U20810 (N_20810,N_19345,N_16102);
and U20811 (N_20811,N_18003,N_16136);
xnor U20812 (N_20812,N_19936,N_16823);
nand U20813 (N_20813,N_16483,N_19748);
nand U20814 (N_20814,N_19501,N_17341);
nor U20815 (N_20815,N_15663,N_19226);
xnor U20816 (N_20816,N_15433,N_17585);
or U20817 (N_20817,N_19827,N_18190);
nor U20818 (N_20818,N_18844,N_18762);
or U20819 (N_20819,N_18879,N_17948);
or U20820 (N_20820,N_17887,N_18455);
nor U20821 (N_20821,N_18575,N_18426);
nand U20822 (N_20822,N_16383,N_19032);
and U20823 (N_20823,N_18604,N_19030);
and U20824 (N_20824,N_19015,N_15236);
or U20825 (N_20825,N_16258,N_17969);
or U20826 (N_20826,N_18420,N_19128);
nor U20827 (N_20827,N_19911,N_17291);
and U20828 (N_20828,N_19920,N_15380);
nor U20829 (N_20829,N_18256,N_15206);
or U20830 (N_20830,N_16724,N_18957);
nor U20831 (N_20831,N_18814,N_15394);
or U20832 (N_20832,N_16323,N_16177);
and U20833 (N_20833,N_16429,N_19175);
xnor U20834 (N_20834,N_18158,N_18739);
and U20835 (N_20835,N_18641,N_16192);
and U20836 (N_20836,N_18200,N_18777);
nand U20837 (N_20837,N_19833,N_18742);
or U20838 (N_20838,N_19652,N_19826);
xnor U20839 (N_20839,N_17136,N_15910);
nand U20840 (N_20840,N_17850,N_17402);
nor U20841 (N_20841,N_15760,N_19088);
or U20842 (N_20842,N_19873,N_15579);
and U20843 (N_20843,N_18770,N_17505);
xor U20844 (N_20844,N_16278,N_17344);
or U20845 (N_20845,N_16836,N_19386);
or U20846 (N_20846,N_18300,N_19836);
or U20847 (N_20847,N_15547,N_18261);
nor U20848 (N_20848,N_18854,N_15048);
xor U20849 (N_20849,N_18564,N_19898);
and U20850 (N_20850,N_16312,N_15861);
nor U20851 (N_20851,N_18726,N_19539);
nand U20852 (N_20852,N_16257,N_16427);
or U20853 (N_20853,N_16885,N_18827);
and U20854 (N_20854,N_16451,N_18153);
nor U20855 (N_20855,N_17059,N_17565);
and U20856 (N_20856,N_16437,N_15954);
xor U20857 (N_20857,N_16110,N_17231);
nand U20858 (N_20858,N_19684,N_18050);
nor U20859 (N_20859,N_15740,N_17977);
nor U20860 (N_20860,N_16407,N_18789);
nor U20861 (N_20861,N_16456,N_17649);
nand U20862 (N_20862,N_16225,N_19401);
nand U20863 (N_20863,N_16078,N_16779);
nor U20864 (N_20864,N_17552,N_16990);
nand U20865 (N_20865,N_16172,N_16122);
nor U20866 (N_20866,N_17774,N_17532);
and U20867 (N_20867,N_15678,N_18211);
or U20868 (N_20868,N_18185,N_15063);
and U20869 (N_20869,N_16868,N_16417);
nand U20870 (N_20870,N_19996,N_19971);
xnor U20871 (N_20871,N_17855,N_19517);
nand U20872 (N_20872,N_15087,N_16178);
and U20873 (N_20873,N_16845,N_17314);
nand U20874 (N_20874,N_16444,N_15528);
nand U20875 (N_20875,N_17342,N_19646);
or U20876 (N_20876,N_17448,N_17092);
or U20877 (N_20877,N_17794,N_15450);
or U20878 (N_20878,N_19291,N_18632);
nand U20879 (N_20879,N_18642,N_19284);
nand U20880 (N_20880,N_16763,N_16777);
xnor U20881 (N_20881,N_16284,N_15358);
or U20882 (N_20882,N_15336,N_16590);
nor U20883 (N_20883,N_15076,N_17841);
nand U20884 (N_20884,N_17528,N_15887);
xnor U20885 (N_20885,N_15612,N_15308);
and U20886 (N_20886,N_18155,N_17737);
nor U20887 (N_20887,N_15460,N_18005);
xnor U20888 (N_20888,N_15892,N_15333);
and U20889 (N_20889,N_15305,N_16300);
nand U20890 (N_20890,N_19013,N_15043);
and U20891 (N_20891,N_19034,N_16632);
xor U20892 (N_20892,N_19107,N_15150);
xnor U20893 (N_20893,N_19509,N_17631);
nand U20894 (N_20894,N_16524,N_16126);
nor U20895 (N_20895,N_15687,N_19494);
nor U20896 (N_20896,N_16014,N_19161);
or U20897 (N_20897,N_17257,N_19299);
or U20898 (N_20898,N_17274,N_18570);
or U20899 (N_20899,N_17303,N_17713);
or U20900 (N_20900,N_17091,N_18791);
nand U20901 (N_20901,N_17123,N_15627);
and U20902 (N_20902,N_18684,N_18415);
and U20903 (N_20903,N_15927,N_19482);
xnor U20904 (N_20904,N_19962,N_19811);
nor U20905 (N_20905,N_18652,N_18521);
and U20906 (N_20906,N_19659,N_19687);
xnor U20907 (N_20907,N_18780,N_18062);
xnor U20908 (N_20908,N_15582,N_18741);
xor U20909 (N_20909,N_17929,N_19574);
nor U20910 (N_20910,N_16887,N_17979);
xor U20911 (N_20911,N_16135,N_18695);
xnor U20912 (N_20912,N_17926,N_15730);
nand U20913 (N_20913,N_15738,N_16716);
and U20914 (N_20914,N_19506,N_18939);
or U20915 (N_20915,N_17975,N_17112);
xnor U20916 (N_20916,N_19670,N_16610);
or U20917 (N_20917,N_17635,N_15609);
xor U20918 (N_20918,N_16782,N_18671);
nand U20919 (N_20919,N_19077,N_16450);
nor U20920 (N_20920,N_18423,N_17687);
nor U20921 (N_20921,N_17917,N_17078);
xnor U20922 (N_20922,N_17613,N_17431);
nand U20923 (N_20923,N_17683,N_17387);
or U20924 (N_20924,N_16115,N_16306);
and U20925 (N_20925,N_17357,N_19041);
or U20926 (N_20926,N_15269,N_16415);
xnor U20927 (N_20927,N_18014,N_16349);
or U20928 (N_20928,N_18806,N_19060);
and U20929 (N_20929,N_19166,N_17641);
or U20930 (N_20930,N_16397,N_17662);
nand U20931 (N_20931,N_19818,N_19679);
or U20932 (N_20932,N_17670,N_19503);
or U20933 (N_20933,N_16519,N_19531);
nand U20934 (N_20934,N_17348,N_19002);
or U20935 (N_20935,N_18297,N_19563);
nor U20936 (N_20936,N_18397,N_16567);
nor U20937 (N_20937,N_19071,N_15478);
or U20938 (N_20938,N_19132,N_17265);
xnor U20939 (N_20939,N_17518,N_18531);
nand U20940 (N_20940,N_15386,N_17297);
nor U20941 (N_20941,N_18093,N_16495);
nor U20942 (N_20942,N_16564,N_17914);
nor U20943 (N_20943,N_15536,N_19520);
nand U20944 (N_20944,N_18930,N_18287);
nor U20945 (N_20945,N_19983,N_15141);
or U20946 (N_20946,N_15576,N_16164);
or U20947 (N_20947,N_15081,N_17506);
nor U20948 (N_20948,N_17986,N_16408);
and U20949 (N_20949,N_18676,N_17809);
xnor U20950 (N_20950,N_15367,N_17454);
nand U20951 (N_20951,N_15100,N_17028);
nor U20952 (N_20952,N_15726,N_19377);
or U20953 (N_20953,N_15903,N_16285);
nor U20954 (N_20954,N_15676,N_15069);
nor U20955 (N_20955,N_19471,N_17714);
xnor U20956 (N_20956,N_17157,N_17717);
nor U20957 (N_20957,N_15408,N_17406);
or U20958 (N_20958,N_16662,N_15869);
xnor U20959 (N_20959,N_19151,N_17458);
and U20960 (N_20960,N_19919,N_19375);
or U20961 (N_20961,N_18023,N_18394);
xnor U20962 (N_20962,N_16335,N_18938);
and U20963 (N_20963,N_17776,N_15911);
xnor U20964 (N_20964,N_18131,N_15029);
nand U20965 (N_20965,N_18526,N_18829);
nand U20966 (N_20966,N_17334,N_18754);
xnor U20967 (N_20967,N_16549,N_16302);
nand U20968 (N_20968,N_16954,N_16118);
and U20969 (N_20969,N_19799,N_17997);
and U20970 (N_20970,N_18578,N_18454);
nor U20971 (N_20971,N_17829,N_17922);
xnor U20972 (N_20972,N_18559,N_19775);
or U20973 (N_20973,N_18830,N_15731);
xnor U20974 (N_20974,N_16027,N_15870);
nand U20975 (N_20975,N_19302,N_18268);
nand U20976 (N_20976,N_19062,N_19150);
and U20977 (N_20977,N_19609,N_19883);
and U20978 (N_20978,N_16784,N_17952);
nand U20979 (N_20979,N_18851,N_17478);
nand U20980 (N_20980,N_18222,N_19591);
nor U20981 (N_20981,N_19976,N_15899);
nand U20982 (N_20982,N_18228,N_17305);
nor U20983 (N_20983,N_15686,N_17477);
and U20984 (N_20984,N_17536,N_18475);
or U20985 (N_20985,N_19098,N_19769);
or U20986 (N_20986,N_19802,N_17718);
or U20987 (N_20987,N_16554,N_17056);
and U20988 (N_20988,N_15325,N_18986);
and U20989 (N_20989,N_17564,N_15854);
nand U20990 (N_20990,N_15897,N_16333);
nor U20991 (N_20991,N_18431,N_16865);
nand U20992 (N_20992,N_16776,N_18845);
or U20993 (N_20993,N_18330,N_17350);
or U20994 (N_20994,N_16382,N_18111);
xnor U20995 (N_20995,N_15053,N_18254);
and U20996 (N_20996,N_16568,N_16150);
or U20997 (N_20997,N_19419,N_18721);
xor U20998 (N_20998,N_17459,N_18639);
or U20999 (N_20999,N_19655,N_16765);
and U21000 (N_21000,N_16080,N_17166);
nor U21001 (N_21001,N_15976,N_17954);
and U21002 (N_21002,N_17775,N_15758);
or U21003 (N_21003,N_17218,N_19773);
and U21004 (N_21004,N_17655,N_18203);
or U21005 (N_21005,N_15237,N_17698);
xor U21006 (N_21006,N_18218,N_16327);
nor U21007 (N_21007,N_19869,N_16131);
nor U21008 (N_21008,N_18988,N_15169);
nand U21009 (N_21009,N_17881,N_16669);
or U21010 (N_21010,N_17739,N_16550);
xor U21011 (N_21011,N_19148,N_19865);
nor U21012 (N_21012,N_17047,N_19330);
nand U21013 (N_21013,N_16700,N_17481);
or U21014 (N_21014,N_17945,N_15974);
or U21015 (N_21015,N_15045,N_17127);
and U21016 (N_21016,N_17756,N_17634);
nand U21017 (N_21017,N_18132,N_19374);
or U21018 (N_21018,N_15189,N_17254);
or U21019 (N_21019,N_15987,N_15613);
and U21020 (N_21020,N_19237,N_16325);
nand U21021 (N_21021,N_18100,N_17227);
nor U21022 (N_21022,N_16713,N_15867);
and U21023 (N_21023,N_18504,N_17836);
and U21024 (N_21024,N_19435,N_16183);
nor U21025 (N_21025,N_17339,N_17953);
nand U21026 (N_21026,N_19910,N_15713);
nor U21027 (N_21027,N_18380,N_19385);
xnor U21028 (N_21028,N_18592,N_17865);
or U21029 (N_21029,N_19510,N_18267);
and U21030 (N_21030,N_15250,N_19834);
nand U21031 (N_21031,N_15776,N_18029);
or U21032 (N_21032,N_17637,N_19433);
nand U21033 (N_21033,N_16548,N_19219);
xnor U21034 (N_21034,N_17499,N_19253);
or U21035 (N_21035,N_17399,N_17694);
nand U21036 (N_21036,N_16983,N_17053);
or U21037 (N_21037,N_18490,N_16199);
nand U21038 (N_21038,N_16819,N_16389);
nand U21039 (N_21039,N_19803,N_18776);
nor U21040 (N_21040,N_17500,N_19637);
xnor U21041 (N_21041,N_18305,N_17770);
nand U21042 (N_21042,N_15060,N_17884);
or U21043 (N_21043,N_15535,N_19681);
nor U21044 (N_21044,N_15652,N_16045);
and U21045 (N_21045,N_18796,N_15916);
nor U21046 (N_21046,N_16778,N_19004);
and U21047 (N_21047,N_19318,N_18077);
nand U21048 (N_21048,N_19031,N_16764);
nand U21049 (N_21049,N_16063,N_18116);
and U21050 (N_21050,N_18664,N_17746);
and U21051 (N_21051,N_17871,N_19418);
nand U21052 (N_21052,N_15502,N_19535);
nor U21053 (N_21053,N_18820,N_17216);
and U21054 (N_21054,N_16860,N_15830);
or U21055 (N_21055,N_18413,N_15468);
or U21056 (N_21056,N_15008,N_16565);
xnor U21057 (N_21057,N_18949,N_18506);
nand U21058 (N_21058,N_16469,N_16004);
and U21059 (N_21059,N_18904,N_18402);
nor U21060 (N_21060,N_18591,N_17055);
xnor U21061 (N_21061,N_15785,N_18361);
nor U21062 (N_21062,N_17815,N_19129);
nand U21063 (N_21063,N_19766,N_17375);
xor U21064 (N_21064,N_18707,N_17608);
xor U21065 (N_21065,N_15443,N_18978);
or U21066 (N_21066,N_17203,N_18543);
nand U21067 (N_21067,N_16337,N_18327);
and U21068 (N_21068,N_15257,N_15574);
and U21069 (N_21069,N_19696,N_16463);
nor U21070 (N_21070,N_15442,N_19857);
and U21071 (N_21071,N_15885,N_19774);
and U21072 (N_21072,N_15698,N_15210);
and U21073 (N_21073,N_17874,N_16200);
nand U21074 (N_21074,N_17188,N_16338);
or U21075 (N_21075,N_16952,N_17545);
nand U21076 (N_21076,N_17711,N_19606);
and U21077 (N_21077,N_19474,N_15736);
xnor U21078 (N_21078,N_16484,N_18513);
and U21079 (N_21079,N_16682,N_15016);
nand U21080 (N_21080,N_19189,N_18941);
xnor U21081 (N_21081,N_16082,N_15837);
and U21082 (N_21082,N_15403,N_19674);
or U21083 (N_21083,N_19244,N_15158);
and U21084 (N_21084,N_16342,N_15880);
or U21085 (N_21085,N_18241,N_17703);
and U21086 (N_21086,N_18603,N_15709);
and U21087 (N_21087,N_15767,N_16053);
xnor U21088 (N_21088,N_16616,N_19616);
nor U21089 (N_21089,N_17898,N_18784);
xor U21090 (N_21090,N_15986,N_19059);
and U21091 (N_21091,N_17606,N_16188);
nor U21092 (N_21092,N_19250,N_16354);
nand U21093 (N_21093,N_17276,N_19283);
nand U21094 (N_21094,N_16459,N_19719);
nand U21095 (N_21095,N_17169,N_16294);
and U21096 (N_21096,N_19723,N_16447);
nor U21097 (N_21097,N_15353,N_18198);
nand U21098 (N_21098,N_18441,N_15035);
nor U21099 (N_21099,N_18147,N_19091);
nand U21100 (N_21100,N_15618,N_17543);
and U21101 (N_21101,N_16142,N_16690);
or U21102 (N_21102,N_19497,N_19115);
nand U21103 (N_21103,N_18075,N_19228);
nor U21104 (N_21104,N_19946,N_19339);
nor U21105 (N_21105,N_19528,N_19724);
or U21106 (N_21106,N_18265,N_15155);
nand U21107 (N_21107,N_15184,N_17194);
or U21108 (N_21108,N_18291,N_17333);
or U21109 (N_21109,N_15845,N_18990);
and U21110 (N_21110,N_19634,N_17102);
nor U21111 (N_21111,N_19690,N_18460);
and U21112 (N_21112,N_16232,N_17789);
nor U21113 (N_21113,N_17921,N_19518);
nand U21114 (N_21114,N_19298,N_19040);
or U21115 (N_21115,N_19714,N_15965);
or U21116 (N_21116,N_19281,N_17579);
nand U21117 (N_21117,N_17050,N_19085);
nor U21118 (N_21118,N_15471,N_16106);
and U21119 (N_21119,N_16788,N_16088);
and U21120 (N_21120,N_17643,N_15819);
xnor U21121 (N_21121,N_17041,N_19094);
nor U21122 (N_21122,N_17251,N_19561);
and U21123 (N_21123,N_16527,N_17951);
and U21124 (N_21124,N_15467,N_19767);
or U21125 (N_21125,N_18745,N_19697);
nor U21126 (N_21126,N_16518,N_19763);
nor U21127 (N_21127,N_19548,N_19513);
or U21128 (N_21128,N_19741,N_16368);
or U21129 (N_21129,N_16895,N_16074);
and U21130 (N_21130,N_18510,N_18440);
nor U21131 (N_21131,N_18912,N_16770);
or U21132 (N_21132,N_19489,N_16873);
nor U21133 (N_21133,N_16838,N_18662);
or U21134 (N_21134,N_16570,N_17527);
nor U21135 (N_21135,N_19373,N_17609);
or U21136 (N_21136,N_17482,N_16265);
nor U21137 (N_21137,N_19376,N_18064);
nor U21138 (N_21138,N_18497,N_16329);
and U21139 (N_21139,N_15872,N_15492);
or U21140 (N_21140,N_17213,N_17627);
nor U21141 (N_21141,N_19498,N_16672);
and U21142 (N_21142,N_18815,N_19673);
nand U21143 (N_21143,N_15806,N_19817);
nor U21144 (N_21144,N_17270,N_16534);
nand U21145 (N_21145,N_19751,N_18201);
or U21146 (N_21146,N_15982,N_16820);
or U21147 (N_21147,N_17022,N_19654);
xnor U21148 (N_21148,N_16740,N_19998);
xnor U21149 (N_21149,N_18262,N_15238);
nor U21150 (N_21150,N_19841,N_19658);
nor U21151 (N_21151,N_19078,N_19447);
nor U21152 (N_21152,N_16101,N_19319);
nor U21153 (N_21153,N_16256,N_17240);
nor U21154 (N_21154,N_16701,N_19334);
or U21155 (N_21155,N_16226,N_18479);
nand U21156 (N_21156,N_17911,N_15234);
or U21157 (N_21157,N_17968,N_16358);
nor U21158 (N_21158,N_19047,N_18425);
or U21159 (N_21159,N_19007,N_15377);
xnor U21160 (N_21160,N_19370,N_15288);
nand U21161 (N_21161,N_19577,N_16402);
nor U21162 (N_21162,N_17383,N_15161);
or U21163 (N_21163,N_17086,N_15886);
xor U21164 (N_21164,N_15180,N_19205);
or U21165 (N_21165,N_16035,N_17033);
nor U21166 (N_21166,N_19759,N_16496);
nand U21167 (N_21167,N_19087,N_15654);
nor U21168 (N_21168,N_16001,N_15256);
xor U21169 (N_21169,N_15679,N_17155);
nor U21170 (N_21170,N_19733,N_18383);
nand U21171 (N_21171,N_18658,N_18500);
or U21172 (N_21172,N_15507,N_19080);
or U21173 (N_21173,N_17051,N_18839);
nor U21174 (N_21174,N_19341,N_15120);
nand U21175 (N_21175,N_19312,N_19516);
or U21176 (N_21176,N_15151,N_18876);
or U21177 (N_21177,N_16636,N_19084);
or U21178 (N_21178,N_19215,N_16213);
xor U21179 (N_21179,N_16356,N_19198);
nor U21180 (N_21180,N_17800,N_19044);
or U21181 (N_21181,N_15865,N_18704);
nand U21182 (N_21182,N_15355,N_18372);
nand U21183 (N_21183,N_17374,N_15979);
xnor U21184 (N_21184,N_17526,N_15821);
nand U21185 (N_21185,N_15835,N_18898);
nand U21186 (N_21186,N_19993,N_16234);
nand U21187 (N_21187,N_16664,N_16851);
nand U21188 (N_21188,N_15193,N_18512);
or U21189 (N_21189,N_17017,N_18429);
nand U21190 (N_21190,N_16840,N_18483);
xor U21191 (N_21191,N_15462,N_19701);
nor U21192 (N_21192,N_16458,N_17958);
nor U21193 (N_21193,N_17205,N_17845);
and U21194 (N_21194,N_18768,N_17419);
and U21195 (N_21195,N_18605,N_15479);
nor U21196 (N_21196,N_17101,N_18299);
and U21197 (N_21197,N_17811,N_16656);
nor U21198 (N_21198,N_16350,N_16502);
nand U21199 (N_21199,N_19607,N_15347);
and U21200 (N_21200,N_17411,N_16768);
or U21201 (N_21201,N_19365,N_17495);
nor U21202 (N_21202,N_15525,N_17749);
and U21203 (N_21203,N_15825,N_16592);
xnor U21204 (N_21204,N_15233,N_19393);
or U21205 (N_21205,N_18347,N_19761);
or U21206 (N_21206,N_16538,N_16311);
nor U21207 (N_21207,N_15196,N_15221);
xnor U21208 (N_21208,N_16347,N_15959);
or U21209 (N_21209,N_18292,N_19014);
nand U21210 (N_21210,N_17317,N_15243);
nor U21211 (N_21211,N_19800,N_18333);
nor U21212 (N_21212,N_17569,N_15390);
or U21213 (N_21213,N_15070,N_15383);
or U21214 (N_21214,N_16175,N_18428);
and U21215 (N_21215,N_15904,N_15860);
and U21216 (N_21216,N_19233,N_15229);
nand U21217 (N_21217,N_18465,N_16238);
or U21218 (N_21218,N_17754,N_15692);
nor U21219 (N_21219,N_19193,N_17872);
nor U21220 (N_21220,N_15822,N_19017);
and U21221 (N_21221,N_19323,N_16961);
and U21222 (N_21222,N_15947,N_17492);
nand U21223 (N_21223,N_15893,N_17434);
and U21224 (N_21224,N_15643,N_18969);
and U21225 (N_21225,N_15459,N_17823);
nor U21226 (N_21226,N_16627,N_18154);
and U21227 (N_21227,N_17819,N_16543);
nand U21228 (N_21228,N_15089,N_16563);
nand U21229 (N_21229,N_19191,N_18323);
nand U21230 (N_21230,N_18853,N_15943);
or U21231 (N_21231,N_18907,N_19160);
or U21232 (N_21232,N_19838,N_15064);
or U21233 (N_21233,N_16086,N_16742);
or U21234 (N_21234,N_16660,N_18708);
and U21235 (N_21235,N_16454,N_16608);
and U21236 (N_21236,N_19355,N_17173);
nor U21237 (N_21237,N_16821,N_16266);
xor U21238 (N_21238,N_16239,N_18960);
nor U21239 (N_21239,N_18250,N_17295);
nor U21240 (N_21240,N_17178,N_18146);
nor U21241 (N_21241,N_17351,N_17353);
or U21242 (N_21242,N_16100,N_18709);
xor U21243 (N_21243,N_18461,N_18316);
and U21244 (N_21244,N_16072,N_19760);
and U21245 (N_21245,N_16044,N_19728);
nand U21246 (N_21246,N_15766,N_16360);
nand U21247 (N_21247,N_19110,N_16230);
or U21248 (N_21248,N_16455,N_19554);
nor U21249 (N_21249,N_18634,N_19121);
nand U21250 (N_21250,N_15778,N_19874);
xnor U21251 (N_21251,N_17562,N_16824);
nand U21252 (N_21252,N_16032,N_18775);
nand U21253 (N_21253,N_17757,N_16718);
and U21254 (N_21254,N_15079,N_15013);
and U21255 (N_21255,N_17002,N_16920);
nand U21256 (N_21256,N_18367,N_16591);
nor U21257 (N_21257,N_18285,N_16998);
or U21258 (N_21258,N_19639,N_18481);
nor U21259 (N_21259,N_15197,N_19989);
nor U21260 (N_21260,N_15047,N_18857);
or U21261 (N_21261,N_18606,N_15583);
and U21262 (N_21262,N_19286,N_17099);
or U21263 (N_21263,N_17779,N_17151);
and U21264 (N_21264,N_17445,N_18530);
and U21265 (N_21265,N_18424,N_17306);
or U21266 (N_21266,N_17284,N_19130);
xnor U21267 (N_21267,N_15075,N_18821);
or U21268 (N_21268,N_18349,N_16497);
nand U21269 (N_21269,N_16292,N_19234);
and U21270 (N_21270,N_15978,N_16003);
and U21271 (N_21271,N_16066,N_15090);
or U21272 (N_21272,N_17932,N_15940);
nor U21273 (N_21273,N_15025,N_15923);
and U21274 (N_21274,N_18152,N_15848);
nand U21275 (N_21275,N_18808,N_15810);
and U21276 (N_21276,N_17250,N_18697);
or U21277 (N_21277,N_18302,N_15164);
nand U21278 (N_21278,N_19194,N_15291);
or U21279 (N_21279,N_15205,N_19680);
nor U21280 (N_21280,N_15929,N_18503);
and U21281 (N_21281,N_18286,N_19204);
xor U21282 (N_21282,N_15937,N_15721);
nor U21283 (N_21283,N_16446,N_15324);
nor U21284 (N_21284,N_16545,N_19285);
or U21285 (N_21285,N_17176,N_16925);
or U21286 (N_21286,N_15416,N_16544);
or U21287 (N_21287,N_15039,N_19781);
or U21288 (N_21288,N_19065,N_17869);
or U21289 (N_21289,N_15504,N_15365);
and U21290 (N_21290,N_19707,N_16445);
or U21291 (N_21291,N_16848,N_19125);
or U21292 (N_21292,N_17018,N_17447);
xnor U21293 (N_21293,N_16521,N_15153);
or U21294 (N_21294,N_17430,N_19307);
nand U21295 (N_21295,N_15426,N_17391);
or U21296 (N_21296,N_17971,N_15014);
or U21297 (N_21297,N_19854,N_19045);
nor U21298 (N_21298,N_17577,N_16148);
nand U21299 (N_21299,N_16167,N_16468);
xor U21300 (N_21300,N_17804,N_15898);
and U21301 (N_21301,N_15046,N_18554);
nand U21302 (N_21302,N_18766,N_16166);
or U21303 (N_21303,N_18686,N_17116);
xnor U21304 (N_21304,N_18880,N_16432);
nand U21305 (N_21305,N_18317,N_18039);
nor U21306 (N_21306,N_15990,N_18555);
xor U21307 (N_21307,N_19146,N_18069);
and U21308 (N_21308,N_15103,N_19008);
nor U21309 (N_21309,N_18648,N_16703);
or U21310 (N_21310,N_16275,N_19003);
or U21311 (N_21311,N_18149,N_15334);
xor U21312 (N_21312,N_19932,N_17412);
nand U21313 (N_21313,N_18071,N_19734);
xnor U21314 (N_21314,N_15034,N_15635);
and U21315 (N_21315,N_19249,N_18546);
nand U21316 (N_21316,N_16320,N_15135);
or U21317 (N_21317,N_16807,N_18536);
and U21318 (N_21318,N_17441,N_18089);
nand U21319 (N_21319,N_18464,N_15790);
or U21320 (N_21320,N_19785,N_18488);
nand U21321 (N_21321,N_15107,N_18783);
or U21322 (N_21322,N_19027,N_15359);
nor U21323 (N_21323,N_16935,N_15337);
and U21324 (N_21324,N_15862,N_15647);
nand U21325 (N_21325,N_17900,N_15341);
nand U21326 (N_21326,N_18998,N_16140);
nand U21327 (N_21327,N_15091,N_16037);
nand U21328 (N_21328,N_15284,N_16228);
and U21329 (N_21329,N_16856,N_15311);
and U21330 (N_21330,N_19280,N_16973);
or U21331 (N_21331,N_19534,N_18370);
or U21332 (N_21332,N_15343,N_17115);
nand U21333 (N_21333,N_17835,N_17016);
and U21334 (N_21334,N_16698,N_19172);
or U21335 (N_21335,N_16749,N_18130);
and U21336 (N_21336,N_18160,N_19588);
xnor U21337 (N_21337,N_19559,N_16571);
xor U21338 (N_21338,N_17368,N_17686);
or U21339 (N_21339,N_18216,N_16747);
and U21340 (N_21340,N_16344,N_15160);
xnor U21341 (N_21341,N_16487,N_17019);
nand U21342 (N_21342,N_18918,N_18354);
or U21343 (N_21343,N_18520,N_19594);
or U21344 (N_21344,N_15441,N_15795);
nor U21345 (N_21345,N_19023,N_18169);
or U21346 (N_21346,N_18217,N_16744);
or U21347 (N_21347,N_18787,N_17036);
and U21348 (N_21348,N_16028,N_18080);
nand U21349 (N_21349,N_18128,N_19756);
nand U21350 (N_21350,N_18569,N_15309);
nand U21351 (N_21351,N_15967,N_15306);
and U21352 (N_21352,N_15513,N_15890);
or U21353 (N_21353,N_15261,N_18757);
xnor U21354 (N_21354,N_17282,N_16107);
nand U21355 (N_21355,N_15566,N_17665);
or U21356 (N_21356,N_18313,N_17497);
xor U21357 (N_21357,N_18514,N_15684);
or U21358 (N_21358,N_15784,N_19668);
nor U21359 (N_21359,N_15473,N_15364);
nor U21360 (N_21360,N_18233,N_16085);
or U21361 (N_21361,N_15127,N_18026);
or U21362 (N_21362,N_18540,N_18828);
nand U21363 (N_21363,N_16370,N_17784);
nor U21364 (N_21364,N_17862,N_18859);
nand U21365 (N_21365,N_17725,N_17407);
and U21366 (N_21366,N_15203,N_15073);
and U21367 (N_21367,N_16163,N_15147);
and U21368 (N_21368,N_18501,N_18967);
or U21369 (N_21369,N_17813,N_19768);
and U21370 (N_21370,N_17471,N_16799);
nand U21371 (N_21371,N_17519,N_17738);
or U21372 (N_21372,N_19965,N_15198);
and U21373 (N_21373,N_17465,N_18727);
nor U21374 (N_21374,N_19493,N_15735);
nand U21375 (N_21375,N_19753,N_16606);
or U21376 (N_21376,N_19455,N_16825);
and U21377 (N_21377,N_17287,N_18997);
nor U21378 (N_21378,N_15017,N_17965);
nor U21379 (N_21379,N_17673,N_18436);
and U21380 (N_21380,N_18862,N_19815);
or U21381 (N_21381,N_17132,N_17318);
and U21382 (N_21382,N_18438,N_15844);
or U21383 (N_21383,N_17755,N_19052);
and U21384 (N_21384,N_17762,N_16288);
nand U21385 (N_21385,N_17576,N_15842);
and U21386 (N_21386,N_15518,N_19424);
and U21387 (N_21387,N_17212,N_16859);
xor U21388 (N_21388,N_18101,N_17464);
nor U21389 (N_21389,N_19487,N_19515);
or U21390 (N_21390,N_15023,N_19336);
nor U21391 (N_21391,N_17795,N_15667);
nor U21392 (N_21392,N_16882,N_16395);
nor U21393 (N_21393,N_15826,N_17745);
and U21394 (N_21394,N_17628,N_17923);
nand U21395 (N_21395,N_16351,N_18038);
or U21396 (N_21396,N_16061,N_15701);
nand U21397 (N_21397,N_18414,N_15868);
and U21398 (N_21398,N_18418,N_19750);
and U21399 (N_21399,N_15078,N_17415);
xor U21400 (N_21400,N_18273,N_16863);
and U21401 (N_21401,N_17273,N_18729);
nand U21402 (N_21402,N_17632,N_15902);
nand U21403 (N_21403,N_17322,N_15915);
nand U21404 (N_21404,N_19479,N_17196);
nand U21405 (N_21405,N_15488,N_19593);
nand U21406 (N_21406,N_15640,N_15734);
and U21407 (N_21407,N_18129,N_16505);
nor U21408 (N_21408,N_15949,N_17590);
and U21409 (N_21409,N_17913,N_16542);
nor U21410 (N_21410,N_19656,N_16516);
and U21411 (N_21411,N_17625,N_19202);
and U21412 (N_21412,N_19822,N_19514);
or U21413 (N_21413,N_19116,N_17802);
nand U21414 (N_21414,N_17365,N_16363);
and U21415 (N_21415,N_19157,N_19809);
nand U21416 (N_21416,N_17788,N_17128);
nand U21417 (N_21417,N_19572,N_19871);
nor U21418 (N_21418,N_18549,N_19884);
or U21419 (N_21419,N_17935,N_17421);
xor U21420 (N_21420,N_16423,N_19892);
nand U21421 (N_21421,N_18328,N_15744);
nor U21422 (N_21422,N_19114,N_17425);
and U21423 (N_21423,N_18322,N_16796);
nand U21424 (N_21424,N_18975,N_16443);
nor U21425 (N_21425,N_15255,N_19000);
xnor U21426 (N_21426,N_15322,N_19968);
nand U21427 (N_21427,N_16811,N_17617);
nor U21428 (N_21428,N_16390,N_16194);
or U21429 (N_21429,N_16513,N_16928);
nor U21430 (N_21430,N_16854,N_17331);
nor U21431 (N_21431,N_15952,N_17107);
nand U21432 (N_21432,N_19139,N_19480);
or U21433 (N_21433,N_18407,N_19562);
nor U21434 (N_21434,N_19955,N_18563);
or U21435 (N_21435,N_18338,N_16581);
xor U21436 (N_21436,N_15746,N_16041);
and U21437 (N_21437,N_19421,N_19885);
or U21438 (N_21438,N_18629,N_19504);
or U21439 (N_21439,N_19459,N_16457);
nand U21440 (N_21440,N_15615,N_15211);
xor U21441 (N_21441,N_18027,N_18271);
or U21442 (N_21442,N_15106,N_18849);
nand U21443 (N_21443,N_19924,N_15114);
nor U21444 (N_21444,N_17925,N_18191);
xor U21445 (N_21445,N_16318,N_17692);
nor U21446 (N_21446,N_18389,N_15133);
nor U21447 (N_21447,N_16517,N_16948);
xor U21448 (N_21448,N_18011,N_16975);
or U21449 (N_21449,N_15214,N_18807);
xnor U21450 (N_21450,N_15273,N_17309);
or U21451 (N_21451,N_18593,N_16413);
or U21452 (N_21452,N_17886,N_17162);
and U21453 (N_21453,N_19523,N_18030);
and U21454 (N_21454,N_19006,N_15629);
xnor U21455 (N_21455,N_18221,N_16876);
and U21456 (N_21456,N_15710,N_17347);
nor U21457 (N_21457,N_16588,N_19565);
nand U21458 (N_21458,N_17093,N_16355);
or U21459 (N_21459,N_17090,N_18452);
or U21460 (N_21460,N_15590,N_17397);
and U21461 (N_21461,N_19943,N_18207);
and U21462 (N_21462,N_15839,N_18722);
or U21463 (N_21463,N_15171,N_17066);
nor U21464 (N_21464,N_16864,N_18478);
nor U21465 (N_21465,N_19778,N_17817);
xnor U21466 (N_21466,N_18779,N_17515);
and U21467 (N_21467,N_19613,N_16641);
nor U21468 (N_21468,N_17378,N_16960);
xnor U21469 (N_21469,N_19918,N_17121);
and U21470 (N_21470,N_16229,N_16684);
and U21471 (N_21471,N_15714,N_15344);
and U21472 (N_21472,N_15575,N_15379);
nand U21473 (N_21473,N_19717,N_17983);
nor U21474 (N_21474,N_18522,N_19267);
and U21475 (N_21475,N_19163,N_19173);
or U21476 (N_21476,N_15935,N_18619);
xor U21477 (N_21477,N_18735,N_16750);
nand U21478 (N_21478,N_17404,N_19740);
nor U21479 (N_21479,N_19923,N_16026);
nor U21480 (N_21480,N_15362,N_16006);
nor U21481 (N_21481,N_16971,N_19889);
and U21482 (N_21482,N_15065,N_16205);
nor U21483 (N_21483,N_19196,N_17075);
nand U21484 (N_21484,N_17901,N_17355);
and U21485 (N_21485,N_15564,N_16364);
nor U21486 (N_21486,N_19991,N_18833);
nor U21487 (N_21487,N_15188,N_17586);
nand U21488 (N_21488,N_18950,N_16800);
nor U21489 (N_21489,N_15074,N_16555);
nand U21490 (N_21490,N_17964,N_17186);
and U21491 (N_21491,N_15175,N_17294);
and U21492 (N_21492,N_16692,N_15457);
nor U21493 (N_21493,N_16585,N_18826);
or U21494 (N_21494,N_18022,N_17362);
or U21495 (N_21495,N_17679,N_19470);
nand U21496 (N_21496,N_15418,N_19938);
and U21497 (N_21497,N_15708,N_18303);
or U21498 (N_21498,N_18903,N_18060);
or U21499 (N_21499,N_18400,N_15606);
or U21500 (N_21500,N_19816,N_18580);
nand U21501 (N_21501,N_17766,N_15077);
or U21502 (N_21502,N_18020,N_16215);
or U21503 (N_21503,N_15116,N_19676);
nand U21504 (N_21504,N_15656,N_15108);
xor U21505 (N_21505,N_17100,N_15567);
nor U21506 (N_21506,N_17142,N_18145);
or U21507 (N_21507,N_19212,N_18212);
and U21508 (N_21508,N_17597,N_19076);
or U21509 (N_21509,N_15768,N_19450);
or U21510 (N_21510,N_15435,N_18294);
and U21511 (N_21511,N_17946,N_18635);
nand U21512 (N_21512,N_16812,N_18197);
nand U21513 (N_21513,N_16223,N_17301);
nor U21514 (N_21514,N_15568,N_18247);
or U21515 (N_21515,N_16295,N_16817);
nand U21516 (N_21516,N_19779,N_17004);
nor U21517 (N_21517,N_17328,N_17939);
or U21518 (N_21518,N_15006,N_16057);
and U21519 (N_21519,N_18163,N_16372);
and U21520 (N_21520,N_16916,N_18332);
and U21521 (N_21521,N_18804,N_18650);
nor U21522 (N_21522,N_17555,N_15569);
or U21523 (N_21523,N_15716,N_17691);
or U21524 (N_21524,N_16079,N_17281);
or U21525 (N_21525,N_16940,N_18192);
nor U21526 (N_21526,N_19082,N_15370);
nor U21527 (N_21527,N_17902,N_15172);
and U21528 (N_21528,N_16720,N_15984);
nand U21529 (N_21529,N_19449,N_18645);
and U21530 (N_21530,N_16688,N_16626);
and U21531 (N_21531,N_17781,N_15314);
and U21532 (N_21532,N_17422,N_17190);
xnor U21533 (N_21533,N_17768,N_17476);
or U21534 (N_21534,N_19399,N_17095);
nor U21535 (N_21535,N_15718,N_16654);
and U21536 (N_21536,N_15977,N_16869);
or U21537 (N_21537,N_19904,N_16986);
xor U21538 (N_21538,N_15143,N_15301);
nor U21539 (N_21539,N_17144,N_16659);
nand U21540 (N_21540,N_15316,N_15187);
or U21541 (N_21541,N_15972,N_15463);
or U21542 (N_21542,N_17489,N_15434);
nor U21543 (N_21543,N_17699,N_18987);
or U21544 (N_21544,N_18936,N_19576);
and U21545 (N_21545,N_17930,N_17263);
nand U21546 (N_21546,N_19230,N_15119);
nand U21547 (N_21547,N_17381,N_17225);
or U21548 (N_21548,N_17325,N_18926);
nand U21549 (N_21549,N_15033,N_15209);
nor U21550 (N_21550,N_19557,N_19629);
nor U21551 (N_21551,N_16227,N_16391);
nor U21552 (N_21552,N_17286,N_16280);
or U21553 (N_21553,N_17340,N_15757);
and U21554 (N_21554,N_19984,N_18872);
nor U21555 (N_21555,N_19445,N_17595);
nand U21556 (N_21556,N_19243,N_19035);
and U21557 (N_21557,N_18090,N_19140);
and U21558 (N_21558,N_17130,N_18682);
and U21559 (N_21559,N_19530,N_19066);
or U21560 (N_21560,N_15889,N_18371);
nor U21561 (N_21561,N_15038,N_15503);
xnor U21562 (N_21562,N_15137,N_15796);
nor U21563 (N_21563,N_19894,N_17783);
nor U21564 (N_21564,N_19408,N_19597);
and U21565 (N_21565,N_17432,N_17690);
nor U21566 (N_21566,N_17452,N_19807);
nor U21567 (N_21567,N_18057,N_16677);
nor U21568 (N_21568,N_17848,N_19939);
nor U21569 (N_21569,N_16658,N_17011);
and U21570 (N_21570,N_15407,N_16984);
and U21571 (N_21571,N_18009,N_18895);
nand U21572 (N_21572,N_19549,N_18981);
nand U21573 (N_21573,N_17437,N_17596);
and U21574 (N_21574,N_17337,N_15086);
nand U21575 (N_21575,N_19127,N_16842);
nand U21576 (N_21576,N_15397,N_18711);
xor U21577 (N_21577,N_18649,N_19279);
nand U21578 (N_21578,N_16373,N_18617);
nand U21579 (N_21579,N_18403,N_19454);
or U21580 (N_21580,N_16512,N_19974);
and U21581 (N_21581,N_17893,N_19154);
nor U21582 (N_21582,N_16785,N_17256);
and U21583 (N_21583,N_18234,N_17444);
and U21584 (N_21584,N_17433,N_16655);
nand U21585 (N_21585,N_19207,N_19912);
nand U21586 (N_21586,N_18793,N_18016);
or U21587 (N_21587,N_15932,N_18565);
nand U21588 (N_21588,N_19120,N_17927);
or U21589 (N_21589,N_16757,N_19603);
nor U21590 (N_21590,N_19325,N_18738);
or U21591 (N_21591,N_16794,N_19682);
nand U21592 (N_21592,N_15745,N_16477);
and U21593 (N_21593,N_17542,N_18342);
nor U21594 (N_21594,N_18877,N_15414);
or U21595 (N_21595,N_19387,N_18983);
and U21596 (N_21596,N_19780,N_15700);
or U21597 (N_21597,N_19050,N_19608);
or U21598 (N_21598,N_19743,N_17639);
nand U21599 (N_21599,N_19074,N_18989);
and U21600 (N_21600,N_16932,N_19070);
or U21601 (N_21601,N_17880,N_17995);
nor U21602 (N_21602,N_17604,N_16328);
xnor U21603 (N_21603,N_18088,N_15600);
or U21604 (N_21604,N_19022,N_18325);
xor U21605 (N_21605,N_19878,N_19713);
xnor U21606 (N_21606,N_17700,N_19311);
nand U21607 (N_21607,N_16727,N_15803);
nand U21608 (N_21608,N_16943,N_16736);
or U21609 (N_21609,N_18572,N_18666);
or U21610 (N_21610,N_19633,N_18355);
nor U21611 (N_21611,N_19273,N_18482);
nand U21612 (N_21612,N_19086,N_15593);
or U21613 (N_21613,N_17485,N_18976);
or U21614 (N_21614,N_16366,N_16498);
and U21615 (N_21615,N_16099,N_19466);
nand U21616 (N_21616,N_19596,N_15595);
or U21617 (N_21617,N_17744,N_17761);
and U21618 (N_21618,N_15818,N_17985);
and U21619 (N_21619,N_15997,N_19765);
and U21620 (N_21620,N_17797,N_17733);
nand U21621 (N_21621,N_18037,N_16198);
xnor U21622 (N_21622,N_15357,N_18035);
or U21623 (N_21623,N_15675,N_15149);
or U21624 (N_21624,N_19764,N_18607);
xnor U21625 (N_21625,N_17349,N_16104);
xnor U21626 (N_21626,N_15571,N_15944);
nand U21627 (N_21627,N_17390,N_15633);
nand U21628 (N_21628,N_18694,N_16151);
nand U21629 (N_21629,N_16015,N_19973);
or U21630 (N_21630,N_16010,N_19695);
xnor U21631 (N_21631,N_19692,N_15425);
nand U21632 (N_21632,N_19564,N_15042);
and U21633 (N_21633,N_19152,N_16293);
xnor U21634 (N_21634,N_18782,N_15548);
xor U21635 (N_21635,N_16359,N_19739);
nor U21636 (N_21636,N_16378,N_18213);
nor U21637 (N_21637,N_15174,N_17689);
nor U21638 (N_21638,N_15610,N_17740);
and U21639 (N_21639,N_16911,N_17537);
nand U21640 (N_21640,N_18810,N_15146);
nor U21641 (N_21641,N_15368,N_19598);
nor U21642 (N_21642,N_19221,N_19638);
or U21643 (N_21643,N_18719,N_18730);
nand U21644 (N_21644,N_17592,N_18240);
and U21645 (N_21645,N_16731,N_15850);
and U21646 (N_21646,N_19306,N_18553);
nand U21647 (N_21647,N_15405,N_18638);
or U21648 (N_21648,N_15587,N_16715);
nor U21649 (N_21649,N_15543,N_15906);
nand U21650 (N_21650,N_19061,N_18002);
nor U21651 (N_21651,N_16196,N_15431);
or U21652 (N_21652,N_16008,N_17764);
nand U21653 (N_21653,N_15495,N_19949);
or U21654 (N_21654,N_15410,N_18601);
nand U21655 (N_21655,N_19560,N_17849);
nor U21656 (N_21656,N_18091,N_19309);
nor U21657 (N_21657,N_17833,N_15447);
nor U21658 (N_21658,N_18610,N_15749);
and U21659 (N_21659,N_19720,N_15345);
nand U21660 (N_21660,N_18897,N_18538);
nor U21661 (N_21661,N_18948,N_17393);
nor U21662 (N_21662,N_15808,N_16334);
or U21663 (N_21663,N_17896,N_15134);
nor U21664 (N_21664,N_16904,N_16119);
nor U21665 (N_21665,N_17363,N_15231);
nand U21666 (N_21666,N_19582,N_15351);
xnor U21667 (N_21667,N_15423,N_19197);
or U21668 (N_21668,N_18175,N_15112);
xnor U21669 (N_21669,N_19891,N_19213);
or U21670 (N_21670,N_16424,N_17546);
xor U21671 (N_21671,N_16900,N_15727);
nor U21672 (N_21672,N_15529,N_17138);
nor U21673 (N_21673,N_19848,N_15814);
nand U21674 (N_21674,N_16559,N_17972);
nand U21675 (N_21675,N_19018,N_17621);
and U21676 (N_21676,N_15356,N_16019);
nor U21677 (N_21677,N_17940,N_19344);
nand U21678 (N_21678,N_15772,N_16201);
or U21679 (N_21679,N_18934,N_19610);
or U21680 (N_21680,N_19642,N_17726);
or U21681 (N_21681,N_18072,N_15634);
or U21682 (N_21682,N_17040,N_16144);
nand U21683 (N_21683,N_15573,N_18985);
and U21684 (N_21684,N_15514,N_17192);
nor U21685 (N_21685,N_17522,N_16603);
nand U21686 (N_21686,N_17416,N_17864);
nor U21687 (N_21687,N_17805,N_17063);
nand U21688 (N_21688,N_19009,N_16756);
and U21689 (N_21689,N_18687,N_18865);
xor U21690 (N_21690,N_18318,N_18858);
or U21691 (N_21691,N_19368,N_17561);
or U21692 (N_21692,N_18193,N_18248);
nor U21693 (N_21693,N_16068,N_17863);
nand U21694 (N_21694,N_18427,N_15037);
and U21695 (N_21695,N_15451,N_15580);
and U21696 (N_21696,N_16937,N_18558);
xor U21697 (N_21697,N_15620,N_19167);
or U21698 (N_21698,N_16263,N_17695);
nand U21699 (N_21699,N_19863,N_18576);
xor U21700 (N_21700,N_15823,N_18311);
nor U21701 (N_21701,N_18232,N_19546);
nand U21702 (N_21702,N_17064,N_16855);
or U21703 (N_21703,N_19389,N_19496);
nor U21704 (N_21704,N_18599,N_19405);
nor U21705 (N_21705,N_18237,N_17156);
nand U21706 (N_21706,N_18817,N_19624);
nand U21707 (N_21707,N_16946,N_19067);
nor U21708 (N_21708,N_17852,N_17837);
nor U21709 (N_21709,N_18786,N_18737);
nand U21710 (N_21710,N_18841,N_18937);
nor U21711 (N_21711,N_17891,N_18946);
or U21712 (N_21712,N_18251,N_16087);
nor U21713 (N_21713,N_19011,N_19278);
nand U21714 (N_21714,N_16927,N_19452);
nand U21715 (N_21715,N_16241,N_17087);
or U21716 (N_21716,N_19417,N_17941);
nor U21717 (N_21717,N_15671,N_15755);
nand U21718 (N_21718,N_17584,N_17798);
nand U21719 (N_21719,N_16628,N_19356);
nand U21720 (N_21720,N_18148,N_18051);
or U21721 (N_21721,N_18800,N_15852);
or U21722 (N_21722,N_16880,N_18151);
nand U21723 (N_21723,N_18208,N_17530);
nand U21724 (N_21724,N_19064,N_18015);
or U21725 (N_21725,N_15296,N_16539);
or U21726 (N_21726,N_19754,N_16005);
nor U21727 (N_21727,N_15328,N_18260);
or U21728 (N_21728,N_15373,N_18675);
nor U21729 (N_21729,N_17524,N_15877);
xor U21730 (N_21730,N_15326,N_18612);
nand U21731 (N_21731,N_16343,N_18725);
or U21732 (N_21732,N_17928,N_17599);
or U21733 (N_21733,N_17268,N_17209);
nand U21734 (N_21734,N_18469,N_18778);
nor U21735 (N_21735,N_18623,N_18269);
or U21736 (N_21736,N_16958,N_17044);
nand U21737 (N_21737,N_16442,N_19322);
xnor U21738 (N_21738,N_19337,N_19122);
or U21739 (N_21739,N_16251,N_15192);
and U21740 (N_21740,N_16849,N_16705);
nand U21741 (N_21741,N_16966,N_18571);
nor U21742 (N_21742,N_16501,N_18194);
nand U21743 (N_21743,N_16687,N_16783);
nor U21744 (N_21744,N_18124,N_18236);
xnor U21745 (N_21745,N_18045,N_16680);
and U21746 (N_21746,N_15638,N_17283);
and U21747 (N_21747,N_19731,N_18025);
nand U21748 (N_21748,N_16915,N_19569);
nor U21749 (N_21749,N_17356,N_16055);
xor U21750 (N_21750,N_16299,N_19649);
nand U21751 (N_21751,N_16723,N_18331);
and U21752 (N_21752,N_15691,N_19206);
and U21753 (N_21753,N_16959,N_15743);
nand U21754 (N_21754,N_15438,N_16425);
and U21755 (N_21755,N_16452,N_17248);
or U21756 (N_21756,N_17648,N_18882);
nand U21757 (N_21757,N_15494,N_19201);
xor U21758 (N_21758,N_17966,N_15335);
and U21759 (N_21759,N_19897,N_15456);
and U21760 (N_21760,N_17076,N_18566);
nand U21761 (N_21761,N_19820,N_17943);
nor U21762 (N_21762,N_18670,N_16890);
or U21763 (N_21763,N_17516,N_17602);
nand U21764 (N_21764,N_15816,N_17587);
xnor U21765 (N_21765,N_19349,N_16050);
nor U21766 (N_21766,N_15592,N_15510);
nand U21767 (N_21767,N_16686,N_16392);
nand U21768 (N_21768,N_16376,N_17307);
xnor U21769 (N_21769,N_19958,N_16016);
or U21770 (N_21770,N_16629,N_18893);
nor U21771 (N_21771,N_15249,N_17252);
nand U21772 (N_21772,N_15170,N_18953);
nor U21773 (N_21773,N_19964,N_19521);
or U21774 (N_21774,N_15907,N_15139);
nand U21775 (N_21775,N_18472,N_18108);
and U21776 (N_21776,N_18680,N_15761);
and U21777 (N_21777,N_18700,N_15472);
or U21778 (N_21778,N_17961,N_19722);
nand U21779 (N_21779,N_15552,N_15512);
xnor U21780 (N_21780,N_19540,N_15641);
or U21781 (N_21781,N_16509,N_19663);
xnor U21782 (N_21782,N_15179,N_16412);
or U21783 (N_21783,N_16297,N_18373);
xnor U21784 (N_21784,N_18227,N_18943);
nand U21785 (N_21785,N_16898,N_16721);
or U21786 (N_21786,N_18416,N_18891);
or U21787 (N_21787,N_16269,N_18736);
nand U21788 (N_21788,N_19689,N_17853);
or U21789 (N_21789,N_16870,N_17909);
nand U21790 (N_21790,N_18699,N_15126);
or U21791 (N_21791,N_15787,N_18798);
and U21792 (N_21792,N_16872,N_15226);
or U21793 (N_21793,N_16374,N_17682);
or U21794 (N_21794,N_16587,N_15802);
and U21795 (N_21795,N_19320,N_17236);
and U21796 (N_21796,N_19096,N_18398);
nand U21797 (N_21797,N_17549,N_18343);
nor U21798 (N_21798,N_16944,N_19960);
nand U21799 (N_21799,N_16643,N_16138);
or U21800 (N_21800,N_18239,N_16739);
nand U21801 (N_21801,N_15799,N_15399);
and U21802 (N_21802,N_15644,N_19641);
or U21803 (N_21803,N_19846,N_17559);
and U21804 (N_21804,N_15307,N_18801);
nor U21805 (N_21805,N_17377,N_17131);
nand U21806 (N_21806,N_17005,N_18785);
and U21807 (N_21807,N_18923,N_17566);
and U21808 (N_21808,N_16472,N_15939);
nor U21809 (N_21809,N_16252,N_15021);
or U21810 (N_21810,N_18613,N_19131);
nor U21811 (N_21811,N_18086,N_16422);
and U21812 (N_21812,N_18683,N_16048);
and U21813 (N_21813,N_15777,N_17658);
or U21814 (N_21814,N_18382,N_16380);
and U21815 (N_21815,N_15742,N_15500);
nand U21816 (N_21816,N_16938,N_15439);
and U21817 (N_21817,N_15449,N_15110);
or U21818 (N_21818,N_18492,N_16254);
or U21819 (N_21819,N_15836,N_17401);
nor U21820 (N_21820,N_19819,N_16332);
and U21821 (N_21821,N_19630,N_19460);
and U21822 (N_21822,N_17701,N_19265);
nand U21823 (N_21823,N_16939,N_17707);
and U21824 (N_21824,N_19224,N_17616);
nor U21825 (N_21825,N_18723,N_15921);
nand U21826 (N_21826,N_16781,N_16369);
nor U21827 (N_21827,N_16271,N_17550);
xor U21828 (N_21828,N_15841,N_16858);
nor U21829 (N_21829,N_18195,N_16386);
and U21830 (N_21830,N_19046,N_17578);
nor U21831 (N_21831,N_18264,N_16272);
nand U21832 (N_21832,N_15223,N_16092);
nand U21833 (N_21833,N_15832,N_18385);
and U21834 (N_21834,N_18456,N_18295);
and U21835 (N_21835,N_18614,N_15453);
and U21836 (N_21836,N_16298,N_19256);
xor U21837 (N_21837,N_16634,N_18545);
and U21838 (N_21838,N_18548,N_16210);
and U21839 (N_21839,N_16648,N_16530);
nand U21840 (N_21840,N_15254,N_15542);
or U21841 (N_21841,N_16123,N_15598);
nor U21842 (N_21842,N_15406,N_19461);
xnor U21843 (N_21843,N_16170,N_18033);
and U21844 (N_21844,N_16038,N_18329);
nor U21845 (N_21845,N_15310,N_17693);
or U21846 (N_21846,N_17696,N_15505);
nand U21847 (N_21847,N_15101,N_16012);
xnor U21848 (N_21848,N_15657,N_17292);
nor U21849 (N_21849,N_15834,N_17237);
nor U21850 (N_21850,N_16062,N_18280);
and U21851 (N_21851,N_18902,N_18971);
xor U21852 (N_21852,N_18258,N_19950);
and U21853 (N_21853,N_16801,N_17185);
xnor U21854 (N_21854,N_16584,N_18181);
and U21855 (N_21855,N_16888,N_19928);
and U21856 (N_21856,N_15707,N_17712);
xor U21857 (N_21857,N_16209,N_18832);
and U21858 (N_21858,N_17899,N_18972);
nor U21859 (N_21859,N_16098,N_17759);
nor U21860 (N_21860,N_19568,N_15270);
nand U21861 (N_21861,N_15720,N_18087);
nand U21862 (N_21862,N_15616,N_19448);
xnor U21863 (N_21863,N_16179,N_15891);
nor U21864 (N_21864,N_18369,N_17591);
nand U21865 (N_21865,N_18931,N_16249);
and U21866 (N_21866,N_15285,N_15539);
or U21867 (N_21867,N_15413,N_17791);
nor U21868 (N_21868,N_16575,N_18847);
nand U21869 (N_21869,N_16353,N_16105);
xor U21870 (N_21870,N_16891,N_15752);
and U21871 (N_21871,N_15317,N_19209);
nor U21872 (N_21872,N_19813,N_16798);
and U21873 (N_21873,N_17122,N_17161);
and U21874 (N_21874,N_19364,N_16901);
or U21875 (N_21875,N_18515,N_17110);
and U21876 (N_21876,N_19155,N_19675);
and U21877 (N_21877,N_16301,N_15673);
nor U21878 (N_21878,N_19353,N_16214);
xnor U21879 (N_21879,N_15085,N_18861);
nor U21880 (N_21880,N_17371,N_15105);
or U21881 (N_21881,N_18321,N_18657);
nand U21882 (N_21882,N_18945,N_16802);
and U21883 (N_21883,N_18107,N_16489);
and U21884 (N_21884,N_15391,N_19028);
nand U21885 (N_21885,N_18792,N_17238);
nor U21886 (N_21886,N_19953,N_17398);
nor U21887 (N_21887,N_17685,N_18485);
nor U21888 (N_21888,N_16371,N_16470);
and U21889 (N_21889,N_19227,N_16847);
nand U21890 (N_21890,N_19636,N_15372);
nor U21891 (N_21891,N_19440,N_15925);
nor U21892 (N_21892,N_18021,N_19438);
or U21893 (N_21893,N_17773,N_17302);
and U21894 (N_21894,N_16208,N_15173);
and U21895 (N_21895,N_16953,N_15585);
and U21896 (N_21896,N_19282,N_16693);
xnor U21897 (N_21897,N_15874,N_16022);
and U21898 (N_21898,N_17229,N_18733);
or U21899 (N_21899,N_17235,N_15546);
nand U21900 (N_21900,N_16691,N_18209);
nor U21901 (N_21901,N_15682,N_19839);
and U21902 (N_21902,N_18348,N_16881);
or U21903 (N_21903,N_18466,N_15384);
nand U21904 (N_21904,N_16792,N_19214);
nor U21905 (N_21905,N_17070,N_19332);
nand U21906 (N_21906,N_19143,N_16637);
nand U21907 (N_21907,N_16411,N_16793);
or U21908 (N_21908,N_19055,N_18447);
and U21909 (N_21909,N_15176,N_18123);
nand U21910 (N_21910,N_16436,N_16157);
or U21911 (N_21911,N_17780,N_18993);
nor U21912 (N_21912,N_15917,N_18177);
nor U21913 (N_21913,N_16419,N_15623);
and U21914 (N_21914,N_17496,N_19247);
xnor U21915 (N_21915,N_16507,N_16618);
xnor U21916 (N_21916,N_19893,N_18958);
nor U21917 (N_21917,N_16430,N_15601);
nand U21918 (N_21918,N_19261,N_15712);
and U21919 (N_21919,N_18894,N_17440);
nor U21920 (N_21920,N_17152,N_17245);
or U21921 (N_21921,N_17409,N_17198);
and U21922 (N_21922,N_16741,N_18388);
or U21923 (N_21923,N_18135,N_17165);
nand U21924 (N_21924,N_18266,N_18661);
nor U21925 (N_21925,N_16169,N_19749);
nand U21926 (N_21926,N_16473,N_19257);
or U21927 (N_21927,N_19416,N_15050);
and U21928 (N_21928,N_17753,N_15690);
nor U21929 (N_21929,N_17885,N_17636);
nor U21930 (N_21930,N_15036,N_15470);
and U21931 (N_21931,N_17903,N_15866);
nand U21932 (N_21932,N_19324,N_16493);
nor U21933 (N_21933,N_15111,N_19260);
nand U21934 (N_21934,N_16218,N_15058);
and U21935 (N_21935,N_19862,N_15551);
or U21936 (N_21936,N_19051,N_16866);
and U21937 (N_21937,N_19653,N_17521);
nand U21938 (N_21938,N_18306,N_19972);
nand U21939 (N_21939,N_16771,N_18141);
or U21940 (N_21940,N_18819,N_19093);
or U21941 (N_21941,N_16492,N_19703);
or U21942 (N_21942,N_16319,N_15055);
and U21943 (N_21943,N_15227,N_19177);
nand U21944 (N_21944,N_18731,N_19507);
nor U21945 (N_21945,N_19439,N_19442);
and U21946 (N_21946,N_18556,N_17624);
nand U21947 (N_21947,N_18063,N_19948);
nand U21948 (N_21948,N_15138,N_18242);
nor U21949 (N_21949,N_17919,N_19566);
or U21950 (N_21950,N_19425,N_16231);
or U21951 (N_21951,N_16387,N_17184);
nand U21952 (N_21952,N_18834,N_15474);
or U21953 (N_21953,N_18162,N_17369);
nand U21954 (N_21954,N_19644,N_19555);
or U21955 (N_21955,N_19156,N_19188);
nand U21956 (N_21956,N_16675,N_18358);
or U21957 (N_21957,N_17008,N_16270);
nand U21958 (N_21958,N_17215,N_17395);
and U21959 (N_21959,N_15247,N_17423);
nor U21960 (N_21960,N_16069,N_15297);
or U21961 (N_21961,N_17082,N_19810);
nor U21962 (N_21962,N_16719,N_16965);
nand U21963 (N_21963,N_15733,N_16460);
nand U21964 (N_21964,N_17705,N_18618);
or U21965 (N_21965,N_18525,N_17414);
xor U21966 (N_21966,N_18869,N_18767);
nor U21967 (N_21967,N_16936,N_15382);
nor U21968 (N_21968,N_15697,N_19388);
nand U21969 (N_21969,N_16287,N_17364);
or U21970 (N_21970,N_18377,N_15275);
nand U21971 (N_21971,N_16712,N_15093);
or U21972 (N_21972,N_18822,N_15581);
nand U21973 (N_21973,N_16652,N_15942);
and U21974 (N_21974,N_19536,N_19170);
and U21975 (N_21975,N_16441,N_18246);
xnor U21976 (N_21976,N_17074,N_19426);
or U21977 (N_21977,N_17633,N_17644);
nor U21978 (N_21978,N_17061,N_16767);
nor U21979 (N_21979,N_15555,N_19988);
and U21980 (N_21980,N_19947,N_16481);
and U21981 (N_21981,N_18166,N_19294);
nand U21982 (N_21982,N_15339,N_17310);
nand U21983 (N_21983,N_19705,N_19266);
and U21984 (N_21984,N_17336,N_17361);
nand U21985 (N_21985,N_18157,N_18127);
nand U21986 (N_21986,N_15168,N_16830);
or U21987 (N_21987,N_19095,N_17910);
or U21988 (N_21988,N_18740,N_19620);
and U21989 (N_21989,N_15348,N_15831);
or U21990 (N_21990,N_16996,N_17671);
nor U21991 (N_21991,N_19667,N_16694);
nand U21992 (N_21992,N_18006,N_19404);
or U21993 (N_21993,N_18688,N_15685);
nand U21994 (N_21994,N_18187,N_18908);
nand U21995 (N_21995,N_17723,N_18231);
nand U21996 (N_21996,N_17230,N_16639);
nor U21997 (N_21997,N_19400,N_18979);
or U21998 (N_21998,N_19486,N_15968);
nor U21999 (N_21999,N_17202,N_15537);
nor U22000 (N_22000,N_18344,N_17605);
xor U22001 (N_22001,N_16216,N_15152);
xnor U22002 (N_22002,N_18636,N_19036);
nand U22003 (N_22003,N_18445,N_19853);
or U22004 (N_22004,N_17517,N_19664);
nor U22005 (N_22005,N_17366,N_18133);
nor U22006 (N_22006,N_18746,N_18056);
or U22007 (N_22007,N_16503,N_19601);
and U22008 (N_22008,N_19648,N_18860);
and U22009 (N_22009,N_16461,N_17736);
or U22010 (N_22010,N_18085,N_15264);
and U22011 (N_22011,N_15294,N_16296);
or U22012 (N_22012,N_17743,N_16500);
nor U22013 (N_22013,N_16410,N_16653);
and U22014 (N_22014,N_16816,N_17207);
xor U22015 (N_22015,N_16180,N_15793);
or U22016 (N_22016,N_17719,N_16448);
or U22017 (N_22017,N_17262,N_18714);
xnor U22018 (N_22018,N_15040,N_15122);
nor U22019 (N_22019,N_16670,N_18899);
nor U22020 (N_22020,N_16595,N_16097);
nand U22021 (N_22021,N_17352,N_19573);
nor U22022 (N_22022,N_16862,N_15999);
or U22023 (N_22023,N_16197,N_19429);
xor U22024 (N_22024,N_15516,N_15004);
nor U22025 (N_22025,N_19737,N_19316);
or U22026 (N_22026,N_16941,N_16154);
or U22027 (N_22027,N_17242,N_15948);
nand U22028 (N_22028,N_17844,N_15509);
nor U22029 (N_22029,N_19963,N_18446);
and U22030 (N_22030,N_18109,N_16049);
xor U22031 (N_22031,N_16406,N_15446);
or U22032 (N_22032,N_15131,N_17001);
nand U22033 (N_22033,N_16846,N_19492);
nand U22034 (N_22034,N_17259,N_17957);
nand U22035 (N_22035,N_15597,N_17668);
nand U22036 (N_22036,N_16339,N_16537);
xnor U22037 (N_22037,N_19276,N_19691);
and U22038 (N_22038,N_18781,N_18668);
or U22039 (N_22039,N_16471,N_16438);
nor U22040 (N_22040,N_18836,N_15163);
nand U22041 (N_22041,N_15469,N_17851);
and U22042 (N_22042,N_15983,N_19446);
nor U22043 (N_22043,N_15320,N_17529);
nor U22044 (N_22044,N_19804,N_17934);
or U22045 (N_22045,N_17386,N_18760);
nand U22046 (N_22046,N_18032,N_18010);
and U22047 (N_22047,N_17081,N_19544);
xnor U22048 (N_22048,N_16011,N_16276);
or U22049 (N_22049,N_17103,N_18973);
and U22050 (N_22050,N_15791,N_19174);
nand U22051 (N_22051,N_15969,N_15630);
and U22052 (N_22052,N_19746,N_15315);
nor U22053 (N_22053,N_19145,N_15354);
nand U22054 (N_22054,N_18432,N_18223);
nor U22055 (N_22055,N_17493,N_18410);
nand U22056 (N_22056,N_17640,N_17806);
nor U22057 (N_22057,N_19477,N_18179);
or U22058 (N_22058,N_15010,N_18336);
or U22059 (N_22059,N_19709,N_15878);
xnor U22060 (N_22060,N_17763,N_18412);
and U22061 (N_22061,N_17629,N_19119);
or U22062 (N_22062,N_15669,N_15241);
nor U22063 (N_22063,N_16111,N_17883);
xor U22064 (N_22064,N_19926,N_18140);
nor U22065 (N_22065,N_17507,N_19420);
and U22066 (N_22066,N_17620,N_19072);
nor U22067 (N_22067,N_19626,N_15894);
nand U22068 (N_22068,N_18253,N_19777);
nor U22069 (N_22069,N_18214,N_16995);
nor U22070 (N_22070,N_16007,N_19381);
and U22071 (N_22071,N_16758,N_17167);
nor U22072 (N_22072,N_18337,N_17950);
nand U22073 (N_22073,N_15798,N_17139);
nand U22074 (N_22074,N_19277,N_19832);
nand U22075 (N_22075,N_17790,N_18041);
or U22076 (N_22076,N_15888,N_17164);
or U22077 (N_22077,N_16070,N_19343);
nor U22078 (N_22078,N_16607,N_16240);
or U22079 (N_22079,N_16222,N_19527);
nor U22080 (N_22080,N_19350,N_17410);
nor U22081 (N_22081,N_17413,N_17553);
nand U22082 (N_22082,N_18916,N_17793);
nor U22083 (N_22083,N_19012,N_18334);
nand U22084 (N_22084,N_15863,N_15224);
nand U22085 (N_22085,N_18244,N_15651);
and U22086 (N_22086,N_18842,N_16729);
nand U22087 (N_22087,N_17808,N_18712);
nor U22088 (N_22088,N_18230,N_15007);
or U22089 (N_22089,N_16336,N_18692);
or U22090 (N_22090,N_15366,N_19289);
xor U22091 (N_22091,N_19136,N_15864);
nor U22092 (N_22092,N_19288,N_15602);
and U22093 (N_22093,N_15558,N_15204);
nand U22094 (N_22094,N_16279,N_15655);
and U22095 (N_22095,N_18921,N_19837);
and U22096 (N_22096,N_18390,N_15591);
xor U22097 (N_22097,N_17455,N_19702);
or U22098 (N_22098,N_18024,N_17048);
or U22099 (N_22099,N_16748,N_15563);
nand U22100 (N_22100,N_18283,N_19432);
or U22101 (N_22101,N_15632,N_16161);
nand U22102 (N_22102,N_15195,N_18034);
nor U22103 (N_22103,N_18560,N_16957);
nor U22104 (N_22104,N_18112,N_18486);
and U22105 (N_22105,N_15763,N_15486);
nand U22106 (N_22106,N_19473,N_19409);
and U22107 (N_22107,N_17239,N_16844);
or U22108 (N_22108,N_15144,N_16931);
nand U22109 (N_22109,N_18049,N_15022);
or U22110 (N_22110,N_16556,N_16315);
and U22111 (N_22111,N_19829,N_18259);
and U22112 (N_22112,N_15465,N_18659);
and U22113 (N_22113,N_19317,N_18550);
nand U22114 (N_22114,N_16635,N_17672);
and U22115 (N_22115,N_19340,N_17285);
or U22116 (N_22116,N_16945,N_15588);
or U22117 (N_22117,N_15794,N_17073);
nand U22118 (N_22118,N_15084,N_19293);
and U22119 (N_22119,N_15097,N_15689);
nor U22120 (N_22120,N_16305,N_15092);
or U22121 (N_22121,N_16805,N_18099);
and U22122 (N_22122,N_16617,N_17201);
or U22123 (N_22123,N_17191,N_18886);
or U22124 (N_22124,N_16523,N_18366);
or U22125 (N_22125,N_15001,N_15626);
nand U22126 (N_22126,N_18084,N_18048);
nor U22127 (N_22127,N_15295,N_17816);
nor U22128 (N_22128,N_16642,N_16433);
xnor U22129 (N_22129,N_17931,N_15895);
or U22130 (N_22130,N_16657,N_18611);
or U22131 (N_22131,N_19412,N_16734);
nand U22132 (N_22132,N_19700,N_15699);
or U22133 (N_22133,N_16348,N_17840);
or U22134 (N_22134,N_17141,N_18710);
nor U22135 (N_22135,N_18004,N_17916);
and U22136 (N_22136,N_15338,N_17513);
and U22137 (N_22137,N_19431,N_17104);
and U22138 (N_22138,N_19788,N_15913);
and U22139 (N_22139,N_18587,N_15985);
nand U22140 (N_22140,N_15553,N_19600);
nand U22141 (N_22141,N_16185,N_19925);
and U22142 (N_22142,N_15286,N_18672);
nand U22143 (N_22143,N_16103,N_15964);
or U22144 (N_22144,N_15751,N_19541);
or U22145 (N_22145,N_16667,N_19900);
nor U22146 (N_22146,N_19335,N_16377);
and U22147 (N_22147,N_17180,N_15614);
nor U22148 (N_22148,N_16009,N_18017);
or U22149 (N_22149,N_15268,N_19327);
nor U22150 (N_22150,N_17539,N_18304);
nor U22151 (N_22151,N_15128,N_17246);
xor U22152 (N_22152,N_16773,N_18749);
and U22153 (N_22153,N_19383,N_17510);
or U22154 (N_22154,N_19579,N_19300);
nor U22155 (N_22155,N_19790,N_15124);
or U22156 (N_22156,N_17269,N_16303);
nor U22157 (N_22157,N_19190,N_16018);
or U22158 (N_22158,N_19434,N_18094);
nand U22159 (N_22159,N_15931,N_18598);
nand U22160 (N_22160,N_16676,N_16551);
nor U22161 (N_22161,N_18404,N_16875);
or U22162 (N_22162,N_15995,N_15374);
nor U22163 (N_22163,N_18356,N_16562);
and U22164 (N_22164,N_17096,N_19835);
xnor U22165 (N_22165,N_15183,N_19451);
and U22166 (N_22166,N_17234,N_19558);
nor U22167 (N_22167,N_16396,N_18551);
or U22168 (N_22168,N_17170,N_16633);
nand U22169 (N_22169,N_15454,N_19025);
nand U22170 (N_22170,N_15811,N_18747);
and U22171 (N_22171,N_17330,N_16907);
nor U22172 (N_22172,N_15589,N_18621);
and U22173 (N_22173,N_16689,N_17068);
and U22174 (N_22174,N_15319,N_17856);
or U22175 (N_22175,N_16910,N_18384);
or U22176 (N_22176,N_16769,N_17145);
nor U22177 (N_22177,N_17588,N_18954);
and U22178 (N_22178,N_18951,N_15577);
or U22179 (N_22179,N_18220,N_16220);
xnor U22180 (N_22180,N_18974,N_16340);
nand U22181 (N_22181,N_19099,N_19363);
or U22182 (N_22182,N_15329,N_17907);
and U22183 (N_22183,N_18473,N_16398);
or U22184 (N_22184,N_19699,N_18748);
nand U22185 (N_22185,N_15901,N_17014);
nand U22186 (N_22186,N_19369,N_15031);
or U22187 (N_22187,N_18589,N_16893);
nor U22188 (N_22188,N_18113,N_19180);
and U22189 (N_22189,N_15252,N_18136);
or U22190 (N_22190,N_15717,N_17426);
or U22191 (N_22191,N_18170,N_15765);
and U22192 (N_22192,N_15540,N_18159);
or U22193 (N_22193,N_18991,N_19635);
and U22194 (N_22194,N_16043,N_19940);
nand U22195 (N_22195,N_18320,N_19789);
xor U22196 (N_22196,N_16569,N_19830);
xnor U22197 (N_22197,N_18927,N_19101);
nand U22198 (N_22198,N_15083,N_18944);
nand U22199 (N_22199,N_16462,N_17135);
nand U22200 (N_22200,N_18681,N_17716);
nor U22201 (N_22201,N_18646,N_15464);
nor U22202 (N_22202,N_19229,N_19921);
or U22203 (N_22203,N_17825,N_16160);
or U22204 (N_22204,N_18078,N_15960);
or U22205 (N_22205,N_19617,N_18204);
or U22206 (N_22206,N_18999,N_15624);
nand U22207 (N_22207,N_18315,N_17030);
xor U22208 (N_22208,N_15421,N_17013);
nor U22209 (N_22209,N_19043,N_18794);
nor U22210 (N_22210,N_19467,N_17989);
nor U22211 (N_22211,N_17877,N_16029);
or U22212 (N_22212,N_18393,N_16540);
nand U22213 (N_22213,N_16557,N_15559);
nand U22214 (N_22214,N_15554,N_16058);
and U22215 (N_22215,N_18516,N_18058);
nor U22216 (N_22216,N_16730,N_19296);
and U22217 (N_22217,N_18691,N_17372);
and U22218 (N_22218,N_18065,N_17657);
nor U22219 (N_22219,N_19805,N_19704);
or U22220 (N_22220,N_15181,N_17912);
nand U22221 (N_22221,N_16933,N_15534);
or U22222 (N_22222,N_15222,N_16264);
nand U22223 (N_22223,N_17296,N_15958);
and U22224 (N_22224,N_19581,N_16696);
and U22225 (N_22225,N_18509,N_18144);
nand U22226 (N_22226,N_18996,N_18105);
or U22227 (N_22227,N_15650,N_19729);
xnor U22228 (N_22228,N_18932,N_16532);
nand U22229 (N_22229,N_16612,N_18138);
or U22230 (N_22230,N_16685,N_15220);
nand U22231 (N_22231,N_19782,N_15683);
nand U22232 (N_22232,N_18359,N_16708);
and U22233 (N_22233,N_17782,N_15672);
or U22234 (N_22234,N_18326,N_15068);
nand U22235 (N_22235,N_16002,N_18887);
or U22236 (N_22236,N_18289,N_16491);
nor U22237 (N_22237,N_17015,N_19220);
and U22238 (N_22238,N_17970,N_16576);
or U22239 (N_22239,N_19199,N_16791);
nor U22240 (N_22240,N_19678,N_17870);
or U22241 (N_22241,N_18119,N_19238);
xor U22242 (N_22242,N_17080,N_17981);
or U22243 (N_22243,N_15276,N_17615);
or U22244 (N_22244,N_19571,N_17563);
or U22245 (N_22245,N_17548,N_19909);
nor U22246 (N_22246,N_19512,N_17778);
nand U22247 (N_22247,N_17149,N_15427);
or U22248 (N_22248,N_17826,N_19465);
and U22249 (N_22249,N_15920,N_16510);
and U22250 (N_22250,N_17462,N_16128);
or U22251 (N_22251,N_18252,N_15190);
or U22252 (N_22252,N_15385,N_19758);
nand U22253 (N_22253,N_16117,N_17313);
nor U22254 (N_22254,N_15444,N_18276);
or U22255 (N_22255,N_18396,N_15732);
nor U22256 (N_22256,N_18186,N_17647);
nand U22257 (N_22257,N_19033,N_19137);
nor U22258 (N_22258,N_19258,N_18487);
nor U22259 (N_22259,N_17818,N_16942);
nor U22260 (N_22260,N_17674,N_19437);
and U22261 (N_22261,N_16084,N_18463);
nor U22262 (N_22262,N_16314,N_17760);
nor U22263 (N_22263,N_18665,N_18183);
nand U22264 (N_22264,N_17126,N_19796);
and U22265 (N_22265,N_16267,N_15980);
xnor U22266 (N_22266,N_19104,N_16964);
xor U22267 (N_22267,N_17888,N_15266);
nor U22268 (N_22268,N_16709,N_15549);
or U22269 (N_22269,N_17905,N_19619);
nand U22270 (N_22270,N_17894,N_18451);
and U22271 (N_22271,N_16528,N_17065);
and U22272 (N_22272,N_16601,N_15998);
and U22273 (N_22273,N_18171,N_19123);
nor U22274 (N_22274,N_17039,N_17991);
and U22275 (N_22275,N_16520,N_17541);
or U22276 (N_22276,N_16706,N_16023);
or U22277 (N_22277,N_19914,N_19144);
or U22278 (N_22278,N_15242,N_19575);
xor U22279 (N_22279,N_16245,N_19808);
nand U22280 (N_22280,N_19942,N_18875);
nand U22281 (N_22281,N_17684,N_17812);
nand U22282 (N_22282,N_19937,N_15668);
and U22283 (N_22283,N_16809,N_19683);
nand U22284 (N_22284,N_18378,N_17405);
or U22285 (N_22285,N_19444,N_15282);
or U22286 (N_22286,N_16988,N_15186);
nand U22287 (N_22287,N_18053,N_15628);
nand U22288 (N_22288,N_18624,N_17583);
and U22289 (N_22289,N_19295,N_16999);
and U22290 (N_22290,N_17859,N_16843);
nor U22291 (N_22291,N_19456,N_15781);
xnor U22292 (N_22292,N_15843,N_15461);
xnor U22293 (N_22293,N_18282,N_18816);
nor U22294 (N_22294,N_18626,N_19430);
and U22295 (N_22295,N_16149,N_16732);
or U22296 (N_22296,N_17676,N_17456);
or U22297 (N_22297,N_17214,N_17461);
or U22298 (N_22298,N_17029,N_19712);
nand U22299 (N_22299,N_18054,N_19647);
nand U22300 (N_22300,N_16884,N_17153);
and U22301 (N_22301,N_18224,N_19411);
nand U22302 (N_22302,N_19135,N_17370);
and U22303 (N_22303,N_16806,N_19814);
and U22304 (N_22304,N_18102,N_17473);
and U22305 (N_22305,N_19218,N_18467);
nor U22306 (N_22306,N_16894,N_17373);
and U22307 (N_22307,N_16533,N_17315);
or U22308 (N_22308,N_18759,N_15858);
nor U22309 (N_22309,N_17032,N_15376);
nor U22310 (N_22310,N_19519,N_15398);
and U22311 (N_22311,N_17735,N_15145);
nand U22312 (N_22312,N_19694,N_15015);
and U22313 (N_22313,N_15218,N_19812);
nor U22314 (N_22314,N_15278,N_18594);
nor U22315 (N_22315,N_16651,N_17751);
nor U22316 (N_22316,N_17654,N_17226);
nand U22317 (N_22317,N_17895,N_17533);
nor U22318 (N_22318,N_19248,N_15956);
nor U22319 (N_22319,N_15201,N_17298);
and U22320 (N_22320,N_16152,N_16711);
xnor U22321 (N_22321,N_18743,N_16886);
nor U22322 (N_22322,N_19933,N_19488);
nor U22323 (N_22323,N_15950,N_16121);
nand U22324 (N_22324,N_19361,N_16717);
nor U22325 (N_22325,N_16326,N_15389);
nand U22326 (N_22326,N_19977,N_17831);
or U22327 (N_22327,N_19039,N_18477);
and U22328 (N_22328,N_17568,N_18896);
or U22329 (N_22329,N_17502,N_17915);
or U22330 (N_22330,N_16797,N_17572);
nor U22331 (N_22331,N_15281,N_19380);
or U22332 (N_22332,N_18012,N_16867);
or U22333 (N_22333,N_17868,N_18557);
nor U22334 (N_22334,N_16963,N_18103);
nor U22335 (N_22335,N_15521,N_16580);
nand U22336 (N_22336,N_17054,N_17098);
and U22337 (N_22337,N_15966,N_19485);
nand U22338 (N_22338,N_16951,N_17379);
nor U22339 (N_22339,N_15185,N_15125);
or U22340 (N_22340,N_17487,N_16613);
nand U22341 (N_22341,N_16810,N_17873);
xnor U22342 (N_22342,N_15259,N_17210);
or U22343 (N_22343,N_15289,N_15933);
nand U22344 (N_22344,N_15262,N_15117);
nand U22345 (N_22345,N_15723,N_17359);
xnor U22346 (N_22346,N_19124,N_16440);
nand U22347 (N_22347,N_19662,N_15118);
nor U22348 (N_22348,N_17278,N_17882);
nor U22349 (N_22349,N_19770,N_15445);
xnor U22350 (N_22350,N_16322,N_16418);
and U22351 (N_22351,N_18911,N_15225);
or U22352 (N_22352,N_18275,N_15596);
nand U22353 (N_22353,N_15476,N_15953);
nand U22354 (N_22354,N_19650,N_19164);
or U22355 (N_22355,N_17801,N_19590);
nand U22356 (N_22356,N_19367,N_18210);
xnor U22357 (N_22357,N_18753,N_17319);
and U22358 (N_22358,N_16330,N_17024);
nand U22359 (N_22359,N_19372,N_17732);
nor U22360 (N_22360,N_15677,N_15560);
or U22361 (N_22361,N_15304,N_18706);
xor U22362 (N_22362,N_17244,N_15971);
nand U22363 (N_22363,N_17293,N_19628);
or U22364 (N_22364,N_19545,N_17959);
nor U22365 (N_22365,N_17000,N_18450);
or U22366 (N_22366,N_15728,N_15951);
nand U22367 (N_22367,N_17400,N_16725);
nor U22368 (N_22368,N_15248,N_16837);
nor U22369 (N_22369,N_16815,N_17469);
nand U22370 (N_22370,N_15340,N_17146);
nand U22371 (N_22371,N_18527,N_15005);
or U22372 (N_22372,N_18837,N_19511);
nand U22373 (N_22373,N_19378,N_19428);
or U22374 (N_22374,N_17290,N_15605);
and U22375 (N_22375,N_19967,N_16431);
xor U22376 (N_22376,N_16155,N_19500);
and U22377 (N_22377,N_16839,N_18856);
nand U22378 (N_22378,N_18848,N_18616);
nor U22379 (N_22379,N_15996,N_19264);
nor U22380 (N_22380,N_17182,N_18667);
or U22381 (N_22381,N_18346,N_19823);
or U22382 (N_22382,N_16930,N_16260);
or U22383 (N_22383,N_19069,N_15775);
and U22384 (N_22384,N_18567,N_18878);
and U22385 (N_22385,N_17598,N_15722);
and U22386 (N_22386,N_16277,N_17626);
nand U22387 (N_22387,N_18161,N_19842);
nor U22388 (N_22388,N_15388,N_15400);
xor U22389 (N_22389,N_17253,N_19097);
nor U22390 (N_22390,N_15533,N_17556);
xnor U22391 (N_22391,N_17933,N_18120);
nand U22392 (N_22392,N_19464,N_17785);
nand U22393 (N_22393,N_15027,N_16993);
or U22394 (N_22394,N_16745,N_15637);
or U22395 (N_22395,N_17376,N_19944);
nor U22396 (N_22396,N_15121,N_19270);
and U22397 (N_22397,N_18824,N_19275);
and U22398 (N_22398,N_15693,N_19896);
and U22399 (N_22399,N_18379,N_16929);
and U22400 (N_22400,N_18470,N_19706);
nor U22401 (N_22401,N_17046,N_19192);
and U22402 (N_22402,N_19902,N_19390);
and U22403 (N_22403,N_17523,N_16760);
nor U22404 (N_22404,N_15293,N_19877);
nor U22405 (N_22405,N_19806,N_16486);
or U22406 (N_22406,N_19024,N_18395);
and U22407 (N_22407,N_19876,N_17177);
nor U22408 (N_22408,N_18577,N_16529);
nor U22409 (N_22409,N_18401,N_15665);
nor U22410 (N_22410,N_16921,N_17508);
or U22411 (N_22411,N_18143,N_18679);
nor U22412 (N_22412,N_18335,N_17117);
or U22413 (N_22413,N_18812,N_18901);
xnor U22414 (N_22414,N_18494,N_15480);
nand U22415 (N_22415,N_15695,N_15490);
and U22416 (N_22416,N_19866,N_18771);
nand U22417 (N_22417,N_17538,N_15782);
nor U22418 (N_22418,N_18910,N_16602);
or U22419 (N_22419,N_19643,N_18350);
xor U22420 (N_22420,N_18756,N_17750);
or U22421 (N_22421,N_18172,N_16075);
nand U22422 (N_22422,N_18970,N_18552);
nand U22423 (N_22423,N_19727,N_19049);
xnor U22424 (N_22424,N_17677,N_17133);
and U22425 (N_22425,N_19159,N_18920);
nor U22426 (N_22426,N_15136,N_15156);
or U22427 (N_22427,N_16611,N_17020);
and U22428 (N_22428,N_16478,N_16054);
nand U22429 (N_22429,N_19742,N_19263);
and U22430 (N_22430,N_16977,N_19915);
nand U22431 (N_22431,N_19715,N_16790);
nand U22432 (N_22432,N_18584,N_15557);
and U22433 (N_22433,N_19407,N_19969);
nor U22434 (N_22434,N_15253,N_18581);
and U22435 (N_22435,N_18582,N_19186);
nand U22436 (N_22436,N_15936,N_16261);
nand U22437 (N_22437,N_17908,N_17535);
nand U22438 (N_22438,N_17942,N_15532);
or U22439 (N_22439,N_15026,N_19744);
and U22440 (N_22440,N_16761,N_17702);
and U22441 (N_22441,N_15838,N_15202);
nand U22442 (N_22442,N_18811,N_19907);
xor U22443 (N_22443,N_15130,N_17830);
nand U22444 (N_22444,N_18802,N_18442);
and U22445 (N_22445,N_17741,N_17594);
nand U22446 (N_22446,N_16176,N_16381);
xnor U22447 (N_22447,N_19246,N_15646);
or U22448 (N_22448,N_18174,N_15991);
and U22449 (N_22449,N_18835,N_19685);
and U22450 (N_22450,N_19314,N_18597);
xnor U22451 (N_22451,N_18761,N_19149);
nand U22452 (N_22452,N_19686,N_17299);
or U22453 (N_22453,N_15072,N_17467);
nand U22454 (N_22454,N_15957,N_17488);
and U22455 (N_22455,N_17420,N_17223);
and U22456 (N_22456,N_19481,N_18914);
xnor U22457 (N_22457,N_17653,N_15094);
and U22458 (N_22458,N_15041,N_15970);
nor U22459 (N_22459,N_16913,N_18929);
nand U22460 (N_22460,N_19537,N_19879);
nand U22461 (N_22461,N_17498,N_18913);
or U22462 (N_22462,N_18360,N_15827);
and U22463 (N_22463,N_19547,N_15396);
nand U22464 (N_22464,N_16308,N_15437);
or U22465 (N_22465,N_17443,N_15724);
or U22466 (N_22466,N_19118,N_15759);
nor U22467 (N_22467,N_18118,N_16474);
or U22468 (N_22468,N_17767,N_18732);
nand U22469 (N_22469,N_19908,N_15562);
nor U22470 (N_22470,N_15485,N_17026);
and U22471 (N_22471,N_18773,N_18693);
or U22472 (N_22472,N_19584,N_16031);
or U22473 (N_22473,N_17638,N_18178);
and U22474 (N_22474,N_18375,N_16589);
nor U22475 (N_22475,N_19272,N_18788);
nor U22476 (N_22476,N_15217,N_18541);
or U22477 (N_22477,N_15165,N_16341);
nor U22478 (N_22478,N_17219,N_16803);
nor U22479 (N_22479,N_17697,N_19592);
nor U22480 (N_22480,N_15458,N_15018);
nor U22481 (N_22481,N_16046,N_18164);
or U22482 (N_22482,N_16421,N_19090);
and U22483 (N_22483,N_15662,N_15371);
nor U22484 (N_22484,N_16994,N_18061);
or U22485 (N_22485,N_18018,N_19599);
nand U22486 (N_22486,N_19625,N_19079);
and U22487 (N_22487,N_17058,N_17974);
nor U22488 (N_22488,N_19888,N_17799);
xor U22489 (N_22489,N_16116,N_18114);
or U22490 (N_22490,N_17289,N_18281);
and U22491 (N_22491,N_18888,N_19111);
or U22492 (N_22492,N_18728,N_16547);
nor U22493 (N_22493,N_18752,N_19899);
or U22494 (N_22494,N_18319,N_16674);
and U22495 (N_22495,N_19752,N_17436);
or U22496 (N_22496,N_16600,N_17097);
nor U22497 (N_22497,N_16804,N_18106);
nor U22498 (N_22498,N_15817,N_17512);
nand U22499 (N_22499,N_19262,N_17280);
and U22500 (N_22500,N_19506,N_18915);
nor U22501 (N_22501,N_15188,N_16063);
or U22502 (N_22502,N_15841,N_18533);
and U22503 (N_22503,N_15308,N_17195);
and U22504 (N_22504,N_19279,N_17856);
and U22505 (N_22505,N_18023,N_16954);
nand U22506 (N_22506,N_17241,N_18621);
or U22507 (N_22507,N_18847,N_17546);
and U22508 (N_22508,N_16884,N_19178);
nor U22509 (N_22509,N_16709,N_19107);
nor U22510 (N_22510,N_18461,N_18115);
nor U22511 (N_22511,N_16655,N_18712);
xnor U22512 (N_22512,N_17849,N_15564);
and U22513 (N_22513,N_17534,N_18096);
and U22514 (N_22514,N_18272,N_17072);
nand U22515 (N_22515,N_17677,N_15061);
xor U22516 (N_22516,N_16979,N_17423);
nand U22517 (N_22517,N_15458,N_15596);
or U22518 (N_22518,N_17891,N_19525);
nor U22519 (N_22519,N_19969,N_16347);
or U22520 (N_22520,N_18405,N_15876);
and U22521 (N_22521,N_16921,N_19760);
nor U22522 (N_22522,N_17305,N_15339);
nor U22523 (N_22523,N_19587,N_19968);
nand U22524 (N_22524,N_17911,N_16050);
nand U22525 (N_22525,N_18870,N_19789);
and U22526 (N_22526,N_18077,N_16546);
or U22527 (N_22527,N_18657,N_18024);
nand U22528 (N_22528,N_19838,N_16578);
and U22529 (N_22529,N_15867,N_15804);
or U22530 (N_22530,N_18290,N_16486);
nand U22531 (N_22531,N_17027,N_17371);
or U22532 (N_22532,N_16323,N_17147);
or U22533 (N_22533,N_15591,N_15515);
or U22534 (N_22534,N_16536,N_18723);
or U22535 (N_22535,N_15203,N_15016);
nand U22536 (N_22536,N_18516,N_15740);
or U22537 (N_22537,N_17844,N_15795);
and U22538 (N_22538,N_15634,N_19342);
and U22539 (N_22539,N_17296,N_15940);
and U22540 (N_22540,N_15812,N_16266);
nand U22541 (N_22541,N_18691,N_18376);
and U22542 (N_22542,N_17731,N_18133);
xnor U22543 (N_22543,N_18408,N_19498);
and U22544 (N_22544,N_18691,N_17773);
and U22545 (N_22545,N_16253,N_15736);
or U22546 (N_22546,N_16356,N_16022);
and U22547 (N_22547,N_19932,N_15760);
nor U22548 (N_22548,N_17859,N_18103);
xnor U22549 (N_22549,N_18224,N_19149);
and U22550 (N_22550,N_19089,N_17457);
nand U22551 (N_22551,N_19697,N_15922);
or U22552 (N_22552,N_16912,N_18859);
and U22553 (N_22553,N_16863,N_15632);
nor U22554 (N_22554,N_15501,N_16783);
nand U22555 (N_22555,N_18274,N_18625);
or U22556 (N_22556,N_19517,N_18940);
nor U22557 (N_22557,N_19258,N_18865);
and U22558 (N_22558,N_19572,N_19557);
nor U22559 (N_22559,N_18614,N_17445);
nand U22560 (N_22560,N_18344,N_16793);
nand U22561 (N_22561,N_16983,N_18922);
or U22562 (N_22562,N_17103,N_16890);
xor U22563 (N_22563,N_15846,N_18762);
xor U22564 (N_22564,N_19208,N_18804);
xnor U22565 (N_22565,N_16925,N_18878);
and U22566 (N_22566,N_15805,N_18318);
or U22567 (N_22567,N_15230,N_19453);
and U22568 (N_22568,N_16665,N_16960);
nand U22569 (N_22569,N_18031,N_19572);
nor U22570 (N_22570,N_17178,N_18697);
nor U22571 (N_22571,N_16517,N_18290);
or U22572 (N_22572,N_18908,N_18560);
or U22573 (N_22573,N_19899,N_19666);
nand U22574 (N_22574,N_17144,N_18860);
and U22575 (N_22575,N_16348,N_19340);
and U22576 (N_22576,N_19075,N_18217);
or U22577 (N_22577,N_15575,N_16452);
xnor U22578 (N_22578,N_18006,N_15662);
or U22579 (N_22579,N_15662,N_17452);
nand U22580 (N_22580,N_19239,N_17528);
xnor U22581 (N_22581,N_15592,N_15818);
nor U22582 (N_22582,N_15169,N_15311);
nor U22583 (N_22583,N_15294,N_16815);
nand U22584 (N_22584,N_15533,N_16137);
nand U22585 (N_22585,N_19137,N_19369);
nand U22586 (N_22586,N_15087,N_16119);
nor U22587 (N_22587,N_17830,N_16074);
nor U22588 (N_22588,N_19586,N_17613);
and U22589 (N_22589,N_15581,N_18144);
nor U22590 (N_22590,N_17477,N_19491);
or U22591 (N_22591,N_19395,N_19280);
nor U22592 (N_22592,N_17752,N_15557);
nand U22593 (N_22593,N_16661,N_17054);
nor U22594 (N_22594,N_18090,N_18149);
nor U22595 (N_22595,N_17433,N_16602);
and U22596 (N_22596,N_17067,N_19243);
and U22597 (N_22597,N_17286,N_18984);
xor U22598 (N_22598,N_17556,N_17044);
nand U22599 (N_22599,N_19259,N_15273);
nand U22600 (N_22600,N_18924,N_18734);
nor U22601 (N_22601,N_17253,N_18046);
nor U22602 (N_22602,N_16907,N_18845);
nand U22603 (N_22603,N_16257,N_19250);
or U22604 (N_22604,N_16054,N_17252);
xnor U22605 (N_22605,N_15292,N_18577);
nand U22606 (N_22606,N_19603,N_18974);
nor U22607 (N_22607,N_17044,N_18969);
and U22608 (N_22608,N_16998,N_15729);
and U22609 (N_22609,N_18298,N_17097);
nand U22610 (N_22610,N_15193,N_19453);
xor U22611 (N_22611,N_18128,N_19492);
or U22612 (N_22612,N_17950,N_15618);
xnor U22613 (N_22613,N_18956,N_16194);
and U22614 (N_22614,N_17083,N_16666);
nand U22615 (N_22615,N_19614,N_19469);
nand U22616 (N_22616,N_17088,N_18187);
nand U22617 (N_22617,N_15778,N_16099);
xor U22618 (N_22618,N_18022,N_19049);
and U22619 (N_22619,N_16369,N_15888);
xnor U22620 (N_22620,N_17028,N_18729);
nand U22621 (N_22621,N_16034,N_15699);
nand U22622 (N_22622,N_17861,N_17127);
nor U22623 (N_22623,N_17065,N_19954);
or U22624 (N_22624,N_18931,N_19437);
nand U22625 (N_22625,N_15472,N_18883);
nor U22626 (N_22626,N_15643,N_16834);
and U22627 (N_22627,N_17287,N_17558);
nand U22628 (N_22628,N_18362,N_19694);
and U22629 (N_22629,N_16074,N_18284);
nor U22630 (N_22630,N_18361,N_19753);
xnor U22631 (N_22631,N_18191,N_19686);
nor U22632 (N_22632,N_17898,N_16736);
xor U22633 (N_22633,N_17457,N_17515);
or U22634 (N_22634,N_19147,N_18470);
nand U22635 (N_22635,N_18977,N_19848);
nand U22636 (N_22636,N_19093,N_15269);
and U22637 (N_22637,N_18271,N_19412);
xor U22638 (N_22638,N_19539,N_18627);
nor U22639 (N_22639,N_18419,N_18045);
and U22640 (N_22640,N_15914,N_18453);
nor U22641 (N_22641,N_17278,N_18290);
nor U22642 (N_22642,N_19226,N_18086);
or U22643 (N_22643,N_18716,N_19448);
and U22644 (N_22644,N_17300,N_16888);
and U22645 (N_22645,N_15817,N_19990);
and U22646 (N_22646,N_18443,N_16028);
or U22647 (N_22647,N_19066,N_16226);
nand U22648 (N_22648,N_19016,N_19489);
and U22649 (N_22649,N_19237,N_18625);
nor U22650 (N_22650,N_18066,N_15331);
nor U22651 (N_22651,N_19816,N_19524);
nor U22652 (N_22652,N_15327,N_15268);
and U22653 (N_22653,N_18199,N_15855);
nor U22654 (N_22654,N_17437,N_17343);
nand U22655 (N_22655,N_15079,N_17057);
and U22656 (N_22656,N_18137,N_16435);
xnor U22657 (N_22657,N_15507,N_18476);
nor U22658 (N_22658,N_16191,N_19502);
xor U22659 (N_22659,N_17119,N_15321);
nand U22660 (N_22660,N_15103,N_16089);
and U22661 (N_22661,N_19146,N_18431);
and U22662 (N_22662,N_19202,N_16826);
nor U22663 (N_22663,N_16038,N_16646);
or U22664 (N_22664,N_18090,N_16989);
xor U22665 (N_22665,N_18519,N_19720);
and U22666 (N_22666,N_15590,N_15188);
or U22667 (N_22667,N_18813,N_16144);
nor U22668 (N_22668,N_15847,N_15073);
or U22669 (N_22669,N_19858,N_16384);
nor U22670 (N_22670,N_18543,N_15053);
xor U22671 (N_22671,N_15527,N_17609);
and U22672 (N_22672,N_15326,N_16921);
xnor U22673 (N_22673,N_18967,N_16663);
and U22674 (N_22674,N_18068,N_18808);
xor U22675 (N_22675,N_19399,N_19337);
nand U22676 (N_22676,N_16849,N_17131);
nand U22677 (N_22677,N_15300,N_15237);
or U22678 (N_22678,N_19207,N_17370);
nand U22679 (N_22679,N_16853,N_18604);
xor U22680 (N_22680,N_18090,N_16344);
or U22681 (N_22681,N_18847,N_18310);
and U22682 (N_22682,N_16668,N_16137);
nor U22683 (N_22683,N_18532,N_17694);
nand U22684 (N_22684,N_17729,N_16435);
and U22685 (N_22685,N_17721,N_17660);
nand U22686 (N_22686,N_19365,N_19850);
and U22687 (N_22687,N_18462,N_17815);
xnor U22688 (N_22688,N_15387,N_15246);
or U22689 (N_22689,N_18413,N_18805);
nor U22690 (N_22690,N_15098,N_16313);
nor U22691 (N_22691,N_18748,N_16005);
nand U22692 (N_22692,N_16954,N_18163);
nand U22693 (N_22693,N_19341,N_15433);
nor U22694 (N_22694,N_18164,N_17891);
or U22695 (N_22695,N_15315,N_15785);
and U22696 (N_22696,N_16581,N_15306);
nor U22697 (N_22697,N_16040,N_17970);
nor U22698 (N_22698,N_16736,N_15636);
nor U22699 (N_22699,N_19406,N_19498);
or U22700 (N_22700,N_15010,N_18642);
and U22701 (N_22701,N_19867,N_17450);
and U22702 (N_22702,N_18807,N_15725);
or U22703 (N_22703,N_18651,N_17549);
or U22704 (N_22704,N_15379,N_16938);
and U22705 (N_22705,N_15514,N_17906);
or U22706 (N_22706,N_18289,N_18669);
nor U22707 (N_22707,N_19834,N_18909);
nand U22708 (N_22708,N_17332,N_15311);
xor U22709 (N_22709,N_15971,N_17506);
xnor U22710 (N_22710,N_18715,N_17069);
and U22711 (N_22711,N_19133,N_18306);
nand U22712 (N_22712,N_19531,N_17435);
nor U22713 (N_22713,N_18520,N_16290);
or U22714 (N_22714,N_17635,N_17090);
or U22715 (N_22715,N_15056,N_17836);
nor U22716 (N_22716,N_19638,N_17998);
or U22717 (N_22717,N_15255,N_17112);
and U22718 (N_22718,N_16037,N_16704);
and U22719 (N_22719,N_19227,N_18800);
nor U22720 (N_22720,N_18975,N_18904);
nand U22721 (N_22721,N_19084,N_18686);
or U22722 (N_22722,N_19130,N_16798);
and U22723 (N_22723,N_17703,N_16684);
or U22724 (N_22724,N_19350,N_16354);
or U22725 (N_22725,N_17359,N_16232);
nor U22726 (N_22726,N_16112,N_17921);
and U22727 (N_22727,N_17900,N_18660);
or U22728 (N_22728,N_17365,N_15649);
or U22729 (N_22729,N_16435,N_17043);
or U22730 (N_22730,N_19589,N_17814);
and U22731 (N_22731,N_17209,N_18413);
or U22732 (N_22732,N_16353,N_19942);
or U22733 (N_22733,N_17934,N_18223);
nand U22734 (N_22734,N_18411,N_19821);
nand U22735 (N_22735,N_19831,N_17375);
xnor U22736 (N_22736,N_15867,N_15780);
and U22737 (N_22737,N_18247,N_15558);
and U22738 (N_22738,N_19808,N_19357);
nor U22739 (N_22739,N_16895,N_16084);
and U22740 (N_22740,N_16072,N_15476);
nand U22741 (N_22741,N_18688,N_15285);
and U22742 (N_22742,N_16906,N_16613);
and U22743 (N_22743,N_16096,N_16156);
or U22744 (N_22744,N_15395,N_17189);
and U22745 (N_22745,N_18174,N_16178);
or U22746 (N_22746,N_18809,N_19475);
and U22747 (N_22747,N_15194,N_18682);
nand U22748 (N_22748,N_19339,N_19532);
and U22749 (N_22749,N_17165,N_17696);
or U22750 (N_22750,N_18122,N_15459);
nor U22751 (N_22751,N_16429,N_19658);
and U22752 (N_22752,N_18377,N_17711);
xnor U22753 (N_22753,N_15458,N_16255);
and U22754 (N_22754,N_19689,N_17454);
nand U22755 (N_22755,N_18925,N_19038);
nor U22756 (N_22756,N_16516,N_15149);
and U22757 (N_22757,N_15834,N_18505);
or U22758 (N_22758,N_18241,N_15859);
and U22759 (N_22759,N_18566,N_16298);
nand U22760 (N_22760,N_17761,N_16479);
nand U22761 (N_22761,N_18747,N_17188);
and U22762 (N_22762,N_18935,N_15701);
nand U22763 (N_22763,N_19735,N_19161);
or U22764 (N_22764,N_17363,N_19194);
nor U22765 (N_22765,N_19463,N_16664);
xor U22766 (N_22766,N_15980,N_16536);
xor U22767 (N_22767,N_19409,N_19216);
xor U22768 (N_22768,N_15864,N_18415);
and U22769 (N_22769,N_15521,N_15695);
or U22770 (N_22770,N_17210,N_19460);
and U22771 (N_22771,N_16230,N_17589);
nand U22772 (N_22772,N_19292,N_17296);
nand U22773 (N_22773,N_16498,N_15017);
or U22774 (N_22774,N_17727,N_17763);
or U22775 (N_22775,N_19237,N_19391);
and U22776 (N_22776,N_18589,N_16636);
and U22777 (N_22777,N_16004,N_18562);
and U22778 (N_22778,N_16187,N_17027);
nand U22779 (N_22779,N_16544,N_18664);
nor U22780 (N_22780,N_19480,N_16469);
nor U22781 (N_22781,N_15635,N_17010);
nand U22782 (N_22782,N_15513,N_16157);
nand U22783 (N_22783,N_15307,N_18521);
or U22784 (N_22784,N_15620,N_15737);
and U22785 (N_22785,N_15557,N_19647);
nor U22786 (N_22786,N_19412,N_19227);
nor U22787 (N_22787,N_17882,N_15636);
xnor U22788 (N_22788,N_16421,N_15705);
and U22789 (N_22789,N_15648,N_18949);
nand U22790 (N_22790,N_17666,N_16506);
and U22791 (N_22791,N_19235,N_18932);
and U22792 (N_22792,N_18798,N_17008);
or U22793 (N_22793,N_18701,N_19511);
nor U22794 (N_22794,N_16923,N_19441);
and U22795 (N_22795,N_17855,N_18860);
nand U22796 (N_22796,N_15231,N_17033);
or U22797 (N_22797,N_16833,N_18160);
and U22798 (N_22798,N_17381,N_15697);
or U22799 (N_22799,N_16690,N_18321);
nand U22800 (N_22800,N_15868,N_16964);
or U22801 (N_22801,N_16653,N_16778);
and U22802 (N_22802,N_17859,N_18786);
nand U22803 (N_22803,N_19869,N_15413);
nor U22804 (N_22804,N_15050,N_15149);
or U22805 (N_22805,N_17603,N_17275);
and U22806 (N_22806,N_19003,N_16148);
nand U22807 (N_22807,N_16253,N_19254);
nand U22808 (N_22808,N_15157,N_15755);
nand U22809 (N_22809,N_17970,N_19841);
and U22810 (N_22810,N_15220,N_15123);
and U22811 (N_22811,N_17280,N_15175);
nor U22812 (N_22812,N_19064,N_17213);
or U22813 (N_22813,N_19288,N_19868);
nand U22814 (N_22814,N_16211,N_16755);
or U22815 (N_22815,N_19965,N_16626);
xnor U22816 (N_22816,N_17072,N_19521);
and U22817 (N_22817,N_18388,N_19243);
nand U22818 (N_22818,N_19300,N_17264);
and U22819 (N_22819,N_19969,N_16699);
and U22820 (N_22820,N_19848,N_18658);
nand U22821 (N_22821,N_15348,N_19665);
xnor U22822 (N_22822,N_17637,N_19685);
or U22823 (N_22823,N_19615,N_17571);
nand U22824 (N_22824,N_17680,N_18211);
or U22825 (N_22825,N_19741,N_15255);
nor U22826 (N_22826,N_17097,N_15356);
xor U22827 (N_22827,N_15748,N_19451);
or U22828 (N_22828,N_16163,N_16072);
nor U22829 (N_22829,N_16962,N_17565);
nand U22830 (N_22830,N_16752,N_18121);
nor U22831 (N_22831,N_18590,N_15992);
nor U22832 (N_22832,N_15040,N_16780);
or U22833 (N_22833,N_18586,N_16382);
or U22834 (N_22834,N_17443,N_16438);
nand U22835 (N_22835,N_15129,N_17094);
xnor U22836 (N_22836,N_15321,N_17635);
nor U22837 (N_22837,N_18874,N_18112);
or U22838 (N_22838,N_19627,N_18359);
and U22839 (N_22839,N_19627,N_17218);
and U22840 (N_22840,N_15326,N_18987);
nand U22841 (N_22841,N_17807,N_19868);
nand U22842 (N_22842,N_16152,N_17047);
or U22843 (N_22843,N_17457,N_15492);
xor U22844 (N_22844,N_15565,N_19220);
nor U22845 (N_22845,N_16676,N_15886);
xnor U22846 (N_22846,N_15621,N_15652);
and U22847 (N_22847,N_15093,N_16958);
or U22848 (N_22848,N_18260,N_16999);
xor U22849 (N_22849,N_18295,N_16532);
or U22850 (N_22850,N_18901,N_19103);
nor U22851 (N_22851,N_15065,N_15737);
and U22852 (N_22852,N_17654,N_17766);
nor U22853 (N_22853,N_19396,N_16988);
and U22854 (N_22854,N_17552,N_16170);
and U22855 (N_22855,N_16498,N_16581);
xor U22856 (N_22856,N_19526,N_17400);
xnor U22857 (N_22857,N_16066,N_15507);
and U22858 (N_22858,N_17538,N_16940);
and U22859 (N_22859,N_19542,N_17847);
nand U22860 (N_22860,N_18049,N_16256);
nand U22861 (N_22861,N_18054,N_15569);
nor U22862 (N_22862,N_17107,N_16090);
nor U22863 (N_22863,N_18048,N_18100);
xnor U22864 (N_22864,N_17492,N_15376);
nand U22865 (N_22865,N_16643,N_15620);
or U22866 (N_22866,N_16125,N_18366);
and U22867 (N_22867,N_18079,N_15834);
nand U22868 (N_22868,N_17297,N_17401);
and U22869 (N_22869,N_17896,N_16115);
nor U22870 (N_22870,N_17899,N_16497);
and U22871 (N_22871,N_19710,N_16653);
or U22872 (N_22872,N_17334,N_15999);
nand U22873 (N_22873,N_16135,N_15838);
and U22874 (N_22874,N_19838,N_17943);
or U22875 (N_22875,N_15292,N_18259);
nor U22876 (N_22876,N_15066,N_16006);
nand U22877 (N_22877,N_16715,N_17485);
and U22878 (N_22878,N_15753,N_19860);
and U22879 (N_22879,N_17730,N_17919);
nand U22880 (N_22880,N_19456,N_16217);
or U22881 (N_22881,N_19764,N_19962);
or U22882 (N_22882,N_15608,N_18849);
or U22883 (N_22883,N_15931,N_17417);
nor U22884 (N_22884,N_15208,N_16912);
and U22885 (N_22885,N_17943,N_17610);
or U22886 (N_22886,N_18425,N_18963);
or U22887 (N_22887,N_18228,N_15610);
nor U22888 (N_22888,N_16112,N_17578);
nand U22889 (N_22889,N_15677,N_17221);
nand U22890 (N_22890,N_15946,N_17648);
nor U22891 (N_22891,N_19517,N_19191);
or U22892 (N_22892,N_19216,N_15083);
nor U22893 (N_22893,N_18686,N_19540);
nor U22894 (N_22894,N_15289,N_18681);
nand U22895 (N_22895,N_15109,N_16984);
and U22896 (N_22896,N_17719,N_18512);
nand U22897 (N_22897,N_18941,N_17380);
nand U22898 (N_22898,N_16915,N_19302);
and U22899 (N_22899,N_19346,N_16661);
or U22900 (N_22900,N_17016,N_16839);
nor U22901 (N_22901,N_15030,N_16082);
nor U22902 (N_22902,N_18140,N_17636);
xnor U22903 (N_22903,N_17729,N_15843);
nand U22904 (N_22904,N_17498,N_17484);
nand U22905 (N_22905,N_15116,N_16667);
or U22906 (N_22906,N_17278,N_18744);
nor U22907 (N_22907,N_18136,N_19526);
and U22908 (N_22908,N_19593,N_19196);
or U22909 (N_22909,N_17040,N_15398);
nor U22910 (N_22910,N_18068,N_16394);
nand U22911 (N_22911,N_19268,N_16565);
nand U22912 (N_22912,N_19044,N_17931);
or U22913 (N_22913,N_16001,N_19481);
and U22914 (N_22914,N_19750,N_19094);
nor U22915 (N_22915,N_15058,N_16325);
or U22916 (N_22916,N_15767,N_17591);
nor U22917 (N_22917,N_16414,N_18210);
and U22918 (N_22918,N_17091,N_19175);
nand U22919 (N_22919,N_19803,N_17041);
and U22920 (N_22920,N_16759,N_18333);
and U22921 (N_22921,N_15855,N_17649);
nand U22922 (N_22922,N_16904,N_19551);
nor U22923 (N_22923,N_17648,N_17226);
or U22924 (N_22924,N_16945,N_19679);
and U22925 (N_22925,N_17030,N_16709);
or U22926 (N_22926,N_19551,N_17747);
and U22927 (N_22927,N_19365,N_17315);
nor U22928 (N_22928,N_19718,N_19175);
or U22929 (N_22929,N_17250,N_19729);
xor U22930 (N_22930,N_16972,N_15479);
nand U22931 (N_22931,N_18903,N_17343);
or U22932 (N_22932,N_17667,N_16935);
and U22933 (N_22933,N_16012,N_18964);
and U22934 (N_22934,N_17343,N_15645);
xor U22935 (N_22935,N_19801,N_15032);
or U22936 (N_22936,N_17910,N_16127);
and U22937 (N_22937,N_16806,N_17049);
or U22938 (N_22938,N_18510,N_17395);
xnor U22939 (N_22939,N_19908,N_17274);
nor U22940 (N_22940,N_15174,N_19502);
or U22941 (N_22941,N_17402,N_19147);
xnor U22942 (N_22942,N_18601,N_16028);
or U22943 (N_22943,N_19744,N_16016);
nand U22944 (N_22944,N_15025,N_17913);
or U22945 (N_22945,N_19367,N_17410);
xnor U22946 (N_22946,N_19533,N_17603);
nand U22947 (N_22947,N_15488,N_19288);
nor U22948 (N_22948,N_17378,N_16838);
or U22949 (N_22949,N_17802,N_15522);
and U22950 (N_22950,N_15545,N_16503);
nor U22951 (N_22951,N_19079,N_15856);
and U22952 (N_22952,N_18569,N_18982);
nor U22953 (N_22953,N_15019,N_17936);
nand U22954 (N_22954,N_15975,N_17485);
or U22955 (N_22955,N_19648,N_18184);
and U22956 (N_22956,N_15489,N_17898);
nand U22957 (N_22957,N_19428,N_16211);
xor U22958 (N_22958,N_17208,N_17233);
and U22959 (N_22959,N_19959,N_19586);
nor U22960 (N_22960,N_18070,N_15981);
and U22961 (N_22961,N_17776,N_16788);
xor U22962 (N_22962,N_17559,N_15849);
and U22963 (N_22963,N_18173,N_18261);
nand U22964 (N_22964,N_15770,N_18758);
and U22965 (N_22965,N_15832,N_16889);
nor U22966 (N_22966,N_16523,N_18420);
nand U22967 (N_22967,N_18886,N_19583);
or U22968 (N_22968,N_16856,N_19123);
xnor U22969 (N_22969,N_19509,N_17424);
nor U22970 (N_22970,N_17339,N_17335);
nand U22971 (N_22971,N_16464,N_15479);
or U22972 (N_22972,N_19400,N_15741);
or U22973 (N_22973,N_15726,N_16674);
and U22974 (N_22974,N_19403,N_18445);
nor U22975 (N_22975,N_16849,N_19742);
nand U22976 (N_22976,N_17895,N_17801);
nor U22977 (N_22977,N_18338,N_17828);
and U22978 (N_22978,N_18476,N_18309);
or U22979 (N_22979,N_19548,N_16613);
or U22980 (N_22980,N_19807,N_19006);
or U22981 (N_22981,N_16422,N_17974);
or U22982 (N_22982,N_17588,N_18342);
nor U22983 (N_22983,N_19679,N_15538);
nand U22984 (N_22984,N_15361,N_16525);
xnor U22985 (N_22985,N_18535,N_18149);
and U22986 (N_22986,N_15236,N_19896);
or U22987 (N_22987,N_19664,N_18923);
xor U22988 (N_22988,N_19180,N_19892);
nand U22989 (N_22989,N_18424,N_16966);
or U22990 (N_22990,N_19897,N_16831);
nand U22991 (N_22991,N_15296,N_18490);
nor U22992 (N_22992,N_15125,N_17169);
and U22993 (N_22993,N_17202,N_18641);
or U22994 (N_22994,N_16341,N_18175);
and U22995 (N_22995,N_16555,N_19046);
nor U22996 (N_22996,N_17916,N_17265);
and U22997 (N_22997,N_16128,N_15995);
xor U22998 (N_22998,N_18070,N_19539);
xor U22999 (N_22999,N_17317,N_18978);
or U23000 (N_23000,N_16531,N_19213);
or U23001 (N_23001,N_19470,N_15507);
nor U23002 (N_23002,N_16121,N_18781);
nand U23003 (N_23003,N_17237,N_17511);
and U23004 (N_23004,N_17686,N_15269);
nand U23005 (N_23005,N_15977,N_19408);
xnor U23006 (N_23006,N_17054,N_19883);
xor U23007 (N_23007,N_17709,N_15679);
nor U23008 (N_23008,N_15053,N_17845);
nand U23009 (N_23009,N_18923,N_19336);
nor U23010 (N_23010,N_16491,N_15019);
nor U23011 (N_23011,N_18557,N_16687);
or U23012 (N_23012,N_15630,N_15118);
or U23013 (N_23013,N_18412,N_15909);
nand U23014 (N_23014,N_19697,N_18072);
and U23015 (N_23015,N_16236,N_15241);
or U23016 (N_23016,N_18448,N_17518);
nor U23017 (N_23017,N_16586,N_17685);
and U23018 (N_23018,N_19201,N_16263);
xnor U23019 (N_23019,N_19485,N_16144);
and U23020 (N_23020,N_19697,N_16701);
or U23021 (N_23021,N_16623,N_17532);
nand U23022 (N_23022,N_17526,N_18492);
or U23023 (N_23023,N_19661,N_17722);
nand U23024 (N_23024,N_18796,N_17258);
or U23025 (N_23025,N_15807,N_15888);
nand U23026 (N_23026,N_19820,N_19332);
nor U23027 (N_23027,N_15239,N_19790);
and U23028 (N_23028,N_19264,N_17473);
nor U23029 (N_23029,N_15133,N_16625);
or U23030 (N_23030,N_16456,N_16067);
nor U23031 (N_23031,N_16026,N_15333);
xnor U23032 (N_23032,N_15484,N_19816);
nor U23033 (N_23033,N_15698,N_15133);
xor U23034 (N_23034,N_17199,N_16070);
or U23035 (N_23035,N_15417,N_18166);
nor U23036 (N_23036,N_19649,N_16717);
nand U23037 (N_23037,N_16321,N_15709);
nand U23038 (N_23038,N_19372,N_17387);
and U23039 (N_23039,N_15501,N_19502);
and U23040 (N_23040,N_16772,N_18000);
or U23041 (N_23041,N_19320,N_15953);
nand U23042 (N_23042,N_19014,N_19012);
and U23043 (N_23043,N_15967,N_16856);
and U23044 (N_23044,N_16013,N_18425);
xnor U23045 (N_23045,N_18915,N_17927);
and U23046 (N_23046,N_18987,N_18688);
xor U23047 (N_23047,N_19503,N_19865);
nor U23048 (N_23048,N_15425,N_17351);
or U23049 (N_23049,N_18017,N_15786);
or U23050 (N_23050,N_18860,N_19607);
nor U23051 (N_23051,N_17889,N_17115);
or U23052 (N_23052,N_19242,N_17090);
or U23053 (N_23053,N_19557,N_16382);
nor U23054 (N_23054,N_19070,N_18547);
and U23055 (N_23055,N_17296,N_15763);
nor U23056 (N_23056,N_17960,N_16935);
and U23057 (N_23057,N_17540,N_18868);
nand U23058 (N_23058,N_18586,N_16478);
xnor U23059 (N_23059,N_16378,N_16825);
and U23060 (N_23060,N_17922,N_19628);
nor U23061 (N_23061,N_19337,N_19257);
xnor U23062 (N_23062,N_17950,N_16353);
and U23063 (N_23063,N_15744,N_18615);
nand U23064 (N_23064,N_19183,N_17010);
and U23065 (N_23065,N_17256,N_17522);
xnor U23066 (N_23066,N_17088,N_19709);
or U23067 (N_23067,N_15671,N_15011);
nand U23068 (N_23068,N_17723,N_16633);
and U23069 (N_23069,N_16971,N_15170);
and U23070 (N_23070,N_18786,N_16785);
or U23071 (N_23071,N_15729,N_18848);
and U23072 (N_23072,N_18296,N_19224);
and U23073 (N_23073,N_18138,N_15578);
and U23074 (N_23074,N_17956,N_16298);
or U23075 (N_23075,N_18898,N_19313);
nand U23076 (N_23076,N_15210,N_15924);
nor U23077 (N_23077,N_18772,N_19980);
or U23078 (N_23078,N_16268,N_15486);
or U23079 (N_23079,N_15367,N_17003);
nor U23080 (N_23080,N_17863,N_17131);
nand U23081 (N_23081,N_15069,N_18893);
or U23082 (N_23082,N_15198,N_16333);
nand U23083 (N_23083,N_19844,N_16493);
nand U23084 (N_23084,N_16056,N_17989);
nor U23085 (N_23085,N_16877,N_15437);
nor U23086 (N_23086,N_18662,N_19266);
and U23087 (N_23087,N_16028,N_17002);
or U23088 (N_23088,N_17665,N_16832);
nor U23089 (N_23089,N_17716,N_19074);
nand U23090 (N_23090,N_18751,N_18837);
nand U23091 (N_23091,N_19227,N_18207);
nand U23092 (N_23092,N_16958,N_17091);
or U23093 (N_23093,N_19090,N_17673);
nor U23094 (N_23094,N_17702,N_15344);
nand U23095 (N_23095,N_18668,N_15083);
or U23096 (N_23096,N_17789,N_16271);
nor U23097 (N_23097,N_16805,N_15594);
and U23098 (N_23098,N_19292,N_17856);
and U23099 (N_23099,N_16257,N_15896);
or U23100 (N_23100,N_15374,N_15647);
nand U23101 (N_23101,N_17903,N_19729);
or U23102 (N_23102,N_19790,N_19248);
or U23103 (N_23103,N_16931,N_17198);
nand U23104 (N_23104,N_16469,N_19627);
nor U23105 (N_23105,N_17271,N_16805);
xnor U23106 (N_23106,N_19378,N_17810);
or U23107 (N_23107,N_18727,N_17769);
or U23108 (N_23108,N_17811,N_16331);
and U23109 (N_23109,N_16986,N_15724);
or U23110 (N_23110,N_16122,N_18135);
nor U23111 (N_23111,N_16714,N_18028);
or U23112 (N_23112,N_19021,N_15347);
nor U23113 (N_23113,N_16973,N_17889);
or U23114 (N_23114,N_15014,N_15839);
nor U23115 (N_23115,N_17947,N_17788);
nor U23116 (N_23116,N_15862,N_19905);
nor U23117 (N_23117,N_16616,N_19084);
xor U23118 (N_23118,N_19064,N_17959);
nand U23119 (N_23119,N_18331,N_19196);
nand U23120 (N_23120,N_17600,N_19119);
or U23121 (N_23121,N_15987,N_15917);
nand U23122 (N_23122,N_18622,N_16801);
nand U23123 (N_23123,N_18491,N_19498);
or U23124 (N_23124,N_18794,N_15436);
xnor U23125 (N_23125,N_17791,N_16787);
or U23126 (N_23126,N_18341,N_15598);
nand U23127 (N_23127,N_15366,N_16502);
or U23128 (N_23128,N_17581,N_15280);
nand U23129 (N_23129,N_17826,N_16011);
nor U23130 (N_23130,N_16934,N_16389);
nand U23131 (N_23131,N_19680,N_19541);
and U23132 (N_23132,N_19192,N_15851);
nor U23133 (N_23133,N_19459,N_19300);
nand U23134 (N_23134,N_16591,N_17185);
nand U23135 (N_23135,N_16334,N_15332);
or U23136 (N_23136,N_16738,N_19996);
nor U23137 (N_23137,N_19839,N_16159);
or U23138 (N_23138,N_15141,N_16703);
or U23139 (N_23139,N_15189,N_17827);
and U23140 (N_23140,N_18924,N_16829);
nand U23141 (N_23141,N_16692,N_15547);
nand U23142 (N_23142,N_18070,N_16063);
nand U23143 (N_23143,N_19836,N_16436);
or U23144 (N_23144,N_15611,N_18112);
nand U23145 (N_23145,N_17177,N_17108);
and U23146 (N_23146,N_17021,N_18379);
and U23147 (N_23147,N_17705,N_18125);
nand U23148 (N_23148,N_15179,N_16856);
nand U23149 (N_23149,N_17889,N_18423);
or U23150 (N_23150,N_15063,N_17464);
nand U23151 (N_23151,N_15860,N_18771);
or U23152 (N_23152,N_17860,N_16950);
xnor U23153 (N_23153,N_16012,N_19397);
nor U23154 (N_23154,N_19640,N_16370);
nand U23155 (N_23155,N_16440,N_18020);
nand U23156 (N_23156,N_16253,N_18786);
nand U23157 (N_23157,N_15117,N_16932);
nand U23158 (N_23158,N_18160,N_16528);
or U23159 (N_23159,N_19166,N_19121);
or U23160 (N_23160,N_18853,N_16918);
or U23161 (N_23161,N_19394,N_16539);
nor U23162 (N_23162,N_16525,N_16857);
and U23163 (N_23163,N_19900,N_17563);
and U23164 (N_23164,N_19242,N_17137);
or U23165 (N_23165,N_16370,N_17709);
and U23166 (N_23166,N_15116,N_18795);
and U23167 (N_23167,N_16025,N_17490);
and U23168 (N_23168,N_15715,N_17919);
or U23169 (N_23169,N_17158,N_15841);
and U23170 (N_23170,N_17276,N_17415);
and U23171 (N_23171,N_15134,N_19158);
nor U23172 (N_23172,N_19705,N_15718);
or U23173 (N_23173,N_18766,N_15628);
and U23174 (N_23174,N_17098,N_18806);
nand U23175 (N_23175,N_19507,N_15379);
nor U23176 (N_23176,N_15284,N_17909);
and U23177 (N_23177,N_15217,N_17930);
or U23178 (N_23178,N_18904,N_15205);
or U23179 (N_23179,N_16238,N_17761);
nand U23180 (N_23180,N_19029,N_16647);
nand U23181 (N_23181,N_17813,N_18617);
nand U23182 (N_23182,N_18508,N_17507);
or U23183 (N_23183,N_18542,N_15976);
nand U23184 (N_23184,N_15457,N_16338);
or U23185 (N_23185,N_18558,N_17498);
or U23186 (N_23186,N_19205,N_18514);
nand U23187 (N_23187,N_19452,N_18565);
nor U23188 (N_23188,N_17844,N_16849);
or U23189 (N_23189,N_18955,N_16876);
xor U23190 (N_23190,N_17622,N_16729);
nor U23191 (N_23191,N_15453,N_18007);
or U23192 (N_23192,N_18492,N_18818);
nor U23193 (N_23193,N_17843,N_18455);
nor U23194 (N_23194,N_15414,N_18956);
nor U23195 (N_23195,N_18840,N_15433);
nor U23196 (N_23196,N_18734,N_19237);
or U23197 (N_23197,N_16439,N_15427);
and U23198 (N_23198,N_18588,N_18993);
nor U23199 (N_23199,N_19163,N_19598);
nand U23200 (N_23200,N_19554,N_16263);
nand U23201 (N_23201,N_19824,N_16274);
and U23202 (N_23202,N_15010,N_15820);
nand U23203 (N_23203,N_15445,N_18012);
nor U23204 (N_23204,N_18713,N_18900);
or U23205 (N_23205,N_17603,N_17634);
or U23206 (N_23206,N_16002,N_16555);
nand U23207 (N_23207,N_17914,N_17649);
or U23208 (N_23208,N_16684,N_15886);
xnor U23209 (N_23209,N_17733,N_17425);
and U23210 (N_23210,N_19426,N_15341);
nand U23211 (N_23211,N_17246,N_18820);
and U23212 (N_23212,N_17422,N_19645);
and U23213 (N_23213,N_19091,N_19859);
and U23214 (N_23214,N_18025,N_17095);
or U23215 (N_23215,N_16984,N_17654);
nor U23216 (N_23216,N_15090,N_19200);
or U23217 (N_23217,N_18309,N_15104);
nand U23218 (N_23218,N_17622,N_15920);
or U23219 (N_23219,N_15420,N_16918);
xnor U23220 (N_23220,N_15815,N_19002);
and U23221 (N_23221,N_17715,N_16439);
nand U23222 (N_23222,N_15170,N_19102);
xor U23223 (N_23223,N_19700,N_16792);
or U23224 (N_23224,N_16966,N_15176);
and U23225 (N_23225,N_17835,N_18495);
and U23226 (N_23226,N_16556,N_16198);
nor U23227 (N_23227,N_19313,N_19624);
and U23228 (N_23228,N_17597,N_18973);
or U23229 (N_23229,N_16940,N_19424);
and U23230 (N_23230,N_15975,N_16697);
xnor U23231 (N_23231,N_17588,N_16398);
nor U23232 (N_23232,N_15920,N_19499);
or U23233 (N_23233,N_18186,N_18295);
or U23234 (N_23234,N_17502,N_17114);
and U23235 (N_23235,N_15075,N_17924);
or U23236 (N_23236,N_17035,N_18633);
or U23237 (N_23237,N_16589,N_19405);
nor U23238 (N_23238,N_18777,N_18413);
nor U23239 (N_23239,N_17260,N_18310);
and U23240 (N_23240,N_16563,N_19475);
nor U23241 (N_23241,N_19951,N_17994);
or U23242 (N_23242,N_19031,N_16358);
or U23243 (N_23243,N_18202,N_16189);
or U23244 (N_23244,N_17224,N_18575);
or U23245 (N_23245,N_16515,N_16974);
nor U23246 (N_23246,N_19291,N_15450);
nor U23247 (N_23247,N_17946,N_16090);
or U23248 (N_23248,N_15058,N_18768);
nand U23249 (N_23249,N_15055,N_16936);
xnor U23250 (N_23250,N_17360,N_15607);
xnor U23251 (N_23251,N_17934,N_18054);
nor U23252 (N_23252,N_19964,N_18983);
and U23253 (N_23253,N_16855,N_15456);
and U23254 (N_23254,N_17693,N_16331);
and U23255 (N_23255,N_19561,N_18765);
or U23256 (N_23256,N_16520,N_16677);
nor U23257 (N_23257,N_18352,N_18912);
and U23258 (N_23258,N_17080,N_17653);
and U23259 (N_23259,N_19233,N_17192);
nor U23260 (N_23260,N_16078,N_19324);
nand U23261 (N_23261,N_19027,N_18771);
nor U23262 (N_23262,N_16586,N_19726);
and U23263 (N_23263,N_18815,N_18992);
xor U23264 (N_23264,N_18673,N_17179);
and U23265 (N_23265,N_17581,N_16134);
and U23266 (N_23266,N_18799,N_18834);
and U23267 (N_23267,N_15118,N_18040);
nand U23268 (N_23268,N_15572,N_19767);
nor U23269 (N_23269,N_17472,N_17336);
nand U23270 (N_23270,N_15512,N_16851);
and U23271 (N_23271,N_15135,N_15571);
and U23272 (N_23272,N_18561,N_19501);
nor U23273 (N_23273,N_18953,N_17473);
and U23274 (N_23274,N_19935,N_16624);
and U23275 (N_23275,N_16946,N_16133);
or U23276 (N_23276,N_18918,N_15523);
nand U23277 (N_23277,N_18393,N_16181);
or U23278 (N_23278,N_17507,N_15721);
and U23279 (N_23279,N_18708,N_16055);
xnor U23280 (N_23280,N_19136,N_18395);
nor U23281 (N_23281,N_15812,N_17422);
nand U23282 (N_23282,N_15852,N_18624);
or U23283 (N_23283,N_16799,N_16498);
or U23284 (N_23284,N_17124,N_17776);
nand U23285 (N_23285,N_18118,N_19037);
nor U23286 (N_23286,N_16153,N_17182);
nand U23287 (N_23287,N_19893,N_18469);
nand U23288 (N_23288,N_15539,N_15234);
xor U23289 (N_23289,N_17319,N_17008);
or U23290 (N_23290,N_19391,N_15686);
or U23291 (N_23291,N_18511,N_15297);
nor U23292 (N_23292,N_17163,N_17193);
or U23293 (N_23293,N_19647,N_18532);
xnor U23294 (N_23294,N_15855,N_18967);
nor U23295 (N_23295,N_15383,N_19379);
and U23296 (N_23296,N_16516,N_16988);
and U23297 (N_23297,N_15274,N_16196);
or U23298 (N_23298,N_17802,N_17239);
nand U23299 (N_23299,N_17970,N_19442);
and U23300 (N_23300,N_19281,N_17815);
nor U23301 (N_23301,N_15472,N_17704);
xnor U23302 (N_23302,N_19323,N_15732);
or U23303 (N_23303,N_15614,N_15302);
nor U23304 (N_23304,N_18532,N_18594);
and U23305 (N_23305,N_16038,N_19719);
nand U23306 (N_23306,N_16186,N_18205);
xor U23307 (N_23307,N_15586,N_17539);
or U23308 (N_23308,N_19101,N_17683);
xor U23309 (N_23309,N_17002,N_15777);
nand U23310 (N_23310,N_18812,N_18529);
nor U23311 (N_23311,N_18984,N_19097);
xnor U23312 (N_23312,N_16725,N_17238);
and U23313 (N_23313,N_15393,N_16833);
and U23314 (N_23314,N_16409,N_17226);
and U23315 (N_23315,N_17031,N_16683);
and U23316 (N_23316,N_18247,N_15703);
or U23317 (N_23317,N_17690,N_18686);
and U23318 (N_23318,N_19098,N_16449);
nand U23319 (N_23319,N_19364,N_15993);
nand U23320 (N_23320,N_17395,N_17764);
nand U23321 (N_23321,N_18907,N_16691);
or U23322 (N_23322,N_19201,N_17575);
nor U23323 (N_23323,N_17738,N_16902);
and U23324 (N_23324,N_18393,N_15365);
or U23325 (N_23325,N_18591,N_16506);
or U23326 (N_23326,N_16777,N_15339);
and U23327 (N_23327,N_18117,N_18744);
or U23328 (N_23328,N_17316,N_17399);
nand U23329 (N_23329,N_16158,N_18184);
and U23330 (N_23330,N_16396,N_15291);
xnor U23331 (N_23331,N_16364,N_15915);
nor U23332 (N_23332,N_19970,N_17136);
and U23333 (N_23333,N_15820,N_15143);
nor U23334 (N_23334,N_15159,N_18292);
xnor U23335 (N_23335,N_19328,N_15061);
nor U23336 (N_23336,N_19751,N_17618);
or U23337 (N_23337,N_17052,N_19621);
nand U23338 (N_23338,N_17076,N_18848);
and U23339 (N_23339,N_17670,N_16562);
or U23340 (N_23340,N_17026,N_17665);
and U23341 (N_23341,N_15951,N_18495);
nor U23342 (N_23342,N_15578,N_15120);
and U23343 (N_23343,N_17741,N_16079);
nor U23344 (N_23344,N_16548,N_17972);
or U23345 (N_23345,N_17579,N_16148);
nor U23346 (N_23346,N_16469,N_15600);
and U23347 (N_23347,N_15307,N_15381);
nand U23348 (N_23348,N_17926,N_18623);
nor U23349 (N_23349,N_18988,N_19991);
nor U23350 (N_23350,N_19994,N_17818);
nor U23351 (N_23351,N_16431,N_19713);
or U23352 (N_23352,N_17956,N_16286);
or U23353 (N_23353,N_15994,N_16331);
and U23354 (N_23354,N_19693,N_19412);
and U23355 (N_23355,N_18274,N_18719);
xor U23356 (N_23356,N_17140,N_17744);
or U23357 (N_23357,N_15092,N_16796);
nor U23358 (N_23358,N_15385,N_17826);
or U23359 (N_23359,N_18058,N_17910);
nor U23360 (N_23360,N_15985,N_16060);
nand U23361 (N_23361,N_15439,N_18257);
or U23362 (N_23362,N_16787,N_16775);
xnor U23363 (N_23363,N_18757,N_19279);
nor U23364 (N_23364,N_17894,N_17149);
nor U23365 (N_23365,N_16210,N_15357);
nand U23366 (N_23366,N_16784,N_17809);
nor U23367 (N_23367,N_16941,N_18105);
or U23368 (N_23368,N_17028,N_15968);
or U23369 (N_23369,N_17806,N_16446);
nor U23370 (N_23370,N_18850,N_19661);
nand U23371 (N_23371,N_18194,N_18349);
nand U23372 (N_23372,N_16849,N_19662);
nor U23373 (N_23373,N_15432,N_15365);
and U23374 (N_23374,N_16138,N_18428);
xor U23375 (N_23375,N_19618,N_19854);
and U23376 (N_23376,N_18815,N_17128);
xnor U23377 (N_23377,N_18839,N_18815);
nand U23378 (N_23378,N_16318,N_16615);
nand U23379 (N_23379,N_17777,N_19738);
and U23380 (N_23380,N_17391,N_17865);
or U23381 (N_23381,N_16308,N_17826);
or U23382 (N_23382,N_19113,N_18081);
and U23383 (N_23383,N_18089,N_19427);
and U23384 (N_23384,N_17940,N_17755);
and U23385 (N_23385,N_17247,N_17119);
nand U23386 (N_23386,N_18298,N_19511);
nor U23387 (N_23387,N_17141,N_18404);
nand U23388 (N_23388,N_18976,N_17480);
and U23389 (N_23389,N_15376,N_17332);
nor U23390 (N_23390,N_18598,N_19138);
or U23391 (N_23391,N_16015,N_19284);
nor U23392 (N_23392,N_15736,N_18341);
nand U23393 (N_23393,N_16075,N_16023);
and U23394 (N_23394,N_19557,N_15185);
or U23395 (N_23395,N_16824,N_16788);
and U23396 (N_23396,N_18810,N_17081);
nor U23397 (N_23397,N_18555,N_16171);
and U23398 (N_23398,N_15872,N_19690);
nand U23399 (N_23399,N_16939,N_19408);
or U23400 (N_23400,N_15198,N_18973);
nand U23401 (N_23401,N_17674,N_18609);
or U23402 (N_23402,N_15530,N_15393);
and U23403 (N_23403,N_18802,N_15182);
or U23404 (N_23404,N_16300,N_18614);
or U23405 (N_23405,N_16926,N_19381);
xor U23406 (N_23406,N_17245,N_17478);
nor U23407 (N_23407,N_17843,N_15058);
or U23408 (N_23408,N_19021,N_19378);
xor U23409 (N_23409,N_16032,N_15121);
or U23410 (N_23410,N_19218,N_17343);
and U23411 (N_23411,N_16033,N_17866);
nand U23412 (N_23412,N_19578,N_18649);
xor U23413 (N_23413,N_18750,N_19442);
or U23414 (N_23414,N_15228,N_17817);
nand U23415 (N_23415,N_15094,N_18084);
nand U23416 (N_23416,N_16636,N_15343);
nand U23417 (N_23417,N_19443,N_18046);
and U23418 (N_23418,N_15655,N_15255);
or U23419 (N_23419,N_19950,N_15338);
or U23420 (N_23420,N_18136,N_17764);
or U23421 (N_23421,N_18811,N_15787);
or U23422 (N_23422,N_17339,N_18797);
or U23423 (N_23423,N_19527,N_15916);
and U23424 (N_23424,N_15833,N_16130);
nand U23425 (N_23425,N_18228,N_17394);
nand U23426 (N_23426,N_19938,N_19015);
and U23427 (N_23427,N_18067,N_19908);
nand U23428 (N_23428,N_16987,N_16676);
nor U23429 (N_23429,N_17435,N_19214);
or U23430 (N_23430,N_16650,N_17817);
or U23431 (N_23431,N_17247,N_17521);
nor U23432 (N_23432,N_16737,N_19597);
or U23433 (N_23433,N_16689,N_17202);
and U23434 (N_23434,N_16711,N_17606);
xnor U23435 (N_23435,N_16117,N_17419);
or U23436 (N_23436,N_16465,N_15764);
and U23437 (N_23437,N_18769,N_18639);
or U23438 (N_23438,N_16208,N_19537);
xnor U23439 (N_23439,N_18682,N_16835);
nor U23440 (N_23440,N_17309,N_16598);
nor U23441 (N_23441,N_19136,N_19121);
xnor U23442 (N_23442,N_16116,N_19934);
nand U23443 (N_23443,N_16081,N_17589);
or U23444 (N_23444,N_17266,N_18594);
and U23445 (N_23445,N_19169,N_15204);
xor U23446 (N_23446,N_16686,N_18233);
nand U23447 (N_23447,N_17564,N_17453);
and U23448 (N_23448,N_16531,N_17318);
and U23449 (N_23449,N_16058,N_16520);
nand U23450 (N_23450,N_16900,N_17033);
nor U23451 (N_23451,N_17862,N_15220);
or U23452 (N_23452,N_16874,N_19714);
or U23453 (N_23453,N_18206,N_19255);
and U23454 (N_23454,N_16129,N_17667);
nand U23455 (N_23455,N_19793,N_16439);
and U23456 (N_23456,N_16422,N_18681);
and U23457 (N_23457,N_16443,N_19601);
and U23458 (N_23458,N_18359,N_19738);
nor U23459 (N_23459,N_17816,N_17210);
nand U23460 (N_23460,N_15578,N_16271);
or U23461 (N_23461,N_16846,N_16671);
and U23462 (N_23462,N_18720,N_17646);
nor U23463 (N_23463,N_16412,N_19613);
or U23464 (N_23464,N_16863,N_15275);
nand U23465 (N_23465,N_18463,N_15939);
or U23466 (N_23466,N_17904,N_17033);
nor U23467 (N_23467,N_15563,N_17429);
or U23468 (N_23468,N_19463,N_18170);
nand U23469 (N_23469,N_15324,N_18559);
nand U23470 (N_23470,N_18883,N_15946);
xor U23471 (N_23471,N_15628,N_17810);
nand U23472 (N_23472,N_19625,N_19428);
xnor U23473 (N_23473,N_16936,N_19992);
nand U23474 (N_23474,N_17212,N_18771);
and U23475 (N_23475,N_16219,N_16664);
nor U23476 (N_23476,N_15705,N_19755);
or U23477 (N_23477,N_18360,N_16814);
nor U23478 (N_23478,N_15348,N_19045);
or U23479 (N_23479,N_15142,N_15895);
and U23480 (N_23480,N_16303,N_17391);
nand U23481 (N_23481,N_19892,N_19304);
nand U23482 (N_23482,N_16835,N_17842);
or U23483 (N_23483,N_17228,N_19074);
xnor U23484 (N_23484,N_17878,N_19369);
nand U23485 (N_23485,N_17345,N_15935);
nand U23486 (N_23486,N_19409,N_18424);
xnor U23487 (N_23487,N_15964,N_16730);
or U23488 (N_23488,N_15079,N_19151);
or U23489 (N_23489,N_15019,N_16054);
or U23490 (N_23490,N_16852,N_15647);
or U23491 (N_23491,N_17567,N_19998);
nand U23492 (N_23492,N_16650,N_15964);
nand U23493 (N_23493,N_15954,N_16540);
xor U23494 (N_23494,N_16715,N_18838);
and U23495 (N_23495,N_17029,N_16663);
xnor U23496 (N_23496,N_15387,N_16191);
nor U23497 (N_23497,N_15436,N_15831);
nor U23498 (N_23498,N_18849,N_15172);
and U23499 (N_23499,N_19832,N_18642);
or U23500 (N_23500,N_19205,N_15363);
or U23501 (N_23501,N_18079,N_15027);
xnor U23502 (N_23502,N_16016,N_16174);
nand U23503 (N_23503,N_16610,N_19996);
nor U23504 (N_23504,N_18097,N_19026);
or U23505 (N_23505,N_17629,N_19469);
nand U23506 (N_23506,N_19276,N_17421);
nand U23507 (N_23507,N_15325,N_19991);
and U23508 (N_23508,N_15751,N_16381);
nor U23509 (N_23509,N_16287,N_16912);
nand U23510 (N_23510,N_15047,N_17402);
and U23511 (N_23511,N_16568,N_17357);
xnor U23512 (N_23512,N_17845,N_16367);
or U23513 (N_23513,N_16177,N_16330);
nand U23514 (N_23514,N_16383,N_17707);
nand U23515 (N_23515,N_19615,N_16449);
nand U23516 (N_23516,N_16557,N_19073);
or U23517 (N_23517,N_19025,N_19686);
nand U23518 (N_23518,N_18959,N_18464);
nor U23519 (N_23519,N_15638,N_17591);
nor U23520 (N_23520,N_15713,N_19273);
and U23521 (N_23521,N_17910,N_19057);
nor U23522 (N_23522,N_15408,N_15619);
nor U23523 (N_23523,N_18287,N_16883);
nand U23524 (N_23524,N_18842,N_18961);
or U23525 (N_23525,N_18551,N_19423);
nor U23526 (N_23526,N_18752,N_18985);
xor U23527 (N_23527,N_17398,N_17326);
and U23528 (N_23528,N_16391,N_16473);
and U23529 (N_23529,N_16004,N_19742);
nor U23530 (N_23530,N_15940,N_18754);
nor U23531 (N_23531,N_17387,N_18851);
nor U23532 (N_23532,N_16594,N_15294);
xor U23533 (N_23533,N_15126,N_16326);
nor U23534 (N_23534,N_18017,N_18372);
nor U23535 (N_23535,N_18926,N_19666);
and U23536 (N_23536,N_15008,N_15228);
and U23537 (N_23537,N_17513,N_15062);
nand U23538 (N_23538,N_19016,N_17709);
and U23539 (N_23539,N_18560,N_18213);
xor U23540 (N_23540,N_15147,N_17683);
and U23541 (N_23541,N_16790,N_18321);
or U23542 (N_23542,N_16403,N_15007);
and U23543 (N_23543,N_17438,N_17003);
xnor U23544 (N_23544,N_18669,N_19896);
and U23545 (N_23545,N_15815,N_18244);
nand U23546 (N_23546,N_19888,N_19177);
and U23547 (N_23547,N_15154,N_18460);
and U23548 (N_23548,N_15459,N_16445);
nand U23549 (N_23549,N_16272,N_16373);
nor U23550 (N_23550,N_17141,N_18626);
nor U23551 (N_23551,N_16961,N_19504);
nor U23552 (N_23552,N_18478,N_17356);
or U23553 (N_23553,N_17062,N_15785);
xor U23554 (N_23554,N_19442,N_15134);
and U23555 (N_23555,N_17595,N_16152);
nor U23556 (N_23556,N_15359,N_16887);
nand U23557 (N_23557,N_15459,N_16468);
xnor U23558 (N_23558,N_16772,N_17260);
or U23559 (N_23559,N_16601,N_18643);
nand U23560 (N_23560,N_19256,N_19479);
and U23561 (N_23561,N_17924,N_19911);
and U23562 (N_23562,N_16233,N_19411);
or U23563 (N_23563,N_16055,N_16676);
nor U23564 (N_23564,N_15071,N_18198);
and U23565 (N_23565,N_16564,N_17401);
and U23566 (N_23566,N_15139,N_19326);
nand U23567 (N_23567,N_15703,N_16351);
or U23568 (N_23568,N_15519,N_16272);
or U23569 (N_23569,N_17820,N_19719);
nand U23570 (N_23570,N_15099,N_15113);
or U23571 (N_23571,N_16607,N_15409);
and U23572 (N_23572,N_15548,N_18760);
or U23573 (N_23573,N_17304,N_16720);
nand U23574 (N_23574,N_17212,N_18706);
nor U23575 (N_23575,N_18585,N_17788);
and U23576 (N_23576,N_15999,N_19362);
and U23577 (N_23577,N_16647,N_18657);
or U23578 (N_23578,N_16016,N_16843);
and U23579 (N_23579,N_19613,N_17373);
nand U23580 (N_23580,N_18452,N_19531);
and U23581 (N_23581,N_15277,N_15450);
nor U23582 (N_23582,N_17758,N_15245);
and U23583 (N_23583,N_15038,N_16382);
xor U23584 (N_23584,N_17825,N_19766);
nor U23585 (N_23585,N_16568,N_19433);
or U23586 (N_23586,N_15615,N_19239);
and U23587 (N_23587,N_18178,N_16556);
nand U23588 (N_23588,N_15262,N_19202);
and U23589 (N_23589,N_15692,N_19136);
nand U23590 (N_23590,N_18018,N_15529);
nor U23591 (N_23591,N_19276,N_15179);
nor U23592 (N_23592,N_17694,N_15343);
nand U23593 (N_23593,N_16087,N_19105);
nand U23594 (N_23594,N_18695,N_17596);
nor U23595 (N_23595,N_17007,N_19646);
nor U23596 (N_23596,N_19681,N_19772);
or U23597 (N_23597,N_15355,N_17153);
or U23598 (N_23598,N_18336,N_18714);
and U23599 (N_23599,N_18434,N_19300);
nand U23600 (N_23600,N_19114,N_16961);
or U23601 (N_23601,N_18821,N_17849);
and U23602 (N_23602,N_19605,N_18765);
and U23603 (N_23603,N_17442,N_18805);
xor U23604 (N_23604,N_17724,N_17155);
nand U23605 (N_23605,N_16742,N_19730);
or U23606 (N_23606,N_15868,N_18115);
nor U23607 (N_23607,N_16147,N_15316);
nand U23608 (N_23608,N_15661,N_16247);
nand U23609 (N_23609,N_18373,N_16264);
or U23610 (N_23610,N_18845,N_18263);
or U23611 (N_23611,N_19772,N_16734);
or U23612 (N_23612,N_16917,N_18368);
or U23613 (N_23613,N_15423,N_16615);
nand U23614 (N_23614,N_15168,N_17819);
nor U23615 (N_23615,N_18969,N_18209);
nor U23616 (N_23616,N_18743,N_17130);
and U23617 (N_23617,N_18571,N_15285);
and U23618 (N_23618,N_15912,N_15839);
nand U23619 (N_23619,N_16853,N_17184);
nor U23620 (N_23620,N_15144,N_19754);
nand U23621 (N_23621,N_16874,N_18381);
nor U23622 (N_23622,N_16653,N_15170);
and U23623 (N_23623,N_19328,N_17750);
xnor U23624 (N_23624,N_17115,N_19413);
nand U23625 (N_23625,N_19399,N_17187);
or U23626 (N_23626,N_15153,N_19380);
xnor U23627 (N_23627,N_19379,N_19753);
xor U23628 (N_23628,N_19849,N_15241);
nand U23629 (N_23629,N_15604,N_19677);
or U23630 (N_23630,N_19760,N_18331);
or U23631 (N_23631,N_16566,N_17311);
nand U23632 (N_23632,N_15196,N_17488);
xor U23633 (N_23633,N_16982,N_15507);
nand U23634 (N_23634,N_19134,N_15921);
nand U23635 (N_23635,N_19161,N_15033);
and U23636 (N_23636,N_15863,N_16685);
or U23637 (N_23637,N_16939,N_15302);
nor U23638 (N_23638,N_15642,N_15670);
or U23639 (N_23639,N_18639,N_19225);
and U23640 (N_23640,N_18661,N_16912);
nand U23641 (N_23641,N_15356,N_18793);
xnor U23642 (N_23642,N_16590,N_17247);
nand U23643 (N_23643,N_17641,N_15951);
nor U23644 (N_23644,N_15456,N_19504);
or U23645 (N_23645,N_18436,N_18172);
or U23646 (N_23646,N_15577,N_18038);
and U23647 (N_23647,N_16293,N_19196);
nand U23648 (N_23648,N_19285,N_17869);
or U23649 (N_23649,N_19347,N_18660);
xor U23650 (N_23650,N_15595,N_17785);
or U23651 (N_23651,N_18813,N_15510);
nor U23652 (N_23652,N_17147,N_18332);
and U23653 (N_23653,N_15377,N_16335);
xor U23654 (N_23654,N_19927,N_18590);
and U23655 (N_23655,N_18884,N_19459);
or U23656 (N_23656,N_18665,N_19628);
or U23657 (N_23657,N_16065,N_19199);
nand U23658 (N_23658,N_15477,N_18749);
and U23659 (N_23659,N_15446,N_19895);
and U23660 (N_23660,N_17086,N_18848);
and U23661 (N_23661,N_17373,N_19866);
nor U23662 (N_23662,N_17138,N_19812);
and U23663 (N_23663,N_15304,N_15648);
nor U23664 (N_23664,N_18930,N_16624);
nor U23665 (N_23665,N_16284,N_18157);
xor U23666 (N_23666,N_15107,N_18839);
and U23667 (N_23667,N_19367,N_15711);
xor U23668 (N_23668,N_19642,N_19622);
xnor U23669 (N_23669,N_15457,N_16704);
nor U23670 (N_23670,N_17394,N_18248);
or U23671 (N_23671,N_18051,N_17194);
nand U23672 (N_23672,N_16668,N_17267);
xnor U23673 (N_23673,N_16035,N_17546);
and U23674 (N_23674,N_18003,N_18453);
xor U23675 (N_23675,N_17345,N_16474);
nor U23676 (N_23676,N_17598,N_15690);
nand U23677 (N_23677,N_19090,N_17334);
nor U23678 (N_23678,N_16875,N_17275);
xnor U23679 (N_23679,N_16357,N_15505);
nand U23680 (N_23680,N_16722,N_15272);
and U23681 (N_23681,N_17249,N_18575);
or U23682 (N_23682,N_18029,N_17131);
nor U23683 (N_23683,N_18048,N_16231);
and U23684 (N_23684,N_17445,N_16400);
xor U23685 (N_23685,N_17470,N_16590);
or U23686 (N_23686,N_19406,N_18061);
xnor U23687 (N_23687,N_16938,N_18442);
and U23688 (N_23688,N_18558,N_19036);
nand U23689 (N_23689,N_18466,N_17825);
or U23690 (N_23690,N_19682,N_15091);
or U23691 (N_23691,N_18644,N_16315);
nand U23692 (N_23692,N_18857,N_18538);
or U23693 (N_23693,N_17417,N_19190);
or U23694 (N_23694,N_17235,N_15277);
nor U23695 (N_23695,N_15395,N_19202);
nor U23696 (N_23696,N_16853,N_16333);
nand U23697 (N_23697,N_16071,N_18670);
nand U23698 (N_23698,N_17801,N_16768);
and U23699 (N_23699,N_18845,N_16556);
nor U23700 (N_23700,N_18572,N_15560);
or U23701 (N_23701,N_19644,N_15180);
nor U23702 (N_23702,N_19513,N_15467);
nor U23703 (N_23703,N_16434,N_19576);
xor U23704 (N_23704,N_18909,N_18464);
nor U23705 (N_23705,N_18971,N_19307);
nand U23706 (N_23706,N_19258,N_19130);
and U23707 (N_23707,N_16540,N_16311);
and U23708 (N_23708,N_15471,N_18650);
and U23709 (N_23709,N_15753,N_15928);
and U23710 (N_23710,N_16410,N_17889);
nand U23711 (N_23711,N_16287,N_18357);
nand U23712 (N_23712,N_18116,N_19432);
nand U23713 (N_23713,N_17757,N_19436);
nor U23714 (N_23714,N_17451,N_16480);
and U23715 (N_23715,N_18449,N_17282);
nand U23716 (N_23716,N_16986,N_17579);
nand U23717 (N_23717,N_19278,N_16804);
xor U23718 (N_23718,N_16000,N_15101);
or U23719 (N_23719,N_19952,N_15521);
nor U23720 (N_23720,N_17102,N_15642);
nand U23721 (N_23721,N_19976,N_19990);
nor U23722 (N_23722,N_15811,N_19905);
xnor U23723 (N_23723,N_17154,N_16298);
xnor U23724 (N_23724,N_15118,N_19341);
nand U23725 (N_23725,N_18627,N_17615);
nor U23726 (N_23726,N_16722,N_17053);
nor U23727 (N_23727,N_17228,N_15573);
nand U23728 (N_23728,N_19198,N_18743);
xor U23729 (N_23729,N_18813,N_15132);
nor U23730 (N_23730,N_18055,N_18703);
nor U23731 (N_23731,N_18091,N_18137);
and U23732 (N_23732,N_16054,N_16886);
and U23733 (N_23733,N_19796,N_19762);
nand U23734 (N_23734,N_19525,N_17282);
or U23735 (N_23735,N_15972,N_17245);
nor U23736 (N_23736,N_19171,N_17666);
or U23737 (N_23737,N_19915,N_17249);
or U23738 (N_23738,N_18335,N_18331);
nor U23739 (N_23739,N_17129,N_18402);
nand U23740 (N_23740,N_15723,N_16639);
or U23741 (N_23741,N_19537,N_17247);
nand U23742 (N_23742,N_17384,N_17802);
nor U23743 (N_23743,N_15209,N_18862);
nor U23744 (N_23744,N_17225,N_18359);
or U23745 (N_23745,N_19344,N_18126);
or U23746 (N_23746,N_15906,N_17860);
nor U23747 (N_23747,N_19823,N_19260);
nor U23748 (N_23748,N_16424,N_19554);
nor U23749 (N_23749,N_17994,N_16041);
or U23750 (N_23750,N_18011,N_15490);
and U23751 (N_23751,N_15212,N_19828);
or U23752 (N_23752,N_18601,N_17815);
nand U23753 (N_23753,N_16489,N_15729);
xor U23754 (N_23754,N_15211,N_15201);
or U23755 (N_23755,N_18979,N_19091);
nand U23756 (N_23756,N_15208,N_17093);
or U23757 (N_23757,N_15458,N_16588);
nand U23758 (N_23758,N_19300,N_17047);
nor U23759 (N_23759,N_17266,N_17228);
nand U23760 (N_23760,N_16033,N_15497);
nand U23761 (N_23761,N_15409,N_19727);
nand U23762 (N_23762,N_16315,N_15329);
nor U23763 (N_23763,N_17502,N_18440);
nor U23764 (N_23764,N_19816,N_16580);
xor U23765 (N_23765,N_18126,N_15264);
nand U23766 (N_23766,N_15005,N_17438);
nor U23767 (N_23767,N_17515,N_15605);
or U23768 (N_23768,N_16617,N_16379);
nand U23769 (N_23769,N_15325,N_17679);
nor U23770 (N_23770,N_18911,N_18218);
nand U23771 (N_23771,N_19163,N_19950);
nand U23772 (N_23772,N_19887,N_18659);
nand U23773 (N_23773,N_15978,N_19579);
and U23774 (N_23774,N_19790,N_17422);
and U23775 (N_23775,N_17782,N_19207);
or U23776 (N_23776,N_18497,N_16578);
nand U23777 (N_23777,N_19845,N_19561);
nor U23778 (N_23778,N_15077,N_15751);
and U23779 (N_23779,N_19556,N_16716);
xnor U23780 (N_23780,N_19155,N_15949);
or U23781 (N_23781,N_19718,N_16619);
and U23782 (N_23782,N_19543,N_16259);
nand U23783 (N_23783,N_17062,N_18822);
nor U23784 (N_23784,N_17066,N_18726);
nor U23785 (N_23785,N_17396,N_15951);
nand U23786 (N_23786,N_16455,N_17889);
xor U23787 (N_23787,N_18318,N_16973);
xor U23788 (N_23788,N_17235,N_17572);
and U23789 (N_23789,N_18498,N_16989);
or U23790 (N_23790,N_17011,N_16246);
nand U23791 (N_23791,N_16327,N_19829);
nor U23792 (N_23792,N_15539,N_18532);
or U23793 (N_23793,N_16155,N_17515);
nor U23794 (N_23794,N_19214,N_16077);
and U23795 (N_23795,N_17038,N_17311);
nor U23796 (N_23796,N_19195,N_15474);
xnor U23797 (N_23797,N_17598,N_15768);
or U23798 (N_23798,N_16803,N_16892);
and U23799 (N_23799,N_15423,N_18694);
nor U23800 (N_23800,N_16536,N_19543);
nor U23801 (N_23801,N_16264,N_15553);
and U23802 (N_23802,N_16777,N_16788);
nand U23803 (N_23803,N_15939,N_15010);
nand U23804 (N_23804,N_15406,N_15262);
and U23805 (N_23805,N_18590,N_18786);
nand U23806 (N_23806,N_15413,N_17854);
nand U23807 (N_23807,N_17056,N_16101);
or U23808 (N_23808,N_16211,N_18774);
nor U23809 (N_23809,N_18982,N_16597);
or U23810 (N_23810,N_19389,N_17106);
and U23811 (N_23811,N_19133,N_19530);
or U23812 (N_23812,N_15028,N_15427);
nand U23813 (N_23813,N_16138,N_17817);
nor U23814 (N_23814,N_18572,N_17330);
or U23815 (N_23815,N_19081,N_15909);
nand U23816 (N_23816,N_18154,N_19170);
and U23817 (N_23817,N_18823,N_16910);
nor U23818 (N_23818,N_18944,N_19807);
or U23819 (N_23819,N_17290,N_15536);
xnor U23820 (N_23820,N_18504,N_15728);
or U23821 (N_23821,N_17921,N_16834);
or U23822 (N_23822,N_19421,N_17401);
and U23823 (N_23823,N_16222,N_16323);
nand U23824 (N_23824,N_16559,N_16000);
xnor U23825 (N_23825,N_16889,N_16805);
nand U23826 (N_23826,N_18989,N_16403);
xor U23827 (N_23827,N_15020,N_15585);
and U23828 (N_23828,N_19817,N_15137);
nand U23829 (N_23829,N_19567,N_19486);
nor U23830 (N_23830,N_18618,N_17833);
and U23831 (N_23831,N_15388,N_16373);
or U23832 (N_23832,N_15691,N_16956);
and U23833 (N_23833,N_17231,N_16212);
nand U23834 (N_23834,N_16871,N_16026);
nand U23835 (N_23835,N_15295,N_17662);
or U23836 (N_23836,N_19199,N_16705);
xor U23837 (N_23837,N_19049,N_19149);
or U23838 (N_23838,N_16111,N_19806);
or U23839 (N_23839,N_17774,N_19177);
nor U23840 (N_23840,N_19615,N_19107);
or U23841 (N_23841,N_16042,N_19177);
nand U23842 (N_23842,N_18337,N_18232);
xnor U23843 (N_23843,N_19065,N_15093);
nand U23844 (N_23844,N_16124,N_17369);
or U23845 (N_23845,N_18532,N_18109);
and U23846 (N_23846,N_18894,N_16014);
and U23847 (N_23847,N_19967,N_19537);
nand U23848 (N_23848,N_19769,N_15044);
and U23849 (N_23849,N_18953,N_15500);
or U23850 (N_23850,N_19245,N_19643);
nand U23851 (N_23851,N_18017,N_15448);
nand U23852 (N_23852,N_19082,N_15586);
nor U23853 (N_23853,N_16504,N_16323);
nand U23854 (N_23854,N_19313,N_16871);
and U23855 (N_23855,N_16653,N_17979);
nand U23856 (N_23856,N_17243,N_16534);
and U23857 (N_23857,N_19716,N_15597);
nand U23858 (N_23858,N_15203,N_17947);
nor U23859 (N_23859,N_19634,N_18646);
xor U23860 (N_23860,N_18703,N_19968);
nor U23861 (N_23861,N_17359,N_18097);
or U23862 (N_23862,N_18712,N_15746);
or U23863 (N_23863,N_16663,N_18775);
nand U23864 (N_23864,N_15529,N_18800);
nand U23865 (N_23865,N_15153,N_17740);
nand U23866 (N_23866,N_16232,N_17542);
nand U23867 (N_23867,N_17723,N_15041);
nand U23868 (N_23868,N_19720,N_17619);
nand U23869 (N_23869,N_17252,N_17125);
or U23870 (N_23870,N_15182,N_16691);
or U23871 (N_23871,N_18957,N_17131);
nand U23872 (N_23872,N_19152,N_19901);
or U23873 (N_23873,N_18479,N_18990);
or U23874 (N_23874,N_15656,N_18431);
and U23875 (N_23875,N_18290,N_15910);
or U23876 (N_23876,N_17829,N_18840);
nand U23877 (N_23877,N_19976,N_16576);
nor U23878 (N_23878,N_17544,N_17479);
or U23879 (N_23879,N_15135,N_18162);
xor U23880 (N_23880,N_15175,N_17820);
or U23881 (N_23881,N_19075,N_17707);
and U23882 (N_23882,N_15872,N_16280);
nand U23883 (N_23883,N_15382,N_16439);
and U23884 (N_23884,N_18160,N_16485);
and U23885 (N_23885,N_18675,N_17736);
or U23886 (N_23886,N_17400,N_19850);
nor U23887 (N_23887,N_17723,N_16762);
nand U23888 (N_23888,N_19749,N_15165);
nor U23889 (N_23889,N_15559,N_18418);
and U23890 (N_23890,N_19128,N_15329);
xor U23891 (N_23891,N_15307,N_16999);
nor U23892 (N_23892,N_19775,N_16235);
nand U23893 (N_23893,N_17914,N_15588);
and U23894 (N_23894,N_17053,N_19993);
or U23895 (N_23895,N_18918,N_18923);
nor U23896 (N_23896,N_16520,N_17952);
xnor U23897 (N_23897,N_17232,N_18023);
nand U23898 (N_23898,N_15617,N_15494);
xnor U23899 (N_23899,N_15366,N_15382);
nand U23900 (N_23900,N_15340,N_19748);
xnor U23901 (N_23901,N_18707,N_17741);
or U23902 (N_23902,N_15343,N_18815);
and U23903 (N_23903,N_16827,N_18724);
or U23904 (N_23904,N_16000,N_19837);
or U23905 (N_23905,N_17541,N_16281);
and U23906 (N_23906,N_17670,N_17325);
nor U23907 (N_23907,N_18861,N_15244);
nand U23908 (N_23908,N_18601,N_19209);
nand U23909 (N_23909,N_19052,N_15440);
or U23910 (N_23910,N_16274,N_17262);
nor U23911 (N_23911,N_18175,N_19738);
xnor U23912 (N_23912,N_18759,N_16455);
nor U23913 (N_23913,N_19448,N_15108);
nor U23914 (N_23914,N_18194,N_16774);
or U23915 (N_23915,N_16427,N_18050);
nor U23916 (N_23916,N_15413,N_15067);
nand U23917 (N_23917,N_18158,N_15505);
xor U23918 (N_23918,N_15931,N_18568);
or U23919 (N_23919,N_16083,N_18660);
nor U23920 (N_23920,N_15933,N_19744);
nor U23921 (N_23921,N_18844,N_17308);
or U23922 (N_23922,N_19209,N_19712);
and U23923 (N_23923,N_19624,N_17080);
nand U23924 (N_23924,N_18532,N_18494);
nor U23925 (N_23925,N_17063,N_17767);
xnor U23926 (N_23926,N_15450,N_18214);
nor U23927 (N_23927,N_16490,N_16308);
nor U23928 (N_23928,N_18831,N_18959);
nor U23929 (N_23929,N_17148,N_15039);
and U23930 (N_23930,N_17044,N_16968);
nor U23931 (N_23931,N_15386,N_17377);
and U23932 (N_23932,N_18333,N_19968);
and U23933 (N_23933,N_18609,N_15485);
or U23934 (N_23934,N_16380,N_18912);
and U23935 (N_23935,N_19738,N_16380);
and U23936 (N_23936,N_17252,N_19932);
and U23937 (N_23937,N_18049,N_19747);
and U23938 (N_23938,N_19628,N_16949);
and U23939 (N_23939,N_19468,N_16521);
nor U23940 (N_23940,N_19938,N_16149);
or U23941 (N_23941,N_18520,N_16181);
nand U23942 (N_23942,N_17641,N_17886);
xnor U23943 (N_23943,N_16107,N_19575);
nand U23944 (N_23944,N_18363,N_18606);
xor U23945 (N_23945,N_15187,N_15487);
nor U23946 (N_23946,N_16642,N_19542);
nor U23947 (N_23947,N_18104,N_17299);
nor U23948 (N_23948,N_17579,N_15567);
or U23949 (N_23949,N_18754,N_19793);
nand U23950 (N_23950,N_16641,N_17963);
xnor U23951 (N_23951,N_19797,N_19690);
nand U23952 (N_23952,N_16990,N_19406);
nand U23953 (N_23953,N_17647,N_18236);
and U23954 (N_23954,N_16785,N_16557);
nor U23955 (N_23955,N_16686,N_18895);
and U23956 (N_23956,N_19346,N_17183);
or U23957 (N_23957,N_16558,N_15557);
nor U23958 (N_23958,N_19346,N_18018);
xor U23959 (N_23959,N_18671,N_17099);
nand U23960 (N_23960,N_17328,N_17932);
nor U23961 (N_23961,N_17300,N_16578);
xnor U23962 (N_23962,N_16137,N_17834);
nand U23963 (N_23963,N_15827,N_15245);
nor U23964 (N_23964,N_16088,N_16534);
or U23965 (N_23965,N_15518,N_15763);
nand U23966 (N_23966,N_19601,N_18629);
or U23967 (N_23967,N_18022,N_16055);
nor U23968 (N_23968,N_15568,N_17269);
nand U23969 (N_23969,N_17785,N_18160);
nor U23970 (N_23970,N_16921,N_19090);
and U23971 (N_23971,N_16544,N_17738);
and U23972 (N_23972,N_16168,N_15693);
nand U23973 (N_23973,N_19097,N_17638);
or U23974 (N_23974,N_17665,N_18076);
and U23975 (N_23975,N_15223,N_15044);
nand U23976 (N_23976,N_18227,N_18717);
nand U23977 (N_23977,N_15601,N_18092);
and U23978 (N_23978,N_19932,N_19812);
nand U23979 (N_23979,N_17284,N_19591);
and U23980 (N_23980,N_15621,N_17066);
nor U23981 (N_23981,N_17016,N_19283);
nand U23982 (N_23982,N_15305,N_19753);
xor U23983 (N_23983,N_15050,N_19950);
and U23984 (N_23984,N_18153,N_16784);
xor U23985 (N_23985,N_18189,N_17907);
and U23986 (N_23986,N_19134,N_18064);
or U23987 (N_23987,N_16651,N_15239);
and U23988 (N_23988,N_15840,N_17261);
nor U23989 (N_23989,N_16866,N_16474);
xor U23990 (N_23990,N_15505,N_16756);
and U23991 (N_23991,N_17444,N_19785);
nand U23992 (N_23992,N_19679,N_15589);
or U23993 (N_23993,N_19384,N_17143);
and U23994 (N_23994,N_15842,N_19335);
and U23995 (N_23995,N_17716,N_16036);
or U23996 (N_23996,N_19172,N_17288);
nor U23997 (N_23997,N_15857,N_16736);
nor U23998 (N_23998,N_19587,N_16295);
or U23999 (N_23999,N_18285,N_19950);
nand U24000 (N_24000,N_19841,N_16960);
nor U24001 (N_24001,N_18333,N_17208);
or U24002 (N_24002,N_17165,N_17067);
xnor U24003 (N_24003,N_15899,N_16253);
nand U24004 (N_24004,N_19321,N_19922);
nor U24005 (N_24005,N_15788,N_18761);
and U24006 (N_24006,N_17808,N_18861);
and U24007 (N_24007,N_18664,N_17563);
and U24008 (N_24008,N_15415,N_15920);
xor U24009 (N_24009,N_18321,N_17122);
or U24010 (N_24010,N_17520,N_19032);
and U24011 (N_24011,N_18473,N_18388);
nand U24012 (N_24012,N_18816,N_16513);
or U24013 (N_24013,N_16002,N_15081);
or U24014 (N_24014,N_16353,N_16244);
and U24015 (N_24015,N_15204,N_17976);
and U24016 (N_24016,N_16227,N_19148);
nor U24017 (N_24017,N_18864,N_17011);
and U24018 (N_24018,N_18353,N_15017);
xor U24019 (N_24019,N_19306,N_18401);
xor U24020 (N_24020,N_17936,N_16173);
xnor U24021 (N_24021,N_18041,N_16841);
nor U24022 (N_24022,N_16574,N_17392);
nand U24023 (N_24023,N_16625,N_19820);
nand U24024 (N_24024,N_19842,N_16140);
nand U24025 (N_24025,N_16266,N_17202);
nand U24026 (N_24026,N_19173,N_16682);
and U24027 (N_24027,N_19295,N_15984);
or U24028 (N_24028,N_16091,N_16217);
nand U24029 (N_24029,N_15165,N_16342);
nor U24030 (N_24030,N_15956,N_17588);
or U24031 (N_24031,N_17448,N_19300);
or U24032 (N_24032,N_17104,N_18288);
nor U24033 (N_24033,N_19150,N_15795);
nor U24034 (N_24034,N_19556,N_15383);
nor U24035 (N_24035,N_19622,N_18079);
xnor U24036 (N_24036,N_19315,N_15982);
and U24037 (N_24037,N_15620,N_19217);
and U24038 (N_24038,N_15441,N_18739);
and U24039 (N_24039,N_15003,N_17651);
and U24040 (N_24040,N_17519,N_17762);
nand U24041 (N_24041,N_15142,N_15492);
nand U24042 (N_24042,N_17883,N_15508);
and U24043 (N_24043,N_15369,N_15772);
nor U24044 (N_24044,N_17860,N_16162);
nor U24045 (N_24045,N_18286,N_16470);
nand U24046 (N_24046,N_19641,N_16230);
nor U24047 (N_24047,N_15597,N_15436);
nand U24048 (N_24048,N_18593,N_16075);
nand U24049 (N_24049,N_15759,N_19210);
and U24050 (N_24050,N_15008,N_15583);
nand U24051 (N_24051,N_18004,N_19494);
nand U24052 (N_24052,N_18494,N_15675);
nand U24053 (N_24053,N_17285,N_16734);
and U24054 (N_24054,N_15970,N_16172);
xnor U24055 (N_24055,N_15075,N_19264);
nor U24056 (N_24056,N_16773,N_16052);
nand U24057 (N_24057,N_18358,N_17228);
or U24058 (N_24058,N_18679,N_17923);
nand U24059 (N_24059,N_16759,N_16069);
or U24060 (N_24060,N_17800,N_19220);
nand U24061 (N_24061,N_18780,N_16884);
and U24062 (N_24062,N_18022,N_16814);
nor U24063 (N_24063,N_16701,N_16755);
nor U24064 (N_24064,N_19599,N_17830);
nand U24065 (N_24065,N_18272,N_16985);
and U24066 (N_24066,N_17900,N_16778);
xnor U24067 (N_24067,N_19084,N_15714);
nand U24068 (N_24068,N_18060,N_16922);
and U24069 (N_24069,N_15906,N_17945);
or U24070 (N_24070,N_18378,N_15565);
xnor U24071 (N_24071,N_19048,N_15640);
xnor U24072 (N_24072,N_19373,N_18749);
nor U24073 (N_24073,N_19270,N_19066);
and U24074 (N_24074,N_17004,N_15570);
nand U24075 (N_24075,N_17813,N_17560);
and U24076 (N_24076,N_17221,N_18009);
nor U24077 (N_24077,N_19615,N_16140);
or U24078 (N_24078,N_16437,N_17662);
or U24079 (N_24079,N_16120,N_17817);
and U24080 (N_24080,N_19806,N_15486);
nand U24081 (N_24081,N_19021,N_17721);
and U24082 (N_24082,N_17876,N_18502);
and U24083 (N_24083,N_18029,N_16460);
or U24084 (N_24084,N_15165,N_17928);
or U24085 (N_24085,N_16320,N_17197);
or U24086 (N_24086,N_18815,N_18784);
nor U24087 (N_24087,N_18370,N_17751);
or U24088 (N_24088,N_18184,N_15137);
or U24089 (N_24089,N_19332,N_15348);
or U24090 (N_24090,N_15610,N_19803);
nor U24091 (N_24091,N_19582,N_19179);
nor U24092 (N_24092,N_15540,N_19982);
or U24093 (N_24093,N_15097,N_17026);
and U24094 (N_24094,N_17302,N_15863);
xnor U24095 (N_24095,N_17236,N_18154);
nand U24096 (N_24096,N_18947,N_15049);
nor U24097 (N_24097,N_16352,N_18233);
nand U24098 (N_24098,N_17632,N_17965);
nor U24099 (N_24099,N_17975,N_18835);
nor U24100 (N_24100,N_16438,N_19087);
nor U24101 (N_24101,N_18644,N_15027);
or U24102 (N_24102,N_15950,N_18994);
nor U24103 (N_24103,N_18505,N_19965);
and U24104 (N_24104,N_19792,N_15059);
xor U24105 (N_24105,N_18184,N_19212);
or U24106 (N_24106,N_18035,N_19166);
or U24107 (N_24107,N_17671,N_16698);
nor U24108 (N_24108,N_18927,N_15276);
or U24109 (N_24109,N_18102,N_18479);
and U24110 (N_24110,N_17001,N_16722);
nand U24111 (N_24111,N_16539,N_15002);
xor U24112 (N_24112,N_18656,N_18366);
xor U24113 (N_24113,N_15558,N_17421);
or U24114 (N_24114,N_19568,N_15300);
nor U24115 (N_24115,N_19987,N_19030);
or U24116 (N_24116,N_16032,N_19559);
nor U24117 (N_24117,N_17197,N_17232);
nor U24118 (N_24118,N_16960,N_19580);
and U24119 (N_24119,N_17448,N_18407);
xor U24120 (N_24120,N_18321,N_16011);
xnor U24121 (N_24121,N_19956,N_19289);
xnor U24122 (N_24122,N_18453,N_17557);
nand U24123 (N_24123,N_15129,N_19143);
xor U24124 (N_24124,N_17505,N_16614);
nand U24125 (N_24125,N_17470,N_15496);
nor U24126 (N_24126,N_16699,N_18844);
or U24127 (N_24127,N_16741,N_19226);
nand U24128 (N_24128,N_18567,N_18699);
or U24129 (N_24129,N_18726,N_17145);
nor U24130 (N_24130,N_18509,N_17818);
nor U24131 (N_24131,N_17547,N_16138);
and U24132 (N_24132,N_18902,N_18705);
nand U24133 (N_24133,N_17819,N_15785);
or U24134 (N_24134,N_18817,N_16807);
nand U24135 (N_24135,N_15915,N_17535);
nand U24136 (N_24136,N_18938,N_17770);
nor U24137 (N_24137,N_15100,N_17389);
nor U24138 (N_24138,N_15210,N_17875);
or U24139 (N_24139,N_16672,N_16734);
or U24140 (N_24140,N_16707,N_17614);
or U24141 (N_24141,N_16176,N_15503);
nand U24142 (N_24142,N_15590,N_18589);
nand U24143 (N_24143,N_18166,N_19761);
nor U24144 (N_24144,N_16964,N_17982);
xnor U24145 (N_24145,N_19028,N_18466);
nor U24146 (N_24146,N_16019,N_19514);
xnor U24147 (N_24147,N_18867,N_19881);
and U24148 (N_24148,N_16412,N_15223);
nor U24149 (N_24149,N_15333,N_16548);
or U24150 (N_24150,N_16823,N_19796);
or U24151 (N_24151,N_16746,N_19260);
or U24152 (N_24152,N_17345,N_17254);
xor U24153 (N_24153,N_15130,N_15185);
nor U24154 (N_24154,N_18090,N_17996);
nand U24155 (N_24155,N_15865,N_17308);
xor U24156 (N_24156,N_19958,N_18339);
nor U24157 (N_24157,N_19940,N_19767);
or U24158 (N_24158,N_15393,N_17282);
nor U24159 (N_24159,N_18170,N_18750);
or U24160 (N_24160,N_19247,N_15369);
nand U24161 (N_24161,N_17508,N_19728);
and U24162 (N_24162,N_18432,N_16011);
or U24163 (N_24163,N_17619,N_17123);
or U24164 (N_24164,N_16609,N_17417);
or U24165 (N_24165,N_18819,N_16486);
xor U24166 (N_24166,N_15709,N_18671);
nand U24167 (N_24167,N_17506,N_15760);
and U24168 (N_24168,N_17888,N_18024);
and U24169 (N_24169,N_19257,N_18951);
and U24170 (N_24170,N_18016,N_15217);
and U24171 (N_24171,N_18435,N_18691);
and U24172 (N_24172,N_18986,N_15242);
nor U24173 (N_24173,N_19885,N_16626);
nor U24174 (N_24174,N_17215,N_18998);
or U24175 (N_24175,N_19906,N_16094);
and U24176 (N_24176,N_19506,N_16371);
nand U24177 (N_24177,N_19383,N_15280);
nand U24178 (N_24178,N_15565,N_17795);
xor U24179 (N_24179,N_18339,N_18932);
and U24180 (N_24180,N_17973,N_15590);
and U24181 (N_24181,N_15632,N_17718);
or U24182 (N_24182,N_19159,N_15167);
or U24183 (N_24183,N_15034,N_17842);
or U24184 (N_24184,N_16644,N_19257);
xnor U24185 (N_24185,N_19150,N_16144);
or U24186 (N_24186,N_17419,N_16171);
or U24187 (N_24187,N_18781,N_15679);
and U24188 (N_24188,N_16237,N_17938);
and U24189 (N_24189,N_17967,N_17287);
or U24190 (N_24190,N_15739,N_19065);
nor U24191 (N_24191,N_18215,N_17944);
or U24192 (N_24192,N_17282,N_19542);
nor U24193 (N_24193,N_17239,N_15929);
nor U24194 (N_24194,N_17143,N_19837);
or U24195 (N_24195,N_16086,N_19076);
or U24196 (N_24196,N_17655,N_18989);
nand U24197 (N_24197,N_19511,N_15486);
and U24198 (N_24198,N_15714,N_19970);
and U24199 (N_24199,N_16384,N_17086);
and U24200 (N_24200,N_19674,N_16918);
nand U24201 (N_24201,N_15917,N_16679);
nor U24202 (N_24202,N_17828,N_17304);
and U24203 (N_24203,N_17568,N_18686);
xor U24204 (N_24204,N_17437,N_19247);
nand U24205 (N_24205,N_15223,N_18734);
nor U24206 (N_24206,N_15443,N_19878);
nand U24207 (N_24207,N_18801,N_15720);
or U24208 (N_24208,N_16604,N_19532);
and U24209 (N_24209,N_16828,N_16567);
nand U24210 (N_24210,N_15993,N_17279);
or U24211 (N_24211,N_19417,N_18431);
nor U24212 (N_24212,N_16685,N_17927);
xnor U24213 (N_24213,N_19587,N_17570);
and U24214 (N_24214,N_16735,N_17649);
and U24215 (N_24215,N_15693,N_18592);
and U24216 (N_24216,N_16760,N_19946);
or U24217 (N_24217,N_16675,N_18472);
nor U24218 (N_24218,N_16984,N_17551);
nand U24219 (N_24219,N_18729,N_16149);
and U24220 (N_24220,N_15073,N_17034);
and U24221 (N_24221,N_18780,N_15003);
or U24222 (N_24222,N_17971,N_19256);
or U24223 (N_24223,N_17218,N_16772);
or U24224 (N_24224,N_18730,N_17587);
nor U24225 (N_24225,N_17609,N_18103);
nand U24226 (N_24226,N_16562,N_19793);
nand U24227 (N_24227,N_18368,N_19066);
nor U24228 (N_24228,N_16550,N_17124);
nor U24229 (N_24229,N_18722,N_17570);
nand U24230 (N_24230,N_18273,N_19972);
or U24231 (N_24231,N_17078,N_17645);
and U24232 (N_24232,N_16694,N_17326);
and U24233 (N_24233,N_19787,N_15815);
nor U24234 (N_24234,N_18943,N_18455);
nand U24235 (N_24235,N_17435,N_15053);
nor U24236 (N_24236,N_18686,N_19986);
and U24237 (N_24237,N_16505,N_15177);
nand U24238 (N_24238,N_16826,N_15738);
nand U24239 (N_24239,N_15141,N_18561);
nor U24240 (N_24240,N_15685,N_16946);
nand U24241 (N_24241,N_16499,N_19290);
or U24242 (N_24242,N_15852,N_15238);
and U24243 (N_24243,N_18992,N_16275);
nor U24244 (N_24244,N_17099,N_15563);
or U24245 (N_24245,N_18778,N_16816);
or U24246 (N_24246,N_17679,N_17139);
or U24247 (N_24247,N_17438,N_15204);
nand U24248 (N_24248,N_19436,N_18768);
xor U24249 (N_24249,N_15118,N_16079);
and U24250 (N_24250,N_17316,N_17267);
or U24251 (N_24251,N_16387,N_16902);
and U24252 (N_24252,N_16186,N_17049);
xor U24253 (N_24253,N_18946,N_16144);
or U24254 (N_24254,N_17794,N_19780);
or U24255 (N_24255,N_15172,N_15344);
and U24256 (N_24256,N_17739,N_16898);
nand U24257 (N_24257,N_19655,N_19408);
or U24258 (N_24258,N_17209,N_19219);
xor U24259 (N_24259,N_16060,N_17839);
or U24260 (N_24260,N_18670,N_16217);
xnor U24261 (N_24261,N_19183,N_16084);
nor U24262 (N_24262,N_19345,N_18751);
or U24263 (N_24263,N_16720,N_18533);
nor U24264 (N_24264,N_15953,N_16612);
nor U24265 (N_24265,N_17700,N_15744);
and U24266 (N_24266,N_15711,N_15888);
nand U24267 (N_24267,N_15724,N_16135);
and U24268 (N_24268,N_19505,N_19887);
and U24269 (N_24269,N_18750,N_18958);
nand U24270 (N_24270,N_16280,N_16477);
and U24271 (N_24271,N_17236,N_17439);
nand U24272 (N_24272,N_17187,N_16105);
nand U24273 (N_24273,N_18407,N_17324);
or U24274 (N_24274,N_18179,N_15764);
nand U24275 (N_24275,N_15918,N_16568);
or U24276 (N_24276,N_18719,N_15422);
and U24277 (N_24277,N_18759,N_18573);
and U24278 (N_24278,N_17946,N_19472);
nor U24279 (N_24279,N_17041,N_18519);
and U24280 (N_24280,N_18248,N_18040);
or U24281 (N_24281,N_18801,N_18162);
nand U24282 (N_24282,N_18663,N_16457);
nand U24283 (N_24283,N_16818,N_16986);
nor U24284 (N_24284,N_19748,N_18562);
nor U24285 (N_24285,N_17934,N_17799);
nor U24286 (N_24286,N_15690,N_17320);
or U24287 (N_24287,N_17573,N_16525);
or U24288 (N_24288,N_17977,N_18927);
and U24289 (N_24289,N_16278,N_19764);
xor U24290 (N_24290,N_19461,N_16588);
or U24291 (N_24291,N_18298,N_18287);
nor U24292 (N_24292,N_19321,N_17774);
nor U24293 (N_24293,N_16532,N_16665);
xnor U24294 (N_24294,N_18896,N_15700);
and U24295 (N_24295,N_15058,N_15563);
nand U24296 (N_24296,N_15884,N_15731);
nor U24297 (N_24297,N_15919,N_15102);
or U24298 (N_24298,N_15967,N_18137);
xor U24299 (N_24299,N_17681,N_19727);
or U24300 (N_24300,N_17504,N_17103);
or U24301 (N_24301,N_17404,N_15911);
nand U24302 (N_24302,N_15775,N_19904);
nor U24303 (N_24303,N_19482,N_18698);
nor U24304 (N_24304,N_17431,N_18768);
nor U24305 (N_24305,N_15009,N_16129);
and U24306 (N_24306,N_18444,N_19827);
xor U24307 (N_24307,N_15549,N_16433);
or U24308 (N_24308,N_18624,N_19265);
or U24309 (N_24309,N_15966,N_16995);
xor U24310 (N_24310,N_17698,N_17067);
xnor U24311 (N_24311,N_16557,N_17807);
nor U24312 (N_24312,N_15706,N_17736);
or U24313 (N_24313,N_16647,N_18921);
and U24314 (N_24314,N_19395,N_19474);
or U24315 (N_24315,N_18682,N_16466);
xor U24316 (N_24316,N_19301,N_15203);
and U24317 (N_24317,N_18356,N_18583);
nand U24318 (N_24318,N_18349,N_18154);
xor U24319 (N_24319,N_18801,N_17530);
nand U24320 (N_24320,N_18312,N_16576);
nor U24321 (N_24321,N_15520,N_15635);
or U24322 (N_24322,N_19194,N_19935);
or U24323 (N_24323,N_17529,N_15403);
or U24324 (N_24324,N_18418,N_16696);
nand U24325 (N_24325,N_16091,N_18737);
nor U24326 (N_24326,N_19111,N_17234);
nand U24327 (N_24327,N_15661,N_18013);
and U24328 (N_24328,N_15245,N_17117);
nand U24329 (N_24329,N_17043,N_16611);
nand U24330 (N_24330,N_15886,N_19089);
and U24331 (N_24331,N_16637,N_16804);
or U24332 (N_24332,N_15676,N_18753);
xor U24333 (N_24333,N_16733,N_15602);
nor U24334 (N_24334,N_16138,N_16974);
nor U24335 (N_24335,N_19501,N_18543);
or U24336 (N_24336,N_15268,N_17616);
nand U24337 (N_24337,N_19985,N_17086);
nor U24338 (N_24338,N_16866,N_17344);
and U24339 (N_24339,N_18770,N_19222);
nor U24340 (N_24340,N_15673,N_18547);
and U24341 (N_24341,N_15864,N_19389);
or U24342 (N_24342,N_17201,N_16943);
or U24343 (N_24343,N_18061,N_17217);
xor U24344 (N_24344,N_19976,N_18704);
xnor U24345 (N_24345,N_17439,N_15814);
and U24346 (N_24346,N_16158,N_18307);
nand U24347 (N_24347,N_17245,N_18209);
or U24348 (N_24348,N_19275,N_16789);
nand U24349 (N_24349,N_19229,N_16454);
or U24350 (N_24350,N_19019,N_15174);
and U24351 (N_24351,N_16379,N_16400);
nor U24352 (N_24352,N_18634,N_17311);
nor U24353 (N_24353,N_16438,N_19016);
nor U24354 (N_24354,N_15278,N_17267);
nor U24355 (N_24355,N_19797,N_15227);
and U24356 (N_24356,N_18126,N_16787);
and U24357 (N_24357,N_19640,N_16568);
nand U24358 (N_24358,N_18419,N_16283);
nor U24359 (N_24359,N_18716,N_18531);
nor U24360 (N_24360,N_18953,N_15190);
nand U24361 (N_24361,N_17885,N_16530);
and U24362 (N_24362,N_19863,N_15508);
or U24363 (N_24363,N_18342,N_18267);
xnor U24364 (N_24364,N_17416,N_17284);
nor U24365 (N_24365,N_19089,N_18997);
and U24366 (N_24366,N_17801,N_17897);
nor U24367 (N_24367,N_16454,N_19969);
nand U24368 (N_24368,N_16128,N_17865);
or U24369 (N_24369,N_18569,N_17360);
nand U24370 (N_24370,N_18293,N_18128);
or U24371 (N_24371,N_17305,N_16761);
or U24372 (N_24372,N_18568,N_17711);
or U24373 (N_24373,N_18503,N_19544);
and U24374 (N_24374,N_17716,N_17249);
or U24375 (N_24375,N_17989,N_16914);
nor U24376 (N_24376,N_18210,N_18709);
nor U24377 (N_24377,N_18188,N_15612);
and U24378 (N_24378,N_18251,N_16656);
or U24379 (N_24379,N_18573,N_17404);
nand U24380 (N_24380,N_17538,N_17610);
nand U24381 (N_24381,N_15111,N_15825);
nor U24382 (N_24382,N_16796,N_15585);
nand U24383 (N_24383,N_18236,N_17217);
nor U24384 (N_24384,N_16148,N_15372);
and U24385 (N_24385,N_16676,N_19576);
or U24386 (N_24386,N_16129,N_16747);
nor U24387 (N_24387,N_18189,N_19966);
nor U24388 (N_24388,N_18834,N_19676);
nand U24389 (N_24389,N_19261,N_15887);
nor U24390 (N_24390,N_18124,N_17229);
and U24391 (N_24391,N_15460,N_16126);
nor U24392 (N_24392,N_15133,N_17085);
and U24393 (N_24393,N_15765,N_16224);
nand U24394 (N_24394,N_15948,N_15090);
nand U24395 (N_24395,N_18970,N_17592);
or U24396 (N_24396,N_15252,N_15228);
or U24397 (N_24397,N_16781,N_17693);
nand U24398 (N_24398,N_17062,N_19827);
or U24399 (N_24399,N_15219,N_19464);
nand U24400 (N_24400,N_15466,N_17461);
or U24401 (N_24401,N_19681,N_17009);
or U24402 (N_24402,N_16442,N_17224);
nand U24403 (N_24403,N_18325,N_16780);
xor U24404 (N_24404,N_18840,N_17550);
xnor U24405 (N_24405,N_19495,N_15760);
nand U24406 (N_24406,N_18069,N_18481);
nand U24407 (N_24407,N_19456,N_15185);
and U24408 (N_24408,N_18064,N_19789);
nand U24409 (N_24409,N_19280,N_16059);
nand U24410 (N_24410,N_15634,N_16427);
or U24411 (N_24411,N_19862,N_16550);
xor U24412 (N_24412,N_18538,N_18100);
or U24413 (N_24413,N_16244,N_19624);
nand U24414 (N_24414,N_18938,N_16102);
and U24415 (N_24415,N_18290,N_15488);
or U24416 (N_24416,N_17692,N_18530);
nor U24417 (N_24417,N_16671,N_19536);
nand U24418 (N_24418,N_18256,N_19829);
or U24419 (N_24419,N_17879,N_15939);
nand U24420 (N_24420,N_19940,N_16632);
and U24421 (N_24421,N_18350,N_18621);
nor U24422 (N_24422,N_18529,N_18985);
nor U24423 (N_24423,N_18439,N_17990);
xnor U24424 (N_24424,N_15859,N_18052);
or U24425 (N_24425,N_17762,N_18683);
and U24426 (N_24426,N_18620,N_18696);
xnor U24427 (N_24427,N_16236,N_15534);
or U24428 (N_24428,N_18691,N_16157);
nand U24429 (N_24429,N_18932,N_18221);
and U24430 (N_24430,N_19107,N_17805);
or U24431 (N_24431,N_19961,N_18187);
nor U24432 (N_24432,N_16395,N_16315);
nor U24433 (N_24433,N_16877,N_16097);
and U24434 (N_24434,N_19630,N_17365);
or U24435 (N_24435,N_18545,N_17217);
nor U24436 (N_24436,N_19942,N_19844);
and U24437 (N_24437,N_18588,N_16875);
and U24438 (N_24438,N_19327,N_17461);
xor U24439 (N_24439,N_17417,N_17276);
xor U24440 (N_24440,N_17150,N_19731);
nor U24441 (N_24441,N_15876,N_18928);
or U24442 (N_24442,N_18669,N_18098);
nand U24443 (N_24443,N_19746,N_16317);
xnor U24444 (N_24444,N_17774,N_17204);
or U24445 (N_24445,N_15013,N_16605);
nand U24446 (N_24446,N_15681,N_18718);
or U24447 (N_24447,N_15828,N_19957);
xnor U24448 (N_24448,N_18643,N_19187);
nor U24449 (N_24449,N_19437,N_15309);
xnor U24450 (N_24450,N_16342,N_16768);
nor U24451 (N_24451,N_17449,N_15348);
nand U24452 (N_24452,N_16457,N_17700);
and U24453 (N_24453,N_18311,N_16198);
nor U24454 (N_24454,N_18331,N_18791);
nand U24455 (N_24455,N_19095,N_16336);
or U24456 (N_24456,N_18669,N_18310);
xnor U24457 (N_24457,N_16774,N_17967);
and U24458 (N_24458,N_15878,N_17937);
nor U24459 (N_24459,N_18768,N_16795);
nor U24460 (N_24460,N_15601,N_19348);
nor U24461 (N_24461,N_15054,N_16828);
or U24462 (N_24462,N_17481,N_16464);
or U24463 (N_24463,N_17493,N_16940);
nand U24464 (N_24464,N_17474,N_18676);
nand U24465 (N_24465,N_16031,N_19400);
nand U24466 (N_24466,N_16926,N_15450);
and U24467 (N_24467,N_19330,N_16521);
nor U24468 (N_24468,N_15917,N_17919);
and U24469 (N_24469,N_16784,N_16083);
nand U24470 (N_24470,N_19897,N_19755);
xnor U24471 (N_24471,N_17530,N_19053);
nor U24472 (N_24472,N_17987,N_18722);
nand U24473 (N_24473,N_16464,N_18619);
nor U24474 (N_24474,N_19306,N_15114);
and U24475 (N_24475,N_17123,N_16391);
nand U24476 (N_24476,N_15934,N_15276);
nand U24477 (N_24477,N_16178,N_18676);
nor U24478 (N_24478,N_18377,N_15216);
xnor U24479 (N_24479,N_18308,N_16630);
and U24480 (N_24480,N_15053,N_17115);
nor U24481 (N_24481,N_18955,N_16009);
and U24482 (N_24482,N_15121,N_18447);
nand U24483 (N_24483,N_15652,N_18049);
nand U24484 (N_24484,N_18214,N_17116);
or U24485 (N_24485,N_17022,N_19990);
and U24486 (N_24486,N_15586,N_18008);
nor U24487 (N_24487,N_19873,N_16097);
nand U24488 (N_24488,N_18791,N_16799);
xnor U24489 (N_24489,N_19591,N_16321);
nand U24490 (N_24490,N_17787,N_18802);
or U24491 (N_24491,N_19718,N_19716);
xnor U24492 (N_24492,N_19674,N_19580);
nand U24493 (N_24493,N_19962,N_15805);
nor U24494 (N_24494,N_19549,N_16579);
or U24495 (N_24495,N_15360,N_17486);
and U24496 (N_24496,N_16314,N_16918);
nor U24497 (N_24497,N_18210,N_18054);
or U24498 (N_24498,N_16198,N_19096);
nor U24499 (N_24499,N_15359,N_15746);
nand U24500 (N_24500,N_16166,N_19556);
nor U24501 (N_24501,N_15364,N_18753);
nand U24502 (N_24502,N_15568,N_19045);
nand U24503 (N_24503,N_19238,N_15779);
xnor U24504 (N_24504,N_15270,N_18006);
nor U24505 (N_24505,N_16728,N_19731);
and U24506 (N_24506,N_19843,N_18090);
and U24507 (N_24507,N_15614,N_16245);
xor U24508 (N_24508,N_15182,N_19538);
nand U24509 (N_24509,N_17952,N_15172);
or U24510 (N_24510,N_15345,N_19954);
nor U24511 (N_24511,N_19235,N_18217);
or U24512 (N_24512,N_15797,N_15537);
nand U24513 (N_24513,N_15554,N_15264);
or U24514 (N_24514,N_19741,N_17236);
and U24515 (N_24515,N_15202,N_15620);
nand U24516 (N_24516,N_19051,N_19111);
or U24517 (N_24517,N_19739,N_16186);
nand U24518 (N_24518,N_18122,N_18203);
nor U24519 (N_24519,N_18119,N_17873);
or U24520 (N_24520,N_15155,N_15914);
nor U24521 (N_24521,N_15950,N_15917);
nor U24522 (N_24522,N_15029,N_17166);
nand U24523 (N_24523,N_15273,N_16016);
or U24524 (N_24524,N_17748,N_15403);
or U24525 (N_24525,N_19816,N_16700);
nand U24526 (N_24526,N_16925,N_16897);
nand U24527 (N_24527,N_17542,N_19081);
or U24528 (N_24528,N_15821,N_18619);
nand U24529 (N_24529,N_19379,N_15638);
nor U24530 (N_24530,N_15994,N_19912);
nand U24531 (N_24531,N_17721,N_16107);
nor U24532 (N_24532,N_18602,N_16874);
nor U24533 (N_24533,N_16860,N_19871);
nor U24534 (N_24534,N_18767,N_19850);
and U24535 (N_24535,N_19515,N_18373);
nand U24536 (N_24536,N_17534,N_18841);
or U24537 (N_24537,N_19373,N_19857);
nor U24538 (N_24538,N_18495,N_15876);
or U24539 (N_24539,N_16555,N_16842);
and U24540 (N_24540,N_16307,N_17954);
and U24541 (N_24541,N_15741,N_18722);
or U24542 (N_24542,N_16504,N_17733);
or U24543 (N_24543,N_18901,N_18913);
or U24544 (N_24544,N_17029,N_16620);
xnor U24545 (N_24545,N_15827,N_19884);
or U24546 (N_24546,N_15456,N_17246);
or U24547 (N_24547,N_19915,N_18680);
nor U24548 (N_24548,N_18261,N_18757);
or U24549 (N_24549,N_16766,N_16599);
or U24550 (N_24550,N_15640,N_17618);
or U24551 (N_24551,N_18814,N_19795);
nand U24552 (N_24552,N_17030,N_17236);
and U24553 (N_24553,N_18257,N_15621);
nand U24554 (N_24554,N_19418,N_18176);
and U24555 (N_24555,N_16627,N_18376);
nand U24556 (N_24556,N_17419,N_18473);
or U24557 (N_24557,N_19569,N_17653);
and U24558 (N_24558,N_16059,N_19101);
or U24559 (N_24559,N_16868,N_15068);
nor U24560 (N_24560,N_19831,N_18123);
or U24561 (N_24561,N_15410,N_17757);
nand U24562 (N_24562,N_18141,N_16052);
and U24563 (N_24563,N_19617,N_16283);
and U24564 (N_24564,N_16100,N_15750);
nor U24565 (N_24565,N_19572,N_15490);
xnor U24566 (N_24566,N_15400,N_18446);
xnor U24567 (N_24567,N_19728,N_17991);
nand U24568 (N_24568,N_17041,N_18592);
nand U24569 (N_24569,N_15564,N_19042);
and U24570 (N_24570,N_17305,N_18340);
nor U24571 (N_24571,N_17844,N_19778);
nand U24572 (N_24572,N_15539,N_18361);
nand U24573 (N_24573,N_18209,N_19862);
nor U24574 (N_24574,N_17475,N_19435);
nor U24575 (N_24575,N_17867,N_18457);
xnor U24576 (N_24576,N_17151,N_19451);
or U24577 (N_24577,N_16858,N_17901);
and U24578 (N_24578,N_16364,N_19119);
xor U24579 (N_24579,N_15225,N_16102);
nand U24580 (N_24580,N_15685,N_16317);
nand U24581 (N_24581,N_16952,N_18374);
nand U24582 (N_24582,N_18050,N_18821);
and U24583 (N_24583,N_16239,N_16199);
nand U24584 (N_24584,N_19786,N_18220);
xor U24585 (N_24585,N_18958,N_18631);
nor U24586 (N_24586,N_19867,N_18773);
nand U24587 (N_24587,N_15730,N_17484);
or U24588 (N_24588,N_18295,N_19977);
nand U24589 (N_24589,N_17691,N_18756);
nor U24590 (N_24590,N_18535,N_17953);
or U24591 (N_24591,N_19138,N_18440);
or U24592 (N_24592,N_16746,N_15356);
xnor U24593 (N_24593,N_18704,N_16262);
or U24594 (N_24594,N_16532,N_19133);
and U24595 (N_24595,N_19492,N_16790);
or U24596 (N_24596,N_16106,N_19069);
or U24597 (N_24597,N_17563,N_17676);
nor U24598 (N_24598,N_18765,N_15461);
or U24599 (N_24599,N_18086,N_15431);
and U24600 (N_24600,N_19468,N_16147);
and U24601 (N_24601,N_15140,N_19828);
nor U24602 (N_24602,N_15940,N_16738);
nor U24603 (N_24603,N_16129,N_17157);
nand U24604 (N_24604,N_16083,N_18220);
and U24605 (N_24605,N_15523,N_17295);
xor U24606 (N_24606,N_17379,N_15296);
and U24607 (N_24607,N_19980,N_17757);
nor U24608 (N_24608,N_17980,N_16174);
or U24609 (N_24609,N_18267,N_15566);
nor U24610 (N_24610,N_17680,N_15370);
and U24611 (N_24611,N_16539,N_16589);
nor U24612 (N_24612,N_19114,N_16982);
nor U24613 (N_24613,N_19382,N_16075);
nor U24614 (N_24614,N_15523,N_17139);
and U24615 (N_24615,N_18056,N_17009);
nand U24616 (N_24616,N_19648,N_17743);
nor U24617 (N_24617,N_15465,N_18908);
or U24618 (N_24618,N_19926,N_18748);
or U24619 (N_24619,N_15452,N_19303);
and U24620 (N_24620,N_17293,N_18764);
nor U24621 (N_24621,N_18218,N_19390);
nand U24622 (N_24622,N_16083,N_18330);
nand U24623 (N_24623,N_15035,N_15025);
or U24624 (N_24624,N_19897,N_18337);
nand U24625 (N_24625,N_19637,N_16070);
nor U24626 (N_24626,N_17862,N_17934);
or U24627 (N_24627,N_15017,N_19801);
nand U24628 (N_24628,N_17158,N_19081);
and U24629 (N_24629,N_17230,N_16064);
or U24630 (N_24630,N_19145,N_16743);
xnor U24631 (N_24631,N_19895,N_15180);
nand U24632 (N_24632,N_15916,N_17980);
and U24633 (N_24633,N_18349,N_18943);
and U24634 (N_24634,N_19622,N_18999);
or U24635 (N_24635,N_17360,N_15264);
and U24636 (N_24636,N_15102,N_16274);
or U24637 (N_24637,N_16472,N_16663);
or U24638 (N_24638,N_19077,N_18217);
nand U24639 (N_24639,N_18654,N_18845);
or U24640 (N_24640,N_18964,N_17727);
and U24641 (N_24641,N_19240,N_19238);
or U24642 (N_24642,N_15736,N_18934);
or U24643 (N_24643,N_17991,N_17679);
nand U24644 (N_24644,N_18198,N_15365);
or U24645 (N_24645,N_19874,N_15071);
and U24646 (N_24646,N_17550,N_19560);
and U24647 (N_24647,N_15097,N_19485);
or U24648 (N_24648,N_18473,N_18038);
and U24649 (N_24649,N_18146,N_15304);
xnor U24650 (N_24650,N_18753,N_16997);
nor U24651 (N_24651,N_15448,N_17084);
or U24652 (N_24652,N_15281,N_15966);
nor U24653 (N_24653,N_18834,N_18873);
and U24654 (N_24654,N_17566,N_15602);
nand U24655 (N_24655,N_18197,N_17040);
and U24656 (N_24656,N_19934,N_18792);
nor U24657 (N_24657,N_18750,N_15284);
nand U24658 (N_24658,N_15047,N_19187);
nand U24659 (N_24659,N_15250,N_16118);
nand U24660 (N_24660,N_18368,N_16594);
nand U24661 (N_24661,N_19153,N_17590);
nand U24662 (N_24662,N_16990,N_16369);
or U24663 (N_24663,N_18339,N_17043);
nor U24664 (N_24664,N_19697,N_15375);
or U24665 (N_24665,N_18313,N_18194);
nand U24666 (N_24666,N_19705,N_18421);
or U24667 (N_24667,N_18632,N_17451);
and U24668 (N_24668,N_15528,N_18271);
nor U24669 (N_24669,N_16241,N_16663);
or U24670 (N_24670,N_17454,N_18734);
nor U24671 (N_24671,N_16456,N_17451);
nor U24672 (N_24672,N_18608,N_15570);
nand U24673 (N_24673,N_18179,N_15609);
and U24674 (N_24674,N_18158,N_15915);
nand U24675 (N_24675,N_17919,N_17664);
and U24676 (N_24676,N_19660,N_19046);
nand U24677 (N_24677,N_16957,N_19477);
or U24678 (N_24678,N_17239,N_18847);
nand U24679 (N_24679,N_15631,N_18932);
and U24680 (N_24680,N_18983,N_17003);
xor U24681 (N_24681,N_16828,N_17108);
nor U24682 (N_24682,N_16250,N_16493);
nand U24683 (N_24683,N_19092,N_19088);
or U24684 (N_24684,N_18032,N_19424);
and U24685 (N_24685,N_18241,N_17921);
or U24686 (N_24686,N_17446,N_15088);
or U24687 (N_24687,N_17966,N_17894);
and U24688 (N_24688,N_17453,N_18314);
or U24689 (N_24689,N_18029,N_17556);
or U24690 (N_24690,N_17376,N_18476);
or U24691 (N_24691,N_19440,N_15586);
nand U24692 (N_24692,N_16526,N_16093);
and U24693 (N_24693,N_17622,N_15982);
nor U24694 (N_24694,N_16794,N_17445);
and U24695 (N_24695,N_19411,N_16148);
and U24696 (N_24696,N_19255,N_17856);
nand U24697 (N_24697,N_15070,N_17923);
or U24698 (N_24698,N_16908,N_16113);
and U24699 (N_24699,N_19644,N_19281);
xnor U24700 (N_24700,N_18427,N_17285);
and U24701 (N_24701,N_16724,N_15696);
nand U24702 (N_24702,N_17766,N_18895);
and U24703 (N_24703,N_16072,N_16326);
nand U24704 (N_24704,N_18679,N_16207);
and U24705 (N_24705,N_17981,N_19997);
and U24706 (N_24706,N_17086,N_15085);
nor U24707 (N_24707,N_17015,N_18196);
nor U24708 (N_24708,N_19016,N_18191);
and U24709 (N_24709,N_16480,N_15903);
xor U24710 (N_24710,N_15294,N_15846);
nand U24711 (N_24711,N_17527,N_15921);
nand U24712 (N_24712,N_16199,N_17571);
nand U24713 (N_24713,N_17985,N_16038);
nor U24714 (N_24714,N_18344,N_17731);
nand U24715 (N_24715,N_17056,N_16601);
or U24716 (N_24716,N_16993,N_19127);
nor U24717 (N_24717,N_18735,N_16339);
and U24718 (N_24718,N_19714,N_18142);
nand U24719 (N_24719,N_17864,N_15439);
nor U24720 (N_24720,N_17423,N_15000);
nand U24721 (N_24721,N_18522,N_19934);
nand U24722 (N_24722,N_16462,N_15586);
and U24723 (N_24723,N_17310,N_15254);
or U24724 (N_24724,N_18197,N_16158);
xor U24725 (N_24725,N_15504,N_17529);
nor U24726 (N_24726,N_18501,N_15460);
and U24727 (N_24727,N_17735,N_16897);
or U24728 (N_24728,N_18969,N_17549);
or U24729 (N_24729,N_18335,N_16816);
or U24730 (N_24730,N_17926,N_19636);
or U24731 (N_24731,N_18866,N_19661);
and U24732 (N_24732,N_17425,N_16295);
and U24733 (N_24733,N_17749,N_19942);
and U24734 (N_24734,N_17093,N_15296);
nor U24735 (N_24735,N_17305,N_17408);
xor U24736 (N_24736,N_16858,N_19519);
or U24737 (N_24737,N_19088,N_18637);
nand U24738 (N_24738,N_16226,N_16635);
or U24739 (N_24739,N_16588,N_19791);
nand U24740 (N_24740,N_17654,N_15199);
nor U24741 (N_24741,N_19225,N_15491);
xor U24742 (N_24742,N_17907,N_18875);
or U24743 (N_24743,N_17254,N_18683);
and U24744 (N_24744,N_19255,N_15080);
and U24745 (N_24745,N_16894,N_15682);
and U24746 (N_24746,N_17343,N_18802);
nor U24747 (N_24747,N_19790,N_18570);
nand U24748 (N_24748,N_19650,N_19245);
and U24749 (N_24749,N_16215,N_19858);
nor U24750 (N_24750,N_16238,N_18627);
nand U24751 (N_24751,N_19062,N_17740);
xnor U24752 (N_24752,N_17728,N_15274);
or U24753 (N_24753,N_17891,N_17085);
and U24754 (N_24754,N_19634,N_17243);
or U24755 (N_24755,N_19290,N_15208);
and U24756 (N_24756,N_18962,N_16396);
nor U24757 (N_24757,N_18241,N_19817);
and U24758 (N_24758,N_18137,N_18243);
xor U24759 (N_24759,N_16315,N_19962);
nand U24760 (N_24760,N_19014,N_15044);
or U24761 (N_24761,N_18348,N_16145);
or U24762 (N_24762,N_19253,N_15507);
and U24763 (N_24763,N_15614,N_18992);
or U24764 (N_24764,N_15588,N_17431);
nor U24765 (N_24765,N_17216,N_18363);
nand U24766 (N_24766,N_18792,N_17468);
nand U24767 (N_24767,N_18625,N_18306);
nor U24768 (N_24768,N_16070,N_17250);
or U24769 (N_24769,N_16424,N_17329);
nand U24770 (N_24770,N_16487,N_18314);
or U24771 (N_24771,N_18406,N_17256);
nand U24772 (N_24772,N_15604,N_18114);
xor U24773 (N_24773,N_19132,N_15207);
and U24774 (N_24774,N_15083,N_16898);
nand U24775 (N_24775,N_18292,N_18284);
or U24776 (N_24776,N_15453,N_17630);
nand U24777 (N_24777,N_16450,N_15203);
nor U24778 (N_24778,N_15687,N_19998);
and U24779 (N_24779,N_19986,N_18275);
nor U24780 (N_24780,N_16701,N_15076);
or U24781 (N_24781,N_16634,N_17960);
or U24782 (N_24782,N_18561,N_19078);
or U24783 (N_24783,N_16299,N_19964);
or U24784 (N_24784,N_17191,N_19174);
nand U24785 (N_24785,N_15996,N_16789);
and U24786 (N_24786,N_16242,N_18763);
nor U24787 (N_24787,N_17012,N_16173);
or U24788 (N_24788,N_16254,N_19374);
or U24789 (N_24789,N_18028,N_19251);
or U24790 (N_24790,N_19699,N_16608);
nor U24791 (N_24791,N_15962,N_19276);
nand U24792 (N_24792,N_19667,N_18585);
nand U24793 (N_24793,N_18042,N_18125);
or U24794 (N_24794,N_15581,N_19450);
nand U24795 (N_24795,N_17162,N_17521);
nand U24796 (N_24796,N_15788,N_18406);
or U24797 (N_24797,N_19019,N_18435);
and U24798 (N_24798,N_17181,N_16641);
xnor U24799 (N_24799,N_18806,N_19685);
nor U24800 (N_24800,N_15959,N_16477);
nand U24801 (N_24801,N_15262,N_16099);
and U24802 (N_24802,N_17079,N_19396);
and U24803 (N_24803,N_17936,N_19247);
or U24804 (N_24804,N_17813,N_16061);
nor U24805 (N_24805,N_18016,N_19598);
and U24806 (N_24806,N_16613,N_19453);
nand U24807 (N_24807,N_17749,N_18530);
nand U24808 (N_24808,N_17201,N_17491);
or U24809 (N_24809,N_17985,N_17802);
nand U24810 (N_24810,N_15820,N_17117);
nor U24811 (N_24811,N_16023,N_19478);
or U24812 (N_24812,N_18832,N_15432);
xor U24813 (N_24813,N_17588,N_19621);
or U24814 (N_24814,N_18312,N_19707);
nor U24815 (N_24815,N_19025,N_19907);
or U24816 (N_24816,N_19012,N_17995);
nand U24817 (N_24817,N_15599,N_16791);
nor U24818 (N_24818,N_17008,N_17196);
and U24819 (N_24819,N_19425,N_19086);
or U24820 (N_24820,N_16583,N_19977);
nor U24821 (N_24821,N_15912,N_17667);
or U24822 (N_24822,N_18225,N_16308);
and U24823 (N_24823,N_19295,N_18918);
or U24824 (N_24824,N_19334,N_19272);
xor U24825 (N_24825,N_15231,N_19477);
nor U24826 (N_24826,N_18853,N_15241);
nor U24827 (N_24827,N_17903,N_17408);
or U24828 (N_24828,N_19820,N_19463);
and U24829 (N_24829,N_17124,N_19179);
nor U24830 (N_24830,N_17295,N_16184);
and U24831 (N_24831,N_17426,N_19082);
and U24832 (N_24832,N_19432,N_16721);
and U24833 (N_24833,N_16510,N_15621);
nor U24834 (N_24834,N_19284,N_15417);
or U24835 (N_24835,N_19390,N_19912);
nand U24836 (N_24836,N_17887,N_19581);
nor U24837 (N_24837,N_16047,N_19989);
nand U24838 (N_24838,N_16594,N_19037);
nand U24839 (N_24839,N_15122,N_19912);
nand U24840 (N_24840,N_16745,N_18494);
nand U24841 (N_24841,N_16054,N_16884);
nor U24842 (N_24842,N_16615,N_16236);
and U24843 (N_24843,N_18986,N_16910);
and U24844 (N_24844,N_19631,N_18702);
nand U24845 (N_24845,N_16668,N_17292);
or U24846 (N_24846,N_19838,N_16554);
nor U24847 (N_24847,N_16491,N_19916);
nor U24848 (N_24848,N_16538,N_17212);
nand U24849 (N_24849,N_16548,N_18627);
nor U24850 (N_24850,N_18069,N_17707);
or U24851 (N_24851,N_17852,N_16389);
xnor U24852 (N_24852,N_19358,N_17506);
nand U24853 (N_24853,N_19843,N_15604);
nor U24854 (N_24854,N_18988,N_18387);
or U24855 (N_24855,N_15251,N_18964);
and U24856 (N_24856,N_17219,N_19120);
and U24857 (N_24857,N_16812,N_17941);
or U24858 (N_24858,N_16293,N_19670);
and U24859 (N_24859,N_17019,N_19519);
nor U24860 (N_24860,N_19083,N_17263);
or U24861 (N_24861,N_18787,N_17604);
nor U24862 (N_24862,N_18362,N_18577);
nand U24863 (N_24863,N_15261,N_19436);
and U24864 (N_24864,N_17258,N_19139);
nand U24865 (N_24865,N_19362,N_18729);
or U24866 (N_24866,N_18491,N_15439);
or U24867 (N_24867,N_16030,N_18004);
and U24868 (N_24868,N_18788,N_17794);
or U24869 (N_24869,N_19069,N_15996);
nor U24870 (N_24870,N_18546,N_15227);
and U24871 (N_24871,N_18828,N_18001);
nor U24872 (N_24872,N_15996,N_15560);
and U24873 (N_24873,N_15732,N_15666);
xor U24874 (N_24874,N_16373,N_15421);
and U24875 (N_24875,N_16501,N_18343);
and U24876 (N_24876,N_17158,N_19314);
and U24877 (N_24877,N_18798,N_18685);
nand U24878 (N_24878,N_18391,N_17431);
and U24879 (N_24879,N_17167,N_17857);
and U24880 (N_24880,N_16166,N_15026);
nor U24881 (N_24881,N_19329,N_19748);
and U24882 (N_24882,N_18777,N_19959);
nor U24883 (N_24883,N_19673,N_18724);
nor U24884 (N_24884,N_15394,N_17263);
nand U24885 (N_24885,N_17831,N_15009);
and U24886 (N_24886,N_18180,N_17509);
and U24887 (N_24887,N_16379,N_15520);
nor U24888 (N_24888,N_19996,N_15947);
nand U24889 (N_24889,N_15035,N_16140);
nor U24890 (N_24890,N_15119,N_17751);
and U24891 (N_24891,N_18627,N_19547);
nand U24892 (N_24892,N_18614,N_17530);
nor U24893 (N_24893,N_18252,N_15909);
or U24894 (N_24894,N_15979,N_15400);
or U24895 (N_24895,N_16732,N_18744);
or U24896 (N_24896,N_17442,N_17303);
nor U24897 (N_24897,N_18677,N_15679);
and U24898 (N_24898,N_16298,N_18972);
nand U24899 (N_24899,N_16436,N_19663);
and U24900 (N_24900,N_15241,N_19387);
or U24901 (N_24901,N_17329,N_15647);
nand U24902 (N_24902,N_19298,N_15139);
and U24903 (N_24903,N_16176,N_15675);
nand U24904 (N_24904,N_17752,N_16750);
and U24905 (N_24905,N_15219,N_18794);
nor U24906 (N_24906,N_16152,N_19771);
or U24907 (N_24907,N_19916,N_17568);
or U24908 (N_24908,N_18960,N_17881);
nor U24909 (N_24909,N_17344,N_18420);
or U24910 (N_24910,N_19123,N_18105);
nand U24911 (N_24911,N_17099,N_16482);
nand U24912 (N_24912,N_19730,N_15893);
or U24913 (N_24913,N_18647,N_17206);
nand U24914 (N_24914,N_18681,N_15306);
nor U24915 (N_24915,N_15325,N_17282);
nand U24916 (N_24916,N_17923,N_15542);
and U24917 (N_24917,N_15018,N_15370);
nor U24918 (N_24918,N_16211,N_19704);
nand U24919 (N_24919,N_16205,N_16661);
nand U24920 (N_24920,N_16123,N_16553);
and U24921 (N_24921,N_19836,N_15324);
and U24922 (N_24922,N_18366,N_15275);
and U24923 (N_24923,N_17507,N_19041);
xor U24924 (N_24924,N_17384,N_18926);
nand U24925 (N_24925,N_15778,N_19980);
or U24926 (N_24926,N_17826,N_15826);
nand U24927 (N_24927,N_16856,N_17911);
and U24928 (N_24928,N_16712,N_17358);
nor U24929 (N_24929,N_17414,N_18549);
and U24930 (N_24930,N_15908,N_18106);
nand U24931 (N_24931,N_15076,N_19138);
and U24932 (N_24932,N_15198,N_18757);
nand U24933 (N_24933,N_15939,N_19690);
nand U24934 (N_24934,N_15467,N_15105);
nand U24935 (N_24935,N_18089,N_15563);
nor U24936 (N_24936,N_15967,N_18698);
or U24937 (N_24937,N_16842,N_17079);
nand U24938 (N_24938,N_19374,N_18024);
nor U24939 (N_24939,N_19255,N_17205);
and U24940 (N_24940,N_17677,N_19769);
nand U24941 (N_24941,N_19973,N_15475);
nand U24942 (N_24942,N_17271,N_17406);
xnor U24943 (N_24943,N_19022,N_19268);
nand U24944 (N_24944,N_16690,N_19752);
or U24945 (N_24945,N_16379,N_16142);
or U24946 (N_24946,N_19091,N_17410);
and U24947 (N_24947,N_18481,N_19885);
nor U24948 (N_24948,N_17604,N_17588);
or U24949 (N_24949,N_19420,N_15035);
or U24950 (N_24950,N_18733,N_19407);
nand U24951 (N_24951,N_18334,N_16801);
xor U24952 (N_24952,N_17349,N_19548);
or U24953 (N_24953,N_17279,N_17929);
and U24954 (N_24954,N_15635,N_18403);
and U24955 (N_24955,N_17642,N_16766);
and U24956 (N_24956,N_18243,N_15869);
or U24957 (N_24957,N_15477,N_16346);
and U24958 (N_24958,N_19969,N_19836);
nor U24959 (N_24959,N_19572,N_19203);
or U24960 (N_24960,N_17997,N_15532);
nor U24961 (N_24961,N_15536,N_16091);
nor U24962 (N_24962,N_15496,N_17202);
or U24963 (N_24963,N_19343,N_18337);
and U24964 (N_24964,N_15726,N_15420);
nand U24965 (N_24965,N_15403,N_19210);
and U24966 (N_24966,N_16270,N_16242);
and U24967 (N_24967,N_18901,N_15889);
or U24968 (N_24968,N_15256,N_18418);
or U24969 (N_24969,N_17209,N_16950);
nor U24970 (N_24970,N_15550,N_16078);
nand U24971 (N_24971,N_18875,N_16983);
nor U24972 (N_24972,N_18801,N_16976);
xor U24973 (N_24973,N_16537,N_19126);
or U24974 (N_24974,N_16900,N_19706);
nand U24975 (N_24975,N_16292,N_18171);
nor U24976 (N_24976,N_17937,N_16534);
or U24977 (N_24977,N_15293,N_16075);
xnor U24978 (N_24978,N_15120,N_19845);
nor U24979 (N_24979,N_18582,N_16992);
nand U24980 (N_24980,N_19509,N_17650);
and U24981 (N_24981,N_17369,N_19787);
xor U24982 (N_24982,N_18638,N_19470);
nand U24983 (N_24983,N_18699,N_17697);
and U24984 (N_24984,N_15303,N_19789);
nor U24985 (N_24985,N_17488,N_17717);
nand U24986 (N_24986,N_17920,N_16183);
xor U24987 (N_24987,N_17458,N_15332);
nand U24988 (N_24988,N_19346,N_16929);
nand U24989 (N_24989,N_15453,N_19643);
nand U24990 (N_24990,N_15596,N_15506);
and U24991 (N_24991,N_19232,N_15476);
nand U24992 (N_24992,N_19931,N_17896);
or U24993 (N_24993,N_18455,N_15681);
nand U24994 (N_24994,N_19028,N_18207);
nand U24995 (N_24995,N_18862,N_16131);
nor U24996 (N_24996,N_15992,N_19748);
nand U24997 (N_24997,N_18820,N_18597);
nand U24998 (N_24998,N_19902,N_16612);
xnor U24999 (N_24999,N_18504,N_17273);
nor U25000 (N_25000,N_22833,N_23124);
nor U25001 (N_25001,N_23614,N_20605);
and U25002 (N_25002,N_21495,N_22211);
or U25003 (N_25003,N_20918,N_23023);
and U25004 (N_25004,N_23956,N_24641);
nand U25005 (N_25005,N_20854,N_24594);
nor U25006 (N_25006,N_20792,N_23423);
nand U25007 (N_25007,N_23960,N_21879);
and U25008 (N_25008,N_22981,N_20823);
nor U25009 (N_25009,N_24194,N_23586);
or U25010 (N_25010,N_24884,N_23888);
or U25011 (N_25011,N_24976,N_21679);
and U25012 (N_25012,N_23912,N_24896);
and U25013 (N_25013,N_21740,N_20153);
and U25014 (N_25014,N_20195,N_22939);
xnor U25015 (N_25015,N_24313,N_20194);
or U25016 (N_25016,N_20016,N_24882);
nor U25017 (N_25017,N_21512,N_22373);
nand U25018 (N_25018,N_21791,N_21023);
or U25019 (N_25019,N_21712,N_23833);
xor U25020 (N_25020,N_24687,N_23549);
xnor U25021 (N_25021,N_23851,N_21442);
nand U25022 (N_25022,N_23872,N_22481);
and U25023 (N_25023,N_24578,N_21190);
or U25024 (N_25024,N_22327,N_21052);
nor U25025 (N_25025,N_24166,N_23232);
nor U25026 (N_25026,N_21282,N_22271);
or U25027 (N_25027,N_21876,N_24052);
xnor U25028 (N_25028,N_22583,N_22463);
or U25029 (N_25029,N_23498,N_21539);
and U25030 (N_25030,N_22112,N_21426);
nor U25031 (N_25031,N_21746,N_23506);
nor U25032 (N_25032,N_23137,N_23234);
and U25033 (N_25033,N_23043,N_23926);
nand U25034 (N_25034,N_22850,N_22267);
nor U25035 (N_25035,N_23184,N_21720);
or U25036 (N_25036,N_21467,N_22356);
nor U25037 (N_25037,N_23138,N_22558);
nand U25038 (N_25038,N_22176,N_20866);
nor U25039 (N_25039,N_21962,N_21762);
xor U25040 (N_25040,N_24139,N_21311);
nor U25041 (N_25041,N_24541,N_22174);
nand U25042 (N_25042,N_23490,N_22553);
and U25043 (N_25043,N_23028,N_23091);
xnor U25044 (N_25044,N_20317,N_21880);
nand U25045 (N_25045,N_22477,N_20112);
nor U25046 (N_25046,N_21155,N_23323);
or U25047 (N_25047,N_23180,N_24036);
or U25048 (N_25048,N_21298,N_23420);
xor U25049 (N_25049,N_24010,N_22923);
xnor U25050 (N_25050,N_22437,N_20452);
or U25051 (N_25051,N_20429,N_23869);
or U25052 (N_25052,N_20995,N_21258);
and U25053 (N_25053,N_23082,N_24106);
or U25054 (N_25054,N_24350,N_24653);
or U25055 (N_25055,N_24928,N_23394);
or U25056 (N_25056,N_24588,N_23487);
nand U25057 (N_25057,N_20865,N_21218);
or U25058 (N_25058,N_20569,N_20223);
and U25059 (N_25059,N_24963,N_22368);
and U25060 (N_25060,N_23532,N_20040);
xnor U25061 (N_25061,N_23416,N_24191);
and U25062 (N_25062,N_21915,N_21095);
or U25063 (N_25063,N_21947,N_21663);
and U25064 (N_25064,N_21186,N_21891);
and U25065 (N_25065,N_24116,N_23330);
and U25066 (N_25066,N_20680,N_21295);
and U25067 (N_25067,N_20484,N_20954);
or U25068 (N_25068,N_22246,N_21728);
nand U25069 (N_25069,N_20777,N_20697);
nor U25070 (N_25070,N_20896,N_24266);
and U25071 (N_25071,N_23999,N_20034);
nand U25072 (N_25072,N_22045,N_24247);
and U25073 (N_25073,N_21597,N_22650);
xor U25074 (N_25074,N_20568,N_22040);
nand U25075 (N_25075,N_22216,N_21751);
nor U25076 (N_25076,N_22126,N_23930);
nand U25077 (N_25077,N_21197,N_22053);
nand U25078 (N_25078,N_23117,N_22351);
nand U25079 (N_25079,N_22046,N_24576);
nand U25080 (N_25080,N_23353,N_24842);
nor U25081 (N_25081,N_24899,N_24377);
or U25082 (N_25082,N_21261,N_24316);
or U25083 (N_25083,N_22128,N_23040);
nand U25084 (N_25084,N_22704,N_24544);
and U25085 (N_25085,N_20883,N_24535);
and U25086 (N_25086,N_22210,N_23044);
or U25087 (N_25087,N_20873,N_21669);
nand U25088 (N_25088,N_23431,N_22465);
or U25089 (N_25089,N_20991,N_23795);
nor U25090 (N_25090,N_20276,N_20330);
nand U25091 (N_25091,N_22906,N_22123);
xor U25092 (N_25092,N_23349,N_22333);
nor U25093 (N_25093,N_24584,N_23895);
or U25094 (N_25094,N_21318,N_20156);
or U25095 (N_25095,N_24823,N_20100);
xor U25096 (N_25096,N_21673,N_24930);
or U25097 (N_25097,N_23565,N_20011);
xor U25098 (N_25098,N_22688,N_22849);
or U25099 (N_25099,N_20344,N_21797);
nand U25100 (N_25100,N_21622,N_20655);
or U25101 (N_25101,N_21476,N_20685);
xor U25102 (N_25102,N_24102,N_21341);
and U25103 (N_25103,N_22291,N_24378);
or U25104 (N_25104,N_22404,N_22431);
and U25105 (N_25105,N_23003,N_24000);
nand U25106 (N_25106,N_23271,N_23205);
xnor U25107 (N_25107,N_21711,N_23317);
nor U25108 (N_25108,N_23211,N_24722);
and U25109 (N_25109,N_22446,N_21838);
or U25110 (N_25110,N_24860,N_21180);
nand U25111 (N_25111,N_23988,N_20711);
nor U25112 (N_25112,N_24839,N_24336);
or U25113 (N_25113,N_24071,N_21451);
nand U25114 (N_25114,N_21061,N_21105);
nor U25115 (N_25115,N_23266,N_22440);
xor U25116 (N_25116,N_22843,N_23355);
xor U25117 (N_25117,N_20635,N_21253);
nor U25118 (N_25118,N_24064,N_20949);
or U25119 (N_25119,N_23708,N_23756);
nor U25120 (N_25120,N_20270,N_22582);
nor U25121 (N_25121,N_22584,N_23937);
or U25122 (N_25122,N_20465,N_20474);
xnor U25123 (N_25123,N_22468,N_24327);
and U25124 (N_25124,N_23611,N_22902);
or U25125 (N_25125,N_20536,N_22748);
nor U25126 (N_25126,N_24994,N_23972);
nand U25127 (N_25127,N_20510,N_24179);
nand U25128 (N_25128,N_21538,N_21111);
xor U25129 (N_25129,N_24443,N_24728);
nand U25130 (N_25130,N_24513,N_23789);
and U25131 (N_25131,N_20084,N_24618);
nand U25132 (N_25132,N_21233,N_24439);
nand U25133 (N_25133,N_21054,N_22590);
or U25134 (N_25134,N_23664,N_23048);
nor U25135 (N_25135,N_21036,N_20583);
and U25136 (N_25136,N_23996,N_23594);
or U25137 (N_25137,N_23993,N_22731);
nand U25138 (N_25138,N_21400,N_20424);
nor U25139 (N_25139,N_23806,N_22682);
and U25140 (N_25140,N_21011,N_20996);
xnor U25141 (N_25141,N_22049,N_23547);
nand U25142 (N_25142,N_22576,N_24789);
nor U25143 (N_25143,N_24863,N_21148);
nor U25144 (N_25144,N_21455,N_24561);
xnor U25145 (N_25145,N_22377,N_23891);
or U25146 (N_25146,N_21939,N_20633);
nand U25147 (N_25147,N_20796,N_23537);
xor U25148 (N_25148,N_22239,N_22771);
or U25149 (N_25149,N_22213,N_24430);
xor U25150 (N_25150,N_22522,N_23623);
nand U25151 (N_25151,N_22117,N_21403);
nand U25152 (N_25152,N_23062,N_20733);
or U25153 (N_25153,N_23244,N_23782);
or U25154 (N_25154,N_21901,N_20416);
xnor U25155 (N_25155,N_22672,N_21971);
or U25156 (N_25156,N_22552,N_23274);
nand U25157 (N_25157,N_22766,N_23267);
or U25158 (N_25158,N_23797,N_24250);
or U25159 (N_25159,N_24840,N_21884);
nor U25160 (N_25160,N_21114,N_22196);
nand U25161 (N_25161,N_20190,N_21732);
or U25162 (N_25162,N_23826,N_21758);
or U25163 (N_25163,N_20606,N_23684);
or U25164 (N_25164,N_21119,N_24821);
or U25165 (N_25165,N_22941,N_24375);
nor U25166 (N_25166,N_22234,N_22918);
or U25167 (N_25167,N_23298,N_20130);
xnor U25168 (N_25168,N_20877,N_23591);
nand U25169 (N_25169,N_23958,N_22625);
nor U25170 (N_25170,N_22494,N_21280);
xor U25171 (N_25171,N_20335,N_22560);
nor U25172 (N_25172,N_21672,N_22168);
or U25173 (N_25173,N_20673,N_23245);
and U25174 (N_25174,N_21245,N_20286);
nor U25175 (N_25175,N_23468,N_21055);
nand U25176 (N_25176,N_24745,N_23172);
and U25177 (N_25177,N_23899,N_23000);
nor U25178 (N_25178,N_21260,N_22253);
and U25179 (N_25179,N_20980,N_22806);
nand U25180 (N_25180,N_22348,N_24615);
or U25181 (N_25181,N_22005,N_20997);
xor U25182 (N_25182,N_24288,N_22060);
and U25183 (N_25183,N_22739,N_22258);
or U25184 (N_25184,N_24132,N_21184);
and U25185 (N_25185,N_23314,N_22914);
or U25186 (N_25186,N_23706,N_22893);
nor U25187 (N_25187,N_22765,N_24537);
nor U25188 (N_25188,N_23750,N_24931);
nor U25189 (N_25189,N_23595,N_23470);
xnor U25190 (N_25190,N_20644,N_24729);
nand U25191 (N_25191,N_24173,N_24766);
nand U25192 (N_25192,N_23990,N_20707);
and U25193 (N_25193,N_21920,N_20594);
nand U25194 (N_25194,N_22572,N_21766);
nand U25195 (N_25195,N_24264,N_24293);
and U25196 (N_25196,N_23372,N_24580);
nor U25197 (N_25197,N_24919,N_24509);
nand U25198 (N_25198,N_21759,N_22891);
or U25199 (N_25199,N_24637,N_22782);
or U25200 (N_25200,N_22834,N_23603);
and U25201 (N_25201,N_24868,N_22082);
and U25202 (N_25202,N_21032,N_24150);
nor U25203 (N_25203,N_20072,N_22366);
nand U25204 (N_25204,N_21178,N_22394);
or U25205 (N_25205,N_23253,N_20201);
and U25206 (N_25206,N_23497,N_20002);
or U25207 (N_25207,N_20386,N_24330);
nand U25208 (N_25208,N_20621,N_23011);
or U25209 (N_25209,N_21832,N_22881);
and U25210 (N_25210,N_24302,N_20876);
xor U25211 (N_25211,N_21957,N_23788);
xnor U25212 (N_25212,N_22542,N_20841);
nor U25213 (N_25213,N_23814,N_21739);
nand U25214 (N_25214,N_21808,N_23521);
xor U25215 (N_25215,N_21588,N_23808);
or U25216 (N_25216,N_22303,N_20458);
nor U25217 (N_25217,N_20313,N_24398);
nand U25218 (N_25218,N_21583,N_23248);
and U25219 (N_25219,N_24679,N_20860);
or U25220 (N_25220,N_23607,N_23156);
xnor U25221 (N_25221,N_22249,N_20445);
nor U25222 (N_25222,N_24359,N_24888);
or U25223 (N_25223,N_23592,N_22455);
and U25224 (N_25224,N_22986,N_23387);
or U25225 (N_25225,N_24373,N_22164);
or U25226 (N_25226,N_20132,N_23859);
xnor U25227 (N_25227,N_24143,N_24086);
and U25228 (N_25228,N_22081,N_24680);
xor U25229 (N_25229,N_24958,N_20942);
or U25230 (N_25230,N_23214,N_21196);
and U25231 (N_25231,N_22710,N_21478);
nand U25232 (N_25232,N_23458,N_24569);
or U25233 (N_25233,N_24392,N_23747);
nor U25234 (N_25234,N_20303,N_21733);
nor U25235 (N_25235,N_23280,N_24796);
or U25236 (N_25236,N_21151,N_20282);
nand U25237 (N_25237,N_24354,N_22120);
or U25238 (N_25238,N_24490,N_21639);
or U25239 (N_25239,N_22163,N_22429);
xor U25240 (N_25240,N_21642,N_20588);
nand U25241 (N_25241,N_21270,N_23982);
xnor U25242 (N_25242,N_22577,N_24235);
or U25243 (N_25243,N_24943,N_24297);
xor U25244 (N_25244,N_20501,N_22664);
and U25245 (N_25245,N_20831,N_20010);
nor U25246 (N_25246,N_24164,N_20610);
and U25247 (N_25247,N_22639,N_21420);
or U25248 (N_25248,N_22727,N_22756);
xnor U25249 (N_25249,N_20682,N_24944);
nand U25250 (N_25250,N_22406,N_21968);
and U25251 (N_25251,N_20477,N_23906);
or U25252 (N_25252,N_24441,N_21089);
or U25253 (N_25253,N_23948,N_23358);
nor U25254 (N_25254,N_24220,N_24131);
and U25255 (N_25255,N_20328,N_22593);
or U25256 (N_25256,N_22221,N_20521);
or U25257 (N_25257,N_21100,N_24085);
nor U25258 (N_25258,N_23342,N_21296);
and U25259 (N_25259,N_23697,N_24609);
nor U25260 (N_25260,N_24393,N_24855);
and U25261 (N_25261,N_21816,N_20720);
or U25262 (N_25262,N_23392,N_20451);
or U25263 (N_25263,N_20053,N_24467);
and U25264 (N_25264,N_21993,N_24001);
nor U25265 (N_25265,N_22416,N_21415);
xnor U25266 (N_25266,N_22815,N_20784);
and U25267 (N_25267,N_20773,N_21950);
or U25268 (N_25268,N_22821,N_21696);
nor U25269 (N_25269,N_20783,N_21976);
and U25270 (N_25270,N_20350,N_23831);
and U25271 (N_25271,N_22975,N_22565);
and U25272 (N_25272,N_23668,N_21685);
nor U25273 (N_25273,N_24686,N_20717);
nor U25274 (N_25274,N_21108,N_22617);
and U25275 (N_25275,N_21173,N_22361);
nand U25276 (N_25276,N_20913,N_21368);
nand U25277 (N_25277,N_23111,N_21041);
and U25278 (N_25278,N_20738,N_24444);
xor U25279 (N_25279,N_23954,N_24877);
and U25280 (N_25280,N_23889,N_21386);
nand U25281 (N_25281,N_21885,N_24021);
nand U25282 (N_25282,N_23503,N_21408);
or U25283 (N_25283,N_23792,N_22957);
and U25284 (N_25284,N_24739,N_22033);
and U25285 (N_25285,N_22869,N_24560);
and U25286 (N_25286,N_22293,N_20261);
and U25287 (N_25287,N_20279,N_20242);
nor U25288 (N_25288,N_24898,N_21125);
nand U25289 (N_25289,N_24254,N_22812);
xor U25290 (N_25290,N_22200,N_20000);
nor U25291 (N_25291,N_22130,N_21038);
and U25292 (N_25292,N_22894,N_24818);
and U25293 (N_25293,N_20272,N_21571);
nor U25294 (N_25294,N_23629,N_20800);
and U25295 (N_25295,N_24205,N_24111);
and U25296 (N_25296,N_23434,N_24291);
or U25297 (N_25297,N_22344,N_20653);
nand U25298 (N_25298,N_24160,N_20497);
nor U25299 (N_25299,N_23634,N_24070);
or U25300 (N_25300,N_22959,N_20619);
and U25301 (N_25301,N_20539,N_21050);
nor U25302 (N_25302,N_20979,N_24167);
nand U25303 (N_25303,N_23628,N_21080);
or U25304 (N_25304,N_23015,N_20262);
or U25305 (N_25305,N_24420,N_22927);
xnor U25306 (N_25306,N_22479,N_21690);
and U25307 (N_25307,N_21877,N_21213);
or U25308 (N_25308,N_24915,N_22025);
nor U25309 (N_25309,N_24465,N_21508);
nor U25310 (N_25310,N_21567,N_22832);
or U25311 (N_25311,N_22282,N_22011);
and U25312 (N_25312,N_22744,N_21674);
or U25313 (N_25313,N_24685,N_21207);
nand U25314 (N_25314,N_22460,N_21342);
nor U25315 (N_25315,N_20086,N_22274);
nand U25316 (N_25316,N_22855,N_23440);
and U25317 (N_25317,N_21098,N_23288);
xor U25318 (N_25318,N_23905,N_23659);
or U25319 (N_25319,N_23730,N_23528);
nand U25320 (N_25320,N_21743,N_21164);
nand U25321 (N_25321,N_23545,N_20781);
nand U25322 (N_25322,N_22759,N_21666);
or U25323 (N_25323,N_20938,N_21444);
nand U25324 (N_25324,N_23325,N_23173);
and U25325 (N_25325,N_22219,N_21202);
xnor U25326 (N_25326,N_21314,N_22945);
or U25327 (N_25327,N_24017,N_21506);
nand U25328 (N_25328,N_20150,N_20441);
nor U25329 (N_25329,N_20125,N_21162);
and U25330 (N_25330,N_21077,N_23114);
xnor U25331 (N_25331,N_24920,N_22714);
xor U25332 (N_25332,N_23983,N_20074);
or U25333 (N_25333,N_20334,N_21479);
nand U25334 (N_25334,N_24464,N_23804);
or U25335 (N_25335,N_24407,N_22061);
nor U25336 (N_25336,N_22605,N_24110);
or U25337 (N_25337,N_23500,N_22359);
or U25338 (N_25338,N_23026,N_23694);
or U25339 (N_25339,N_23714,N_23239);
or U25340 (N_25340,N_20546,N_21012);
and U25341 (N_25341,N_24602,N_22086);
nor U25342 (N_25342,N_22983,N_20907);
xor U25343 (N_25343,N_22156,N_20558);
nor U25344 (N_25344,N_20809,N_20983);
and U25345 (N_25345,N_23981,N_21736);
nor U25346 (N_25346,N_20020,N_21263);
nand U25347 (N_25347,N_21596,N_21550);
nand U25348 (N_25348,N_24575,N_21128);
nand U25349 (N_25349,N_22773,N_21170);
nor U25350 (N_25350,N_21124,N_21545);
xnor U25351 (N_25351,N_21922,N_24523);
or U25352 (N_25352,N_21987,N_20404);
nand U25353 (N_25353,N_23332,N_23039);
and U25354 (N_25354,N_24962,N_21820);
nor U25355 (N_25355,N_21328,N_22382);
and U25356 (N_25356,N_21387,N_21051);
or U25357 (N_25357,N_24923,N_23335);
nor U25358 (N_25358,N_21355,N_23965);
xor U25359 (N_25359,N_20387,N_21088);
or U25360 (N_25360,N_21831,N_21842);
or U25361 (N_25361,N_20992,N_21874);
nand U25362 (N_25362,N_23508,N_22533);
nor U25363 (N_25363,N_22390,N_22925);
nand U25364 (N_25364,N_20482,N_21570);
nand U25365 (N_25365,N_22331,N_24995);
and U25366 (N_25366,N_20993,N_23907);
nor U25367 (N_25367,N_23422,N_24648);
nand U25368 (N_25368,N_24451,N_22814);
xnor U25369 (N_25369,N_22952,N_24874);
nand U25370 (N_25370,N_24300,N_20397);
and U25371 (N_25371,N_24469,N_21755);
and U25372 (N_25372,N_21299,N_24127);
nor U25373 (N_25373,N_23933,N_23702);
nor U25374 (N_25374,N_24304,N_23371);
nand U25375 (N_25375,N_20599,N_24579);
and U25376 (N_25376,N_23775,N_24557);
nand U25377 (N_25377,N_21285,N_22330);
or U25378 (N_25378,N_20500,N_22669);
xnor U25379 (N_25379,N_23834,N_22228);
nand U25380 (N_25380,N_22804,N_23226);
nand U25381 (N_25381,N_24075,N_22640);
nor U25382 (N_25382,N_20590,N_20897);
nand U25383 (N_25383,N_22441,N_22124);
xor U25384 (N_25384,N_22751,N_22009);
or U25385 (N_25385,N_22616,N_21416);
or U25386 (N_25386,N_20198,N_20975);
nor U25387 (N_25387,N_21424,N_22847);
nand U25388 (N_25388,N_21737,N_23771);
nor U25389 (N_25389,N_21802,N_22649);
nor U25390 (N_25390,N_20687,N_20540);
xnor U25391 (N_25391,N_24934,N_21074);
nand U25392 (N_25392,N_20495,N_22971);
and U25393 (N_25393,N_20880,N_21306);
xnor U25394 (N_25394,N_23718,N_20419);
nand U25395 (N_25395,N_24966,N_24140);
nor U25396 (N_25396,N_23976,N_23832);
nor U25397 (N_25397,N_24754,N_21425);
or U25398 (N_25398,N_21255,N_20776);
nor U25399 (N_25399,N_20830,N_24664);
or U25400 (N_25400,N_23210,N_20952);
or U25401 (N_25401,N_20339,N_24508);
or U25402 (N_25402,N_23203,N_21433);
nand U25403 (N_25403,N_24060,N_22929);
and U25404 (N_25404,N_22829,N_22524);
nor U25405 (N_25405,N_24084,N_22116);
or U25406 (N_25406,N_22694,N_23050);
xor U25407 (N_25407,N_20167,N_22601);
nor U25408 (N_25408,N_24011,N_23622);
nand U25409 (N_25409,N_22544,N_20485);
nand U25410 (N_25410,N_21738,N_23240);
xnor U25411 (N_25411,N_24760,N_23146);
xnor U25412 (N_25412,N_22093,N_24362);
or U25413 (N_25413,N_23390,N_24222);
nand U25414 (N_25414,N_20658,N_21106);
nor U25415 (N_25415,N_23548,N_22127);
nor U25416 (N_25416,N_20185,N_20355);
and U25417 (N_25417,N_24517,N_21064);
nand U25418 (N_25418,N_22670,N_20129);
and U25419 (N_25419,N_21703,N_22871);
and U25420 (N_25420,N_20889,N_21026);
and U25421 (N_25421,N_24244,N_22875);
or U25422 (N_25422,N_24324,N_22618);
xor U25423 (N_25423,N_23557,N_22725);
xor U25424 (N_25424,N_24847,N_24031);
nor U25425 (N_25425,N_20326,N_23336);
xnor U25426 (N_25426,N_22141,N_20088);
and U25427 (N_25427,N_22421,N_22398);
nand U25428 (N_25428,N_24651,N_23292);
nor U25429 (N_25429,N_20461,N_21345);
or U25430 (N_25430,N_22944,N_21322);
and U25431 (N_25431,N_24295,N_21945);
nor U25432 (N_25432,N_21211,N_24276);
and U25433 (N_25433,N_20677,N_23721);
or U25434 (N_25434,N_24281,N_21069);
nand U25435 (N_25435,N_22492,N_21134);
and U25436 (N_25436,N_23057,N_22596);
or U25437 (N_25437,N_20535,N_23080);
nor U25438 (N_25438,N_20693,N_23686);
nand U25439 (N_25439,N_21916,N_23469);
or U25440 (N_25440,N_23699,N_21194);
or U25441 (N_25441,N_21087,N_22963);
nand U25442 (N_25442,N_22525,N_21520);
and U25443 (N_25443,N_21401,N_21323);
xor U25444 (N_25444,N_24364,N_23901);
or U25445 (N_25445,N_23916,N_22317);
nand U25446 (N_25446,N_20499,N_23561);
and U25447 (N_25447,N_20176,N_21025);
xor U25448 (N_25448,N_21259,N_22177);
nor U25449 (N_25449,N_24768,N_21572);
nor U25450 (N_25450,N_23307,N_23363);
nor U25451 (N_25451,N_21562,N_22750);
and U25452 (N_25452,N_21407,N_20814);
and U25453 (N_25453,N_21302,N_22798);
or U25454 (N_25454,N_20067,N_23185);
and U25455 (N_25455,N_20265,N_22289);
or U25456 (N_25456,N_22497,N_24015);
and U25457 (N_25457,N_24023,N_23587);
and U25458 (N_25458,N_23546,N_21232);
and U25459 (N_25459,N_20926,N_22559);
or U25460 (N_25460,N_21191,N_23709);
nor U25461 (N_25461,N_24128,N_24639);
nor U25462 (N_25462,N_24411,N_23612);
nor U25463 (N_25463,N_21671,N_22961);
nand U25464 (N_25464,N_22449,N_24113);
or U25465 (N_25465,N_21395,N_21174);
nor U25466 (N_25466,N_20799,N_23737);
nand U25467 (N_25467,N_24503,N_20819);
and U25468 (N_25468,N_22186,N_23734);
nand U25469 (N_25469,N_20453,N_23558);
nor U25470 (N_25470,N_24296,N_22658);
nor U25471 (N_25471,N_21068,N_20280);
and U25472 (N_25472,N_20353,N_21843);
nand U25473 (N_25473,N_24193,N_20049);
or U25474 (N_25474,N_23516,N_21856);
and U25475 (N_25475,N_24619,N_24376);
or U25476 (N_25476,N_20371,N_22973);
or U25477 (N_25477,N_23078,N_20632);
and U25478 (N_25478,N_24546,N_22325);
and U25479 (N_25479,N_22058,N_21057);
nand U25480 (N_25480,N_24762,N_23896);
nand U25481 (N_25481,N_22212,N_20565);
xor U25482 (N_25482,N_23934,N_23250);
and U25483 (N_25483,N_21300,N_21560);
nand U25484 (N_25484,N_23817,N_24916);
nor U25485 (N_25485,N_23564,N_23915);
and U25486 (N_25486,N_20835,N_24960);
nand U25487 (N_25487,N_21139,N_21573);
nor U25488 (N_25488,N_22529,N_22423);
and U25489 (N_25489,N_20848,N_23282);
and U25490 (N_25490,N_22436,N_22048);
xor U25491 (N_25491,N_23550,N_23984);
and U25492 (N_25492,N_20244,N_21189);
or U25493 (N_25493,N_20931,N_22439);
nor U25494 (N_25494,N_21153,N_20963);
nand U25495 (N_25495,N_21798,N_20026);
xnor U25496 (N_25496,N_24769,N_21557);
and U25497 (N_25497,N_24628,N_21313);
or U25498 (N_25498,N_21684,N_21385);
nand U25499 (N_25499,N_20252,N_24526);
and U25500 (N_25500,N_23295,N_21231);
or U25501 (N_25501,N_20472,N_23157);
nand U25502 (N_25502,N_20612,N_20764);
nand U25503 (N_25503,N_23106,N_24879);
xor U25504 (N_25504,N_22919,N_24487);
nand U25505 (N_25505,N_22510,N_22690);
nor U25506 (N_25506,N_20691,N_21882);
nor U25507 (N_25507,N_24846,N_23898);
and U25508 (N_25508,N_23511,N_20912);
and U25509 (N_25509,N_21973,N_21655);
nor U25510 (N_25510,N_22237,N_24701);
nand U25511 (N_25511,N_21205,N_21866);
xor U25512 (N_25512,N_20439,N_22599);
nor U25513 (N_25513,N_20204,N_20669);
nand U25514 (N_25514,N_24092,N_21470);
nor U25515 (N_25515,N_21195,N_24691);
and U25516 (N_25516,N_22292,N_23149);
nand U25517 (N_25517,N_24683,N_22109);
nor U25518 (N_25518,N_21549,N_20713);
nor U25519 (N_25519,N_22953,N_20972);
xnor U25520 (N_25520,N_23141,N_21719);
nand U25521 (N_25521,N_24123,N_23190);
xnor U25522 (N_25522,N_21953,N_20810);
and U25523 (N_25523,N_22612,N_20791);
and U25524 (N_25524,N_23081,N_21131);
or U25525 (N_25525,N_23609,N_21801);
and U25526 (N_25526,N_20686,N_23989);
and U25527 (N_25527,N_20217,N_20778);
nor U25528 (N_25528,N_21783,N_20173);
or U25529 (N_25529,N_23932,N_21181);
xnor U25530 (N_25530,N_21946,N_21770);
nand U25531 (N_25531,N_21465,N_21157);
and U25532 (N_25532,N_22733,N_22837);
xnor U25533 (N_25533,N_23328,N_22098);
nor U25534 (N_25534,N_23496,N_22085);
xor U25535 (N_25535,N_20358,N_22064);
or U25536 (N_25536,N_24016,N_21615);
nor U25537 (N_25537,N_22991,N_21986);
nand U25538 (N_25538,N_21163,N_24682);
or U25539 (N_25539,N_24308,N_22346);
or U25540 (N_25540,N_22335,N_20164);
nand U25541 (N_25541,N_20166,N_21459);
nor U25542 (N_25542,N_23308,N_22826);
or U25543 (N_25543,N_23327,N_22385);
nand U25544 (N_25544,N_24219,N_23179);
nand U25545 (N_25545,N_21500,N_20742);
nor U25546 (N_25546,N_20449,N_21552);
nand U25547 (N_25547,N_22448,N_21037);
nor U25548 (N_25548,N_20861,N_21492);
or U25549 (N_25549,N_23324,N_20113);
or U25550 (N_25550,N_21595,N_20023);
and U25551 (N_25551,N_20464,N_20255);
nand U25552 (N_25552,N_24640,N_22614);
nand U25553 (N_25553,N_21653,N_23602);
nand U25554 (N_25554,N_23258,N_24456);
or U25555 (N_25555,N_22801,N_23339);
nor U25556 (N_25556,N_22379,N_20695);
or U25557 (N_25557,N_21564,N_23158);
nor U25558 (N_25558,N_23405,N_22089);
and U25559 (N_25559,N_21179,N_24942);
or U25560 (N_25560,N_23066,N_21018);
and U25561 (N_25561,N_24187,N_21132);
xor U25562 (N_25562,N_21099,N_20920);
or U25563 (N_25563,N_21351,N_24929);
and U25564 (N_25564,N_24022,N_22541);
nor U25565 (N_25565,N_21498,N_23689);
nand U25566 (N_25566,N_23876,N_22171);
nor U25567 (N_25567,N_20797,N_20118);
and U25568 (N_25568,N_22286,N_24521);
nand U25569 (N_25569,N_23783,N_20595);
nand U25570 (N_25570,N_21610,N_21568);
nand U25571 (N_25571,N_20417,N_21347);
and U25572 (N_25572,N_20824,N_21223);
or U25573 (N_25573,N_22570,N_20066);
nand U25574 (N_25574,N_23456,N_22467);
and U25575 (N_25575,N_24183,N_21242);
or U25576 (N_25576,N_22946,N_24791);
nand U25577 (N_25577,N_23058,N_24834);
xnor U25578 (N_25578,N_24172,N_24352);
nand U25579 (N_25579,N_20758,N_24518);
or U25580 (N_25580,N_23919,N_24852);
nand U25581 (N_25581,N_22712,N_24667);
and U25582 (N_25582,N_24059,N_22504);
and U25583 (N_25583,N_22738,N_23223);
nor U25584 (N_25584,N_22554,N_24974);
nor U25585 (N_25585,N_20999,N_23882);
nand U25586 (N_25586,N_20988,N_20575);
nor U25587 (N_25587,N_20122,N_20479);
nand U25588 (N_25588,N_21217,N_20904);
nand U25589 (N_25589,N_24644,N_21225);
and U25590 (N_25590,N_23204,N_23202);
nand U25591 (N_25591,N_21103,N_22091);
nand U25592 (N_25592,N_23432,N_21118);
or U25593 (N_25593,N_23928,N_21254);
nor U25594 (N_25594,N_24115,N_22592);
and U25595 (N_25595,N_23751,N_23719);
or U25596 (N_25596,N_23819,N_21485);
nor U25597 (N_25597,N_20301,N_22442);
xor U25598 (N_25598,N_21445,N_22789);
and U25599 (N_25599,N_21555,N_20227);
or U25600 (N_25600,N_21772,N_20712);
nor U25601 (N_25601,N_22452,N_20447);
nor U25602 (N_25602,N_24385,N_24321);
nor U25603 (N_25603,N_24180,N_24299);
and U25604 (N_25604,N_20019,N_22024);
nand U25605 (N_25605,N_24340,N_23032);
or U25606 (N_25606,N_20807,N_24216);
and U25607 (N_25607,N_20647,N_24759);
and U25608 (N_25608,N_22323,N_20718);
nand U25609 (N_25609,N_23429,N_20863);
or U25610 (N_25610,N_23463,N_24472);
nand U25611 (N_25611,N_22195,N_20249);
nand U25612 (N_25612,N_23921,N_22280);
and U25613 (N_25613,N_24409,N_23024);
and U25614 (N_25614,N_22236,N_22706);
nor U25615 (N_25615,N_24389,N_23970);
or U25616 (N_25616,N_24214,N_21219);
nor U25617 (N_25617,N_24824,N_22043);
nor U25618 (N_25618,N_22666,N_20361);
nand U25619 (N_25619,N_24658,N_20577);
nor U25620 (N_25620,N_21835,N_23563);
or U25621 (N_25621,N_21286,N_20945);
or U25622 (N_25622,N_22932,N_22707);
or U25623 (N_25623,N_22791,N_20769);
nand U25624 (N_25624,N_22378,N_24067);
and U25625 (N_25625,N_23523,N_23260);
nand U25626 (N_25626,N_23660,N_22063);
or U25627 (N_25627,N_23123,N_23121);
and U25628 (N_25628,N_22030,N_21350);
and U25629 (N_25629,N_20480,N_23908);
nand U25630 (N_25630,N_23009,N_21951);
xnor U25631 (N_25631,N_22907,N_24417);
nand U25632 (N_25632,N_22571,N_20133);
xor U25633 (N_25633,N_24935,N_21984);
and U25634 (N_25634,N_22092,N_22732);
nor U25635 (N_25635,N_22321,N_23480);
or U25636 (N_25636,N_21989,N_20700);
nor U25637 (N_25637,N_23018,N_20205);
nor U25638 (N_25638,N_23192,N_21632);
nor U25639 (N_25639,N_24710,N_20478);
and U25640 (N_25640,N_24097,N_23485);
nor U25641 (N_25641,N_22934,N_23740);
nor U25642 (N_25642,N_20545,N_20930);
or U25643 (N_25643,N_22051,N_22624);
or U25644 (N_25644,N_22708,N_24582);
nor U25645 (N_25645,N_24955,N_22050);
nor U25646 (N_25646,N_24862,N_24450);
nand U25647 (N_25647,N_22107,N_21629);
nor U25648 (N_25648,N_22140,N_21049);
nor U25649 (N_25649,N_23777,N_24119);
or U25650 (N_25650,N_21393,N_23213);
nor U25651 (N_25651,N_24024,N_22375);
nand U25652 (N_25652,N_24624,N_23688);
nor U25653 (N_25653,N_24795,N_23909);
and U25654 (N_25654,N_20348,N_22065);
nor U25655 (N_25655,N_23581,N_24066);
or U25656 (N_25656,N_22659,N_20079);
or U25657 (N_25657,N_22100,N_21965);
and U25658 (N_25658,N_24591,N_21767);
and U25659 (N_25659,N_22476,N_23412);
xor U25660 (N_25660,N_20574,N_23604);
nand U25661 (N_25661,N_23509,N_21079);
xnor U25662 (N_25662,N_22685,N_20729);
or U25663 (N_25663,N_22161,N_22352);
nand U25664 (N_25664,N_21094,N_21692);
nand U25665 (N_25665,N_23847,N_22471);
and U25666 (N_25666,N_23035,N_24989);
nand U25667 (N_25667,N_21826,N_21461);
nand U25668 (N_25668,N_20354,N_24440);
and U25669 (N_25669,N_20529,N_20843);
nand U25670 (N_25670,N_24379,N_21329);
or U25671 (N_25671,N_24061,N_22762);
nor U25672 (N_25672,N_23535,N_22222);
or U25673 (N_25673,N_20774,N_20618);
nor U25674 (N_25674,N_24857,N_22886);
nor U25675 (N_25675,N_22059,N_23312);
nor U25676 (N_25676,N_21643,N_22122);
nor U25677 (N_25677,N_21857,N_20381);
nand U25678 (N_25678,N_24474,N_24985);
or U25679 (N_25679,N_21366,N_21053);
nand U25680 (N_25680,N_22501,N_23864);
and U25681 (N_25681,N_23566,N_23092);
nor U25682 (N_25682,N_21252,N_24524);
nor U25683 (N_25683,N_20378,N_20329);
xnor U25684 (N_25684,N_22247,N_20391);
and U25685 (N_25685,N_23060,N_22967);
nand U25686 (N_25686,N_22469,N_24121);
and U25687 (N_25687,N_23268,N_23389);
xor U25688 (N_25688,N_24053,N_20767);
nand U25689 (N_25689,N_21764,N_24318);
nand U25690 (N_25690,N_24570,N_23341);
xnor U25691 (N_25691,N_22300,N_22686);
nor U25692 (N_25692,N_20165,N_22668);
nand U25693 (N_25693,N_21988,N_23757);
or U25694 (N_25694,N_22193,N_21411);
nor U25695 (N_25695,N_22989,N_20116);
nand U25696 (N_25696,N_21587,N_24290);
and U25697 (N_25697,N_22155,N_23770);
nor U25698 (N_25698,N_22447,N_20298);
and U25699 (N_25699,N_22676,N_21071);
nor U25700 (N_25700,N_21172,N_22817);
or U25701 (N_25701,N_21226,N_24372);
and U25702 (N_25702,N_24395,N_21398);
xnor U25703 (N_25703,N_22717,N_22555);
or U25704 (N_25704,N_24197,N_23145);
nor U25705 (N_25705,N_22106,N_21936);
and U25706 (N_25706,N_24181,N_21405);
nand U25707 (N_25707,N_20174,N_20874);
xor U25708 (N_25708,N_23108,N_21126);
and U25709 (N_25709,N_24705,N_22662);
nand U25710 (N_25710,N_23212,N_22962);
nor U25711 (N_25711,N_23251,N_20512);
or U25712 (N_25712,N_20857,N_21853);
nor U25713 (N_25713,N_22638,N_22285);
nor U25714 (N_25714,N_21959,N_21358);
and U25715 (N_25715,N_24695,N_24032);
or U25716 (N_25716,N_21625,N_24043);
nor U25717 (N_25717,N_23310,N_22786);
nand U25718 (N_25718,N_23388,N_22936);
nor U25719 (N_25719,N_22697,N_24735);
nor U25720 (N_25720,N_23624,N_20380);
nand U25721 (N_25721,N_23633,N_21239);
or U25722 (N_25722,N_22242,N_21530);
nand U25723 (N_25723,N_22793,N_20550);
nand U25724 (N_25724,N_20425,N_23135);
nor U25725 (N_25725,N_20413,N_23601);
nor U25726 (N_25726,N_23839,N_21609);
and U25727 (N_25727,N_20645,N_23753);
nand U25728 (N_25728,N_23583,N_20188);
xor U25729 (N_25729,N_21035,N_20015);
or U25730 (N_25730,N_22924,N_24319);
xnor U25731 (N_25731,N_22790,N_20177);
or U25732 (N_25732,N_21360,N_24153);
nand U25733 (N_25733,N_24702,N_24926);
nand U25734 (N_25734,N_24617,N_24170);
and U25735 (N_25735,N_24771,N_20723);
nor U25736 (N_25736,N_24952,N_21700);
nor U25737 (N_25737,N_22261,N_21378);
or U25738 (N_25738,N_24087,N_21943);
xnor U25739 (N_25739,N_24156,N_22597);
nor U25740 (N_25740,N_23890,N_21897);
nand U25741 (N_25741,N_21418,N_20193);
and U25742 (N_25742,N_23885,N_23283);
or U25743 (N_25743,N_23229,N_24638);
xnor U25744 (N_25744,N_20143,N_22250);
nor U25745 (N_25745,N_24289,N_20184);
or U25746 (N_25746,N_23316,N_23103);
and U25747 (N_25747,N_22667,N_24812);
and U25748 (N_25748,N_22495,N_21660);
nor U25749 (N_25749,N_20037,N_23075);
or U25750 (N_25750,N_22438,N_20524);
and U25751 (N_25751,N_21975,N_20273);
and U25752 (N_25752,N_20502,N_23529);
nand U25753 (N_25753,N_22265,N_23553);
or U25754 (N_25754,N_21379,N_23723);
and U25755 (N_25755,N_21204,N_22151);
nor U25756 (N_25756,N_21464,N_21869);
or U25757 (N_25757,N_20243,N_23690);
nor U25758 (N_25758,N_21698,N_23873);
nor U25759 (N_25759,N_22878,N_22129);
nor U25760 (N_25760,N_20951,N_24257);
nand U25761 (N_25761,N_24305,N_21929);
nand U25762 (N_25762,N_23536,N_21811);
or U25763 (N_25763,N_23648,N_20801);
nand U25764 (N_25764,N_23575,N_23863);
nand U25765 (N_25765,N_20128,N_24231);
nand U25766 (N_25766,N_24063,N_24777);
xor U25767 (N_25767,N_23365,N_24232);
nor U25768 (N_25768,N_20071,N_22631);
or U25769 (N_25769,N_21705,N_23029);
and U25770 (N_25770,N_20821,N_20703);
nand U25771 (N_25771,N_24104,N_22889);
or U25772 (N_25772,N_21494,N_20316);
nor U25773 (N_25773,N_22110,N_22768);
and U25774 (N_25774,N_23656,N_21117);
and U25775 (N_25775,N_20838,N_24833);
nor U25776 (N_25776,N_23674,N_22337);
or U25777 (N_25777,N_24422,N_22974);
nor U25778 (N_25778,N_24844,N_23764);
and U25779 (N_25779,N_20170,N_21717);
xnor U25780 (N_25780,N_20956,N_20965);
nor U25781 (N_25781,N_23247,N_22512);
xor U25782 (N_25782,N_24100,N_24787);
nor U25783 (N_25783,N_23874,N_23687);
and U25784 (N_25784,N_23947,N_22132);
or U25785 (N_25785,N_23980,N_22646);
or U25786 (N_25786,N_23552,N_24815);
and U25787 (N_25787,N_23918,N_23437);
or U25788 (N_25788,N_22969,N_24099);
nand U25789 (N_25789,N_24347,N_20234);
nand U25790 (N_25790,N_22742,N_21683);
or U25791 (N_25791,N_22233,N_22018);
or U25792 (N_25792,N_23713,N_23054);
nor U25793 (N_25793,N_23348,N_21185);
nand U25794 (N_25794,N_21156,N_21291);
nor U25795 (N_25795,N_24437,N_24148);
nor U25796 (N_25796,N_21824,N_23761);
and U25797 (N_25797,N_23269,N_20611);
or U25798 (N_25798,N_20739,N_23790);
or U25799 (N_25799,N_24399,N_20388);
nand U25800 (N_25800,N_20368,N_21447);
nor U25801 (N_25801,N_23849,N_20525);
nor U25802 (N_25802,N_21579,N_20728);
nand U25803 (N_25803,N_21917,N_23744);
or U25804 (N_25804,N_24360,N_20957);
nor U25805 (N_25805,N_20976,N_23334);
or U25806 (N_25806,N_24583,N_22964);
or U25807 (N_25807,N_22816,N_20440);
nor U25808 (N_25808,N_22860,N_20247);
nor U25809 (N_25809,N_21507,N_23279);
or U25810 (N_25810,N_22266,N_20825);
nor U25811 (N_25811,N_21889,N_21014);
nand U25812 (N_25812,N_21898,N_23287);
or U25813 (N_25813,N_23850,N_24954);
or U25814 (N_25814,N_23554,N_20189);
nand U25815 (N_25815,N_24149,N_24635);
nor U25816 (N_25816,N_21353,N_20620);
and U25817 (N_25817,N_24185,N_23183);
and U25818 (N_25818,N_20491,N_22270);
and U25819 (N_25819,N_20159,N_23063);
and U25820 (N_25820,N_24724,N_20580);
nand U25821 (N_25821,N_21534,N_24406);
and U25822 (N_25822,N_22620,N_21556);
nor U25823 (N_25823,N_20586,N_20598);
or U25824 (N_25824,N_22935,N_23733);
nand U25825 (N_25825,N_23652,N_22741);
xor U25826 (N_25826,N_21136,N_23477);
nor U25827 (N_25827,N_21283,N_22078);
and U25828 (N_25828,N_22550,N_23522);
and U25829 (N_25829,N_22904,N_24343);
nand U25830 (N_25830,N_20853,N_24917);
or U25831 (N_25831,N_23119,N_20716);
or U25832 (N_25832,N_22154,N_22800);
nand U25833 (N_25833,N_21201,N_23171);
nand U25834 (N_25834,N_23964,N_23577);
nand U25835 (N_25835,N_21496,N_24421);
nor U25836 (N_25836,N_22142,N_21473);
nor U25837 (N_25837,N_24936,N_22119);
nor U25838 (N_25838,N_24845,N_21369);
nor U25839 (N_25839,N_23518,N_21215);
and U25840 (N_25840,N_23022,N_21578);
xnor U25841 (N_25841,N_22496,N_21359);
xor U25842 (N_25842,N_23914,N_22077);
and U25843 (N_25843,N_21076,N_24008);
or U25844 (N_25844,N_23049,N_21646);
or U25845 (N_25845,N_21007,N_23020);
nand U25846 (N_25846,N_20833,N_23163);
or U25847 (N_25847,N_23820,N_24269);
xor U25848 (N_25848,N_20837,N_21844);
nor U25849 (N_25849,N_24809,N_20001);
nor U25850 (N_25850,N_21086,N_20622);
and U25851 (N_25851,N_20726,N_24887);
nand U25852 (N_25852,N_24174,N_23065);
nand U25853 (N_25853,N_24287,N_21354);
nand U25854 (N_25854,N_21841,N_23130);
nor U25855 (N_25855,N_20937,N_23768);
and U25856 (N_25856,N_23491,N_24082);
and U25857 (N_25857,N_21540,N_24573);
or U25858 (N_25858,N_23643,N_22622);
nand U25859 (N_25859,N_24656,N_22519);
nand U25860 (N_25860,N_21310,N_21812);
nand U25861 (N_25861,N_24961,N_23286);
nand U25862 (N_25862,N_22118,N_23599);
xor U25863 (N_25863,N_23313,N_23679);
nor U25864 (N_25864,N_24741,N_22966);
nor U25865 (N_25865,N_20967,N_20410);
xor U25866 (N_25866,N_24652,N_23331);
xnor U25867 (N_25867,N_23127,N_21166);
or U25868 (N_25868,N_24038,N_24013);
nor U25869 (N_25869,N_24366,N_23128);
and U25870 (N_25870,N_22999,N_22692);
nor U25871 (N_25871,N_20457,N_21474);
and U25872 (N_25872,N_23867,N_21734);
or U25873 (N_25873,N_24209,N_23161);
or U25874 (N_25874,N_23871,N_20487);
and U25875 (N_25875,N_20870,N_21029);
nand U25876 (N_25876,N_22774,N_24550);
and U25877 (N_25877,N_21017,N_20320);
or U25878 (N_25878,N_20106,N_23155);
or U25879 (N_25879,N_24820,N_22034);
nor U25880 (N_25880,N_22165,N_22288);
nor U25881 (N_25881,N_22458,N_20259);
xor U25882 (N_25882,N_20640,N_23488);
nor U25883 (N_25883,N_22036,N_23290);
nor U25884 (N_25884,N_22008,N_24718);
nor U25885 (N_25885,N_22125,N_22055);
and U25886 (N_25886,N_22681,N_24719);
nand U25887 (N_25887,N_22456,N_21913);
xor U25888 (N_25888,N_20052,N_24382);
or U25889 (N_25889,N_22811,N_20278);
and U25890 (N_25890,N_23370,N_21697);
or U25891 (N_25891,N_20562,N_22430);
or U25892 (N_25892,N_24309,N_20947);
nand U25893 (N_25893,N_24800,N_22099);
nand U25894 (N_25894,N_23068,N_20542);
or U25895 (N_25895,N_21544,N_24457);
nand U25896 (N_25896,N_22278,N_24761);
nand U25897 (N_25897,N_20637,N_23868);
nand U25898 (N_25898,N_20109,N_20077);
and U25899 (N_25899,N_22763,N_24757);
and U25900 (N_25900,N_20970,N_21633);
nand U25901 (N_25901,N_22673,N_24326);
and U25902 (N_25902,N_22851,N_22980);
nor U25903 (N_25903,N_24612,N_23099);
or U25904 (N_25904,N_24495,N_23395);
or U25905 (N_25905,N_22858,N_21788);
or U25906 (N_25906,N_22937,N_21575);
nor U25907 (N_25907,N_24114,N_24186);
nand U25908 (N_25908,N_23033,N_21890);
nand U25909 (N_25909,N_24587,N_22632);
and U25910 (N_25910,N_22502,N_23544);
xor U25911 (N_25911,N_23584,N_23769);
nor U25912 (N_25912,N_23354,N_23110);
nor U25913 (N_25913,N_20342,N_20033);
nor U25914 (N_25914,N_24538,N_21397);
nor U25915 (N_25915,N_23705,N_22134);
and U25916 (N_25916,N_20839,N_22340);
nor U25917 (N_25917,N_21900,N_23252);
or U25918 (N_25918,N_24665,N_23259);
and U25919 (N_25919,N_24567,N_22121);
nor U25920 (N_25920,N_24122,N_23105);
and U25921 (N_25921,N_24776,N_20299);
nand U25922 (N_25922,N_24904,N_24897);
nor U25923 (N_25923,N_23922,N_24556);
and U25924 (N_25924,N_24981,N_21192);
and U25925 (N_25925,N_21248,N_21175);
nand U25926 (N_25926,N_21948,N_20114);
or U25927 (N_25927,N_23727,N_22730);
nand U25928 (N_25928,N_23381,N_21430);
xor U25929 (N_25929,N_21644,N_23653);
and U25930 (N_25930,N_20815,N_23169);
nor U25931 (N_25931,N_21435,N_24418);
or U25932 (N_25932,N_23739,N_23071);
or U25933 (N_25933,N_22339,N_23272);
xor U25934 (N_25934,N_23333,N_24873);
nor U25935 (N_25935,N_22209,N_23900);
nand U25936 (N_25936,N_24913,N_23228);
nand U25937 (N_25937,N_23840,N_23630);
nor U25938 (N_25938,N_24112,N_24836);
nand U25939 (N_25939,N_22283,N_23047);
nand U25940 (N_25940,N_24229,N_24221);
nand U25941 (N_25941,N_24322,N_24826);
xor U25942 (N_25942,N_21039,N_20105);
or U25943 (N_25943,N_24262,N_24853);
nand U25944 (N_25944,N_24374,N_21009);
and U25945 (N_25945,N_21316,N_21336);
nand U25946 (N_25946,N_20063,N_20236);
nor U25947 (N_25947,N_24566,N_20393);
xnor U25948 (N_25948,N_23798,N_24607);
or U25949 (N_25949,N_23425,N_20846);
nand U25950 (N_25950,N_22805,N_24764);
and U25951 (N_25951,N_20055,N_21450);
nor U25952 (N_25952,N_21851,N_21486);
or U25953 (N_25953,N_21264,N_23373);
or U25954 (N_25954,N_21636,N_24212);
and U25955 (N_25955,N_21399,N_24348);
and U25956 (N_25956,N_24415,N_20924);
or U25957 (N_25957,N_22810,N_24325);
or U25958 (N_25958,N_24162,N_24646);
and U25959 (N_25959,N_23217,N_24892);
and U25960 (N_25960,N_24120,N_20324);
nor U25961 (N_25961,N_22206,N_22758);
and U25962 (N_25962,N_21062,N_21301);
or U25963 (N_25963,N_21338,N_23678);
or U25964 (N_25964,N_24419,N_20469);
or U25965 (N_25965,N_23610,N_22302);
or U25966 (N_25966,N_21293,N_22393);
xnor U25967 (N_25967,N_24522,N_20083);
nand U25968 (N_25968,N_20559,N_24380);
nand U25969 (N_25969,N_22518,N_24642);
xor U25970 (N_25970,N_21104,N_21756);
and U25971 (N_25971,N_22573,N_24144);
or U25972 (N_25972,N_22890,N_24386);
nor U25973 (N_25973,N_20409,N_21631);
nand U25974 (N_25974,N_20916,N_23109);
nand U25975 (N_25975,N_22785,N_22947);
nand U25976 (N_25976,N_21875,N_24206);
nor U25977 (N_25977,N_24540,N_24057);
nand U25978 (N_25978,N_24323,N_22928);
and U25979 (N_25979,N_21159,N_23994);
nor U25980 (N_25980,N_22466,N_24520);
or U25981 (N_25981,N_22305,N_21412);
nor U25982 (N_25982,N_22530,N_23472);
and U25983 (N_25983,N_22689,N_21852);
and U25984 (N_25984,N_20859,N_21849);
or U25985 (N_25985,N_23366,N_22031);
and U25986 (N_25986,N_22840,N_24306);
nand U25987 (N_25987,N_20310,N_22022);
xnor U25988 (N_25988,N_20675,N_20375);
xnor U25989 (N_25989,N_22532,N_23927);
nand U25990 (N_25990,N_24048,N_24041);
xor U25991 (N_25991,N_21865,N_24218);
and U25992 (N_25992,N_24941,N_21774);
nand U25993 (N_25993,N_22995,N_24723);
xor U25994 (N_25994,N_22231,N_24089);
or U25995 (N_25995,N_21761,N_21101);
nor U25996 (N_25996,N_22802,N_20646);
or U25997 (N_25997,N_20233,N_22679);
nor U25998 (N_25998,N_20757,N_21093);
nand U25999 (N_25999,N_24654,N_20958);
nand U26000 (N_26000,N_23821,N_21290);
and U26001 (N_26001,N_23220,N_24447);
and U26002 (N_26002,N_21715,N_23693);
and U26003 (N_26003,N_24611,N_23326);
nand U26004 (N_26004,N_23100,N_20210);
and U26005 (N_26005,N_20139,N_22691);
nor U26006 (N_26006,N_22695,N_24026);
and U26007 (N_26007,N_20104,N_21097);
nor U26008 (N_26008,N_21115,N_20030);
and U26009 (N_26009,N_20119,N_22068);
nor U26010 (N_26010,N_23419,N_23555);
nand U26011 (N_26011,N_21475,N_21505);
nand U26012 (N_26012,N_20456,N_22574);
nor U26013 (N_26013,N_23862,N_22876);
and U26014 (N_26014,N_23017,N_20402);
nor U26015 (N_26015,N_20422,N_22316);
or U26016 (N_26016,N_24674,N_24661);
or U26017 (N_26017,N_24650,N_21789);
or U26018 (N_26018,N_24717,N_22844);
nand U26019 (N_26019,N_21724,N_22551);
xnor U26020 (N_26020,N_24252,N_23216);
nand U26021 (N_26021,N_20450,N_21985);
and U26022 (N_26022,N_24633,N_23238);
nor U26023 (N_26023,N_22087,N_23303);
and U26024 (N_26024,N_23973,N_20507);
xor U26025 (N_26025,N_23237,N_23368);
xnor U26026 (N_26026,N_23102,N_23181);
and U26027 (N_26027,N_23445,N_21868);
and U26028 (N_26028,N_24571,N_22260);
or U26029 (N_26029,N_20763,N_20305);
or U26030 (N_26030,N_24914,N_20579);
nand U26031 (N_26031,N_20470,N_20625);
nor U26032 (N_26032,N_20211,N_22580);
or U26033 (N_26033,N_22426,N_21121);
nor U26034 (N_26034,N_20110,N_21519);
nand U26035 (N_26035,N_21352,N_22543);
or U26036 (N_26036,N_24554,N_20840);
and U26037 (N_26037,N_23802,N_22764);
nand U26038 (N_26038,N_24731,N_23696);
or U26039 (N_26039,N_23655,N_22108);
or U26040 (N_26040,N_23430,N_20107);
or U26041 (N_26041,N_23464,N_24458);
nand U26042 (N_26042,N_23070,N_20933);
nor U26043 (N_26043,N_22726,N_24693);
xor U26044 (N_26044,N_20961,N_22648);
nand U26045 (N_26045,N_24310,N_21276);
xor U26046 (N_26046,N_23681,N_23883);
nor U26047 (N_26047,N_21614,N_21749);
xnor U26048 (N_26048,N_21744,N_20182);
nand U26049 (N_26049,N_22480,N_22038);
and U26050 (N_26050,N_21165,N_21613);
xor U26051 (N_26051,N_20462,N_20898);
nor U26052 (N_26052,N_23570,N_23360);
or U26053 (N_26053,N_22054,N_24978);
or U26054 (N_26054,N_23378,N_20731);
or U26055 (N_26055,N_22521,N_21315);
nand U26056 (N_26056,N_20141,N_24527);
or U26057 (N_26057,N_24045,N_20029);
and U26058 (N_26058,N_21059,N_21208);
nor U26059 (N_26059,N_20035,N_20827);
nor U26060 (N_26060,N_20561,N_22147);
and U26061 (N_26061,N_22955,N_20571);
nand U26062 (N_26062,N_23076,N_20082);
nand U26063 (N_26063,N_24435,N_21488);
nor U26064 (N_26064,N_24502,N_23069);
or U26065 (N_26065,N_22079,N_20494);
nor U26066 (N_26066,N_22841,N_20221);
and U26067 (N_26067,N_20438,N_24631);
and U26068 (N_26068,N_20901,N_23542);
nand U26069 (N_26069,N_24886,N_22488);
nand U26070 (N_26070,N_23424,N_23182);
or U26071 (N_26071,N_22749,N_22432);
and U26072 (N_26072,N_20089,N_24480);
and U26073 (N_26073,N_20553,N_24471);
xor U26074 (N_26074,N_22954,N_24479);
nor U26075 (N_26075,N_24614,N_20987);
nand U26076 (N_26076,N_24808,N_22041);
and U26077 (N_26077,N_24251,N_24867);
nand U26078 (N_26078,N_23125,N_22514);
nand U26079 (N_26079,N_20349,N_23540);
nand U26080 (N_26080,N_23627,N_22201);
or U26081 (N_26081,N_21060,N_24466);
nand U26082 (N_26082,N_23941,N_21085);
and U26083 (N_26083,N_20971,N_20314);
nor U26084 (N_26084,N_20054,N_23741);
or U26085 (N_26085,N_21961,N_22813);
nand U26086 (N_26086,N_23087,N_22257);
or U26087 (N_26087,N_22701,N_22032);
and U26088 (N_26088,N_23573,N_21477);
nor U26089 (N_26089,N_20881,N_20587);
nand U26090 (N_26090,N_22415,N_22678);
nand U26091 (N_26091,N_23006,N_20531);
nor U26092 (N_26092,N_24049,N_21908);
and U26093 (N_26093,N_23853,N_22796);
xnor U26094 (N_26094,N_24804,N_21361);
nor U26095 (N_26095,N_22000,N_22752);
and U26096 (N_26096,N_23846,N_22734);
nor U26097 (N_26097,N_21434,N_23435);
nand U26098 (N_26098,N_21680,N_20097);
nor U26099 (N_26099,N_20179,N_21070);
or U26100 (N_26100,N_23957,N_21129);
nand U26101 (N_26101,N_21490,N_24058);
nand U26102 (N_26102,N_20013,N_22493);
nand U26103 (N_26103,N_22433,N_24514);
or U26104 (N_26104,N_22114,N_24147);
or U26105 (N_26105,N_24312,N_22218);
and U26106 (N_26106,N_22487,N_20929);
or U26107 (N_26107,N_22548,N_23961);
nand U26108 (N_26108,N_21589,N_23902);
nand U26109 (N_26109,N_21974,N_21503);
nor U26110 (N_26110,N_21991,N_21307);
and U26111 (N_26111,N_23801,N_23977);
and U26112 (N_26112,N_21246,N_23159);
and U26113 (N_26113,N_20850,N_20744);
or U26114 (N_26114,N_23059,N_20775);
nand U26115 (N_26115,N_24829,N_23374);
nand U26116 (N_26116,N_22419,N_21067);
nor U26117 (N_26117,N_21458,N_20294);
nand U26118 (N_26118,N_24907,N_23710);
and U26119 (N_26119,N_20552,N_20448);
and U26120 (N_26120,N_20795,N_22080);
or U26121 (N_26121,N_20538,N_23013);
xnor U26122 (N_26122,N_22037,N_20503);
and U26123 (N_26123,N_22511,N_23301);
nand U26124 (N_26124,N_20080,N_23337);
nor U26125 (N_26125,N_20124,N_20994);
nand U26126 (N_26126,N_23246,N_23446);
nand U26127 (N_26127,N_20615,N_22647);
nor U26128 (N_26128,N_24263,N_23036);
or U26129 (N_26129,N_24188,N_21436);
and U26130 (N_26130,N_21930,N_23089);
and U26131 (N_26131,N_24712,N_24199);
xor U26132 (N_26132,N_23943,N_22019);
and U26133 (N_26133,N_20936,N_23767);
and U26134 (N_26134,N_22149,N_23893);
and U26135 (N_26135,N_22405,N_24999);
and U26136 (N_26136,N_21333,N_21371);
and U26137 (N_26137,N_24811,N_20341);
and U26138 (N_26138,N_24154,N_21873);
or U26139 (N_26139,N_23177,N_20921);
and U26140 (N_26140,N_22520,N_21269);
xor U26141 (N_26141,N_22410,N_21637);
or U26142 (N_26142,N_22958,N_22227);
or U26143 (N_26143,N_23153,N_22047);
nand U26144 (N_26144,N_21709,N_23836);
or U26145 (N_26145,N_20572,N_24224);
and U26146 (N_26146,N_20263,N_22338);
nand U26147 (N_26147,N_22882,N_21996);
nor U26148 (N_26148,N_24630,N_21586);
nand U26149 (N_26149,N_21647,N_21977);
and U26150 (N_26150,N_24158,N_20842);
nand U26151 (N_26151,N_23042,N_24384);
xor U26152 (N_26152,N_22716,N_20008);
nand U26153 (N_26153,N_24753,N_20822);
nor U26154 (N_26154,N_21998,N_20385);
and U26155 (N_26155,N_24645,N_20338);
nor U26156 (N_26156,N_20708,N_23530);
nand U26157 (N_26157,N_20851,N_23673);
nand U26158 (N_26158,N_21082,N_24331);
or U26159 (N_26159,N_20288,N_20508);
nor U26160 (N_26160,N_20309,N_22016);
or U26161 (N_26161,N_22857,N_23309);
or U26162 (N_26162,N_20092,N_20284);
and U26163 (N_26163,N_20973,N_21150);
nand U26164 (N_26164,N_22276,N_24211);
or U26165 (N_26165,N_23787,N_23671);
nor U26166 (N_26166,N_24905,N_20534);
nor U26167 (N_26167,N_21431,N_20974);
nor U26168 (N_26168,N_20732,N_24613);
or U26169 (N_26169,N_24329,N_23762);
xor U26170 (N_26170,N_21370,N_24979);
and U26171 (N_26171,N_22729,N_23311);
or U26172 (N_26172,N_20427,N_21796);
and U26173 (N_26173,N_21787,N_22852);
and U26174 (N_26174,N_21548,N_20702);
nor U26175 (N_26175,N_24298,N_24233);
and U26176 (N_26176,N_22898,N_23276);
and U26177 (N_26177,N_22336,N_23582);
and U26178 (N_26178,N_21840,N_20683);
nor U26179 (N_26179,N_20098,N_23857);
nand U26180 (N_26180,N_20366,N_22979);
xnor U26181 (N_26181,N_23828,N_20607);
or U26182 (N_26182,N_23255,N_22799);
xnor U26183 (N_26183,N_20578,N_21367);
and U26184 (N_26184,N_20352,N_24165);
or U26185 (N_26185,N_20556,N_20157);
and U26186 (N_26186,N_20073,N_24807);
nand U26187 (N_26187,N_23559,N_22371);
and U26188 (N_26188,N_20679,N_21502);
and U26189 (N_26189,N_22754,N_21410);
or U26190 (N_26190,N_21394,N_22252);
nand U26191 (N_26191,N_20384,N_22435);
and U26192 (N_26192,N_23541,N_24881);
xor U26193 (N_26193,N_24029,N_24623);
or U26194 (N_26194,N_23598,N_20629);
or U26195 (N_26195,N_24077,N_24752);
nand U26196 (N_26196,N_21978,N_22824);
nor U26197 (N_26197,N_20435,N_20196);
nor U26198 (N_26198,N_21933,N_22627);
nand U26199 (N_26199,N_24511,N_23386);
nand U26200 (N_26200,N_20140,N_23649);
nand U26201 (N_26201,N_20798,N_20293);
or U26202 (N_26202,N_23227,N_21383);
and U26203 (N_26203,N_22178,N_24828);
nor U26204 (N_26204,N_22254,N_20081);
nor U26205 (N_26205,N_24822,N_21404);
nor U26206 (N_26206,N_24080,N_20332);
nand U26207 (N_26207,N_24529,N_21542);
or U26208 (N_26208,N_20694,N_20789);
nand U26209 (N_26209,N_22635,N_22781);
or U26210 (N_26210,N_21598,N_22783);
nand U26211 (N_26211,N_21525,N_24758);
nand U26212 (N_26212,N_21675,N_22880);
nor U26213 (N_26213,N_21529,N_24893);
or U26214 (N_26214,N_24714,N_21380);
or U26215 (N_26215,N_24969,N_23030);
nand U26216 (N_26216,N_23164,N_21906);
or U26217 (N_26217,N_20858,N_21982);
or U26218 (N_26218,N_23270,N_22067);
nor U26219 (N_26219,N_20161,N_22343);
xnor U26220 (N_26220,N_21803,N_23254);
nand U26221 (N_26221,N_24774,N_20828);
or U26222 (N_26222,N_23088,N_22723);
xnor U26223 (N_26223,N_23072,N_21272);
nor U26224 (N_26224,N_21382,N_23439);
and U26225 (N_26225,N_24697,N_20111);
and U26226 (N_26226,N_24986,N_20476);
or U26227 (N_26227,N_24367,N_24433);
or U26228 (N_26228,N_24725,N_24161);
or U26229 (N_26229,N_21522,N_20785);
and U26230 (N_26230,N_24255,N_21152);
nor U26231 (N_26231,N_24094,N_22459);
nand U26232 (N_26232,N_21904,N_24657);
nand U26233 (N_26233,N_22943,N_21523);
nor U26234 (N_26234,N_22629,N_24987);
or U26235 (N_26235,N_22324,N_23041);
nand U26236 (N_26236,N_22443,N_20420);
and U26237 (N_26237,N_20101,N_24478);
nor U26238 (N_26238,N_23824,N_20199);
nand U26239 (N_26239,N_24204,N_24670);
or U26240 (N_26240,N_24046,N_22357);
or U26241 (N_26241,N_20662,N_24971);
xor U26242 (N_26242,N_21923,N_21224);
nand U26243 (N_26243,N_23763,N_22113);
nand U26244 (N_26244,N_23136,N_23150);
nand U26245 (N_26245,N_21096,N_23479);
or U26246 (N_26246,N_23654,N_23329);
nand U26247 (N_26247,N_21257,N_22537);
or U26248 (N_26248,N_22621,N_20977);
nor U26249 (N_26249,N_20533,N_20704);
or U26250 (N_26250,N_23707,N_21543);
nand U26251 (N_26251,N_23829,N_24848);
and U26252 (N_26252,N_20398,N_21845);
and U26253 (N_26253,N_20319,N_21515);
or U26254 (N_26254,N_20616,N_24706);
and U26255 (N_26255,N_21599,N_20289);
nor U26256 (N_26256,N_22722,N_20882);
nor U26257 (N_26257,N_20549,N_22942);
and U26258 (N_26258,N_23700,N_24563);
xnor U26259 (N_26259,N_20820,N_21292);
nand U26260 (N_26260,N_20246,N_23385);
or U26261 (N_26261,N_22345,N_22241);
nand U26262 (N_26262,N_24095,N_21648);
or U26263 (N_26263,N_20617,N_24589);
nand U26264 (N_26264,N_21249,N_21147);
nor U26265 (N_26265,N_21221,N_24436);
nor U26266 (N_26266,N_23357,N_22262);
xnor U26267 (N_26267,N_20095,N_20115);
or U26268 (N_26268,N_20689,N_24548);
nand U26269 (N_26269,N_20428,N_24361);
nand U26270 (N_26270,N_24885,N_21227);
nand U26271 (N_26271,N_24698,N_22095);
or U26272 (N_26272,N_23452,N_22607);
nor U26273 (N_26273,N_24856,N_23460);
nand U26274 (N_26274,N_20186,N_22454);
or U26275 (N_26275,N_21034,N_23118);
nor U26276 (N_26276,N_24201,N_20245);
and U26277 (N_26277,N_23097,N_22281);
or U26278 (N_26278,N_23886,N_21716);
nor U26279 (N_26279,N_22131,N_23019);
xor U26280 (N_26280,N_23728,N_23493);
and U26281 (N_26281,N_24669,N_23682);
and U26282 (N_26282,N_22397,N_20787);
xnor U26283 (N_26283,N_21768,N_20948);
or U26284 (N_26284,N_22776,N_23402);
xnor U26285 (N_26285,N_24707,N_22921);
xnor U26286 (N_26286,N_21251,N_23224);
nand U26287 (N_26287,N_22863,N_22372);
xnor U26288 (N_26288,N_21472,N_20207);
xor U26289 (N_26289,N_21776,N_23257);
nand U26290 (N_26290,N_23474,N_23515);
nor U26291 (N_26291,N_23305,N_21334);
nand U26292 (N_26292,N_20614,N_20044);
or U26293 (N_26293,N_21140,N_24349);
nand U26294 (N_26294,N_21863,N_24107);
xor U26295 (N_26295,N_22998,N_20254);
nor U26296 (N_26296,N_21116,N_21695);
nor U26297 (N_26297,N_22162,N_23129);
and U26298 (N_26298,N_22103,N_21848);
nand U26299 (N_26299,N_23551,N_23188);
or U26300 (N_26300,N_24632,N_23672);
and U26301 (N_26301,N_24342,N_22845);
and U26302 (N_26302,N_22503,N_20762);
nand U26303 (N_26303,N_24565,N_23666);
or U26304 (N_26304,N_21804,N_20911);
nand U26305 (N_26305,N_22803,N_22674);
nor U26306 (N_26306,N_21693,N_24091);
nand U26307 (N_26307,N_21309,N_22071);
and U26308 (N_26308,N_21177,N_21970);
or U26309 (N_26309,N_21003,N_22135);
nand U26310 (N_26310,N_23780,N_20471);
nor U26311 (N_26311,N_22332,N_21273);
and U26312 (N_26312,N_24189,N_20923);
or U26313 (N_26313,N_24039,N_22506);
xnor U26314 (N_26314,N_24751,N_22445);
nor U26315 (N_26315,N_22505,N_24736);
nor U26316 (N_26316,N_22848,N_22655);
xor U26317 (N_26317,N_24079,N_23315);
nor U26318 (N_26318,N_20959,N_22540);
or U26319 (N_26319,N_24236,N_22306);
nor U26320 (N_26320,N_21002,N_22897);
or U26321 (N_26321,N_24694,N_23382);
or U26322 (N_26322,N_21621,N_21994);
nor U26323 (N_26323,N_20808,N_24891);
or U26324 (N_26324,N_21084,N_22587);
and U26325 (N_26325,N_24634,N_20688);
or U26326 (N_26326,N_22900,N_22978);
and U26327 (N_26327,N_23784,N_20727);
xnor U26328 (N_26328,N_23852,N_23992);
nand U26329 (N_26329,N_21576,N_21109);
nand U26330 (N_26330,N_22204,N_22585);
nand U26331 (N_26331,N_23187,N_24788);
nor U26332 (N_26332,N_24426,N_24675);
nor U26333 (N_26333,N_24286,N_21340);
nand U26334 (N_26334,N_21829,N_22069);
nor U26335 (N_26335,N_20915,N_21083);
and U26336 (N_26336,N_23635,N_24230);
nand U26337 (N_26337,N_23510,N_20698);
or U26338 (N_26338,N_22846,N_23519);
xnor U26339 (N_26339,N_20004,N_24740);
and U26340 (N_26340,N_20197,N_23426);
xor U26341 (N_26341,N_22434,N_22696);
xnor U26342 (N_26342,N_22720,N_22740);
and U26343 (N_26343,N_23695,N_20816);
nand U26344 (N_26344,N_23507,N_20523);
nor U26345 (N_26345,N_24678,N_24484);
or U26346 (N_26346,N_22075,N_21439);
nor U26347 (N_26347,N_23760,N_23860);
xnor U26348 (N_26348,N_20557,N_24176);
and U26349 (N_26349,N_23569,N_20878);
and U26350 (N_26350,N_21457,N_20365);
xnor U26351 (N_26351,N_21122,N_21827);
and U26352 (N_26352,N_24505,N_21337);
xor U26353 (N_26353,N_22606,N_20879);
or U26354 (N_26354,N_21102,N_20146);
nor U26355 (N_26355,N_20057,N_24234);
or U26356 (N_26356,N_22198,N_20264);
nand U26357 (N_26357,N_22035,N_24983);
nor U26358 (N_26358,N_24311,N_23935);
xor U26359 (N_26359,N_24413,N_24870);
nor U26360 (N_26360,N_20364,N_24599);
nor U26361 (N_26361,N_20505,N_20667);
nand U26362 (N_26362,N_24608,N_21212);
nand U26363 (N_26363,N_20943,N_23884);
and U26364 (N_26364,N_23524,N_21748);
nand U26365 (N_26365,N_21817,N_22515);
nand U26366 (N_26366,N_21577,N_24858);
or U26367 (N_26367,N_23475,N_23538);
nor U26368 (N_26368,N_23241,N_24096);
or U26369 (N_26369,N_21837,N_23494);
and U26370 (N_26370,N_23256,N_20226);
nand U26371 (N_26371,N_21203,N_24932);
xor U26372 (N_26372,N_22004,N_24475);
nor U26373 (N_26373,N_21854,N_20027);
and U26374 (N_26374,N_23637,N_22901);
and U26375 (N_26375,N_23619,N_21938);
and U26376 (N_26376,N_24355,N_24785);
or U26377 (N_26377,N_21501,N_23571);
nor U26378 (N_26378,N_23512,N_23870);
nor U26379 (N_26379,N_23646,N_21678);
nor U26380 (N_26380,N_23004,N_20902);
or U26381 (N_26381,N_20300,N_20181);
or U26382 (N_26382,N_23966,N_23249);
and U26383 (N_26383,N_21604,N_24586);
and U26384 (N_26384,N_20291,N_24977);
or U26385 (N_26385,N_22425,N_24088);
nand U26386 (N_26386,N_20307,N_23218);
nand U26387 (N_26387,N_20061,N_20705);
and U26388 (N_26388,N_22173,N_22229);
xor U26389 (N_26389,N_24733,N_24069);
xnor U26390 (N_26390,N_22486,N_23746);
nand U26391 (N_26391,N_23572,N_24258);
or U26392 (N_26392,N_24346,N_22391);
or U26393 (N_26393,N_20434,N_24790);
and U26394 (N_26394,N_21926,N_21066);
and U26395 (N_26395,N_22719,N_21275);
and U26396 (N_26396,N_24253,N_20087);
nand U26397 (N_26397,N_22187,N_22268);
nor U26398 (N_26398,N_23892,N_21078);
and U26399 (N_26399,N_21809,N_22819);
xor U26400 (N_26400,N_24534,N_24315);
nand U26401 (N_26401,N_23848,N_24198);
nor U26402 (N_26402,N_20761,N_22909);
and U26403 (N_26403,N_21830,N_22746);
and U26404 (N_26404,N_20379,N_24098);
nand U26405 (N_26405,N_20985,N_24709);
or U26406 (N_26406,N_22396,N_21325);
nand U26407 (N_26407,N_24980,N_24074);
nor U26408 (N_26408,N_22988,N_21489);
nand U26409 (N_26409,N_22578,N_24245);
nand U26410 (N_26410,N_21481,N_20017);
nor U26411 (N_26411,N_23779,N_22527);
nand U26412 (N_26412,N_21658,N_24854);
nor U26413 (N_26413,N_21935,N_22809);
or U26414 (N_26414,N_24345,N_21043);
or U26415 (N_26415,N_23404,N_20396);
or U26416 (N_26416,N_20903,N_22992);
and U26417 (N_26417,N_24108,N_20802);
nand U26418 (N_26418,N_22224,N_24547);
or U26419 (N_26419,N_24483,N_20108);
and U26420 (N_26420,N_22328,N_24659);
and U26421 (N_26421,N_23651,N_22354);
and U26422 (N_26422,N_24228,N_20436);
nand U26423 (N_26423,N_24203,N_24763);
and U26424 (N_26424,N_20039,N_22698);
and U26425 (N_26425,N_22428,N_22166);
xnor U26426 (N_26426,N_23923,N_23376);
or U26427 (N_26427,N_23411,N_24703);
nor U26428 (N_26428,N_23067,N_20152);
nand U26429 (N_26429,N_22972,N_20737);
nand U26430 (N_26430,N_20064,N_23803);
xor U26431 (N_26431,N_24152,N_22994);
or U26432 (N_26432,N_21954,N_24912);
nor U26433 (N_26433,N_23207,N_23796);
nand U26434 (N_26434,N_23618,N_21800);
or U26435 (N_26435,N_23897,N_24688);
xor U26436 (N_26436,N_23144,N_23356);
nand U26437 (N_26437,N_24009,N_21547);
or U26438 (N_26438,N_24014,N_22483);
nor U26439 (N_26439,N_22591,N_23486);
or U26440 (N_26440,N_24677,N_22770);
and U26441 (N_26441,N_24446,N_21594);
nand U26442 (N_26442,N_20369,N_21565);
nor U26443 (N_26443,N_21331,N_22023);
or U26444 (N_26444,N_23526,N_23196);
or U26445 (N_26445,N_22136,N_22408);
nand U26446 (N_26446,N_24792,N_20235);
and U26447 (N_26447,N_22015,N_21063);
nand U26448 (N_26448,N_24213,N_20909);
nand U26449 (N_26449,N_20519,N_24925);
and U26450 (N_26450,N_21541,N_22825);
or U26451 (N_26451,N_20681,N_20287);
or U26452 (N_26452,N_24040,N_22420);
xor U26453 (N_26453,N_23197,N_22400);
or U26454 (N_26454,N_21514,N_24459);
or U26455 (N_26455,N_24827,N_24938);
or U26456 (N_26456,N_21626,N_22538);
nand U26457 (N_26457,N_22175,N_24453);
nor U26458 (N_26458,N_22478,N_22567);
xnor U26459 (N_26459,N_23991,N_21775);
nor U26460 (N_26460,N_24414,N_20408);
xor U26461 (N_26461,N_24721,N_21228);
and U26462 (N_26462,N_22562,N_23056);
or U26463 (N_26463,N_24700,N_23951);
or U26464 (N_26464,N_21944,N_21707);
nor U26465 (N_26465,N_24090,N_20543);
and U26466 (N_26466,N_24078,N_24237);
xor U26467 (N_26467,N_24425,N_20817);
and U26468 (N_26468,N_23304,N_23986);
and U26469 (N_26469,N_21220,N_22528);
or U26470 (N_26470,N_22076,N_21168);
or U26471 (N_26471,N_23805,N_24238);
and U26472 (N_26472,N_23698,N_24906);
nand U26473 (N_26473,N_20530,N_22090);
or U26474 (N_26474,N_20032,N_24817);
or U26475 (N_26475,N_23176,N_23613);
nor U26476 (N_26476,N_22619,N_22226);
nor U26477 (N_26477,N_24223,N_22320);
or U26478 (N_26478,N_22643,N_22062);
nor U26479 (N_26479,N_21421,N_22220);
nand U26480 (N_26480,N_20481,N_21375);
or U26481 (N_26481,N_23338,N_23632);
or U26482 (N_26482,N_23436,N_20202);
nand U26483 (N_26483,N_23265,N_20636);
nand U26484 (N_26484,N_24655,N_20582);
and U26485 (N_26485,N_21903,N_20759);
and U26486 (N_26486,N_24390,N_24831);
nand U26487 (N_26487,N_24190,N_21046);
or U26488 (N_26488,N_21584,N_22531);
and U26489 (N_26489,N_24668,N_20567);
xor U26490 (N_26490,N_21000,N_23638);
nand U26491 (N_26491,N_21305,N_20660);
nand U26492 (N_26492,N_20006,N_22411);
or U26493 (N_26493,N_20906,N_22401);
xnor U26494 (N_26494,N_23359,N_21819);
or U26495 (N_26495,N_21130,N_24984);
nand U26496 (N_26496,N_23407,N_24488);
xor U26497 (N_26497,N_23393,N_20144);
or U26498 (N_26498,N_24512,N_23351);
xnor U26499 (N_26499,N_23318,N_22490);
nand U26500 (N_26500,N_23534,N_21362);
or U26501 (N_26501,N_23944,N_24397);
or U26502 (N_26502,N_23670,N_22042);
and U26503 (N_26503,N_22409,N_21659);
or U26504 (N_26504,N_24696,N_20304);
or U26505 (N_26505,N_21638,N_20331);
or U26506 (N_26506,N_21045,N_22517);
xnor U26507 (N_26507,N_21454,N_24900);
nor U26508 (N_26508,N_20135,N_20290);
or U26509 (N_26509,N_23827,N_20661);
or U26510 (N_26510,N_24543,N_23658);
nor U26511 (N_26511,N_23722,N_23012);
and U26512 (N_26512,N_24600,N_21344);
and U26513 (N_26513,N_22353,N_20584);
nor U26514 (N_26514,N_23556,N_23567);
nor U26515 (N_26515,N_21905,N_23143);
and U26516 (N_26516,N_24445,N_24610);
xnor U26517 (N_26517,N_20389,N_24240);
and U26518 (N_26518,N_23663,N_20171);
and U26519 (N_26519,N_23726,N_21389);
or U26520 (N_26520,N_24195,N_23285);
xor U26521 (N_26521,N_24832,N_24734);
nor U26522 (N_26522,N_24939,N_22308);
nand U26523 (N_26523,N_21199,N_21236);
and U26524 (N_26524,N_24797,N_20794);
nand U26525 (N_26525,N_20297,N_24671);
or U26526 (N_26526,N_22461,N_20984);
or U26527 (N_26527,N_23098,N_21001);
xor U26528 (N_26528,N_24948,N_20554);
and U26529 (N_26529,N_21713,N_23104);
and U26530 (N_26530,N_22183,N_24793);
and U26531 (N_26531,N_23650,N_20147);
and U26532 (N_26532,N_22778,N_24460);
nor U26533 (N_26533,N_21652,N_20241);
or U26534 (N_26534,N_23946,N_20120);
nand U26535 (N_26535,N_23910,N_21883);
and U26536 (N_26536,N_22027,N_22913);
or U26537 (N_26537,N_24536,N_22215);
nand U26538 (N_26538,N_21805,N_22052);
nor U26539 (N_26539,N_21952,N_22568);
nand U26540 (N_26540,N_24396,N_24555);
and U26541 (N_26541,N_24991,N_23716);
nor U26542 (N_26542,N_21384,N_23809);
or U26543 (N_26543,N_24146,N_23096);
or U26544 (N_26544,N_23807,N_20513);
nand U26545 (N_26545,N_21990,N_22777);
xnor U26546 (N_26546,N_20407,N_20463);
or U26547 (N_26547,N_22029,N_22295);
and U26548 (N_26548,N_21429,N_20684);
or U26549 (N_26549,N_22747,N_20910);
nand U26550 (N_26550,N_24770,N_22403);
nor U26551 (N_26551,N_22602,N_21858);
and U26552 (N_26552,N_22787,N_23887);
nand U26553 (N_26553,N_21044,N_23122);
nand U26554 (N_26554,N_21727,N_21510);
nor U26555 (N_26555,N_21004,N_24317);
nor U26556 (N_26556,N_21821,N_20443);
nor U26557 (N_26557,N_23302,N_24957);
xnor U26558 (N_26558,N_24876,N_22199);
nor U26559 (N_26559,N_21590,N_21365);
and U26560 (N_26560,N_21019,N_22595);
and U26561 (N_26561,N_21483,N_21887);
or U26562 (N_26562,N_20935,N_20075);
nor U26563 (N_26563,N_24044,N_21092);
xor U26564 (N_26564,N_21941,N_20145);
and U26565 (N_26565,N_23038,N_20322);
nand U26566 (N_26566,N_22651,N_20748);
nor U26567 (N_26567,N_20544,N_24968);
nor U26568 (N_26568,N_22364,N_21907);
nand U26569 (N_26569,N_24872,N_21617);
or U26570 (N_26570,N_21899,N_23492);
or U26571 (N_26571,N_23278,N_21013);
and U26572 (N_26572,N_23597,N_24427);
nor U26573 (N_26573,N_23499,N_22794);
or U26574 (N_26574,N_21460,N_24260);
xnor U26575 (N_26575,N_22388,N_21825);
and U26576 (N_26576,N_23403,N_21528);
nor U26577 (N_26577,N_23952,N_24970);
or U26578 (N_26578,N_21769,N_21815);
nand U26579 (N_26579,N_20187,N_23574);
xor U26580 (N_26580,N_24303,N_21284);
or U26581 (N_26581,N_23929,N_23517);
or U26582 (N_26582,N_24062,N_20117);
nand U26583 (N_26583,N_22508,N_21925);
nand U26584 (N_26584,N_23685,N_24519);
nand U26585 (N_26585,N_22545,N_21343);
xor U26586 (N_26586,N_21142,N_24405);
nor U26587 (N_26587,N_22105,N_23639);
nand U26588 (N_26588,N_23209,N_24019);
nor U26589 (N_26589,N_22304,N_24138);
nor U26590 (N_26590,N_21406,N_22240);
and U26591 (N_26591,N_22414,N_20968);
nand U26592 (N_26592,N_20946,N_23045);
nor U26593 (N_26593,N_20012,N_21754);
and U26594 (N_26594,N_21422,N_24175);
or U26595 (N_26595,N_20696,N_24636);
and U26596 (N_26596,N_23838,N_24462);
and U26597 (N_26597,N_20219,N_21006);
nand U26598 (N_26598,N_20414,N_23527);
nand U26599 (N_26599,N_23858,N_23415);
xor U26600 (N_26600,N_20022,N_20932);
nor U26601 (N_26601,N_21850,N_20460);
or U26602 (N_26602,N_20005,N_21704);
xor U26603 (N_26603,N_23837,N_20154);
and U26604 (N_26604,N_20400,N_24813);
xnor U26605 (N_26605,N_24129,N_21861);
or U26606 (N_26606,N_22862,N_24755);
and U26607 (N_26607,N_23589,N_20832);
and U26608 (N_26608,N_21966,N_22926);
or U26609 (N_26609,N_24182,N_22111);
or U26610 (N_26610,N_22598,N_20492);
or U26611 (N_26611,N_23380,N_20426);
and U26612 (N_26612,N_20169,N_20172);
or U26613 (N_26613,N_23815,N_22355);
nand U26614 (N_26614,N_23772,N_21005);
and U26615 (N_26615,N_24552,N_21138);
nor U26616 (N_26616,N_20648,N_22499);
nand U26617 (N_26617,N_21532,N_22569);
nor U26618 (N_26618,N_21997,N_21591);
or U26619 (N_26619,N_24081,N_24604);
and U26620 (N_26620,N_21640,N_21558);
nand U26621 (N_26621,N_23786,N_22547);
nand U26622 (N_26622,N_23400,N_23856);
nor U26623 (N_26623,N_22384,N_21010);
and U26624 (N_26624,N_20591,N_20302);
xor U26625 (N_26625,N_23454,N_22820);
and U26626 (N_26626,N_22684,N_22279);
or U26627 (N_26627,N_22792,N_22899);
or U26628 (N_26628,N_24135,N_24625);
nand U26629 (N_26629,N_24408,N_20399);
or U26630 (N_26630,N_24353,N_20065);
nor U26631 (N_26631,N_24780,N_24799);
xnor U26632 (N_26632,N_20867,N_21878);
xnor U26633 (N_26633,N_22711,N_21963);
xnor U26634 (N_26634,N_24933,N_20253);
nor U26635 (N_26635,N_24184,N_22637);
nor U26636 (N_26636,N_23005,N_22102);
nor U26637 (N_26637,N_24387,N_24501);
and U26638 (N_26638,N_20760,N_22399);
and U26639 (N_26639,N_24225,N_22298);
nand U26640 (N_26640,N_21551,N_22713);
and U26641 (N_26641,N_23021,N_21607);
nand U26642 (N_26642,N_24489,N_21554);
and U26643 (N_26643,N_21670,N_21872);
nor U26644 (N_26644,N_23785,N_22633);
and U26645 (N_26645,N_20978,N_21265);
or U26646 (N_26646,N_24003,N_21580);
and U26647 (N_26647,N_21356,N_21919);
or U26648 (N_26648,N_20337,N_20372);
and U26649 (N_26649,N_22735,N_23617);
and U26650 (N_26650,N_23879,N_24779);
and U26651 (N_26651,N_22417,N_24320);
nor U26652 (N_26652,N_22534,N_22188);
nand U26653 (N_26653,N_23676,N_24902);
xor U26654 (N_26654,N_21710,N_24109);
and U26655 (N_26655,N_23418,N_22230);
xor U26656 (N_26656,N_20811,N_21888);
xnor U26657 (N_26657,N_24909,N_21438);
and U26658 (N_26658,N_20628,N_21127);
nor U26659 (N_26659,N_22660,N_22780);
xor U26660 (N_26660,N_23383,N_20526);
or U26661 (N_26661,N_22350,N_21169);
or U26662 (N_26662,N_23364,N_20312);
xnor U26663 (N_26663,N_20532,N_20650);
xnor U26664 (N_26664,N_21559,N_22208);
nor U26665 (N_26665,N_22671,N_23086);
nor U26666 (N_26666,N_23084,N_20891);
nand U26667 (N_26667,N_21912,N_20069);
nand U26668 (N_26668,N_20306,N_20137);
or U26669 (N_26669,N_21193,N_24279);
xor U26670 (N_26670,N_24055,N_21860);
and U26671 (N_26671,N_20444,N_20927);
nor U26672 (N_26672,N_23667,N_21056);
or U26673 (N_26673,N_21627,N_20323);
nand U26674 (N_26674,N_20772,N_21417);
or U26675 (N_26675,N_21753,N_21964);
nor U26676 (N_26676,N_22703,N_24037);
nor U26677 (N_26677,N_22312,N_22677);
or U26678 (N_26678,N_23367,N_21497);
nor U26679 (N_26679,N_23969,N_24864);
nor U26680 (N_26680,N_24998,N_22322);
or U26681 (N_26681,N_20051,N_24545);
nand U26682 (N_26682,N_21020,N_20248);
nand U26683 (N_26683,N_24620,N_20674);
nor U26684 (N_26684,N_21833,N_23101);
or U26685 (N_26685,N_22808,N_21075);
nand U26686 (N_26686,N_22475,N_22159);
nand U26687 (N_26687,N_21437,N_20657);
or U26688 (N_26688,N_24692,N_22549);
nand U26689 (N_26689,N_20624,N_22101);
and U26690 (N_26690,N_24226,N_22895);
nor U26691 (N_26691,N_22683,N_23513);
nor U26692 (N_26692,N_22950,N_22938);
or U26693 (N_26693,N_20382,N_20036);
or U26694 (N_26694,N_24371,N_23031);
nand U26695 (N_26695,N_21167,N_21701);
and U26696 (N_26696,N_24468,N_20347);
or U26697 (N_26697,N_23115,N_23725);
nand U26698 (N_26698,N_21531,N_24485);
xor U26699 (N_26699,N_21274,N_22313);
or U26700 (N_26700,N_22309,N_23199);
nand U26701 (N_26701,N_23142,N_20076);
and U26702 (N_26702,N_21894,N_23813);
nand U26703 (N_26703,N_21321,N_23151);
and U26704 (N_26704,N_20269,N_24510);
and U26705 (N_26705,N_21981,N_21327);
xor U26706 (N_26706,N_24400,N_24559);
and U26707 (N_26707,N_23998,N_24277);
nand U26708 (N_26708,N_23978,N_22523);
or U26709 (N_26709,N_20327,N_21521);
nand U26710 (N_26710,N_20875,N_24908);
nor U26711 (N_26711,N_24072,N_20343);
nand U26712 (N_26712,N_21113,N_20158);
and U26713 (N_26713,N_23133,N_21645);
and U26714 (N_26714,N_20028,N_21730);
xnor U26715 (N_26715,N_21834,N_24551);
nor U26716 (N_26716,N_24532,N_21304);
or U26717 (N_26717,N_22191,N_22144);
nand U26718 (N_26718,N_21718,N_20631);
and U26719 (N_26719,N_20741,N_24337);
nor U26720 (N_26720,N_20676,N_23776);
and U26721 (N_26721,N_23344,N_21471);
nand U26722 (N_26722,N_24950,N_20941);
xnor U26723 (N_26723,N_20493,N_20281);
and U26724 (N_26724,N_21608,N_21241);
nand U26725 (N_26725,N_22057,N_20024);
xnor U26726 (N_26726,N_23732,N_21216);
and U26727 (N_26727,N_23221,N_21446);
xnor U26728 (N_26728,N_20862,N_20218);
or U26729 (N_26729,N_22613,N_20730);
nand U26730 (N_26730,N_20014,N_21681);
xnor U26731 (N_26731,N_20849,N_23793);
nor U26732 (N_26732,N_23626,N_23568);
or U26733 (N_26733,N_20090,N_23942);
or U26734 (N_26734,N_21691,N_23979);
and U26735 (N_26735,N_23758,N_23263);
and U26736 (N_26736,N_24805,N_20517);
nand U26737 (N_26737,N_20813,N_24940);
and U26738 (N_26738,N_22269,N_24410);
and U26739 (N_26739,N_24783,N_21612);
or U26740 (N_26740,N_20886,N_20415);
or U26741 (N_26741,N_22169,N_24155);
nor U26742 (N_26742,N_23409,N_24034);
or U26743 (N_26743,N_20953,N_22290);
xor U26744 (N_26744,N_21983,N_21624);
nor U26745 (N_26745,N_23645,N_20232);
nor U26746 (N_26746,N_20392,N_20257);
or U26747 (N_26747,N_22888,N_22807);
and U26748 (N_26748,N_21972,N_22922);
and U26749 (N_26749,N_21654,N_20374);
nand U26750 (N_26750,N_23703,N_24292);
nor U26751 (N_26751,N_23139,N_24585);
nor U26752 (N_26752,N_22296,N_22450);
nor U26753 (N_26753,N_23865,N_22370);
nor U26754 (N_26754,N_21391,N_22526);
nor U26755 (N_26755,N_22143,N_20766);
nor U26756 (N_26756,N_22920,N_24504);
or U26757 (N_26757,N_24243,N_21778);
or U26758 (N_26758,N_22115,N_20377);
nor U26759 (N_26759,N_20277,N_21016);
nand U26760 (N_26760,N_24027,N_24101);
and U26761 (N_26761,N_22003,N_20925);
and U26762 (N_26762,N_21813,N_23955);
or U26763 (N_26763,N_20701,N_21662);
nor U26764 (N_26764,N_21630,N_21480);
nor U26765 (N_26765,N_21955,N_21999);
nand U26766 (N_26766,N_24169,N_20192);
and U26767 (N_26767,N_21268,N_21427);
xnor U26768 (N_26768,N_22600,N_22628);
or U26769 (N_26769,N_22993,N_22873);
nand U26770 (N_26770,N_24333,N_24889);
or U26771 (N_26771,N_22853,N_23861);
or U26772 (N_26772,N_22728,N_24137);
nand U26773 (N_26773,N_21814,N_21795);
nand U26774 (N_26774,N_21133,N_24171);
or U26775 (N_26775,N_24937,N_22185);
nor U26776 (N_26776,N_24959,N_21235);
nor U26777 (N_26777,N_21771,N_22145);
nand U26778 (N_26778,N_20038,N_24491);
nand U26779 (N_26779,N_20782,N_21847);
nor U26780 (N_26780,N_20812,N_20753);
nand U26781 (N_26781,N_23016,N_24515);
nand U26782 (N_26782,N_23968,N_23219);
or U26783 (N_26783,N_22996,N_21807);
nand U26784 (N_26784,N_21741,N_20403);
and U26785 (N_26785,N_23731,N_24737);
xor U26786 (N_26786,N_23320,N_23168);
nand U26787 (N_26787,N_23116,N_22997);
nand U26788 (N_26788,N_22736,N_21750);
nand U26789 (N_26789,N_21517,N_21281);
nor U26790 (N_26790,N_24494,N_20721);
nor U26791 (N_26791,N_21651,N_22297);
or U26792 (N_26792,N_24429,N_24339);
xnor U26793 (N_26793,N_24217,N_24145);
nor U26794 (N_26794,N_20747,N_24363);
or U26795 (N_26795,N_20834,N_22013);
and U26796 (N_26796,N_20589,N_22985);
nand U26797 (N_26797,N_21794,N_23433);
nand U26798 (N_26798,N_23608,N_24338);
nor U26799 (N_26799,N_21757,N_20370);
or U26800 (N_26800,N_23346,N_22709);
nor U26801 (N_26801,N_20672,N_22104);
xnor U26802 (N_26802,N_22797,N_23296);
xor U26803 (N_26803,N_24481,N_21511);
or U26804 (N_26804,N_23165,N_20670);
or U26805 (N_26805,N_24431,N_24124);
nor U26806 (N_26806,N_20560,N_22170);
nor U26807 (N_26807,N_20046,N_24699);
or U26808 (N_26808,N_20486,N_23450);
or U26809 (N_26809,N_22301,N_22930);
or U26810 (N_26810,N_21042,N_22380);
and U26811 (N_26811,N_23428,N_24383);
nand U26812 (N_26812,N_20845,N_20224);
or U26813 (N_26813,N_24404,N_24018);
or U26814 (N_26814,N_22146,N_22482);
or U26815 (N_26815,N_21171,N_20719);
nor U26816 (N_26816,N_23691,N_21790);
and U26817 (N_26817,N_22866,N_22642);
nand U26818 (N_26818,N_20206,N_22158);
or U26819 (N_26819,N_23189,N_22329);
nor U26820 (N_26820,N_22152,N_23742);
nor U26821 (N_26821,N_24553,N_23306);
nor U26822 (N_26822,N_24151,N_24806);
xor U26823 (N_26823,N_23167,N_21793);
nand U26824 (N_26824,N_20268,N_20939);
or U26825 (N_26825,N_22014,N_23830);
xnor U26826 (N_26826,N_23077,N_22172);
or U26827 (N_26827,N_24126,N_21332);
or U26828 (N_26828,N_24403,N_20496);
and U26829 (N_26829,N_21818,N_22556);
nand U26830 (N_26830,N_22259,N_21448);
nand U26831 (N_26831,N_22307,N_23369);
or U26832 (N_26832,N_21110,N_24242);
nand U26833 (N_26833,N_21349,N_22157);
nor U26834 (N_26834,N_22137,N_24825);
and U26835 (N_26835,N_21779,N_21611);
and U26836 (N_26836,N_21846,N_23112);
nor U26837 (N_26837,N_24894,N_22884);
and U26838 (N_26838,N_21881,N_24814);
or U26839 (N_26839,N_23484,N_22887);
and U26840 (N_26840,N_20070,N_24947);
nor U26841 (N_26841,N_20048,N_21688);
nand U26842 (N_26842,N_22743,N_24903);
nor U26843 (N_26843,N_22001,N_20740);
nand U26844 (N_26844,N_23642,N_20966);
xor U26845 (N_26845,N_23079,N_24918);
nand U26846 (N_26846,N_22006,N_22012);
xor U26847 (N_26847,N_24772,N_20292);
nand U26848 (N_26848,N_20274,N_23665);
xor U26849 (N_26849,N_22464,N_21909);
nand U26850 (N_26850,N_22579,N_24030);
nor U26851 (N_26851,N_22294,N_24720);
and U26852 (N_26852,N_20581,N_20981);
nand U26853 (N_26853,N_21689,N_24051);
nor U26854 (N_26854,N_24819,N_23046);
xnor U26855 (N_26855,N_20639,N_23384);
and U26856 (N_26856,N_20597,N_23361);
nor U26857 (N_26857,N_24134,N_24742);
and U26858 (N_26858,N_20360,N_20045);
or U26859 (N_26859,N_23293,N_23154);
and U26860 (N_26860,N_20256,N_22917);
and U26861 (N_26861,N_20437,N_22795);
and U26862 (N_26862,N_20654,N_24616);
or U26863 (N_26863,N_24732,N_21927);
and U26864 (N_26864,N_24965,N_20656);
and U26865 (N_26865,N_23938,N_24992);
nor U26866 (N_26866,N_22026,N_22769);
or U26867 (N_26867,N_21346,N_21956);
or U26868 (N_26868,N_20570,N_23677);
or U26869 (N_26869,N_24117,N_24301);
or U26870 (N_26870,N_22594,N_24595);
nor U26871 (N_26871,N_20804,N_23174);
and U26872 (N_26872,N_23410,N_21641);
nor U26873 (N_26873,N_20151,N_21143);
or U26874 (N_26874,N_20134,N_24344);
nand U26875 (N_26875,N_23924,N_21441);
nor U26876 (N_26876,N_20203,N_23455);
or U26877 (N_26877,N_20395,N_24626);
or U26878 (N_26878,N_23453,N_24530);
nor U26879 (N_26879,N_20209,N_20818);
or U26880 (N_26880,N_21934,N_22788);
nor U26881 (N_26881,N_20836,N_21649);
or U26882 (N_26882,N_24975,N_20142);
and U26883 (N_26883,N_23596,N_22225);
or U26884 (N_26884,N_20917,N_24434);
nand U26885 (N_26885,N_24215,N_20638);
xor U26886 (N_26886,N_23720,N_22761);
nand U26887 (N_26887,N_23949,N_20944);
and U26888 (N_26888,N_22190,N_24020);
nand U26889 (N_26889,N_21785,N_24946);
nand U26890 (N_26890,N_22867,N_20214);
or U26891 (N_26891,N_24261,N_23443);
or U26892 (N_26892,N_24076,N_21449);
and U26893 (N_26893,N_24765,N_23417);
nand U26894 (N_26894,N_20258,N_20050);
or U26895 (N_26895,N_22872,N_21980);
nand U26896 (N_26896,N_21288,N_20752);
xor U26897 (N_26897,N_20592,N_21048);
and U26898 (N_26898,N_21176,N_21603);
and U26899 (N_26899,N_23027,N_23085);
or U26900 (N_26900,N_20266,N_21120);
or U26901 (N_26901,N_20191,N_20608);
nand U26902 (N_26902,N_20351,N_22987);
nand U26903 (N_26903,N_21605,N_20239);
nand U26904 (N_26904,N_22784,N_24275);
xnor U26905 (N_26905,N_22314,N_22094);
or U26906 (N_26906,N_21535,N_21289);
or U26907 (N_26907,N_20062,N_21209);
and U26908 (N_26908,N_23481,N_21040);
xor U26909 (N_26909,N_22916,N_20715);
nor U26910 (N_26910,N_24025,N_23717);
nand U26911 (N_26911,N_22539,N_24461);
or U26912 (N_26912,N_20950,N_20373);
nor U26913 (N_26913,N_23692,N_23759);
or U26914 (N_26914,N_24357,N_20168);
nand U26915 (N_26915,N_24449,N_22661);
or U26916 (N_26916,N_24622,N_21024);
nand U26917 (N_26917,N_22223,N_22473);
and U26918 (N_26918,N_24778,N_21033);
nand U26919 (N_26919,N_23636,N_23483);
nand U26920 (N_26920,N_21188,N_22586);
or U26921 (N_26921,N_22700,N_22264);
nor U26922 (N_26922,N_22299,N_24949);
or U26923 (N_26923,N_23752,N_21714);
nand U26924 (N_26924,N_24663,N_23230);
xor U26925 (N_26925,N_24794,N_20585);
and U26926 (N_26926,N_24568,N_22626);
nor U26927 (N_26927,N_23215,N_21214);
or U26928 (N_26928,N_22184,N_23774);
or U26929 (N_26929,N_23543,N_21244);
or U26930 (N_26930,N_21297,N_21149);
nor U26931 (N_26931,N_22516,N_23198);
and U26932 (N_26932,N_20765,N_23640);
xor U26933 (N_26933,N_23735,N_22066);
or U26934 (N_26934,N_24516,N_24871);
or U26935 (N_26935,N_21924,N_23616);
nor U26936 (N_26936,N_24141,N_21240);
or U26937 (N_26937,N_21031,N_21686);
and U26938 (N_26938,N_24358,N_21661);
nor U26939 (N_26939,N_20504,N_20596);
or U26940 (N_26940,N_20475,N_21468);
or U26941 (N_26941,N_23997,N_20922);
or U26942 (N_26942,N_23438,N_20751);
or U26943 (N_26943,N_24428,N_21230);
nand U26944 (N_26944,N_24956,N_20613);
xnor U26945 (N_26945,N_24007,N_22933);
nor U26946 (N_26946,N_24973,N_24901);
nor U26947 (N_26947,N_22150,N_24964);
and U26948 (N_26948,N_21308,N_21402);
nand U26949 (N_26949,N_20905,N_23008);
or U26950 (N_26950,N_22836,N_24278);
nor U26951 (N_26951,N_20336,N_20755);
nand U26952 (N_26952,N_23406,N_20131);
nand U26953 (N_26953,N_22491,N_20668);
and U26954 (N_26954,N_24993,N_22948);
xor U26955 (N_26955,N_24666,N_20627);
xnor U26956 (N_26956,N_22277,N_22272);
nor U26957 (N_26957,N_22982,N_21499);
xor U26958 (N_26958,N_24890,N_21735);
nand U26959 (N_26959,N_22772,N_21319);
or U26960 (N_26960,N_24895,N_23822);
nor U26961 (N_26961,N_21533,N_21462);
nand U26962 (N_26962,N_22581,N_21509);
xor U26963 (N_26963,N_22039,N_23396);
nor U26964 (N_26964,N_21992,N_20969);
or U26965 (N_26965,N_24596,N_21524);
nor U26966 (N_26966,N_20890,N_20573);
or U26967 (N_26967,N_23148,N_22474);
nand U26968 (N_26968,N_21892,N_24280);
nor U26969 (N_26969,N_23319,N_22608);
nor U26970 (N_26970,N_20178,N_24621);
nand U26971 (N_26971,N_22413,N_24861);
nor U26972 (N_26972,N_22513,N_20894);
nor U26973 (N_26973,N_20318,N_22365);
or U26974 (N_26974,N_23505,N_23132);
nor U26975 (N_26975,N_23281,N_21456);
and U26976 (N_26976,N_22207,N_21895);
and U26977 (N_26977,N_20664,N_20405);
or U26978 (N_26978,N_21072,N_20651);
or U26979 (N_26979,N_24715,N_23606);
and U26980 (N_26980,N_23975,N_22360);
and U26981 (N_26981,N_22326,N_21022);
nor U26982 (N_26982,N_20509,N_20919);
nand U26983 (N_26983,N_21324,N_23397);
nor U26984 (N_26984,N_22965,N_23823);
nand U26985 (N_26985,N_20960,N_22070);
or U26986 (N_26986,N_20215,N_20564);
or U26987 (N_26987,N_20025,N_20216);
or U26988 (N_26988,N_20459,N_20623);
or U26989 (N_26989,N_21569,N_23037);
nand U26990 (N_26990,N_23377,N_20750);
nand U26991 (N_26991,N_22864,N_20421);
nor U26992 (N_26992,N_20068,N_24967);
and U26993 (N_26993,N_22705,N_24756);
nand U26994 (N_26994,N_24767,N_23471);
nand U26995 (N_26995,N_21141,N_20699);
nor U26996 (N_26996,N_24477,N_23818);
xnor U26997 (N_26997,N_21773,N_21335);
or U26998 (N_26998,N_24412,N_24259);
nand U26999 (N_26999,N_22915,N_22842);
xor U27000 (N_27000,N_22693,N_22760);
or U27001 (N_27001,N_20826,N_21482);
or U27002 (N_27002,N_22903,N_20982);
or U27003 (N_27003,N_24249,N_22535);
nand U27004 (N_27004,N_24133,N_21958);
nand U27005 (N_27005,N_23447,N_20522);
nor U27006 (N_27006,N_23810,N_21518);
or U27007 (N_27007,N_24866,N_20149);
or U27008 (N_27008,N_23816,N_24207);
and U27009 (N_27009,N_21931,N_24601);
and U27010 (N_27010,N_21780,N_22854);
nor U27011 (N_27011,N_23261,N_20043);
nand U27012 (N_27012,N_23010,N_24365);
nor U27013 (N_27013,N_24157,N_24549);
or U27014 (N_27014,N_21144,N_21726);
or U27015 (N_27015,N_20467,N_22636);
and U27016 (N_27016,N_22395,N_21763);
nor U27017 (N_27017,N_20283,N_20788);
and U27018 (N_27018,N_20641,N_20285);
nand U27019 (N_27019,N_21330,N_24368);
or U27020 (N_27020,N_22374,N_22830);
nand U27021 (N_27021,N_20357,N_23277);
nor U27022 (N_27022,N_23894,N_21516);
or U27023 (N_27023,N_22203,N_22949);
or U27024 (N_27024,N_21487,N_21781);
nor U27025 (N_27025,N_20123,N_24227);
nand U27026 (N_27026,N_22868,N_21694);
nor U27027 (N_27027,N_22634,N_20240);
or U27028 (N_27028,N_24598,N_21413);
xnor U27029 (N_27029,N_23950,N_20237);
and U27030 (N_27030,N_23967,N_20430);
nor U27031 (N_27031,N_23971,N_21271);
xor U27032 (N_27032,N_23812,N_22718);
and U27033 (N_27033,N_24328,N_22656);
nor U27034 (N_27034,N_21326,N_23585);
nand U27035 (N_27035,N_22263,N_20418);
nor U27036 (N_27036,N_22133,N_23715);
and U27037 (N_27037,N_21723,N_23520);
nor U27038 (N_27038,N_21267,N_22757);
or U27039 (N_27039,N_24351,N_20829);
or U27040 (N_27040,N_22334,N_23350);
nor U27041 (N_27041,N_22444,N_23755);
or U27042 (N_27042,N_24972,N_20527);
nand U27043 (N_27043,N_21995,N_24528);
nor U27044 (N_27044,N_24455,N_24068);
nand U27045 (N_27045,N_23917,N_21030);
xor U27046 (N_27046,N_22007,N_23094);
xor U27047 (N_27047,N_21668,N_24865);
nand U27048 (N_27048,N_20790,N_21960);
xnor U27049 (N_27049,N_20663,N_24356);
nor U27050 (N_27050,N_24103,N_24716);
nor U27051 (N_27051,N_21810,N_20401);
nor U27052 (N_27052,N_22341,N_21760);
and U27053 (N_27053,N_22273,N_21392);
nor U27054 (N_27054,N_22908,N_21969);
nor U27055 (N_27055,N_20003,N_21452);
nand U27056 (N_27056,N_22831,N_24486);
nand U27057 (N_27057,N_24525,N_21725);
nor U27058 (N_27058,N_21414,N_24256);
nor U27059 (N_27059,N_23140,N_20630);
nand U27060 (N_27060,N_23236,N_20060);
and U27061 (N_27061,N_20021,N_22874);
nor U27062 (N_27062,N_24951,N_21886);
nand U27063 (N_27063,N_21582,N_23421);
nor U27064 (N_27064,N_23704,N_20735);
nand U27065 (N_27065,N_20212,N_20899);
or U27066 (N_27066,N_20231,N_21942);
or U27067 (N_27067,N_21910,N_24073);
nand U27068 (N_27068,N_23427,N_24042);
or U27069 (N_27069,N_20163,N_22044);
nand U27070 (N_27070,N_22663,N_21357);
nand U27071 (N_27071,N_20514,N_22318);
nor U27072 (N_27072,N_24738,N_23931);
nor U27073 (N_27073,N_21200,N_23152);
nand U27074 (N_27074,N_24883,N_21600);
or U27075 (N_27075,N_20652,N_24163);
or U27076 (N_27076,N_20743,N_20346);
nand U27077 (N_27077,N_23262,N_22737);
and U27078 (N_27078,N_23945,N_24593);
nand U27079 (N_27079,N_22968,N_20749);
and U27080 (N_27080,N_20990,N_23242);
or U27081 (N_27081,N_24841,N_21967);
xnor U27082 (N_27082,N_22182,N_23052);
or U27083 (N_27083,N_24802,N_24629);
nand U27084 (N_27084,N_24402,N_20126);
nor U27085 (N_27085,N_22179,N_21183);
and U27086 (N_27086,N_23625,N_23126);
xnor U27087 (N_27087,N_24647,N_23473);
nand U27088 (N_27088,N_21618,N_22702);
xor U27089 (N_27089,N_21198,N_24268);
nor U27090 (N_27090,N_22779,N_23913);
and U27091 (N_27091,N_23284,N_21028);
nand U27092 (N_27092,N_21243,N_22485);
and U27093 (N_27093,N_24285,N_23074);
nand U27094 (N_27094,N_24506,N_21667);
or U27095 (N_27095,N_22604,N_21893);
nand U27096 (N_27096,N_21463,N_20175);
or U27097 (N_27097,N_20432,N_24200);
xor U27098 (N_27098,N_24676,N_22940);
nor U27099 (N_27099,N_22232,N_20709);
nand U27100 (N_27100,N_22235,N_23170);
nand U27101 (N_27101,N_24065,N_24835);
and U27102 (N_27102,N_24748,N_22148);
nand U27103 (N_27103,N_21708,N_23962);
and U27104 (N_27104,N_20872,N_20267);
or U27105 (N_27105,N_23222,N_20483);
nor U27106 (N_27106,N_23749,N_22383);
nor U27107 (N_27107,N_24533,N_21161);
nor U27108 (N_27108,N_24726,N_24334);
and U27109 (N_27109,N_21593,N_22192);
nand U27110 (N_27110,N_20238,N_24922);
xnor U27111 (N_27111,N_22470,N_23051);
nand U27112 (N_27112,N_20692,N_20659);
and U27113 (N_27113,N_21372,N_22838);
and U27114 (N_27114,N_22879,N_20102);
nor U27115 (N_27115,N_24482,N_24033);
nand U27116 (N_27116,N_23661,N_23662);
nand U27117 (N_27117,N_20551,N_23401);
and U27118 (N_27118,N_23352,N_20604);
or U27119 (N_27119,N_23773,N_22767);
nand U27120 (N_27120,N_22181,N_24093);
and U27121 (N_27121,N_22362,N_24816);
nor U27122 (N_27122,N_22020,N_23444);
nand U27123 (N_27123,N_23233,N_24370);
and U27124 (N_27124,N_21864,N_23034);
or U27125 (N_27125,N_23835,N_21836);
xor U27126 (N_27126,N_20155,N_22097);
nand U27127 (N_27127,N_21932,N_22588);
or U27128 (N_27128,N_21278,N_24837);
and U27129 (N_27129,N_23061,N_23745);
nand U27130 (N_27130,N_22074,N_21493);
and U27131 (N_27131,N_24246,N_24267);
and U27132 (N_27132,N_22319,N_20666);
or U27133 (N_27133,N_24603,N_24649);
nor U27134 (N_27134,N_23791,N_23476);
nand U27135 (N_27135,N_22451,N_23398);
and U27136 (N_27136,N_20888,N_23600);
xor U27137 (N_27137,N_22856,N_23995);
and U27138 (N_27138,N_22699,N_22462);
nor U27139 (N_27139,N_22536,N_24492);
or U27140 (N_27140,N_24572,N_20042);
and U27141 (N_27141,N_20914,N_23131);
nand U27142 (N_27142,N_20466,N_20555);
nand U27143 (N_27143,N_24577,N_21158);
nor U27144 (N_27144,N_20803,N_24997);
xor U27145 (N_27145,N_23743,N_24473);
or U27146 (N_27146,N_22951,N_22589);
and U27147 (N_27147,N_24878,N_24202);
or U27148 (N_27148,N_23501,N_22823);
or U27149 (N_27149,N_20093,N_23880);
nand U27150 (N_27150,N_23275,N_20665);
xor U27151 (N_27151,N_22347,N_24054);
nor U27152 (N_27152,N_24452,N_21440);
and U27153 (N_27153,N_21015,N_22745);
xnor U27154 (N_27154,N_24274,N_24283);
nand U27155 (N_27155,N_21921,N_24945);
xnor U27156 (N_27156,N_20468,N_21513);
nand U27157 (N_27157,N_21765,N_20780);
nor U27158 (N_27158,N_23193,N_23781);
xnor U27159 (N_27159,N_22389,N_24136);
xor U27160 (N_27160,N_22194,N_21466);
and U27161 (N_27161,N_24592,N_22610);
nor U27162 (N_27162,N_22827,N_23495);
or U27163 (N_27163,N_20511,N_20096);
or U27164 (N_27164,N_24801,N_20725);
nor U27165 (N_27165,N_24982,N_22358);
nand U27166 (N_27166,N_24005,N_22564);
nand U27167 (N_27167,N_20887,N_21566);
and U27168 (N_27168,N_23766,N_24681);
and U27169 (N_27169,N_22017,N_20446);
and U27170 (N_27170,N_22238,N_23531);
or U27171 (N_27171,N_22153,N_20411);
and U27172 (N_27172,N_22202,N_20768);
nand U27173 (N_27173,N_24454,N_21623);
nor U27174 (N_27174,N_21546,N_24178);
xor U27175 (N_27175,N_24463,N_23399);
nand U27176 (N_27176,N_24859,N_23489);
or U27177 (N_27177,N_20678,N_23844);
nand U27178 (N_27178,N_24730,N_24798);
nor U27179 (N_27179,N_22387,N_21687);
nand U27180 (N_27180,N_21388,N_22287);
or U27181 (N_27181,N_23878,N_23297);
nand U27182 (N_27182,N_20547,N_24498);
nor U27183 (N_27183,N_24564,N_24838);
and U27184 (N_27184,N_20722,N_22453);
or U27185 (N_27185,N_24990,N_23134);
xnor U27186 (N_27186,N_23701,N_21266);
nand U27187 (N_27187,N_23794,N_22381);
xnor U27188 (N_27188,N_20690,N_20771);
nand U27189 (N_27189,N_24142,N_20423);
and U27190 (N_27190,N_21428,N_23680);
or U27191 (N_27191,N_22255,N_24341);
nand U27192 (N_27192,N_20213,N_21453);
nand U27193 (N_27193,N_23939,N_22412);
nand U27194 (N_27194,N_24690,N_23683);
and U27195 (N_27195,N_22675,N_23615);
or U27196 (N_27196,N_23590,N_24499);
and U27197 (N_27197,N_23641,N_24307);
nand U27198 (N_27198,N_23845,N_21628);
nor U27199 (N_27199,N_24432,N_20473);
and U27200 (N_27200,N_21806,N_20222);
nor U27201 (N_27201,N_24270,N_21021);
or U27202 (N_27202,N_23194,N_20078);
xor U27203 (N_27203,N_21504,N_22615);
xor U27204 (N_27204,N_20325,N_21656);
or U27205 (N_27205,N_23881,N_21409);
nor U27206 (N_27206,N_21682,N_20634);
and U27207 (N_27207,N_24083,N_24953);
nor U27208 (N_27208,N_20390,N_23235);
xnor U27209 (N_27209,N_24727,N_24192);
and U27210 (N_27210,N_21747,N_24369);
or U27211 (N_27211,N_23765,N_22424);
and U27212 (N_27212,N_22641,N_23904);
nor U27213 (N_27213,N_20311,N_23007);
and U27214 (N_27214,N_24689,N_21702);
xor U27215 (N_27215,N_23025,N_23842);
and U27216 (N_27216,N_20018,N_20892);
or U27217 (N_27217,N_22687,N_23448);
and U27218 (N_27218,N_20383,N_22392);
nor U27219 (N_27219,N_21870,N_24749);
nor U27220 (N_27220,N_24168,N_21145);
nor U27221 (N_27221,N_22073,N_22083);
and U27222 (N_27222,N_21047,N_22376);
nand U27223 (N_27223,N_20734,N_22160);
and U27224 (N_27224,N_21635,N_20200);
nor U27225 (N_27225,N_21657,N_24558);
and U27226 (N_27226,N_20786,N_24747);
or U27227 (N_27227,N_23200,N_24875);
nor U27228 (N_27228,N_23903,N_23855);
or U27229 (N_27229,N_20745,N_23504);
and U27230 (N_27230,N_20433,N_23647);
xor U27231 (N_27231,N_21073,N_20230);
and U27232 (N_27232,N_24208,N_21862);
and U27233 (N_27233,N_21058,N_23525);
xnor U27234 (N_27234,N_21423,N_22557);
and U27235 (N_27235,N_22457,N_23090);
or U27236 (N_27236,N_24539,N_20756);
and U27237 (N_27237,N_24047,N_22753);
nand U27238 (N_27238,N_24401,N_23621);
nor U27239 (N_27239,N_24210,N_24507);
xor U27240 (N_27240,N_20516,N_23593);
and U27241 (N_27241,N_23669,N_21782);
nand U27242 (N_27242,N_20356,N_23843);
nand U27243 (N_27243,N_21381,N_20649);
xnor U27244 (N_27244,N_20091,N_21665);
nor U27245 (N_27245,N_20489,N_21553);
or U27246 (N_27246,N_23166,N_24750);
nor U27247 (N_27247,N_24424,N_22563);
and U27248 (N_27248,N_22870,N_24332);
xnor U27249 (N_27249,N_21091,N_20031);
nand U27250 (N_27250,N_23273,N_20998);
and U27251 (N_27251,N_21238,N_23291);
nor U27252 (N_27252,N_22877,N_22311);
nor U27253 (N_27253,N_23778,N_23321);
and U27254 (N_27254,N_23502,N_24470);
xnor U27255 (N_27255,N_21601,N_21859);
or U27256 (N_27256,N_21234,N_23014);
xor U27257 (N_27257,N_20855,N_22715);
or U27258 (N_27258,N_23514,N_24130);
nand U27259 (N_27259,N_23208,N_24012);
and U27260 (N_27260,N_20225,N_22609);
and U27261 (N_27261,N_20779,N_23539);
or U27262 (N_27262,N_24581,N_23449);
xor U27263 (N_27263,N_22256,N_22665);
and U27264 (N_27264,N_21828,N_22509);
nor U27265 (N_27265,N_23748,N_24927);
nand U27266 (N_27266,N_20548,N_20964);
nor U27267 (N_27267,N_21364,N_24849);
or U27268 (N_27268,N_22028,N_22072);
or U27269 (N_27269,N_22977,N_23620);
or U27270 (N_27270,N_23841,N_21706);
nand U27271 (N_27271,N_23379,N_24196);
nand U27272 (N_27272,N_23186,N_22931);
and U27273 (N_27273,N_20180,N_20805);
and U27274 (N_27274,N_21250,N_22205);
nand U27275 (N_27275,N_20138,N_24996);
xor U27276 (N_27276,N_23225,N_23343);
nand U27277 (N_27277,N_20566,N_22566);
nor U27278 (N_27278,N_23875,N_21871);
nor U27279 (N_27279,N_21699,N_22386);
nand U27280 (N_27280,N_22484,N_21592);
nand U27281 (N_27281,N_21123,N_24880);
xnor U27282 (N_27282,N_21786,N_22912);
nor U27283 (N_27283,N_23195,N_22630);
nand U27284 (N_27284,N_23936,N_22657);
nor U27285 (N_27285,N_21896,N_23987);
nand U27286 (N_27286,N_23724,N_20602);
or U27287 (N_27287,N_24830,N_20333);
nand U27288 (N_27288,N_24531,N_21537);
nand U27289 (N_27289,N_22010,N_24744);
nand U27290 (N_27290,N_24708,N_24388);
or U27291 (N_27291,N_23300,N_22472);
and U27292 (N_27292,N_21823,N_22507);
nor U27293 (N_27293,N_21160,N_20041);
nand U27294 (N_27294,N_24988,N_22407);
nor U27295 (N_27295,N_24850,N_22197);
xor U27296 (N_27296,N_20593,N_23712);
and U27297 (N_27297,N_24056,N_20454);
nor U27298 (N_27298,N_21210,N_20706);
nand U27299 (N_27299,N_23442,N_23462);
or U27300 (N_27300,N_23533,N_24803);
nand U27301 (N_27301,N_24050,N_21784);
xnor U27302 (N_27302,N_23466,N_20359);
nor U27303 (N_27303,N_23160,N_22422);
or U27304 (N_27304,N_21918,N_22892);
nand U27305 (N_27305,N_21619,N_20746);
nand U27306 (N_27306,N_24911,N_20885);
or U27307 (N_27307,N_23940,N_22180);
and U27308 (N_27308,N_23073,N_20601);
or U27309 (N_27309,N_20609,N_22623);
or U27310 (N_27310,N_23754,N_24542);
nor U27311 (N_27311,N_21320,N_22828);
and U27312 (N_27312,N_22755,N_20315);
and U27313 (N_27313,N_21914,N_24590);
nand U27314 (N_27314,N_21606,N_23963);
and U27315 (N_27315,N_22427,N_21940);
and U27316 (N_27316,N_20296,N_23264);
nor U27317 (N_27317,N_21721,N_21722);
xor U27318 (N_27318,N_20099,N_23294);
and U27319 (N_27319,N_21949,N_23738);
nor U27320 (N_27320,N_24476,N_24248);
and U27321 (N_27321,N_24493,N_21616);
nand U27322 (N_27322,N_20059,N_21526);
nand U27323 (N_27323,N_21112,N_24684);
nor U27324 (N_27324,N_20528,N_22835);
or U27325 (N_27325,N_20498,N_20376);
nand U27326 (N_27326,N_20576,N_22603);
and U27327 (N_27327,N_20518,N_24416);
nor U27328 (N_27328,N_23578,N_21742);
or U27329 (N_27329,N_23736,N_24781);
and U27330 (N_27330,N_20136,N_21432);
and U27331 (N_27331,N_24746,N_21137);
or U27332 (N_27332,N_23605,N_21928);
or U27333 (N_27333,N_23391,N_20868);
and U27334 (N_27334,N_22284,N_24381);
nor U27335 (N_27335,N_20455,N_23478);
xor U27336 (N_27336,N_21419,N_23093);
xnor U27337 (N_27337,N_20162,N_21563);
nor U27338 (N_27338,N_23459,N_23107);
or U27339 (N_27339,N_24851,N_21777);
and U27340 (N_27340,N_20260,N_24704);
and U27341 (N_27341,N_24265,N_22310);
or U27342 (N_27342,N_24605,N_20724);
nand U27343 (N_27343,N_23825,N_23347);
nand U27344 (N_27344,N_24125,N_20714);
nor U27345 (N_27345,N_24627,N_22214);
and U27346 (N_27346,N_21902,N_21256);
nor U27347 (N_27347,N_23465,N_23001);
nor U27348 (N_27348,N_21279,N_20895);
and U27349 (N_27349,N_24273,N_23322);
nand U27350 (N_27350,N_20148,N_20345);
nand U27351 (N_27351,N_21731,N_23191);
nor U27352 (N_27352,N_24004,N_24660);
or U27353 (N_27353,N_23457,N_22896);
and U27354 (N_27354,N_24177,N_23467);
nand U27355 (N_27355,N_24448,N_23560);
or U27356 (N_27356,N_23299,N_23408);
nor U27357 (N_27357,N_21536,N_23959);
and U27358 (N_27358,N_23974,N_23985);
and U27359 (N_27359,N_24574,N_22865);
nand U27360 (N_27360,N_22363,N_23451);
nand U27361 (N_27361,N_22217,N_20056);
xor U27362 (N_27362,N_21585,N_22243);
nor U27363 (N_27363,N_22905,N_20940);
or U27364 (N_27364,N_23162,N_20363);
nor U27365 (N_27365,N_22883,N_20806);
and U27366 (N_27366,N_21008,N_23631);
and U27367 (N_27367,N_23799,N_23413);
and U27368 (N_27368,N_20220,N_22369);
nor U27369 (N_27369,N_20962,N_24028);
or U27370 (N_27370,N_23729,N_21303);
nand U27371 (N_27371,N_24438,N_21574);
and U27372 (N_27372,N_21229,N_20047);
nor U27373 (N_27373,N_20490,N_22653);
xnor U27374 (N_27374,N_20986,N_21339);
xor U27375 (N_27375,N_22984,N_24423);
nor U27376 (N_27376,N_20603,N_22680);
nand U27377 (N_27377,N_20864,N_24314);
nor U27378 (N_27378,N_23800,N_21065);
nand U27379 (N_27379,N_21650,N_22911);
nor U27380 (N_27380,N_22349,N_20770);
and U27381 (N_27381,N_23201,N_24843);
or U27382 (N_27382,N_20989,N_24562);
nand U27383 (N_27383,N_24786,N_23113);
nor U27384 (N_27384,N_23206,N_24035);
nor U27385 (N_27385,N_24500,N_23289);
nand U27386 (N_27386,N_24910,N_21277);
nand U27387 (N_27387,N_20406,N_22575);
and U27388 (N_27388,N_21937,N_21634);
and U27389 (N_27389,N_21581,N_20367);
nand U27390 (N_27390,N_21187,N_22839);
xor U27391 (N_27391,N_21294,N_21799);
nand U27392 (N_27392,N_23231,N_20271);
nor U27393 (N_27393,N_20520,N_20007);
and U27394 (N_27394,N_22910,N_20412);
nor U27395 (N_27395,N_20900,N_23877);
and U27396 (N_27396,N_21182,N_24496);
or U27397 (N_27397,N_21822,N_22056);
or U27398 (N_27398,N_21911,N_21491);
and U27399 (N_27399,N_21443,N_24271);
nor U27400 (N_27400,N_24294,N_23345);
nor U27401 (N_27401,N_22644,N_24282);
xnor U27402 (N_27402,N_21620,N_20754);
xor U27403 (N_27403,N_21107,N_21027);
or U27404 (N_27404,N_22652,N_24606);
nand U27405 (N_27405,N_22956,N_20229);
nor U27406 (N_27406,N_20394,N_21561);
and U27407 (N_27407,N_23340,N_23243);
or U27408 (N_27408,N_20893,N_24239);
and U27409 (N_27409,N_20183,N_21373);
nor U27410 (N_27410,N_21374,N_20869);
nor U27411 (N_27411,N_22818,N_20884);
and U27412 (N_27412,N_23482,N_20275);
or U27413 (N_27413,N_23175,N_24006);
and U27414 (N_27414,N_23095,N_20228);
xor U27415 (N_27415,N_20844,N_22859);
or U27416 (N_27416,N_22021,N_20094);
and U27417 (N_27417,N_20362,N_20515);
nor U27418 (N_27418,N_24743,N_20793);
nor U27419 (N_27419,N_24241,N_21839);
nor U27420 (N_27420,N_22500,N_20160);
xnor U27421 (N_27421,N_20710,N_24105);
nor U27422 (N_27422,N_22138,N_20295);
or U27423 (N_27423,N_20563,N_20671);
nor U27424 (N_27424,N_20852,N_23866);
or U27425 (N_27425,N_22976,N_21676);
and U27426 (N_27426,N_23083,N_24775);
and U27427 (N_27427,N_23178,N_24673);
and U27428 (N_27428,N_20321,N_22342);
nor U27429 (N_27429,N_21247,N_24159);
and U27430 (N_27430,N_23002,N_21677);
nand U27431 (N_27431,N_22498,N_22139);
nor U27432 (N_27432,N_22402,N_23580);
nand U27433 (N_27433,N_23120,N_21664);
nor U27434 (N_27434,N_21348,N_20847);
or U27435 (N_27435,N_24391,N_20121);
and U27436 (N_27436,N_23562,N_21287);
and U27437 (N_27437,N_21745,N_22244);
nand U27438 (N_27438,N_22645,N_21317);
or U27439 (N_27439,N_21206,N_20934);
nor U27440 (N_27440,N_23588,N_21792);
nand U27441 (N_27441,N_24272,N_24643);
or U27442 (N_27442,N_21135,N_21527);
and U27443 (N_27443,N_22546,N_22251);
or U27444 (N_27444,N_23854,N_24118);
and U27445 (N_27445,N_21081,N_23441);
xnor U27446 (N_27446,N_23644,N_23375);
xor U27447 (N_27447,N_23711,N_21390);
nand U27448 (N_27448,N_20251,N_24002);
and U27449 (N_27449,N_22561,N_20488);
and U27450 (N_27450,N_22654,N_22822);
nor U27451 (N_27451,N_20442,N_21312);
and U27452 (N_27452,N_21376,N_22096);
and U27453 (N_27453,N_20626,N_23920);
nand U27454 (N_27454,N_20642,N_21090);
or U27455 (N_27455,N_23953,N_24784);
or U27456 (N_27456,N_22611,N_21396);
or U27457 (N_27457,N_24662,N_21154);
nand U27458 (N_27458,N_24869,N_22724);
and U27459 (N_27459,N_20600,N_23576);
xor U27460 (N_27460,N_23053,N_22084);
and U27461 (N_27461,N_24672,N_23461);
nand U27462 (N_27462,N_21729,N_22721);
nand U27463 (N_27463,N_22088,N_20643);
xnor U27464 (N_27464,N_23911,N_20058);
or U27465 (N_27465,N_22960,N_23362);
or U27466 (N_27466,N_22315,N_24782);
or U27467 (N_27467,N_20928,N_24284);
and U27468 (N_27468,N_24597,N_22990);
and U27469 (N_27469,N_22861,N_20537);
nor U27470 (N_27470,N_23657,N_20955);
nand U27471 (N_27471,N_24711,N_21867);
nor U27472 (N_27472,N_20208,N_22275);
and U27473 (N_27473,N_21262,N_20250);
nor U27474 (N_27474,N_20856,N_22885);
and U27475 (N_27475,N_23925,N_23675);
and U27476 (N_27476,N_21146,N_21855);
or U27477 (N_27477,N_24773,N_23414);
nand U27478 (N_27478,N_22367,N_20308);
and U27479 (N_27479,N_20871,N_22002);
or U27480 (N_27480,N_22248,N_24394);
and U27481 (N_27481,N_21484,N_21222);
xor U27482 (N_27482,N_22489,N_22167);
nor U27483 (N_27483,N_21363,N_23811);
or U27484 (N_27484,N_24921,N_20431);
nand U27485 (N_27485,N_20340,N_23147);
nor U27486 (N_27486,N_23055,N_24810);
nand U27487 (N_27487,N_20908,N_24924);
nor U27488 (N_27488,N_20103,N_20736);
and U27489 (N_27489,N_21237,N_24713);
or U27490 (N_27490,N_21602,N_24335);
nor U27491 (N_27491,N_23064,N_20085);
or U27492 (N_27492,N_22245,N_20541);
nor U27493 (N_27493,N_22970,N_21752);
and U27494 (N_27494,N_24442,N_21377);
nand U27495 (N_27495,N_23579,N_22189);
or U27496 (N_27496,N_21469,N_20506);
or U27497 (N_27497,N_20127,N_20009);
nor U27498 (N_27498,N_24497,N_22775);
nand U27499 (N_27499,N_21979,N_22418);
nand U27500 (N_27500,N_23437,N_21731);
nand U27501 (N_27501,N_20388,N_24922);
or U27502 (N_27502,N_22940,N_23633);
or U27503 (N_27503,N_20647,N_21852);
nand U27504 (N_27504,N_24787,N_23121);
or U27505 (N_27505,N_23852,N_22617);
or U27506 (N_27506,N_23236,N_20902);
or U27507 (N_27507,N_20280,N_21475);
and U27508 (N_27508,N_24919,N_23815);
xnor U27509 (N_27509,N_21329,N_24958);
or U27510 (N_27510,N_24484,N_21505);
and U27511 (N_27511,N_22361,N_20679);
or U27512 (N_27512,N_22732,N_24437);
nand U27513 (N_27513,N_20376,N_24312);
xor U27514 (N_27514,N_21936,N_24199);
and U27515 (N_27515,N_21339,N_21926);
nor U27516 (N_27516,N_20050,N_20237);
or U27517 (N_27517,N_22277,N_24525);
nor U27518 (N_27518,N_21481,N_24688);
nor U27519 (N_27519,N_22612,N_24675);
or U27520 (N_27520,N_21764,N_21827);
nand U27521 (N_27521,N_23471,N_20410);
nand U27522 (N_27522,N_23382,N_21595);
nand U27523 (N_27523,N_22338,N_24722);
nor U27524 (N_27524,N_22859,N_21806);
nand U27525 (N_27525,N_23215,N_21105);
or U27526 (N_27526,N_23017,N_24578);
nor U27527 (N_27527,N_23395,N_23291);
and U27528 (N_27528,N_20662,N_21100);
nand U27529 (N_27529,N_23751,N_21749);
and U27530 (N_27530,N_24898,N_23509);
xnor U27531 (N_27531,N_20583,N_23481);
or U27532 (N_27532,N_22569,N_21340);
and U27533 (N_27533,N_23535,N_24481);
and U27534 (N_27534,N_22129,N_24371);
nand U27535 (N_27535,N_24655,N_20606);
or U27536 (N_27536,N_23129,N_20400);
xor U27537 (N_27537,N_23305,N_24712);
nand U27538 (N_27538,N_24178,N_24954);
nor U27539 (N_27539,N_22818,N_24125);
nor U27540 (N_27540,N_24296,N_23765);
nand U27541 (N_27541,N_24897,N_20113);
nand U27542 (N_27542,N_23823,N_24318);
nand U27543 (N_27543,N_23390,N_20377);
nor U27544 (N_27544,N_20637,N_22519);
xor U27545 (N_27545,N_24326,N_21106);
or U27546 (N_27546,N_21958,N_23609);
and U27547 (N_27547,N_21518,N_22697);
nand U27548 (N_27548,N_20163,N_24527);
nand U27549 (N_27549,N_23322,N_22661);
nor U27550 (N_27550,N_21062,N_21443);
nor U27551 (N_27551,N_21075,N_24108);
or U27552 (N_27552,N_20615,N_20273);
and U27553 (N_27553,N_23622,N_24204);
nor U27554 (N_27554,N_24348,N_20581);
nand U27555 (N_27555,N_24895,N_21531);
and U27556 (N_27556,N_21772,N_20696);
or U27557 (N_27557,N_24429,N_22110);
nand U27558 (N_27558,N_21048,N_23049);
or U27559 (N_27559,N_23994,N_21414);
nor U27560 (N_27560,N_21034,N_21011);
or U27561 (N_27561,N_20109,N_24571);
or U27562 (N_27562,N_23375,N_24223);
xor U27563 (N_27563,N_22807,N_20443);
and U27564 (N_27564,N_23767,N_23978);
and U27565 (N_27565,N_22567,N_20644);
nor U27566 (N_27566,N_22485,N_21552);
and U27567 (N_27567,N_22078,N_22301);
nand U27568 (N_27568,N_21316,N_24016);
or U27569 (N_27569,N_20711,N_21331);
and U27570 (N_27570,N_23784,N_23417);
and U27571 (N_27571,N_22745,N_21754);
nand U27572 (N_27572,N_21545,N_22009);
and U27573 (N_27573,N_22277,N_20729);
xnor U27574 (N_27574,N_24459,N_21100);
and U27575 (N_27575,N_24728,N_23517);
and U27576 (N_27576,N_21714,N_21137);
nor U27577 (N_27577,N_21070,N_24001);
or U27578 (N_27578,N_22912,N_23369);
or U27579 (N_27579,N_21251,N_22955);
and U27580 (N_27580,N_23630,N_24743);
nand U27581 (N_27581,N_24777,N_24219);
and U27582 (N_27582,N_20269,N_21007);
xnor U27583 (N_27583,N_20132,N_24159);
and U27584 (N_27584,N_22331,N_23398);
nand U27585 (N_27585,N_21702,N_22301);
nor U27586 (N_27586,N_22506,N_21046);
nand U27587 (N_27587,N_24848,N_24244);
nand U27588 (N_27588,N_21998,N_22650);
nand U27589 (N_27589,N_21354,N_24885);
xnor U27590 (N_27590,N_21568,N_22983);
nor U27591 (N_27591,N_21089,N_23997);
nand U27592 (N_27592,N_20057,N_22031);
or U27593 (N_27593,N_20480,N_23598);
nand U27594 (N_27594,N_23765,N_24939);
and U27595 (N_27595,N_20634,N_22364);
nand U27596 (N_27596,N_23410,N_24958);
and U27597 (N_27597,N_22121,N_22211);
nor U27598 (N_27598,N_21189,N_21183);
nand U27599 (N_27599,N_23753,N_23513);
or U27600 (N_27600,N_23120,N_20247);
nand U27601 (N_27601,N_21849,N_20402);
or U27602 (N_27602,N_23505,N_20475);
or U27603 (N_27603,N_24916,N_24268);
nand U27604 (N_27604,N_22213,N_23040);
nor U27605 (N_27605,N_20604,N_20635);
or U27606 (N_27606,N_24539,N_23055);
nor U27607 (N_27607,N_21142,N_23473);
or U27608 (N_27608,N_22526,N_22062);
or U27609 (N_27609,N_24565,N_24645);
or U27610 (N_27610,N_23615,N_20144);
and U27611 (N_27611,N_22096,N_23919);
nand U27612 (N_27612,N_23315,N_23986);
and U27613 (N_27613,N_21011,N_20367);
or U27614 (N_27614,N_20673,N_20942);
or U27615 (N_27615,N_21768,N_22957);
nor U27616 (N_27616,N_23911,N_22199);
nand U27617 (N_27617,N_20855,N_23038);
or U27618 (N_27618,N_24444,N_20656);
nand U27619 (N_27619,N_20818,N_22050);
nand U27620 (N_27620,N_21564,N_24853);
and U27621 (N_27621,N_24724,N_20396);
or U27622 (N_27622,N_20370,N_21764);
or U27623 (N_27623,N_23095,N_20753);
or U27624 (N_27624,N_20447,N_22701);
nand U27625 (N_27625,N_23032,N_22143);
and U27626 (N_27626,N_21740,N_20404);
nand U27627 (N_27627,N_21226,N_20098);
or U27628 (N_27628,N_23384,N_20851);
xnor U27629 (N_27629,N_23410,N_21607);
nor U27630 (N_27630,N_23091,N_23555);
nor U27631 (N_27631,N_21102,N_23309);
and U27632 (N_27632,N_24838,N_22433);
nand U27633 (N_27633,N_21444,N_23325);
xor U27634 (N_27634,N_20337,N_24226);
and U27635 (N_27635,N_23812,N_20589);
nor U27636 (N_27636,N_20521,N_21619);
nand U27637 (N_27637,N_23076,N_21404);
or U27638 (N_27638,N_21475,N_22858);
nand U27639 (N_27639,N_22077,N_20217);
nand U27640 (N_27640,N_22593,N_23174);
xnor U27641 (N_27641,N_21995,N_23590);
or U27642 (N_27642,N_22428,N_24654);
or U27643 (N_27643,N_23677,N_24409);
nor U27644 (N_27644,N_21304,N_21843);
nand U27645 (N_27645,N_20336,N_21734);
xnor U27646 (N_27646,N_20380,N_21488);
nand U27647 (N_27647,N_21435,N_22138);
nand U27648 (N_27648,N_20474,N_20109);
or U27649 (N_27649,N_20188,N_22494);
or U27650 (N_27650,N_23756,N_22885);
nand U27651 (N_27651,N_22657,N_22410);
and U27652 (N_27652,N_20227,N_20105);
or U27653 (N_27653,N_21907,N_23924);
or U27654 (N_27654,N_20143,N_20852);
xor U27655 (N_27655,N_21244,N_21092);
or U27656 (N_27656,N_22696,N_24786);
nor U27657 (N_27657,N_22120,N_23708);
or U27658 (N_27658,N_23583,N_23574);
nand U27659 (N_27659,N_20869,N_23227);
or U27660 (N_27660,N_21825,N_22118);
or U27661 (N_27661,N_23718,N_24854);
or U27662 (N_27662,N_20317,N_21620);
and U27663 (N_27663,N_21090,N_20694);
nor U27664 (N_27664,N_20475,N_23628);
nand U27665 (N_27665,N_23362,N_22825);
nand U27666 (N_27666,N_22332,N_22429);
xor U27667 (N_27667,N_20406,N_21401);
or U27668 (N_27668,N_24268,N_21167);
or U27669 (N_27669,N_23641,N_21153);
nor U27670 (N_27670,N_23732,N_24564);
nand U27671 (N_27671,N_23146,N_23858);
nand U27672 (N_27672,N_24543,N_24414);
or U27673 (N_27673,N_24653,N_21699);
or U27674 (N_27674,N_23293,N_21482);
nand U27675 (N_27675,N_23832,N_24631);
or U27676 (N_27676,N_21080,N_21333);
nor U27677 (N_27677,N_23772,N_20417);
nand U27678 (N_27678,N_20416,N_20694);
nor U27679 (N_27679,N_22350,N_20250);
nor U27680 (N_27680,N_24370,N_24488);
and U27681 (N_27681,N_24697,N_23253);
or U27682 (N_27682,N_24921,N_23950);
nor U27683 (N_27683,N_20709,N_20348);
nand U27684 (N_27684,N_24452,N_20555);
and U27685 (N_27685,N_23945,N_20984);
nor U27686 (N_27686,N_24548,N_23373);
xor U27687 (N_27687,N_23562,N_23742);
nor U27688 (N_27688,N_23432,N_23738);
nor U27689 (N_27689,N_23662,N_23048);
nand U27690 (N_27690,N_20832,N_21285);
and U27691 (N_27691,N_20632,N_24241);
and U27692 (N_27692,N_22514,N_21466);
or U27693 (N_27693,N_20317,N_21252);
or U27694 (N_27694,N_23682,N_23821);
or U27695 (N_27695,N_21461,N_23228);
nand U27696 (N_27696,N_23929,N_21365);
nand U27697 (N_27697,N_24245,N_20587);
and U27698 (N_27698,N_22243,N_22080);
nand U27699 (N_27699,N_21836,N_23256);
xor U27700 (N_27700,N_20223,N_20810);
nor U27701 (N_27701,N_22310,N_22529);
nand U27702 (N_27702,N_21296,N_21878);
and U27703 (N_27703,N_20870,N_22394);
or U27704 (N_27704,N_20320,N_22130);
nand U27705 (N_27705,N_22740,N_20234);
nand U27706 (N_27706,N_21053,N_23916);
or U27707 (N_27707,N_24899,N_21384);
and U27708 (N_27708,N_23899,N_22039);
or U27709 (N_27709,N_24425,N_22351);
or U27710 (N_27710,N_23993,N_23404);
nand U27711 (N_27711,N_23655,N_20090);
xnor U27712 (N_27712,N_23648,N_21000);
nand U27713 (N_27713,N_22610,N_22489);
nand U27714 (N_27714,N_23422,N_23826);
xnor U27715 (N_27715,N_20938,N_24075);
nand U27716 (N_27716,N_20612,N_22845);
nand U27717 (N_27717,N_20925,N_24370);
xnor U27718 (N_27718,N_22891,N_20712);
nand U27719 (N_27719,N_20147,N_22891);
nor U27720 (N_27720,N_20522,N_20672);
nand U27721 (N_27721,N_20424,N_22768);
or U27722 (N_27722,N_22755,N_24311);
nand U27723 (N_27723,N_21126,N_20964);
or U27724 (N_27724,N_23639,N_23479);
nor U27725 (N_27725,N_22299,N_23412);
nand U27726 (N_27726,N_24208,N_20546);
or U27727 (N_27727,N_22928,N_21233);
or U27728 (N_27728,N_23829,N_21192);
nand U27729 (N_27729,N_24038,N_22054);
nand U27730 (N_27730,N_23824,N_23552);
or U27731 (N_27731,N_20241,N_23530);
or U27732 (N_27732,N_23478,N_22337);
nor U27733 (N_27733,N_23003,N_24800);
nor U27734 (N_27734,N_22198,N_23518);
nor U27735 (N_27735,N_20543,N_24002);
and U27736 (N_27736,N_21228,N_24205);
and U27737 (N_27737,N_20347,N_21167);
xnor U27738 (N_27738,N_20965,N_22084);
and U27739 (N_27739,N_22120,N_20073);
or U27740 (N_27740,N_20535,N_20906);
nor U27741 (N_27741,N_20338,N_22447);
nand U27742 (N_27742,N_20572,N_24330);
nor U27743 (N_27743,N_22141,N_22275);
nand U27744 (N_27744,N_20507,N_20259);
or U27745 (N_27745,N_24825,N_24216);
and U27746 (N_27746,N_20322,N_22267);
or U27747 (N_27747,N_24208,N_21909);
nor U27748 (N_27748,N_21825,N_22360);
nor U27749 (N_27749,N_22928,N_20348);
nand U27750 (N_27750,N_21854,N_20791);
nand U27751 (N_27751,N_23570,N_23144);
nor U27752 (N_27752,N_24279,N_23557);
or U27753 (N_27753,N_21964,N_20720);
and U27754 (N_27754,N_24018,N_20089);
nor U27755 (N_27755,N_23291,N_24601);
and U27756 (N_27756,N_24322,N_23476);
or U27757 (N_27757,N_22267,N_22584);
and U27758 (N_27758,N_24644,N_22250);
or U27759 (N_27759,N_23724,N_24102);
or U27760 (N_27760,N_24129,N_22843);
or U27761 (N_27761,N_20438,N_20235);
or U27762 (N_27762,N_22765,N_21573);
and U27763 (N_27763,N_21322,N_21630);
xor U27764 (N_27764,N_20420,N_21943);
nand U27765 (N_27765,N_22875,N_20792);
or U27766 (N_27766,N_22955,N_24628);
or U27767 (N_27767,N_22042,N_21952);
and U27768 (N_27768,N_20612,N_22294);
or U27769 (N_27769,N_20220,N_21847);
nand U27770 (N_27770,N_23337,N_21986);
or U27771 (N_27771,N_22895,N_23732);
or U27772 (N_27772,N_23630,N_21504);
nand U27773 (N_27773,N_23857,N_21473);
nand U27774 (N_27774,N_24702,N_24503);
nor U27775 (N_27775,N_20453,N_20307);
nor U27776 (N_27776,N_23354,N_22366);
nor U27777 (N_27777,N_22360,N_23186);
and U27778 (N_27778,N_22648,N_20906);
and U27779 (N_27779,N_20071,N_23854);
and U27780 (N_27780,N_24633,N_22080);
nor U27781 (N_27781,N_23553,N_21390);
nor U27782 (N_27782,N_23904,N_21754);
nand U27783 (N_27783,N_22232,N_23151);
or U27784 (N_27784,N_20688,N_22893);
and U27785 (N_27785,N_21755,N_22795);
or U27786 (N_27786,N_22792,N_22347);
nand U27787 (N_27787,N_21803,N_21628);
nand U27788 (N_27788,N_22324,N_20744);
nor U27789 (N_27789,N_20894,N_23216);
or U27790 (N_27790,N_21699,N_20288);
or U27791 (N_27791,N_21534,N_22102);
or U27792 (N_27792,N_20102,N_24393);
xnor U27793 (N_27793,N_24591,N_23481);
or U27794 (N_27794,N_21064,N_22079);
and U27795 (N_27795,N_24523,N_24941);
nand U27796 (N_27796,N_23534,N_21009);
nor U27797 (N_27797,N_23377,N_22523);
or U27798 (N_27798,N_20301,N_24670);
or U27799 (N_27799,N_23370,N_22440);
or U27800 (N_27800,N_21293,N_24627);
xnor U27801 (N_27801,N_21202,N_24378);
nor U27802 (N_27802,N_20459,N_20743);
and U27803 (N_27803,N_21870,N_20810);
nand U27804 (N_27804,N_22701,N_23539);
nand U27805 (N_27805,N_21397,N_23732);
nor U27806 (N_27806,N_21222,N_23863);
and U27807 (N_27807,N_20014,N_21914);
nand U27808 (N_27808,N_20177,N_23787);
or U27809 (N_27809,N_20740,N_21417);
nand U27810 (N_27810,N_22459,N_21574);
nand U27811 (N_27811,N_22182,N_23648);
nor U27812 (N_27812,N_23783,N_22926);
nand U27813 (N_27813,N_22817,N_23896);
or U27814 (N_27814,N_21484,N_24260);
or U27815 (N_27815,N_21571,N_21367);
nor U27816 (N_27816,N_24974,N_21962);
xnor U27817 (N_27817,N_22254,N_22568);
or U27818 (N_27818,N_24656,N_23400);
and U27819 (N_27819,N_24560,N_23529);
and U27820 (N_27820,N_22962,N_23163);
nand U27821 (N_27821,N_23183,N_20825);
xor U27822 (N_27822,N_23800,N_22923);
and U27823 (N_27823,N_21526,N_24660);
nand U27824 (N_27824,N_23738,N_22628);
xor U27825 (N_27825,N_21979,N_22863);
and U27826 (N_27826,N_24450,N_24639);
and U27827 (N_27827,N_22938,N_24133);
nor U27828 (N_27828,N_22377,N_20360);
and U27829 (N_27829,N_21918,N_24380);
and U27830 (N_27830,N_22520,N_22562);
and U27831 (N_27831,N_24296,N_24135);
and U27832 (N_27832,N_22371,N_24612);
and U27833 (N_27833,N_24953,N_24623);
nand U27834 (N_27834,N_20471,N_24637);
nor U27835 (N_27835,N_20716,N_20091);
and U27836 (N_27836,N_20497,N_21000);
or U27837 (N_27837,N_22758,N_24112);
nor U27838 (N_27838,N_24539,N_24261);
and U27839 (N_27839,N_24403,N_22475);
or U27840 (N_27840,N_22956,N_22553);
or U27841 (N_27841,N_24706,N_20566);
or U27842 (N_27842,N_22296,N_23653);
or U27843 (N_27843,N_22741,N_22868);
xnor U27844 (N_27844,N_22324,N_21152);
nor U27845 (N_27845,N_20156,N_24385);
nor U27846 (N_27846,N_23083,N_20819);
or U27847 (N_27847,N_23324,N_24280);
and U27848 (N_27848,N_20919,N_21055);
or U27849 (N_27849,N_21710,N_21317);
nand U27850 (N_27850,N_24863,N_24559);
nand U27851 (N_27851,N_22139,N_20315);
and U27852 (N_27852,N_21348,N_23701);
and U27853 (N_27853,N_20967,N_21233);
or U27854 (N_27854,N_23357,N_22426);
nor U27855 (N_27855,N_23289,N_21836);
and U27856 (N_27856,N_21412,N_21125);
nor U27857 (N_27857,N_20125,N_20682);
and U27858 (N_27858,N_22785,N_23504);
and U27859 (N_27859,N_24064,N_21852);
nand U27860 (N_27860,N_21130,N_22613);
nand U27861 (N_27861,N_20325,N_21366);
nor U27862 (N_27862,N_21175,N_22107);
and U27863 (N_27863,N_23982,N_22574);
nor U27864 (N_27864,N_20753,N_23808);
xnor U27865 (N_27865,N_21473,N_20602);
or U27866 (N_27866,N_22787,N_23029);
nand U27867 (N_27867,N_20036,N_23264);
nor U27868 (N_27868,N_21001,N_24364);
or U27869 (N_27869,N_23653,N_21622);
xor U27870 (N_27870,N_24814,N_22936);
and U27871 (N_27871,N_22942,N_24247);
and U27872 (N_27872,N_20279,N_21704);
nor U27873 (N_27873,N_21517,N_22716);
and U27874 (N_27874,N_23797,N_22485);
nor U27875 (N_27875,N_21425,N_24121);
nand U27876 (N_27876,N_22847,N_20014);
nor U27877 (N_27877,N_20730,N_20306);
nor U27878 (N_27878,N_24281,N_23535);
and U27879 (N_27879,N_24491,N_23510);
and U27880 (N_27880,N_20372,N_21115);
and U27881 (N_27881,N_21020,N_20192);
and U27882 (N_27882,N_20105,N_23226);
nand U27883 (N_27883,N_22047,N_24873);
or U27884 (N_27884,N_23877,N_23102);
and U27885 (N_27885,N_20033,N_21172);
or U27886 (N_27886,N_24862,N_22803);
nor U27887 (N_27887,N_24289,N_23271);
or U27888 (N_27888,N_22399,N_22443);
or U27889 (N_27889,N_24937,N_20175);
nand U27890 (N_27890,N_22426,N_24594);
nor U27891 (N_27891,N_20470,N_22997);
nor U27892 (N_27892,N_23626,N_20445);
xor U27893 (N_27893,N_21106,N_20265);
nand U27894 (N_27894,N_22947,N_21435);
xnor U27895 (N_27895,N_24954,N_20763);
xnor U27896 (N_27896,N_24597,N_22481);
nor U27897 (N_27897,N_24645,N_24180);
or U27898 (N_27898,N_21069,N_20193);
or U27899 (N_27899,N_22696,N_21962);
nor U27900 (N_27900,N_24661,N_21687);
or U27901 (N_27901,N_20981,N_22622);
xor U27902 (N_27902,N_24993,N_22075);
or U27903 (N_27903,N_21237,N_24010);
and U27904 (N_27904,N_23262,N_23171);
and U27905 (N_27905,N_22980,N_21167);
xnor U27906 (N_27906,N_20307,N_21337);
nor U27907 (N_27907,N_23800,N_23615);
and U27908 (N_27908,N_22463,N_24410);
nor U27909 (N_27909,N_23886,N_23858);
nor U27910 (N_27910,N_20142,N_20069);
xor U27911 (N_27911,N_24458,N_23902);
or U27912 (N_27912,N_21045,N_23166);
nand U27913 (N_27913,N_21810,N_23833);
nand U27914 (N_27914,N_22582,N_20242);
nor U27915 (N_27915,N_20304,N_24351);
nand U27916 (N_27916,N_21397,N_20242);
and U27917 (N_27917,N_21181,N_23373);
xor U27918 (N_27918,N_22053,N_24331);
nor U27919 (N_27919,N_24703,N_22135);
or U27920 (N_27920,N_22389,N_22092);
nor U27921 (N_27921,N_22558,N_23768);
nor U27922 (N_27922,N_21723,N_20690);
or U27923 (N_27923,N_21651,N_20057);
nor U27924 (N_27924,N_21856,N_24123);
or U27925 (N_27925,N_21498,N_24145);
and U27926 (N_27926,N_23063,N_22691);
and U27927 (N_27927,N_22590,N_23204);
xnor U27928 (N_27928,N_21443,N_23927);
and U27929 (N_27929,N_23523,N_23563);
nand U27930 (N_27930,N_22665,N_23123);
nand U27931 (N_27931,N_24000,N_22596);
nand U27932 (N_27932,N_21560,N_24128);
and U27933 (N_27933,N_23519,N_24343);
xnor U27934 (N_27934,N_20453,N_20675);
and U27935 (N_27935,N_21881,N_22639);
and U27936 (N_27936,N_20120,N_21402);
nor U27937 (N_27937,N_21711,N_23071);
or U27938 (N_27938,N_20096,N_23993);
nor U27939 (N_27939,N_20562,N_20947);
or U27940 (N_27940,N_24071,N_21842);
nand U27941 (N_27941,N_23621,N_23018);
and U27942 (N_27942,N_20472,N_22382);
and U27943 (N_27943,N_22817,N_24355);
xor U27944 (N_27944,N_21634,N_21906);
nor U27945 (N_27945,N_24080,N_22078);
nor U27946 (N_27946,N_22171,N_21651);
and U27947 (N_27947,N_22913,N_21088);
nand U27948 (N_27948,N_20027,N_22671);
xor U27949 (N_27949,N_24709,N_20640);
nand U27950 (N_27950,N_22061,N_20890);
nor U27951 (N_27951,N_23234,N_22191);
and U27952 (N_27952,N_22967,N_22174);
and U27953 (N_27953,N_22286,N_20373);
or U27954 (N_27954,N_23140,N_24802);
xor U27955 (N_27955,N_21695,N_22867);
nand U27956 (N_27956,N_21238,N_21134);
nor U27957 (N_27957,N_23873,N_24333);
nand U27958 (N_27958,N_21300,N_23790);
nand U27959 (N_27959,N_23278,N_21149);
and U27960 (N_27960,N_23785,N_21397);
nor U27961 (N_27961,N_20855,N_23356);
or U27962 (N_27962,N_21522,N_23160);
nand U27963 (N_27963,N_23462,N_23805);
nand U27964 (N_27964,N_22999,N_24889);
and U27965 (N_27965,N_24751,N_21811);
nand U27966 (N_27966,N_22910,N_20489);
nor U27967 (N_27967,N_24699,N_20503);
nand U27968 (N_27968,N_24861,N_20447);
or U27969 (N_27969,N_20349,N_22392);
xor U27970 (N_27970,N_23028,N_22025);
or U27971 (N_27971,N_21004,N_23683);
nor U27972 (N_27972,N_20353,N_20560);
nand U27973 (N_27973,N_23476,N_22239);
nor U27974 (N_27974,N_20061,N_22781);
and U27975 (N_27975,N_24337,N_22751);
or U27976 (N_27976,N_22263,N_22293);
nand U27977 (N_27977,N_20056,N_21417);
xnor U27978 (N_27978,N_23999,N_22224);
and U27979 (N_27979,N_24468,N_20285);
and U27980 (N_27980,N_22708,N_23118);
or U27981 (N_27981,N_22541,N_21390);
nor U27982 (N_27982,N_22562,N_22832);
nand U27983 (N_27983,N_20080,N_24924);
nand U27984 (N_27984,N_23502,N_24029);
and U27985 (N_27985,N_21225,N_23270);
and U27986 (N_27986,N_24869,N_24624);
nand U27987 (N_27987,N_22736,N_24824);
nor U27988 (N_27988,N_20645,N_20122);
nor U27989 (N_27989,N_23668,N_23666);
or U27990 (N_27990,N_22193,N_23918);
or U27991 (N_27991,N_21698,N_23355);
or U27992 (N_27992,N_21145,N_20745);
nand U27993 (N_27993,N_22999,N_24599);
or U27994 (N_27994,N_21573,N_23479);
or U27995 (N_27995,N_20495,N_20697);
and U27996 (N_27996,N_23633,N_20882);
and U27997 (N_27997,N_21242,N_23522);
nand U27998 (N_27998,N_21754,N_23004);
xor U27999 (N_27999,N_22951,N_21986);
and U28000 (N_28000,N_22646,N_23647);
nand U28001 (N_28001,N_22009,N_23591);
and U28002 (N_28002,N_22170,N_22219);
nand U28003 (N_28003,N_24687,N_20208);
or U28004 (N_28004,N_20044,N_22240);
or U28005 (N_28005,N_23602,N_21927);
nor U28006 (N_28006,N_23748,N_24035);
xnor U28007 (N_28007,N_20150,N_23141);
and U28008 (N_28008,N_23917,N_23951);
and U28009 (N_28009,N_20611,N_24887);
nor U28010 (N_28010,N_22542,N_23110);
and U28011 (N_28011,N_24674,N_20858);
nor U28012 (N_28012,N_23415,N_21710);
nand U28013 (N_28013,N_20417,N_24798);
or U28014 (N_28014,N_24735,N_24251);
nand U28015 (N_28015,N_21999,N_23030);
nand U28016 (N_28016,N_20172,N_21138);
nand U28017 (N_28017,N_21315,N_24258);
and U28018 (N_28018,N_23898,N_23829);
nand U28019 (N_28019,N_24504,N_20792);
xnor U28020 (N_28020,N_20468,N_23685);
and U28021 (N_28021,N_20543,N_23116);
and U28022 (N_28022,N_22539,N_20697);
and U28023 (N_28023,N_20328,N_24923);
and U28024 (N_28024,N_23189,N_21844);
nand U28025 (N_28025,N_23605,N_22528);
nand U28026 (N_28026,N_21272,N_22961);
nor U28027 (N_28027,N_22475,N_24179);
nor U28028 (N_28028,N_24808,N_22607);
nor U28029 (N_28029,N_22086,N_24795);
nand U28030 (N_28030,N_21070,N_21640);
or U28031 (N_28031,N_22147,N_22890);
xnor U28032 (N_28032,N_20134,N_23167);
nor U28033 (N_28033,N_22433,N_21503);
nor U28034 (N_28034,N_23060,N_24200);
nand U28035 (N_28035,N_21954,N_22037);
or U28036 (N_28036,N_22057,N_24622);
and U28037 (N_28037,N_24056,N_22128);
nand U28038 (N_28038,N_21266,N_24962);
nor U28039 (N_28039,N_23840,N_24908);
nand U28040 (N_28040,N_22746,N_21991);
and U28041 (N_28041,N_23886,N_22303);
or U28042 (N_28042,N_23767,N_21409);
nand U28043 (N_28043,N_23312,N_20696);
or U28044 (N_28044,N_24879,N_23974);
nand U28045 (N_28045,N_22691,N_20867);
or U28046 (N_28046,N_20610,N_24039);
nor U28047 (N_28047,N_23045,N_22332);
or U28048 (N_28048,N_22246,N_22976);
and U28049 (N_28049,N_21343,N_22904);
xor U28050 (N_28050,N_20720,N_24351);
nor U28051 (N_28051,N_21881,N_22309);
or U28052 (N_28052,N_21574,N_20753);
nor U28053 (N_28053,N_22096,N_20428);
nand U28054 (N_28054,N_20768,N_21887);
nor U28055 (N_28055,N_21663,N_22795);
nand U28056 (N_28056,N_21509,N_24259);
and U28057 (N_28057,N_20794,N_21644);
or U28058 (N_28058,N_21289,N_20990);
or U28059 (N_28059,N_22919,N_23233);
or U28060 (N_28060,N_23827,N_23092);
and U28061 (N_28061,N_22861,N_23592);
or U28062 (N_28062,N_24226,N_22535);
nor U28063 (N_28063,N_20186,N_21606);
or U28064 (N_28064,N_20532,N_24685);
nand U28065 (N_28065,N_23405,N_22392);
or U28066 (N_28066,N_23505,N_23119);
xor U28067 (N_28067,N_20156,N_21483);
nor U28068 (N_28068,N_24873,N_22481);
xnor U28069 (N_28069,N_24811,N_23134);
nand U28070 (N_28070,N_23341,N_23517);
and U28071 (N_28071,N_22061,N_22686);
nand U28072 (N_28072,N_24564,N_20134);
nand U28073 (N_28073,N_21445,N_20682);
nor U28074 (N_28074,N_23666,N_22285);
nor U28075 (N_28075,N_24487,N_23380);
nand U28076 (N_28076,N_24372,N_20124);
and U28077 (N_28077,N_23273,N_21833);
and U28078 (N_28078,N_22393,N_21687);
xnor U28079 (N_28079,N_22314,N_22443);
or U28080 (N_28080,N_24260,N_24943);
and U28081 (N_28081,N_22105,N_22118);
or U28082 (N_28082,N_23609,N_20879);
nor U28083 (N_28083,N_24932,N_24186);
nor U28084 (N_28084,N_24101,N_21808);
nand U28085 (N_28085,N_23224,N_22269);
xnor U28086 (N_28086,N_21151,N_20800);
nand U28087 (N_28087,N_24613,N_21234);
nand U28088 (N_28088,N_22706,N_22219);
or U28089 (N_28089,N_24612,N_21033);
or U28090 (N_28090,N_21961,N_22854);
xor U28091 (N_28091,N_21317,N_21701);
and U28092 (N_28092,N_20407,N_24523);
nor U28093 (N_28093,N_20886,N_21536);
nor U28094 (N_28094,N_22057,N_20743);
nand U28095 (N_28095,N_20843,N_22845);
nor U28096 (N_28096,N_22391,N_24392);
or U28097 (N_28097,N_23354,N_22763);
xor U28098 (N_28098,N_22402,N_21858);
nor U28099 (N_28099,N_23853,N_21303);
nand U28100 (N_28100,N_23066,N_21601);
or U28101 (N_28101,N_22387,N_21040);
nand U28102 (N_28102,N_24071,N_20826);
or U28103 (N_28103,N_21999,N_21735);
xor U28104 (N_28104,N_24882,N_23540);
and U28105 (N_28105,N_24265,N_22434);
nor U28106 (N_28106,N_21803,N_24248);
nor U28107 (N_28107,N_20695,N_20503);
or U28108 (N_28108,N_24355,N_22235);
and U28109 (N_28109,N_22601,N_23331);
nand U28110 (N_28110,N_24848,N_21633);
and U28111 (N_28111,N_22603,N_21752);
and U28112 (N_28112,N_23709,N_21500);
or U28113 (N_28113,N_20765,N_23243);
xnor U28114 (N_28114,N_23436,N_24504);
or U28115 (N_28115,N_24485,N_23587);
or U28116 (N_28116,N_23680,N_21003);
nand U28117 (N_28117,N_23915,N_22135);
nor U28118 (N_28118,N_24187,N_21969);
or U28119 (N_28119,N_21163,N_21907);
and U28120 (N_28120,N_22502,N_22658);
nand U28121 (N_28121,N_22095,N_24308);
nand U28122 (N_28122,N_21168,N_23359);
or U28123 (N_28123,N_21146,N_20615);
nand U28124 (N_28124,N_21876,N_21709);
nand U28125 (N_28125,N_22078,N_23488);
nand U28126 (N_28126,N_23032,N_21378);
nand U28127 (N_28127,N_23942,N_21186);
nor U28128 (N_28128,N_24322,N_24708);
nor U28129 (N_28129,N_23713,N_24428);
and U28130 (N_28130,N_22435,N_24474);
nor U28131 (N_28131,N_22641,N_21439);
nor U28132 (N_28132,N_23839,N_24579);
nor U28133 (N_28133,N_23607,N_24905);
nand U28134 (N_28134,N_21397,N_24627);
nand U28135 (N_28135,N_24826,N_24547);
nor U28136 (N_28136,N_21052,N_24668);
nor U28137 (N_28137,N_23006,N_23927);
nor U28138 (N_28138,N_22180,N_22386);
nand U28139 (N_28139,N_24113,N_21094);
nor U28140 (N_28140,N_21456,N_22376);
nand U28141 (N_28141,N_20223,N_23381);
nor U28142 (N_28142,N_21644,N_20460);
or U28143 (N_28143,N_22669,N_20739);
xnor U28144 (N_28144,N_21480,N_21289);
and U28145 (N_28145,N_24306,N_24823);
xnor U28146 (N_28146,N_22725,N_23054);
nand U28147 (N_28147,N_24784,N_23426);
and U28148 (N_28148,N_22656,N_24765);
or U28149 (N_28149,N_23213,N_20538);
nand U28150 (N_28150,N_23114,N_22979);
nor U28151 (N_28151,N_21503,N_23957);
nor U28152 (N_28152,N_20270,N_24445);
nor U28153 (N_28153,N_21713,N_22113);
nand U28154 (N_28154,N_21330,N_22738);
nor U28155 (N_28155,N_21266,N_21038);
nand U28156 (N_28156,N_21692,N_21360);
and U28157 (N_28157,N_23657,N_21945);
xnor U28158 (N_28158,N_21796,N_23155);
or U28159 (N_28159,N_23649,N_24873);
and U28160 (N_28160,N_22954,N_24727);
nand U28161 (N_28161,N_23411,N_21374);
or U28162 (N_28162,N_24721,N_23387);
nand U28163 (N_28163,N_21856,N_20105);
nand U28164 (N_28164,N_22820,N_21650);
nand U28165 (N_28165,N_22837,N_21701);
nand U28166 (N_28166,N_23052,N_24303);
xor U28167 (N_28167,N_22540,N_20859);
xnor U28168 (N_28168,N_22170,N_20708);
and U28169 (N_28169,N_20271,N_24108);
nand U28170 (N_28170,N_21912,N_20747);
and U28171 (N_28171,N_24210,N_24687);
nor U28172 (N_28172,N_24658,N_21159);
nand U28173 (N_28173,N_21096,N_24954);
xor U28174 (N_28174,N_23634,N_20608);
and U28175 (N_28175,N_23180,N_22370);
xnor U28176 (N_28176,N_23953,N_20328);
or U28177 (N_28177,N_24813,N_22322);
or U28178 (N_28178,N_23816,N_24878);
and U28179 (N_28179,N_20386,N_23635);
nand U28180 (N_28180,N_21139,N_22015);
nor U28181 (N_28181,N_20296,N_22884);
nand U28182 (N_28182,N_21338,N_24105);
or U28183 (N_28183,N_23751,N_22403);
and U28184 (N_28184,N_20626,N_21322);
and U28185 (N_28185,N_22060,N_24223);
and U28186 (N_28186,N_20950,N_20665);
nor U28187 (N_28187,N_22182,N_21984);
nand U28188 (N_28188,N_23675,N_22345);
nor U28189 (N_28189,N_20578,N_22609);
nand U28190 (N_28190,N_21409,N_24086);
nor U28191 (N_28191,N_20689,N_23080);
nand U28192 (N_28192,N_24453,N_24671);
or U28193 (N_28193,N_21165,N_22304);
and U28194 (N_28194,N_23478,N_23136);
nand U28195 (N_28195,N_22423,N_24732);
or U28196 (N_28196,N_23429,N_20139);
or U28197 (N_28197,N_21581,N_22319);
nand U28198 (N_28198,N_21087,N_22295);
and U28199 (N_28199,N_22721,N_20775);
nand U28200 (N_28200,N_22286,N_21918);
and U28201 (N_28201,N_23255,N_22170);
nor U28202 (N_28202,N_21934,N_23322);
and U28203 (N_28203,N_21030,N_22853);
and U28204 (N_28204,N_24099,N_21034);
or U28205 (N_28205,N_21560,N_22065);
or U28206 (N_28206,N_22789,N_23745);
and U28207 (N_28207,N_21828,N_22210);
xor U28208 (N_28208,N_20802,N_20171);
xor U28209 (N_28209,N_21575,N_21868);
nor U28210 (N_28210,N_21063,N_23222);
or U28211 (N_28211,N_21488,N_20688);
and U28212 (N_28212,N_23054,N_24995);
nor U28213 (N_28213,N_22787,N_23506);
or U28214 (N_28214,N_22534,N_22718);
or U28215 (N_28215,N_20896,N_21722);
nand U28216 (N_28216,N_22211,N_22116);
or U28217 (N_28217,N_24421,N_21259);
nor U28218 (N_28218,N_22631,N_22414);
or U28219 (N_28219,N_24669,N_21697);
nor U28220 (N_28220,N_24057,N_21983);
nor U28221 (N_28221,N_21068,N_23637);
nor U28222 (N_28222,N_22309,N_24933);
or U28223 (N_28223,N_23722,N_20909);
and U28224 (N_28224,N_23253,N_24930);
or U28225 (N_28225,N_24528,N_24230);
nor U28226 (N_28226,N_22777,N_23998);
or U28227 (N_28227,N_23837,N_24215);
nand U28228 (N_28228,N_20761,N_21544);
and U28229 (N_28229,N_20834,N_20386);
nand U28230 (N_28230,N_21267,N_22616);
and U28231 (N_28231,N_23588,N_21493);
nor U28232 (N_28232,N_23770,N_20014);
and U28233 (N_28233,N_22771,N_24172);
and U28234 (N_28234,N_22460,N_20894);
nand U28235 (N_28235,N_24577,N_21366);
xor U28236 (N_28236,N_22321,N_23743);
xor U28237 (N_28237,N_23832,N_21967);
or U28238 (N_28238,N_21058,N_23637);
xor U28239 (N_28239,N_22172,N_24448);
and U28240 (N_28240,N_21916,N_24504);
nand U28241 (N_28241,N_20725,N_23817);
or U28242 (N_28242,N_22807,N_20934);
or U28243 (N_28243,N_21895,N_22252);
nor U28244 (N_28244,N_23581,N_24383);
and U28245 (N_28245,N_21622,N_21789);
nor U28246 (N_28246,N_24994,N_23078);
or U28247 (N_28247,N_22686,N_21700);
nand U28248 (N_28248,N_24810,N_20385);
and U28249 (N_28249,N_23239,N_23077);
nor U28250 (N_28250,N_23942,N_22986);
nand U28251 (N_28251,N_24245,N_24337);
or U28252 (N_28252,N_24420,N_20547);
nor U28253 (N_28253,N_21975,N_23937);
and U28254 (N_28254,N_24398,N_20472);
nand U28255 (N_28255,N_24040,N_21269);
nand U28256 (N_28256,N_21313,N_22896);
xor U28257 (N_28257,N_21827,N_24160);
and U28258 (N_28258,N_21564,N_23031);
nand U28259 (N_28259,N_24306,N_22208);
and U28260 (N_28260,N_23473,N_22827);
nor U28261 (N_28261,N_24541,N_24022);
and U28262 (N_28262,N_20570,N_20012);
nand U28263 (N_28263,N_23557,N_24350);
nor U28264 (N_28264,N_24849,N_20118);
and U28265 (N_28265,N_21780,N_22404);
nand U28266 (N_28266,N_24970,N_20590);
or U28267 (N_28267,N_20060,N_24168);
nand U28268 (N_28268,N_21248,N_24895);
nor U28269 (N_28269,N_21412,N_22590);
nand U28270 (N_28270,N_22856,N_21022);
nand U28271 (N_28271,N_22480,N_21901);
nand U28272 (N_28272,N_20367,N_23125);
and U28273 (N_28273,N_20575,N_22306);
nand U28274 (N_28274,N_20814,N_21297);
xor U28275 (N_28275,N_23848,N_24839);
nor U28276 (N_28276,N_22791,N_24696);
and U28277 (N_28277,N_22961,N_23681);
nor U28278 (N_28278,N_20909,N_23354);
or U28279 (N_28279,N_22861,N_24203);
and U28280 (N_28280,N_22720,N_23220);
xnor U28281 (N_28281,N_20777,N_21004);
and U28282 (N_28282,N_24200,N_21434);
nor U28283 (N_28283,N_22479,N_20158);
and U28284 (N_28284,N_20256,N_20306);
nand U28285 (N_28285,N_22043,N_24599);
and U28286 (N_28286,N_22959,N_20229);
nor U28287 (N_28287,N_21584,N_20738);
nand U28288 (N_28288,N_21807,N_24922);
or U28289 (N_28289,N_21043,N_20757);
nor U28290 (N_28290,N_20583,N_23081);
and U28291 (N_28291,N_23169,N_20737);
nand U28292 (N_28292,N_20727,N_24992);
xnor U28293 (N_28293,N_22973,N_24521);
nand U28294 (N_28294,N_24326,N_23448);
nand U28295 (N_28295,N_23321,N_23231);
nor U28296 (N_28296,N_21299,N_20241);
and U28297 (N_28297,N_20658,N_24864);
and U28298 (N_28298,N_21541,N_22265);
nor U28299 (N_28299,N_23382,N_21654);
nor U28300 (N_28300,N_22388,N_23083);
nor U28301 (N_28301,N_20815,N_23842);
or U28302 (N_28302,N_23952,N_22443);
xor U28303 (N_28303,N_22982,N_20966);
nand U28304 (N_28304,N_22893,N_21946);
xor U28305 (N_28305,N_22589,N_21031);
nor U28306 (N_28306,N_20709,N_22971);
and U28307 (N_28307,N_20476,N_24682);
and U28308 (N_28308,N_23306,N_22968);
or U28309 (N_28309,N_21969,N_22049);
xnor U28310 (N_28310,N_24979,N_23234);
nor U28311 (N_28311,N_22574,N_24493);
nand U28312 (N_28312,N_23866,N_23490);
nor U28313 (N_28313,N_23211,N_20347);
nand U28314 (N_28314,N_20750,N_21671);
or U28315 (N_28315,N_20935,N_24801);
nor U28316 (N_28316,N_22346,N_20935);
and U28317 (N_28317,N_24737,N_24014);
nand U28318 (N_28318,N_20145,N_24663);
nand U28319 (N_28319,N_23724,N_23065);
nand U28320 (N_28320,N_20035,N_22484);
nor U28321 (N_28321,N_21799,N_20917);
nor U28322 (N_28322,N_24198,N_23123);
or U28323 (N_28323,N_24995,N_24783);
xor U28324 (N_28324,N_22984,N_21716);
and U28325 (N_28325,N_21337,N_21931);
and U28326 (N_28326,N_20109,N_24742);
and U28327 (N_28327,N_21964,N_24202);
and U28328 (N_28328,N_24872,N_23166);
xnor U28329 (N_28329,N_20261,N_24341);
and U28330 (N_28330,N_21951,N_24039);
nand U28331 (N_28331,N_21745,N_22650);
and U28332 (N_28332,N_20055,N_23874);
or U28333 (N_28333,N_21892,N_23861);
and U28334 (N_28334,N_24727,N_22856);
nand U28335 (N_28335,N_24660,N_22978);
xnor U28336 (N_28336,N_20374,N_22914);
and U28337 (N_28337,N_21134,N_20956);
and U28338 (N_28338,N_22260,N_21461);
nand U28339 (N_28339,N_22445,N_23948);
or U28340 (N_28340,N_20572,N_20676);
nor U28341 (N_28341,N_24579,N_20190);
nor U28342 (N_28342,N_22299,N_21447);
nand U28343 (N_28343,N_21695,N_23271);
and U28344 (N_28344,N_20257,N_24194);
xor U28345 (N_28345,N_22305,N_22784);
nor U28346 (N_28346,N_23958,N_20396);
or U28347 (N_28347,N_23996,N_24246);
and U28348 (N_28348,N_23274,N_22190);
nor U28349 (N_28349,N_23488,N_21041);
nand U28350 (N_28350,N_23824,N_22422);
xor U28351 (N_28351,N_22975,N_22129);
nand U28352 (N_28352,N_22058,N_20911);
nor U28353 (N_28353,N_23357,N_21450);
or U28354 (N_28354,N_22144,N_23190);
nor U28355 (N_28355,N_24672,N_23360);
and U28356 (N_28356,N_24194,N_24284);
nor U28357 (N_28357,N_21479,N_24671);
or U28358 (N_28358,N_21205,N_23930);
and U28359 (N_28359,N_23960,N_23374);
and U28360 (N_28360,N_20767,N_24840);
nor U28361 (N_28361,N_23635,N_21939);
nand U28362 (N_28362,N_22190,N_23138);
or U28363 (N_28363,N_20710,N_23390);
or U28364 (N_28364,N_23548,N_20047);
and U28365 (N_28365,N_20632,N_21227);
and U28366 (N_28366,N_23203,N_22160);
or U28367 (N_28367,N_23183,N_24120);
nand U28368 (N_28368,N_24088,N_22446);
xor U28369 (N_28369,N_21630,N_22380);
and U28370 (N_28370,N_22703,N_20245);
xor U28371 (N_28371,N_23544,N_22769);
xnor U28372 (N_28372,N_24394,N_20261);
nand U28373 (N_28373,N_24139,N_22023);
or U28374 (N_28374,N_20265,N_21824);
nor U28375 (N_28375,N_22962,N_24984);
or U28376 (N_28376,N_22742,N_24474);
nor U28377 (N_28377,N_21452,N_20173);
or U28378 (N_28378,N_23581,N_20653);
nor U28379 (N_28379,N_21100,N_20233);
nand U28380 (N_28380,N_20018,N_22140);
xor U28381 (N_28381,N_21449,N_20279);
nand U28382 (N_28382,N_21495,N_23812);
nand U28383 (N_28383,N_24782,N_21085);
nor U28384 (N_28384,N_20411,N_23480);
nand U28385 (N_28385,N_23747,N_24233);
and U28386 (N_28386,N_20395,N_24917);
nand U28387 (N_28387,N_24850,N_21328);
xnor U28388 (N_28388,N_23345,N_20631);
xor U28389 (N_28389,N_23477,N_24263);
nor U28390 (N_28390,N_22413,N_24231);
and U28391 (N_28391,N_21491,N_20398);
nand U28392 (N_28392,N_21535,N_22173);
and U28393 (N_28393,N_24731,N_23112);
nand U28394 (N_28394,N_21260,N_23353);
xnor U28395 (N_28395,N_23543,N_24373);
and U28396 (N_28396,N_21989,N_20987);
or U28397 (N_28397,N_21205,N_21650);
or U28398 (N_28398,N_22522,N_24678);
xor U28399 (N_28399,N_20280,N_22246);
or U28400 (N_28400,N_22806,N_24802);
xor U28401 (N_28401,N_22875,N_20761);
nand U28402 (N_28402,N_20700,N_21224);
nor U28403 (N_28403,N_24887,N_23561);
nand U28404 (N_28404,N_23820,N_20460);
and U28405 (N_28405,N_23654,N_24913);
or U28406 (N_28406,N_21155,N_23831);
or U28407 (N_28407,N_23179,N_20926);
xnor U28408 (N_28408,N_20887,N_20364);
nor U28409 (N_28409,N_24907,N_23888);
and U28410 (N_28410,N_20560,N_21044);
nand U28411 (N_28411,N_23040,N_20076);
nor U28412 (N_28412,N_22078,N_21519);
and U28413 (N_28413,N_20211,N_20881);
or U28414 (N_28414,N_20292,N_20963);
xnor U28415 (N_28415,N_24891,N_24077);
or U28416 (N_28416,N_20305,N_23749);
nand U28417 (N_28417,N_20721,N_23996);
nand U28418 (N_28418,N_22901,N_21842);
or U28419 (N_28419,N_23725,N_21894);
and U28420 (N_28420,N_23578,N_21104);
and U28421 (N_28421,N_24383,N_21699);
nor U28422 (N_28422,N_21679,N_20246);
and U28423 (N_28423,N_23899,N_21494);
or U28424 (N_28424,N_23841,N_21771);
nand U28425 (N_28425,N_21099,N_24119);
nor U28426 (N_28426,N_24744,N_21398);
xnor U28427 (N_28427,N_20173,N_24228);
or U28428 (N_28428,N_21778,N_20742);
nor U28429 (N_28429,N_23723,N_20478);
xnor U28430 (N_28430,N_23467,N_24396);
or U28431 (N_28431,N_23722,N_23493);
nand U28432 (N_28432,N_24212,N_20084);
nand U28433 (N_28433,N_20799,N_21921);
nand U28434 (N_28434,N_22314,N_24669);
xor U28435 (N_28435,N_21631,N_20532);
and U28436 (N_28436,N_21700,N_20119);
and U28437 (N_28437,N_21216,N_23458);
or U28438 (N_28438,N_23287,N_21184);
or U28439 (N_28439,N_21838,N_24991);
or U28440 (N_28440,N_24559,N_23470);
and U28441 (N_28441,N_24779,N_22321);
and U28442 (N_28442,N_24431,N_21773);
and U28443 (N_28443,N_23836,N_21297);
nand U28444 (N_28444,N_22901,N_20906);
nand U28445 (N_28445,N_24721,N_23135);
nand U28446 (N_28446,N_24663,N_22154);
and U28447 (N_28447,N_24449,N_20678);
and U28448 (N_28448,N_23376,N_22538);
nor U28449 (N_28449,N_20940,N_22968);
nor U28450 (N_28450,N_22047,N_21252);
and U28451 (N_28451,N_24101,N_24959);
nand U28452 (N_28452,N_24770,N_20160);
or U28453 (N_28453,N_23679,N_22091);
and U28454 (N_28454,N_21328,N_22686);
nor U28455 (N_28455,N_20721,N_23261);
nand U28456 (N_28456,N_22468,N_22489);
xnor U28457 (N_28457,N_20908,N_21854);
or U28458 (N_28458,N_20371,N_20423);
nor U28459 (N_28459,N_21616,N_21647);
nor U28460 (N_28460,N_21760,N_23976);
and U28461 (N_28461,N_24558,N_22316);
xor U28462 (N_28462,N_20217,N_21392);
nor U28463 (N_28463,N_22311,N_20806);
nand U28464 (N_28464,N_23053,N_22305);
or U28465 (N_28465,N_23910,N_21049);
and U28466 (N_28466,N_20875,N_22523);
and U28467 (N_28467,N_20836,N_22101);
nor U28468 (N_28468,N_23183,N_20830);
and U28469 (N_28469,N_24153,N_22600);
nor U28470 (N_28470,N_24848,N_22717);
or U28471 (N_28471,N_20095,N_24227);
xnor U28472 (N_28472,N_24930,N_21234);
xnor U28473 (N_28473,N_20414,N_21465);
and U28474 (N_28474,N_24097,N_20735);
nor U28475 (N_28475,N_20049,N_21011);
nand U28476 (N_28476,N_20439,N_21297);
nor U28477 (N_28477,N_23625,N_24133);
nand U28478 (N_28478,N_23573,N_24345);
and U28479 (N_28479,N_21903,N_21664);
nand U28480 (N_28480,N_22294,N_20122);
nand U28481 (N_28481,N_24859,N_22857);
nor U28482 (N_28482,N_24022,N_20215);
or U28483 (N_28483,N_21000,N_22132);
or U28484 (N_28484,N_23555,N_23843);
xor U28485 (N_28485,N_23486,N_21366);
nor U28486 (N_28486,N_24840,N_22960);
or U28487 (N_28487,N_23850,N_23447);
nand U28488 (N_28488,N_23021,N_22025);
nor U28489 (N_28489,N_20784,N_23916);
nand U28490 (N_28490,N_22366,N_20275);
nor U28491 (N_28491,N_23947,N_23434);
nand U28492 (N_28492,N_21297,N_20584);
nand U28493 (N_28493,N_24393,N_22332);
xor U28494 (N_28494,N_21265,N_21687);
or U28495 (N_28495,N_22999,N_23212);
nand U28496 (N_28496,N_21179,N_22975);
nor U28497 (N_28497,N_24526,N_21614);
or U28498 (N_28498,N_23624,N_24373);
nor U28499 (N_28499,N_22698,N_21440);
or U28500 (N_28500,N_24441,N_22203);
nor U28501 (N_28501,N_23391,N_21736);
nor U28502 (N_28502,N_24594,N_23692);
or U28503 (N_28503,N_20460,N_24255);
or U28504 (N_28504,N_20952,N_23991);
and U28505 (N_28505,N_23641,N_21308);
or U28506 (N_28506,N_20124,N_24246);
and U28507 (N_28507,N_21856,N_21426);
and U28508 (N_28508,N_20922,N_20553);
nand U28509 (N_28509,N_20807,N_23668);
or U28510 (N_28510,N_21642,N_23762);
and U28511 (N_28511,N_20831,N_24189);
or U28512 (N_28512,N_22787,N_21256);
nor U28513 (N_28513,N_20857,N_23193);
or U28514 (N_28514,N_23821,N_22691);
or U28515 (N_28515,N_24535,N_21576);
nor U28516 (N_28516,N_21926,N_24268);
and U28517 (N_28517,N_20428,N_23474);
or U28518 (N_28518,N_20194,N_22077);
and U28519 (N_28519,N_24268,N_24461);
nor U28520 (N_28520,N_24693,N_20950);
or U28521 (N_28521,N_21929,N_20195);
nor U28522 (N_28522,N_24302,N_22873);
nand U28523 (N_28523,N_20587,N_24362);
nand U28524 (N_28524,N_23843,N_24597);
xor U28525 (N_28525,N_21332,N_24125);
nand U28526 (N_28526,N_21438,N_21439);
and U28527 (N_28527,N_23894,N_20775);
nand U28528 (N_28528,N_24532,N_24073);
or U28529 (N_28529,N_21021,N_22638);
and U28530 (N_28530,N_24899,N_20239);
and U28531 (N_28531,N_20337,N_23381);
nor U28532 (N_28532,N_21411,N_24651);
or U28533 (N_28533,N_23949,N_22913);
or U28534 (N_28534,N_22370,N_24776);
and U28535 (N_28535,N_20487,N_23288);
nor U28536 (N_28536,N_22232,N_20153);
and U28537 (N_28537,N_24095,N_23059);
and U28538 (N_28538,N_22568,N_23438);
and U28539 (N_28539,N_23465,N_21378);
nor U28540 (N_28540,N_22385,N_24112);
nand U28541 (N_28541,N_21190,N_24620);
or U28542 (N_28542,N_23682,N_21914);
nor U28543 (N_28543,N_24631,N_20185);
or U28544 (N_28544,N_23670,N_24853);
or U28545 (N_28545,N_22940,N_24382);
xnor U28546 (N_28546,N_20432,N_22396);
or U28547 (N_28547,N_23704,N_24467);
and U28548 (N_28548,N_22825,N_24594);
xor U28549 (N_28549,N_21116,N_23268);
and U28550 (N_28550,N_20534,N_20971);
or U28551 (N_28551,N_21205,N_24361);
nand U28552 (N_28552,N_21871,N_20647);
nand U28553 (N_28553,N_22108,N_24037);
nor U28554 (N_28554,N_20827,N_21997);
nand U28555 (N_28555,N_24498,N_20284);
nand U28556 (N_28556,N_20885,N_24968);
nor U28557 (N_28557,N_24204,N_20314);
or U28558 (N_28558,N_22723,N_20977);
nor U28559 (N_28559,N_21589,N_21141);
nand U28560 (N_28560,N_20920,N_22449);
nor U28561 (N_28561,N_22736,N_22576);
and U28562 (N_28562,N_20433,N_20107);
nand U28563 (N_28563,N_21460,N_21632);
nand U28564 (N_28564,N_22679,N_21821);
and U28565 (N_28565,N_23086,N_22435);
and U28566 (N_28566,N_21396,N_20137);
and U28567 (N_28567,N_21054,N_23406);
nand U28568 (N_28568,N_21919,N_24767);
and U28569 (N_28569,N_22459,N_23478);
nand U28570 (N_28570,N_23792,N_22213);
xnor U28571 (N_28571,N_23529,N_20947);
and U28572 (N_28572,N_20634,N_21954);
nand U28573 (N_28573,N_20530,N_24703);
or U28574 (N_28574,N_22726,N_20831);
and U28575 (N_28575,N_22893,N_22845);
nand U28576 (N_28576,N_22060,N_21147);
nor U28577 (N_28577,N_22682,N_20074);
nor U28578 (N_28578,N_22275,N_21076);
nand U28579 (N_28579,N_23071,N_23187);
nor U28580 (N_28580,N_23137,N_21475);
nand U28581 (N_28581,N_22248,N_21812);
nor U28582 (N_28582,N_24207,N_20186);
nand U28583 (N_28583,N_23953,N_20512);
nand U28584 (N_28584,N_21871,N_22423);
nand U28585 (N_28585,N_21979,N_24589);
nor U28586 (N_28586,N_20039,N_24570);
nand U28587 (N_28587,N_23639,N_23297);
nor U28588 (N_28588,N_22681,N_21329);
nor U28589 (N_28589,N_21976,N_23660);
nand U28590 (N_28590,N_22897,N_24775);
or U28591 (N_28591,N_24109,N_20954);
nor U28592 (N_28592,N_24127,N_21700);
and U28593 (N_28593,N_20243,N_22415);
or U28594 (N_28594,N_22645,N_21387);
and U28595 (N_28595,N_23037,N_22283);
nor U28596 (N_28596,N_21767,N_21091);
and U28597 (N_28597,N_20675,N_20578);
and U28598 (N_28598,N_20063,N_23758);
and U28599 (N_28599,N_21328,N_22737);
and U28600 (N_28600,N_21542,N_22085);
nand U28601 (N_28601,N_21477,N_20291);
or U28602 (N_28602,N_21605,N_23792);
nor U28603 (N_28603,N_20157,N_24447);
and U28604 (N_28604,N_23775,N_20957);
or U28605 (N_28605,N_20478,N_20624);
xnor U28606 (N_28606,N_20467,N_20799);
nor U28607 (N_28607,N_24407,N_23445);
nor U28608 (N_28608,N_24705,N_22121);
or U28609 (N_28609,N_24865,N_20478);
and U28610 (N_28610,N_20370,N_24442);
and U28611 (N_28611,N_24604,N_21273);
and U28612 (N_28612,N_22023,N_22037);
and U28613 (N_28613,N_22738,N_20105);
and U28614 (N_28614,N_23343,N_20694);
and U28615 (N_28615,N_23302,N_21423);
xnor U28616 (N_28616,N_22002,N_24389);
nand U28617 (N_28617,N_22638,N_22023);
xnor U28618 (N_28618,N_20446,N_23241);
nand U28619 (N_28619,N_21354,N_24408);
xnor U28620 (N_28620,N_22633,N_23848);
nand U28621 (N_28621,N_22713,N_24529);
nor U28622 (N_28622,N_20976,N_21038);
or U28623 (N_28623,N_20918,N_20714);
nand U28624 (N_28624,N_23673,N_24800);
and U28625 (N_28625,N_22638,N_23674);
and U28626 (N_28626,N_20185,N_21839);
or U28627 (N_28627,N_20794,N_20268);
nand U28628 (N_28628,N_22931,N_24383);
or U28629 (N_28629,N_23716,N_21495);
nor U28630 (N_28630,N_21381,N_24411);
or U28631 (N_28631,N_21481,N_21747);
nand U28632 (N_28632,N_24925,N_21599);
and U28633 (N_28633,N_21176,N_23250);
or U28634 (N_28634,N_21988,N_22051);
and U28635 (N_28635,N_20520,N_22897);
nor U28636 (N_28636,N_20877,N_22093);
and U28637 (N_28637,N_22484,N_23467);
nor U28638 (N_28638,N_20352,N_22775);
and U28639 (N_28639,N_23428,N_21089);
xor U28640 (N_28640,N_23695,N_22939);
nand U28641 (N_28641,N_20055,N_20592);
or U28642 (N_28642,N_22141,N_23929);
nand U28643 (N_28643,N_21429,N_20198);
nand U28644 (N_28644,N_20661,N_22338);
nand U28645 (N_28645,N_22542,N_24877);
and U28646 (N_28646,N_24878,N_23504);
and U28647 (N_28647,N_20110,N_22585);
nand U28648 (N_28648,N_21127,N_24963);
xor U28649 (N_28649,N_23120,N_20200);
or U28650 (N_28650,N_20394,N_24047);
nand U28651 (N_28651,N_23714,N_22217);
nor U28652 (N_28652,N_23989,N_22892);
nor U28653 (N_28653,N_20232,N_23274);
or U28654 (N_28654,N_21857,N_23239);
or U28655 (N_28655,N_24849,N_21388);
nand U28656 (N_28656,N_22079,N_21139);
nand U28657 (N_28657,N_24857,N_21288);
nand U28658 (N_28658,N_21823,N_23628);
nand U28659 (N_28659,N_20325,N_20826);
or U28660 (N_28660,N_23245,N_23717);
and U28661 (N_28661,N_23115,N_21978);
nand U28662 (N_28662,N_22943,N_24927);
nor U28663 (N_28663,N_20790,N_23455);
nor U28664 (N_28664,N_23258,N_20493);
and U28665 (N_28665,N_24494,N_24793);
and U28666 (N_28666,N_23529,N_21699);
and U28667 (N_28667,N_23742,N_20630);
xor U28668 (N_28668,N_22726,N_20430);
and U28669 (N_28669,N_22118,N_22240);
and U28670 (N_28670,N_23180,N_22920);
or U28671 (N_28671,N_22224,N_23196);
and U28672 (N_28672,N_24558,N_20915);
or U28673 (N_28673,N_24912,N_24623);
or U28674 (N_28674,N_22288,N_24327);
and U28675 (N_28675,N_22366,N_21980);
nor U28676 (N_28676,N_23664,N_20953);
or U28677 (N_28677,N_20434,N_22344);
nand U28678 (N_28678,N_20640,N_23082);
nand U28679 (N_28679,N_20752,N_20640);
nand U28680 (N_28680,N_22425,N_21892);
and U28681 (N_28681,N_21642,N_21761);
or U28682 (N_28682,N_24298,N_21668);
nor U28683 (N_28683,N_20327,N_20554);
and U28684 (N_28684,N_22020,N_21778);
or U28685 (N_28685,N_22440,N_22264);
and U28686 (N_28686,N_21450,N_24300);
xnor U28687 (N_28687,N_24993,N_22099);
nor U28688 (N_28688,N_24194,N_22694);
and U28689 (N_28689,N_21315,N_23583);
and U28690 (N_28690,N_20135,N_20035);
xnor U28691 (N_28691,N_21357,N_24630);
nand U28692 (N_28692,N_24980,N_24142);
nor U28693 (N_28693,N_23329,N_21907);
or U28694 (N_28694,N_23589,N_23475);
and U28695 (N_28695,N_24786,N_21815);
or U28696 (N_28696,N_23811,N_22133);
and U28697 (N_28697,N_23218,N_21340);
or U28698 (N_28698,N_24656,N_20502);
nor U28699 (N_28699,N_24904,N_20629);
nor U28700 (N_28700,N_24509,N_20493);
or U28701 (N_28701,N_22329,N_24677);
nor U28702 (N_28702,N_22758,N_24135);
and U28703 (N_28703,N_24162,N_22022);
and U28704 (N_28704,N_23074,N_22821);
and U28705 (N_28705,N_21637,N_23943);
xor U28706 (N_28706,N_21581,N_21099);
nor U28707 (N_28707,N_24686,N_22550);
nand U28708 (N_28708,N_21851,N_21106);
or U28709 (N_28709,N_22917,N_22814);
xnor U28710 (N_28710,N_23689,N_22041);
and U28711 (N_28711,N_22759,N_24037);
or U28712 (N_28712,N_23278,N_21999);
xor U28713 (N_28713,N_21799,N_23500);
or U28714 (N_28714,N_21202,N_20389);
or U28715 (N_28715,N_23613,N_20985);
and U28716 (N_28716,N_22187,N_22717);
nand U28717 (N_28717,N_21033,N_24889);
xnor U28718 (N_28718,N_22801,N_21699);
xnor U28719 (N_28719,N_22476,N_22669);
or U28720 (N_28720,N_22188,N_24781);
nand U28721 (N_28721,N_20029,N_24921);
and U28722 (N_28722,N_20706,N_22935);
or U28723 (N_28723,N_23974,N_23269);
or U28724 (N_28724,N_24171,N_22718);
and U28725 (N_28725,N_23302,N_24531);
xnor U28726 (N_28726,N_24896,N_23648);
or U28727 (N_28727,N_24131,N_20564);
or U28728 (N_28728,N_23476,N_21411);
or U28729 (N_28729,N_22439,N_21609);
nand U28730 (N_28730,N_24084,N_20740);
nand U28731 (N_28731,N_24846,N_24222);
and U28732 (N_28732,N_23257,N_22676);
and U28733 (N_28733,N_22688,N_21240);
and U28734 (N_28734,N_21085,N_24034);
nand U28735 (N_28735,N_24946,N_21879);
xor U28736 (N_28736,N_22637,N_20449);
and U28737 (N_28737,N_21106,N_24040);
and U28738 (N_28738,N_22101,N_22565);
nor U28739 (N_28739,N_22818,N_20166);
nor U28740 (N_28740,N_20893,N_22588);
or U28741 (N_28741,N_21643,N_22937);
xnor U28742 (N_28742,N_20185,N_22512);
and U28743 (N_28743,N_20979,N_23388);
and U28744 (N_28744,N_20928,N_20767);
or U28745 (N_28745,N_22168,N_23750);
or U28746 (N_28746,N_20339,N_21093);
and U28747 (N_28747,N_23701,N_24822);
xnor U28748 (N_28748,N_24782,N_20374);
nand U28749 (N_28749,N_22642,N_22782);
or U28750 (N_28750,N_22971,N_24531);
nor U28751 (N_28751,N_21317,N_20695);
xnor U28752 (N_28752,N_20469,N_23186);
and U28753 (N_28753,N_24268,N_22929);
nor U28754 (N_28754,N_20569,N_21819);
nor U28755 (N_28755,N_21511,N_20333);
xnor U28756 (N_28756,N_21061,N_20689);
and U28757 (N_28757,N_20389,N_21978);
nor U28758 (N_28758,N_23429,N_21734);
or U28759 (N_28759,N_20712,N_23218);
and U28760 (N_28760,N_22006,N_24420);
and U28761 (N_28761,N_23038,N_20743);
or U28762 (N_28762,N_21240,N_22003);
nand U28763 (N_28763,N_22339,N_20311);
and U28764 (N_28764,N_24335,N_22546);
nand U28765 (N_28765,N_23928,N_24689);
nand U28766 (N_28766,N_20382,N_23483);
or U28767 (N_28767,N_21676,N_23848);
and U28768 (N_28768,N_24967,N_22050);
nor U28769 (N_28769,N_23265,N_23654);
xnor U28770 (N_28770,N_24470,N_24202);
and U28771 (N_28771,N_20300,N_23752);
and U28772 (N_28772,N_20586,N_23948);
nand U28773 (N_28773,N_22854,N_20726);
nor U28774 (N_28774,N_22845,N_23161);
xnor U28775 (N_28775,N_20382,N_21019);
nor U28776 (N_28776,N_20691,N_21444);
nor U28777 (N_28777,N_20079,N_22755);
nand U28778 (N_28778,N_21022,N_21587);
or U28779 (N_28779,N_22879,N_20882);
xnor U28780 (N_28780,N_24445,N_20019);
nor U28781 (N_28781,N_23387,N_21465);
nor U28782 (N_28782,N_21510,N_22350);
nor U28783 (N_28783,N_23498,N_23213);
or U28784 (N_28784,N_24612,N_21992);
nor U28785 (N_28785,N_22587,N_20217);
and U28786 (N_28786,N_23194,N_21831);
xnor U28787 (N_28787,N_24905,N_22130);
or U28788 (N_28788,N_22499,N_20413);
xor U28789 (N_28789,N_21429,N_21474);
nor U28790 (N_28790,N_20590,N_24391);
nor U28791 (N_28791,N_23623,N_24498);
and U28792 (N_28792,N_20427,N_20141);
xnor U28793 (N_28793,N_24600,N_21078);
or U28794 (N_28794,N_23014,N_22947);
nand U28795 (N_28795,N_24373,N_22651);
nand U28796 (N_28796,N_23436,N_21927);
xor U28797 (N_28797,N_24571,N_20424);
xor U28798 (N_28798,N_20749,N_24015);
and U28799 (N_28799,N_24417,N_20030);
nor U28800 (N_28800,N_22062,N_21167);
or U28801 (N_28801,N_24172,N_20773);
nor U28802 (N_28802,N_23314,N_23689);
and U28803 (N_28803,N_23026,N_20792);
and U28804 (N_28804,N_24830,N_23293);
nor U28805 (N_28805,N_21889,N_23231);
and U28806 (N_28806,N_20709,N_23050);
nor U28807 (N_28807,N_23260,N_21458);
and U28808 (N_28808,N_21021,N_21135);
nand U28809 (N_28809,N_22017,N_24442);
nand U28810 (N_28810,N_22709,N_20573);
nor U28811 (N_28811,N_21377,N_24935);
nand U28812 (N_28812,N_24253,N_22469);
nand U28813 (N_28813,N_21189,N_23895);
nor U28814 (N_28814,N_22187,N_24569);
nand U28815 (N_28815,N_23631,N_22901);
nand U28816 (N_28816,N_21839,N_22757);
nand U28817 (N_28817,N_23313,N_23907);
xnor U28818 (N_28818,N_20423,N_23503);
and U28819 (N_28819,N_20980,N_20856);
or U28820 (N_28820,N_21719,N_23643);
and U28821 (N_28821,N_20718,N_21157);
nand U28822 (N_28822,N_20484,N_23403);
xnor U28823 (N_28823,N_22941,N_21448);
nor U28824 (N_28824,N_20229,N_21372);
nand U28825 (N_28825,N_20104,N_22488);
nor U28826 (N_28826,N_24509,N_21994);
and U28827 (N_28827,N_23296,N_22105);
or U28828 (N_28828,N_24588,N_24424);
nor U28829 (N_28829,N_22127,N_22084);
and U28830 (N_28830,N_24017,N_22651);
or U28831 (N_28831,N_20416,N_22328);
nor U28832 (N_28832,N_20906,N_24261);
nand U28833 (N_28833,N_21394,N_20447);
nand U28834 (N_28834,N_20246,N_20211);
or U28835 (N_28835,N_20551,N_21510);
nand U28836 (N_28836,N_23229,N_23441);
nand U28837 (N_28837,N_23254,N_23871);
nor U28838 (N_28838,N_21410,N_21329);
and U28839 (N_28839,N_20307,N_20940);
and U28840 (N_28840,N_23840,N_24198);
nor U28841 (N_28841,N_22161,N_22743);
xor U28842 (N_28842,N_23190,N_21734);
and U28843 (N_28843,N_20373,N_23648);
or U28844 (N_28844,N_20810,N_21240);
nand U28845 (N_28845,N_24870,N_21335);
nand U28846 (N_28846,N_24790,N_21256);
nor U28847 (N_28847,N_21086,N_24531);
xor U28848 (N_28848,N_22837,N_24484);
nor U28849 (N_28849,N_22582,N_22799);
or U28850 (N_28850,N_24489,N_20500);
nor U28851 (N_28851,N_24434,N_23393);
or U28852 (N_28852,N_23054,N_20937);
nand U28853 (N_28853,N_22583,N_21466);
and U28854 (N_28854,N_20793,N_23991);
nand U28855 (N_28855,N_23506,N_21901);
and U28856 (N_28856,N_24348,N_20384);
nor U28857 (N_28857,N_21912,N_23487);
and U28858 (N_28858,N_23134,N_23161);
nor U28859 (N_28859,N_24949,N_20219);
and U28860 (N_28860,N_22411,N_23499);
nor U28861 (N_28861,N_23458,N_21436);
nand U28862 (N_28862,N_22081,N_22049);
nand U28863 (N_28863,N_24545,N_21349);
nand U28864 (N_28864,N_22300,N_24920);
nor U28865 (N_28865,N_20727,N_24080);
nor U28866 (N_28866,N_20675,N_22911);
nand U28867 (N_28867,N_21204,N_22101);
xnor U28868 (N_28868,N_23765,N_24494);
nor U28869 (N_28869,N_21657,N_23405);
and U28870 (N_28870,N_23524,N_22052);
nand U28871 (N_28871,N_24642,N_24389);
nand U28872 (N_28872,N_21486,N_20990);
and U28873 (N_28873,N_20778,N_24110);
and U28874 (N_28874,N_21376,N_23690);
and U28875 (N_28875,N_23406,N_23549);
or U28876 (N_28876,N_23896,N_24591);
nand U28877 (N_28877,N_23323,N_21432);
and U28878 (N_28878,N_20452,N_20079);
xnor U28879 (N_28879,N_23973,N_24000);
nand U28880 (N_28880,N_21888,N_23085);
or U28881 (N_28881,N_24874,N_22274);
nor U28882 (N_28882,N_21737,N_23031);
nand U28883 (N_28883,N_24122,N_23047);
or U28884 (N_28884,N_24331,N_24353);
nor U28885 (N_28885,N_22776,N_22328);
nand U28886 (N_28886,N_24359,N_20282);
nor U28887 (N_28887,N_21909,N_23857);
nand U28888 (N_28888,N_21459,N_24607);
nor U28889 (N_28889,N_24360,N_21442);
and U28890 (N_28890,N_22806,N_20016);
nand U28891 (N_28891,N_21955,N_20759);
nor U28892 (N_28892,N_21471,N_24939);
nor U28893 (N_28893,N_22514,N_23839);
and U28894 (N_28894,N_22308,N_21997);
nand U28895 (N_28895,N_22391,N_20430);
or U28896 (N_28896,N_24572,N_24079);
nor U28897 (N_28897,N_22320,N_22108);
and U28898 (N_28898,N_20593,N_23276);
nor U28899 (N_28899,N_23874,N_20671);
or U28900 (N_28900,N_24234,N_22198);
nand U28901 (N_28901,N_24920,N_24619);
nor U28902 (N_28902,N_24518,N_20078);
nor U28903 (N_28903,N_23853,N_21760);
nand U28904 (N_28904,N_24503,N_20508);
nor U28905 (N_28905,N_22600,N_24350);
or U28906 (N_28906,N_23020,N_24397);
nand U28907 (N_28907,N_23802,N_23458);
nor U28908 (N_28908,N_24614,N_20824);
nand U28909 (N_28909,N_23957,N_20347);
nor U28910 (N_28910,N_20863,N_22818);
nor U28911 (N_28911,N_22608,N_20074);
or U28912 (N_28912,N_20830,N_20854);
or U28913 (N_28913,N_22981,N_22835);
or U28914 (N_28914,N_24312,N_24613);
nand U28915 (N_28915,N_23027,N_20415);
nor U28916 (N_28916,N_21435,N_20115);
xor U28917 (N_28917,N_24749,N_24210);
nand U28918 (N_28918,N_23542,N_22876);
nor U28919 (N_28919,N_24112,N_21299);
and U28920 (N_28920,N_23129,N_24364);
or U28921 (N_28921,N_20438,N_24612);
nor U28922 (N_28922,N_23679,N_22650);
or U28923 (N_28923,N_24132,N_23965);
and U28924 (N_28924,N_22166,N_21009);
nor U28925 (N_28925,N_21894,N_23314);
nand U28926 (N_28926,N_20290,N_23829);
nor U28927 (N_28927,N_24083,N_23348);
or U28928 (N_28928,N_22838,N_23523);
or U28929 (N_28929,N_20957,N_20722);
xor U28930 (N_28930,N_21898,N_20446);
or U28931 (N_28931,N_22536,N_22502);
or U28932 (N_28932,N_20038,N_23874);
nand U28933 (N_28933,N_23778,N_21883);
nor U28934 (N_28934,N_24356,N_22643);
nand U28935 (N_28935,N_20517,N_21857);
nand U28936 (N_28936,N_23334,N_23532);
or U28937 (N_28937,N_20163,N_21113);
and U28938 (N_28938,N_20189,N_21599);
nand U28939 (N_28939,N_22698,N_22901);
nand U28940 (N_28940,N_22920,N_20485);
and U28941 (N_28941,N_21477,N_20277);
or U28942 (N_28942,N_20431,N_22104);
or U28943 (N_28943,N_21500,N_22381);
nand U28944 (N_28944,N_22804,N_21951);
nor U28945 (N_28945,N_24197,N_21508);
nand U28946 (N_28946,N_22400,N_22566);
or U28947 (N_28947,N_24466,N_23712);
nand U28948 (N_28948,N_20341,N_20698);
nand U28949 (N_28949,N_22707,N_20695);
or U28950 (N_28950,N_24912,N_22218);
and U28951 (N_28951,N_24057,N_22626);
or U28952 (N_28952,N_23760,N_24266);
nand U28953 (N_28953,N_23713,N_22105);
nand U28954 (N_28954,N_23149,N_23788);
or U28955 (N_28955,N_21202,N_22070);
nand U28956 (N_28956,N_21667,N_24913);
and U28957 (N_28957,N_21844,N_23748);
nor U28958 (N_28958,N_22495,N_21997);
or U28959 (N_28959,N_21054,N_22548);
or U28960 (N_28960,N_20233,N_23779);
nor U28961 (N_28961,N_23294,N_20671);
nand U28962 (N_28962,N_23269,N_22283);
or U28963 (N_28963,N_21504,N_22696);
xnor U28964 (N_28964,N_24859,N_23014);
or U28965 (N_28965,N_21946,N_23214);
or U28966 (N_28966,N_22196,N_24998);
or U28967 (N_28967,N_22172,N_21678);
or U28968 (N_28968,N_24782,N_22080);
nor U28969 (N_28969,N_22269,N_23430);
nand U28970 (N_28970,N_21036,N_20797);
and U28971 (N_28971,N_20512,N_20798);
nor U28972 (N_28972,N_22128,N_23866);
nor U28973 (N_28973,N_22594,N_23480);
and U28974 (N_28974,N_22533,N_22557);
nand U28975 (N_28975,N_22079,N_20096);
or U28976 (N_28976,N_24106,N_21351);
nor U28977 (N_28977,N_24726,N_23023);
or U28978 (N_28978,N_23579,N_21941);
nand U28979 (N_28979,N_21691,N_22456);
nor U28980 (N_28980,N_24765,N_24042);
and U28981 (N_28981,N_20164,N_21086);
nor U28982 (N_28982,N_20162,N_22116);
and U28983 (N_28983,N_20568,N_21120);
xnor U28984 (N_28984,N_23564,N_24894);
nor U28985 (N_28985,N_24516,N_22392);
or U28986 (N_28986,N_22931,N_20143);
nand U28987 (N_28987,N_21874,N_22309);
xor U28988 (N_28988,N_21637,N_24526);
xnor U28989 (N_28989,N_23744,N_23211);
and U28990 (N_28990,N_20475,N_24860);
nand U28991 (N_28991,N_24110,N_24541);
or U28992 (N_28992,N_23330,N_23031);
or U28993 (N_28993,N_21413,N_21664);
nor U28994 (N_28994,N_23344,N_23831);
or U28995 (N_28995,N_21209,N_20979);
or U28996 (N_28996,N_20069,N_21803);
nor U28997 (N_28997,N_21712,N_22039);
nor U28998 (N_28998,N_24013,N_24337);
or U28999 (N_28999,N_21791,N_21115);
nor U29000 (N_29000,N_23882,N_20621);
nor U29001 (N_29001,N_20539,N_24375);
nand U29002 (N_29002,N_20938,N_22921);
or U29003 (N_29003,N_23535,N_23247);
and U29004 (N_29004,N_20705,N_21963);
and U29005 (N_29005,N_21204,N_20694);
and U29006 (N_29006,N_22787,N_21807);
or U29007 (N_29007,N_21558,N_22344);
nor U29008 (N_29008,N_21402,N_22553);
or U29009 (N_29009,N_21001,N_20434);
or U29010 (N_29010,N_24095,N_24756);
nor U29011 (N_29011,N_24637,N_22357);
or U29012 (N_29012,N_20345,N_24130);
and U29013 (N_29013,N_23139,N_24464);
or U29014 (N_29014,N_21883,N_24383);
nand U29015 (N_29015,N_21175,N_22676);
or U29016 (N_29016,N_21685,N_24841);
nand U29017 (N_29017,N_23807,N_24693);
and U29018 (N_29018,N_22645,N_21366);
and U29019 (N_29019,N_24836,N_22383);
nor U29020 (N_29020,N_20297,N_20064);
or U29021 (N_29021,N_20141,N_23422);
nor U29022 (N_29022,N_23138,N_23646);
and U29023 (N_29023,N_20005,N_23396);
or U29024 (N_29024,N_24500,N_21931);
nor U29025 (N_29025,N_24863,N_23324);
nand U29026 (N_29026,N_20204,N_22126);
or U29027 (N_29027,N_21015,N_22002);
nand U29028 (N_29028,N_23109,N_20483);
nor U29029 (N_29029,N_22444,N_23011);
and U29030 (N_29030,N_23494,N_22705);
or U29031 (N_29031,N_23205,N_22903);
nor U29032 (N_29032,N_22043,N_24512);
xnor U29033 (N_29033,N_23536,N_24995);
and U29034 (N_29034,N_24998,N_23866);
or U29035 (N_29035,N_22154,N_22669);
nand U29036 (N_29036,N_22646,N_20427);
nor U29037 (N_29037,N_23459,N_20647);
xnor U29038 (N_29038,N_23047,N_23016);
and U29039 (N_29039,N_20601,N_21882);
and U29040 (N_29040,N_20592,N_20919);
and U29041 (N_29041,N_20746,N_21276);
nor U29042 (N_29042,N_24518,N_23697);
or U29043 (N_29043,N_23962,N_24613);
xnor U29044 (N_29044,N_21463,N_23804);
xnor U29045 (N_29045,N_20856,N_20246);
or U29046 (N_29046,N_24607,N_22207);
nand U29047 (N_29047,N_22282,N_23936);
nand U29048 (N_29048,N_21895,N_21468);
and U29049 (N_29049,N_23322,N_20206);
nand U29050 (N_29050,N_22938,N_20435);
nand U29051 (N_29051,N_21029,N_20094);
nand U29052 (N_29052,N_23635,N_22574);
nor U29053 (N_29053,N_21643,N_24364);
and U29054 (N_29054,N_24519,N_20404);
or U29055 (N_29055,N_23938,N_24946);
nand U29056 (N_29056,N_23982,N_23706);
and U29057 (N_29057,N_21184,N_21492);
xnor U29058 (N_29058,N_21743,N_20508);
nand U29059 (N_29059,N_20031,N_20767);
xor U29060 (N_29060,N_21596,N_23145);
and U29061 (N_29061,N_22463,N_22349);
nand U29062 (N_29062,N_23727,N_21652);
nand U29063 (N_29063,N_20621,N_21557);
nand U29064 (N_29064,N_23705,N_22647);
or U29065 (N_29065,N_24060,N_23210);
nor U29066 (N_29066,N_20703,N_21435);
nand U29067 (N_29067,N_20335,N_23799);
nand U29068 (N_29068,N_23944,N_24692);
nand U29069 (N_29069,N_20828,N_21220);
nor U29070 (N_29070,N_22112,N_24501);
xor U29071 (N_29071,N_23827,N_22593);
nand U29072 (N_29072,N_24233,N_23654);
nand U29073 (N_29073,N_21119,N_22235);
nand U29074 (N_29074,N_20896,N_24042);
or U29075 (N_29075,N_21767,N_24340);
or U29076 (N_29076,N_22593,N_24503);
nand U29077 (N_29077,N_23454,N_20213);
and U29078 (N_29078,N_23475,N_22835);
nand U29079 (N_29079,N_22648,N_20110);
or U29080 (N_29080,N_21880,N_23931);
nand U29081 (N_29081,N_24377,N_20080);
nand U29082 (N_29082,N_21483,N_23444);
and U29083 (N_29083,N_21723,N_23349);
xnor U29084 (N_29084,N_24067,N_23739);
and U29085 (N_29085,N_21650,N_20271);
nand U29086 (N_29086,N_24707,N_24081);
and U29087 (N_29087,N_23413,N_23657);
or U29088 (N_29088,N_24569,N_22472);
or U29089 (N_29089,N_23248,N_24362);
xnor U29090 (N_29090,N_20874,N_24207);
nor U29091 (N_29091,N_21827,N_20259);
or U29092 (N_29092,N_24065,N_21975);
xor U29093 (N_29093,N_21234,N_22322);
and U29094 (N_29094,N_24105,N_22363);
or U29095 (N_29095,N_21796,N_22613);
nand U29096 (N_29096,N_22892,N_22200);
nand U29097 (N_29097,N_23925,N_24650);
nor U29098 (N_29098,N_24020,N_22398);
nand U29099 (N_29099,N_24749,N_24781);
xnor U29100 (N_29100,N_22462,N_23676);
or U29101 (N_29101,N_22391,N_20816);
nor U29102 (N_29102,N_21365,N_23021);
nor U29103 (N_29103,N_22931,N_21291);
nand U29104 (N_29104,N_22039,N_23169);
nor U29105 (N_29105,N_22651,N_23430);
or U29106 (N_29106,N_20194,N_21692);
nor U29107 (N_29107,N_21317,N_22996);
xor U29108 (N_29108,N_24154,N_21212);
nor U29109 (N_29109,N_22672,N_24006);
nand U29110 (N_29110,N_21016,N_21706);
or U29111 (N_29111,N_21170,N_22876);
or U29112 (N_29112,N_23796,N_20880);
and U29113 (N_29113,N_23633,N_21148);
or U29114 (N_29114,N_23570,N_22458);
or U29115 (N_29115,N_24474,N_21966);
xor U29116 (N_29116,N_21675,N_21572);
and U29117 (N_29117,N_20738,N_20858);
nor U29118 (N_29118,N_20437,N_23358);
nor U29119 (N_29119,N_23956,N_23505);
and U29120 (N_29120,N_20700,N_23257);
nor U29121 (N_29121,N_24717,N_23556);
and U29122 (N_29122,N_24908,N_24325);
or U29123 (N_29123,N_23630,N_22314);
nand U29124 (N_29124,N_22710,N_20114);
nor U29125 (N_29125,N_24334,N_23353);
or U29126 (N_29126,N_22841,N_21938);
nand U29127 (N_29127,N_20011,N_23450);
and U29128 (N_29128,N_20951,N_20400);
or U29129 (N_29129,N_20004,N_22803);
nor U29130 (N_29130,N_24685,N_23911);
nor U29131 (N_29131,N_23159,N_21097);
nor U29132 (N_29132,N_21944,N_21940);
or U29133 (N_29133,N_24073,N_23645);
or U29134 (N_29134,N_23207,N_23833);
or U29135 (N_29135,N_22125,N_20651);
or U29136 (N_29136,N_24327,N_23770);
or U29137 (N_29137,N_21859,N_22720);
xor U29138 (N_29138,N_21448,N_24670);
and U29139 (N_29139,N_20400,N_24581);
nor U29140 (N_29140,N_21556,N_21978);
nand U29141 (N_29141,N_20341,N_24913);
xor U29142 (N_29142,N_22527,N_24486);
and U29143 (N_29143,N_23662,N_23699);
nor U29144 (N_29144,N_20891,N_21081);
nand U29145 (N_29145,N_20268,N_23601);
or U29146 (N_29146,N_24313,N_22051);
or U29147 (N_29147,N_22334,N_20458);
nor U29148 (N_29148,N_20715,N_22968);
and U29149 (N_29149,N_24390,N_20484);
xor U29150 (N_29150,N_24840,N_22884);
nor U29151 (N_29151,N_21509,N_21706);
or U29152 (N_29152,N_22578,N_22025);
and U29153 (N_29153,N_20185,N_22941);
nor U29154 (N_29154,N_21592,N_21801);
and U29155 (N_29155,N_20008,N_24885);
and U29156 (N_29156,N_21699,N_22886);
or U29157 (N_29157,N_23749,N_21323);
or U29158 (N_29158,N_24579,N_20928);
nand U29159 (N_29159,N_21550,N_21553);
nor U29160 (N_29160,N_20429,N_24181);
nor U29161 (N_29161,N_24339,N_24626);
nor U29162 (N_29162,N_24546,N_24176);
nor U29163 (N_29163,N_21289,N_24304);
nand U29164 (N_29164,N_20407,N_23435);
nand U29165 (N_29165,N_24024,N_23423);
and U29166 (N_29166,N_21999,N_24924);
xor U29167 (N_29167,N_21639,N_23191);
or U29168 (N_29168,N_20189,N_21776);
nor U29169 (N_29169,N_22409,N_20357);
xnor U29170 (N_29170,N_21169,N_20684);
and U29171 (N_29171,N_24565,N_20898);
and U29172 (N_29172,N_23586,N_24601);
nor U29173 (N_29173,N_22086,N_20085);
xnor U29174 (N_29174,N_22679,N_24090);
nand U29175 (N_29175,N_21483,N_20787);
nor U29176 (N_29176,N_22434,N_21223);
or U29177 (N_29177,N_20205,N_23432);
or U29178 (N_29178,N_21195,N_23036);
nor U29179 (N_29179,N_21672,N_20828);
or U29180 (N_29180,N_20414,N_23298);
or U29181 (N_29181,N_22168,N_23111);
or U29182 (N_29182,N_24604,N_24364);
nand U29183 (N_29183,N_23720,N_24004);
or U29184 (N_29184,N_23317,N_24780);
nand U29185 (N_29185,N_20369,N_22237);
and U29186 (N_29186,N_20309,N_20564);
and U29187 (N_29187,N_24222,N_24161);
or U29188 (N_29188,N_22606,N_22183);
and U29189 (N_29189,N_24972,N_24867);
nor U29190 (N_29190,N_22186,N_23405);
nand U29191 (N_29191,N_24008,N_20754);
or U29192 (N_29192,N_21616,N_24028);
and U29193 (N_29193,N_24803,N_22132);
or U29194 (N_29194,N_20343,N_22223);
nand U29195 (N_29195,N_20115,N_24654);
xnor U29196 (N_29196,N_23645,N_20823);
nand U29197 (N_29197,N_21750,N_21095);
and U29198 (N_29198,N_21053,N_20367);
nor U29199 (N_29199,N_20379,N_20662);
and U29200 (N_29200,N_21714,N_24365);
nand U29201 (N_29201,N_23514,N_23902);
or U29202 (N_29202,N_22164,N_24212);
nand U29203 (N_29203,N_23527,N_23587);
and U29204 (N_29204,N_21578,N_23967);
and U29205 (N_29205,N_22991,N_24915);
and U29206 (N_29206,N_20712,N_23341);
or U29207 (N_29207,N_21003,N_22217);
nand U29208 (N_29208,N_23892,N_22720);
or U29209 (N_29209,N_24204,N_21996);
xor U29210 (N_29210,N_22223,N_24202);
and U29211 (N_29211,N_24406,N_21707);
and U29212 (N_29212,N_21091,N_20246);
or U29213 (N_29213,N_22894,N_22588);
or U29214 (N_29214,N_22142,N_23581);
or U29215 (N_29215,N_22882,N_21386);
and U29216 (N_29216,N_20830,N_23711);
nand U29217 (N_29217,N_20490,N_20794);
nand U29218 (N_29218,N_20776,N_21602);
or U29219 (N_29219,N_24933,N_20976);
nand U29220 (N_29220,N_23999,N_20176);
and U29221 (N_29221,N_24573,N_24903);
xor U29222 (N_29222,N_23786,N_23646);
or U29223 (N_29223,N_24290,N_20557);
or U29224 (N_29224,N_22181,N_23136);
nor U29225 (N_29225,N_20681,N_20321);
xor U29226 (N_29226,N_21536,N_21598);
nand U29227 (N_29227,N_23311,N_24781);
and U29228 (N_29228,N_20812,N_22443);
and U29229 (N_29229,N_23222,N_20911);
xnor U29230 (N_29230,N_24164,N_22461);
nor U29231 (N_29231,N_23789,N_24898);
and U29232 (N_29232,N_22324,N_23035);
xor U29233 (N_29233,N_24047,N_23995);
or U29234 (N_29234,N_23434,N_22482);
xor U29235 (N_29235,N_23084,N_24915);
or U29236 (N_29236,N_20090,N_23864);
and U29237 (N_29237,N_24447,N_22865);
nand U29238 (N_29238,N_21315,N_23455);
or U29239 (N_29239,N_23746,N_22280);
nor U29240 (N_29240,N_21311,N_22983);
nor U29241 (N_29241,N_20603,N_23390);
xor U29242 (N_29242,N_20817,N_20380);
and U29243 (N_29243,N_20965,N_22025);
or U29244 (N_29244,N_21627,N_21103);
nor U29245 (N_29245,N_24002,N_21656);
or U29246 (N_29246,N_24956,N_23973);
and U29247 (N_29247,N_22082,N_22414);
nand U29248 (N_29248,N_24801,N_24507);
nor U29249 (N_29249,N_23440,N_21507);
nor U29250 (N_29250,N_24436,N_24697);
and U29251 (N_29251,N_23185,N_23221);
or U29252 (N_29252,N_23643,N_24036);
or U29253 (N_29253,N_20411,N_20835);
or U29254 (N_29254,N_23134,N_23590);
or U29255 (N_29255,N_20368,N_22574);
and U29256 (N_29256,N_24777,N_23962);
and U29257 (N_29257,N_21497,N_23137);
nor U29258 (N_29258,N_24694,N_20240);
or U29259 (N_29259,N_21435,N_20887);
and U29260 (N_29260,N_21001,N_21592);
nor U29261 (N_29261,N_21680,N_20742);
nor U29262 (N_29262,N_20752,N_21794);
nand U29263 (N_29263,N_20906,N_22158);
nor U29264 (N_29264,N_22595,N_22705);
or U29265 (N_29265,N_20413,N_21608);
and U29266 (N_29266,N_21780,N_21790);
or U29267 (N_29267,N_23850,N_23521);
nor U29268 (N_29268,N_21583,N_23857);
and U29269 (N_29269,N_21681,N_24459);
nor U29270 (N_29270,N_21153,N_23104);
or U29271 (N_29271,N_23445,N_24977);
or U29272 (N_29272,N_20973,N_23107);
nand U29273 (N_29273,N_22578,N_24918);
and U29274 (N_29274,N_20854,N_21037);
or U29275 (N_29275,N_20826,N_24092);
nand U29276 (N_29276,N_20801,N_20424);
nor U29277 (N_29277,N_24829,N_20630);
xnor U29278 (N_29278,N_23160,N_23260);
or U29279 (N_29279,N_24699,N_23019);
nor U29280 (N_29280,N_24318,N_23176);
and U29281 (N_29281,N_20362,N_23073);
nor U29282 (N_29282,N_24004,N_20173);
or U29283 (N_29283,N_21223,N_24631);
nor U29284 (N_29284,N_23826,N_24608);
nand U29285 (N_29285,N_20765,N_22024);
nand U29286 (N_29286,N_20880,N_20988);
and U29287 (N_29287,N_20076,N_24103);
or U29288 (N_29288,N_22003,N_20600);
nand U29289 (N_29289,N_20251,N_24843);
or U29290 (N_29290,N_21464,N_23183);
xnor U29291 (N_29291,N_23177,N_22724);
and U29292 (N_29292,N_22098,N_24336);
nor U29293 (N_29293,N_20445,N_22335);
and U29294 (N_29294,N_21564,N_22761);
and U29295 (N_29295,N_23789,N_20515);
and U29296 (N_29296,N_24651,N_22199);
nand U29297 (N_29297,N_23295,N_24672);
or U29298 (N_29298,N_21087,N_20230);
or U29299 (N_29299,N_23336,N_20497);
and U29300 (N_29300,N_22326,N_20207);
nand U29301 (N_29301,N_22045,N_24408);
or U29302 (N_29302,N_20009,N_20137);
and U29303 (N_29303,N_22914,N_20693);
xnor U29304 (N_29304,N_24999,N_21895);
or U29305 (N_29305,N_24352,N_22461);
or U29306 (N_29306,N_24161,N_24936);
or U29307 (N_29307,N_24976,N_20240);
and U29308 (N_29308,N_21605,N_20812);
or U29309 (N_29309,N_23477,N_23389);
nand U29310 (N_29310,N_22737,N_20265);
nor U29311 (N_29311,N_21364,N_22334);
nand U29312 (N_29312,N_24806,N_22643);
and U29313 (N_29313,N_21007,N_22111);
nand U29314 (N_29314,N_22417,N_24854);
nor U29315 (N_29315,N_20333,N_23458);
or U29316 (N_29316,N_20361,N_23208);
nor U29317 (N_29317,N_21782,N_23630);
nand U29318 (N_29318,N_21062,N_20264);
or U29319 (N_29319,N_22576,N_23873);
or U29320 (N_29320,N_22866,N_20317);
or U29321 (N_29321,N_20118,N_21592);
nor U29322 (N_29322,N_21626,N_20518);
nor U29323 (N_29323,N_21822,N_23012);
nor U29324 (N_29324,N_20645,N_22042);
and U29325 (N_29325,N_21514,N_23633);
nor U29326 (N_29326,N_23082,N_20794);
nand U29327 (N_29327,N_21045,N_24686);
and U29328 (N_29328,N_20968,N_23045);
nor U29329 (N_29329,N_24352,N_20244);
nand U29330 (N_29330,N_24440,N_20112);
or U29331 (N_29331,N_23925,N_22732);
nor U29332 (N_29332,N_22747,N_23511);
nand U29333 (N_29333,N_22682,N_24955);
or U29334 (N_29334,N_22925,N_21219);
nand U29335 (N_29335,N_23537,N_20347);
and U29336 (N_29336,N_23386,N_23968);
nor U29337 (N_29337,N_21954,N_22823);
and U29338 (N_29338,N_22285,N_22173);
nand U29339 (N_29339,N_20575,N_23655);
and U29340 (N_29340,N_22628,N_21255);
or U29341 (N_29341,N_20813,N_21381);
nor U29342 (N_29342,N_21072,N_22678);
or U29343 (N_29343,N_20808,N_23533);
nand U29344 (N_29344,N_20078,N_22897);
xnor U29345 (N_29345,N_22607,N_23110);
or U29346 (N_29346,N_22183,N_21775);
and U29347 (N_29347,N_24316,N_22246);
nand U29348 (N_29348,N_20864,N_20088);
or U29349 (N_29349,N_20262,N_21523);
or U29350 (N_29350,N_24785,N_20871);
nor U29351 (N_29351,N_22549,N_21881);
xor U29352 (N_29352,N_21088,N_23646);
nand U29353 (N_29353,N_24075,N_24983);
and U29354 (N_29354,N_22260,N_23723);
and U29355 (N_29355,N_24944,N_24330);
nor U29356 (N_29356,N_21571,N_21834);
nor U29357 (N_29357,N_24400,N_23851);
nor U29358 (N_29358,N_23597,N_23262);
and U29359 (N_29359,N_22086,N_20115);
and U29360 (N_29360,N_23584,N_22770);
and U29361 (N_29361,N_20400,N_20686);
nor U29362 (N_29362,N_21682,N_21955);
nor U29363 (N_29363,N_20966,N_24072);
or U29364 (N_29364,N_23084,N_21959);
or U29365 (N_29365,N_23408,N_20173);
nand U29366 (N_29366,N_20280,N_24376);
nor U29367 (N_29367,N_21825,N_23591);
and U29368 (N_29368,N_22677,N_22817);
and U29369 (N_29369,N_20953,N_20779);
nor U29370 (N_29370,N_24253,N_22998);
nor U29371 (N_29371,N_23851,N_20246);
or U29372 (N_29372,N_22431,N_24181);
and U29373 (N_29373,N_22299,N_24481);
or U29374 (N_29374,N_21343,N_20640);
nand U29375 (N_29375,N_21056,N_22911);
or U29376 (N_29376,N_21806,N_22621);
and U29377 (N_29377,N_23946,N_21208);
xor U29378 (N_29378,N_24333,N_21214);
nand U29379 (N_29379,N_23449,N_21448);
nor U29380 (N_29380,N_21119,N_24602);
and U29381 (N_29381,N_21058,N_20960);
or U29382 (N_29382,N_23221,N_22005);
xnor U29383 (N_29383,N_24111,N_22646);
or U29384 (N_29384,N_21617,N_23707);
and U29385 (N_29385,N_22141,N_21915);
or U29386 (N_29386,N_24749,N_22629);
nand U29387 (N_29387,N_22355,N_24389);
nor U29388 (N_29388,N_24704,N_23832);
nand U29389 (N_29389,N_21442,N_24793);
and U29390 (N_29390,N_21010,N_22098);
or U29391 (N_29391,N_22581,N_20956);
nor U29392 (N_29392,N_24880,N_21353);
and U29393 (N_29393,N_22200,N_22241);
and U29394 (N_29394,N_23233,N_20208);
and U29395 (N_29395,N_23741,N_22359);
nand U29396 (N_29396,N_23171,N_22821);
nor U29397 (N_29397,N_23633,N_20773);
nand U29398 (N_29398,N_20492,N_21692);
or U29399 (N_29399,N_24110,N_24112);
nor U29400 (N_29400,N_22020,N_21096);
or U29401 (N_29401,N_24561,N_21031);
or U29402 (N_29402,N_24189,N_22131);
xnor U29403 (N_29403,N_21293,N_20278);
and U29404 (N_29404,N_24222,N_20058);
nand U29405 (N_29405,N_24552,N_21234);
or U29406 (N_29406,N_24357,N_24253);
or U29407 (N_29407,N_21622,N_20554);
nand U29408 (N_29408,N_21563,N_24575);
or U29409 (N_29409,N_20782,N_20628);
nor U29410 (N_29410,N_23307,N_22194);
nor U29411 (N_29411,N_22919,N_23215);
or U29412 (N_29412,N_20896,N_22560);
or U29413 (N_29413,N_22577,N_21420);
and U29414 (N_29414,N_20362,N_24138);
nand U29415 (N_29415,N_21300,N_21371);
or U29416 (N_29416,N_20540,N_21593);
xor U29417 (N_29417,N_23704,N_24400);
or U29418 (N_29418,N_23514,N_20851);
xnor U29419 (N_29419,N_20672,N_21037);
or U29420 (N_29420,N_23386,N_21853);
nor U29421 (N_29421,N_22378,N_23833);
or U29422 (N_29422,N_22977,N_21245);
xnor U29423 (N_29423,N_22117,N_24280);
or U29424 (N_29424,N_23209,N_24397);
xnor U29425 (N_29425,N_20468,N_23209);
or U29426 (N_29426,N_23339,N_21624);
nand U29427 (N_29427,N_23211,N_21305);
xnor U29428 (N_29428,N_22708,N_23835);
or U29429 (N_29429,N_23178,N_23049);
or U29430 (N_29430,N_24253,N_21321);
and U29431 (N_29431,N_20703,N_22991);
nor U29432 (N_29432,N_22213,N_23449);
nand U29433 (N_29433,N_23392,N_23766);
or U29434 (N_29434,N_24804,N_24442);
or U29435 (N_29435,N_22786,N_21190);
nor U29436 (N_29436,N_21686,N_24710);
or U29437 (N_29437,N_24460,N_24584);
or U29438 (N_29438,N_20596,N_24956);
or U29439 (N_29439,N_20233,N_20722);
nor U29440 (N_29440,N_20230,N_21451);
nor U29441 (N_29441,N_22242,N_24753);
or U29442 (N_29442,N_24885,N_23443);
xnor U29443 (N_29443,N_20757,N_20168);
nor U29444 (N_29444,N_23452,N_24881);
xor U29445 (N_29445,N_24991,N_21865);
nand U29446 (N_29446,N_21801,N_22476);
nand U29447 (N_29447,N_20755,N_22942);
nor U29448 (N_29448,N_21952,N_22459);
nor U29449 (N_29449,N_21468,N_20368);
or U29450 (N_29450,N_20900,N_20151);
nor U29451 (N_29451,N_24770,N_23962);
xnor U29452 (N_29452,N_23388,N_24652);
or U29453 (N_29453,N_20937,N_21949);
and U29454 (N_29454,N_21844,N_20480);
or U29455 (N_29455,N_23642,N_23470);
xor U29456 (N_29456,N_22699,N_21003);
nor U29457 (N_29457,N_22521,N_21394);
and U29458 (N_29458,N_23311,N_20540);
nand U29459 (N_29459,N_21627,N_21912);
and U29460 (N_29460,N_21998,N_20506);
and U29461 (N_29461,N_23981,N_21327);
and U29462 (N_29462,N_23848,N_20887);
and U29463 (N_29463,N_24582,N_24448);
and U29464 (N_29464,N_20418,N_23695);
nand U29465 (N_29465,N_23002,N_21177);
and U29466 (N_29466,N_24192,N_23412);
nor U29467 (N_29467,N_24504,N_23226);
and U29468 (N_29468,N_23106,N_21857);
or U29469 (N_29469,N_21372,N_20669);
nand U29470 (N_29470,N_24834,N_21588);
xnor U29471 (N_29471,N_20548,N_24064);
nor U29472 (N_29472,N_24512,N_21622);
nand U29473 (N_29473,N_21807,N_21756);
nand U29474 (N_29474,N_20570,N_22812);
and U29475 (N_29475,N_20293,N_22092);
and U29476 (N_29476,N_21401,N_23102);
nand U29477 (N_29477,N_24468,N_23367);
nor U29478 (N_29478,N_20492,N_21315);
nor U29479 (N_29479,N_24108,N_24966);
nor U29480 (N_29480,N_22311,N_20773);
nand U29481 (N_29481,N_23673,N_22747);
and U29482 (N_29482,N_24963,N_23640);
nor U29483 (N_29483,N_21240,N_24209);
nor U29484 (N_29484,N_21330,N_21631);
nand U29485 (N_29485,N_24975,N_20848);
nor U29486 (N_29486,N_20628,N_23348);
nor U29487 (N_29487,N_22706,N_21870);
or U29488 (N_29488,N_21571,N_20818);
nand U29489 (N_29489,N_20587,N_21468);
and U29490 (N_29490,N_20033,N_21357);
nand U29491 (N_29491,N_23290,N_24758);
nand U29492 (N_29492,N_21361,N_21520);
and U29493 (N_29493,N_24486,N_22004);
nor U29494 (N_29494,N_20269,N_20272);
and U29495 (N_29495,N_24243,N_21617);
nand U29496 (N_29496,N_24320,N_20004);
nand U29497 (N_29497,N_23465,N_21867);
or U29498 (N_29498,N_21811,N_23566);
or U29499 (N_29499,N_21252,N_24984);
nor U29500 (N_29500,N_21691,N_21024);
nand U29501 (N_29501,N_24186,N_22890);
nor U29502 (N_29502,N_24889,N_22230);
nor U29503 (N_29503,N_24110,N_21266);
nand U29504 (N_29504,N_23587,N_20308);
nor U29505 (N_29505,N_23882,N_20635);
or U29506 (N_29506,N_24937,N_22474);
and U29507 (N_29507,N_23006,N_21565);
nand U29508 (N_29508,N_22937,N_21651);
nor U29509 (N_29509,N_24279,N_21070);
nor U29510 (N_29510,N_24511,N_20382);
and U29511 (N_29511,N_20731,N_20236);
nand U29512 (N_29512,N_22509,N_21110);
or U29513 (N_29513,N_22895,N_22698);
or U29514 (N_29514,N_23208,N_24507);
nand U29515 (N_29515,N_21718,N_22777);
or U29516 (N_29516,N_24966,N_21266);
nor U29517 (N_29517,N_21364,N_21715);
nor U29518 (N_29518,N_21875,N_20852);
or U29519 (N_29519,N_20288,N_21025);
and U29520 (N_29520,N_23126,N_23406);
nand U29521 (N_29521,N_24318,N_22318);
xor U29522 (N_29522,N_23272,N_23128);
nor U29523 (N_29523,N_22523,N_23366);
or U29524 (N_29524,N_23978,N_20341);
nand U29525 (N_29525,N_20301,N_20165);
and U29526 (N_29526,N_20767,N_21090);
or U29527 (N_29527,N_22827,N_23508);
or U29528 (N_29528,N_24536,N_24961);
or U29529 (N_29529,N_20848,N_21694);
or U29530 (N_29530,N_24922,N_22896);
nand U29531 (N_29531,N_24728,N_23104);
nand U29532 (N_29532,N_24313,N_24681);
nand U29533 (N_29533,N_24849,N_21901);
nor U29534 (N_29534,N_20686,N_22601);
nor U29535 (N_29535,N_20160,N_21453);
nand U29536 (N_29536,N_21976,N_22195);
or U29537 (N_29537,N_24833,N_24991);
nor U29538 (N_29538,N_24539,N_22558);
nand U29539 (N_29539,N_22713,N_20560);
and U29540 (N_29540,N_22129,N_21736);
xor U29541 (N_29541,N_23799,N_21111);
nor U29542 (N_29542,N_23263,N_24330);
nand U29543 (N_29543,N_24255,N_24825);
or U29544 (N_29544,N_20541,N_20295);
nand U29545 (N_29545,N_20896,N_20048);
or U29546 (N_29546,N_21062,N_20954);
xnor U29547 (N_29547,N_24621,N_21920);
or U29548 (N_29548,N_24396,N_22064);
nand U29549 (N_29549,N_21612,N_20783);
nor U29550 (N_29550,N_20387,N_22521);
xor U29551 (N_29551,N_22402,N_23689);
nand U29552 (N_29552,N_23170,N_20379);
or U29553 (N_29553,N_21650,N_24370);
nand U29554 (N_29554,N_20531,N_24176);
nand U29555 (N_29555,N_20763,N_22343);
nor U29556 (N_29556,N_23610,N_23130);
or U29557 (N_29557,N_21239,N_24501);
and U29558 (N_29558,N_20448,N_21060);
xor U29559 (N_29559,N_24977,N_21883);
nor U29560 (N_29560,N_21788,N_22787);
nand U29561 (N_29561,N_23346,N_20090);
or U29562 (N_29562,N_24815,N_20218);
and U29563 (N_29563,N_24717,N_24704);
nand U29564 (N_29564,N_21244,N_24770);
xnor U29565 (N_29565,N_23858,N_24398);
or U29566 (N_29566,N_24922,N_24195);
and U29567 (N_29567,N_23242,N_21338);
and U29568 (N_29568,N_22096,N_22910);
or U29569 (N_29569,N_22672,N_24171);
xnor U29570 (N_29570,N_21669,N_21012);
nor U29571 (N_29571,N_24901,N_24337);
nor U29572 (N_29572,N_24191,N_22173);
nand U29573 (N_29573,N_23905,N_22751);
or U29574 (N_29574,N_22791,N_24051);
and U29575 (N_29575,N_22790,N_23119);
nand U29576 (N_29576,N_20700,N_22429);
nor U29577 (N_29577,N_24179,N_22302);
or U29578 (N_29578,N_21542,N_20324);
nor U29579 (N_29579,N_24129,N_22113);
or U29580 (N_29580,N_24089,N_21769);
and U29581 (N_29581,N_20878,N_21869);
nor U29582 (N_29582,N_24056,N_20232);
and U29583 (N_29583,N_23800,N_22853);
and U29584 (N_29584,N_24636,N_23312);
or U29585 (N_29585,N_22385,N_23364);
nor U29586 (N_29586,N_23278,N_23620);
nor U29587 (N_29587,N_22698,N_24585);
nand U29588 (N_29588,N_20327,N_24913);
or U29589 (N_29589,N_21654,N_20828);
nor U29590 (N_29590,N_21858,N_21017);
or U29591 (N_29591,N_23297,N_21316);
or U29592 (N_29592,N_24620,N_24941);
xor U29593 (N_29593,N_23587,N_23089);
or U29594 (N_29594,N_23487,N_24914);
and U29595 (N_29595,N_21437,N_20484);
or U29596 (N_29596,N_20706,N_20113);
xor U29597 (N_29597,N_22521,N_24413);
or U29598 (N_29598,N_23764,N_20636);
nor U29599 (N_29599,N_21820,N_24390);
xnor U29600 (N_29600,N_24100,N_20386);
nor U29601 (N_29601,N_23553,N_24198);
nor U29602 (N_29602,N_23337,N_24859);
and U29603 (N_29603,N_22109,N_24618);
and U29604 (N_29604,N_20963,N_20817);
nand U29605 (N_29605,N_21204,N_21691);
or U29606 (N_29606,N_20450,N_22599);
or U29607 (N_29607,N_20326,N_21840);
and U29608 (N_29608,N_20213,N_22186);
nor U29609 (N_29609,N_23554,N_22994);
nor U29610 (N_29610,N_24874,N_23694);
nor U29611 (N_29611,N_20024,N_24313);
nand U29612 (N_29612,N_20704,N_22466);
and U29613 (N_29613,N_24359,N_23243);
or U29614 (N_29614,N_20593,N_21075);
and U29615 (N_29615,N_20253,N_24851);
and U29616 (N_29616,N_20869,N_21416);
nor U29617 (N_29617,N_20129,N_23498);
or U29618 (N_29618,N_20379,N_22397);
or U29619 (N_29619,N_24204,N_23406);
nand U29620 (N_29620,N_23151,N_21663);
nor U29621 (N_29621,N_22189,N_21534);
nor U29622 (N_29622,N_24495,N_23836);
and U29623 (N_29623,N_22451,N_24070);
or U29624 (N_29624,N_22036,N_24273);
nor U29625 (N_29625,N_20867,N_22146);
and U29626 (N_29626,N_24851,N_23108);
nor U29627 (N_29627,N_23729,N_21483);
nor U29628 (N_29628,N_23962,N_24738);
nor U29629 (N_29629,N_20528,N_20841);
nand U29630 (N_29630,N_23827,N_22286);
xnor U29631 (N_29631,N_23347,N_20788);
nor U29632 (N_29632,N_23859,N_20011);
nand U29633 (N_29633,N_22475,N_22556);
nand U29634 (N_29634,N_23207,N_21734);
nor U29635 (N_29635,N_21314,N_20164);
nand U29636 (N_29636,N_24425,N_21525);
or U29637 (N_29637,N_21530,N_22425);
nor U29638 (N_29638,N_20703,N_20617);
or U29639 (N_29639,N_22218,N_23160);
xor U29640 (N_29640,N_20094,N_21410);
or U29641 (N_29641,N_22300,N_23572);
nor U29642 (N_29642,N_20481,N_22358);
nor U29643 (N_29643,N_23302,N_23256);
nor U29644 (N_29644,N_21557,N_23793);
xnor U29645 (N_29645,N_21467,N_20662);
or U29646 (N_29646,N_24868,N_21936);
xor U29647 (N_29647,N_20333,N_24267);
nand U29648 (N_29648,N_20399,N_20382);
nand U29649 (N_29649,N_21248,N_23243);
or U29650 (N_29650,N_21496,N_21280);
nor U29651 (N_29651,N_23742,N_24632);
and U29652 (N_29652,N_24911,N_23259);
and U29653 (N_29653,N_21305,N_24860);
and U29654 (N_29654,N_20107,N_23118);
and U29655 (N_29655,N_22480,N_22572);
or U29656 (N_29656,N_23734,N_20035);
xor U29657 (N_29657,N_23004,N_23209);
and U29658 (N_29658,N_21038,N_24641);
or U29659 (N_29659,N_23981,N_21165);
nor U29660 (N_29660,N_24247,N_20860);
and U29661 (N_29661,N_21788,N_22850);
xor U29662 (N_29662,N_24040,N_20673);
and U29663 (N_29663,N_21813,N_23169);
nand U29664 (N_29664,N_22949,N_23660);
and U29665 (N_29665,N_24535,N_24262);
nand U29666 (N_29666,N_22621,N_21445);
nor U29667 (N_29667,N_24593,N_22859);
nor U29668 (N_29668,N_21528,N_20165);
nor U29669 (N_29669,N_21248,N_22831);
or U29670 (N_29670,N_23495,N_24760);
xor U29671 (N_29671,N_23924,N_23124);
nor U29672 (N_29672,N_23472,N_24055);
and U29673 (N_29673,N_23143,N_21912);
and U29674 (N_29674,N_21792,N_20286);
or U29675 (N_29675,N_24395,N_23228);
or U29676 (N_29676,N_24177,N_23837);
nand U29677 (N_29677,N_23085,N_23918);
and U29678 (N_29678,N_22859,N_22398);
or U29679 (N_29679,N_20904,N_21876);
and U29680 (N_29680,N_22239,N_23944);
nand U29681 (N_29681,N_23926,N_22281);
xor U29682 (N_29682,N_24097,N_21799);
xnor U29683 (N_29683,N_20212,N_21350);
nor U29684 (N_29684,N_21395,N_21766);
nand U29685 (N_29685,N_21474,N_21145);
nand U29686 (N_29686,N_20112,N_20339);
nor U29687 (N_29687,N_24591,N_24354);
nor U29688 (N_29688,N_20303,N_20886);
nand U29689 (N_29689,N_21765,N_20616);
nand U29690 (N_29690,N_20774,N_24959);
nor U29691 (N_29691,N_20601,N_22710);
and U29692 (N_29692,N_22647,N_20474);
nor U29693 (N_29693,N_20796,N_21603);
and U29694 (N_29694,N_24282,N_20265);
nand U29695 (N_29695,N_22857,N_22205);
nand U29696 (N_29696,N_21694,N_24062);
nor U29697 (N_29697,N_22750,N_20514);
nand U29698 (N_29698,N_20246,N_24701);
or U29699 (N_29699,N_22205,N_23398);
or U29700 (N_29700,N_22369,N_20860);
nand U29701 (N_29701,N_21589,N_22498);
or U29702 (N_29702,N_20340,N_24968);
nand U29703 (N_29703,N_24062,N_20112);
nand U29704 (N_29704,N_23726,N_20742);
xor U29705 (N_29705,N_21843,N_24462);
nor U29706 (N_29706,N_24861,N_21395);
and U29707 (N_29707,N_21471,N_20536);
nand U29708 (N_29708,N_23867,N_21313);
or U29709 (N_29709,N_24012,N_23144);
nand U29710 (N_29710,N_21168,N_21086);
nor U29711 (N_29711,N_22749,N_22062);
nand U29712 (N_29712,N_21926,N_21954);
and U29713 (N_29713,N_23418,N_23714);
and U29714 (N_29714,N_21838,N_24924);
and U29715 (N_29715,N_23081,N_21432);
or U29716 (N_29716,N_22071,N_24347);
and U29717 (N_29717,N_20559,N_20963);
nand U29718 (N_29718,N_20713,N_22523);
nand U29719 (N_29719,N_21861,N_22152);
and U29720 (N_29720,N_23314,N_22101);
or U29721 (N_29721,N_23347,N_21464);
nor U29722 (N_29722,N_20448,N_20479);
and U29723 (N_29723,N_22993,N_22677);
and U29724 (N_29724,N_22865,N_24483);
nor U29725 (N_29725,N_20614,N_21295);
and U29726 (N_29726,N_24651,N_21698);
nand U29727 (N_29727,N_20523,N_24040);
nor U29728 (N_29728,N_20124,N_23748);
or U29729 (N_29729,N_23491,N_24083);
nand U29730 (N_29730,N_21063,N_22201);
xnor U29731 (N_29731,N_20220,N_20145);
nor U29732 (N_29732,N_20358,N_22879);
xor U29733 (N_29733,N_24991,N_23721);
nand U29734 (N_29734,N_22287,N_21028);
nand U29735 (N_29735,N_21353,N_24926);
xnor U29736 (N_29736,N_21504,N_22365);
or U29737 (N_29737,N_22379,N_20144);
or U29738 (N_29738,N_23687,N_21336);
and U29739 (N_29739,N_22453,N_20910);
nor U29740 (N_29740,N_22271,N_20626);
or U29741 (N_29741,N_23358,N_24652);
nor U29742 (N_29742,N_21126,N_23912);
xnor U29743 (N_29743,N_24625,N_21710);
nand U29744 (N_29744,N_21355,N_21333);
nand U29745 (N_29745,N_23799,N_20323);
and U29746 (N_29746,N_20761,N_24039);
nor U29747 (N_29747,N_23267,N_23759);
nor U29748 (N_29748,N_23856,N_21181);
xnor U29749 (N_29749,N_20197,N_22225);
and U29750 (N_29750,N_20137,N_20118);
xnor U29751 (N_29751,N_22922,N_21442);
and U29752 (N_29752,N_22273,N_21666);
or U29753 (N_29753,N_20194,N_22605);
and U29754 (N_29754,N_20775,N_21756);
and U29755 (N_29755,N_20690,N_24325);
nand U29756 (N_29756,N_24995,N_22926);
and U29757 (N_29757,N_20166,N_23258);
nand U29758 (N_29758,N_24067,N_22610);
nand U29759 (N_29759,N_24719,N_23872);
nand U29760 (N_29760,N_20316,N_20648);
and U29761 (N_29761,N_20072,N_22352);
nand U29762 (N_29762,N_22446,N_22654);
and U29763 (N_29763,N_24937,N_23843);
xnor U29764 (N_29764,N_22615,N_23819);
nor U29765 (N_29765,N_23878,N_21423);
nor U29766 (N_29766,N_21585,N_22195);
nand U29767 (N_29767,N_22318,N_24211);
nor U29768 (N_29768,N_23302,N_23100);
nor U29769 (N_29769,N_22698,N_24784);
nor U29770 (N_29770,N_21070,N_20679);
and U29771 (N_29771,N_23279,N_22874);
nand U29772 (N_29772,N_21132,N_23378);
nor U29773 (N_29773,N_23726,N_21565);
nand U29774 (N_29774,N_20859,N_24819);
nand U29775 (N_29775,N_22940,N_21581);
or U29776 (N_29776,N_20759,N_24952);
nand U29777 (N_29777,N_20673,N_22650);
nand U29778 (N_29778,N_21717,N_21710);
and U29779 (N_29779,N_21094,N_20736);
nor U29780 (N_29780,N_24927,N_20702);
nand U29781 (N_29781,N_23603,N_24267);
nand U29782 (N_29782,N_24179,N_22963);
nor U29783 (N_29783,N_21425,N_20312);
xor U29784 (N_29784,N_22623,N_24598);
or U29785 (N_29785,N_23964,N_20913);
and U29786 (N_29786,N_22205,N_21899);
nand U29787 (N_29787,N_24176,N_23775);
nand U29788 (N_29788,N_22853,N_20670);
nand U29789 (N_29789,N_20646,N_23653);
or U29790 (N_29790,N_23222,N_20292);
and U29791 (N_29791,N_24706,N_23669);
xnor U29792 (N_29792,N_24450,N_22707);
or U29793 (N_29793,N_20983,N_22763);
or U29794 (N_29794,N_20397,N_20593);
and U29795 (N_29795,N_22244,N_20223);
nand U29796 (N_29796,N_20919,N_22731);
or U29797 (N_29797,N_21911,N_22479);
and U29798 (N_29798,N_24335,N_22979);
nor U29799 (N_29799,N_24425,N_21578);
xnor U29800 (N_29800,N_20754,N_24067);
and U29801 (N_29801,N_20536,N_23357);
or U29802 (N_29802,N_20129,N_24812);
or U29803 (N_29803,N_22976,N_23266);
nor U29804 (N_29804,N_21674,N_20144);
nand U29805 (N_29805,N_23872,N_20647);
nand U29806 (N_29806,N_24418,N_23318);
or U29807 (N_29807,N_23696,N_21588);
or U29808 (N_29808,N_24901,N_23035);
nor U29809 (N_29809,N_22790,N_22181);
xnor U29810 (N_29810,N_20434,N_21872);
nand U29811 (N_29811,N_23136,N_21358);
nor U29812 (N_29812,N_24960,N_24422);
or U29813 (N_29813,N_23922,N_23830);
nor U29814 (N_29814,N_21764,N_23259);
nand U29815 (N_29815,N_24076,N_20272);
nor U29816 (N_29816,N_21955,N_23597);
xor U29817 (N_29817,N_23950,N_22942);
nand U29818 (N_29818,N_22826,N_24331);
nor U29819 (N_29819,N_23546,N_24902);
nand U29820 (N_29820,N_22876,N_20025);
and U29821 (N_29821,N_24401,N_23534);
xnor U29822 (N_29822,N_21804,N_20306);
or U29823 (N_29823,N_24117,N_23634);
and U29824 (N_29824,N_22809,N_22983);
xnor U29825 (N_29825,N_20782,N_23492);
nor U29826 (N_29826,N_20142,N_24568);
or U29827 (N_29827,N_23298,N_23264);
nand U29828 (N_29828,N_21710,N_23374);
xor U29829 (N_29829,N_23079,N_22691);
nor U29830 (N_29830,N_20028,N_21069);
and U29831 (N_29831,N_23749,N_24927);
nor U29832 (N_29832,N_20993,N_24607);
or U29833 (N_29833,N_20232,N_21784);
nand U29834 (N_29834,N_21932,N_21533);
or U29835 (N_29835,N_22349,N_22528);
and U29836 (N_29836,N_20498,N_24123);
and U29837 (N_29837,N_24402,N_23579);
nand U29838 (N_29838,N_21889,N_24407);
xor U29839 (N_29839,N_22458,N_22547);
nand U29840 (N_29840,N_20538,N_21877);
nor U29841 (N_29841,N_24418,N_20263);
and U29842 (N_29842,N_23527,N_20433);
nand U29843 (N_29843,N_22164,N_20618);
nor U29844 (N_29844,N_22913,N_23247);
nor U29845 (N_29845,N_24936,N_22300);
xor U29846 (N_29846,N_23268,N_24488);
nand U29847 (N_29847,N_22894,N_23698);
or U29848 (N_29848,N_24971,N_20220);
or U29849 (N_29849,N_20705,N_23432);
nand U29850 (N_29850,N_22275,N_24366);
or U29851 (N_29851,N_24679,N_24569);
nand U29852 (N_29852,N_20317,N_23005);
and U29853 (N_29853,N_23617,N_21682);
and U29854 (N_29854,N_23893,N_23661);
or U29855 (N_29855,N_24802,N_22875);
or U29856 (N_29856,N_21616,N_24753);
nand U29857 (N_29857,N_23744,N_20183);
nor U29858 (N_29858,N_20419,N_23933);
xnor U29859 (N_29859,N_23977,N_20358);
xor U29860 (N_29860,N_22626,N_20999);
nand U29861 (N_29861,N_22322,N_24531);
or U29862 (N_29862,N_24288,N_22633);
and U29863 (N_29863,N_22697,N_24353);
and U29864 (N_29864,N_22549,N_21665);
nand U29865 (N_29865,N_24008,N_20165);
or U29866 (N_29866,N_21122,N_21481);
nand U29867 (N_29867,N_22706,N_23015);
nor U29868 (N_29868,N_21042,N_24922);
or U29869 (N_29869,N_21981,N_20838);
nor U29870 (N_29870,N_22822,N_23791);
or U29871 (N_29871,N_22424,N_22844);
or U29872 (N_29872,N_22505,N_22211);
or U29873 (N_29873,N_22743,N_21050);
nor U29874 (N_29874,N_23284,N_23675);
and U29875 (N_29875,N_21121,N_20846);
nor U29876 (N_29876,N_23047,N_22272);
nor U29877 (N_29877,N_23995,N_21024);
and U29878 (N_29878,N_24180,N_22543);
xor U29879 (N_29879,N_22467,N_21174);
xnor U29880 (N_29880,N_20909,N_21964);
nor U29881 (N_29881,N_23060,N_20302);
nor U29882 (N_29882,N_20073,N_23787);
and U29883 (N_29883,N_23614,N_24967);
and U29884 (N_29884,N_23259,N_20137);
or U29885 (N_29885,N_24951,N_21483);
nor U29886 (N_29886,N_20158,N_20935);
and U29887 (N_29887,N_24652,N_22910);
or U29888 (N_29888,N_24932,N_22596);
nor U29889 (N_29889,N_24212,N_22380);
and U29890 (N_29890,N_24227,N_21293);
and U29891 (N_29891,N_22646,N_22663);
or U29892 (N_29892,N_20595,N_23112);
nand U29893 (N_29893,N_22427,N_20493);
nand U29894 (N_29894,N_20085,N_21788);
nor U29895 (N_29895,N_20405,N_22036);
or U29896 (N_29896,N_22996,N_21697);
nor U29897 (N_29897,N_21778,N_24059);
nor U29898 (N_29898,N_24007,N_22354);
xnor U29899 (N_29899,N_22290,N_23339);
nand U29900 (N_29900,N_23228,N_23182);
or U29901 (N_29901,N_22744,N_23261);
nand U29902 (N_29902,N_21783,N_22372);
and U29903 (N_29903,N_22042,N_22822);
xor U29904 (N_29904,N_22703,N_22017);
and U29905 (N_29905,N_23846,N_21206);
nor U29906 (N_29906,N_23036,N_22461);
nand U29907 (N_29907,N_21034,N_20625);
nand U29908 (N_29908,N_23658,N_24244);
and U29909 (N_29909,N_23364,N_21187);
or U29910 (N_29910,N_23303,N_21856);
and U29911 (N_29911,N_21327,N_24280);
and U29912 (N_29912,N_20398,N_21246);
xnor U29913 (N_29913,N_23857,N_20382);
nor U29914 (N_29914,N_23601,N_24639);
and U29915 (N_29915,N_21582,N_22238);
and U29916 (N_29916,N_20816,N_22140);
nor U29917 (N_29917,N_24003,N_21721);
and U29918 (N_29918,N_22111,N_20090);
xnor U29919 (N_29919,N_22541,N_20622);
nand U29920 (N_29920,N_23691,N_23582);
and U29921 (N_29921,N_20550,N_24217);
nor U29922 (N_29922,N_21786,N_23811);
nor U29923 (N_29923,N_24385,N_20218);
and U29924 (N_29924,N_21996,N_21707);
nor U29925 (N_29925,N_21172,N_23570);
xor U29926 (N_29926,N_22209,N_23119);
nand U29927 (N_29927,N_23481,N_20024);
nor U29928 (N_29928,N_21914,N_20128);
or U29929 (N_29929,N_21849,N_23854);
nand U29930 (N_29930,N_21317,N_20981);
and U29931 (N_29931,N_23482,N_22697);
nor U29932 (N_29932,N_20451,N_24526);
nor U29933 (N_29933,N_23796,N_23458);
nor U29934 (N_29934,N_22116,N_24719);
xnor U29935 (N_29935,N_24389,N_20981);
nor U29936 (N_29936,N_21037,N_24212);
xnor U29937 (N_29937,N_22759,N_24365);
or U29938 (N_29938,N_22772,N_23713);
nand U29939 (N_29939,N_23536,N_21628);
and U29940 (N_29940,N_23319,N_21468);
nor U29941 (N_29941,N_22287,N_20223);
and U29942 (N_29942,N_20597,N_20421);
and U29943 (N_29943,N_22274,N_22634);
and U29944 (N_29944,N_24578,N_23815);
nor U29945 (N_29945,N_22381,N_22316);
nand U29946 (N_29946,N_21220,N_22545);
nand U29947 (N_29947,N_23158,N_21057);
nor U29948 (N_29948,N_24837,N_24206);
or U29949 (N_29949,N_22130,N_21375);
nand U29950 (N_29950,N_23498,N_21795);
or U29951 (N_29951,N_23221,N_21734);
nor U29952 (N_29952,N_20488,N_22439);
nand U29953 (N_29953,N_22607,N_23381);
nand U29954 (N_29954,N_21281,N_24492);
xnor U29955 (N_29955,N_21283,N_22053);
and U29956 (N_29956,N_21460,N_20012);
nor U29957 (N_29957,N_21698,N_23923);
nand U29958 (N_29958,N_22931,N_24926);
or U29959 (N_29959,N_24504,N_22611);
nand U29960 (N_29960,N_24249,N_20236);
or U29961 (N_29961,N_23716,N_24651);
and U29962 (N_29962,N_22621,N_22093);
or U29963 (N_29963,N_24670,N_21182);
and U29964 (N_29964,N_23380,N_23080);
and U29965 (N_29965,N_23365,N_22011);
or U29966 (N_29966,N_23677,N_23126);
nor U29967 (N_29967,N_22062,N_20890);
and U29968 (N_29968,N_24545,N_20871);
nand U29969 (N_29969,N_22089,N_20944);
nand U29970 (N_29970,N_20325,N_22280);
nand U29971 (N_29971,N_23045,N_20746);
nand U29972 (N_29972,N_20317,N_22136);
nor U29973 (N_29973,N_20397,N_23383);
xnor U29974 (N_29974,N_23849,N_21407);
nor U29975 (N_29975,N_20836,N_21631);
xnor U29976 (N_29976,N_23177,N_21901);
nand U29977 (N_29977,N_22511,N_24543);
nor U29978 (N_29978,N_20924,N_20171);
nand U29979 (N_29979,N_21997,N_24710);
or U29980 (N_29980,N_20603,N_23191);
or U29981 (N_29981,N_24049,N_21405);
and U29982 (N_29982,N_21783,N_21584);
and U29983 (N_29983,N_23590,N_20668);
xor U29984 (N_29984,N_21944,N_24482);
nand U29985 (N_29985,N_23008,N_21218);
nor U29986 (N_29986,N_21841,N_22985);
and U29987 (N_29987,N_20651,N_23057);
nand U29988 (N_29988,N_23174,N_23490);
nand U29989 (N_29989,N_20694,N_22756);
xor U29990 (N_29990,N_22982,N_22859);
xnor U29991 (N_29991,N_24500,N_21209);
nor U29992 (N_29992,N_24382,N_22649);
and U29993 (N_29993,N_23488,N_23757);
nand U29994 (N_29994,N_21495,N_23751);
and U29995 (N_29995,N_22961,N_22623);
nor U29996 (N_29996,N_21338,N_22912);
nand U29997 (N_29997,N_24582,N_20125);
or U29998 (N_29998,N_23764,N_21489);
xnor U29999 (N_29999,N_20882,N_21259);
and UO_0 (O_0,N_29847,N_27312);
and UO_1 (O_1,N_25498,N_26851);
and UO_2 (O_2,N_27795,N_26329);
and UO_3 (O_3,N_27623,N_29232);
or UO_4 (O_4,N_25426,N_26543);
nor UO_5 (O_5,N_27401,N_26977);
or UO_6 (O_6,N_28270,N_29124);
nor UO_7 (O_7,N_26043,N_26101);
or UO_8 (O_8,N_26441,N_29323);
nand UO_9 (O_9,N_25326,N_28758);
or UO_10 (O_10,N_27322,N_25155);
nand UO_11 (O_11,N_29955,N_26860);
nor UO_12 (O_12,N_27993,N_29205);
nor UO_13 (O_13,N_26203,N_26169);
nand UO_14 (O_14,N_25462,N_26031);
or UO_15 (O_15,N_26708,N_25022);
nand UO_16 (O_16,N_25555,N_27581);
xnor UO_17 (O_17,N_25605,N_26554);
xor UO_18 (O_18,N_25826,N_25986);
and UO_19 (O_19,N_26471,N_27622);
or UO_20 (O_20,N_29372,N_27550);
xnor UO_21 (O_21,N_27371,N_25355);
xnor UO_22 (O_22,N_27030,N_29929);
and UO_23 (O_23,N_28787,N_29636);
and UO_24 (O_24,N_29255,N_26296);
xor UO_25 (O_25,N_27023,N_28467);
xor UO_26 (O_26,N_29111,N_29374);
nand UO_27 (O_27,N_28286,N_25726);
nand UO_28 (O_28,N_25730,N_26493);
or UO_29 (O_29,N_27725,N_26552);
and UO_30 (O_30,N_28916,N_25580);
nand UO_31 (O_31,N_26350,N_25131);
or UO_32 (O_32,N_26082,N_27280);
and UO_33 (O_33,N_25535,N_28862);
nand UO_34 (O_34,N_28114,N_25338);
nand UO_35 (O_35,N_28069,N_28778);
and UO_36 (O_36,N_28927,N_25375);
and UO_37 (O_37,N_28018,N_27566);
and UO_38 (O_38,N_29197,N_28344);
nor UO_39 (O_39,N_27712,N_29959);
nand UO_40 (O_40,N_27574,N_27285);
or UO_41 (O_41,N_29334,N_25886);
and UO_42 (O_42,N_28715,N_28164);
and UO_43 (O_43,N_27932,N_28724);
xor UO_44 (O_44,N_27181,N_28345);
or UO_45 (O_45,N_29495,N_27502);
and UO_46 (O_46,N_26556,N_29917);
nand UO_47 (O_47,N_29531,N_27422);
or UO_48 (O_48,N_28499,N_29503);
xnor UO_49 (O_49,N_27443,N_29622);
nor UO_50 (O_50,N_25383,N_28054);
nand UO_51 (O_51,N_26728,N_29360);
xnor UO_52 (O_52,N_25269,N_28472);
nor UO_53 (O_53,N_28953,N_28510);
or UO_54 (O_54,N_25560,N_25884);
nand UO_55 (O_55,N_26260,N_28740);
and UO_56 (O_56,N_28731,N_27708);
and UO_57 (O_57,N_28213,N_27817);
nor UO_58 (O_58,N_28530,N_28451);
xor UO_59 (O_59,N_26666,N_27626);
and UO_60 (O_60,N_27888,N_27334);
or UO_61 (O_61,N_25296,N_27608);
or UO_62 (O_62,N_29530,N_25585);
and UO_63 (O_63,N_25740,N_26980);
nor UO_64 (O_64,N_25564,N_26963);
xnor UO_65 (O_65,N_25311,N_25033);
nand UO_66 (O_66,N_29728,N_25302);
nor UO_67 (O_67,N_27904,N_25157);
and UO_68 (O_68,N_25396,N_25569);
nand UO_69 (O_69,N_28151,N_27995);
nand UO_70 (O_70,N_25032,N_26608);
and UO_71 (O_71,N_25662,N_25325);
or UO_72 (O_72,N_25331,N_26369);
nand UO_73 (O_73,N_26995,N_28584);
nor UO_74 (O_74,N_26946,N_26660);
or UO_75 (O_75,N_29156,N_25103);
nand UO_76 (O_76,N_25016,N_29328);
xor UO_77 (O_77,N_29267,N_28420);
and UO_78 (O_78,N_28762,N_28661);
and UO_79 (O_79,N_25360,N_28839);
xor UO_80 (O_80,N_26420,N_29435);
or UO_81 (O_81,N_28232,N_28032);
nor UO_82 (O_82,N_25420,N_29534);
nor UO_83 (O_83,N_27053,N_25076);
xnor UO_84 (O_84,N_28958,N_28921);
or UO_85 (O_85,N_25552,N_25673);
xnor UO_86 (O_86,N_27718,N_26771);
and UO_87 (O_87,N_28131,N_28195);
nand UO_88 (O_88,N_29674,N_26920);
nand UO_89 (O_89,N_29085,N_29220);
or UO_90 (O_90,N_27269,N_27816);
nor UO_91 (O_91,N_27770,N_26242);
and UO_92 (O_92,N_26815,N_26450);
xnor UO_93 (O_93,N_26205,N_25418);
nand UO_94 (O_94,N_28609,N_26249);
or UO_95 (O_95,N_28265,N_28328);
nor UO_96 (O_96,N_29543,N_25688);
xor UO_97 (O_97,N_27548,N_28247);
or UO_98 (O_98,N_28269,N_29906);
xor UO_99 (O_99,N_28261,N_27853);
nand UO_100 (O_100,N_28040,N_29765);
or UO_101 (O_101,N_25994,N_25461);
or UO_102 (O_102,N_26687,N_26872);
and UO_103 (O_103,N_29392,N_28111);
nor UO_104 (O_104,N_28144,N_28375);
or UO_105 (O_105,N_29373,N_27735);
nand UO_106 (O_106,N_25260,N_29501);
nor UO_107 (O_107,N_25822,N_25273);
and UO_108 (O_108,N_25433,N_29966);
or UO_109 (O_109,N_25636,N_25758);
nand UO_110 (O_110,N_25637,N_29285);
and UO_111 (O_111,N_27954,N_27777);
nand UO_112 (O_112,N_27951,N_26558);
nor UO_113 (O_113,N_28325,N_26185);
and UO_114 (O_114,N_26596,N_29427);
and UO_115 (O_115,N_27056,N_26367);
and UO_116 (O_116,N_25698,N_27873);
nor UO_117 (O_117,N_25253,N_27402);
nor UO_118 (O_118,N_27721,N_27674);
or UO_119 (O_119,N_26497,N_26217);
nand UO_120 (O_120,N_25832,N_29398);
and UO_121 (O_121,N_29590,N_28821);
or UO_122 (O_122,N_25322,N_25916);
and UO_123 (O_123,N_27769,N_25339);
nand UO_124 (O_124,N_28105,N_29597);
and UO_125 (O_125,N_29110,N_26459);
and UO_126 (O_126,N_27406,N_26675);
or UO_127 (O_127,N_25149,N_26914);
xnor UO_128 (O_128,N_26679,N_27826);
or UO_129 (O_129,N_27753,N_27155);
nand UO_130 (O_130,N_28448,N_27306);
nor UO_131 (O_131,N_26211,N_28932);
nand UO_132 (O_132,N_28877,N_27169);
nand UO_133 (O_133,N_28129,N_26958);
and UO_134 (O_134,N_27541,N_28575);
and UO_135 (O_135,N_26125,N_29602);
nor UO_136 (O_136,N_26682,N_26491);
nor UO_137 (O_137,N_28760,N_26099);
nand UO_138 (O_138,N_25600,N_26225);
or UO_139 (O_139,N_25573,N_29785);
nand UO_140 (O_140,N_27653,N_29062);
or UO_141 (O_141,N_29594,N_29292);
nor UO_142 (O_142,N_27834,N_29146);
nand UO_143 (O_143,N_29720,N_25723);
nand UO_144 (O_144,N_25438,N_28332);
and UO_145 (O_145,N_28314,N_26723);
xor UO_146 (O_146,N_26346,N_26128);
xor UO_147 (O_147,N_26146,N_25905);
nand UO_148 (O_148,N_27913,N_26653);
and UO_149 (O_149,N_28718,N_29225);
nand UO_150 (O_150,N_27097,N_28602);
and UO_151 (O_151,N_25531,N_26711);
or UO_152 (O_152,N_25490,N_26172);
nor UO_153 (O_153,N_25306,N_28540);
nor UO_154 (O_154,N_28736,N_27824);
nand UO_155 (O_155,N_26956,N_25896);
or UO_156 (O_156,N_26859,N_27166);
xnor UO_157 (O_157,N_26353,N_26607);
or UO_158 (O_158,N_29043,N_27438);
or UO_159 (O_159,N_25778,N_28356);
nand UO_160 (O_160,N_26754,N_27462);
nor UO_161 (O_161,N_25198,N_28555);
nor UO_162 (O_162,N_25393,N_26198);
and UO_163 (O_163,N_29015,N_29248);
or UO_164 (O_164,N_28140,N_27710);
nor UO_165 (O_165,N_28985,N_27969);
nand UO_166 (O_166,N_28145,N_29642);
nand UO_167 (O_167,N_28596,N_27270);
and UO_168 (O_168,N_27185,N_27743);
xnor UO_169 (O_169,N_26718,N_27737);
or UO_170 (O_170,N_29990,N_26566);
nand UO_171 (O_171,N_28469,N_26466);
and UO_172 (O_172,N_29281,N_26009);
xor UO_173 (O_173,N_28662,N_26278);
xnor UO_174 (O_174,N_25912,N_27364);
nor UO_175 (O_175,N_26720,N_27054);
xor UO_176 (O_176,N_27872,N_27950);
nand UO_177 (O_177,N_29224,N_27953);
and UO_178 (O_178,N_27599,N_28371);
nor UO_179 (O_179,N_26981,N_25709);
nor UO_180 (O_180,N_27660,N_26818);
nand UO_181 (O_181,N_26505,N_29660);
xnor UO_182 (O_182,N_28322,N_26953);
and UO_183 (O_183,N_29535,N_25679);
nor UO_184 (O_184,N_29083,N_27144);
xor UO_185 (O_185,N_29241,N_27781);
nor UO_186 (O_186,N_28674,N_28378);
or UO_187 (O_187,N_27271,N_25417);
and UO_188 (O_188,N_26574,N_25368);
nor UO_189 (O_189,N_26620,N_27176);
xnor UO_190 (O_190,N_27890,N_25392);
nor UO_191 (O_191,N_27063,N_26640);
and UO_192 (O_192,N_25116,N_29358);
nor UO_193 (O_193,N_28576,N_25004);
or UO_194 (O_194,N_26819,N_29216);
nor UO_195 (O_195,N_26943,N_26999);
nand UO_196 (O_196,N_27646,N_29128);
nand UO_197 (O_197,N_25722,N_26308);
nand UO_198 (O_198,N_26651,N_29551);
and UO_199 (O_199,N_28041,N_27846);
nor UO_200 (O_200,N_28123,N_25352);
and UO_201 (O_201,N_27374,N_25687);
or UO_202 (O_202,N_29889,N_28682);
or UO_203 (O_203,N_28414,N_26562);
nor UO_204 (O_204,N_26791,N_25348);
and UO_205 (O_205,N_26313,N_26157);
and UO_206 (O_206,N_29382,N_28075);
xnor UO_207 (O_207,N_29206,N_25554);
nand UO_208 (O_208,N_28970,N_26616);
nand UO_209 (O_209,N_26438,N_25411);
nand UO_210 (O_210,N_28687,N_25652);
and UO_211 (O_211,N_29848,N_29724);
xor UO_212 (O_212,N_25397,N_29617);
and UO_213 (O_213,N_26922,N_28854);
nand UO_214 (O_214,N_27908,N_29817);
nor UO_215 (O_215,N_27731,N_26287);
xnor UO_216 (O_216,N_29059,N_28616);
and UO_217 (O_217,N_25812,N_29129);
nand UO_218 (O_218,N_25363,N_28090);
nand UO_219 (O_219,N_25820,N_25448);
nand UO_220 (O_220,N_27507,N_27766);
and UO_221 (O_221,N_29411,N_28125);
nor UO_222 (O_222,N_28719,N_25310);
xor UO_223 (O_223,N_29734,N_27659);
nand UO_224 (O_224,N_29237,N_25772);
nand UO_225 (O_225,N_27936,N_29598);
nand UO_226 (O_226,N_29485,N_29448);
or UO_227 (O_227,N_27874,N_27159);
or UO_228 (O_228,N_25574,N_27642);
or UO_229 (O_229,N_26394,N_29027);
or UO_230 (O_230,N_29486,N_28087);
or UO_231 (O_231,N_25817,N_25145);
and UO_232 (O_232,N_28506,N_28606);
and UO_233 (O_233,N_26811,N_26749);
nor UO_234 (O_234,N_27996,N_29303);
nor UO_235 (O_235,N_27043,N_28016);
or UO_236 (O_236,N_28465,N_26677);
nand UO_237 (O_237,N_27449,N_28360);
nor UO_238 (O_238,N_29175,N_26569);
and UO_239 (O_239,N_25732,N_26453);
and UO_240 (O_240,N_27121,N_26785);
nor UO_241 (O_241,N_29553,N_28203);
and UO_242 (O_242,N_29747,N_28299);
or UO_243 (O_243,N_28341,N_28438);
nor UO_244 (O_244,N_28235,N_26780);
xnor UO_245 (O_245,N_28827,N_28691);
nor UO_246 (O_246,N_27609,N_25347);
xnor UO_247 (O_247,N_25452,N_26865);
nand UO_248 (O_248,N_29091,N_27376);
or UO_249 (O_249,N_29329,N_28436);
nor UO_250 (O_250,N_28374,N_28189);
nand UO_251 (O_251,N_27864,N_29671);
and UO_252 (O_252,N_29465,N_26843);
nand UO_253 (O_253,N_26189,N_25836);
nand UO_254 (O_254,N_26582,N_27394);
nor UO_255 (O_255,N_28968,N_25953);
nor UO_256 (O_256,N_26973,N_27621);
and UO_257 (O_257,N_29322,N_29631);
and UO_258 (O_258,N_27597,N_25431);
nand UO_259 (O_259,N_25281,N_25694);
nor UO_260 (O_260,N_28473,N_27860);
or UO_261 (O_261,N_28194,N_26143);
nor UO_262 (O_262,N_29922,N_27190);
nand UO_263 (O_263,N_27959,N_28914);
nand UO_264 (O_264,N_26764,N_25596);
nor UO_265 (O_265,N_28885,N_25428);
and UO_266 (O_266,N_26145,N_27935);
and UO_267 (O_267,N_28826,N_27758);
xnor UO_268 (O_268,N_29638,N_28882);
nand UO_269 (O_269,N_28831,N_27087);
or UO_270 (O_270,N_28370,N_25171);
nand UO_271 (O_271,N_29314,N_27511);
and UO_272 (O_272,N_26700,N_27984);
nand UO_273 (O_273,N_28033,N_28775);
xor UO_274 (O_274,N_29673,N_29996);
xnor UO_275 (O_275,N_26656,N_25685);
and UO_276 (O_276,N_26040,N_29182);
nor UO_277 (O_277,N_29291,N_26545);
xor UO_278 (O_278,N_26159,N_29344);
or UO_279 (O_279,N_29945,N_25266);
nand UO_280 (O_280,N_25805,N_26229);
nand UO_281 (O_281,N_29440,N_25388);
nor UO_282 (O_282,N_25249,N_26557);
nor UO_283 (O_283,N_25774,N_29058);
nand UO_284 (O_284,N_26023,N_27052);
and UO_285 (O_285,N_28899,N_29130);
or UO_286 (O_286,N_28770,N_28879);
or UO_287 (O_287,N_27172,N_29213);
nor UO_288 (O_288,N_29429,N_29540);
nand UO_289 (O_289,N_28729,N_26488);
nor UO_290 (O_290,N_26489,N_27474);
nor UO_291 (O_291,N_26520,N_27578);
nand UO_292 (O_292,N_28912,N_25749);
or UO_293 (O_293,N_29188,N_28909);
and UO_294 (O_294,N_28065,N_29227);
and UO_295 (O_295,N_25903,N_26743);
or UO_296 (O_296,N_25707,N_29295);
nor UO_297 (O_297,N_27384,N_25752);
or UO_298 (O_298,N_28700,N_27093);
or UO_299 (O_299,N_26611,N_28329);
nor UO_300 (O_300,N_26934,N_28005);
and UO_301 (O_301,N_29093,N_29259);
or UO_302 (O_302,N_27831,N_26364);
nor UO_303 (O_303,N_27862,N_26415);
and UO_304 (O_304,N_28588,N_26120);
nand UO_305 (O_305,N_29307,N_29489);
nand UO_306 (O_306,N_25522,N_29716);
nor UO_307 (O_307,N_29230,N_26096);
nor UO_308 (O_308,N_27879,N_26898);
nand UO_309 (O_309,N_26684,N_26991);
and UO_310 (O_310,N_28264,N_28429);
nor UO_311 (O_311,N_28285,N_29737);
or UO_312 (O_312,N_27757,N_28004);
and UO_313 (O_313,N_27627,N_26761);
nand UO_314 (O_314,N_27124,N_28253);
nand UO_315 (O_315,N_28126,N_28186);
and UO_316 (O_316,N_27763,N_27547);
nand UO_317 (O_317,N_25842,N_27484);
and UO_318 (O_318,N_28814,N_27414);
xnor UO_319 (O_319,N_25138,N_28401);
nor UO_320 (O_320,N_26309,N_25293);
and UO_321 (O_321,N_25001,N_27783);
or UO_322 (O_322,N_27080,N_29976);
nor UO_323 (O_323,N_28385,N_25624);
nor UO_324 (O_324,N_28765,N_26810);
nor UO_325 (O_325,N_28254,N_29731);
nand UO_326 (O_326,N_25191,N_29529);
nand UO_327 (O_327,N_25919,N_28135);
nand UO_328 (O_328,N_28024,N_25756);
nand UO_329 (O_329,N_26162,N_27409);
or UO_330 (O_330,N_28352,N_29125);
nand UO_331 (O_331,N_27435,N_26766);
and UO_332 (O_332,N_29558,N_28504);
or UO_333 (O_333,N_27255,N_26911);
and UO_334 (O_334,N_25159,N_25497);
nor UO_335 (O_335,N_28376,N_27786);
nor UO_336 (O_336,N_26072,N_29278);
or UO_337 (O_337,N_26853,N_27819);
and UO_338 (O_338,N_25520,N_27018);
nor UO_339 (O_339,N_25721,N_25027);
and UO_340 (O_340,N_29041,N_28394);
and UO_341 (O_341,N_28300,N_27196);
or UO_342 (O_342,N_27698,N_28160);
or UO_343 (O_343,N_28888,N_27563);
or UO_344 (O_344,N_29449,N_29888);
nor UO_345 (O_345,N_26330,N_28003);
nor UO_346 (O_346,N_29297,N_26404);
xor UO_347 (O_347,N_25255,N_26053);
and UO_348 (O_348,N_29866,N_28335);
nor UO_349 (O_349,N_27290,N_25925);
xor UO_350 (O_350,N_27289,N_26074);
or UO_351 (O_351,N_25133,N_25282);
nor UO_352 (O_352,N_29759,N_27752);
and UO_353 (O_353,N_29585,N_25118);
nand UO_354 (O_354,N_26685,N_26635);
or UO_355 (O_355,N_25505,N_29261);
xnor UO_356 (O_356,N_25119,N_29532);
nor UO_357 (O_357,N_25747,N_27342);
nor UO_358 (O_358,N_25455,N_25214);
nor UO_359 (O_359,N_29050,N_27472);
nand UO_360 (O_360,N_25317,N_26797);
xor UO_361 (O_361,N_25813,N_28938);
and UO_362 (O_362,N_26388,N_26294);
and UO_363 (O_363,N_26643,N_27488);
and UO_364 (O_364,N_25250,N_29753);
or UO_365 (O_365,N_27207,N_28172);
xnor UO_366 (O_366,N_26318,N_26020);
and UO_367 (O_367,N_26515,N_26787);
and UO_368 (O_368,N_25324,N_26654);
nand UO_369 (O_369,N_28563,N_26650);
or UO_370 (O_370,N_29943,N_29378);
nor UO_371 (O_371,N_27034,N_25079);
nand UO_372 (O_372,N_28533,N_27191);
nand UO_373 (O_373,N_28789,N_25811);
and UO_374 (O_374,N_25235,N_28613);
nor UO_375 (O_375,N_29797,N_26924);
nand UO_376 (O_376,N_25835,N_27286);
nand UO_377 (O_377,N_27701,N_29176);
and UO_378 (O_378,N_29482,N_26735);
nand UO_379 (O_379,N_29108,N_29928);
nand UO_380 (O_380,N_25425,N_28531);
xnor UO_381 (O_381,N_25495,N_26927);
nand UO_382 (O_382,N_25309,N_26414);
nand UO_383 (O_383,N_25714,N_28222);
nor UO_384 (O_384,N_29567,N_25582);
xnor UO_385 (O_385,N_27517,N_29923);
nor UO_386 (O_386,N_29726,N_29353);
xnor UO_387 (O_387,N_29647,N_28689);
nand UO_388 (O_388,N_26292,N_29987);
nor UO_389 (O_389,N_29466,N_27135);
nor UO_390 (O_390,N_26021,N_25185);
nand UO_391 (O_391,N_27806,N_27638);
or UO_392 (O_392,N_25734,N_27569);
xnor UO_393 (O_393,N_25868,N_25923);
and UO_394 (O_394,N_27146,N_29949);
and UO_395 (O_395,N_25446,N_27902);
or UO_396 (O_396,N_27441,N_27423);
or UO_397 (O_397,N_29394,N_28417);
xor UO_398 (O_398,N_25394,N_26445);
or UO_399 (O_399,N_28157,N_29807);
and UO_400 (O_400,N_26713,N_25879);
or UO_401 (O_401,N_28078,N_26659);
xor UO_402 (O_402,N_29732,N_26396);
nand UO_403 (O_403,N_25951,N_29226);
or UO_404 (O_404,N_27980,N_29704);
and UO_405 (O_405,N_26097,N_26672);
xnor UO_406 (O_406,N_29745,N_26965);
or UO_407 (O_407,N_26918,N_29873);
nor UO_408 (O_408,N_29190,N_28746);
or UO_409 (O_409,N_28389,N_29719);
nand UO_410 (O_410,N_27390,N_25254);
or UO_411 (O_411,N_26647,N_27988);
and UO_412 (O_412,N_25158,N_27477);
and UO_413 (O_413,N_27006,N_25809);
xnor UO_414 (O_414,N_29306,N_29640);
and UO_415 (O_415,N_28259,N_28184);
and UO_416 (O_416,N_27369,N_25271);
nor UO_417 (O_417,N_29781,N_26123);
nor UO_418 (O_418,N_26435,N_28188);
or UO_419 (O_419,N_26579,N_25511);
nor UO_420 (O_420,N_25938,N_27327);
nor UO_421 (O_421,N_28863,N_27920);
nand UO_422 (O_422,N_28427,N_26447);
nor UO_423 (O_423,N_27564,N_26059);
nor UO_424 (O_424,N_27776,N_26714);
nor UO_425 (O_425,N_26816,N_25287);
and UO_426 (O_426,N_29180,N_25952);
or UO_427 (O_427,N_27604,N_29727);
or UO_428 (O_428,N_27764,N_29702);
nand UO_429 (O_429,N_28367,N_29506);
or UO_430 (O_430,N_28838,N_27415);
and UO_431 (O_431,N_26850,N_25230);
nand UO_432 (O_432,N_27068,N_28017);
xor UO_433 (O_433,N_25403,N_26966);
nor UO_434 (O_434,N_26832,N_26055);
or UO_435 (O_435,N_27227,N_25207);
or UO_436 (O_436,N_28987,N_26486);
nand UO_437 (O_437,N_26532,N_26054);
and UO_438 (O_438,N_29989,N_29915);
or UO_439 (O_439,N_28260,N_28302);
and UO_440 (O_440,N_26235,N_28544);
and UO_441 (O_441,N_28699,N_29249);
and UO_442 (O_442,N_29950,N_28644);
nand UO_443 (O_443,N_28320,N_29971);
nor UO_444 (O_444,N_26495,N_29764);
nand UO_445 (O_445,N_25000,N_28056);
or UO_446 (O_446,N_29164,N_27542);
nand UO_447 (O_447,N_28867,N_29243);
nand UO_448 (O_448,N_25010,N_26932);
xnor UO_449 (O_449,N_26972,N_28437);
and UO_450 (O_450,N_29834,N_27212);
nor UO_451 (O_451,N_29891,N_28406);
nand UO_452 (O_452,N_26088,N_27664);
or UO_453 (O_453,N_25151,N_26553);
nor UO_454 (O_454,N_26703,N_29983);
nand UO_455 (O_455,N_29994,N_25139);
nor UO_456 (O_456,N_29454,N_28614);
xor UO_457 (O_457,N_25791,N_27045);
and UO_458 (O_458,N_25150,N_29017);
nand UO_459 (O_459,N_27760,N_27837);
xor UO_460 (O_460,N_28808,N_26193);
nor UO_461 (O_461,N_29018,N_28999);
nand UO_462 (O_462,N_25100,N_26967);
nand UO_463 (O_463,N_27942,N_29251);
or UO_464 (O_464,N_29457,N_26796);
nor UO_465 (O_465,N_26302,N_28524);
nor UO_466 (O_466,N_27670,N_26902);
and UO_467 (O_467,N_26245,N_26176);
nor UO_468 (O_468,N_25940,N_28963);
nand UO_469 (O_469,N_25108,N_27025);
nor UO_470 (O_470,N_28946,N_29002);
or UO_471 (O_471,N_28119,N_28246);
nor UO_472 (O_472,N_26304,N_28634);
nand UO_473 (O_473,N_26039,N_26759);
nand UO_474 (O_474,N_26848,N_27921);
and UO_475 (O_475,N_28846,N_25389);
and UO_476 (O_476,N_25658,N_27797);
nor UO_477 (O_477,N_29831,N_28444);
or UO_478 (O_478,N_28136,N_29443);
xor UO_479 (O_479,N_29321,N_25891);
and UO_480 (O_480,N_29223,N_26641);
xnor UO_481 (O_481,N_25804,N_29755);
nand UO_482 (O_482,N_28411,N_29377);
or UO_483 (O_483,N_25148,N_25285);
nand UO_484 (O_484,N_28974,N_26583);
xnor UO_485 (O_485,N_29412,N_27064);
nor UO_486 (O_486,N_28421,N_26253);
nand UO_487 (O_487,N_27096,N_25996);
nor UO_488 (O_488,N_29566,N_28199);
or UO_489 (O_489,N_25199,N_25391);
and UO_490 (O_490,N_28461,N_27429);
nand UO_491 (O_491,N_27657,N_26200);
and UO_492 (O_492,N_26301,N_29115);
xor UO_493 (O_493,N_27445,N_26188);
nor UO_494 (O_494,N_28275,N_28772);
or UO_495 (O_495,N_25669,N_26744);
nand UO_496 (O_496,N_25908,N_25547);
nor UO_497 (O_497,N_29010,N_25660);
nor UO_498 (O_498,N_26588,N_26430);
and UO_499 (O_499,N_28162,N_25981);
nor UO_500 (O_500,N_28969,N_27863);
nand UO_501 (O_501,N_25910,N_29752);
xor UO_502 (O_502,N_29452,N_29774);
xnor UO_503 (O_503,N_26518,N_29691);
xnor UO_504 (O_504,N_27534,N_27473);
nor UO_505 (O_505,N_28837,N_28624);
and UO_506 (O_506,N_26544,N_28728);
xnor UO_507 (O_507,N_27309,N_29253);
or UO_508 (O_508,N_27949,N_29030);
nor UO_509 (O_509,N_28471,N_28435);
and UO_510 (O_510,N_25308,N_26344);
xor UO_511 (O_511,N_29644,N_26707);
xor UO_512 (O_512,N_29240,N_25176);
and UO_513 (O_513,N_25506,N_25532);
nand UO_514 (O_514,N_27095,N_28847);
and UO_515 (O_515,N_28697,N_27972);
nand UO_516 (O_516,N_27554,N_28404);
or UO_517 (O_517,N_27189,N_25664);
xor UO_518 (O_518,N_26751,N_27671);
or UO_519 (O_519,N_27665,N_28630);
xnor UO_520 (O_520,N_25213,N_29109);
nor UO_521 (O_521,N_29679,N_25366);
and UO_522 (O_522,N_25210,N_25703);
nor UO_523 (O_523,N_25626,N_26772);
nand UO_524 (O_524,N_26239,N_29437);
nand UO_525 (O_525,N_25935,N_26721);
and UO_526 (O_526,N_28156,N_27224);
nand UO_527 (O_527,N_29901,N_27244);
xor UO_528 (O_528,N_27592,N_27464);
nor UO_529 (O_529,N_28106,N_29393);
nand UO_530 (O_530,N_28931,N_26846);
or UO_531 (O_531,N_25012,N_26382);
nand UO_532 (O_532,N_27298,N_28620);
nor UO_533 (O_533,N_27560,N_27198);
or UO_534 (O_534,N_29234,N_26547);
and UO_535 (O_535,N_27361,N_29988);
nand UO_536 (O_536,N_27150,N_25346);
nor UO_537 (O_537,N_29758,N_27497);
nand UO_538 (O_538,N_25979,N_28565);
and UO_539 (O_539,N_27739,N_25135);
nand UO_540 (O_540,N_28572,N_29688);
and UO_541 (O_541,N_29218,N_29462);
or UO_542 (O_542,N_26195,N_25046);
and UO_543 (O_543,N_25657,N_27841);
nand UO_544 (O_544,N_29562,N_27354);
and UO_545 (O_545,N_29818,N_26938);
and UO_546 (O_546,N_26642,N_27506);
or UO_547 (O_547,N_29119,N_26171);
xor UO_548 (O_548,N_27915,N_25299);
xor UO_549 (O_549,N_29997,N_28923);
nand UO_550 (O_550,N_27287,N_27262);
nor UO_551 (O_551,N_28955,N_28183);
and UO_552 (O_552,N_29274,N_28327);
and UO_553 (O_553,N_28021,N_26536);
nand UO_554 (O_554,N_25899,N_25251);
xor UO_555 (O_555,N_26000,N_28781);
xnor UO_556 (O_556,N_25974,N_27118);
nor UO_557 (O_557,N_28911,N_26038);
or UO_558 (O_558,N_25982,N_25515);
nor UO_559 (O_559,N_29113,N_28052);
nor UO_560 (O_560,N_27066,N_25517);
nor UO_561 (O_561,N_29244,N_29368);
nand UO_562 (O_562,N_25502,N_27199);
and UO_563 (O_563,N_28400,N_25437);
nand UO_564 (O_564,N_25733,N_27008);
nand UO_565 (O_565,N_27083,N_26266);
or UO_566 (O_566,N_27179,N_25457);
and UO_567 (O_567,N_26221,N_28625);
and UO_568 (O_568,N_29042,N_29140);
nand UO_569 (O_569,N_25365,N_27705);
xor UO_570 (O_570,N_29635,N_29039);
nor UO_571 (O_571,N_26567,N_26987);
nand UO_572 (O_572,N_25550,N_27630);
and UO_573 (O_573,N_27524,N_26472);
nand UO_574 (O_574,N_28840,N_25866);
nor UO_575 (O_575,N_25632,N_27678);
nor UO_576 (O_576,N_29761,N_26514);
and UO_577 (O_577,N_26270,N_29754);
nor UO_578 (O_578,N_25663,N_25954);
xnor UO_579 (O_579,N_26164,N_27226);
or UO_580 (O_580,N_28959,N_28419);
nand UO_581 (O_581,N_26361,N_28793);
nor UO_582 (O_582,N_26502,N_29592);
nor UO_583 (O_583,N_29627,N_28538);
nand UO_584 (O_584,N_29023,N_28303);
or UO_585 (O_585,N_27754,N_27111);
nand UO_586 (O_586,N_25857,N_25725);
or UO_587 (O_587,N_28901,N_25788);
and UO_588 (O_588,N_28226,N_26929);
xnor UO_589 (O_589,N_26498,N_25622);
or UO_590 (O_590,N_27886,N_26370);
nor UO_591 (O_591,N_25451,N_28262);
and UO_592 (O_592,N_28463,N_25545);
and UO_593 (O_593,N_25706,N_29420);
or UO_594 (O_594,N_29711,N_26150);
or UO_595 (O_595,N_28103,N_26576);
and UO_596 (O_596,N_28339,N_25764);
and UO_597 (O_597,N_28201,N_29659);
or UO_598 (O_598,N_26434,N_29441);
and UO_599 (O_599,N_25386,N_26114);
nand UO_600 (O_600,N_27640,N_28434);
or UO_601 (O_601,N_28548,N_28204);
nor UO_602 (O_602,N_29646,N_25378);
or UO_603 (O_603,N_29383,N_26118);
nor UO_604 (O_604,N_28055,N_29625);
and UO_605 (O_605,N_26628,N_28391);
or UO_606 (O_606,N_29363,N_27442);
nor UO_607 (O_607,N_26337,N_27958);
nor UO_608 (O_608,N_29475,N_27861);
nor UO_609 (O_609,N_28359,N_28238);
xor UO_610 (O_610,N_26612,N_27300);
and UO_611 (O_611,N_25889,N_25421);
or UO_612 (O_612,N_27746,N_27380);
or UO_613 (O_613,N_26826,N_29655);
nand UO_614 (O_614,N_29820,N_29031);
nand UO_615 (O_615,N_29151,N_28598);
xor UO_616 (O_616,N_25167,N_26631);
and UO_617 (O_617,N_29601,N_28407);
and UO_618 (O_618,N_26305,N_25668);
nand UO_619 (O_619,N_29079,N_25351);
nand UO_620 (O_620,N_25286,N_29643);
or UO_621 (O_621,N_26306,N_28155);
xnor UO_622 (O_622,N_25798,N_29975);
and UO_623 (O_623,N_25964,N_29311);
or UO_624 (O_624,N_28979,N_27898);
xor UO_625 (O_625,N_25915,N_29881);
nor UO_626 (O_626,N_28871,N_26481);
and UO_627 (O_627,N_27330,N_26342);
nor UO_628 (O_628,N_26130,N_26463);
and UO_629 (O_629,N_25504,N_28278);
nor UO_630 (O_630,N_28197,N_28681);
nor UO_631 (O_631,N_28558,N_26517);
xnor UO_632 (O_632,N_29693,N_29710);
or UO_633 (O_633,N_25379,N_28284);
xor UO_634 (O_634,N_27614,N_28450);
xnor UO_635 (O_635,N_27595,N_29678);
nand UO_636 (O_636,N_28384,N_25237);
nor UO_637 (O_637,N_29615,N_29878);
nand UO_638 (O_638,N_29035,N_25712);
xnor UO_639 (O_639,N_29619,N_26261);
and UO_640 (O_640,N_26136,N_29157);
and UO_641 (O_641,N_29852,N_26990);
xnor UO_642 (O_642,N_27605,N_27724);
nor UO_643 (O_643,N_26715,N_27440);
and UO_644 (O_644,N_29425,N_25252);
nand UO_645 (O_645,N_28550,N_26492);
nand UO_646 (O_646,N_26692,N_28405);
nor UO_647 (O_647,N_26770,N_26033);
xnor UO_648 (O_648,N_28153,N_26351);
nor UO_649 (O_649,N_26695,N_28211);
or UO_650 (O_650,N_25161,N_29876);
nor UO_651 (O_651,N_28115,N_28245);
nor UO_652 (O_652,N_29528,N_25794);
or UO_653 (O_653,N_27704,N_25305);
xor UO_654 (O_654,N_29336,N_29877);
xor UO_655 (O_655,N_26633,N_28457);
and UO_656 (O_656,N_28089,N_26984);
or UO_657 (O_657,N_26540,N_28063);
nand UO_658 (O_658,N_28440,N_25278);
nand UO_659 (O_659,N_28082,N_25170);
or UO_660 (O_660,N_27767,N_27546);
nand UO_661 (O_661,N_29548,N_26336);
and UO_662 (O_662,N_28649,N_26798);
nor UO_663 (O_663,N_26156,N_25450);
nand UO_664 (O_664,N_27419,N_25692);
nor UO_665 (O_665,N_28956,N_28712);
nor UO_666 (O_666,N_27311,N_29444);
nor UO_667 (O_667,N_27734,N_27251);
and UO_668 (O_668,N_29733,N_25541);
or UO_669 (O_669,N_29283,N_26599);
or UO_670 (O_670,N_27697,N_28460);
or UO_671 (O_671,N_26768,N_28071);
or UO_672 (O_672,N_29842,N_28973);
xnor UO_673 (O_673,N_27293,N_25708);
xnor UO_674 (O_674,N_25948,N_28578);
nand UO_675 (O_675,N_26355,N_27337);
nor UO_676 (O_676,N_25267,N_26568);
or UO_677 (O_677,N_29100,N_25796);
or UO_678 (O_678,N_25247,N_29011);
nand UO_679 (O_679,N_29367,N_25792);
nor UO_680 (O_680,N_25052,N_26110);
or UO_681 (O_681,N_27707,N_26969);
or UO_682 (O_682,N_25060,N_28688);
or UO_683 (O_683,N_26516,N_29618);
nand UO_684 (O_684,N_28030,N_26190);
nand UO_685 (O_685,N_25384,N_28816);
nor UO_686 (O_686,N_27973,N_26484);
nand UO_687 (O_687,N_29954,N_27695);
xor UO_688 (O_688,N_28337,N_29611);
nor UO_689 (O_689,N_27428,N_28967);
and UO_690 (O_690,N_29632,N_25244);
nand UO_691 (O_691,N_26885,N_25190);
and UO_692 (O_692,N_27565,N_27832);
or UO_693 (O_693,N_27941,N_25799);
or UO_694 (O_694,N_27711,N_25565);
nor UO_695 (O_695,N_26437,N_27594);
xnor UO_696 (O_696,N_29127,N_28274);
nor UO_697 (O_697,N_27125,N_26783);
nand UO_698 (O_698,N_29893,N_29439);
and UO_699 (O_699,N_29541,N_25784);
xnor UO_700 (O_700,N_26901,N_29850);
or UO_701 (O_701,N_26177,N_27839);
xnor UO_702 (O_702,N_25641,N_26449);
nor UO_703 (O_703,N_29573,N_29497);
and UO_704 (O_704,N_25702,N_25606);
or UO_705 (O_705,N_28676,N_28933);
nor UO_706 (O_706,N_25888,N_29369);
nand UO_707 (O_707,N_27396,N_29723);
or UO_708 (O_708,N_28554,N_28216);
nor UO_709 (O_709,N_27531,N_28535);
xnor UO_710 (O_710,N_27963,N_29073);
nor UO_711 (O_711,N_25280,N_28971);
nand UO_712 (O_712,N_26283,N_27404);
or UO_713 (O_713,N_26795,N_26483);
and UO_714 (O_714,N_27616,N_28875);
and UO_715 (O_715,N_29359,N_25860);
and UO_716 (O_716,N_25197,N_25156);
nand UO_717 (O_717,N_25609,N_26227);
nor UO_718 (O_718,N_28042,N_29036);
nand UO_719 (O_719,N_26512,N_27126);
and UO_720 (O_720,N_25340,N_28560);
nor UO_721 (O_721,N_29169,N_25594);
or UO_722 (O_722,N_25023,N_25677);
nand UO_723 (O_723,N_28100,N_29846);
nor UO_724 (O_724,N_29401,N_26440);
nor UO_725 (O_725,N_28803,N_26386);
or UO_726 (O_726,N_29520,N_25629);
nor UO_727 (O_727,N_27340,N_29173);
and UO_728 (O_728,N_29488,N_25670);
or UO_729 (O_729,N_25755,N_27385);
nor UO_730 (O_730,N_25895,N_29319);
or UO_731 (O_731,N_27245,N_28398);
and UO_732 (O_732,N_27593,N_27106);
and UO_733 (O_733,N_28859,N_28086);
nor UO_734 (O_734,N_25243,N_29492);
nor UO_735 (O_735,N_26263,N_28545);
nor UO_736 (O_736,N_28828,N_29925);
nor UO_737 (O_737,N_26267,N_25101);
nor UO_738 (O_738,N_26978,N_25072);
nand UO_739 (O_739,N_29064,N_25675);
nor UO_740 (O_740,N_25781,N_29149);
and UO_741 (O_741,N_28592,N_26774);
or UO_742 (O_742,N_27700,N_28823);
or UO_743 (O_743,N_25062,N_28887);
nand UO_744 (O_744,N_27129,N_28272);
or UO_745 (O_745,N_27217,N_29184);
and UO_746 (O_746,N_28593,N_25117);
xor UO_747 (O_747,N_28799,N_27335);
nor UO_748 (O_748,N_26909,N_27570);
xnor UO_749 (O_749,N_26894,N_29187);
and UO_750 (O_750,N_28589,N_27790);
or UO_751 (O_751,N_27591,N_27213);
or UO_752 (O_752,N_25526,N_27110);
nand UO_753 (O_753,N_27641,N_28742);
nand UO_754 (O_754,N_28683,N_28170);
and UO_755 (O_755,N_25094,N_25649);
or UO_756 (O_756,N_29145,N_26107);
or UO_757 (O_757,N_25483,N_29265);
nand UO_758 (O_758,N_27260,N_28281);
nor UO_759 (O_759,N_27625,N_28134);
nand UO_760 (O_760,N_27976,N_27676);
and UO_761 (O_761,N_27382,N_27463);
and UO_762 (O_762,N_29056,N_27060);
or UO_763 (O_763,N_25469,N_25034);
or UO_764 (O_764,N_29572,N_29934);
or UO_765 (O_765,N_29965,N_25203);
nand UO_766 (O_766,N_27346,N_28800);
and UO_767 (O_767,N_27586,N_28813);
or UO_768 (O_768,N_26864,N_27200);
and UO_769 (O_769,N_25054,N_28431);
or UO_770 (O_770,N_25422,N_29969);
nor UO_771 (O_771,N_27157,N_25944);
nor UO_772 (O_772,N_27081,N_27679);
or UO_773 (O_773,N_25719,N_27723);
nor UO_774 (O_774,N_27381,N_27307);
or UO_775 (O_775,N_25315,N_25336);
nor UO_776 (O_776,N_27273,N_25508);
xor UO_777 (O_777,N_27326,N_28424);
and UO_778 (O_778,N_29008,N_25753);
or UO_779 (O_779,N_27149,N_27512);
or UO_780 (O_780,N_25332,N_29730);
nand UO_781 (O_781,N_28496,N_28079);
or UO_782 (O_782,N_28590,N_29516);
and UO_783 (O_783,N_26477,N_28288);
and UO_784 (O_784,N_25834,N_27878);
and UO_785 (O_785,N_28255,N_25513);
or UO_786 (O_786,N_28263,N_29591);
and UO_787 (O_787,N_26729,N_29078);
and UO_788 (O_788,N_28658,N_27632);
or UO_789 (O_789,N_28954,N_29556);
nor UO_790 (O_790,N_29458,N_25743);
nor UO_791 (O_791,N_28647,N_28242);
nand UO_792 (O_792,N_28752,N_27105);
and UO_793 (O_793,N_26140,N_26841);
nand UO_794 (O_794,N_28168,N_27505);
or UO_795 (O_795,N_29616,N_29649);
nor UO_796 (O_796,N_29855,N_26952);
xor UO_797 (O_797,N_29126,N_29884);
or UO_798 (O_798,N_27559,N_26233);
or UO_799 (O_799,N_26115,N_27029);
nand UO_800 (O_800,N_27602,N_29293);
xnor UO_801 (O_801,N_25906,N_26663);
nor UO_802 (O_802,N_27466,N_25892);
nor UO_803 (O_803,N_27090,N_28044);
or UO_804 (O_804,N_25548,N_26745);
or UO_805 (O_805,N_25104,N_25330);
and UO_806 (O_806,N_25126,N_26326);
nor UO_807 (O_807,N_26323,N_28886);
and UO_808 (O_808,N_25918,N_27225);
nand UO_809 (O_809,N_25745,N_27363);
nand UO_810 (O_810,N_28072,N_27331);
or UO_811 (O_811,N_27742,N_29304);
nor UO_812 (O_812,N_28088,N_28468);
and UO_813 (O_813,N_27934,N_29471);
nor UO_814 (O_814,N_28507,N_28845);
and UO_815 (O_815,N_25546,N_27533);
and UO_816 (O_816,N_28920,N_27272);
nor UO_817 (O_817,N_29081,N_29469);
xnor UO_818 (O_818,N_28992,N_27324);
and UO_819 (O_819,N_28217,N_29760);
nand UO_820 (O_820,N_25969,N_28913);
nor UO_821 (O_821,N_28788,N_26598);
or UO_822 (O_822,N_26103,N_29798);
xor UO_823 (O_823,N_25682,N_28951);
or UO_824 (O_824,N_27498,N_28804);
nor UO_825 (O_825,N_29193,N_26658);
and UO_826 (O_826,N_25018,N_28551);
nor UO_827 (O_827,N_29181,N_26087);
or UO_828 (O_828,N_25815,N_26881);
nor UO_829 (O_829,N_29662,N_29174);
and UO_830 (O_830,N_26327,N_26577);
and UO_831 (O_831,N_29236,N_29135);
or UO_832 (O_832,N_25265,N_26839);
xnor UO_833 (O_833,N_29606,N_29178);
nor UO_834 (O_834,N_25294,N_28543);
nor UO_835 (O_835,N_28139,N_25611);
nand UO_836 (O_836,N_26584,N_25699);
and UO_837 (O_837,N_27957,N_27132);
nor UO_838 (O_838,N_26231,N_28453);
nor UO_839 (O_839,N_29784,N_26908);
xnor UO_840 (O_840,N_28801,N_29772);
xor UO_841 (O_841,N_29786,N_26432);
or UO_842 (O_842,N_27065,N_29012);
or UO_843 (O_843,N_28110,N_28915);
xor UO_844 (O_844,N_28966,N_28508);
and UO_845 (O_845,N_25464,N_29512);
nor UO_846 (O_846,N_27139,N_29194);
or UO_847 (O_847,N_29555,N_29480);
or UO_848 (O_848,N_26867,N_26377);
nand UO_849 (O_849,N_27811,N_29599);
nand UO_850 (O_850,N_28998,N_29399);
nor UO_851 (O_851,N_28710,N_27238);
nor UO_852 (O_852,N_29003,N_25169);
nand UO_853 (O_853,N_29748,N_26381);
and UO_854 (O_854,N_27055,N_28735);
or UO_855 (O_855,N_28297,N_28102);
nor UO_856 (O_856,N_29410,N_26668);
nor UO_857 (O_857,N_25482,N_27082);
nand UO_858 (O_858,N_29687,N_27787);
nor UO_859 (O_859,N_25395,N_29381);
nand UO_860 (O_860,N_27789,N_29371);
nand UO_861 (O_861,N_26870,N_28289);
nand UO_862 (O_862,N_28629,N_25748);
or UO_863 (O_863,N_29456,N_29239);
nand UO_864 (O_864,N_26609,N_29034);
and UO_865 (O_865,N_28948,N_28612);
nand UO_866 (O_866,N_29992,N_29298);
xor UO_867 (O_867,N_27109,N_28383);
nand UO_868 (O_868,N_25744,N_25130);
nor UO_869 (O_869,N_26767,N_27962);
and UO_870 (O_870,N_25276,N_29349);
and UO_871 (O_871,N_26921,N_25415);
or UO_872 (O_872,N_26802,N_29523);
or UO_873 (O_873,N_26391,N_25540);
or UO_874 (O_874,N_29902,N_27386);
nor UO_875 (O_875,N_27356,N_27486);
or UO_876 (O_876,N_28240,N_25579);
nand UO_877 (O_877,N_28501,N_27558);
or UO_878 (O_878,N_28393,N_29605);
xnor UO_879 (O_879,N_28169,N_26147);
and UO_880 (O_880,N_28006,N_28241);
xor UO_881 (O_881,N_27254,N_27693);
or UO_882 (O_882,N_26138,N_29813);
nand UO_883 (O_883,N_28843,N_25275);
nor UO_884 (O_884,N_29396,N_29269);
or UO_885 (O_885,N_28868,N_29911);
nand UO_886 (O_886,N_28101,N_28591);
nand UO_887 (O_887,N_29013,N_27427);
or UO_888 (O_888,N_28085,N_29863);
and UO_889 (O_889,N_29186,N_26511);
and UO_890 (O_890,N_29020,N_27802);
and UO_891 (O_891,N_28035,N_29744);
nor UO_892 (O_892,N_26044,N_25066);
nand UO_893 (O_893,N_29795,N_29262);
and UO_894 (O_894,N_29001,N_26444);
nand UO_895 (O_895,N_25318,N_26402);
or UO_896 (O_896,N_25962,N_29517);
nand UO_897 (O_897,N_27654,N_27232);
and UO_898 (O_898,N_25650,N_27214);
and UO_899 (O_899,N_25024,N_26716);
nand UO_900 (O_900,N_26880,N_25187);
nor UO_901 (O_901,N_26688,N_27820);
nand UO_902 (O_902,N_26001,N_26446);
nand UO_903 (O_903,N_26078,N_26197);
nand UO_904 (O_904,N_28092,N_28517);
nand UO_905 (O_905,N_25053,N_26276);
nor UO_906 (O_906,N_29266,N_29246);
xnor UO_907 (O_907,N_27320,N_27572);
nand UO_908 (O_908,N_26222,N_27476);
or UO_909 (O_909,N_26812,N_26428);
and UO_910 (O_910,N_29460,N_26575);
xor UO_911 (O_911,N_29951,N_26676);
and UO_912 (O_912,N_27156,N_29854);
xor UO_913 (O_913,N_25931,N_26374);
xor UO_914 (O_914,N_27818,N_29101);
xor UO_915 (O_915,N_28307,N_25705);
nor UO_916 (O_916,N_29839,N_29310);
nor UO_917 (O_917,N_27002,N_26691);
nor UO_918 (O_918,N_25638,N_25222);
nor UO_919 (O_919,N_29634,N_28493);
nor UO_920 (O_920,N_28397,N_26218);
or UO_921 (O_921,N_26585,N_27321);
nand UO_922 (O_922,N_29650,N_28792);
nand UO_923 (O_923,N_25581,N_25028);
or UO_924 (O_924,N_26892,N_28903);
or UO_925 (O_925,N_27392,N_29947);
or UO_926 (O_926,N_25742,N_29708);
xnor UO_927 (O_927,N_25398,N_26476);
nand UO_928 (O_928,N_29519,N_28957);
and UO_929 (O_929,N_28485,N_29029);
and UO_930 (O_930,N_27123,N_28373);
nand UO_931 (O_931,N_27343,N_29245);
nor UO_932 (O_932,N_27788,N_28856);
and UO_933 (O_933,N_25690,N_29047);
nor UO_934 (O_934,N_26490,N_26368);
and UO_935 (O_935,N_26947,N_25667);
nand UO_936 (O_936,N_29654,N_29782);
nor UO_937 (O_937,N_27315,N_27400);
nor UO_938 (O_938,N_29565,N_25372);
or UO_939 (O_939,N_29603,N_27259);
xor UO_940 (O_940,N_25056,N_29690);
xnor UO_941 (O_941,N_28898,N_26570);
or UO_942 (O_942,N_26244,N_26572);
or UO_943 (O_943,N_25193,N_25890);
and UO_944 (O_944,N_28002,N_28621);
and UO_945 (O_945,N_26539,N_29827);
or UO_946 (O_946,N_28646,N_25303);
and UO_947 (O_947,N_25037,N_28013);
nand UO_948 (O_948,N_26343,N_27989);
or UO_949 (O_949,N_27297,N_26998);
nor UO_950 (O_950,N_29857,N_27883);
nand UO_951 (O_951,N_27044,N_25551);
or UO_952 (O_952,N_28773,N_28568);
and UO_953 (O_953,N_28635,N_27552);
or UO_954 (O_954,N_27618,N_29788);
nor UO_955 (O_955,N_27033,N_25189);
nand UO_956 (O_956,N_25175,N_26600);
or UO_957 (O_957,N_26855,N_25598);
nor UO_958 (O_958,N_28806,N_29474);
or UO_959 (O_959,N_27836,N_26015);
or UO_960 (O_960,N_27650,N_28491);
nor UO_961 (O_961,N_27613,N_28271);
xnor UO_962 (O_962,N_29680,N_28282);
nor UO_963 (O_963,N_27823,N_29467);
nor UO_964 (O_964,N_26124,N_29057);
or UO_965 (O_965,N_26950,N_27071);
nand UO_966 (O_966,N_29498,N_27930);
xor UO_967 (O_967,N_25576,N_29964);
nor UO_968 (O_968,N_28696,N_29511);
and UO_969 (O_969,N_27761,N_26251);
nand UO_970 (O_970,N_29009,N_29963);
or UO_971 (O_971,N_29561,N_27600);
xor UO_972 (O_972,N_26126,N_28362);
and UO_973 (O_973,N_28007,N_28505);
xor UO_974 (O_974,N_29767,N_25640);
nand UO_975 (O_975,N_29570,N_28466);
and UO_976 (O_976,N_27134,N_26834);
or UO_977 (O_977,N_27360,N_27738);
nand UO_978 (O_978,N_29593,N_27078);
xnor UO_979 (O_979,N_27411,N_27170);
xnor UO_980 (O_980,N_25571,N_25718);
and UO_981 (O_981,N_28585,N_27069);
and UO_982 (O_982,N_28150,N_25454);
and UO_983 (O_983,N_29579,N_26474);
nand UO_984 (O_984,N_25406,N_27113);
xor UO_985 (O_985,N_27912,N_27900);
nand UO_986 (O_986,N_25713,N_25153);
nor UO_987 (O_987,N_29749,N_25779);
nand UO_988 (O_988,N_29134,N_29433);
or UO_989 (O_989,N_25205,N_29794);
xor UO_990 (O_990,N_27964,N_29851);
or UO_991 (O_991,N_26104,N_27635);
nor UO_992 (O_992,N_25586,N_26213);
and UO_993 (O_993,N_26828,N_28495);
nand UO_994 (O_994,N_26763,N_25316);
and UO_995 (O_995,N_28749,N_26380);
nor UO_996 (O_996,N_25627,N_25288);
nor UO_997 (O_997,N_25978,N_25911);
xnor UO_998 (O_998,N_25323,N_25876);
nor UO_999 (O_999,N_29525,N_28433);
nor UO_1000 (O_1000,N_29568,N_29330);
or UO_1001 (O_1001,N_25852,N_28701);
and UO_1002 (O_1002,N_29426,N_28477);
xnor UO_1003 (O_1003,N_28166,N_28750);
nor UO_1004 (O_1004,N_26487,N_28884);
and UO_1005 (O_1005,N_28012,N_25771);
and UO_1006 (O_1006,N_29473,N_27647);
nor UO_1007 (O_1007,N_26762,N_26636);
xnor UO_1008 (O_1008,N_29342,N_29131);
nor UO_1009 (O_1009,N_29932,N_26944);
nor UO_1010 (O_1010,N_26027,N_25655);
or UO_1011 (O_1011,N_29419,N_25810);
and UO_1012 (O_1012,N_29651,N_26601);
nand UO_1013 (O_1013,N_27412,N_26537);
or UO_1014 (O_1014,N_29509,N_29777);
xor UO_1015 (O_1015,N_25983,N_27177);
or UO_1016 (O_1016,N_25382,N_29515);
or UO_1017 (O_1017,N_25929,N_25179);
xnor UO_1018 (O_1018,N_29022,N_26893);
nand UO_1019 (O_1019,N_29066,N_27849);
or UO_1020 (O_1020,N_27779,N_27793);
nor UO_1021 (O_1021,N_26457,N_28776);
nand UO_1022 (O_1022,N_29835,N_29271);
and UO_1023 (O_1023,N_27929,N_26202);
and UO_1024 (O_1024,N_27910,N_28000);
and UO_1025 (O_1025,N_27514,N_27745);
or UO_1026 (O_1026,N_29666,N_29325);
and UO_1027 (O_1027,N_29400,N_29264);
and UO_1028 (O_1028,N_28659,N_28641);
and UO_1029 (O_1029,N_25099,N_29301);
xnor UO_1030 (O_1030,N_29872,N_27961);
nor UO_1031 (O_1031,N_29544,N_28768);
and UO_1032 (O_1032,N_28392,N_27020);
nor UO_1033 (O_1033,N_29860,N_29552);
or UO_1034 (O_1034,N_25327,N_27495);
nor UO_1035 (O_1035,N_26578,N_25659);
or UO_1036 (O_1036,N_29446,N_26400);
nor UO_1037 (O_1037,N_27336,N_28663);
nor UO_1038 (O_1038,N_26265,N_29580);
and UO_1039 (O_1039,N_29152,N_29575);
or UO_1040 (O_1040,N_26779,N_26731);
and UO_1041 (O_1041,N_27719,N_25795);
or UO_1042 (O_1042,N_25468,N_29499);
nand UO_1043 (O_1043,N_29138,N_27407);
nand UO_1044 (O_1044,N_25177,N_28480);
xnor UO_1045 (O_1045,N_26187,N_25936);
and UO_1046 (O_1046,N_27276,N_26955);
nand UO_1047 (O_1047,N_25124,N_28426);
nor UO_1048 (O_1048,N_27329,N_25204);
or UO_1049 (O_1049,N_27525,N_28008);
or UO_1050 (O_1050,N_29204,N_29641);
nor UO_1051 (O_1051,N_26338,N_27903);
and UO_1052 (O_1052,N_26291,N_29663);
nor UO_1053 (O_1053,N_27133,N_27265);
and UO_1054 (O_1054,N_25440,N_28961);
and UO_1055 (O_1055,N_29914,N_29924);
nand UO_1056 (O_1056,N_28317,N_28706);
nor UO_1057 (O_1057,N_28601,N_28777);
nand UO_1058 (O_1058,N_28368,N_25578);
nand UO_1059 (O_1059,N_27303,N_26738);
xnor UO_1060 (O_1060,N_26372,N_27047);
nand UO_1061 (O_1061,N_29004,N_28148);
and UO_1062 (O_1062,N_29849,N_25463);
and UO_1063 (O_1063,N_28672,N_27379);
nor UO_1064 (O_1064,N_28096,N_25773);
nor UO_1065 (O_1065,N_29811,N_25674);
or UO_1066 (O_1066,N_25846,N_29461);
nand UO_1067 (O_1067,N_26769,N_28902);
nor UO_1068 (O_1068,N_26605,N_28185);
and UO_1069 (O_1069,N_25091,N_27117);
xor UO_1070 (O_1070,N_27193,N_26499);
or UO_1071 (O_1071,N_26904,N_25376);
nand UO_1072 (O_1072,N_25955,N_25009);
and UO_1073 (O_1073,N_25941,N_28964);
nand UO_1074 (O_1074,N_27518,N_28812);
xnor UO_1075 (O_1075,N_26638,N_25828);
and UO_1076 (O_1076,N_27986,N_27805);
and UO_1077 (O_1077,N_26259,N_25013);
or UO_1078 (O_1078,N_28986,N_26931);
or UO_1079 (O_1079,N_26209,N_27540);
nand UO_1080 (O_1080,N_28309,N_29123);
or UO_1081 (O_1081,N_29087,N_29946);
xnor UO_1082 (O_1082,N_29814,N_29326);
or UO_1083 (O_1083,N_27545,N_27946);
nor UO_1084 (O_1084,N_28498,N_26137);
and UO_1085 (O_1085,N_28797,N_28693);
and UO_1086 (O_1086,N_28536,N_28527);
or UO_1087 (O_1087,N_29610,N_26519);
nor UO_1088 (O_1088,N_27210,N_25084);
nor UO_1089 (O_1089,N_29669,N_27945);
nor UO_1090 (O_1090,N_25933,N_29898);
xnor UO_1091 (O_1091,N_26709,N_25816);
xor UO_1092 (O_1092,N_28364,N_25928);
nand UO_1093 (O_1093,N_29341,N_29089);
nor UO_1094 (O_1094,N_29074,N_29703);
or UO_1095 (O_1095,N_28409,N_25430);
and UO_1096 (O_1096,N_29095,N_26108);
nor UO_1097 (O_1097,N_28830,N_28523);
nand UO_1098 (O_1098,N_27870,N_26727);
and UO_1099 (O_1099,N_25466,N_29604);
or UO_1100 (O_1100,N_25575,N_26228);
or UO_1101 (O_1101,N_25841,N_27730);
xnor UO_1102 (O_1102,N_26644,N_28889);
and UO_1103 (O_1103,N_27075,N_26903);
or UO_1104 (O_1104,N_28739,N_27822);
and UO_1105 (O_1105,N_25814,N_29909);
nor UO_1106 (O_1106,N_29417,N_26070);
or UO_1107 (O_1107,N_26726,N_27278);
nor UO_1108 (O_1108,N_27607,N_26293);
and UO_1109 (O_1109,N_29069,N_25897);
xor UO_1110 (O_1110,N_29139,N_25570);
and UO_1111 (O_1111,N_27282,N_28784);
or UO_1112 (O_1112,N_26007,N_27504);
or UO_1113 (O_1113,N_25845,N_29289);
nand UO_1114 (O_1114,N_28324,N_25562);
nor UO_1115 (O_1115,N_26670,N_26613);
and UO_1116 (O_1116,N_25077,N_25516);
or UO_1117 (O_1117,N_28388,N_25147);
nor UO_1118 (O_1118,N_25830,N_25058);
xnor UO_1119 (O_1119,N_25854,N_26551);
or UO_1120 (O_1120,N_25473,N_28811);
nor UO_1121 (O_1121,N_25656,N_26900);
and UO_1122 (O_1122,N_28542,N_25824);
nand UO_1123 (O_1123,N_28610,N_26823);
nand UO_1124 (O_1124,N_27573,N_26760);
xor UO_1125 (O_1125,N_26945,N_25603);
nor UO_1126 (O_1126,N_26992,N_26247);
nor UO_1127 (O_1127,N_28023,N_27733);
nor UO_1128 (O_1128,N_26624,N_28618);
and UO_1129 (O_1129,N_28878,N_28512);
or UO_1130 (O_1130,N_28723,N_27800);
nand UO_1131 (O_1131,N_27643,N_27703);
nand UO_1132 (O_1132,N_25608,N_29320);
nor UO_1133 (O_1133,N_27673,N_25209);
or UO_1134 (O_1134,N_27583,N_25112);
nand UO_1135 (O_1135,N_28481,N_26923);
and UO_1136 (O_1136,N_28048,N_25107);
and UO_1137 (O_1137,N_28494,N_28611);
and UO_1138 (O_1138,N_27794,N_28632);
nor UO_1139 (O_1139,N_25301,N_26454);
and UO_1140 (O_1140,N_28236,N_26408);
nand UO_1141 (O_1141,N_27651,N_28177);
nor UO_1142 (O_1142,N_29793,N_26152);
nand UO_1143 (O_1143,N_28755,N_27122);
nand UO_1144 (O_1144,N_29995,N_26105);
nand UO_1145 (O_1145,N_28528,N_25566);
xor UO_1146 (O_1146,N_26976,N_27182);
nand UO_1147 (O_1147,N_29757,N_25858);
and UO_1148 (O_1148,N_25232,N_28073);
nor UO_1149 (O_1149,N_28142,N_29912);
or UO_1150 (O_1150,N_25435,N_27645);
and UO_1151 (O_1151,N_25797,N_29870);
nand UO_1152 (O_1152,N_28342,N_28704);
or UO_1153 (O_1153,N_26085,N_27567);
and UO_1154 (O_1154,N_26220,N_25011);
and UO_1155 (O_1155,N_29768,N_26436);
nor UO_1156 (O_1156,N_25038,N_29385);
and UO_1157 (O_1157,N_27319,N_27866);
and UO_1158 (O_1158,N_25711,N_25510);
and UO_1159 (O_1159,N_27098,N_29277);
nor UO_1160 (O_1160,N_26013,N_28234);
or UO_1161 (O_1161,N_27765,N_29463);
or UO_1162 (O_1162,N_28763,N_26319);
and UO_1163 (O_1163,N_28252,N_28643);
xor UO_1164 (O_1164,N_27871,N_25870);
nand UO_1165 (O_1165,N_28751,N_26896);
or UO_1166 (O_1166,N_27798,N_28330);
and UO_1167 (O_1167,N_28764,N_28231);
and UO_1168 (O_1168,N_26022,N_25958);
nor UO_1169 (O_1169,N_27612,N_28780);
nor UO_1170 (O_1170,N_29539,N_27677);
xor UO_1171 (O_1171,N_25592,N_27856);
nand UO_1172 (O_1172,N_28412,N_29335);
and UO_1173 (O_1173,N_28984,N_29683);
and UO_1174 (O_1174,N_29736,N_25746);
nand UO_1175 (O_1175,N_27981,N_29607);
nand UO_1176 (O_1176,N_29316,N_28734);
nand UO_1177 (O_1177,N_29006,N_25610);
nor UO_1178 (O_1178,N_25220,N_27228);
or UO_1179 (O_1179,N_29941,N_29933);
and UO_1180 (O_1180,N_25988,N_29490);
nand UO_1181 (O_1181,N_28574,N_28215);
xor UO_1182 (O_1182,N_29546,N_28109);
or UO_1183 (O_1183,N_28227,N_26733);
and UO_1184 (O_1184,N_28462,N_26411);
nor UO_1185 (O_1185,N_29144,N_25530);
nand UO_1186 (O_1186,N_27520,N_25456);
or UO_1187 (O_1187,N_28027,N_29065);
or UO_1188 (O_1188,N_27814,N_26699);
xnor UO_1189 (O_1189,N_27686,N_25127);
nor UO_1190 (O_1190,N_29268,N_28483);
or UO_1191 (O_1191,N_26919,N_25123);
or UO_1192 (O_1192,N_28489,N_27799);
or UO_1193 (O_1193,N_26689,N_27656);
and UO_1194 (O_1194,N_25212,N_26094);
xor UO_1195 (O_1195,N_25007,N_29484);
xor UO_1196 (O_1196,N_26063,N_26765);
nor UO_1197 (O_1197,N_25279,N_27014);
nand UO_1198 (O_1198,N_25587,N_28896);
or UO_1199 (O_1199,N_25843,N_25307);
xnor UO_1200 (O_1200,N_25172,N_25537);
nand UO_1201 (O_1201,N_27308,N_28458);
nor UO_1202 (O_1202,N_27299,N_29773);
nand UO_1203 (O_1203,N_25992,N_27010);
xnor UO_1204 (O_1204,N_25387,N_28894);
and UO_1205 (O_1205,N_27174,N_29402);
or UO_1206 (O_1206,N_25274,N_27905);
nor UO_1207 (O_1207,N_26373,N_26281);
or UO_1208 (O_1208,N_27136,N_28441);
nor UO_1209 (O_1209,N_29832,N_28552);
xnor UO_1210 (O_1210,N_27751,N_26462);
or UO_1211 (O_1211,N_25907,N_27154);
nand UO_1212 (O_1212,N_29365,N_26561);
nor UO_1213 (O_1213,N_27974,N_26116);
xor UO_1214 (O_1214,N_29697,N_25525);
or UO_1215 (O_1215,N_28841,N_29479);
nand UO_1216 (O_1216,N_29201,N_25651);
and UO_1217 (O_1217,N_26916,N_27467);
nand UO_1218 (O_1218,N_26182,N_27611);
or UO_1219 (O_1219,N_28703,N_25128);
and UO_1220 (O_1220,N_27535,N_26794);
nand UO_1221 (O_1221,N_26005,N_27828);
nor UO_1222 (O_1222,N_28600,N_27771);
or UO_1223 (O_1223,N_27243,N_25644);
nand UO_1224 (O_1224,N_26875,N_28053);
nand UO_1225 (O_1225,N_25818,N_29068);
nand UO_1226 (O_1226,N_25041,N_27891);
and UO_1227 (O_1227,N_27370,N_27658);
nor UO_1228 (O_1228,N_26236,N_28766);
and UO_1229 (O_1229,N_28141,N_26530);
and UO_1230 (O_1230,N_25257,N_27792);
and UO_1231 (O_1231,N_29999,N_29282);
nand UO_1232 (O_1232,N_26928,N_27436);
and UO_1233 (O_1233,N_27393,N_26257);
and UO_1234 (O_1234,N_27310,N_27631);
nand UO_1235 (O_1235,N_29621,N_26429);
nor UO_1236 (O_1236,N_28557,N_25604);
or UO_1237 (O_1237,N_29290,N_26595);
nor UO_1238 (O_1238,N_27352,N_27717);
and UO_1239 (O_1239,N_26284,N_27747);
and UO_1240 (O_1240,N_27274,N_26655);
and UO_1241 (O_1241,N_28022,N_26949);
or UO_1242 (O_1242,N_25070,N_27430);
and UO_1243 (O_1243,N_26062,N_27694);
and UO_1244 (O_1244,N_28187,N_28895);
xnor UO_1245 (O_1245,N_28581,N_26362);
or UO_1246 (O_1246,N_26258,N_27530);
or UO_1247 (O_1247,N_28664,N_26122);
and UO_1248 (O_1248,N_25620,N_26117);
nand UO_1249 (O_1249,N_29464,N_28336);
nor UO_1250 (O_1250,N_27005,N_29957);
and UO_1251 (O_1251,N_26451,N_27858);
or UO_1252 (O_1252,N_25248,N_28147);
nor UO_1253 (O_1253,N_25487,N_27926);
nor UO_1254 (O_1254,N_25258,N_26232);
nand UO_1255 (O_1255,N_27918,N_29810);
or UO_1256 (O_1256,N_29172,N_25538);
nor UO_1257 (O_1257,N_26084,N_27897);
or UO_1258 (O_1258,N_28318,N_25484);
or UO_1259 (O_1259,N_29620,N_27387);
and UO_1260 (O_1260,N_25887,N_26081);
xnor UO_1261 (O_1261,N_27292,N_29407);
xor UO_1262 (O_1262,N_29163,N_29209);
or UO_1263 (O_1263,N_27944,N_29510);
nor UO_1264 (O_1264,N_26809,N_27281);
nand UO_1265 (O_1265,N_27876,N_25216);
nand UO_1266 (O_1266,N_29536,N_26746);
nand UO_1267 (O_1267,N_29867,N_25998);
nor UO_1268 (O_1268,N_26439,N_28815);
and UO_1269 (O_1269,N_29981,N_27967);
xor UO_1270 (O_1270,N_28721,N_26158);
xnor UO_1271 (O_1271,N_25102,N_26328);
or UO_1272 (O_1272,N_29395,N_28220);
and UO_1273 (O_1273,N_28490,N_29885);
or UO_1274 (O_1274,N_25264,N_26888);
nor UO_1275 (O_1275,N_26534,N_27584);
and UO_1276 (O_1276,N_28539,N_29118);
nand UO_1277 (O_1277,N_26111,N_28754);
nor UO_1278 (O_1278,N_27202,N_27741);
and UO_1279 (O_1279,N_25136,N_28893);
or UO_1280 (O_1280,N_29148,N_25088);
nor UO_1281 (O_1281,N_28121,N_29345);
and UO_1282 (O_1282,N_28873,N_27809);
xor UO_1283 (O_1283,N_28057,N_25424);
or UO_1284 (O_1284,N_25577,N_27358);
or UO_1285 (O_1285,N_29859,N_27516);
nand UO_1286 (O_1286,N_27223,N_29159);
nand UO_1287 (O_1287,N_29775,N_25943);
nand UO_1288 (O_1288,N_25591,N_27924);
or UO_1289 (O_1289,N_27161,N_25724);
or UO_1290 (O_1290,N_25434,N_25003);
xnor UO_1291 (O_1291,N_26160,N_29905);
or UO_1292 (O_1292,N_25840,N_26571);
and UO_1293 (O_1293,N_28518,N_26403);
nand UO_1294 (O_1294,N_27041,N_26906);
nand UO_1295 (O_1295,N_27830,N_28117);
nor UO_1296 (O_1296,N_27112,N_28537);
nor UO_1297 (O_1297,N_29588,N_25314);
and UO_1298 (O_1298,N_27907,N_27532);
and UO_1299 (O_1299,N_25471,N_28757);
nand UO_1300 (O_1300,N_29455,N_25859);
nand UO_1301 (O_1301,N_27732,N_25984);
and UO_1302 (O_1302,N_26448,N_26788);
and UO_1303 (O_1303,N_26050,N_27636);
nand UO_1304 (O_1304,N_29158,N_26852);
or UO_1305 (O_1305,N_28413,N_29315);
nand UO_1306 (O_1306,N_26856,N_26139);
nand UO_1307 (O_1307,N_28047,N_29356);
nor UO_1308 (O_1308,N_29630,N_28446);
nand UO_1309 (O_1309,N_29046,N_26680);
or UO_1310 (O_1310,N_29664,N_26405);
nand UO_1311 (O_1311,N_28939,N_27195);
nand UO_1312 (O_1312,N_25999,N_28167);
and UO_1313 (O_1313,N_29390,N_25631);
nor UO_1314 (O_1314,N_27620,N_27948);
or UO_1315 (O_1315,N_29203,N_26181);
xor UO_1316 (O_1316,N_26662,N_26219);
or UO_1317 (O_1317,N_27688,N_27294);
nor UO_1318 (O_1318,N_28313,N_29524);
or UO_1319 (O_1319,N_25950,N_26496);
or UO_1320 (O_1320,N_25739,N_28753);
and UO_1321 (O_1321,N_28511,N_26422);
nand UO_1322 (O_1322,N_28010,N_29280);
or UO_1323 (O_1323,N_27494,N_29386);
and UO_1324 (O_1324,N_27696,N_29409);
or UO_1325 (O_1325,N_28066,N_28684);
nand UO_1326 (O_1326,N_27318,N_29185);
nand UO_1327 (O_1327,N_29275,N_29415);
nor UO_1328 (O_1328,N_27383,N_26316);
or UO_1329 (O_1329,N_27201,N_27108);
and UO_1330 (O_1330,N_25404,N_25492);
nand UO_1331 (O_1331,N_26621,N_28965);
nor UO_1332 (O_1332,N_29776,N_25465);
nand UO_1333 (O_1333,N_27058,N_25790);
nor UO_1334 (O_1334,N_26521,N_29537);
nand UO_1335 (O_1335,N_25242,N_28680);
nor UO_1336 (O_1336,N_25134,N_29233);
nand UO_1337 (O_1337,N_25672,N_27515);
or UO_1338 (O_1338,N_27062,N_25977);
xnor UO_1339 (O_1339,N_27399,N_25272);
nor UO_1340 (O_1340,N_28192,N_27803);
nand UO_1341 (O_1341,N_28379,N_28470);
nor UO_1342 (O_1342,N_27887,N_26153);
and UO_1343 (O_1343,N_28865,N_28455);
nor UO_1344 (O_1344,N_27922,N_29284);
and UO_1345 (O_1345,N_26705,N_29653);
xnor UO_1346 (O_1346,N_29442,N_29527);
nor UO_1347 (O_1347,N_26979,N_26161);
nand UO_1348 (O_1348,N_25399,N_29361);
or UO_1349 (O_1349,N_25678,N_29670);
nor UO_1350 (O_1350,N_25039,N_26671);
xor UO_1351 (O_1351,N_29633,N_29526);
nor UO_1352 (O_1352,N_28298,N_28497);
xnor UO_1353 (O_1353,N_29815,N_25423);
and UO_1354 (O_1354,N_26985,N_25035);
or UO_1355 (O_1355,N_26333,N_25031);
or UO_1356 (O_1356,N_26028,N_27355);
nand UO_1357 (O_1357,N_29522,N_27470);
and UO_1358 (O_1358,N_25073,N_29468);
or UO_1359 (O_1359,N_26523,N_28381);
nor UO_1360 (O_1360,N_28782,N_28062);
and UO_1361 (O_1361,N_29903,N_29756);
nor UO_1362 (O_1362,N_27375,N_25872);
nand UO_1363 (O_1363,N_27994,N_27187);
nor UO_1364 (O_1364,N_28904,N_26494);
nor UO_1365 (O_1365,N_26808,N_28361);
or UO_1366 (O_1366,N_27448,N_26192);
nor UO_1367 (O_1367,N_29257,N_29908);
or UO_1368 (O_1368,N_25064,N_27624);
nand UO_1369 (O_1369,N_25831,N_28221);
or UO_1370 (O_1370,N_26528,N_28207);
nor UO_1371 (O_1371,N_26861,N_26121);
and UO_1372 (O_1372,N_28980,N_28502);
nand UO_1373 (O_1373,N_25543,N_25524);
and UO_1374 (O_1374,N_26307,N_25751);
nor UO_1375 (O_1375,N_28315,N_26224);
or UO_1376 (O_1376,N_27775,N_29668);
nand UO_1377 (O_1377,N_26204,N_28233);
nor UO_1378 (O_1378,N_26272,N_26201);
and UO_1379 (O_1379,N_27284,N_27316);
xor UO_1380 (O_1380,N_28319,N_27729);
or UO_1381 (O_1381,N_26298,N_27416);
nor UO_1382 (O_1382,N_25342,N_25559);
or UO_1383 (O_1383,N_28785,N_28311);
and UO_1384 (O_1384,N_26098,N_27555);
or UO_1385 (O_1385,N_28208,N_25973);
nand UO_1386 (O_1386,N_27990,N_26775);
or UO_1387 (O_1387,N_28243,N_28627);
and UO_1388 (O_1388,N_25229,N_25597);
nand UO_1389 (O_1389,N_28791,N_28962);
nand UO_1390 (O_1390,N_29600,N_25328);
and UO_1391 (O_1391,N_28015,N_28937);
or UO_1392 (O_1392,N_27801,N_29189);
or UO_1393 (O_1393,N_27728,N_29263);
and UO_1394 (O_1394,N_25313,N_25481);
or UO_1395 (O_1395,N_25063,N_28977);
nor UO_1396 (O_1396,N_28176,N_26503);
and UO_1397 (O_1397,N_25704,N_28091);
nand UO_1398 (O_1398,N_29780,N_28919);
and UO_1399 (O_1399,N_29504,N_28848);
or UO_1400 (O_1400,N_27844,N_29856);
xor UO_1401 (O_1401,N_27587,N_29142);
and UO_1402 (O_1402,N_28273,N_27471);
and UO_1403 (O_1403,N_29279,N_26790);
nor UO_1404 (O_1404,N_27726,N_29821);
nor UO_1405 (O_1405,N_25357,N_26821);
or UO_1406 (O_1406,N_25068,N_26786);
or UO_1407 (O_1407,N_27923,N_29830);
and UO_1408 (O_1408,N_28645,N_28648);
or UO_1409 (O_1409,N_27985,N_27341);
nor UO_1410 (O_1410,N_26669,N_29584);
nor UO_1411 (O_1411,N_28205,N_26866);
nand UO_1412 (O_1412,N_25025,N_29801);
nand UO_1413 (O_1413,N_28382,N_27357);
nor UO_1414 (O_1414,N_27896,N_25261);
or UO_1415 (O_1415,N_26750,N_27562);
nand UO_1416 (O_1416,N_27288,N_27237);
nand UO_1417 (O_1417,N_27557,N_29907);
nor UO_1418 (O_1418,N_28181,N_29082);
or UO_1419 (O_1419,N_29919,N_27481);
or UO_1420 (O_1420,N_29800,N_29967);
and UO_1421 (O_1421,N_26897,N_26041);
xor UO_1422 (O_1422,N_29300,N_27522);
nor UO_1423 (O_1423,N_26509,N_26975);
xor UO_1424 (O_1424,N_28292,N_26207);
or UO_1425 (O_1425,N_29613,N_28112);
or UO_1426 (O_1426,N_27782,N_27454);
and UO_1427 (O_1427,N_28989,N_27784);
or UO_1428 (O_1428,N_26581,N_29370);
or UO_1429 (O_1429,N_25968,N_27424);
or UO_1430 (O_1430,N_26290,N_27513);
or UO_1431 (O_1431,N_26303,N_26730);
and UO_1432 (O_1432,N_26564,N_29408);
nand UO_1433 (O_1433,N_29500,N_27013);
xnor UO_1434 (O_1434,N_25245,N_29564);
nand UO_1435 (O_1435,N_27048,N_28587);
or UO_1436 (O_1436,N_25590,N_27598);
nand UO_1437 (O_1437,N_28516,N_25494);
and UO_1438 (O_1438,N_26960,N_29077);
or UO_1439 (O_1439,N_28193,N_28358);
nand UO_1440 (O_1440,N_26820,N_27778);
or UO_1441 (O_1441,N_29033,N_28399);
nor UO_1442 (O_1442,N_29858,N_29044);
nand UO_1443 (O_1443,N_25558,N_29899);
nor UO_1444 (O_1444,N_29092,N_29071);
or UO_1445 (O_1445,N_28020,N_25900);
or UO_1446 (O_1446,N_25329,N_25129);
nand UO_1447 (O_1447,N_25297,N_29658);
and UO_1448 (O_1448,N_27851,N_25496);
nand UO_1449 (O_1449,N_29961,N_29982);
or UO_1450 (O_1450,N_26742,N_29608);
nand UO_1451 (O_1451,N_25074,N_28452);
or UO_1452 (O_1452,N_26862,N_29166);
nor UO_1453 (O_1453,N_25681,N_27489);
nand UO_1454 (O_1454,N_26464,N_28947);
and UO_1455 (O_1455,N_29238,N_29339);
and UO_1456 (O_1456,N_29894,N_29286);
or UO_1457 (O_1457,N_26154,N_26665);
nor UO_1458 (O_1458,N_28521,N_28039);
and UO_1459 (O_1459,N_28456,N_25017);
nand UO_1460 (O_1460,N_26506,N_29096);
nand UO_1461 (O_1461,N_28928,N_25367);
and UO_1462 (O_1462,N_26993,N_26757);
xor UO_1463 (O_1463,N_28626,N_29843);
or UO_1464 (O_1464,N_28713,N_28767);
nor UO_1465 (O_1465,N_29717,N_27317);
xnor UO_1466 (O_1466,N_28380,N_27940);
xnor UO_1467 (O_1467,N_28346,N_27049);
and UO_1468 (O_1468,N_26468,N_26939);
nand UO_1469 (O_1469,N_26593,N_25319);
nor UO_1470 (O_1470,N_26546,N_29542);
xnor UO_1471 (O_1471,N_26508,N_28917);
or UO_1472 (O_1472,N_27833,N_26254);
and UO_1473 (O_1473,N_27325,N_29993);
xnor UO_1474 (O_1474,N_25236,N_28686);
and UO_1475 (O_1475,N_27714,N_25183);
nand UO_1476 (O_1476,N_28347,N_25371);
nor UO_1477 (O_1477,N_26857,N_27501);
nor UO_1478 (O_1478,N_29229,N_26887);
nand UO_1479 (O_1479,N_29676,N_25475);
or UO_1480 (O_1480,N_29453,N_27173);
nor UO_1481 (O_1481,N_28059,N_25602);
nand UO_1482 (O_1482,N_27768,N_27885);
nor UO_1483 (O_1483,N_27536,N_26045);
nor UO_1484 (O_1484,N_27715,N_26825);
and UO_1485 (O_1485,N_29829,N_28642);
or UO_1486 (O_1486,N_29487,N_29816);
and UO_1487 (O_1487,N_28025,N_29287);
and UO_1488 (O_1488,N_27175,N_28705);
nand UO_1489 (O_1489,N_29254,N_25333);
nor UO_1490 (O_1490,N_25989,N_25400);
nor UO_1491 (O_1491,N_25121,N_25869);
nor UO_1492 (O_1492,N_26199,N_26625);
xor UO_1493 (O_1493,N_27911,N_28855);
and UO_1494 (O_1494,N_29569,N_26393);
or UO_1495 (O_1495,N_27116,N_25821);
nand UO_1496 (O_1496,N_27479,N_29844);
and UO_1497 (O_1497,N_26563,N_26348);
nor UO_1498 (O_1498,N_27838,N_26268);
and UO_1499 (O_1499,N_28650,N_28130);
and UO_1500 (O_1500,N_26882,N_28583);
xnor UO_1501 (O_1501,N_27649,N_27032);
nand UO_1502 (O_1502,N_28891,N_29272);
or UO_1503 (O_1503,N_26412,N_29648);
nor UO_1504 (O_1504,N_25206,N_25459);
nor UO_1505 (O_1505,N_28930,N_28924);
nor UO_1506 (O_1506,N_26696,N_28857);
nor UO_1507 (O_1507,N_27577,N_27537);
and UO_1508 (O_1508,N_28143,N_28761);
or UO_1509 (O_1509,N_26196,N_26748);
and UO_1510 (O_1510,N_25042,N_27639);
nand UO_1511 (O_1511,N_27478,N_27450);
nor UO_1512 (O_1512,N_27579,N_25043);
nor UO_1513 (O_1513,N_25125,N_26844);
and UO_1514 (O_1514,N_26102,N_29939);
and UO_1515 (O_1515,N_25345,N_25697);
nand UO_1516 (O_1516,N_26035,N_26673);
xnor UO_1517 (O_1517,N_26681,N_26431);
or UO_1518 (O_1518,N_25727,N_28108);
or UO_1519 (O_1519,N_28026,N_27916);
nor UO_1520 (O_1520,N_27843,N_29481);
nor UO_1521 (O_1521,N_28619,N_26335);
or UO_1522 (O_1522,N_27580,N_28122);
xor UO_1523 (O_1523,N_27680,N_25163);
or UO_1524 (O_1524,N_28709,N_28881);
and UO_1525 (O_1525,N_29920,N_26778);
xnor UO_1526 (O_1526,N_26597,N_29404);
xor UO_1527 (O_1527,N_26191,N_29000);
nor UO_1528 (O_1528,N_29380,N_26167);
nand UO_1529 (O_1529,N_27348,N_29722);
or UO_1530 (O_1530,N_26702,N_27003);
or UO_1531 (O_1531,N_29695,N_26179);
xnor UO_1532 (O_1532,N_28633,N_25090);
or UO_1533 (O_1533,N_26314,N_25416);
nand UO_1534 (O_1534,N_27615,N_28519);
nand UO_1535 (O_1535,N_29208,N_29053);
nor UO_1536 (O_1536,N_26216,N_26724);
or UO_1537 (O_1537,N_26359,N_25071);
nand UO_1538 (O_1538,N_29513,N_27186);
nor UO_1539 (O_1539,N_26065,N_29120);
nor UO_1540 (O_1540,N_25447,N_26324);
nand UO_1541 (O_1541,N_26755,N_25195);
and UO_1542 (O_1542,N_28566,N_25217);
or UO_1543 (O_1543,N_29672,N_28408);
or UO_1544 (O_1544,N_28306,N_27829);
nor UO_1545 (O_1545,N_28011,N_27184);
xnor UO_1546 (O_1546,N_29431,N_26151);
and UO_1547 (O_1547,N_28665,N_25111);
nor UO_1548 (O_1548,N_25040,N_27490);
nor UO_1549 (O_1549,N_26971,N_27939);
or UO_1550 (O_1550,N_27339,N_29016);
and UO_1551 (O_1551,N_25567,N_25491);
and UO_1552 (O_1552,N_25093,N_25298);
and UO_1553 (O_1553,N_27016,N_29838);
nor UO_1554 (O_1554,N_29133,N_26320);
nand UO_1555 (O_1555,N_28617,N_25380);
xnor UO_1556 (O_1556,N_28994,N_27403);
or UO_1557 (O_1557,N_28036,N_25601);
nand UO_1558 (O_1558,N_28818,N_27241);
and UO_1559 (O_1559,N_29853,N_29614);
or UO_1560 (O_1560,N_29099,N_27979);
nand UO_1561 (O_1561,N_29696,N_25321);
xnor UO_1562 (O_1562,N_25067,N_25680);
nand UO_1563 (O_1563,N_25863,N_25165);
or UO_1564 (O_1564,N_28595,N_28133);
nand UO_1565 (O_1565,N_25777,N_29879);
or UO_1566 (O_1566,N_26782,N_29533);
or UO_1567 (O_1567,N_26622,N_26100);
nor UO_1568 (O_1568,N_27661,N_29938);
or UO_1569 (O_1569,N_28425,N_25926);
nand UO_1570 (O_1570,N_25614,N_27901);
and UO_1571 (O_1571,N_25642,N_25623);
and UO_1572 (O_1572,N_25096,N_27480);
and UO_1573 (O_1573,N_27469,N_25902);
and UO_1574 (O_1574,N_29741,N_26589);
or UO_1575 (O_1575,N_26410,N_27007);
nand UO_1576 (O_1576,N_28929,N_28654);
and UO_1577 (O_1577,N_29403,N_25188);
nand UO_1578 (O_1578,N_26590,N_26997);
xor UO_1579 (O_1579,N_27239,N_27992);
nand UO_1580 (O_1580,N_28500,N_28149);
or UO_1581 (O_1581,N_29273,N_26698);
or UO_1582 (O_1582,N_26533,N_28640);
nor UO_1583 (O_1583,N_27446,N_29824);
nand UO_1584 (O_1584,N_26704,N_25479);
and UO_1585 (O_1585,N_26926,N_29198);
xor UO_1586 (O_1586,N_26425,N_25917);
nand UO_1587 (O_1587,N_26758,N_27899);
nor UO_1588 (O_1588,N_27875,N_25256);
nand UO_1589 (O_1589,N_27426,N_25635);
nor UO_1590 (O_1590,N_26804,N_25716);
and UO_1591 (O_1591,N_26407,N_27153);
and UO_1592 (O_1592,N_27314,N_27162);
nor UO_1593 (O_1593,N_29121,N_26256);
nor UO_1594 (O_1594,N_26889,N_27461);
and UO_1595 (O_1595,N_25485,N_27235);
nand UO_1596 (O_1596,N_29299,N_25885);
xnor UO_1597 (O_1597,N_26460,N_26241);
xor UO_1598 (O_1598,N_26060,N_25909);
nand UO_1599 (O_1599,N_28492,N_28291);
nor UO_1600 (O_1600,N_29707,N_29958);
or UO_1601 (O_1601,N_28428,N_26527);
nand UO_1602 (O_1602,N_25341,N_25477);
or UO_1603 (O_1603,N_26535,N_28476);
nand UO_1604 (O_1604,N_26878,N_25019);
nand UO_1605 (O_1605,N_26210,N_28864);
or UO_1606 (O_1606,N_27256,N_28058);
nand UO_1607 (O_1607,N_26907,N_25653);
or UO_1608 (O_1608,N_29682,N_29215);
or UO_1609 (O_1609,N_27040,N_25168);
or UO_1610 (O_1610,N_29805,N_25233);
nor UO_1611 (O_1611,N_25373,N_29705);
nand UO_1612 (O_1612,N_26002,N_27551);
or UO_1613 (O_1613,N_25861,N_29837);
nand UO_1614 (O_1614,N_27589,N_27526);
nand UO_1615 (O_1615,N_26071,N_27204);
or UO_1616 (O_1616,N_28569,N_28019);
nand UO_1617 (O_1617,N_25061,N_27762);
xnor UO_1618 (O_1618,N_27692,N_26106);
and UO_1619 (O_1619,N_27323,N_27453);
nand UO_1620 (O_1620,N_28926,N_29294);
and UO_1621 (O_1621,N_26019,N_28001);
or UO_1622 (O_1622,N_25429,N_26061);
nor UO_1623 (O_1623,N_25142,N_26383);
nor UO_1624 (O_1624,N_28060,N_27183);
and UO_1625 (O_1625,N_28037,N_27978);
and UO_1626 (O_1626,N_27061,N_26297);
and UO_1627 (O_1627,N_27222,N_25684);
nand UO_1628 (O_1628,N_28488,N_25871);
xor UO_1629 (O_1629,N_25693,N_27051);
nand UO_1630 (O_1630,N_25731,N_28230);
nand UO_1631 (O_1631,N_26912,N_26935);
nand UO_1632 (O_1632,N_25460,N_27397);
or UO_1633 (O_1633,N_25883,N_25563);
and UO_1634 (O_1634,N_27220,N_28825);
xor UO_1635 (O_1635,N_28331,N_26086);
xor UO_1636 (O_1636,N_29196,N_26068);
nand UO_1637 (O_1637,N_27780,N_25536);
nand UO_1638 (O_1638,N_29250,N_26385);
nor UO_1639 (O_1639,N_27699,N_27807);
nand UO_1640 (O_1640,N_28657,N_28128);
or UO_1641 (O_1641,N_26352,N_26542);
and UO_1642 (O_1642,N_28210,N_29871);
and UO_1643 (O_1643,N_25486,N_25807);
nor UO_1644 (O_1644,N_29375,N_29137);
or UO_1645 (O_1645,N_25277,N_27943);
nor UO_1646 (O_1646,N_27248,N_29984);
nor UO_1647 (O_1647,N_29563,N_28556);
nor UO_1648 (O_1648,N_27675,N_28051);
xnor UO_1649 (O_1649,N_28416,N_25987);
or UO_1650 (O_1650,N_25985,N_29155);
and UO_1651 (O_1651,N_28950,N_28945);
or UO_1652 (O_1652,N_27722,N_27629);
nand UO_1653 (O_1653,N_29459,N_26317);
or UO_1654 (O_1654,N_26427,N_27344);
xor UO_1655 (O_1655,N_25959,N_26522);
and UO_1656 (O_1656,N_29883,N_29192);
or UO_1657 (O_1657,N_29107,N_29086);
and UO_1658 (O_1658,N_29055,N_26559);
nor UO_1659 (O_1659,N_28034,N_28159);
nor UO_1660 (O_1660,N_25853,N_29170);
nor UO_1661 (O_1661,N_25584,N_28802);
nor UO_1662 (O_1662,N_27296,N_27835);
and UO_1663 (O_1663,N_26531,N_29739);
xor UO_1664 (O_1664,N_25478,N_27850);
or UO_1665 (O_1665,N_26295,N_29802);
and UO_1666 (O_1666,N_29986,N_27773);
nor UO_1667 (O_1667,N_25057,N_29869);
nor UO_1668 (O_1668,N_26847,N_27302);
and UO_1669 (O_1669,N_29364,N_27413);
nor UO_1670 (O_1670,N_28852,N_26409);
or UO_1671 (O_1671,N_25356,N_28747);
nor UO_1672 (O_1672,N_26424,N_26423);
and UO_1673 (O_1673,N_27774,N_25829);
or UO_1674 (O_1674,N_29434,N_25353);
or UO_1675 (O_1675,N_29122,N_25173);
nand UO_1676 (O_1676,N_26784,N_26994);
xor UO_1677 (O_1677,N_27492,N_28171);
or UO_1678 (O_1678,N_29779,N_26149);
or UO_1679 (O_1679,N_26248,N_28730);
and UO_1680 (O_1680,N_26937,N_25607);
or UO_1681 (O_1681,N_27998,N_26504);
nor UO_1682 (O_1682,N_27350,N_29578);
and UO_1683 (O_1683,N_25619,N_28351);
or UO_1684 (O_1684,N_27845,N_27681);
or UO_1685 (O_1685,N_29762,N_26032);
or UO_1686 (O_1686,N_25349,N_29200);
nor UO_1687 (O_1687,N_26524,N_26879);
nor UO_1688 (O_1688,N_29918,N_25621);
nor UO_1689 (O_1689,N_27345,N_28892);
and UO_1690 (O_1690,N_27855,N_25527);
nor UO_1691 (O_1691,N_29944,N_29477);
and UO_1692 (O_1692,N_29305,N_25075);
and UO_1693 (O_1693,N_27756,N_29804);
and UO_1694 (O_1694,N_29228,N_28608);
nand UO_1695 (O_1695,N_28308,N_26243);
nand UO_1696 (O_1696,N_25946,N_29352);
nor UO_1697 (O_1697,N_25020,N_27865);
xor UO_1698 (O_1698,N_28836,N_26413);
or UO_1699 (O_1699,N_27215,N_28486);
or UO_1700 (O_1700,N_28068,N_29729);
nor UO_1701 (O_1701,N_27194,N_25738);
or UO_1702 (O_1702,N_29681,N_29840);
or UO_1703 (O_1703,N_26109,N_25320);
nand UO_1704 (O_1704,N_27933,N_26645);
nor UO_1705 (O_1705,N_25358,N_26093);
nor UO_1706 (O_1706,N_27057,N_26057);
xor UO_1707 (O_1707,N_28161,N_29545);
nor UO_1708 (O_1708,N_29177,N_28478);
or UO_1709 (O_1709,N_25838,N_26234);
or UO_1710 (O_1710,N_25202,N_28529);
xnor UO_1711 (O_1711,N_26807,N_29550);
and UO_1712 (O_1712,N_25474,N_28050);
xnor UO_1713 (O_1713,N_28997,N_28196);
nor UO_1714 (O_1714,N_26006,N_28636);
nand UO_1715 (O_1715,N_29904,N_27101);
xnor UO_1716 (O_1716,N_27892,N_27931);
nor UO_1717 (O_1717,N_28182,N_25361);
or UO_1718 (O_1718,N_25523,N_27458);
and UO_1719 (O_1719,N_26208,N_26358);
or UO_1720 (O_1720,N_27004,N_29288);
nand UO_1721 (O_1721,N_29799,N_27919);
nor UO_1722 (O_1722,N_29436,N_28244);
nor UO_1723 (O_1723,N_28454,N_28334);
and UO_1724 (O_1724,N_28695,N_28783);
nand UO_1725 (O_1725,N_28874,N_25164);
nor UO_1726 (O_1726,N_25819,N_27432);
nand UO_1727 (O_1727,N_27585,N_25290);
nor UO_1728 (O_1728,N_26034,N_27038);
and UO_1729 (O_1729,N_28354,N_26288);
and UO_1730 (O_1730,N_29937,N_25671);
nand UO_1731 (O_1731,N_26876,N_25211);
nand UO_1732 (O_1732,N_27977,N_27668);
nor UO_1733 (O_1733,N_28127,N_29787);
xor UO_1734 (O_1734,N_27628,N_27085);
nand UO_1735 (O_1735,N_29324,N_26614);
nor UO_1736 (O_1736,N_25618,N_25808);
or UO_1737 (O_1737,N_25695,N_28395);
nor UO_1738 (O_1738,N_26639,N_28043);
nor UO_1739 (O_1739,N_29970,N_26226);
and UO_1740 (O_1740,N_25337,N_29783);
and UO_1741 (O_1741,N_25181,N_26623);
or UO_1742 (O_1742,N_27938,N_28178);
nor UO_1743 (O_1743,N_28698,N_29423);
or UO_1744 (O_1744,N_26842,N_25008);
or UO_1745 (O_1745,N_28809,N_26629);
and UO_1746 (O_1746,N_25710,N_26840);
xnor UO_1747 (O_1747,N_27036,N_25534);
nand UO_1748 (O_1748,N_26678,N_28279);
and UO_1749 (O_1749,N_29978,N_27046);
or UO_1750 (O_1750,N_28943,N_29991);
and UO_1751 (O_1751,N_25728,N_25700);
nand UO_1752 (O_1752,N_27230,N_26014);
or UO_1753 (O_1753,N_29432,N_25047);
nor UO_1754 (O_1754,N_26083,N_29972);
or UO_1755 (O_1755,N_27388,N_28733);
nor UO_1756 (O_1756,N_25289,N_28671);
and UO_1757 (O_1757,N_25736,N_29868);
or UO_1758 (O_1758,N_29088,N_26813);
and UO_1759 (O_1759,N_28834,N_26264);
or UO_1760 (O_1760,N_26325,N_25932);
and UO_1761 (O_1761,N_28179,N_27785);
xnor UO_1762 (O_1762,N_25374,N_26127);
nor UO_1763 (O_1763,N_29051,N_27854);
nor UO_1764 (O_1764,N_28983,N_26092);
nor UO_1765 (O_1765,N_26064,N_26510);
nor UO_1766 (O_1766,N_29823,N_25801);
or UO_1767 (O_1767,N_26830,N_26479);
nand UO_1768 (O_1768,N_29916,N_27434);
nand UO_1769 (O_1769,N_29713,N_26354);
nand UO_1770 (O_1770,N_27263,N_29235);
or UO_1771 (O_1771,N_27250,N_26467);
nand UO_1772 (O_1772,N_28603,N_25259);
nand UO_1773 (O_1773,N_28993,N_27491);
nor UO_1774 (O_1774,N_26433,N_27086);
or UO_1775 (O_1775,N_29105,N_26058);
or UO_1776 (O_1776,N_29406,N_25166);
or UO_1777 (O_1777,N_26717,N_27804);
nand UO_1778 (O_1778,N_27813,N_26277);
nor UO_1779 (O_1779,N_29841,N_27012);
or UO_1780 (O_1780,N_26173,N_29979);
or UO_1781 (O_1781,N_29699,N_27151);
or UO_1782 (O_1782,N_27590,N_27713);
nand UO_1783 (O_1783,N_27152,N_25827);
nor UO_1784 (O_1784,N_28277,N_25162);
nor UO_1785 (O_1785,N_26246,N_25803);
or UO_1786 (O_1786,N_27205,N_28028);
or UO_1787 (O_1787,N_25381,N_29880);
or UO_1788 (O_1788,N_28638,N_27247);
or UO_1789 (O_1789,N_25666,N_29447);
and UO_1790 (O_1790,N_25414,N_27882);
xor UO_1791 (O_1791,N_29116,N_25881);
and UO_1792 (O_1792,N_26419,N_27333);
nor UO_1793 (O_1793,N_25441,N_26756);
and UO_1794 (O_1794,N_25762,N_26163);
nand UO_1795 (O_1795,N_26384,N_27447);
nor UO_1796 (O_1796,N_26838,N_29333);
xnor UO_1797 (O_1797,N_29388,N_27231);
nand UO_1798 (O_1798,N_29612,N_29384);
nor UO_1799 (O_1799,N_29657,N_26632);
xor UO_1800 (O_1800,N_27468,N_27475);
and UO_1801 (O_1801,N_28228,N_27991);
and UO_1802 (O_1802,N_28678,N_27107);
nand UO_1803 (O_1803,N_25549,N_28796);
and UO_1804 (O_1804,N_29574,N_29331);
xor UO_1805 (O_1805,N_28906,N_27037);
and UO_1806 (O_1806,N_25956,N_27141);
or UO_1807 (O_1807,N_29581,N_26741);
or UO_1808 (O_1808,N_25512,N_28014);
nand UO_1809 (O_1809,N_28677,N_28061);
nor UO_1810 (O_1810,N_28113,N_25782);
and UO_1811 (O_1811,N_26858,N_29478);
and UO_1812 (O_1812,N_25284,N_28655);
or UO_1813 (O_1813,N_25343,N_25407);
nand UO_1814 (O_1814,N_29549,N_29075);
and UO_1815 (O_1815,N_25350,N_25904);
xnor UO_1816 (O_1816,N_27076,N_28716);
nor UO_1817 (O_1817,N_29112,N_25542);
or UO_1818 (O_1818,N_28942,N_27373);
xnor UO_1819 (O_1819,N_27252,N_28995);
or UO_1820 (O_1820,N_27128,N_26962);
xnor UO_1821 (O_1821,N_27840,N_28935);
or UO_1822 (O_1822,N_25021,N_28564);
nand UO_1823 (O_1823,N_29195,N_29494);
or UO_1824 (O_1824,N_26884,N_26829);
and UO_1825 (O_1825,N_25661,N_29661);
nor UO_1826 (O_1826,N_25029,N_26166);
nor UO_1827 (O_1827,N_27496,N_27031);
nor UO_1828 (O_1828,N_29242,N_25612);
or UO_1829 (O_1829,N_27750,N_29809);
or UO_1830 (O_1830,N_29700,N_27021);
nor UO_1831 (O_1831,N_29424,N_26183);
xor UO_1832 (O_1832,N_29037,N_28443);
xor UO_1833 (O_1833,N_25867,N_28224);
nor UO_1834 (O_1834,N_27509,N_28835);
and UO_1835 (O_1835,N_27582,N_28191);
nand UO_1836 (O_1836,N_29609,N_25114);
and UO_1837 (O_1837,N_25055,N_25539);
nor UO_1838 (O_1838,N_25648,N_27880);
or UO_1839 (O_1839,N_25625,N_27145);
and UO_1840 (O_1840,N_27249,N_29072);
and UO_1841 (O_1841,N_25785,N_26719);
and UO_1842 (O_1842,N_26417,N_25335);
nor UO_1843 (O_1843,N_25847,N_28225);
nand UO_1844 (O_1844,N_25993,N_29712);
xnor UO_1845 (O_1845,N_28851,N_29589);
nor UO_1846 (O_1846,N_29554,N_25806);
nand UO_1847 (O_1847,N_25767,N_26732);
or UO_1848 (O_1848,N_28077,N_26262);
and UO_1849 (O_1849,N_29379,N_25141);
or UO_1850 (O_1850,N_27825,N_29665);
and UO_1851 (O_1851,N_26657,N_27421);
or UO_1852 (O_1852,N_28849,N_26837);
or UO_1853 (O_1853,N_28084,N_28976);
nor UO_1854 (O_1854,N_29926,N_26954);
and UO_1855 (O_1855,N_29428,N_26004);
nand UO_1856 (O_1856,N_25225,N_26587);
and UO_1857 (O_1857,N_25837,N_28759);
and UO_1858 (O_1858,N_25647,N_28790);
nor UO_1859 (O_1859,N_29709,N_25262);
nand UO_1860 (O_1860,N_28858,N_29960);
and UO_1861 (O_1861,N_28833,N_27906);
nor UO_1862 (O_1862,N_29191,N_27460);
nor UO_1863 (O_1863,N_27755,N_25224);
nand UO_1864 (O_1864,N_25443,N_28363);
nand UO_1865 (O_1865,N_28107,N_27042);
or UO_1866 (O_1866,N_29725,N_27808);
nand UO_1867 (O_1867,N_28180,N_27211);
or UO_1868 (O_1868,N_29347,N_28293);
and UO_1869 (O_1869,N_25715,N_27258);
nor UO_1870 (O_1870,N_29231,N_29061);
nor UO_1871 (O_1871,N_25082,N_25963);
nand UO_1872 (O_1872,N_27017,N_29864);
or UO_1873 (O_1873,N_26822,N_26398);
nor UO_1874 (O_1874,N_26683,N_28338);
nor UO_1875 (O_1875,N_25639,N_28206);
or UO_1876 (O_1876,N_29685,N_26077);
and UO_1877 (O_1877,N_28982,N_28482);
xnor UO_1878 (O_1878,N_29796,N_27960);
or UO_1879 (O_1879,N_28173,N_28656);
or UO_1880 (O_1880,N_27092,N_27539);
xor UO_1881 (O_1881,N_25683,N_25930);
nor UO_1882 (O_1882,N_29199,N_26321);
nand UO_1883 (O_1883,N_25240,N_26376);
nor UO_1884 (O_1884,N_27894,N_25966);
nand UO_1885 (O_1885,N_28978,N_28675);
nand UO_1886 (O_1886,N_28553,N_25086);
and UO_1887 (O_1887,N_29825,N_28668);
or UO_1888 (O_1888,N_27279,N_26606);
nand UO_1889 (O_1889,N_27483,N_28165);
xnor UO_1890 (O_1890,N_29063,N_28290);
nand UO_1891 (O_1891,N_28251,N_26941);
and UO_1892 (O_1892,N_28158,N_25412);
or UO_1893 (O_1893,N_29547,N_28515);
nand UO_1894 (O_1894,N_26312,N_29389);
and UO_1895 (O_1895,N_28637,N_27633);
or UO_1896 (O_1896,N_29770,N_28479);
and UO_1897 (O_1897,N_26549,N_25246);
nand UO_1898 (O_1898,N_29931,N_26560);
nor UO_1899 (O_1899,N_27666,N_26016);
nand UO_1900 (O_1900,N_28824,N_26895);
or UO_1901 (O_1901,N_27102,N_25390);
nor UO_1902 (O_1902,N_27168,N_25083);
and UO_1903 (O_1903,N_25851,N_25427);
nor UO_1904 (O_1904,N_28447,N_26357);
nor UO_1905 (O_1905,N_26618,N_27970);
nor UO_1906 (O_1906,N_25405,N_29168);
and UO_1907 (O_1907,N_27691,N_26617);
nand UO_1908 (O_1908,N_26793,N_29686);
nand UO_1909 (O_1909,N_25270,N_26637);
and UO_1910 (O_1910,N_25436,N_26056);
nand UO_1911 (O_1911,N_29808,N_27987);
or UO_1912 (O_1912,N_25628,N_28571);
nand UO_1913 (O_1913,N_28296,N_28708);
nor UO_1914 (O_1914,N_27528,N_26443);
and UO_1915 (O_1915,N_28639,N_27485);
and UO_1916 (O_1916,N_25144,N_25965);
nor UO_1917 (O_1917,N_28268,N_25786);
nand UO_1918 (O_1918,N_26910,N_27059);
and UO_1919 (O_1919,N_29935,N_27815);
nand UO_1920 (O_1920,N_27538,N_26089);
nand UO_1921 (O_1921,N_28137,N_26817);
or UO_1922 (O_1922,N_25192,N_26026);
xor UO_1923 (O_1923,N_25215,N_26011);
nand UO_1924 (O_1924,N_26131,N_29445);
and UO_1925 (O_1925,N_25467,N_28872);
nand UO_1926 (O_1926,N_28120,N_28726);
or UO_1927 (O_1927,N_25201,N_27165);
nor UO_1928 (O_1928,N_27072,N_25839);
nand UO_1929 (O_1929,N_29132,N_29746);
nor UO_1930 (O_1930,N_25051,N_27842);
and UO_1931 (O_1931,N_28474,N_26178);
nor UO_1932 (O_1932,N_28475,N_27000);
and UO_1933 (O_1933,N_25445,N_25501);
nand UO_1934 (O_1934,N_27508,N_29806);
nor UO_1935 (O_1935,N_28866,N_28267);
nor UO_1936 (O_1936,N_25617,N_26475);
or UO_1937 (O_1937,N_27812,N_26725);
nor UO_1938 (O_1938,N_27561,N_27208);
nor UO_1939 (O_1939,N_26989,N_25458);
or UO_1940 (O_1940,N_29391,N_25238);
or UO_1941 (O_1941,N_27180,N_27634);
nor UO_1942 (O_1942,N_26275,N_27965);
and UO_1943 (O_1943,N_26833,N_28031);
nand UO_1944 (O_1944,N_27452,N_27088);
and UO_1945 (O_1945,N_25750,N_25239);
and UO_1946 (O_1946,N_29060,N_28732);
and UO_1947 (O_1947,N_29483,N_28365);
nand UO_1948 (O_1948,N_25218,N_26686);
nand UO_1949 (O_1949,N_29430,N_28727);
nand UO_1950 (O_1950,N_29413,N_26541);
nor UO_1951 (O_1951,N_26693,N_28323);
xor UO_1952 (O_1952,N_28737,N_28256);
xor UO_1953 (O_1953,N_27759,N_29715);
and UO_1954 (O_1954,N_29422,N_26646);
nor UO_1955 (O_1955,N_26619,N_25855);
or UO_1956 (O_1956,N_25880,N_26652);
nand UO_1957 (O_1957,N_27291,N_25770);
xor UO_1958 (O_1958,N_27848,N_25893);
or UO_1959 (O_1959,N_29493,N_28944);
or UO_1960 (O_1960,N_27588,N_27459);
nor UO_1961 (O_1961,N_26334,N_26773);
nor UO_1962 (O_1962,N_27455,N_26134);
nand UO_1963 (O_1963,N_28559,N_26452);
and UO_1964 (O_1964,N_29652,N_27648);
nand UO_1965 (O_1965,N_29114,N_25081);
nor UO_1966 (O_1966,N_27523,N_29438);
or UO_1967 (O_1967,N_26951,N_27685);
nand UO_1968 (O_1968,N_26873,N_26803);
nor UO_1969 (O_1969,N_27465,N_25763);
or UO_1970 (O_1970,N_29836,N_28850);
xnor UO_1971 (O_1971,N_27937,N_26465);
nand UO_1972 (O_1972,N_26066,N_25137);
nor UO_1973 (O_1973,N_26079,N_26801);
and UO_1974 (O_1974,N_27094,N_26003);
and UO_1975 (O_1975,N_29738,N_28390);
and UO_1976 (O_1976,N_27167,N_26697);
nor UO_1977 (O_1977,N_25488,N_25783);
or UO_1978 (O_1978,N_25444,N_26667);
xnor UO_1979 (O_1979,N_28526,N_25006);
xor UO_1980 (O_1980,N_27553,N_26418);
or UO_1981 (O_1981,N_29974,N_29927);
and UO_1982 (O_1982,N_26133,N_25823);
and UO_1983 (O_1983,N_28343,N_25544);
xor UO_1984 (O_1984,N_25152,N_25476);
or UO_1985 (O_1985,N_28853,N_28738);
nand UO_1986 (O_1986,N_25759,N_28805);
xnor UO_1987 (O_1987,N_26214,N_27015);
nor UO_1988 (O_1988,N_26615,N_29094);
or UO_1989 (O_1989,N_29104,N_27736);
or UO_1990 (O_1990,N_26690,N_25503);
or UO_1991 (O_1991,N_25701,N_25529);
or UO_1992 (O_1992,N_26170,N_28940);
nor UO_1993 (O_1993,N_26706,N_27706);
nand UO_1994 (O_1994,N_28897,N_27529);
nor UO_1995 (O_1995,N_27389,N_28163);
and UO_1996 (O_1996,N_26461,N_28258);
and UO_1997 (O_1997,N_27997,N_27510);
nor UO_1998 (O_1998,N_26310,N_26899);
nor UO_1999 (O_1999,N_28594,N_26933);
and UO_2000 (O_2000,N_27372,N_25691);
xnor UO_2001 (O_2001,N_25480,N_29032);
or UO_2002 (O_2002,N_28190,N_27305);
nand UO_2003 (O_2003,N_26863,N_29357);
nor UO_2004 (O_2004,N_28257,N_28717);
and UO_2005 (O_2005,N_29067,N_25014);
or UO_2006 (O_2006,N_28372,N_29656);
xnor UO_2007 (O_2007,N_25633,N_26271);
or UO_2008 (O_2008,N_28304,N_27221);
or UO_2009 (O_2009,N_26604,N_28080);
xnor UO_2010 (O_2010,N_29694,N_26340);
or UO_2011 (O_2011,N_25109,N_29698);
and UO_2012 (O_2012,N_25359,N_26891);
nand UO_2013 (O_2013,N_29491,N_27130);
nor UO_2014 (O_2014,N_28223,N_26827);
or UO_2015 (O_2015,N_27881,N_26175);
and UO_2016 (O_2016,N_26456,N_25735);
and UO_2017 (O_2017,N_25761,N_26473);
or UO_2018 (O_2018,N_25186,N_26017);
and UO_2019 (O_2019,N_25087,N_28097);
and UO_2020 (O_2020,N_25939,N_27368);
and UO_2021 (O_2021,N_29296,N_29343);
and UO_2022 (O_2022,N_25226,N_25369);
xor UO_2023 (O_2023,N_29507,N_25862);
and UO_2024 (O_2024,N_27216,N_29962);
or UO_2025 (O_2025,N_25439,N_28415);
or UO_2026 (O_2026,N_28310,N_27026);
xnor UO_2027 (O_2027,N_28702,N_28198);
and UO_2028 (O_2028,N_28076,N_25453);
nor UO_2029 (O_2029,N_27377,N_26223);
nand UO_2030 (O_2030,N_28484,N_26736);
nor UO_2031 (O_2031,N_27966,N_27218);
or UO_2032 (O_2032,N_27456,N_29882);
and UO_2033 (O_2033,N_26626,N_25975);
xnor UO_2034 (O_2034,N_26752,N_29405);
nor UO_2035 (O_2035,N_29948,N_25377);
nor UO_2036 (O_2036,N_29418,N_28822);
nor UO_2037 (O_2037,N_25768,N_25231);
nand UO_2038 (O_2038,N_26299,N_27893);
and UO_2039 (O_2039,N_25634,N_26392);
or UO_2040 (O_2040,N_26868,N_28949);
or UO_2041 (O_2041,N_26925,N_28795);
xnor UO_2042 (O_2042,N_26485,N_28366);
and UO_2043 (O_2043,N_29019,N_27304);
xor UO_2044 (O_2044,N_25787,N_28900);
xor UO_2045 (O_2045,N_25920,N_27164);
or UO_2046 (O_2046,N_26397,N_26674);
xor UO_2047 (O_2047,N_27137,N_25097);
nor UO_2048 (O_2048,N_29886,N_25776);
nand UO_2049 (O_2049,N_27267,N_27847);
or UO_2050 (O_2050,N_26634,N_26538);
and UO_2051 (O_2051,N_25521,N_26215);
nand UO_2052 (O_2052,N_25182,N_28861);
nor UO_2053 (O_2053,N_28146,N_25110);
xor UO_2054 (O_2054,N_26356,N_27909);
xnor UO_2055 (O_2055,N_29874,N_29302);
and UO_2056 (O_2056,N_29270,N_27091);
nor UO_2057 (O_2057,N_26144,N_29518);
and UO_2058 (O_2058,N_26300,N_25856);
xnor UO_2059 (O_2059,N_29980,N_29740);
nand UO_2060 (O_2060,N_29217,N_25894);
nand UO_2061 (O_2061,N_25489,N_25514);
nand UO_2062 (O_2062,N_27009,N_26279);
and UO_2063 (O_2063,N_28074,N_29623);
and UO_2064 (O_2064,N_29778,N_25961);
nor UO_2065 (O_2065,N_27859,N_26877);
or UO_2066 (O_2066,N_29714,N_29309);
xnor UO_2067 (O_2067,N_28276,N_27418);
and UO_2068 (O_2068,N_26250,N_27433);
or UO_2069 (O_2069,N_25942,N_25178);
nand UO_2070 (O_2070,N_28779,N_28819);
nand UO_2071 (O_2071,N_25769,N_28842);
nand UO_2072 (O_2072,N_26942,N_26836);
or UO_2073 (O_2073,N_28599,N_25518);
and UO_2074 (O_2074,N_27353,N_28312);
and UO_2075 (O_2075,N_29913,N_25875);
nor UO_2076 (O_2076,N_26913,N_27999);
or UO_2077 (O_2077,N_29355,N_28349);
nand UO_2078 (O_2078,N_27791,N_25583);
xnor UO_2079 (O_2079,N_27956,N_28104);
or UO_2080 (O_2080,N_27690,N_26142);
or UO_2081 (O_2081,N_25921,N_29890);
nor UO_2082 (O_2082,N_26090,N_25419);
xnor UO_2083 (O_2083,N_28541,N_27684);
or UO_2084 (O_2084,N_29587,N_25304);
xnor UO_2085 (O_2085,N_27499,N_29910);
nand UO_2086 (O_2086,N_28860,N_25065);
nand UO_2087 (O_2087,N_25760,N_29940);
or UO_2088 (O_2088,N_29338,N_26165);
nand UO_2089 (O_2089,N_29366,N_26051);
nand UO_2090 (O_2090,N_25924,N_25997);
or UO_2091 (O_2091,N_28561,N_29639);
nor UO_2092 (O_2092,N_27975,N_29586);
or UO_2093 (O_2093,N_28562,N_26550);
or UO_2094 (O_2094,N_27405,N_26042);
nor UO_2095 (O_2095,N_28741,N_29973);
and UO_2096 (O_2096,N_27596,N_28981);
or UO_2097 (O_2097,N_26455,N_25765);
or UO_2098 (O_2098,N_27242,N_26018);
or UO_2099 (O_2099,N_25030,N_26341);
and UO_2100 (O_2100,N_26936,N_26010);
or UO_2101 (O_2101,N_29766,N_29861);
and UO_2102 (O_2102,N_27437,N_29054);
or UO_2103 (O_2103,N_29595,N_29677);
xor UO_2104 (O_2104,N_27073,N_29179);
nor UO_2105 (O_2105,N_27138,N_26948);
or UO_2106 (O_2106,N_28586,N_25410);
or UO_2107 (O_2107,N_25553,N_29141);
and UO_2108 (O_2108,N_25200,N_27644);
nor UO_2109 (O_2109,N_26592,N_29833);
or UO_2110 (O_2110,N_25991,N_28996);
nor UO_2111 (O_2111,N_28423,N_25802);
nand UO_2112 (O_2112,N_26315,N_27869);
nor UO_2113 (O_2113,N_26649,N_25850);
or UO_2114 (O_2114,N_29956,N_25026);
or UO_2115 (O_2115,N_26525,N_29348);
xnor UO_2116 (O_2116,N_25227,N_28287);
and UO_2117 (O_2117,N_29472,N_26112);
xnor UO_2118 (O_2118,N_27968,N_26664);
or UO_2119 (O_2119,N_26777,N_25120);
nor UO_2120 (O_2120,N_27744,N_29136);
or UO_2121 (O_2121,N_25848,N_29040);
and UO_2122 (O_2122,N_26753,N_28038);
and UO_2123 (O_2123,N_29828,N_28348);
and UO_2124 (O_2124,N_27209,N_25766);
and UO_2125 (O_2125,N_25833,N_28810);
nand UO_2126 (O_2126,N_25645,N_25556);
or UO_2127 (O_2127,N_29812,N_27603);
and UO_2128 (O_2128,N_29038,N_27889);
or UO_2129 (O_2129,N_28333,N_25901);
or UO_2130 (O_2130,N_25947,N_29354);
nor UO_2131 (O_2131,N_29496,N_26339);
nor UO_2132 (O_2132,N_25059,N_25844);
nor UO_2133 (O_2133,N_28679,N_28387);
nand UO_2134 (O_2134,N_25873,N_29791);
nand UO_2135 (O_2135,N_29207,N_28124);
xor UO_2136 (O_2136,N_29161,N_27606);
nor UO_2137 (O_2137,N_28604,N_26194);
or UO_2138 (O_2138,N_27549,N_29045);
nand UO_2139 (O_2139,N_26416,N_29706);
or UO_2140 (O_2140,N_26824,N_27074);
or UO_2141 (O_2141,N_26238,N_25132);
nand UO_2142 (O_2142,N_28152,N_28118);
nand UO_2143 (O_2143,N_28607,N_29628);
xnor UO_2144 (O_2144,N_29936,N_26982);
xnor UO_2145 (O_2145,N_25519,N_29222);
nand UO_2146 (O_2146,N_25557,N_28070);
xnor UO_2147 (O_2147,N_26805,N_28202);
and UO_2148 (O_2148,N_29308,N_27253);
or UO_2149 (O_2149,N_28045,N_28403);
or UO_2150 (O_2150,N_28029,N_29875);
and UO_2151 (O_2151,N_28666,N_29701);
nand UO_2152 (O_2152,N_25757,N_29276);
or UO_2153 (O_2153,N_27682,N_29210);
or UO_2154 (O_2154,N_28653,N_27140);
nand UO_2155 (O_2155,N_25362,N_26529);
xnor UO_2156 (O_2156,N_26940,N_28922);
nand UO_2157 (O_2157,N_29559,N_28745);
nand UO_2158 (O_2158,N_28720,N_25789);
or UO_2159 (O_2159,N_25143,N_27810);
nand UO_2160 (O_2160,N_26095,N_28200);
or UO_2161 (O_2161,N_29514,N_28250);
xnor UO_2162 (O_2162,N_25976,N_29021);
nand UO_2163 (O_2163,N_29626,N_29070);
and UO_2164 (O_2164,N_27720,N_27947);
nand UO_2165 (O_2165,N_29362,N_28577);
and UO_2166 (O_2166,N_28744,N_29313);
and UO_2167 (O_2167,N_29692,N_27233);
nand UO_2168 (O_2168,N_27100,N_29576);
nor UO_2169 (O_2169,N_27351,N_26008);
and UO_2170 (O_2170,N_25780,N_25223);
and UO_2171 (O_2171,N_25080,N_25849);
nand UO_2172 (O_2172,N_29416,N_28503);
and UO_2173 (O_2173,N_25800,N_25595);
nor UO_2174 (O_2174,N_25449,N_26387);
xor UO_2175 (O_2175,N_27114,N_29346);
or UO_2176 (O_2176,N_27914,N_28459);
nand UO_2177 (O_2177,N_26513,N_27772);
and UO_2178 (O_2178,N_28817,N_25221);
xor UO_2179 (O_2179,N_26289,N_26371);
nand UO_2180 (O_2180,N_28316,N_29508);
xor UO_2181 (O_2181,N_26186,N_25971);
or UO_2182 (O_2182,N_27067,N_27366);
nand UO_2183 (O_2183,N_29162,N_28487);
nor UO_2184 (O_2184,N_25589,N_25561);
nor UO_2185 (O_2185,N_28907,N_25970);
nand UO_2186 (O_2186,N_25646,N_27001);
nand UO_2187 (O_2187,N_28547,N_25995);
and UO_2188 (O_2188,N_28748,N_26854);
and UO_2189 (O_2189,N_28774,N_28094);
or UO_2190 (O_2190,N_27952,N_25878);
or UO_2191 (O_2191,N_28660,N_28353);
nand UO_2192 (O_2192,N_26630,N_25967);
or UO_2193 (O_2193,N_27617,N_25005);
xnor UO_2194 (O_2194,N_25533,N_26526);
nand UO_2195 (O_2195,N_26996,N_25219);
or UO_2196 (O_2196,N_28442,N_26580);
nand UO_2197 (O_2197,N_28239,N_26365);
and UO_2198 (O_2198,N_26421,N_27444);
nor UO_2199 (O_2199,N_25312,N_25208);
or UO_2200 (O_2200,N_26174,N_29028);
and UO_2201 (O_2201,N_27332,N_26917);
nor UO_2202 (O_2202,N_29845,N_29763);
nor UO_2203 (O_2203,N_26627,N_28464);
or UO_2204 (O_2204,N_25741,N_26610);
and UO_2205 (O_2205,N_29822,N_28266);
nor UO_2206 (O_2206,N_26184,N_27431);
nand UO_2207 (O_2207,N_25413,N_27925);
nand UO_2208 (O_2208,N_25588,N_28294);
nor UO_2209 (O_2209,N_27261,N_25295);
nor UO_2210 (O_2210,N_26069,N_27084);
xnor UO_2211 (O_2211,N_29953,N_26789);
and UO_2212 (O_2212,N_29684,N_29930);
and UO_2213 (O_2213,N_27971,N_26442);
nand UO_2214 (O_2214,N_25228,N_25729);
nor UO_2215 (O_2215,N_26135,N_28219);
or UO_2216 (O_2216,N_26389,N_26332);
nand UO_2217 (O_2217,N_26091,N_29476);
xnor UO_2218 (O_2218,N_27857,N_28295);
nor UO_2219 (O_2219,N_26360,N_27571);
nor UO_2220 (O_2220,N_29332,N_26781);
or UO_2221 (O_2221,N_27398,N_29735);
and UO_2222 (O_2222,N_28941,N_26067);
nand UO_2223 (O_2223,N_28769,N_27240);
nor UO_2224 (O_2224,N_25408,N_27702);
or UO_2225 (O_2225,N_28418,N_29026);
or UO_2226 (O_2226,N_28573,N_26046);
nor UO_2227 (O_2227,N_25972,N_26701);
nor UO_2228 (O_2228,N_28546,N_27568);
or UO_2229 (O_2229,N_29260,N_29624);
and UO_2230 (O_2230,N_27295,N_27493);
xor UO_2231 (O_2231,N_28326,N_26591);
nor UO_2232 (O_2232,N_25957,N_26273);
nand UO_2233 (O_2233,N_29629,N_26119);
or UO_2234 (O_2234,N_25095,N_25196);
nand UO_2235 (O_2235,N_27171,N_26799);
nor UO_2236 (O_2236,N_26395,N_25913);
nor UO_2237 (O_2237,N_28532,N_28249);
nor UO_2238 (O_2238,N_29750,N_29414);
nand UO_2239 (O_2239,N_28064,N_26959);
nor UO_2240 (O_2240,N_29896,N_29721);
or UO_2241 (O_2241,N_27749,N_27796);
and UO_2242 (O_2242,N_28350,N_26363);
or UO_2243 (O_2243,N_29214,N_26722);
xnor UO_2244 (O_2244,N_27487,N_25980);
and UO_2245 (O_2245,N_29789,N_27347);
nor UO_2246 (O_2246,N_27120,N_28714);
or UO_2247 (O_2247,N_25599,N_28116);
and UO_2248 (O_2248,N_29097,N_27667);
nor UO_2249 (O_2249,N_25945,N_28099);
or UO_2250 (O_2250,N_26957,N_25676);
or UO_2251 (O_2251,N_27417,N_26378);
xnor UO_2252 (O_2252,N_29340,N_28396);
or UO_2253 (O_2253,N_29084,N_29024);
nand UO_2254 (O_2254,N_25401,N_25470);
nor UO_2255 (O_2255,N_29985,N_27395);
and UO_2256 (O_2256,N_25864,N_29900);
nor UO_2257 (O_2257,N_29718,N_25015);
and UO_2258 (O_2258,N_26739,N_26501);
or UO_2259 (O_2259,N_28910,N_27313);
and UO_2260 (O_2260,N_26036,N_25048);
or UO_2261 (O_2261,N_27391,N_26831);
or UO_2262 (O_2262,N_28386,N_26349);
or UO_2263 (O_2263,N_27544,N_25184);
xor UO_2264 (O_2264,N_29952,N_26968);
or UO_2265 (O_2265,N_25616,N_26800);
and UO_2266 (O_2266,N_28549,N_27663);
nand UO_2267 (O_2267,N_28707,N_25268);
nand UO_2268 (O_2268,N_27188,N_29076);
or UO_2269 (O_2269,N_29751,N_25686);
nor UO_2270 (O_2270,N_25385,N_28807);
nand UO_2271 (O_2271,N_27024,N_25689);
or UO_2272 (O_2272,N_28218,N_29005);
nand UO_2273 (O_2273,N_26710,N_29557);
xor UO_2274 (O_2274,N_27264,N_25154);
or UO_2275 (O_2275,N_26322,N_26603);
or UO_2276 (O_2276,N_28301,N_25882);
xnor UO_2277 (O_2277,N_27727,N_26974);
and UO_2278 (O_2278,N_29387,N_29150);
and UO_2279 (O_2279,N_27408,N_27119);
nand UO_2280 (O_2280,N_26594,N_25432);
nand UO_2281 (O_2281,N_29143,N_25174);
nand UO_2282 (O_2282,N_27983,N_25092);
xor UO_2283 (O_2283,N_28049,N_28794);
nor UO_2284 (O_2284,N_28083,N_29790);
or UO_2285 (O_2285,N_27349,N_29103);
nor UO_2286 (O_2286,N_25914,N_27457);
and UO_2287 (O_2287,N_26282,N_28631);
or UO_2288 (O_2288,N_28960,N_26648);
and UO_2289 (O_2289,N_29892,N_26712);
nor UO_2290 (O_2290,N_28694,N_25098);
and UO_2291 (O_2291,N_27131,N_28357);
xor UO_2292 (O_2292,N_29154,N_25106);
xnor UO_2293 (O_2293,N_25937,N_28174);
xnor UO_2294 (O_2294,N_28138,N_25160);
and UO_2295 (O_2295,N_25717,N_25949);
nor UO_2296 (O_2296,N_26252,N_25049);
or UO_2297 (O_2297,N_29102,N_27439);
and UO_2298 (O_2298,N_29577,N_28869);
nand UO_2299 (O_2299,N_25334,N_28786);
nor UO_2300 (O_2300,N_26048,N_25180);
and UO_2301 (O_2301,N_27178,N_28522);
or UO_2302 (O_2302,N_28918,N_29080);
nor UO_2303 (O_2303,N_27219,N_28673);
nor UO_2304 (O_2304,N_26375,N_28690);
or UO_2305 (O_2305,N_26155,N_28237);
and UO_2306 (O_2306,N_28212,N_27127);
nor UO_2307 (O_2307,N_26661,N_25234);
nor UO_2308 (O_2308,N_28685,N_29247);
nor UO_2309 (O_2309,N_29117,N_27378);
and UO_2310 (O_2310,N_25934,N_29252);
and UO_2311 (O_2311,N_27669,N_28692);
nor UO_2312 (O_2312,N_27019,N_26255);
nand UO_2313 (O_2313,N_28095,N_27163);
xnor UO_2314 (O_2314,N_25113,N_26025);
xnor UO_2315 (O_2315,N_28355,N_28798);
nand UO_2316 (O_2316,N_27142,N_26986);
nor UO_2317 (O_2317,N_29968,N_27268);
nand UO_2318 (O_2318,N_28009,N_28067);
or UO_2319 (O_2319,N_25775,N_27500);
and UO_2320 (O_2320,N_28934,N_26480);
nor UO_2321 (O_2321,N_26890,N_26930);
and UO_2322 (O_2322,N_27192,N_26835);
and UO_2323 (O_2323,N_26573,N_27275);
and UO_2324 (O_2324,N_27895,N_27420);
or UO_2325 (O_2325,N_25364,N_27827);
or UO_2326 (O_2326,N_28605,N_28283);
nor UO_2327 (O_2327,N_26080,N_28670);
nand UO_2328 (O_2328,N_27576,N_26886);
nor UO_2329 (O_2329,N_25696,N_29153);
and UO_2330 (O_2330,N_25402,N_29571);
nor UO_2331 (O_2331,N_27246,N_26792);
nor UO_2332 (O_2332,N_28046,N_29183);
or UO_2333 (O_2333,N_28534,N_28098);
nor UO_2334 (O_2334,N_25069,N_28229);
and UO_2335 (O_2335,N_26012,N_27328);
and UO_2336 (O_2336,N_28439,N_29583);
nand UO_2337 (O_2337,N_27039,N_26113);
and UO_2338 (O_2338,N_26548,N_26230);
xnor UO_2339 (O_2339,N_28570,N_25874);
nor UO_2340 (O_2340,N_27543,N_27197);
nand UO_2341 (O_2341,N_25045,N_29337);
nor UO_2342 (O_2342,N_27234,N_28925);
or UO_2343 (O_2343,N_25263,N_28890);
and UO_2344 (O_2344,N_27709,N_26500);
or UO_2345 (O_2345,N_28209,N_25643);
nor UO_2346 (O_2346,N_27301,N_27148);
nor UO_2347 (O_2347,N_27482,N_29221);
and UO_2348 (O_2348,N_27338,N_27527);
nor UO_2349 (O_2349,N_29007,N_28430);
nor UO_2350 (O_2350,N_25085,N_25877);
nor UO_2351 (O_2351,N_28711,N_27683);
and UO_2352 (O_2352,N_27077,N_29167);
xnor UO_2353 (O_2353,N_26052,N_26983);
or UO_2354 (O_2354,N_28990,N_28669);
nand UO_2355 (O_2355,N_25292,N_28132);
xnor UO_2356 (O_2356,N_26964,N_28175);
or UO_2357 (O_2357,N_27610,N_29318);
and UO_2358 (O_2358,N_25370,N_28936);
xnor UO_2359 (O_2359,N_27367,N_26961);
and UO_2360 (O_2360,N_28422,N_28567);
or UO_2361 (O_2361,N_28154,N_27079);
nand UO_2362 (O_2362,N_29327,N_29165);
nor UO_2363 (O_2363,N_25960,N_28756);
and UO_2364 (O_2364,N_29895,N_26030);
or UO_2365 (O_2365,N_27027,N_29521);
nor UO_2366 (O_2366,N_27104,N_28280);
or UO_2367 (O_2367,N_26871,N_27867);
nor UO_2368 (O_2368,N_27877,N_29675);
and UO_2369 (O_2369,N_26478,N_28905);
or UO_2370 (O_2370,N_26507,N_28248);
nor UO_2371 (O_2371,N_29771,N_25036);
or UO_2372 (O_2372,N_26024,N_29397);
and UO_2373 (O_2373,N_27748,N_25300);
nand UO_2374 (O_2374,N_26240,N_28432);
or UO_2375 (O_2375,N_28880,N_26345);
nand UO_2376 (O_2376,N_27519,N_27927);
and UO_2377 (O_2377,N_27556,N_26874);
nand UO_2378 (O_2378,N_25922,N_25572);
nor UO_2379 (O_2379,N_28582,N_29014);
nand UO_2380 (O_2380,N_27050,N_26049);
xor UO_2381 (O_2381,N_29645,N_29803);
nor UO_2382 (O_2382,N_25737,N_26470);
xor UO_2383 (O_2383,N_29052,N_25990);
xnor UO_2384 (O_2384,N_27652,N_29942);
nor UO_2385 (O_2385,N_28972,N_28597);
and UO_2386 (O_2386,N_27115,N_27689);
nor UO_2387 (O_2387,N_25241,N_28377);
or UO_2388 (O_2388,N_29596,N_29049);
or UO_2389 (O_2389,N_26274,N_27716);
and UO_2390 (O_2390,N_29312,N_28876);
nor UO_2391 (O_2391,N_28952,N_29219);
nand UO_2392 (O_2392,N_29538,N_29450);
xnor UO_2393 (O_2393,N_29212,N_26399);
nand UO_2394 (O_2394,N_29743,N_29160);
nand UO_2395 (O_2395,N_29211,N_26883);
or UO_2396 (O_2396,N_25613,N_25825);
and UO_2397 (O_2397,N_26694,N_28651);
nand UO_2398 (O_2398,N_27601,N_26482);
nor UO_2399 (O_2399,N_27257,N_25927);
nor UO_2400 (O_2400,N_27821,N_29317);
and UO_2401 (O_2401,N_28622,N_25002);
or UO_2402 (O_2402,N_26406,N_26905);
nand UO_2403 (O_2403,N_25291,N_26426);
nand UO_2404 (O_2404,N_25344,N_25898);
and UO_2405 (O_2405,N_27203,N_25500);
xnor UO_2406 (O_2406,N_25865,N_29897);
or UO_2407 (O_2407,N_26814,N_25754);
or UO_2408 (O_2408,N_27099,N_29256);
or UO_2409 (O_2409,N_28449,N_26037);
nor UO_2410 (O_2410,N_29865,N_26347);
nor UO_2411 (O_2411,N_28883,N_25140);
nand UO_2412 (O_2412,N_28579,N_27160);
nor UO_2413 (O_2413,N_25615,N_27740);
or UO_2414 (O_2414,N_28321,N_29742);
and UO_2415 (O_2415,N_28652,N_26047);
and UO_2416 (O_2416,N_26311,N_27982);
and UO_2417 (O_2417,N_29202,N_28820);
and UO_2418 (O_2418,N_29470,N_29090);
nor UO_2419 (O_2419,N_28667,N_25105);
nand UO_2420 (O_2420,N_27365,N_29689);
or UO_2421 (O_2421,N_29147,N_29421);
or UO_2422 (O_2422,N_25509,N_27884);
and UO_2423 (O_2423,N_25499,N_27206);
nand UO_2424 (O_2424,N_26555,N_29819);
and UO_2425 (O_2425,N_25528,N_28832);
nor UO_2426 (O_2426,N_26458,N_28743);
and UO_2427 (O_2427,N_29351,N_29451);
or UO_2428 (O_2428,N_26285,N_29106);
and UO_2429 (O_2429,N_27928,N_27410);
nand UO_2430 (O_2430,N_26565,N_26915);
nor UO_2431 (O_2431,N_26379,N_28615);
or UO_2432 (O_2432,N_28628,N_29862);
nor UO_2433 (O_2433,N_27277,N_27070);
or UO_2434 (O_2434,N_27619,N_26206);
nand UO_2435 (O_2435,N_29505,N_28975);
or UO_2436 (O_2436,N_27283,N_29376);
xor UO_2437 (O_2437,N_25568,N_25078);
and UO_2438 (O_2438,N_25593,N_26469);
and UO_2439 (O_2439,N_29637,N_26747);
or UO_2440 (O_2440,N_29826,N_26141);
or UO_2441 (O_2441,N_26806,N_27955);
and UO_2442 (O_2442,N_26776,N_28514);
and UO_2443 (O_2443,N_27425,N_27229);
and UO_2444 (O_2444,N_26129,N_27521);
nand UO_2445 (O_2445,N_27637,N_26132);
nand UO_2446 (O_2446,N_27868,N_27011);
and UO_2447 (O_2447,N_28525,N_28991);
and UO_2448 (O_2448,N_27917,N_28445);
and UO_2449 (O_2449,N_27147,N_27089);
xnor UO_2450 (O_2450,N_26331,N_27451);
or UO_2451 (O_2451,N_25089,N_28513);
or UO_2452 (O_2452,N_25442,N_28829);
and UO_2453 (O_2453,N_27158,N_29921);
nor UO_2454 (O_2454,N_26740,N_27575);
xor UO_2455 (O_2455,N_28870,N_29350);
and UO_2456 (O_2456,N_26734,N_29792);
or UO_2457 (O_2457,N_26286,N_28725);
nor UO_2458 (O_2458,N_27359,N_27103);
or UO_2459 (O_2459,N_29998,N_27362);
nor UO_2460 (O_2460,N_28722,N_25122);
nor UO_2461 (O_2461,N_26148,N_28305);
and UO_2462 (O_2462,N_26849,N_28580);
nand UO_2463 (O_2463,N_29025,N_29171);
and UO_2464 (O_2464,N_25665,N_29887);
nor UO_2465 (O_2465,N_28908,N_28369);
xnor UO_2466 (O_2466,N_25146,N_27672);
and UO_2467 (O_2467,N_25654,N_27022);
and UO_2468 (O_2468,N_28214,N_25472);
xor UO_2469 (O_2469,N_27236,N_27028);
xnor UO_2470 (O_2470,N_29582,N_27655);
and UO_2471 (O_2471,N_29667,N_25409);
or UO_2472 (O_2472,N_27687,N_26970);
nor UO_2473 (O_2473,N_28623,N_26737);
nand UO_2474 (O_2474,N_26869,N_25354);
and UO_2475 (O_2475,N_26602,N_26845);
or UO_2476 (O_2476,N_25050,N_29502);
or UO_2477 (O_2477,N_27035,N_25194);
or UO_2478 (O_2478,N_26401,N_28988);
xor UO_2479 (O_2479,N_25720,N_26029);
and UO_2480 (O_2480,N_28844,N_28520);
and UO_2481 (O_2481,N_28402,N_29258);
xor UO_2482 (O_2482,N_25044,N_27662);
nand UO_2483 (O_2483,N_28081,N_29560);
nand UO_2484 (O_2484,N_26586,N_26280);
xor UO_2485 (O_2485,N_28340,N_26988);
and UO_2486 (O_2486,N_29098,N_28093);
nor UO_2487 (O_2487,N_26212,N_25493);
nor UO_2488 (O_2488,N_27143,N_29769);
nor UO_2489 (O_2489,N_26390,N_25283);
or UO_2490 (O_2490,N_29048,N_26075);
or UO_2491 (O_2491,N_28771,N_26269);
and UO_2492 (O_2492,N_26237,N_29977);
or UO_2493 (O_2493,N_25507,N_27503);
nand UO_2494 (O_2494,N_28410,N_26076);
or UO_2495 (O_2495,N_26073,N_27266);
nor UO_2496 (O_2496,N_28509,N_26168);
or UO_2497 (O_2497,N_25630,N_27852);
and UO_2498 (O_2498,N_25793,N_26366);
and UO_2499 (O_2499,N_25115,N_26180);
nand UO_2500 (O_2500,N_26088,N_29953);
or UO_2501 (O_2501,N_29004,N_26502);
or UO_2502 (O_2502,N_26870,N_29649);
nor UO_2503 (O_2503,N_26172,N_25185);
nand UO_2504 (O_2504,N_27386,N_28700);
nor UO_2505 (O_2505,N_25581,N_26069);
nor UO_2506 (O_2506,N_29194,N_27473);
nand UO_2507 (O_2507,N_25245,N_26427);
nand UO_2508 (O_2508,N_28023,N_25186);
nand UO_2509 (O_2509,N_26285,N_28026);
nor UO_2510 (O_2510,N_26264,N_26416);
nor UO_2511 (O_2511,N_28842,N_27784);
or UO_2512 (O_2512,N_26148,N_27093);
and UO_2513 (O_2513,N_29820,N_27225);
nand UO_2514 (O_2514,N_25716,N_29893);
nor UO_2515 (O_2515,N_25832,N_25957);
and UO_2516 (O_2516,N_28799,N_26411);
and UO_2517 (O_2517,N_29659,N_28203);
or UO_2518 (O_2518,N_29856,N_26417);
and UO_2519 (O_2519,N_28203,N_25286);
and UO_2520 (O_2520,N_25354,N_25981);
and UO_2521 (O_2521,N_25829,N_25264);
nor UO_2522 (O_2522,N_25510,N_28367);
and UO_2523 (O_2523,N_26719,N_28574);
nand UO_2524 (O_2524,N_26094,N_28660);
nand UO_2525 (O_2525,N_27217,N_29045);
or UO_2526 (O_2526,N_28204,N_25309);
nor UO_2527 (O_2527,N_25855,N_29109);
nor UO_2528 (O_2528,N_25923,N_28853);
nand UO_2529 (O_2529,N_29591,N_28616);
xnor UO_2530 (O_2530,N_29181,N_25607);
or UO_2531 (O_2531,N_25833,N_27736);
nand UO_2532 (O_2532,N_25073,N_27019);
xor UO_2533 (O_2533,N_28508,N_26855);
and UO_2534 (O_2534,N_29625,N_26123);
nand UO_2535 (O_2535,N_27531,N_28348);
or UO_2536 (O_2536,N_25975,N_29211);
nand UO_2537 (O_2537,N_29170,N_25626);
and UO_2538 (O_2538,N_27668,N_26804);
and UO_2539 (O_2539,N_26533,N_28814);
nand UO_2540 (O_2540,N_26654,N_28284);
xor UO_2541 (O_2541,N_29249,N_28513);
nor UO_2542 (O_2542,N_27295,N_28820);
nand UO_2543 (O_2543,N_25562,N_27806);
or UO_2544 (O_2544,N_28122,N_28086);
or UO_2545 (O_2545,N_28313,N_26170);
xor UO_2546 (O_2546,N_26534,N_29294);
nand UO_2547 (O_2547,N_27139,N_26631);
and UO_2548 (O_2548,N_25442,N_26967);
nor UO_2549 (O_2549,N_29406,N_25492);
xor UO_2550 (O_2550,N_25485,N_25471);
nand UO_2551 (O_2551,N_29309,N_28618);
and UO_2552 (O_2552,N_25919,N_28619);
and UO_2553 (O_2553,N_29306,N_26982);
xor UO_2554 (O_2554,N_29586,N_28986);
or UO_2555 (O_2555,N_29532,N_27398);
xor UO_2556 (O_2556,N_27629,N_27694);
or UO_2557 (O_2557,N_27521,N_29880);
nor UO_2558 (O_2558,N_29641,N_26854);
nand UO_2559 (O_2559,N_28441,N_25610);
or UO_2560 (O_2560,N_25997,N_26796);
xnor UO_2561 (O_2561,N_29320,N_26307);
and UO_2562 (O_2562,N_26897,N_27296);
xor UO_2563 (O_2563,N_29575,N_25753);
nand UO_2564 (O_2564,N_26764,N_26015);
xnor UO_2565 (O_2565,N_26567,N_26774);
or UO_2566 (O_2566,N_28252,N_27940);
nand UO_2567 (O_2567,N_29100,N_29304);
nor UO_2568 (O_2568,N_26939,N_26936);
nor UO_2569 (O_2569,N_26394,N_25330);
nor UO_2570 (O_2570,N_29887,N_27827);
nor UO_2571 (O_2571,N_28688,N_29918);
or UO_2572 (O_2572,N_25600,N_26391);
nand UO_2573 (O_2573,N_28601,N_26193);
nand UO_2574 (O_2574,N_27286,N_28451);
and UO_2575 (O_2575,N_27357,N_29403);
nor UO_2576 (O_2576,N_27632,N_27145);
nor UO_2577 (O_2577,N_25564,N_28161);
and UO_2578 (O_2578,N_26865,N_25487);
xor UO_2579 (O_2579,N_25400,N_29075);
nor UO_2580 (O_2580,N_25064,N_26325);
or UO_2581 (O_2581,N_27779,N_28703);
xor UO_2582 (O_2582,N_25732,N_29105);
or UO_2583 (O_2583,N_28168,N_28441);
nand UO_2584 (O_2584,N_25046,N_29406);
nand UO_2585 (O_2585,N_26912,N_29174);
nand UO_2586 (O_2586,N_26935,N_27316);
and UO_2587 (O_2587,N_28792,N_26822);
or UO_2588 (O_2588,N_26247,N_27957);
or UO_2589 (O_2589,N_25948,N_26720);
nor UO_2590 (O_2590,N_26059,N_27050);
and UO_2591 (O_2591,N_26264,N_29251);
and UO_2592 (O_2592,N_25008,N_29591);
xnor UO_2593 (O_2593,N_25443,N_29206);
and UO_2594 (O_2594,N_27374,N_29248);
xnor UO_2595 (O_2595,N_26073,N_28435);
nor UO_2596 (O_2596,N_28938,N_25576);
xor UO_2597 (O_2597,N_28495,N_27645);
or UO_2598 (O_2598,N_28816,N_27666);
and UO_2599 (O_2599,N_28544,N_26583);
nor UO_2600 (O_2600,N_29914,N_28895);
and UO_2601 (O_2601,N_27732,N_28245);
nand UO_2602 (O_2602,N_25984,N_27864);
nor UO_2603 (O_2603,N_26309,N_25260);
xnor UO_2604 (O_2604,N_25497,N_29509);
nor UO_2605 (O_2605,N_27904,N_28950);
nor UO_2606 (O_2606,N_27240,N_27096);
xnor UO_2607 (O_2607,N_26923,N_26887);
or UO_2608 (O_2608,N_25505,N_27763);
or UO_2609 (O_2609,N_27725,N_29649);
nand UO_2610 (O_2610,N_25469,N_25782);
xor UO_2611 (O_2611,N_27922,N_29602);
xnor UO_2612 (O_2612,N_26253,N_25866);
or UO_2613 (O_2613,N_29245,N_29333);
and UO_2614 (O_2614,N_28167,N_26257);
and UO_2615 (O_2615,N_26849,N_27989);
and UO_2616 (O_2616,N_29580,N_26063);
nor UO_2617 (O_2617,N_27216,N_29276);
nand UO_2618 (O_2618,N_28174,N_26253);
nor UO_2619 (O_2619,N_27857,N_28302);
or UO_2620 (O_2620,N_27835,N_27941);
nor UO_2621 (O_2621,N_26833,N_28998);
nor UO_2622 (O_2622,N_29340,N_25550);
and UO_2623 (O_2623,N_28034,N_27045);
and UO_2624 (O_2624,N_29566,N_27385);
or UO_2625 (O_2625,N_26998,N_27374);
nor UO_2626 (O_2626,N_26107,N_29780);
nor UO_2627 (O_2627,N_27137,N_27503);
or UO_2628 (O_2628,N_26591,N_26232);
nor UO_2629 (O_2629,N_29434,N_25616);
or UO_2630 (O_2630,N_27060,N_27237);
nor UO_2631 (O_2631,N_28047,N_27871);
nand UO_2632 (O_2632,N_28689,N_25346);
nor UO_2633 (O_2633,N_27083,N_27767);
nor UO_2634 (O_2634,N_27435,N_27535);
nor UO_2635 (O_2635,N_25905,N_27292);
nand UO_2636 (O_2636,N_25799,N_28555);
nor UO_2637 (O_2637,N_28836,N_28079);
and UO_2638 (O_2638,N_29262,N_25372);
nor UO_2639 (O_2639,N_29249,N_25736);
nand UO_2640 (O_2640,N_28274,N_28846);
and UO_2641 (O_2641,N_26849,N_25053);
nand UO_2642 (O_2642,N_27085,N_28050);
nor UO_2643 (O_2643,N_25226,N_28440);
nand UO_2644 (O_2644,N_25190,N_25536);
nor UO_2645 (O_2645,N_26786,N_26422);
xor UO_2646 (O_2646,N_26158,N_26365);
nor UO_2647 (O_2647,N_27459,N_25517);
nand UO_2648 (O_2648,N_29398,N_29665);
or UO_2649 (O_2649,N_25277,N_28452);
and UO_2650 (O_2650,N_28415,N_29082);
nand UO_2651 (O_2651,N_25091,N_27667);
xnor UO_2652 (O_2652,N_26916,N_27491);
nand UO_2653 (O_2653,N_25857,N_28794);
xnor UO_2654 (O_2654,N_25375,N_27448);
or UO_2655 (O_2655,N_26609,N_26135);
nor UO_2656 (O_2656,N_27016,N_28948);
nor UO_2657 (O_2657,N_28510,N_25512);
and UO_2658 (O_2658,N_26593,N_25053);
nand UO_2659 (O_2659,N_28603,N_25125);
xnor UO_2660 (O_2660,N_25450,N_26048);
nor UO_2661 (O_2661,N_28890,N_28444);
nor UO_2662 (O_2662,N_25970,N_28464);
and UO_2663 (O_2663,N_28590,N_27859);
nand UO_2664 (O_2664,N_25425,N_25598);
or UO_2665 (O_2665,N_26371,N_27029);
nand UO_2666 (O_2666,N_28702,N_26086);
and UO_2667 (O_2667,N_26172,N_25739);
nand UO_2668 (O_2668,N_26853,N_26960);
and UO_2669 (O_2669,N_25858,N_29805);
or UO_2670 (O_2670,N_29048,N_25947);
and UO_2671 (O_2671,N_26706,N_28424);
or UO_2672 (O_2672,N_28609,N_27981);
nor UO_2673 (O_2673,N_25752,N_29740);
xor UO_2674 (O_2674,N_26580,N_27321);
and UO_2675 (O_2675,N_26648,N_28697);
and UO_2676 (O_2676,N_26591,N_28371);
and UO_2677 (O_2677,N_28308,N_26010);
xnor UO_2678 (O_2678,N_25576,N_29118);
or UO_2679 (O_2679,N_27432,N_28894);
or UO_2680 (O_2680,N_29996,N_25165);
and UO_2681 (O_2681,N_25128,N_27760);
or UO_2682 (O_2682,N_25613,N_28824);
or UO_2683 (O_2683,N_26514,N_28431);
or UO_2684 (O_2684,N_27595,N_25417);
or UO_2685 (O_2685,N_29074,N_27836);
and UO_2686 (O_2686,N_27731,N_27931);
nor UO_2687 (O_2687,N_29599,N_29608);
and UO_2688 (O_2688,N_26276,N_25554);
nor UO_2689 (O_2689,N_27092,N_27972);
xor UO_2690 (O_2690,N_26813,N_25851);
nor UO_2691 (O_2691,N_29707,N_28775);
and UO_2692 (O_2692,N_26223,N_28372);
or UO_2693 (O_2693,N_25212,N_28220);
nand UO_2694 (O_2694,N_26486,N_25766);
nor UO_2695 (O_2695,N_29303,N_27056);
xor UO_2696 (O_2696,N_25119,N_26961);
nor UO_2697 (O_2697,N_27320,N_25215);
or UO_2698 (O_2698,N_29390,N_29918);
and UO_2699 (O_2699,N_27374,N_28590);
or UO_2700 (O_2700,N_28685,N_27909);
nand UO_2701 (O_2701,N_26984,N_27316);
nand UO_2702 (O_2702,N_26580,N_27678);
xor UO_2703 (O_2703,N_27700,N_29504);
and UO_2704 (O_2704,N_26130,N_25456);
or UO_2705 (O_2705,N_29516,N_26025);
or UO_2706 (O_2706,N_25778,N_26961);
nand UO_2707 (O_2707,N_28760,N_25654);
and UO_2708 (O_2708,N_26640,N_29719);
xor UO_2709 (O_2709,N_26732,N_28925);
or UO_2710 (O_2710,N_25158,N_28426);
or UO_2711 (O_2711,N_27770,N_29480);
nand UO_2712 (O_2712,N_26940,N_25048);
nand UO_2713 (O_2713,N_28463,N_25746);
xor UO_2714 (O_2714,N_28652,N_28618);
and UO_2715 (O_2715,N_25134,N_27954);
nor UO_2716 (O_2716,N_25950,N_28721);
or UO_2717 (O_2717,N_25471,N_26015);
nand UO_2718 (O_2718,N_27464,N_27521);
nand UO_2719 (O_2719,N_26155,N_28592);
or UO_2720 (O_2720,N_26918,N_29606);
nand UO_2721 (O_2721,N_29196,N_29304);
xnor UO_2722 (O_2722,N_27260,N_27208);
nor UO_2723 (O_2723,N_26028,N_29006);
xnor UO_2724 (O_2724,N_25568,N_27111);
nor UO_2725 (O_2725,N_27494,N_27654);
and UO_2726 (O_2726,N_28719,N_25583);
nand UO_2727 (O_2727,N_29808,N_28380);
or UO_2728 (O_2728,N_25464,N_28348);
and UO_2729 (O_2729,N_27468,N_25957);
and UO_2730 (O_2730,N_28230,N_26001);
and UO_2731 (O_2731,N_27740,N_29909);
or UO_2732 (O_2732,N_25131,N_25030);
or UO_2733 (O_2733,N_25595,N_26884);
and UO_2734 (O_2734,N_26480,N_26066);
nand UO_2735 (O_2735,N_25617,N_25932);
nand UO_2736 (O_2736,N_25630,N_29053);
and UO_2737 (O_2737,N_28931,N_25092);
or UO_2738 (O_2738,N_27241,N_27715);
or UO_2739 (O_2739,N_26018,N_29995);
and UO_2740 (O_2740,N_29103,N_29181);
nand UO_2741 (O_2741,N_26181,N_27366);
nand UO_2742 (O_2742,N_29946,N_25093);
and UO_2743 (O_2743,N_25465,N_28469);
nor UO_2744 (O_2744,N_25343,N_27344);
nand UO_2745 (O_2745,N_25119,N_28311);
and UO_2746 (O_2746,N_28690,N_29850);
nand UO_2747 (O_2747,N_28441,N_25430);
nor UO_2748 (O_2748,N_26577,N_26334);
and UO_2749 (O_2749,N_25478,N_27815);
nand UO_2750 (O_2750,N_29548,N_29861);
nand UO_2751 (O_2751,N_27122,N_25082);
and UO_2752 (O_2752,N_28515,N_28739);
and UO_2753 (O_2753,N_29546,N_27311);
nand UO_2754 (O_2754,N_26139,N_29683);
or UO_2755 (O_2755,N_26438,N_28449);
nor UO_2756 (O_2756,N_25100,N_28693);
nand UO_2757 (O_2757,N_29909,N_29590);
and UO_2758 (O_2758,N_29071,N_29415);
nor UO_2759 (O_2759,N_28740,N_28753);
nor UO_2760 (O_2760,N_26561,N_25657);
nand UO_2761 (O_2761,N_25558,N_28565);
and UO_2762 (O_2762,N_29556,N_25807);
nor UO_2763 (O_2763,N_27986,N_29118);
nand UO_2764 (O_2764,N_26643,N_28100);
nor UO_2765 (O_2765,N_26600,N_27553);
nor UO_2766 (O_2766,N_27473,N_27055);
and UO_2767 (O_2767,N_26781,N_26214);
xnor UO_2768 (O_2768,N_28314,N_27388);
and UO_2769 (O_2769,N_28355,N_27537);
and UO_2770 (O_2770,N_28709,N_28576);
xnor UO_2771 (O_2771,N_28425,N_25102);
and UO_2772 (O_2772,N_27482,N_27949);
xor UO_2773 (O_2773,N_25501,N_28295);
and UO_2774 (O_2774,N_29775,N_27177);
nand UO_2775 (O_2775,N_25144,N_27207);
or UO_2776 (O_2776,N_26311,N_25521);
and UO_2777 (O_2777,N_27690,N_25004);
nor UO_2778 (O_2778,N_29505,N_27161);
and UO_2779 (O_2779,N_25678,N_29367);
and UO_2780 (O_2780,N_28122,N_27522);
or UO_2781 (O_2781,N_26279,N_26271);
or UO_2782 (O_2782,N_25317,N_28118);
xnor UO_2783 (O_2783,N_26432,N_26434);
or UO_2784 (O_2784,N_27233,N_26888);
and UO_2785 (O_2785,N_25374,N_26869);
and UO_2786 (O_2786,N_27570,N_28153);
xor UO_2787 (O_2787,N_27339,N_28514);
xor UO_2788 (O_2788,N_25175,N_29826);
nor UO_2789 (O_2789,N_27548,N_26574);
nand UO_2790 (O_2790,N_28365,N_28991);
or UO_2791 (O_2791,N_27237,N_29948);
and UO_2792 (O_2792,N_29514,N_25567);
nor UO_2793 (O_2793,N_25763,N_27822);
xor UO_2794 (O_2794,N_27777,N_29179);
nand UO_2795 (O_2795,N_29079,N_27320);
or UO_2796 (O_2796,N_27117,N_26247);
and UO_2797 (O_2797,N_25428,N_27723);
nand UO_2798 (O_2798,N_26245,N_25851);
or UO_2799 (O_2799,N_27942,N_28022);
nand UO_2800 (O_2800,N_28908,N_26571);
or UO_2801 (O_2801,N_28662,N_27965);
and UO_2802 (O_2802,N_27986,N_27407);
and UO_2803 (O_2803,N_25281,N_28780);
and UO_2804 (O_2804,N_27912,N_26060);
nand UO_2805 (O_2805,N_25554,N_27442);
and UO_2806 (O_2806,N_25843,N_28834);
and UO_2807 (O_2807,N_27048,N_26727);
nor UO_2808 (O_2808,N_27985,N_28327);
or UO_2809 (O_2809,N_27042,N_29406);
or UO_2810 (O_2810,N_27820,N_25897);
nand UO_2811 (O_2811,N_29093,N_25083);
or UO_2812 (O_2812,N_28246,N_29094);
or UO_2813 (O_2813,N_29207,N_29884);
xnor UO_2814 (O_2814,N_26559,N_27775);
or UO_2815 (O_2815,N_29467,N_27058);
nand UO_2816 (O_2816,N_27670,N_28323);
nand UO_2817 (O_2817,N_26923,N_29265);
or UO_2818 (O_2818,N_28425,N_26514);
and UO_2819 (O_2819,N_27174,N_27230);
and UO_2820 (O_2820,N_27160,N_28937);
nand UO_2821 (O_2821,N_29339,N_28579);
and UO_2822 (O_2822,N_29129,N_25127);
nand UO_2823 (O_2823,N_27889,N_25910);
nand UO_2824 (O_2824,N_25880,N_27841);
nand UO_2825 (O_2825,N_27558,N_26621);
and UO_2826 (O_2826,N_25851,N_26033);
nand UO_2827 (O_2827,N_26755,N_29672);
or UO_2828 (O_2828,N_28185,N_26560);
and UO_2829 (O_2829,N_29004,N_26724);
and UO_2830 (O_2830,N_26771,N_26818);
or UO_2831 (O_2831,N_25157,N_25111);
nand UO_2832 (O_2832,N_28319,N_29899);
or UO_2833 (O_2833,N_29027,N_27717);
and UO_2834 (O_2834,N_27533,N_29125);
nand UO_2835 (O_2835,N_29283,N_29723);
and UO_2836 (O_2836,N_26066,N_29910);
xnor UO_2837 (O_2837,N_27823,N_29827);
and UO_2838 (O_2838,N_27423,N_29295);
or UO_2839 (O_2839,N_26946,N_25875);
xnor UO_2840 (O_2840,N_27682,N_26488);
nand UO_2841 (O_2841,N_26077,N_29507);
or UO_2842 (O_2842,N_28753,N_29643);
or UO_2843 (O_2843,N_27770,N_26614);
nand UO_2844 (O_2844,N_25355,N_26687);
nand UO_2845 (O_2845,N_27846,N_27820);
or UO_2846 (O_2846,N_28513,N_26015);
nor UO_2847 (O_2847,N_28218,N_28932);
nor UO_2848 (O_2848,N_26846,N_25001);
nand UO_2849 (O_2849,N_28488,N_25982);
nand UO_2850 (O_2850,N_25415,N_27948);
nand UO_2851 (O_2851,N_28110,N_25268);
nor UO_2852 (O_2852,N_26663,N_28967);
nor UO_2853 (O_2853,N_28945,N_27401);
nand UO_2854 (O_2854,N_25256,N_25516);
nor UO_2855 (O_2855,N_28774,N_27063);
or UO_2856 (O_2856,N_25744,N_26353);
nand UO_2857 (O_2857,N_25134,N_27882);
or UO_2858 (O_2858,N_29123,N_25633);
xnor UO_2859 (O_2859,N_26808,N_26151);
nand UO_2860 (O_2860,N_28575,N_26308);
nand UO_2861 (O_2861,N_29334,N_26706);
nor UO_2862 (O_2862,N_29529,N_26928);
nand UO_2863 (O_2863,N_27439,N_27743);
or UO_2864 (O_2864,N_29901,N_29391);
nor UO_2865 (O_2865,N_27187,N_26656);
or UO_2866 (O_2866,N_26047,N_26855);
and UO_2867 (O_2867,N_26340,N_29960);
and UO_2868 (O_2868,N_25884,N_26039);
or UO_2869 (O_2869,N_25526,N_29671);
nor UO_2870 (O_2870,N_26370,N_25108);
xor UO_2871 (O_2871,N_29401,N_28688);
nand UO_2872 (O_2872,N_27486,N_28679);
and UO_2873 (O_2873,N_29044,N_25543);
nor UO_2874 (O_2874,N_27754,N_27851);
nor UO_2875 (O_2875,N_26939,N_25147);
nand UO_2876 (O_2876,N_29716,N_29888);
nand UO_2877 (O_2877,N_27766,N_29308);
nor UO_2878 (O_2878,N_27017,N_27912);
nand UO_2879 (O_2879,N_26490,N_25740);
xor UO_2880 (O_2880,N_29967,N_29751);
or UO_2881 (O_2881,N_28739,N_29109);
nor UO_2882 (O_2882,N_27853,N_27431);
nand UO_2883 (O_2883,N_27621,N_28245);
nand UO_2884 (O_2884,N_28126,N_29611);
or UO_2885 (O_2885,N_26373,N_27003);
nor UO_2886 (O_2886,N_25987,N_25778);
and UO_2887 (O_2887,N_25746,N_28334);
nand UO_2888 (O_2888,N_29154,N_26782);
nand UO_2889 (O_2889,N_28505,N_27269);
xor UO_2890 (O_2890,N_28695,N_28466);
and UO_2891 (O_2891,N_28029,N_29205);
and UO_2892 (O_2892,N_26836,N_29105);
nor UO_2893 (O_2893,N_25198,N_28994);
xor UO_2894 (O_2894,N_26454,N_25187);
or UO_2895 (O_2895,N_26442,N_26877);
and UO_2896 (O_2896,N_26191,N_28934);
nor UO_2897 (O_2897,N_28811,N_25799);
nand UO_2898 (O_2898,N_28385,N_26668);
or UO_2899 (O_2899,N_28978,N_28913);
or UO_2900 (O_2900,N_27198,N_27994);
xnor UO_2901 (O_2901,N_25175,N_26556);
and UO_2902 (O_2902,N_27922,N_28052);
and UO_2903 (O_2903,N_28854,N_27908);
nor UO_2904 (O_2904,N_25816,N_28385);
nor UO_2905 (O_2905,N_27774,N_28384);
nor UO_2906 (O_2906,N_26295,N_29467);
nand UO_2907 (O_2907,N_29039,N_25988);
xnor UO_2908 (O_2908,N_27125,N_28122);
nand UO_2909 (O_2909,N_26084,N_27553);
or UO_2910 (O_2910,N_27200,N_25352);
or UO_2911 (O_2911,N_28115,N_27583);
or UO_2912 (O_2912,N_29143,N_28634);
nor UO_2913 (O_2913,N_25122,N_25039);
nor UO_2914 (O_2914,N_27204,N_27052);
and UO_2915 (O_2915,N_29573,N_28448);
nand UO_2916 (O_2916,N_28089,N_27400);
or UO_2917 (O_2917,N_28849,N_26986);
nand UO_2918 (O_2918,N_26359,N_28214);
nor UO_2919 (O_2919,N_25481,N_25581);
nor UO_2920 (O_2920,N_25580,N_28391);
or UO_2921 (O_2921,N_29816,N_29390);
nand UO_2922 (O_2922,N_29940,N_28932);
nor UO_2923 (O_2923,N_28802,N_29223);
nor UO_2924 (O_2924,N_25486,N_29944);
xnor UO_2925 (O_2925,N_26182,N_26889);
and UO_2926 (O_2926,N_26345,N_27442);
nand UO_2927 (O_2927,N_26195,N_27136);
nor UO_2928 (O_2928,N_27762,N_29511);
and UO_2929 (O_2929,N_26037,N_29326);
or UO_2930 (O_2930,N_28520,N_28391);
or UO_2931 (O_2931,N_28892,N_25812);
or UO_2932 (O_2932,N_26261,N_28998);
and UO_2933 (O_2933,N_27978,N_26926);
nor UO_2934 (O_2934,N_26992,N_29620);
or UO_2935 (O_2935,N_26786,N_25830);
nor UO_2936 (O_2936,N_29282,N_28827);
nor UO_2937 (O_2937,N_29647,N_28935);
nand UO_2938 (O_2938,N_27329,N_26517);
nand UO_2939 (O_2939,N_27777,N_27176);
xor UO_2940 (O_2940,N_28366,N_27977);
xnor UO_2941 (O_2941,N_26728,N_25219);
nand UO_2942 (O_2942,N_29589,N_25712);
nand UO_2943 (O_2943,N_25394,N_28005);
or UO_2944 (O_2944,N_25272,N_25448);
nand UO_2945 (O_2945,N_25264,N_25778);
nor UO_2946 (O_2946,N_25378,N_29229);
nor UO_2947 (O_2947,N_26122,N_27534);
or UO_2948 (O_2948,N_27627,N_25753);
and UO_2949 (O_2949,N_29563,N_26521);
nor UO_2950 (O_2950,N_26733,N_25428);
or UO_2951 (O_2951,N_27669,N_27183);
nor UO_2952 (O_2952,N_26952,N_26158);
xor UO_2953 (O_2953,N_29007,N_29283);
and UO_2954 (O_2954,N_29679,N_29816);
nand UO_2955 (O_2955,N_26637,N_26621);
xor UO_2956 (O_2956,N_25544,N_26864);
nor UO_2957 (O_2957,N_26933,N_25195);
nand UO_2958 (O_2958,N_26756,N_29938);
nand UO_2959 (O_2959,N_29308,N_27049);
nand UO_2960 (O_2960,N_26900,N_25639);
or UO_2961 (O_2961,N_28608,N_28700);
nand UO_2962 (O_2962,N_25653,N_29593);
or UO_2963 (O_2963,N_28696,N_26446);
or UO_2964 (O_2964,N_26742,N_29715);
nor UO_2965 (O_2965,N_25894,N_27048);
nand UO_2966 (O_2966,N_27728,N_27220);
nor UO_2967 (O_2967,N_27582,N_26389);
nand UO_2968 (O_2968,N_27365,N_27588);
and UO_2969 (O_2969,N_27824,N_27044);
nand UO_2970 (O_2970,N_26931,N_27359);
and UO_2971 (O_2971,N_28854,N_27155);
or UO_2972 (O_2972,N_28013,N_27229);
nor UO_2973 (O_2973,N_28823,N_27024);
or UO_2974 (O_2974,N_28256,N_28406);
nand UO_2975 (O_2975,N_29233,N_29915);
or UO_2976 (O_2976,N_27243,N_28526);
xor UO_2977 (O_2977,N_26967,N_26066);
nand UO_2978 (O_2978,N_25745,N_27262);
nand UO_2979 (O_2979,N_25847,N_26220);
or UO_2980 (O_2980,N_27407,N_28885);
and UO_2981 (O_2981,N_29621,N_27935);
nand UO_2982 (O_2982,N_25221,N_26842);
and UO_2983 (O_2983,N_25509,N_28609);
xnor UO_2984 (O_2984,N_29638,N_28002);
xnor UO_2985 (O_2985,N_28753,N_28418);
and UO_2986 (O_2986,N_28986,N_25622);
and UO_2987 (O_2987,N_25947,N_26092);
nor UO_2988 (O_2988,N_26343,N_26547);
nor UO_2989 (O_2989,N_28838,N_28648);
or UO_2990 (O_2990,N_28682,N_27114);
xnor UO_2991 (O_2991,N_26663,N_28131);
xor UO_2992 (O_2992,N_26580,N_25386);
or UO_2993 (O_2993,N_26594,N_27951);
nand UO_2994 (O_2994,N_29831,N_29252);
nand UO_2995 (O_2995,N_27781,N_29544);
nand UO_2996 (O_2996,N_29187,N_25796);
and UO_2997 (O_2997,N_25908,N_27994);
nand UO_2998 (O_2998,N_25243,N_29644);
and UO_2999 (O_2999,N_28764,N_29725);
nor UO_3000 (O_3000,N_25527,N_26451);
nand UO_3001 (O_3001,N_26607,N_28751);
nor UO_3002 (O_3002,N_26294,N_26839);
or UO_3003 (O_3003,N_26446,N_27098);
or UO_3004 (O_3004,N_27485,N_25866);
nand UO_3005 (O_3005,N_28746,N_28160);
nor UO_3006 (O_3006,N_27677,N_25077);
xor UO_3007 (O_3007,N_25603,N_29867);
nand UO_3008 (O_3008,N_27191,N_25001);
nand UO_3009 (O_3009,N_26464,N_28030);
or UO_3010 (O_3010,N_26112,N_28775);
and UO_3011 (O_3011,N_27053,N_29760);
nand UO_3012 (O_3012,N_26439,N_29105);
nand UO_3013 (O_3013,N_27025,N_25193);
nor UO_3014 (O_3014,N_25734,N_27363);
nand UO_3015 (O_3015,N_29259,N_29792);
and UO_3016 (O_3016,N_26489,N_25299);
nand UO_3017 (O_3017,N_29033,N_26239);
nand UO_3018 (O_3018,N_25006,N_27560);
nor UO_3019 (O_3019,N_29813,N_29973);
or UO_3020 (O_3020,N_27550,N_28634);
nand UO_3021 (O_3021,N_29577,N_29558);
nor UO_3022 (O_3022,N_29627,N_29458);
nor UO_3023 (O_3023,N_25766,N_29546);
and UO_3024 (O_3024,N_26386,N_25017);
or UO_3025 (O_3025,N_25626,N_26987);
xnor UO_3026 (O_3026,N_28282,N_29030);
xnor UO_3027 (O_3027,N_27567,N_29552);
nor UO_3028 (O_3028,N_26777,N_26516);
nand UO_3029 (O_3029,N_26173,N_27891);
nand UO_3030 (O_3030,N_25131,N_29390);
or UO_3031 (O_3031,N_26195,N_29397);
or UO_3032 (O_3032,N_28239,N_28197);
or UO_3033 (O_3033,N_26856,N_26039);
or UO_3034 (O_3034,N_25723,N_25674);
xnor UO_3035 (O_3035,N_28286,N_28950);
and UO_3036 (O_3036,N_25377,N_25930);
or UO_3037 (O_3037,N_29451,N_28444);
xor UO_3038 (O_3038,N_26096,N_26504);
or UO_3039 (O_3039,N_25050,N_27435);
nor UO_3040 (O_3040,N_25974,N_26784);
nor UO_3041 (O_3041,N_25529,N_25393);
and UO_3042 (O_3042,N_29650,N_26618);
and UO_3043 (O_3043,N_29122,N_28675);
nor UO_3044 (O_3044,N_27306,N_28378);
nand UO_3045 (O_3045,N_27533,N_27723);
or UO_3046 (O_3046,N_29740,N_29754);
nand UO_3047 (O_3047,N_28074,N_27196);
nand UO_3048 (O_3048,N_25021,N_25924);
nand UO_3049 (O_3049,N_28140,N_26773);
or UO_3050 (O_3050,N_28003,N_26017);
nor UO_3051 (O_3051,N_28173,N_27472);
and UO_3052 (O_3052,N_25979,N_27630);
xor UO_3053 (O_3053,N_25496,N_25885);
nand UO_3054 (O_3054,N_28725,N_28570);
and UO_3055 (O_3055,N_28907,N_26345);
xnor UO_3056 (O_3056,N_27177,N_26711);
and UO_3057 (O_3057,N_26253,N_25584);
and UO_3058 (O_3058,N_28767,N_25137);
or UO_3059 (O_3059,N_26335,N_29337);
and UO_3060 (O_3060,N_28745,N_26013);
nor UO_3061 (O_3061,N_27738,N_26540);
and UO_3062 (O_3062,N_29159,N_29051);
nor UO_3063 (O_3063,N_27335,N_29975);
or UO_3064 (O_3064,N_26871,N_29170);
and UO_3065 (O_3065,N_28060,N_26337);
nor UO_3066 (O_3066,N_25948,N_25640);
nor UO_3067 (O_3067,N_28971,N_27983);
xor UO_3068 (O_3068,N_25037,N_27453);
and UO_3069 (O_3069,N_25743,N_28277);
nor UO_3070 (O_3070,N_25458,N_27378);
nor UO_3071 (O_3071,N_28024,N_28675);
nor UO_3072 (O_3072,N_28808,N_26335);
nand UO_3073 (O_3073,N_28774,N_26805);
nor UO_3074 (O_3074,N_29152,N_28544);
or UO_3075 (O_3075,N_26415,N_26664);
xor UO_3076 (O_3076,N_26520,N_26192);
nand UO_3077 (O_3077,N_29557,N_28841);
or UO_3078 (O_3078,N_26033,N_29094);
or UO_3079 (O_3079,N_27289,N_29861);
nor UO_3080 (O_3080,N_25254,N_28668);
or UO_3081 (O_3081,N_25817,N_29042);
and UO_3082 (O_3082,N_29884,N_26840);
nor UO_3083 (O_3083,N_26837,N_26409);
or UO_3084 (O_3084,N_27385,N_28427);
nor UO_3085 (O_3085,N_29010,N_27828);
or UO_3086 (O_3086,N_27189,N_29937);
and UO_3087 (O_3087,N_26756,N_29176);
xor UO_3088 (O_3088,N_26579,N_28420);
xnor UO_3089 (O_3089,N_26375,N_27425);
nor UO_3090 (O_3090,N_26811,N_28491);
or UO_3091 (O_3091,N_25858,N_25347);
or UO_3092 (O_3092,N_28731,N_26646);
and UO_3093 (O_3093,N_27310,N_26674);
and UO_3094 (O_3094,N_25237,N_26336);
and UO_3095 (O_3095,N_27250,N_27182);
nor UO_3096 (O_3096,N_26494,N_25201);
nand UO_3097 (O_3097,N_29486,N_29010);
or UO_3098 (O_3098,N_28490,N_27177);
nor UO_3099 (O_3099,N_26329,N_27249);
and UO_3100 (O_3100,N_25424,N_28167);
nand UO_3101 (O_3101,N_26713,N_29963);
nor UO_3102 (O_3102,N_28449,N_25003);
nor UO_3103 (O_3103,N_29842,N_27404);
xor UO_3104 (O_3104,N_26047,N_29626);
and UO_3105 (O_3105,N_26683,N_29271);
nand UO_3106 (O_3106,N_28531,N_27133);
nor UO_3107 (O_3107,N_26393,N_26135);
nand UO_3108 (O_3108,N_28156,N_28278);
or UO_3109 (O_3109,N_26046,N_29299);
nand UO_3110 (O_3110,N_29517,N_28211);
xnor UO_3111 (O_3111,N_28891,N_29049);
and UO_3112 (O_3112,N_26950,N_25778);
nand UO_3113 (O_3113,N_25551,N_28131);
nor UO_3114 (O_3114,N_27291,N_26396);
or UO_3115 (O_3115,N_28146,N_25912);
or UO_3116 (O_3116,N_28822,N_27462);
nor UO_3117 (O_3117,N_25154,N_25033);
nand UO_3118 (O_3118,N_27384,N_29633);
or UO_3119 (O_3119,N_27414,N_29333);
nor UO_3120 (O_3120,N_27194,N_28809);
or UO_3121 (O_3121,N_25424,N_28586);
xnor UO_3122 (O_3122,N_27658,N_27645);
nand UO_3123 (O_3123,N_27286,N_27095);
xnor UO_3124 (O_3124,N_25026,N_26376);
and UO_3125 (O_3125,N_26764,N_27751);
nor UO_3126 (O_3126,N_27488,N_25040);
nor UO_3127 (O_3127,N_27354,N_27633);
or UO_3128 (O_3128,N_28027,N_29140);
and UO_3129 (O_3129,N_27394,N_28447);
xor UO_3130 (O_3130,N_29264,N_29178);
nor UO_3131 (O_3131,N_28428,N_25251);
xnor UO_3132 (O_3132,N_27049,N_25841);
or UO_3133 (O_3133,N_28070,N_27563);
or UO_3134 (O_3134,N_25056,N_26554);
or UO_3135 (O_3135,N_29686,N_28307);
nand UO_3136 (O_3136,N_25172,N_29439);
and UO_3137 (O_3137,N_29826,N_28700);
and UO_3138 (O_3138,N_26169,N_29379);
nor UO_3139 (O_3139,N_25189,N_26608);
or UO_3140 (O_3140,N_27915,N_28034);
nor UO_3141 (O_3141,N_27431,N_28520);
and UO_3142 (O_3142,N_28201,N_27699);
xor UO_3143 (O_3143,N_25887,N_27273);
nor UO_3144 (O_3144,N_25577,N_29889);
xor UO_3145 (O_3145,N_25477,N_28462);
nor UO_3146 (O_3146,N_25156,N_27944);
and UO_3147 (O_3147,N_29936,N_28394);
or UO_3148 (O_3148,N_29093,N_27461);
nand UO_3149 (O_3149,N_28451,N_26065);
nand UO_3150 (O_3150,N_28923,N_26264);
nor UO_3151 (O_3151,N_27146,N_29976);
or UO_3152 (O_3152,N_26027,N_26430);
or UO_3153 (O_3153,N_25872,N_28863);
or UO_3154 (O_3154,N_25909,N_26956);
nand UO_3155 (O_3155,N_27205,N_25563);
or UO_3156 (O_3156,N_28328,N_27620);
and UO_3157 (O_3157,N_27458,N_29412);
and UO_3158 (O_3158,N_29253,N_28405);
nand UO_3159 (O_3159,N_25599,N_25610);
nand UO_3160 (O_3160,N_28318,N_29923);
xnor UO_3161 (O_3161,N_27217,N_27090);
nand UO_3162 (O_3162,N_28833,N_25643);
and UO_3163 (O_3163,N_28065,N_25909);
nor UO_3164 (O_3164,N_26101,N_25266);
nor UO_3165 (O_3165,N_28900,N_28242);
or UO_3166 (O_3166,N_26809,N_29876);
nand UO_3167 (O_3167,N_29998,N_29446);
nand UO_3168 (O_3168,N_28732,N_28539);
nand UO_3169 (O_3169,N_29579,N_27489);
nand UO_3170 (O_3170,N_25069,N_28814);
nand UO_3171 (O_3171,N_27595,N_29499);
nor UO_3172 (O_3172,N_25969,N_28180);
and UO_3173 (O_3173,N_27804,N_29114);
and UO_3174 (O_3174,N_29206,N_28573);
or UO_3175 (O_3175,N_28435,N_28474);
and UO_3176 (O_3176,N_26654,N_28513);
nor UO_3177 (O_3177,N_25667,N_28827);
and UO_3178 (O_3178,N_25982,N_29753);
or UO_3179 (O_3179,N_29573,N_27367);
or UO_3180 (O_3180,N_25685,N_27040);
nor UO_3181 (O_3181,N_27028,N_28892);
nor UO_3182 (O_3182,N_28135,N_25526);
nor UO_3183 (O_3183,N_27578,N_29054);
and UO_3184 (O_3184,N_28188,N_26880);
and UO_3185 (O_3185,N_27210,N_26014);
nor UO_3186 (O_3186,N_29774,N_28713);
or UO_3187 (O_3187,N_27173,N_29038);
and UO_3188 (O_3188,N_28014,N_25836);
xor UO_3189 (O_3189,N_28771,N_25768);
or UO_3190 (O_3190,N_27304,N_25022);
nor UO_3191 (O_3191,N_25374,N_28506);
or UO_3192 (O_3192,N_25082,N_26727);
nand UO_3193 (O_3193,N_25995,N_27579);
and UO_3194 (O_3194,N_25884,N_26115);
xor UO_3195 (O_3195,N_28423,N_25167);
and UO_3196 (O_3196,N_28081,N_29583);
or UO_3197 (O_3197,N_27364,N_29596);
or UO_3198 (O_3198,N_27142,N_27533);
and UO_3199 (O_3199,N_28645,N_25303);
and UO_3200 (O_3200,N_25949,N_25917);
nand UO_3201 (O_3201,N_26417,N_28417);
and UO_3202 (O_3202,N_28788,N_27009);
or UO_3203 (O_3203,N_27204,N_25435);
or UO_3204 (O_3204,N_26049,N_28149);
nand UO_3205 (O_3205,N_27357,N_26693);
nand UO_3206 (O_3206,N_26297,N_26582);
and UO_3207 (O_3207,N_29882,N_25739);
or UO_3208 (O_3208,N_29859,N_27105);
and UO_3209 (O_3209,N_27789,N_27694);
nand UO_3210 (O_3210,N_25315,N_27063);
xnor UO_3211 (O_3211,N_27804,N_28405);
and UO_3212 (O_3212,N_28354,N_28112);
and UO_3213 (O_3213,N_27723,N_28554);
nor UO_3214 (O_3214,N_27163,N_25268);
or UO_3215 (O_3215,N_29755,N_26321);
nand UO_3216 (O_3216,N_29519,N_26941);
xor UO_3217 (O_3217,N_26327,N_26401);
nand UO_3218 (O_3218,N_29451,N_25828);
or UO_3219 (O_3219,N_27726,N_27514);
nor UO_3220 (O_3220,N_25540,N_28290);
and UO_3221 (O_3221,N_25988,N_25066);
and UO_3222 (O_3222,N_25719,N_29328);
and UO_3223 (O_3223,N_29173,N_29640);
and UO_3224 (O_3224,N_26386,N_25832);
nand UO_3225 (O_3225,N_25045,N_29592);
and UO_3226 (O_3226,N_25859,N_26279);
or UO_3227 (O_3227,N_28001,N_26526);
nand UO_3228 (O_3228,N_28049,N_26150);
nor UO_3229 (O_3229,N_29492,N_28890);
and UO_3230 (O_3230,N_26310,N_25437);
nand UO_3231 (O_3231,N_27545,N_26805);
nand UO_3232 (O_3232,N_29351,N_25407);
nand UO_3233 (O_3233,N_25050,N_26925);
nand UO_3234 (O_3234,N_25149,N_29496);
nor UO_3235 (O_3235,N_29922,N_25609);
nor UO_3236 (O_3236,N_28511,N_28445);
or UO_3237 (O_3237,N_25834,N_28906);
or UO_3238 (O_3238,N_26677,N_27831);
xor UO_3239 (O_3239,N_25418,N_28769);
nand UO_3240 (O_3240,N_29565,N_25772);
and UO_3241 (O_3241,N_26508,N_25080);
nand UO_3242 (O_3242,N_25262,N_27990);
and UO_3243 (O_3243,N_27439,N_27293);
nand UO_3244 (O_3244,N_25221,N_25486);
nor UO_3245 (O_3245,N_27431,N_29771);
nor UO_3246 (O_3246,N_28141,N_28496);
nor UO_3247 (O_3247,N_28828,N_26909);
and UO_3248 (O_3248,N_25024,N_28807);
nor UO_3249 (O_3249,N_27922,N_27555);
or UO_3250 (O_3250,N_26830,N_29929);
or UO_3251 (O_3251,N_29971,N_27304);
and UO_3252 (O_3252,N_27449,N_29650);
nor UO_3253 (O_3253,N_25442,N_28465);
or UO_3254 (O_3254,N_28113,N_26594);
nor UO_3255 (O_3255,N_27565,N_28451);
or UO_3256 (O_3256,N_27299,N_28427);
nand UO_3257 (O_3257,N_26698,N_28849);
nor UO_3258 (O_3258,N_29197,N_27281);
nand UO_3259 (O_3259,N_26377,N_25773);
xor UO_3260 (O_3260,N_28558,N_25014);
nor UO_3261 (O_3261,N_25571,N_29370);
nor UO_3262 (O_3262,N_26034,N_29117);
or UO_3263 (O_3263,N_27325,N_25112);
nor UO_3264 (O_3264,N_29461,N_29971);
and UO_3265 (O_3265,N_25569,N_25462);
nand UO_3266 (O_3266,N_28900,N_28771);
and UO_3267 (O_3267,N_28506,N_26644);
or UO_3268 (O_3268,N_25124,N_26140);
and UO_3269 (O_3269,N_28165,N_29706);
nor UO_3270 (O_3270,N_29367,N_28667);
nand UO_3271 (O_3271,N_25053,N_28244);
or UO_3272 (O_3272,N_27844,N_25649);
and UO_3273 (O_3273,N_28547,N_26716);
and UO_3274 (O_3274,N_26746,N_27483);
or UO_3275 (O_3275,N_27349,N_25718);
and UO_3276 (O_3276,N_26299,N_28198);
or UO_3277 (O_3277,N_27049,N_27568);
nand UO_3278 (O_3278,N_26806,N_26245);
nand UO_3279 (O_3279,N_27140,N_26091);
nand UO_3280 (O_3280,N_27220,N_26329);
nor UO_3281 (O_3281,N_27426,N_28992);
nor UO_3282 (O_3282,N_27832,N_28562);
xor UO_3283 (O_3283,N_27543,N_27615);
nand UO_3284 (O_3284,N_26157,N_28806);
nor UO_3285 (O_3285,N_29168,N_28859);
and UO_3286 (O_3286,N_25897,N_27867);
and UO_3287 (O_3287,N_25481,N_29999);
nand UO_3288 (O_3288,N_25459,N_29092);
nor UO_3289 (O_3289,N_27166,N_28484);
nor UO_3290 (O_3290,N_25990,N_29317);
nand UO_3291 (O_3291,N_27288,N_27688);
nand UO_3292 (O_3292,N_29023,N_29684);
nand UO_3293 (O_3293,N_28709,N_29607);
nand UO_3294 (O_3294,N_28804,N_27831);
nor UO_3295 (O_3295,N_28184,N_27976);
or UO_3296 (O_3296,N_26971,N_29407);
nand UO_3297 (O_3297,N_28047,N_25475);
nor UO_3298 (O_3298,N_27059,N_29381);
and UO_3299 (O_3299,N_26720,N_29645);
and UO_3300 (O_3300,N_25084,N_25648);
and UO_3301 (O_3301,N_29389,N_28960);
and UO_3302 (O_3302,N_25395,N_25739);
nand UO_3303 (O_3303,N_27959,N_25475);
nand UO_3304 (O_3304,N_29753,N_28409);
or UO_3305 (O_3305,N_26102,N_26295);
nand UO_3306 (O_3306,N_27113,N_25911);
nor UO_3307 (O_3307,N_27937,N_28685);
nand UO_3308 (O_3308,N_29801,N_29214);
xor UO_3309 (O_3309,N_27515,N_27196);
nand UO_3310 (O_3310,N_28554,N_29220);
and UO_3311 (O_3311,N_27392,N_28669);
nand UO_3312 (O_3312,N_27090,N_28139);
and UO_3313 (O_3313,N_27693,N_25738);
xor UO_3314 (O_3314,N_28034,N_29235);
or UO_3315 (O_3315,N_25843,N_26641);
or UO_3316 (O_3316,N_25014,N_26111);
nand UO_3317 (O_3317,N_29253,N_27481);
and UO_3318 (O_3318,N_27490,N_29592);
nor UO_3319 (O_3319,N_27669,N_26919);
or UO_3320 (O_3320,N_27590,N_29507);
or UO_3321 (O_3321,N_29061,N_27470);
and UO_3322 (O_3322,N_27592,N_26956);
or UO_3323 (O_3323,N_25578,N_27933);
nor UO_3324 (O_3324,N_28868,N_29428);
or UO_3325 (O_3325,N_27563,N_29685);
nor UO_3326 (O_3326,N_25528,N_27654);
nand UO_3327 (O_3327,N_27908,N_25142);
xor UO_3328 (O_3328,N_26052,N_27691);
nor UO_3329 (O_3329,N_26948,N_26733);
nor UO_3330 (O_3330,N_27038,N_29882);
xor UO_3331 (O_3331,N_29238,N_27259);
and UO_3332 (O_3332,N_29754,N_27211);
or UO_3333 (O_3333,N_25362,N_28358);
nand UO_3334 (O_3334,N_26128,N_29517);
and UO_3335 (O_3335,N_25004,N_28357);
or UO_3336 (O_3336,N_27308,N_28841);
or UO_3337 (O_3337,N_25594,N_29545);
nor UO_3338 (O_3338,N_25773,N_25429);
nand UO_3339 (O_3339,N_29544,N_26893);
nand UO_3340 (O_3340,N_29802,N_29403);
and UO_3341 (O_3341,N_29859,N_27754);
and UO_3342 (O_3342,N_25464,N_28768);
or UO_3343 (O_3343,N_27884,N_29605);
nor UO_3344 (O_3344,N_29186,N_28333);
or UO_3345 (O_3345,N_27673,N_26568);
nand UO_3346 (O_3346,N_27648,N_28078);
or UO_3347 (O_3347,N_26049,N_26801);
nor UO_3348 (O_3348,N_26694,N_27005);
xnor UO_3349 (O_3349,N_28458,N_28376);
xor UO_3350 (O_3350,N_25374,N_25249);
and UO_3351 (O_3351,N_28641,N_29181);
xor UO_3352 (O_3352,N_26419,N_29939);
and UO_3353 (O_3353,N_26736,N_25364);
or UO_3354 (O_3354,N_25968,N_29273);
and UO_3355 (O_3355,N_25051,N_25566);
nand UO_3356 (O_3356,N_27841,N_27518);
or UO_3357 (O_3357,N_28097,N_29888);
xnor UO_3358 (O_3358,N_29792,N_27769);
or UO_3359 (O_3359,N_25801,N_29420);
and UO_3360 (O_3360,N_26199,N_26403);
and UO_3361 (O_3361,N_28850,N_27974);
nand UO_3362 (O_3362,N_29195,N_27956);
and UO_3363 (O_3363,N_25253,N_29411);
or UO_3364 (O_3364,N_27501,N_29368);
and UO_3365 (O_3365,N_28278,N_28648);
nor UO_3366 (O_3366,N_25537,N_25888);
and UO_3367 (O_3367,N_29125,N_27251);
nand UO_3368 (O_3368,N_27406,N_25390);
nor UO_3369 (O_3369,N_28231,N_25661);
nor UO_3370 (O_3370,N_28713,N_29203);
nor UO_3371 (O_3371,N_27023,N_25421);
nor UO_3372 (O_3372,N_27789,N_26830);
xor UO_3373 (O_3373,N_27444,N_26737);
xnor UO_3374 (O_3374,N_29978,N_28779);
and UO_3375 (O_3375,N_28574,N_25716);
and UO_3376 (O_3376,N_28142,N_27059);
nor UO_3377 (O_3377,N_28582,N_29341);
nand UO_3378 (O_3378,N_28637,N_25380);
or UO_3379 (O_3379,N_28511,N_25741);
nand UO_3380 (O_3380,N_26369,N_29881);
nand UO_3381 (O_3381,N_28354,N_29436);
and UO_3382 (O_3382,N_25657,N_26304);
nor UO_3383 (O_3383,N_27999,N_28767);
nand UO_3384 (O_3384,N_29624,N_28908);
or UO_3385 (O_3385,N_28162,N_25865);
nand UO_3386 (O_3386,N_28815,N_28201);
and UO_3387 (O_3387,N_25934,N_29851);
nor UO_3388 (O_3388,N_29407,N_29702);
or UO_3389 (O_3389,N_26020,N_29110);
nor UO_3390 (O_3390,N_26318,N_28493);
and UO_3391 (O_3391,N_28021,N_29795);
nand UO_3392 (O_3392,N_25921,N_28394);
and UO_3393 (O_3393,N_27864,N_28489);
nor UO_3394 (O_3394,N_27536,N_29598);
or UO_3395 (O_3395,N_25476,N_26383);
or UO_3396 (O_3396,N_28846,N_29631);
nor UO_3397 (O_3397,N_25485,N_27925);
nand UO_3398 (O_3398,N_28527,N_26439);
nor UO_3399 (O_3399,N_26881,N_27115);
and UO_3400 (O_3400,N_26896,N_29261);
or UO_3401 (O_3401,N_26923,N_25080);
or UO_3402 (O_3402,N_26729,N_25274);
nand UO_3403 (O_3403,N_28934,N_28213);
nand UO_3404 (O_3404,N_29379,N_28711);
and UO_3405 (O_3405,N_29511,N_25819);
nand UO_3406 (O_3406,N_26159,N_26767);
nor UO_3407 (O_3407,N_29795,N_28853);
or UO_3408 (O_3408,N_27742,N_25965);
or UO_3409 (O_3409,N_25419,N_25515);
nand UO_3410 (O_3410,N_29578,N_26303);
and UO_3411 (O_3411,N_27833,N_28597);
nor UO_3412 (O_3412,N_27753,N_29579);
and UO_3413 (O_3413,N_26099,N_26449);
or UO_3414 (O_3414,N_26534,N_26157);
or UO_3415 (O_3415,N_29173,N_29241);
nand UO_3416 (O_3416,N_27111,N_28147);
xor UO_3417 (O_3417,N_29298,N_25336);
nor UO_3418 (O_3418,N_26908,N_26410);
xor UO_3419 (O_3419,N_26800,N_28022);
or UO_3420 (O_3420,N_26928,N_29465);
and UO_3421 (O_3421,N_25188,N_28615);
or UO_3422 (O_3422,N_26268,N_25367);
and UO_3423 (O_3423,N_26629,N_25994);
nand UO_3424 (O_3424,N_26435,N_28426);
and UO_3425 (O_3425,N_28399,N_29161);
nor UO_3426 (O_3426,N_25729,N_28548);
nand UO_3427 (O_3427,N_27808,N_26021);
nand UO_3428 (O_3428,N_26233,N_29444);
nor UO_3429 (O_3429,N_26781,N_25727);
and UO_3430 (O_3430,N_28786,N_28249);
and UO_3431 (O_3431,N_27133,N_26131);
nor UO_3432 (O_3432,N_27508,N_26972);
nand UO_3433 (O_3433,N_29953,N_25312);
nor UO_3434 (O_3434,N_26442,N_29699);
and UO_3435 (O_3435,N_29932,N_26836);
and UO_3436 (O_3436,N_27874,N_25503);
or UO_3437 (O_3437,N_27042,N_28145);
or UO_3438 (O_3438,N_28331,N_29103);
or UO_3439 (O_3439,N_25977,N_25200);
and UO_3440 (O_3440,N_25154,N_25276);
nand UO_3441 (O_3441,N_25431,N_27098);
nor UO_3442 (O_3442,N_28359,N_29948);
and UO_3443 (O_3443,N_27055,N_27342);
or UO_3444 (O_3444,N_28539,N_28731);
nand UO_3445 (O_3445,N_28466,N_28339);
nor UO_3446 (O_3446,N_25633,N_29981);
xor UO_3447 (O_3447,N_25868,N_26172);
or UO_3448 (O_3448,N_25618,N_27007);
or UO_3449 (O_3449,N_29015,N_26599);
nor UO_3450 (O_3450,N_26659,N_28167);
and UO_3451 (O_3451,N_29099,N_28293);
nand UO_3452 (O_3452,N_28695,N_28368);
or UO_3453 (O_3453,N_26771,N_29057);
and UO_3454 (O_3454,N_27320,N_26304);
nor UO_3455 (O_3455,N_27207,N_29230);
nand UO_3456 (O_3456,N_29440,N_28267);
nand UO_3457 (O_3457,N_28690,N_29173);
xor UO_3458 (O_3458,N_25185,N_28924);
xor UO_3459 (O_3459,N_27741,N_29449);
and UO_3460 (O_3460,N_25632,N_25617);
or UO_3461 (O_3461,N_25911,N_29074);
or UO_3462 (O_3462,N_27164,N_28375);
nor UO_3463 (O_3463,N_29517,N_27763);
nor UO_3464 (O_3464,N_27637,N_29858);
nand UO_3465 (O_3465,N_28162,N_25292);
or UO_3466 (O_3466,N_27961,N_25822);
nand UO_3467 (O_3467,N_27797,N_26651);
nand UO_3468 (O_3468,N_25263,N_25504);
and UO_3469 (O_3469,N_27735,N_29224);
or UO_3470 (O_3470,N_28462,N_28634);
nand UO_3471 (O_3471,N_27740,N_29644);
and UO_3472 (O_3472,N_29655,N_28746);
nand UO_3473 (O_3473,N_25686,N_27948);
or UO_3474 (O_3474,N_27079,N_29415);
or UO_3475 (O_3475,N_28143,N_28113);
and UO_3476 (O_3476,N_29277,N_27721);
or UO_3477 (O_3477,N_29802,N_29331);
and UO_3478 (O_3478,N_29788,N_27127);
and UO_3479 (O_3479,N_28890,N_25957);
nand UO_3480 (O_3480,N_29181,N_29342);
xnor UO_3481 (O_3481,N_27584,N_27794);
nor UO_3482 (O_3482,N_25151,N_26419);
and UO_3483 (O_3483,N_25444,N_25520);
or UO_3484 (O_3484,N_27801,N_28674);
or UO_3485 (O_3485,N_29014,N_27037);
nor UO_3486 (O_3486,N_28291,N_26884);
and UO_3487 (O_3487,N_26996,N_27036);
nand UO_3488 (O_3488,N_27397,N_29159);
nand UO_3489 (O_3489,N_27112,N_27644);
or UO_3490 (O_3490,N_26060,N_26118);
nor UO_3491 (O_3491,N_25671,N_28143);
nand UO_3492 (O_3492,N_27268,N_25988);
nor UO_3493 (O_3493,N_27097,N_29011);
nor UO_3494 (O_3494,N_29920,N_25481);
or UO_3495 (O_3495,N_26527,N_27224);
and UO_3496 (O_3496,N_26887,N_28748);
or UO_3497 (O_3497,N_25850,N_26743);
nand UO_3498 (O_3498,N_28128,N_28374);
or UO_3499 (O_3499,N_25278,N_29130);
endmodule