module basic_2000_20000_2500_20_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
or U0 (N_0,In_796,In_714);
and U1 (N_1,In_742,In_385);
and U2 (N_2,In_1657,In_460);
nand U3 (N_3,In_1948,In_1502);
and U4 (N_4,In_1229,In_1631);
xnor U5 (N_5,In_1267,In_336);
xnor U6 (N_6,In_415,In_773);
nand U7 (N_7,In_1049,In_761);
or U8 (N_8,In_456,In_930);
nor U9 (N_9,In_708,In_919);
and U10 (N_10,In_1845,In_366);
nand U11 (N_11,In_795,In_484);
xor U12 (N_12,In_896,In_1121);
nand U13 (N_13,In_1218,In_1817);
xnor U14 (N_14,In_1306,In_1658);
and U15 (N_15,In_443,In_150);
or U16 (N_16,In_269,In_1540);
or U17 (N_17,In_1716,In_1142);
nor U18 (N_18,In_1268,In_405);
nand U19 (N_19,In_1365,In_267);
nor U20 (N_20,In_592,In_662);
or U21 (N_21,In_1271,In_832);
nand U22 (N_22,In_934,In_33);
or U23 (N_23,In_334,In_1659);
and U24 (N_24,In_469,In_684);
nor U25 (N_25,In_863,In_1450);
xnor U26 (N_26,In_120,In_928);
or U27 (N_27,In_828,In_1969);
nand U28 (N_28,In_1602,In_1685);
and U29 (N_29,In_1204,In_817);
and U30 (N_30,In_1115,In_360);
xor U31 (N_31,In_1927,In_1105);
and U32 (N_32,In_1864,In_154);
nand U33 (N_33,In_864,In_1663);
and U34 (N_34,In_1992,In_1059);
and U35 (N_35,In_1582,In_1124);
and U36 (N_36,In_1174,In_1025);
or U37 (N_37,In_537,In_1839);
or U38 (N_38,In_993,In_3);
nand U39 (N_39,In_1870,In_1054);
nor U40 (N_40,In_185,In_705);
xor U41 (N_41,In_1057,In_706);
and U42 (N_42,In_1607,In_1897);
nand U43 (N_43,In_358,In_1606);
xor U44 (N_44,In_1113,In_200);
and U45 (N_45,In_1230,In_695);
or U46 (N_46,In_1064,In_441);
nor U47 (N_47,In_339,In_1881);
or U48 (N_48,In_1160,In_306);
nand U49 (N_49,In_1273,In_1489);
nor U50 (N_50,In_442,In_1186);
nand U51 (N_51,In_99,In_1624);
and U52 (N_52,In_81,In_985);
and U53 (N_53,In_270,In_965);
nand U54 (N_54,In_899,In_1287);
or U55 (N_55,In_80,In_229);
xnor U56 (N_56,In_1648,In_904);
and U57 (N_57,In_858,In_1519);
nor U58 (N_58,In_819,In_660);
and U59 (N_59,In_1537,In_390);
xnor U60 (N_60,In_861,In_21);
nand U61 (N_61,In_1786,In_1783);
xnor U62 (N_62,In_1962,In_472);
or U63 (N_63,In_1684,In_74);
and U64 (N_64,In_918,In_1437);
xnor U65 (N_65,In_398,In_77);
and U66 (N_66,In_1043,In_218);
xor U67 (N_67,In_375,In_184);
and U68 (N_68,In_196,In_1303);
nor U69 (N_69,In_679,In_1534);
or U70 (N_70,In_293,In_807);
nor U71 (N_71,In_1797,In_1697);
and U72 (N_72,In_1690,In_1368);
xnor U73 (N_73,In_1382,In_1076);
nand U74 (N_74,In_1510,In_1411);
or U75 (N_75,In_1472,In_1682);
nand U76 (N_76,In_1676,In_1248);
nand U77 (N_77,In_1806,In_255);
nor U78 (N_78,In_402,In_1002);
nor U79 (N_79,In_1900,In_1921);
nand U80 (N_80,In_459,In_1629);
xor U81 (N_81,In_1324,In_1498);
and U82 (N_82,In_717,In_173);
or U83 (N_83,In_739,In_31);
or U84 (N_84,In_355,In_439);
nand U85 (N_85,In_254,In_300);
nand U86 (N_86,In_1622,In_1162);
xor U87 (N_87,In_161,In_683);
or U88 (N_88,In_1448,In_1392);
xnor U89 (N_89,In_1449,In_1913);
nand U90 (N_90,In_1082,In_1945);
xnor U91 (N_91,In_91,In_356);
xnor U92 (N_92,In_539,In_992);
xor U93 (N_93,In_802,In_926);
or U94 (N_94,In_1352,In_1335);
xnor U95 (N_95,In_948,In_1844);
and U96 (N_96,In_722,In_1099);
or U97 (N_97,In_230,In_117);
nand U98 (N_98,In_262,In_1095);
nor U99 (N_99,In_1356,In_1963);
nand U100 (N_100,In_32,In_462);
nor U101 (N_101,In_1348,In_853);
or U102 (N_102,In_535,In_954);
nor U103 (N_103,In_492,In_1547);
nand U104 (N_104,In_326,In_118);
nor U105 (N_105,In_1092,In_1868);
xnor U106 (N_106,In_105,In_561);
and U107 (N_107,In_1832,In_1642);
xor U108 (N_108,In_503,In_885);
nand U109 (N_109,In_1233,In_1019);
and U110 (N_110,In_40,In_801);
or U111 (N_111,In_1484,In_1102);
or U112 (N_112,In_1778,In_1822);
nand U113 (N_113,In_482,In_1998);
nor U114 (N_114,In_340,In_933);
or U115 (N_115,In_842,In_1120);
xor U116 (N_116,In_1349,In_1184);
xor U117 (N_117,In_639,In_238);
and U118 (N_118,In_157,In_1702);
nor U119 (N_119,In_127,In_1422);
nand U120 (N_120,In_202,In_1570);
or U121 (N_121,In_1488,In_711);
nand U122 (N_122,In_1736,In_752);
and U123 (N_123,In_383,In_97);
nand U124 (N_124,In_524,In_677);
xnor U125 (N_125,In_550,In_1617);
or U126 (N_126,In_1242,In_1136);
and U127 (N_127,In_1545,In_1704);
xnor U128 (N_128,In_1668,In_1699);
or U129 (N_129,In_1956,In_1650);
nor U130 (N_130,In_1444,In_1746);
xor U131 (N_131,In_406,In_692);
nand U132 (N_132,In_1334,In_1987);
xnor U133 (N_133,In_19,In_760);
xnor U134 (N_134,In_1785,In_1048);
and U135 (N_135,In_151,In_653);
and U136 (N_136,In_1988,In_1666);
xor U137 (N_137,In_1143,In_1360);
or U138 (N_138,In_556,In_1199);
nand U139 (N_139,In_1752,In_1386);
xor U140 (N_140,In_75,In_1183);
or U141 (N_141,In_155,In_892);
xnor U142 (N_142,In_477,In_746);
nor U143 (N_143,In_69,In_490);
nand U144 (N_144,In_1427,In_995);
xnor U145 (N_145,In_1369,In_781);
or U146 (N_146,In_106,In_922);
nand U147 (N_147,In_302,In_823);
xor U148 (N_148,In_1171,In_1879);
and U149 (N_149,In_49,In_1880);
and U150 (N_150,In_1140,In_1373);
xor U151 (N_151,In_1920,In_7);
xor U152 (N_152,In_720,In_1601);
nand U153 (N_153,In_1380,In_843);
xor U154 (N_154,In_46,In_295);
or U155 (N_155,In_1563,In_1304);
xor U156 (N_156,In_1342,In_1807);
and U157 (N_157,In_573,In_1841);
xnor U158 (N_158,In_657,In_1029);
nand U159 (N_159,In_841,In_290);
or U160 (N_160,In_371,In_454);
and U161 (N_161,In_719,In_675);
xor U162 (N_162,In_1588,In_1770);
nor U163 (N_163,In_614,In_215);
or U164 (N_164,In_1769,In_1168);
nor U165 (N_165,In_1968,In_1718);
nor U166 (N_166,In_1645,In_1714);
nand U167 (N_167,In_478,In_1237);
nor U168 (N_168,In_710,In_1730);
xnor U169 (N_169,In_17,In_1577);
nand U170 (N_170,In_531,In_1196);
nand U171 (N_171,In_645,In_1083);
xor U172 (N_172,In_13,In_227);
nand U173 (N_173,In_451,In_1201);
xor U174 (N_174,In_652,In_1947);
xor U175 (N_175,In_1619,In_808);
and U176 (N_176,In_1006,In_749);
xnor U177 (N_177,In_1397,In_980);
xnor U178 (N_178,In_538,In_135);
or U179 (N_179,In_586,In_775);
xnor U180 (N_180,In_310,In_1282);
xor U181 (N_181,In_1035,In_1493);
nor U182 (N_182,In_1784,In_1293);
and U183 (N_183,In_1410,In_317);
or U184 (N_184,In_1141,In_1876);
xor U185 (N_185,In_681,In_1132);
nor U186 (N_186,In_1202,In_1023);
xnor U187 (N_187,In_569,In_805);
and U188 (N_188,In_1917,In_1371);
and U189 (N_189,In_1111,In_102);
nand U190 (N_190,In_663,In_1340);
nand U191 (N_191,In_630,In_1464);
or U192 (N_192,In_1852,In_1131);
or U193 (N_193,In_601,In_180);
and U194 (N_194,In_174,In_1991);
nor U195 (N_195,In_1362,In_891);
xor U196 (N_196,In_1753,In_1965);
nand U197 (N_197,In_1625,In_380);
nand U198 (N_198,In_1401,In_1742);
and U199 (N_199,In_1564,In_1862);
or U200 (N_200,In_528,In_836);
nor U201 (N_201,In_214,In_1937);
and U202 (N_202,In_163,In_643);
xnor U203 (N_203,In_359,In_1527);
xor U204 (N_204,In_1418,In_647);
and U205 (N_205,In_1055,In_571);
and U206 (N_206,In_430,In_1614);
nor U207 (N_207,In_1548,In_1737);
or U208 (N_208,In_838,In_1037);
nand U209 (N_209,In_186,In_821);
xnor U210 (N_210,In_1310,In_755);
nand U211 (N_211,In_327,In_789);
nor U212 (N_212,In_1695,In_1262);
nor U213 (N_213,In_622,In_1311);
nor U214 (N_214,In_580,In_597);
xnor U215 (N_215,In_792,In_104);
xor U216 (N_216,In_1958,In_551);
and U217 (N_217,In_1318,In_975);
and U218 (N_218,In_713,In_1731);
nand U219 (N_219,In_712,In_665);
or U220 (N_220,In_1150,In_446);
and U221 (N_221,In_14,In_697);
nor U222 (N_222,In_1180,In_994);
and U223 (N_223,In_1949,In_486);
nand U224 (N_224,In_1156,In_1930);
nor U225 (N_225,In_707,In_208);
nor U226 (N_226,In_266,In_1056);
nor U227 (N_227,In_481,In_1538);
and U228 (N_228,In_1439,In_164);
or U229 (N_229,In_1677,In_670);
xor U230 (N_230,In_1565,In_1584);
xnor U231 (N_231,In_1872,In_136);
xor U232 (N_232,In_1652,In_1686);
xor U233 (N_233,In_1261,In_1573);
and U234 (N_234,In_499,In_878);
or U235 (N_235,In_1317,In_1713);
or U236 (N_236,In_748,In_55);
xnor U237 (N_237,In_198,In_1278);
and U238 (N_238,In_1744,In_1873);
nand U239 (N_239,In_845,In_955);
xor U240 (N_240,In_1192,In_1891);
nand U241 (N_241,In_192,In_1416);
xor U242 (N_242,In_242,In_1728);
nand U243 (N_243,In_834,In_991);
or U244 (N_244,In_1398,In_1031);
nor U245 (N_245,In_455,In_433);
nor U246 (N_246,In_1989,In_1331);
or U247 (N_247,In_541,In_89);
xnor U248 (N_248,In_984,In_536);
and U249 (N_249,In_160,In_134);
nor U250 (N_250,In_1587,In_693);
or U251 (N_251,In_1018,In_1126);
xnor U252 (N_252,In_680,In_1152);
nor U253 (N_253,In_600,In_53);
and U254 (N_254,In_564,In_217);
or U255 (N_255,In_47,In_626);
nand U256 (N_256,In_771,In_1000);
nand U257 (N_257,In_357,In_1297);
and U258 (N_258,In_354,In_696);
nand U259 (N_259,In_401,In_577);
nor U260 (N_260,In_171,In_1263);
and U261 (N_261,In_1066,In_1768);
and U262 (N_262,In_273,In_458);
or U263 (N_263,In_1119,In_1253);
or U264 (N_264,In_566,In_1276);
xnor U265 (N_265,In_1496,In_119);
or U266 (N_266,In_1265,In_1281);
or U267 (N_267,In_855,In_465);
or U268 (N_268,In_1466,In_1129);
nor U269 (N_269,In_352,In_1012);
nor U270 (N_270,In_1720,In_1687);
or U271 (N_271,In_1015,In_778);
or U272 (N_272,In_608,In_282);
nand U273 (N_273,In_931,In_9);
xnor U274 (N_274,In_1457,In_1800);
nor U275 (N_275,In_1755,In_888);
nor U276 (N_276,In_263,In_1553);
xnor U277 (N_277,In_534,In_1478);
xor U278 (N_278,In_1557,In_1258);
nand U279 (N_279,In_413,In_66);
nor U280 (N_280,In_235,In_400);
xnor U281 (N_281,In_318,In_1093);
and U282 (N_282,In_903,In_189);
xnor U283 (N_283,In_743,In_168);
or U284 (N_284,In_1641,In_1298);
xnor U285 (N_285,In_865,In_1300);
and U286 (N_286,In_595,In_1147);
and U287 (N_287,In_1618,In_350);
xnor U288 (N_288,In_392,In_480);
and U289 (N_289,In_1793,In_1149);
or U290 (N_290,In_1995,In_822);
xor U291 (N_291,In_924,In_1222);
nand U292 (N_292,In_1173,In_598);
and U293 (N_293,In_1389,In_624);
nand U294 (N_294,In_374,In_474);
and U295 (N_295,In_1234,In_1094);
and U296 (N_296,In_113,In_314);
and U297 (N_297,In_734,In_1109);
nand U298 (N_298,In_241,In_1080);
and U299 (N_299,In_312,In_345);
nor U300 (N_300,In_784,In_1471);
xor U301 (N_301,In_1904,In_1486);
xnor U302 (N_302,In_297,In_309);
or U303 (N_303,In_36,In_848);
nor U304 (N_304,In_389,In_1100);
nand U305 (N_305,In_814,In_1166);
or U306 (N_306,In_724,In_1309);
nand U307 (N_307,In_8,In_1791);
or U308 (N_308,In_615,In_835);
nor U309 (N_309,In_518,In_1578);
nand U310 (N_310,In_436,In_116);
or U311 (N_311,In_1693,In_1223);
nor U312 (N_312,In_876,In_1435);
nor U313 (N_313,In_1283,In_977);
nor U314 (N_314,In_1594,In_1698);
and U315 (N_315,In_1827,In_1857);
and U316 (N_316,In_915,In_1421);
nand U317 (N_317,In_1347,In_1581);
or U318 (N_318,In_353,In_741);
and U319 (N_319,In_1819,In_50);
or U320 (N_320,In_223,In_783);
nor U321 (N_321,In_377,In_41);
and U322 (N_322,In_974,In_1420);
xor U323 (N_323,In_195,In_289);
nor U324 (N_324,In_1345,In_1837);
nand U325 (N_325,In_893,In_234);
or U326 (N_326,In_611,In_256);
xnor U327 (N_327,In_428,In_1723);
or U328 (N_328,In_1976,In_1754);
and U329 (N_329,In_990,In_1532);
nand U330 (N_330,In_1032,In_424);
nand U331 (N_331,In_671,In_1586);
and U332 (N_332,In_1112,In_635);
or U333 (N_333,In_471,In_1462);
and U334 (N_334,In_1378,In_169);
or U335 (N_335,In_634,In_346);
nor U336 (N_336,In_396,In_1787);
and U337 (N_337,In_1799,In_476);
nand U338 (N_338,In_912,In_1660);
and U339 (N_339,In_938,In_1801);
and U340 (N_340,In_1933,In_1357);
nand U341 (N_341,In_616,In_6);
nand U342 (N_342,In_1951,In_347);
xnor U343 (N_343,In_1216,In_1773);
and U344 (N_344,In_421,In_1321);
or U345 (N_345,In_1181,In_570);
nand U346 (N_346,In_132,In_475);
and U347 (N_347,In_957,In_756);
nand U348 (N_348,In_763,In_610);
nor U349 (N_349,In_372,In_1740);
or U350 (N_350,In_1203,In_26);
nor U351 (N_351,In_1393,In_594);
nor U352 (N_352,In_1200,In_1302);
nand U353 (N_353,In_232,In_1157);
or U354 (N_354,In_1005,In_941);
or U355 (N_355,In_1259,In_798);
and U356 (N_356,In_258,In_762);
nand U357 (N_357,In_1669,In_747);
xnor U358 (N_358,In_1299,In_1932);
nand U359 (N_359,In_895,In_496);
xor U360 (N_360,In_1016,In_628);
nor U361 (N_361,In_517,In_873);
nor U362 (N_362,In_1155,In_505);
and U363 (N_363,In_45,In_1408);
xor U364 (N_364,In_72,In_799);
or U365 (N_365,In_1733,In_1503);
or U366 (N_366,In_250,In_603);
nand U367 (N_367,In_1114,In_1027);
and U368 (N_368,In_1855,In_1853);
and U369 (N_369,In_1325,In_1425);
xnor U370 (N_370,In_177,In_1811);
nor U371 (N_371,In_1456,In_1851);
or U372 (N_372,In_1721,In_498);
or U373 (N_373,In_1243,In_1603);
xnor U374 (N_374,In_76,In_1701);
nor U375 (N_375,In_1159,In_1705);
or U376 (N_376,In_1465,In_125);
nand U377 (N_377,In_1344,In_563);
nor U378 (N_378,In_64,In_613);
and U379 (N_379,In_1122,In_1164);
or U380 (N_380,In_277,In_1759);
and U381 (N_381,In_1492,In_56);
or U382 (N_382,In_1320,In_379);
or U383 (N_383,In_1003,In_709);
xnor U384 (N_384,In_1280,In_58);
nor U385 (N_385,In_726,In_1020);
nor U386 (N_386,In_399,In_1836);
xnor U387 (N_387,In_582,In_1533);
or U388 (N_388,In_549,In_27);
nand U389 (N_389,In_44,In_629);
or U390 (N_390,In_137,In_1172);
or U391 (N_391,In_252,In_987);
nor U392 (N_392,In_1546,In_579);
nand U393 (N_393,In_114,In_514);
nor U394 (N_394,In_1148,In_387);
or U395 (N_395,In_1419,In_1063);
and U396 (N_396,In_1315,In_1580);
and U397 (N_397,In_1907,In_1980);
or U398 (N_398,In_388,In_770);
xor U399 (N_399,In_1552,In_1058);
and U400 (N_400,In_946,In_108);
or U401 (N_401,In_236,In_1810);
xor U402 (N_402,In_1961,In_159);
and U403 (N_403,In_682,In_212);
nor U404 (N_404,In_690,In_1888);
or U405 (N_405,In_1828,In_793);
nor U406 (N_406,In_461,In_249);
xnor U407 (N_407,In_1972,In_1826);
nor U408 (N_408,In_632,In_1116);
or U409 (N_409,In_627,In_1558);
nand U410 (N_410,In_1308,In_1207);
and U411 (N_411,In_1908,In_193);
and U412 (N_412,In_1633,In_1091);
nand U413 (N_413,In_916,In_856);
xor U414 (N_414,In_1643,In_1327);
and U415 (N_415,In_338,In_1191);
xnor U416 (N_416,In_1902,In_434);
nand U417 (N_417,In_544,In_905);
nor U418 (N_418,In_1764,In_907);
nand U419 (N_419,In_1217,In_1244);
and U420 (N_420,In_156,In_1404);
or U421 (N_421,In_153,In_1487);
nor U422 (N_422,In_248,In_1758);
nand U423 (N_423,In_1396,In_1459);
nor U424 (N_424,In_1381,In_1734);
or U425 (N_425,In_138,In_431);
and U426 (N_426,In_844,In_1556);
nor U427 (N_427,In_175,In_1743);
nor U428 (N_428,In_1225,In_88);
nor U429 (N_429,In_902,In_1052);
nor U430 (N_430,In_1585,In_1898);
xor U431 (N_431,In_523,In_1915);
xnor U432 (N_432,In_1906,In_1313);
or U433 (N_433,In_812,In_1535);
nand U434 (N_434,In_606,In_1739);
or U435 (N_435,In_849,In_857);
nor U436 (N_436,In_1195,In_1509);
or U437 (N_437,In_479,In_368);
and U438 (N_438,In_207,In_1615);
and U439 (N_439,In_1964,In_1860);
nor U440 (N_440,In_1610,In_1394);
nor U441 (N_441,In_292,In_605);
and U442 (N_442,In_1804,In_1803);
nor U443 (N_443,In_640,In_1353);
xnor U444 (N_444,In_1228,In_877);
nand U445 (N_445,In_131,In_699);
and U446 (N_446,In_25,In_147);
nand U447 (N_447,In_34,In_1205);
xor U448 (N_448,In_315,In_145);
xnor U449 (N_449,In_687,In_1929);
and U450 (N_450,In_1024,In_378);
nor U451 (N_451,In_1326,In_1825);
nand U452 (N_452,In_553,In_1220);
nor U453 (N_453,In_1361,In_1214);
and U454 (N_454,In_285,In_1446);
or U455 (N_455,In_1522,In_829);
and U456 (N_456,In_109,In_502);
or U457 (N_457,In_1461,In_811);
nor U458 (N_458,In_976,In_167);
or U459 (N_459,In_759,In_927);
and U460 (N_460,In_572,In_429);
xor U461 (N_461,In_565,In_617);
or U462 (N_462,In_1044,In_952);
or U463 (N_463,In_1983,In_311);
xor U464 (N_464,In_576,In_1525);
nand U465 (N_465,In_703,In_1358);
or U466 (N_466,In_633,In_1074);
nand U467 (N_467,In_584,In_951);
nand U468 (N_468,In_700,In_970);
xnor U469 (N_469,In_546,In_1040);
and U470 (N_470,In_349,In_911);
nand U471 (N_471,In_1390,In_209);
nand U472 (N_472,In_111,In_1593);
nand U473 (N_473,In_1821,In_42);
or U474 (N_474,In_1820,In_149);
or U475 (N_475,In_489,In_1475);
nand U476 (N_476,In_1562,In_1474);
nor U477 (N_477,In_324,In_702);
xnor U478 (N_478,In_655,In_1994);
nor U479 (N_479,In_278,In_854);
or U480 (N_480,In_1495,In_1664);
or U481 (N_481,In_1850,In_1689);
xor U482 (N_482,In_337,In_664);
xor U483 (N_483,In_1745,In_1957);
and U484 (N_484,In_1175,In_126);
and U485 (N_485,In_221,In_1046);
nand U486 (N_486,In_1423,In_824);
nand U487 (N_487,In_1213,In_1824);
nor U488 (N_488,In_28,In_1632);
or U489 (N_489,In_1681,In_1706);
xnor U490 (N_490,In_754,In_929);
xor U491 (N_491,In_966,In_790);
and U492 (N_492,In_935,In_1990);
xnor U493 (N_493,In_316,In_1703);
and U494 (N_494,In_419,In_816);
xnor U495 (N_495,In_1067,In_1208);
or U496 (N_496,In_901,In_1065);
nor U497 (N_497,In_1438,In_913);
and U498 (N_498,In_1238,In_1559);
or U499 (N_499,In_68,In_800);
nand U500 (N_500,In_1153,In_659);
nor U501 (N_501,In_704,In_1926);
and U502 (N_502,In_52,In_1424);
and U503 (N_503,In_765,In_1928);
nand U504 (N_504,In_130,In_216);
nor U505 (N_505,In_82,In_727);
or U506 (N_506,In_1123,In_280);
or U507 (N_507,In_129,In_201);
or U508 (N_508,In_958,In_532);
nor U509 (N_509,In_425,In_820);
nand U510 (N_510,In_92,In_1761);
and U511 (N_511,In_1939,In_325);
nor U512 (N_512,In_543,In_1512);
xor U513 (N_513,In_1506,In_331);
nand U514 (N_514,In_1959,In_1374);
xnor U515 (N_515,In_620,In_222);
nand U516 (N_516,In_1236,In_299);
or U517 (N_517,In_1613,In_1226);
or U518 (N_518,In_1252,In_1145);
nand U519 (N_519,In_745,In_1240);
or U520 (N_520,In_1875,In_1823);
or U521 (N_521,In_962,In_1975);
nand U522 (N_522,In_1918,In_1497);
nand U523 (N_523,In_1079,In_779);
and U524 (N_524,In_394,In_738);
nor U525 (N_525,In_1366,In_491);
nand U526 (N_526,In_1925,In_205);
nor U527 (N_527,In_1154,In_341);
nand U528 (N_528,In_1075,In_1290);
nand U529 (N_529,In_494,In_1413);
or U530 (N_530,In_1866,In_204);
xnor U531 (N_531,In_307,In_1185);
and U532 (N_532,In_67,In_1986);
xnor U533 (N_533,In_1877,In_1680);
or U534 (N_534,In_1665,In_1568);
xor U535 (N_535,In_435,In_636);
nand U536 (N_536,In_1595,In_1818);
or U537 (N_537,In_1483,In_1477);
nor U538 (N_538,In_30,In_1288);
nand U539 (N_539,In_57,In_1372);
nand U540 (N_540,In_609,In_1692);
xnor U541 (N_541,In_1979,In_1463);
and U542 (N_542,In_559,In_1194);
or U543 (N_543,In_1574,In_1206);
nand U544 (N_544,In_1653,In_16);
nand U545 (N_545,In_1751,In_251);
xnor U546 (N_546,In_376,In_558);
and U547 (N_547,In_1518,In_23);
nor U548 (N_548,In_448,In_1576);
or U549 (N_549,In_529,In_1071);
nand U550 (N_550,In_1504,In_1878);
nand U551 (N_551,In_1328,In_1127);
nand U552 (N_552,In_846,In_1598);
nor U553 (N_553,In_1623,In_148);
xor U554 (N_554,In_35,In_1004);
nor U555 (N_555,In_859,In_791);
xor U556 (N_556,In_1539,In_276);
nor U557 (N_557,In_464,In_1513);
xor U558 (N_558,In_284,In_384);
xor U559 (N_559,In_1651,In_463);
nand U560 (N_560,In_1480,In_718);
nor U561 (N_561,In_194,In_228);
nor U562 (N_562,In_1848,In_1500);
nor U563 (N_563,In_1443,In_407);
or U564 (N_564,In_1266,In_533);
xor U565 (N_565,In_1940,In_404);
or U566 (N_566,In_581,In_1246);
nand U567 (N_567,In_1813,In_1775);
nand U568 (N_568,In_1333,In_121);
nand U569 (N_569,In_1169,In_203);
or U570 (N_570,In_1882,In_500);
and U571 (N_571,In_894,In_488);
nor U572 (N_572,In_593,In_1749);
nor U573 (N_573,In_418,In_947);
xnor U574 (N_574,In_363,In_240);
xor U575 (N_575,In_1889,In_1712);
xnor U576 (N_576,In_1816,In_226);
nor U577 (N_577,In_1430,In_54);
xor U578 (N_578,In_1802,In_1146);
or U579 (N_579,In_182,In_432);
xor U580 (N_580,In_510,In_989);
or U581 (N_581,In_638,In_777);
or U582 (N_582,In_1104,In_11);
nand U583 (N_583,In_1050,In_766);
and U584 (N_584,In_729,In_444);
nand U585 (N_585,In_1432,In_265);
and U586 (N_586,In_426,In_591);
or U587 (N_587,In_809,In_1520);
nand U588 (N_588,In_1634,In_1885);
or U589 (N_589,In_1984,In_588);
nor U590 (N_590,In_968,In_224);
xor U591 (N_591,In_1391,In_1296);
nor U592 (N_592,In_698,In_243);
or U593 (N_593,In_271,In_1011);
nor U594 (N_594,In_225,In_37);
nor U595 (N_595,In_1700,In_487);
nor U596 (N_596,In_10,In_1399);
nor U597 (N_597,In_1566,In_1943);
xor U598 (N_598,In_1405,In_810);
and U599 (N_599,In_774,In_1501);
and U600 (N_600,In_128,In_322);
nor U601 (N_601,In_210,In_1098);
or U602 (N_602,In_1479,In_1081);
nand U603 (N_603,In_382,In_275);
or U604 (N_604,In_219,In_725);
nor U605 (N_605,In_1384,In_516);
and U606 (N_606,In_1454,In_921);
nand U607 (N_607,In_1717,In_1884);
and U608 (N_608,In_678,In_70);
or U609 (N_609,In_365,In_1089);
nand U610 (N_610,In_468,In_437);
nor U611 (N_611,In_1178,In_1895);
nand U612 (N_612,In_85,In_1523);
nand U613 (N_613,In_953,In_1766);
nor U614 (N_614,In_575,In_560);
xnor U615 (N_615,In_1010,In_1445);
and U616 (N_616,In_879,In_1211);
nand U617 (N_617,In_244,In_1198);
nand U618 (N_618,In_1130,In_1033);
xnor U619 (N_619,In_361,In_1550);
and U620 (N_620,In_1163,In_495);
or U621 (N_621,In_694,In_351);
nand U622 (N_622,In_1224,In_181);
xor U623 (N_623,In_925,In_782);
and U624 (N_624,In_423,In_1400);
or U625 (N_625,In_1190,In_323);
xor U626 (N_626,In_1516,In_590);
nand U627 (N_627,In_1070,In_107);
or U628 (N_628,In_669,In_839);
nor U629 (N_629,In_1591,In_1170);
nor U630 (N_630,In_1077,In_409);
and U631 (N_631,In_1526,In_259);
xnor U632 (N_632,In_1861,In_381);
and U633 (N_633,In_1835,In_1599);
or U634 (N_634,In_604,In_526);
and U635 (N_635,In_764,In_949);
or U636 (N_636,In_279,In_1060);
nand U637 (N_637,In_1227,In_568);
xnor U638 (N_638,In_1028,In_261);
nor U639 (N_639,In_1771,In_1193);
nand U640 (N_640,In_1620,In_1893);
or U641 (N_641,In_1795,In_1307);
xor U642 (N_642,In_1757,In_1429);
nor U643 (N_643,In_1128,In_508);
nor U644 (N_644,In_24,In_1285);
xor U645 (N_645,In_1453,In_39);
nor U646 (N_646,In_386,In_1528);
nor U647 (N_647,In_393,In_144);
nand U648 (N_648,In_1197,In_997);
xnor U649 (N_649,In_651,In_100);
nand U650 (N_650,In_1542,In_542);
or U651 (N_651,In_1843,In_245);
or U652 (N_652,In_60,In_78);
nor U653 (N_653,In_1798,In_1034);
or U654 (N_654,In_12,In_260);
and U655 (N_655,In_1476,In_1865);
or U656 (N_656,In_1455,In_1232);
nor U657 (N_657,In_1499,In_883);
and U658 (N_658,In_788,In_1790);
xor U659 (N_659,In_1747,In_1711);
xnor U660 (N_660,In_1187,In_1715);
xor U661 (N_661,In_715,In_1337);
nand U662 (N_662,In_1774,In_414);
xnor U663 (N_663,In_668,In_1707);
or U664 (N_664,In_1395,In_1294);
nor U665 (N_665,In_522,In_881);
and U666 (N_666,In_1039,In_257);
or U667 (N_667,In_688,In_1997);
xnor U668 (N_668,In_344,In_767);
xnor U669 (N_669,In_1038,In_452);
nand U670 (N_670,In_619,In_1762);
xor U671 (N_671,In_1966,In_466);
or U672 (N_672,In_239,In_959);
xnor U673 (N_673,In_1950,In_827);
or U674 (N_674,In_1541,In_1021);
nor U675 (N_675,In_691,In_1314);
or U676 (N_676,In_1176,In_1135);
and U677 (N_677,In_438,In_914);
xnor U678 (N_678,In_939,In_1363);
or U679 (N_679,In_445,In_1);
and U680 (N_680,In_1045,In_320);
or U681 (N_681,In_1812,In_1467);
nand U682 (N_682,In_871,In_868);
and U683 (N_683,In_1383,In_547);
nor U684 (N_684,In_753,In_945);
xor U685 (N_685,In_983,In_1403);
xor U686 (N_686,In_1815,In_631);
xnor U687 (N_687,In_794,In_94);
nand U688 (N_688,In_1674,In_1385);
nand U689 (N_689,In_1379,In_1376);
xor U690 (N_690,In_1794,In_416);
xnor U691 (N_691,In_1627,In_1249);
xnor U692 (N_692,In_884,In_1735);
or U693 (N_693,In_826,In_1245);
xnor U694 (N_694,In_397,In_898);
or U695 (N_695,In_1167,In_1661);
xnor U696 (N_696,In_1887,In_644);
or U697 (N_697,In_422,In_942);
and U698 (N_698,In_1073,In_1426);
nand U699 (N_699,In_1838,In_1544);
xor U700 (N_700,In_313,In_866);
nor U701 (N_701,In_1727,In_1247);
xnor U702 (N_702,In_847,In_944);
xnor U703 (N_703,In_1732,In_906);
nor U704 (N_704,In_1179,In_1007);
nand U705 (N_705,In_188,In_1831);
nand U706 (N_706,In_1367,In_1428);
nor U707 (N_707,In_1026,In_1008);
or U708 (N_708,In_305,In_960);
and U709 (N_709,In_1788,In_642);
xnor U710 (N_710,In_321,In_1551);
and U711 (N_711,In_1078,In_1894);
or U712 (N_712,In_1600,In_1239);
nor U713 (N_713,In_923,In_1377);
xnor U714 (N_714,In_1182,In_83);
nor U715 (N_715,In_1292,In_1255);
xnor U716 (N_716,In_1279,In_737);
or U717 (N_717,In_112,In_142);
nor U718 (N_718,In_1649,In_1451);
nand U719 (N_719,In_1638,In_889);
or U720 (N_720,In_1289,In_291);
or U721 (N_721,In_650,In_1936);
xor U722 (N_722,In_1014,In_408);
nand U723 (N_723,In_886,In_972);
and U724 (N_724,In_1856,In_1470);
nor U725 (N_725,In_333,In_1886);
xor U726 (N_726,In_685,In_562);
and U727 (N_727,In_772,In_1896);
nor U728 (N_728,In_298,In_1387);
or U729 (N_729,In_483,In_676);
xnor U730 (N_730,In_1388,In_1834);
xnor U731 (N_731,In_1842,In_1605);
nand U732 (N_732,In_917,In_661);
or U733 (N_733,In_803,In_1096);
xnor U734 (N_734,In_1375,In_1286);
xnor U735 (N_735,In_1777,In_1931);
xor U736 (N_736,In_963,In_1106);
or U737 (N_737,In_1053,In_1579);
xor U738 (N_738,In_1829,In_869);
and U739 (N_739,In_1505,In_999);
xnor U740 (N_740,In_728,In_246);
nand U741 (N_741,In_998,In_1952);
and U742 (N_742,In_1993,In_1955);
nor U743 (N_743,In_530,In_335);
or U744 (N_744,In_1679,In_646);
nor U745 (N_745,In_733,In_1341);
and U746 (N_746,In_978,In_84);
or U747 (N_747,In_648,In_837);
or U748 (N_748,In_1254,In_554);
nor U749 (N_749,In_1899,In_1219);
nand U750 (N_750,In_1440,In_880);
and U751 (N_751,In_190,In_1415);
nor U752 (N_752,In_1604,In_890);
nor U753 (N_753,In_1782,In_15);
nor U754 (N_754,In_283,In_1776);
nand U755 (N_755,In_940,In_1189);
nor U756 (N_756,In_589,In_658);
xnor U757 (N_757,In_509,In_199);
nor U758 (N_758,In_29,In_1626);
and U759 (N_759,In_1575,In_231);
nand U760 (N_760,In_1911,In_48);
nor U761 (N_761,In_162,In_1209);
nand U762 (N_762,In_1433,In_110);
or U763 (N_763,In_101,In_417);
nor U764 (N_764,In_540,In_348);
nand U765 (N_765,In_673,In_1909);
xnor U766 (N_766,In_1555,In_1001);
xor U767 (N_767,In_730,In_146);
or U768 (N_768,In_851,In_1890);
nand U769 (N_769,In_1017,In_501);
nor U770 (N_770,In_723,In_330);
or U771 (N_771,In_950,In_512);
nand U772 (N_772,In_1571,In_674);
nor U773 (N_773,In_986,In_1808);
xor U774 (N_774,In_304,In_1536);
or U775 (N_775,In_2,In_1583);
and U776 (N_776,In_98,In_1678);
or U777 (N_777,In_1572,In_716);
or U778 (N_778,In_1779,In_1954);
and U779 (N_779,In_552,In_1772);
xor U780 (N_780,In_1441,In_701);
xor U781 (N_781,In_1137,In_654);
xor U782 (N_782,In_1354,In_797);
nand U783 (N_783,In_1709,In_328);
nor U784 (N_784,In_623,In_268);
nor U785 (N_785,In_1683,In_1062);
or U786 (N_786,In_740,In_1673);
nor U787 (N_787,In_1636,In_1609);
xnor U788 (N_788,In_804,In_96);
and U789 (N_789,In_1531,In_672);
or U790 (N_790,In_165,In_1407);
or U791 (N_791,In_4,In_656);
or U792 (N_792,In_786,In_1654);
nor U793 (N_793,In_22,In_1549);
or U794 (N_794,In_213,In_875);
nor U795 (N_795,In_1295,In_1051);
and U796 (N_796,In_296,In_166);
nor U797 (N_797,In_1630,In_519);
nand U798 (N_798,In_1117,In_574);
nand U799 (N_799,In_768,In_1482);
or U800 (N_800,In_1671,In_1473);
nor U801 (N_801,In_1973,In_1977);
xor U802 (N_802,In_599,In_1511);
nor U803 (N_803,In_583,In_93);
and U804 (N_804,In_504,In_1256);
xnor U805 (N_805,In_1942,In_65);
nand U806 (N_806,In_1215,In_625);
nor U807 (N_807,In_20,In_1967);
xor U808 (N_808,In_506,In_1022);
or U809 (N_809,In_587,In_1833);
and U810 (N_810,In_1529,In_43);
or U811 (N_811,In_815,In_1323);
and U812 (N_812,In_1569,In_937);
nand U813 (N_813,In_1257,In_1941);
xor U814 (N_814,In_139,In_757);
or U815 (N_815,In_343,In_909);
or U816 (N_816,In_1402,In_1922);
nor U817 (N_817,In_1301,In_1892);
xor U818 (N_818,In_1346,In_63);
and U819 (N_819,In_447,In_956);
nor U820 (N_820,In_1656,In_1867);
and U821 (N_821,In_1946,In_818);
and U822 (N_822,In_1696,In_1858);
xnor U823 (N_823,In_1982,In_758);
xor U824 (N_824,In_1494,In_1543);
xor U825 (N_825,In_1767,In_176);
and U826 (N_826,In_1621,In_95);
nand U827 (N_827,In_1710,In_1260);
nand U828 (N_828,In_545,In_287);
nor U829 (N_829,In_1436,In_1490);
or U830 (N_830,In_1781,In_1210);
nand U831 (N_831,In_1590,In_988);
and U832 (N_832,In_1158,In_1640);
nor U833 (N_833,In_1901,In_1725);
or U834 (N_834,In_1364,In_852);
nand U835 (N_835,In_1355,In_1724);
nor U836 (N_836,In_1343,In_1981);
and U837 (N_837,In_641,In_1789);
and U838 (N_838,In_1177,In_1978);
xor U839 (N_839,In_1338,In_1611);
nor U840 (N_840,In_152,In_1009);
or U841 (N_841,In_0,In_1729);
and U842 (N_842,In_1468,In_1069);
nor U843 (N_843,In_1854,In_1241);
nor U844 (N_844,In_178,In_513);
and U845 (N_845,In_527,In_555);
nand U846 (N_846,In_87,In_908);
nor U847 (N_847,In_391,In_440);
and U848 (N_848,In_1748,In_170);
or U849 (N_849,In_1561,In_887);
nand U850 (N_850,In_1919,In_450);
nand U851 (N_851,In_515,In_1597);
and U852 (N_852,In_900,In_1270);
nor U853 (N_853,In_1722,In_1646);
nand U854 (N_854,In_59,In_1305);
nor U855 (N_855,In_79,In_303);
nor U856 (N_856,In_1125,In_1675);
xor U857 (N_857,In_971,In_308);
or U858 (N_858,In_332,In_910);
nor U859 (N_859,In_362,In_825);
nand U860 (N_860,In_1103,In_1974);
nor U861 (N_861,In_1284,In_1805);
nor U862 (N_862,In_751,In_585);
and U863 (N_863,In_1370,In_373);
xnor U864 (N_864,In_1560,In_1934);
nor U865 (N_865,In_1765,In_1068);
and U866 (N_866,In_860,In_806);
or U867 (N_867,In_1869,In_1264);
xor U868 (N_868,In_1985,In_1086);
nand U869 (N_869,In_596,In_1108);
nor U870 (N_870,In_1460,In_667);
nor U871 (N_871,In_342,In_172);
or U872 (N_872,In_5,In_607);
nand U873 (N_873,In_870,In_274);
or U874 (N_874,In_211,In_427);
xor U875 (N_875,In_1662,In_1231);
and U876 (N_876,In_1452,In_521);
or U877 (N_877,In_1417,In_1447);
or U878 (N_878,In_1134,In_1914);
xnor U879 (N_879,In_61,In_1274);
nand U880 (N_880,In_1336,In_1924);
xnor U881 (N_881,In_1097,In_1780);
nor U882 (N_882,In_1507,In_1635);
xnor U883 (N_883,In_882,In_1738);
xnor U884 (N_884,In_1846,In_1809);
xnor U885 (N_885,In_90,In_872);
or U886 (N_886,In_329,In_1275);
xnor U887 (N_887,In_86,In_133);
nand U888 (N_888,In_621,In_1350);
nor U889 (N_889,In_1431,In_1916);
and U890 (N_890,In_1521,In_1508);
or U891 (N_891,In_1041,In_1608);
and U892 (N_892,In_578,In_493);
nand U893 (N_893,In_1874,In_233);
nor U894 (N_894,In_1088,In_1277);
nand U895 (N_895,In_140,In_666);
nand U896 (N_896,In_735,In_979);
nand U897 (N_897,In_1030,In_982);
nor U898 (N_898,In_686,In_1530);
nor U899 (N_899,In_897,In_364);
nor U900 (N_900,In_602,In_38);
or U901 (N_901,In_369,In_1847);
and U902 (N_902,In_1515,In_1272);
nand U903 (N_903,In_286,In_1691);
xnor U904 (N_904,In_485,In_294);
xnor U905 (N_905,In_1061,In_1637);
xor U906 (N_906,In_1036,In_1250);
xnor U907 (N_907,In_411,In_1612);
and U908 (N_908,In_367,In_1330);
nor U909 (N_909,In_1101,In_1406);
nor U910 (N_910,In_1485,In_964);
xor U911 (N_911,In_301,In_187);
and U912 (N_912,In_1554,In_750);
xor U913 (N_913,In_395,In_220);
or U914 (N_914,In_731,In_1750);
xor U915 (N_915,In_197,In_557);
and U916 (N_916,In_1442,In_1953);
or U917 (N_917,In_143,In_1291);
nand U918 (N_918,In_158,In_1359);
or U919 (N_919,In_1616,In_1434);
or U920 (N_920,In_1469,In_141);
nor U921 (N_921,In_967,In_497);
nand U922 (N_922,In_973,In_1814);
or U923 (N_923,In_1351,In_1269);
or U924 (N_924,In_1910,In_649);
xnor U925 (N_925,In_264,In_1085);
nor U926 (N_926,In_831,In_981);
xor U927 (N_927,In_191,In_1409);
nor U928 (N_928,In_467,In_520);
nor U929 (N_929,In_1139,In_71);
and U930 (N_930,In_1796,In_1923);
nand U931 (N_931,In_1332,In_1667);
xor U932 (N_932,In_1694,In_453);
and U933 (N_933,In_1792,In_1107);
or U934 (N_934,In_862,In_932);
and U935 (N_935,In_237,In_1339);
xor U936 (N_936,In_1672,In_732);
or U937 (N_937,In_1414,In_996);
or U938 (N_938,In_1138,In_787);
nor U939 (N_939,In_548,In_830);
and U940 (N_940,In_840,In_179);
nor U941 (N_941,In_1999,In_1971);
nor U942 (N_942,In_1084,In_62);
and U943 (N_943,In_1996,In_1567);
xor U944 (N_944,In_1938,In_1316);
nand U945 (N_945,In_103,In_920);
and U946 (N_946,In_1322,In_943);
xnor U947 (N_947,In_1013,In_1596);
nand U948 (N_948,In_507,In_1491);
or U949 (N_949,In_449,In_473);
and U950 (N_950,In_1760,In_1042);
nand U951 (N_951,In_319,In_1524);
xnor U952 (N_952,In_1647,In_253);
or U953 (N_953,In_1944,In_1329);
xor U954 (N_954,In_1251,In_183);
and U955 (N_955,In_272,In_612);
and U956 (N_956,In_412,In_1090);
xnor U957 (N_957,In_1756,In_1763);
or U958 (N_958,In_1628,In_457);
nor U959 (N_959,In_1849,In_1639);
and U960 (N_960,In_420,In_833);
nor U961 (N_961,In_1840,In_1883);
and U962 (N_962,In_1670,In_1212);
xor U963 (N_963,In_1830,In_961);
xor U964 (N_964,In_1458,In_1592);
or U965 (N_965,In_1859,In_1110);
nand U966 (N_966,In_736,In_1708);
nand U967 (N_967,In_1935,In_689);
nor U968 (N_968,In_1133,In_1144);
or U969 (N_969,In_1970,In_1118);
and U970 (N_970,In_206,In_18);
and U971 (N_971,In_1688,In_1871);
nand U972 (N_972,In_874,In_1644);
xor U973 (N_973,In_1655,In_813);
nand U974 (N_974,In_776,In_785);
xnor U975 (N_975,In_780,In_1087);
nand U976 (N_976,In_1221,In_51);
and U977 (N_977,In_370,In_969);
nand U978 (N_978,In_1188,In_470);
xnor U979 (N_979,In_721,In_525);
xor U980 (N_980,In_1741,In_1161);
and U981 (N_981,In_123,In_1903);
nor U982 (N_982,In_1514,In_1589);
xnor U983 (N_983,In_288,In_744);
nand U984 (N_984,In_1072,In_410);
xor U985 (N_985,In_1960,In_403);
and U986 (N_986,In_1912,In_850);
nor U987 (N_987,In_511,In_1517);
and U988 (N_988,In_867,In_1412);
and U989 (N_989,In_1319,In_1905);
nand U990 (N_990,In_1165,In_115);
xor U991 (N_991,In_936,In_73);
xnor U992 (N_992,In_769,In_618);
nor U993 (N_993,In_247,In_1719);
and U994 (N_994,In_281,In_1312);
or U995 (N_995,In_124,In_1481);
and U996 (N_996,In_122,In_1235);
or U997 (N_997,In_1863,In_1726);
and U998 (N_998,In_637,In_567);
or U999 (N_999,In_1151,In_1047);
xnor U1000 (N_1000,N_507,N_635);
and U1001 (N_1001,N_618,N_363);
nor U1002 (N_1002,N_842,N_819);
nor U1003 (N_1003,N_807,N_371);
xnor U1004 (N_1004,N_833,N_440);
nor U1005 (N_1005,N_595,N_718);
or U1006 (N_1006,N_285,N_661);
nand U1007 (N_1007,N_428,N_152);
nand U1008 (N_1008,N_412,N_598);
or U1009 (N_1009,N_441,N_492);
nand U1010 (N_1010,N_360,N_865);
and U1011 (N_1011,N_17,N_419);
nand U1012 (N_1012,N_940,N_714);
nor U1013 (N_1013,N_463,N_373);
nand U1014 (N_1014,N_794,N_395);
and U1015 (N_1015,N_651,N_534);
nor U1016 (N_1016,N_830,N_526);
nand U1017 (N_1017,N_500,N_973);
or U1018 (N_1018,N_906,N_14);
nand U1019 (N_1019,N_383,N_646);
nand U1020 (N_1020,N_495,N_780);
xnor U1021 (N_1021,N_978,N_509);
nor U1022 (N_1022,N_279,N_685);
or U1023 (N_1023,N_958,N_53);
xor U1024 (N_1024,N_854,N_118);
or U1025 (N_1025,N_359,N_109);
nor U1026 (N_1026,N_178,N_80);
nor U1027 (N_1027,N_394,N_270);
nor U1028 (N_1028,N_572,N_736);
xnor U1029 (N_1029,N_739,N_448);
nor U1030 (N_1030,N_757,N_265);
and U1031 (N_1031,N_792,N_560);
nor U1032 (N_1032,N_793,N_212);
and U1033 (N_1033,N_782,N_147);
xor U1034 (N_1034,N_485,N_219);
nand U1035 (N_1035,N_514,N_486);
and U1036 (N_1036,N_131,N_103);
or U1037 (N_1037,N_624,N_436);
xnor U1038 (N_1038,N_471,N_79);
xor U1039 (N_1039,N_340,N_781);
nand U1040 (N_1040,N_205,N_915);
or U1041 (N_1041,N_771,N_497);
and U1042 (N_1042,N_576,N_614);
xor U1043 (N_1043,N_700,N_216);
or U1044 (N_1044,N_465,N_803);
or U1045 (N_1045,N_133,N_424);
and U1046 (N_1046,N_893,N_350);
nor U1047 (N_1047,N_992,N_63);
nand U1048 (N_1048,N_808,N_970);
xor U1049 (N_1049,N_54,N_923);
nor U1050 (N_1050,N_105,N_564);
nor U1051 (N_1051,N_837,N_774);
xnor U1052 (N_1052,N_400,N_40);
or U1053 (N_1053,N_449,N_277);
or U1054 (N_1054,N_149,N_554);
or U1055 (N_1055,N_206,N_670);
and U1056 (N_1056,N_910,N_20);
and U1057 (N_1057,N_330,N_888);
or U1058 (N_1058,N_242,N_537);
and U1059 (N_1059,N_733,N_744);
nor U1060 (N_1060,N_225,N_846);
or U1061 (N_1061,N_316,N_622);
nand U1062 (N_1062,N_114,N_708);
or U1063 (N_1063,N_121,N_73);
xor U1064 (N_1064,N_386,N_252);
nand U1065 (N_1065,N_664,N_88);
nand U1066 (N_1066,N_106,N_167);
and U1067 (N_1067,N_288,N_155);
nor U1068 (N_1068,N_107,N_305);
nand U1069 (N_1069,N_989,N_160);
and U1070 (N_1070,N_601,N_937);
and U1071 (N_1071,N_84,N_203);
nand U1072 (N_1072,N_318,N_422);
nor U1073 (N_1073,N_697,N_38);
nand U1074 (N_1074,N_444,N_66);
nand U1075 (N_1075,N_229,N_578);
and U1076 (N_1076,N_932,N_291);
or U1077 (N_1077,N_62,N_328);
xor U1078 (N_1078,N_2,N_934);
nand U1079 (N_1079,N_476,N_481);
and U1080 (N_1080,N_358,N_821);
nand U1081 (N_1081,N_672,N_317);
or U1082 (N_1082,N_899,N_687);
or U1083 (N_1083,N_593,N_690);
nor U1084 (N_1084,N_337,N_67);
nand U1085 (N_1085,N_692,N_789);
nor U1086 (N_1086,N_90,N_549);
nor U1087 (N_1087,N_579,N_35);
and U1088 (N_1088,N_420,N_489);
nand U1089 (N_1089,N_283,N_797);
nand U1090 (N_1090,N_312,N_272);
nor U1091 (N_1091,N_136,N_166);
or U1092 (N_1092,N_679,N_768);
nor U1093 (N_1093,N_10,N_960);
or U1094 (N_1094,N_408,N_749);
nor U1095 (N_1095,N_409,N_348);
xnor U1096 (N_1096,N_309,N_108);
nand U1097 (N_1097,N_196,N_342);
and U1098 (N_1098,N_384,N_37);
and U1099 (N_1099,N_880,N_853);
nand U1100 (N_1100,N_901,N_947);
nor U1101 (N_1101,N_473,N_969);
xor U1102 (N_1102,N_477,N_620);
nand U1103 (N_1103,N_49,N_946);
nand U1104 (N_1104,N_873,N_369);
nor U1105 (N_1105,N_584,N_563);
and U1106 (N_1106,N_141,N_851);
nor U1107 (N_1107,N_843,N_723);
nand U1108 (N_1108,N_625,N_680);
nand U1109 (N_1109,N_674,N_326);
xor U1110 (N_1110,N_998,N_126);
or U1111 (N_1111,N_621,N_34);
xor U1112 (N_1112,N_382,N_539);
and U1113 (N_1113,N_188,N_902);
nand U1114 (N_1114,N_855,N_538);
and U1115 (N_1115,N_832,N_182);
nor U1116 (N_1116,N_331,N_30);
or U1117 (N_1117,N_675,N_11);
nor U1118 (N_1118,N_688,N_453);
nor U1119 (N_1119,N_5,N_335);
and U1120 (N_1120,N_239,N_811);
nand U1121 (N_1121,N_245,N_938);
xor U1122 (N_1122,N_24,N_531);
and U1123 (N_1123,N_478,N_323);
or U1124 (N_1124,N_208,N_266);
nor U1125 (N_1125,N_986,N_78);
xnor U1126 (N_1126,N_597,N_583);
nor U1127 (N_1127,N_365,N_804);
and U1128 (N_1128,N_438,N_591);
nor U1129 (N_1129,N_284,N_268);
or U1130 (N_1130,N_362,N_437);
or U1131 (N_1131,N_499,N_559);
xor U1132 (N_1132,N_740,N_553);
and U1133 (N_1133,N_988,N_712);
or U1134 (N_1134,N_728,N_370);
or U1135 (N_1135,N_380,N_673);
nand U1136 (N_1136,N_791,N_926);
nor U1137 (N_1137,N_528,N_931);
and U1138 (N_1138,N_308,N_629);
xor U1139 (N_1139,N_462,N_496);
nor U1140 (N_1140,N_310,N_171);
and U1141 (N_1141,N_678,N_849);
nand U1142 (N_1142,N_125,N_936);
nor U1143 (N_1143,N_707,N_161);
or U1144 (N_1144,N_968,N_154);
and U1145 (N_1145,N_405,N_329);
nand U1146 (N_1146,N_75,N_456);
xor U1147 (N_1147,N_727,N_975);
or U1148 (N_1148,N_996,N_532);
or U1149 (N_1149,N_493,N_825);
nand U1150 (N_1150,N_388,N_871);
nor U1151 (N_1151,N_480,N_443);
nand U1152 (N_1152,N_530,N_72);
xnor U1153 (N_1153,N_168,N_227);
xor U1154 (N_1154,N_282,N_96);
nor U1155 (N_1155,N_795,N_941);
and U1156 (N_1156,N_375,N_693);
and U1157 (N_1157,N_766,N_710);
nand U1158 (N_1158,N_244,N_983);
xor U1159 (N_1159,N_953,N_985);
and U1160 (N_1160,N_209,N_641);
or U1161 (N_1161,N_724,N_758);
and U1162 (N_1162,N_426,N_957);
xnor U1163 (N_1163,N_25,N_117);
nand U1164 (N_1164,N_741,N_713);
or U1165 (N_1165,N_439,N_210);
xnor U1166 (N_1166,N_101,N_751);
and U1167 (N_1167,N_633,N_355);
nor U1168 (N_1168,N_41,N_615);
or U1169 (N_1169,N_974,N_494);
and U1170 (N_1170,N_349,N_776);
nor U1171 (N_1171,N_129,N_609);
or U1172 (N_1172,N_276,N_286);
and U1173 (N_1173,N_22,N_180);
nor U1174 (N_1174,N_430,N_366);
xnor U1175 (N_1175,N_46,N_55);
nand U1176 (N_1176,N_86,N_100);
xnor U1177 (N_1177,N_702,N_181);
or U1178 (N_1178,N_322,N_427);
nand U1179 (N_1179,N_982,N_224);
or U1180 (N_1180,N_396,N_60);
nand U1181 (N_1181,N_634,N_818);
nand U1182 (N_1182,N_385,N_257);
xor U1183 (N_1183,N_201,N_215);
and U1184 (N_1184,N_952,N_176);
or U1185 (N_1185,N_159,N_99);
xor U1186 (N_1186,N_13,N_955);
xor U1187 (N_1187,N_914,N_85);
xnor U1188 (N_1188,N_194,N_894);
or U1189 (N_1189,N_652,N_660);
nor U1190 (N_1190,N_287,N_655);
nand U1191 (N_1191,N_980,N_746);
xor U1192 (N_1192,N_912,N_729);
nor U1193 (N_1193,N_649,N_413);
nor U1194 (N_1194,N_637,N_338);
xnor U1195 (N_1195,N_944,N_4);
nand U1196 (N_1196,N_616,N_484);
or U1197 (N_1197,N_120,N_258);
xor U1198 (N_1198,N_840,N_725);
xor U1199 (N_1199,N_162,N_423);
nor U1200 (N_1200,N_874,N_518);
and U1201 (N_1201,N_645,N_164);
nor U1202 (N_1202,N_275,N_737);
or U1203 (N_1203,N_567,N_142);
and U1204 (N_1204,N_717,N_232);
nor U1205 (N_1205,N_694,N_157);
or U1206 (N_1206,N_701,N_519);
nand U1207 (N_1207,N_71,N_607);
nand U1208 (N_1208,N_93,N_89);
xnor U1209 (N_1209,N_571,N_483);
or U1210 (N_1210,N_524,N_945);
xor U1211 (N_1211,N_964,N_600);
and U1212 (N_1212,N_608,N_457);
nand U1213 (N_1213,N_632,N_542);
xor U1214 (N_1214,N_754,N_927);
and U1215 (N_1215,N_698,N_346);
xnor U1216 (N_1216,N_234,N_805);
nor U1217 (N_1217,N_70,N_812);
and U1218 (N_1218,N_403,N_472);
nor U1219 (N_1219,N_411,N_623);
nand U1220 (N_1220,N_877,N_876);
nand U1221 (N_1221,N_823,N_433);
nor U1222 (N_1222,N_839,N_200);
xor U1223 (N_1223,N_657,N_418);
xnor U1224 (N_1224,N_399,N_407);
and U1225 (N_1225,N_83,N_255);
nand U1226 (N_1226,N_997,N_510);
nand U1227 (N_1227,N_990,N_44);
nand U1228 (N_1228,N_872,N_414);
nand U1229 (N_1229,N_98,N_568);
and U1230 (N_1230,N_59,N_467);
or U1231 (N_1231,N_521,N_379);
or U1232 (N_1232,N_425,N_321);
or U1233 (N_1233,N_529,N_281);
xnor U1234 (N_1234,N_451,N_26);
nor U1235 (N_1235,N_223,N_7);
or U1236 (N_1236,N_214,N_315);
or U1237 (N_1237,N_847,N_606);
xnor U1238 (N_1238,N_347,N_417);
and U1239 (N_1239,N_897,N_881);
nand U1240 (N_1240,N_202,N_838);
and U1241 (N_1241,N_543,N_230);
or U1242 (N_1242,N_140,N_654);
nand U1243 (N_1243,N_314,N_777);
nor U1244 (N_1244,N_306,N_857);
or U1245 (N_1245,N_274,N_762);
nand U1246 (N_1246,N_236,N_924);
and U1247 (N_1247,N_3,N_195);
or U1248 (N_1248,N_612,N_716);
and U1249 (N_1249,N_332,N_192);
or U1250 (N_1250,N_501,N_94);
or U1251 (N_1251,N_45,N_119);
nor U1252 (N_1252,N_642,N_922);
and U1253 (N_1253,N_844,N_296);
or U1254 (N_1254,N_163,N_662);
and U1255 (N_1255,N_683,N_522);
or U1256 (N_1256,N_689,N_742);
or U1257 (N_1257,N_479,N_199);
and U1258 (N_1258,N_0,N_190);
nand U1259 (N_1259,N_619,N_908);
and U1260 (N_1260,N_515,N_204);
nor U1261 (N_1261,N_432,N_21);
or U1262 (N_1262,N_512,N_351);
nand U1263 (N_1263,N_508,N_545);
nand U1264 (N_1264,N_848,N_822);
xnor U1265 (N_1265,N_574,N_248);
nor U1266 (N_1266,N_594,N_172);
xor U1267 (N_1267,N_339,N_752);
nand U1268 (N_1268,N_237,N_706);
nor U1269 (N_1269,N_994,N_302);
and U1270 (N_1270,N_113,N_130);
and U1271 (N_1271,N_148,N_882);
nor U1272 (N_1272,N_977,N_650);
or U1273 (N_1273,N_639,N_189);
or U1274 (N_1274,N_860,N_617);
or U1275 (N_1275,N_381,N_137);
or U1276 (N_1276,N_150,N_919);
and U1277 (N_1277,N_959,N_801);
or U1278 (N_1278,N_77,N_535);
and U1279 (N_1279,N_592,N_111);
or U1280 (N_1280,N_731,N_124);
and U1281 (N_1281,N_604,N_965);
nand U1282 (N_1282,N_682,N_867);
xnor U1283 (N_1283,N_962,N_565);
nand U1284 (N_1284,N_311,N_590);
and U1285 (N_1285,N_469,N_582);
xor U1286 (N_1286,N_64,N_869);
nor U1287 (N_1287,N_896,N_979);
and U1288 (N_1288,N_533,N_561);
or U1289 (N_1289,N_364,N_341);
xor U1290 (N_1290,N_605,N_246);
and U1291 (N_1291,N_570,N_951);
or U1292 (N_1292,N_65,N_353);
nand U1293 (N_1293,N_884,N_813);
nor U1294 (N_1294,N_42,N_372);
nor U1295 (N_1295,N_112,N_784);
xor U1296 (N_1296,N_56,N_640);
nor U1297 (N_1297,N_581,N_263);
and U1298 (N_1298,N_134,N_628);
nand U1299 (N_1299,N_179,N_905);
and U1300 (N_1300,N_779,N_450);
and U1301 (N_1301,N_841,N_763);
nand U1302 (N_1302,N_862,N_447);
and U1303 (N_1303,N_336,N_82);
xnor U1304 (N_1304,N_186,N_971);
or U1305 (N_1305,N_68,N_861);
or U1306 (N_1306,N_866,N_389);
xor U1307 (N_1307,N_446,N_904);
and U1308 (N_1308,N_156,N_787);
nor U1309 (N_1309,N_343,N_961);
and U1310 (N_1310,N_197,N_415);
and U1311 (N_1311,N_930,N_378);
nor U1312 (N_1312,N_913,N_470);
nor U1313 (N_1313,N_146,N_569);
xnor U1314 (N_1314,N_145,N_292);
nand U1315 (N_1315,N_665,N_631);
nor U1316 (N_1316,N_984,N_987);
nand U1317 (N_1317,N_602,N_153);
or U1318 (N_1318,N_260,N_814);
nor U1319 (N_1319,N_290,N_513);
xnor U1320 (N_1320,N_81,N_231);
or U1321 (N_1321,N_404,N_31);
nor U1322 (N_1322,N_852,N_235);
xor U1323 (N_1323,N_885,N_892);
or U1324 (N_1324,N_19,N_183);
nor U1325 (N_1325,N_921,N_956);
xnor U1326 (N_1326,N_264,N_726);
nand U1327 (N_1327,N_516,N_299);
nand U1328 (N_1328,N_6,N_367);
xnor U1329 (N_1329,N_730,N_254);
nor U1330 (N_1330,N_431,N_523);
nor U1331 (N_1331,N_392,N_177);
nand U1332 (N_1332,N_459,N_517);
nor U1333 (N_1333,N_759,N_834);
nand U1334 (N_1334,N_151,N_278);
xnor U1335 (N_1335,N_74,N_464);
nand U1336 (N_1336,N_525,N_760);
nor U1337 (N_1337,N_806,N_699);
and U1338 (N_1338,N_294,N_596);
or U1339 (N_1339,N_859,N_720);
xor U1340 (N_1340,N_703,N_243);
and U1341 (N_1341,N_251,N_935);
nand U1342 (N_1342,N_18,N_556);
and U1343 (N_1343,N_458,N_920);
nand U1344 (N_1344,N_663,N_589);
xnor U1345 (N_1345,N_966,N_50);
or U1346 (N_1346,N_48,N_52);
nor U1347 (N_1347,N_391,N_57);
xor U1348 (N_1348,N_611,N_256);
xor U1349 (N_1349,N_175,N_490);
xor U1350 (N_1350,N_566,N_240);
nand U1351 (N_1351,N_250,N_249);
and U1352 (N_1352,N_705,N_557);
xor U1353 (N_1353,N_738,N_402);
and U1354 (N_1354,N_221,N_856);
nor U1355 (N_1355,N_262,N_536);
or U1356 (N_1356,N_943,N_273);
nand U1357 (N_1357,N_173,N_442);
and U1358 (N_1358,N_357,N_719);
nand U1359 (N_1359,N_743,N_455);
and U1360 (N_1360,N_586,N_233);
nor U1361 (N_1361,N_750,N_217);
xnor U1362 (N_1362,N_226,N_858);
xor U1363 (N_1363,N_573,N_976);
nand U1364 (N_1364,N_58,N_487);
xnor U1365 (N_1365,N_344,N_220);
nor U1366 (N_1366,N_555,N_69);
xor U1367 (N_1367,N_898,N_61);
nand U1368 (N_1368,N_23,N_993);
xor U1369 (N_1369,N_313,N_127);
and U1370 (N_1370,N_585,N_909);
nand U1371 (N_1371,N_135,N_228);
xnor U1372 (N_1372,N_104,N_753);
xnor U1373 (N_1373,N_636,N_667);
and U1374 (N_1374,N_666,N_110);
nor U1375 (N_1375,N_482,N_184);
nor U1376 (N_1376,N_785,N_304);
xor U1377 (N_1377,N_722,N_735);
xnor U1378 (N_1378,N_454,N_303);
xor U1379 (N_1379,N_376,N_831);
and U1380 (N_1380,N_916,N_721);
nor U1381 (N_1381,N_613,N_755);
nor U1382 (N_1382,N_540,N_47);
nor U1383 (N_1383,N_325,N_732);
nand U1384 (N_1384,N_644,N_16);
or U1385 (N_1385,N_468,N_546);
nand U1386 (N_1386,N_656,N_102);
and U1387 (N_1387,N_116,N_826);
and U1388 (N_1388,N_551,N_51);
nand U1389 (N_1389,N_798,N_879);
nand U1390 (N_1390,N_802,N_778);
and U1391 (N_1391,N_460,N_599);
xnor U1392 (N_1392,N_511,N_928);
nor U1393 (N_1393,N_948,N_580);
nand U1394 (N_1394,N_298,N_28);
and U1395 (N_1395,N_289,N_169);
xnor U1396 (N_1396,N_696,N_132);
xnor U1397 (N_1397,N_261,N_1);
nor U1398 (N_1398,N_747,N_981);
xnor U1399 (N_1399,N_950,N_324);
nor U1400 (N_1400,N_558,N_488);
xnor U1401 (N_1401,N_630,N_800);
nand U1402 (N_1402,N_504,N_648);
nor U1403 (N_1403,N_647,N_668);
and U1404 (N_1404,N_374,N_222);
nand U1405 (N_1405,N_92,N_498);
xor U1406 (N_1406,N_191,N_991);
or U1407 (N_1407,N_253,N_827);
and U1408 (N_1408,N_527,N_815);
and U1409 (N_1409,N_474,N_933);
xor U1410 (N_1410,N_452,N_886);
or U1411 (N_1411,N_506,N_627);
nand U1412 (N_1412,N_783,N_170);
nand U1413 (N_1413,N_850,N_461);
nand U1414 (N_1414,N_29,N_320);
or U1415 (N_1415,N_745,N_875);
nand U1416 (N_1416,N_786,N_128);
and U1417 (N_1417,N_835,N_307);
and U1418 (N_1418,N_368,N_939);
nor U1419 (N_1419,N_491,N_158);
nor U1420 (N_1420,N_87,N_676);
or U1421 (N_1421,N_505,N_241);
or U1422 (N_1422,N_809,N_878);
xor U1423 (N_1423,N_577,N_269);
nor U1424 (N_1424,N_942,N_297);
nand U1425 (N_1425,N_772,N_475);
xor U1426 (N_1426,N_575,N_911);
or U1427 (N_1427,N_756,N_377);
nor U1428 (N_1428,N_387,N_870);
nor U1429 (N_1429,N_691,N_211);
and U1430 (N_1430,N_43,N_445);
or U1431 (N_1431,N_868,N_562);
and U1432 (N_1432,N_709,N_15);
nand U1433 (N_1433,N_820,N_185);
or U1434 (N_1434,N_393,N_686);
nand U1435 (N_1435,N_788,N_972);
xnor U1436 (N_1436,N_548,N_406);
nand U1437 (N_1437,N_677,N_12);
or U1438 (N_1438,N_610,N_900);
and U1439 (N_1439,N_32,N_925);
and U1440 (N_1440,N_97,N_280);
xnor U1441 (N_1441,N_889,N_887);
nor U1442 (N_1442,N_817,N_824);
and U1443 (N_1443,N_999,N_207);
nand U1444 (N_1444,N_36,N_883);
and U1445 (N_1445,N_659,N_300);
nand U1446 (N_1446,N_301,N_587);
nand U1447 (N_1447,N_398,N_434);
nor U1448 (N_1448,N_715,N_401);
nand U1449 (N_1449,N_9,N_907);
and U1450 (N_1450,N_352,N_334);
nor U1451 (N_1451,N_416,N_267);
xnor U1452 (N_1452,N_33,N_995);
nor U1453 (N_1453,N_863,N_681);
and U1454 (N_1454,N_773,N_143);
and U1455 (N_1455,N_198,N_421);
xnor U1456 (N_1456,N_193,N_390);
and U1457 (N_1457,N_333,N_238);
xor U1458 (N_1458,N_76,N_653);
and U1459 (N_1459,N_903,N_658);
or U1460 (N_1460,N_541,N_356);
and U1461 (N_1461,N_917,N_864);
nand U1462 (N_1462,N_704,N_123);
nand U1463 (N_1463,N_345,N_115);
nand U1464 (N_1464,N_547,N_218);
or U1465 (N_1465,N_144,N_929);
xor U1466 (N_1466,N_435,N_796);
nor U1467 (N_1467,N_638,N_165);
xnor U1468 (N_1468,N_765,N_27);
nor U1469 (N_1469,N_354,N_671);
and U1470 (N_1470,N_213,N_799);
xnor U1471 (N_1471,N_410,N_836);
and U1472 (N_1472,N_139,N_247);
and U1473 (N_1473,N_748,N_259);
nor U1474 (N_1474,N_544,N_39);
xnor U1475 (N_1475,N_845,N_466);
and U1476 (N_1476,N_327,N_91);
nand U1477 (N_1477,N_122,N_520);
nor U1478 (N_1478,N_550,N_8);
xnor U1479 (N_1479,N_502,N_95);
and U1480 (N_1480,N_603,N_967);
nor U1481 (N_1481,N_963,N_669);
or U1482 (N_1482,N_626,N_828);
or U1483 (N_1483,N_295,N_138);
nand U1484 (N_1484,N_734,N_174);
nor U1485 (N_1485,N_187,N_895);
and U1486 (N_1486,N_361,N_829);
nor U1487 (N_1487,N_775,N_770);
nand U1488 (N_1488,N_890,N_949);
or U1489 (N_1489,N_397,N_790);
and U1490 (N_1490,N_552,N_695);
and U1491 (N_1491,N_643,N_810);
xor U1492 (N_1492,N_588,N_319);
xor U1493 (N_1493,N_891,N_954);
xnor U1494 (N_1494,N_503,N_761);
nand U1495 (N_1495,N_293,N_764);
nor U1496 (N_1496,N_429,N_684);
and U1497 (N_1497,N_816,N_767);
nor U1498 (N_1498,N_711,N_271);
xnor U1499 (N_1499,N_769,N_918);
nor U1500 (N_1500,N_501,N_434);
nor U1501 (N_1501,N_804,N_471);
xnor U1502 (N_1502,N_663,N_463);
nor U1503 (N_1503,N_394,N_239);
nand U1504 (N_1504,N_444,N_7);
nand U1505 (N_1505,N_182,N_735);
nand U1506 (N_1506,N_283,N_473);
nor U1507 (N_1507,N_893,N_484);
xor U1508 (N_1508,N_838,N_436);
nor U1509 (N_1509,N_76,N_378);
xnor U1510 (N_1510,N_162,N_90);
or U1511 (N_1511,N_891,N_650);
and U1512 (N_1512,N_118,N_965);
nand U1513 (N_1513,N_720,N_916);
or U1514 (N_1514,N_257,N_118);
nand U1515 (N_1515,N_742,N_822);
or U1516 (N_1516,N_330,N_529);
xor U1517 (N_1517,N_82,N_581);
nand U1518 (N_1518,N_505,N_874);
nor U1519 (N_1519,N_714,N_160);
xnor U1520 (N_1520,N_589,N_892);
nand U1521 (N_1521,N_279,N_925);
nand U1522 (N_1522,N_594,N_796);
xor U1523 (N_1523,N_388,N_988);
nor U1524 (N_1524,N_785,N_181);
and U1525 (N_1525,N_293,N_238);
or U1526 (N_1526,N_498,N_168);
nor U1527 (N_1527,N_344,N_832);
nand U1528 (N_1528,N_695,N_538);
and U1529 (N_1529,N_402,N_392);
and U1530 (N_1530,N_77,N_958);
or U1531 (N_1531,N_560,N_173);
xor U1532 (N_1532,N_387,N_6);
nand U1533 (N_1533,N_410,N_591);
xnor U1534 (N_1534,N_35,N_364);
xor U1535 (N_1535,N_841,N_343);
nor U1536 (N_1536,N_237,N_555);
xor U1537 (N_1537,N_230,N_427);
nand U1538 (N_1538,N_615,N_893);
xor U1539 (N_1539,N_268,N_447);
nor U1540 (N_1540,N_923,N_626);
or U1541 (N_1541,N_10,N_828);
and U1542 (N_1542,N_821,N_298);
nand U1543 (N_1543,N_660,N_337);
nand U1544 (N_1544,N_290,N_398);
nor U1545 (N_1545,N_192,N_127);
and U1546 (N_1546,N_14,N_861);
or U1547 (N_1547,N_178,N_378);
xnor U1548 (N_1548,N_670,N_793);
and U1549 (N_1549,N_324,N_177);
nor U1550 (N_1550,N_134,N_525);
and U1551 (N_1551,N_959,N_789);
nor U1552 (N_1552,N_940,N_879);
nand U1553 (N_1553,N_860,N_866);
and U1554 (N_1554,N_375,N_24);
xor U1555 (N_1555,N_745,N_668);
nor U1556 (N_1556,N_777,N_115);
or U1557 (N_1557,N_783,N_430);
and U1558 (N_1558,N_914,N_655);
xor U1559 (N_1559,N_437,N_814);
nor U1560 (N_1560,N_294,N_342);
nand U1561 (N_1561,N_75,N_405);
nor U1562 (N_1562,N_948,N_209);
or U1563 (N_1563,N_272,N_4);
nand U1564 (N_1564,N_369,N_103);
or U1565 (N_1565,N_174,N_237);
xnor U1566 (N_1566,N_827,N_297);
nand U1567 (N_1567,N_964,N_521);
and U1568 (N_1568,N_679,N_288);
or U1569 (N_1569,N_311,N_986);
or U1570 (N_1570,N_682,N_527);
nand U1571 (N_1571,N_272,N_350);
nor U1572 (N_1572,N_821,N_721);
xor U1573 (N_1573,N_477,N_708);
nand U1574 (N_1574,N_606,N_540);
and U1575 (N_1575,N_655,N_248);
nor U1576 (N_1576,N_921,N_658);
and U1577 (N_1577,N_756,N_225);
xnor U1578 (N_1578,N_135,N_914);
nor U1579 (N_1579,N_703,N_326);
nor U1580 (N_1580,N_901,N_116);
or U1581 (N_1581,N_978,N_906);
nor U1582 (N_1582,N_497,N_71);
and U1583 (N_1583,N_661,N_2);
nand U1584 (N_1584,N_762,N_814);
nand U1585 (N_1585,N_621,N_334);
nor U1586 (N_1586,N_443,N_887);
nand U1587 (N_1587,N_428,N_115);
xor U1588 (N_1588,N_787,N_23);
nor U1589 (N_1589,N_897,N_999);
nor U1590 (N_1590,N_818,N_301);
xnor U1591 (N_1591,N_816,N_406);
nand U1592 (N_1592,N_990,N_397);
xnor U1593 (N_1593,N_650,N_383);
xnor U1594 (N_1594,N_606,N_491);
nand U1595 (N_1595,N_951,N_633);
or U1596 (N_1596,N_20,N_837);
nor U1597 (N_1597,N_666,N_637);
nand U1598 (N_1598,N_85,N_278);
or U1599 (N_1599,N_171,N_368);
or U1600 (N_1600,N_113,N_343);
or U1601 (N_1601,N_886,N_621);
or U1602 (N_1602,N_828,N_490);
and U1603 (N_1603,N_428,N_715);
nand U1604 (N_1604,N_171,N_336);
xnor U1605 (N_1605,N_762,N_995);
xnor U1606 (N_1606,N_354,N_83);
nor U1607 (N_1607,N_854,N_271);
xnor U1608 (N_1608,N_917,N_779);
xor U1609 (N_1609,N_278,N_734);
or U1610 (N_1610,N_115,N_565);
nor U1611 (N_1611,N_149,N_662);
nand U1612 (N_1612,N_441,N_155);
and U1613 (N_1613,N_842,N_0);
nor U1614 (N_1614,N_112,N_349);
nand U1615 (N_1615,N_526,N_135);
nand U1616 (N_1616,N_416,N_435);
xor U1617 (N_1617,N_167,N_220);
xor U1618 (N_1618,N_384,N_102);
nor U1619 (N_1619,N_729,N_776);
or U1620 (N_1620,N_194,N_641);
xor U1621 (N_1621,N_120,N_691);
nor U1622 (N_1622,N_497,N_540);
xnor U1623 (N_1623,N_771,N_741);
nand U1624 (N_1624,N_516,N_104);
xor U1625 (N_1625,N_654,N_177);
and U1626 (N_1626,N_843,N_920);
nor U1627 (N_1627,N_199,N_684);
nand U1628 (N_1628,N_769,N_362);
nand U1629 (N_1629,N_757,N_286);
nand U1630 (N_1630,N_505,N_837);
and U1631 (N_1631,N_752,N_855);
nand U1632 (N_1632,N_839,N_435);
nor U1633 (N_1633,N_697,N_513);
and U1634 (N_1634,N_273,N_686);
and U1635 (N_1635,N_652,N_445);
or U1636 (N_1636,N_674,N_480);
nand U1637 (N_1637,N_497,N_451);
and U1638 (N_1638,N_700,N_112);
xnor U1639 (N_1639,N_57,N_938);
or U1640 (N_1640,N_718,N_359);
and U1641 (N_1641,N_577,N_797);
and U1642 (N_1642,N_883,N_216);
nor U1643 (N_1643,N_603,N_359);
and U1644 (N_1644,N_336,N_196);
and U1645 (N_1645,N_854,N_144);
xnor U1646 (N_1646,N_615,N_679);
nand U1647 (N_1647,N_971,N_963);
nand U1648 (N_1648,N_598,N_954);
nor U1649 (N_1649,N_401,N_805);
nand U1650 (N_1650,N_192,N_89);
nand U1651 (N_1651,N_512,N_313);
xor U1652 (N_1652,N_301,N_996);
or U1653 (N_1653,N_423,N_194);
nand U1654 (N_1654,N_436,N_236);
nand U1655 (N_1655,N_891,N_918);
nor U1656 (N_1656,N_494,N_933);
and U1657 (N_1657,N_954,N_166);
xor U1658 (N_1658,N_425,N_27);
and U1659 (N_1659,N_679,N_147);
or U1660 (N_1660,N_188,N_972);
nor U1661 (N_1661,N_877,N_510);
nand U1662 (N_1662,N_547,N_73);
nand U1663 (N_1663,N_986,N_35);
nand U1664 (N_1664,N_742,N_793);
nor U1665 (N_1665,N_221,N_485);
nand U1666 (N_1666,N_658,N_504);
and U1667 (N_1667,N_527,N_669);
nand U1668 (N_1668,N_4,N_76);
or U1669 (N_1669,N_604,N_516);
nand U1670 (N_1670,N_63,N_790);
nor U1671 (N_1671,N_170,N_724);
nor U1672 (N_1672,N_910,N_354);
nor U1673 (N_1673,N_508,N_66);
nor U1674 (N_1674,N_873,N_927);
or U1675 (N_1675,N_678,N_50);
xor U1676 (N_1676,N_94,N_610);
xnor U1677 (N_1677,N_919,N_152);
or U1678 (N_1678,N_415,N_876);
nand U1679 (N_1679,N_762,N_501);
nand U1680 (N_1680,N_717,N_417);
or U1681 (N_1681,N_237,N_633);
nor U1682 (N_1682,N_908,N_762);
and U1683 (N_1683,N_934,N_713);
xnor U1684 (N_1684,N_990,N_266);
or U1685 (N_1685,N_458,N_814);
nor U1686 (N_1686,N_881,N_286);
and U1687 (N_1687,N_27,N_440);
or U1688 (N_1688,N_21,N_542);
nand U1689 (N_1689,N_758,N_930);
nand U1690 (N_1690,N_933,N_546);
nand U1691 (N_1691,N_596,N_410);
and U1692 (N_1692,N_981,N_627);
or U1693 (N_1693,N_786,N_978);
nor U1694 (N_1694,N_1,N_694);
nand U1695 (N_1695,N_876,N_243);
and U1696 (N_1696,N_887,N_982);
or U1697 (N_1697,N_175,N_832);
and U1698 (N_1698,N_318,N_165);
or U1699 (N_1699,N_296,N_775);
or U1700 (N_1700,N_901,N_879);
nor U1701 (N_1701,N_984,N_483);
nor U1702 (N_1702,N_102,N_601);
nor U1703 (N_1703,N_822,N_462);
and U1704 (N_1704,N_372,N_485);
nor U1705 (N_1705,N_547,N_999);
nor U1706 (N_1706,N_304,N_348);
nor U1707 (N_1707,N_45,N_645);
or U1708 (N_1708,N_164,N_166);
nand U1709 (N_1709,N_712,N_974);
nor U1710 (N_1710,N_454,N_775);
xor U1711 (N_1711,N_756,N_920);
or U1712 (N_1712,N_859,N_96);
nand U1713 (N_1713,N_43,N_711);
and U1714 (N_1714,N_195,N_348);
and U1715 (N_1715,N_761,N_547);
nand U1716 (N_1716,N_370,N_685);
or U1717 (N_1717,N_537,N_462);
xor U1718 (N_1718,N_170,N_791);
or U1719 (N_1719,N_452,N_845);
and U1720 (N_1720,N_514,N_917);
xor U1721 (N_1721,N_716,N_583);
nor U1722 (N_1722,N_363,N_25);
or U1723 (N_1723,N_112,N_229);
and U1724 (N_1724,N_425,N_858);
xnor U1725 (N_1725,N_513,N_998);
xor U1726 (N_1726,N_125,N_488);
nand U1727 (N_1727,N_287,N_935);
or U1728 (N_1728,N_873,N_303);
or U1729 (N_1729,N_234,N_933);
and U1730 (N_1730,N_374,N_829);
nand U1731 (N_1731,N_693,N_962);
nand U1732 (N_1732,N_83,N_42);
or U1733 (N_1733,N_757,N_574);
or U1734 (N_1734,N_177,N_671);
nor U1735 (N_1735,N_668,N_265);
or U1736 (N_1736,N_760,N_1);
xnor U1737 (N_1737,N_21,N_596);
nor U1738 (N_1738,N_418,N_532);
or U1739 (N_1739,N_4,N_483);
nor U1740 (N_1740,N_873,N_74);
nor U1741 (N_1741,N_597,N_769);
or U1742 (N_1742,N_966,N_389);
and U1743 (N_1743,N_88,N_315);
and U1744 (N_1744,N_741,N_99);
and U1745 (N_1745,N_250,N_701);
xnor U1746 (N_1746,N_974,N_395);
or U1747 (N_1747,N_950,N_672);
and U1748 (N_1748,N_565,N_304);
nor U1749 (N_1749,N_115,N_845);
nand U1750 (N_1750,N_709,N_375);
nor U1751 (N_1751,N_442,N_373);
nand U1752 (N_1752,N_839,N_472);
or U1753 (N_1753,N_437,N_736);
or U1754 (N_1754,N_255,N_533);
or U1755 (N_1755,N_766,N_248);
xnor U1756 (N_1756,N_771,N_164);
nand U1757 (N_1757,N_356,N_355);
xnor U1758 (N_1758,N_594,N_738);
xnor U1759 (N_1759,N_310,N_940);
or U1760 (N_1760,N_74,N_590);
or U1761 (N_1761,N_776,N_565);
or U1762 (N_1762,N_249,N_706);
and U1763 (N_1763,N_557,N_605);
nor U1764 (N_1764,N_977,N_983);
or U1765 (N_1765,N_810,N_331);
xor U1766 (N_1766,N_587,N_24);
nand U1767 (N_1767,N_944,N_389);
nor U1768 (N_1768,N_647,N_4);
nor U1769 (N_1769,N_394,N_877);
xnor U1770 (N_1770,N_332,N_142);
xnor U1771 (N_1771,N_714,N_759);
nor U1772 (N_1772,N_522,N_606);
nand U1773 (N_1773,N_876,N_993);
xnor U1774 (N_1774,N_453,N_541);
and U1775 (N_1775,N_621,N_447);
nand U1776 (N_1776,N_958,N_33);
nor U1777 (N_1777,N_168,N_596);
nand U1778 (N_1778,N_525,N_848);
or U1779 (N_1779,N_533,N_186);
xor U1780 (N_1780,N_459,N_596);
xnor U1781 (N_1781,N_183,N_928);
or U1782 (N_1782,N_433,N_796);
nor U1783 (N_1783,N_948,N_908);
nand U1784 (N_1784,N_977,N_991);
nor U1785 (N_1785,N_24,N_511);
or U1786 (N_1786,N_507,N_5);
xnor U1787 (N_1787,N_228,N_892);
or U1788 (N_1788,N_98,N_831);
and U1789 (N_1789,N_293,N_833);
nor U1790 (N_1790,N_964,N_199);
xnor U1791 (N_1791,N_593,N_295);
nor U1792 (N_1792,N_298,N_810);
xor U1793 (N_1793,N_219,N_639);
or U1794 (N_1794,N_343,N_28);
nand U1795 (N_1795,N_201,N_759);
and U1796 (N_1796,N_908,N_639);
nor U1797 (N_1797,N_227,N_786);
nand U1798 (N_1798,N_722,N_795);
xor U1799 (N_1799,N_938,N_346);
nor U1800 (N_1800,N_796,N_992);
nor U1801 (N_1801,N_118,N_485);
or U1802 (N_1802,N_930,N_553);
nor U1803 (N_1803,N_752,N_359);
and U1804 (N_1804,N_684,N_782);
nor U1805 (N_1805,N_198,N_29);
or U1806 (N_1806,N_86,N_318);
nand U1807 (N_1807,N_989,N_485);
xor U1808 (N_1808,N_903,N_17);
or U1809 (N_1809,N_780,N_683);
or U1810 (N_1810,N_273,N_975);
or U1811 (N_1811,N_291,N_645);
or U1812 (N_1812,N_759,N_627);
or U1813 (N_1813,N_456,N_915);
or U1814 (N_1814,N_606,N_464);
nand U1815 (N_1815,N_404,N_385);
xor U1816 (N_1816,N_857,N_410);
xor U1817 (N_1817,N_772,N_949);
and U1818 (N_1818,N_665,N_845);
xnor U1819 (N_1819,N_837,N_635);
or U1820 (N_1820,N_927,N_714);
and U1821 (N_1821,N_666,N_355);
nand U1822 (N_1822,N_707,N_631);
or U1823 (N_1823,N_724,N_69);
nor U1824 (N_1824,N_632,N_569);
or U1825 (N_1825,N_846,N_218);
and U1826 (N_1826,N_235,N_72);
xnor U1827 (N_1827,N_111,N_32);
nand U1828 (N_1828,N_498,N_962);
xor U1829 (N_1829,N_845,N_181);
nand U1830 (N_1830,N_385,N_512);
xor U1831 (N_1831,N_829,N_587);
xor U1832 (N_1832,N_427,N_298);
nand U1833 (N_1833,N_553,N_624);
nand U1834 (N_1834,N_497,N_948);
xor U1835 (N_1835,N_596,N_107);
and U1836 (N_1836,N_191,N_101);
nor U1837 (N_1837,N_82,N_365);
or U1838 (N_1838,N_401,N_578);
nor U1839 (N_1839,N_444,N_229);
and U1840 (N_1840,N_66,N_417);
and U1841 (N_1841,N_198,N_972);
or U1842 (N_1842,N_673,N_233);
nand U1843 (N_1843,N_672,N_37);
or U1844 (N_1844,N_169,N_474);
or U1845 (N_1845,N_634,N_726);
nand U1846 (N_1846,N_93,N_18);
and U1847 (N_1847,N_82,N_142);
nor U1848 (N_1848,N_463,N_888);
nand U1849 (N_1849,N_751,N_614);
xnor U1850 (N_1850,N_336,N_874);
xor U1851 (N_1851,N_972,N_660);
xor U1852 (N_1852,N_441,N_569);
nor U1853 (N_1853,N_129,N_840);
and U1854 (N_1854,N_374,N_433);
xnor U1855 (N_1855,N_29,N_739);
or U1856 (N_1856,N_495,N_862);
nand U1857 (N_1857,N_258,N_669);
or U1858 (N_1858,N_192,N_399);
nor U1859 (N_1859,N_181,N_969);
and U1860 (N_1860,N_370,N_613);
nor U1861 (N_1861,N_286,N_209);
and U1862 (N_1862,N_93,N_554);
nor U1863 (N_1863,N_495,N_973);
or U1864 (N_1864,N_515,N_848);
or U1865 (N_1865,N_355,N_990);
or U1866 (N_1866,N_725,N_430);
nand U1867 (N_1867,N_986,N_322);
xor U1868 (N_1868,N_290,N_882);
xor U1869 (N_1869,N_208,N_805);
and U1870 (N_1870,N_196,N_731);
nand U1871 (N_1871,N_939,N_558);
and U1872 (N_1872,N_30,N_102);
and U1873 (N_1873,N_393,N_244);
nand U1874 (N_1874,N_200,N_501);
nor U1875 (N_1875,N_774,N_53);
nor U1876 (N_1876,N_11,N_846);
nor U1877 (N_1877,N_199,N_740);
nand U1878 (N_1878,N_50,N_450);
and U1879 (N_1879,N_624,N_971);
nor U1880 (N_1880,N_5,N_603);
nor U1881 (N_1881,N_346,N_741);
and U1882 (N_1882,N_371,N_2);
nor U1883 (N_1883,N_940,N_291);
and U1884 (N_1884,N_79,N_117);
and U1885 (N_1885,N_755,N_563);
or U1886 (N_1886,N_557,N_628);
and U1887 (N_1887,N_611,N_715);
nand U1888 (N_1888,N_222,N_379);
and U1889 (N_1889,N_396,N_174);
xnor U1890 (N_1890,N_177,N_532);
or U1891 (N_1891,N_976,N_128);
or U1892 (N_1892,N_157,N_979);
and U1893 (N_1893,N_75,N_497);
nand U1894 (N_1894,N_270,N_297);
or U1895 (N_1895,N_264,N_745);
nand U1896 (N_1896,N_462,N_768);
and U1897 (N_1897,N_845,N_401);
and U1898 (N_1898,N_529,N_591);
xnor U1899 (N_1899,N_809,N_629);
nand U1900 (N_1900,N_162,N_554);
xnor U1901 (N_1901,N_647,N_218);
xor U1902 (N_1902,N_804,N_130);
nand U1903 (N_1903,N_402,N_939);
or U1904 (N_1904,N_373,N_601);
or U1905 (N_1905,N_853,N_710);
or U1906 (N_1906,N_285,N_539);
and U1907 (N_1907,N_666,N_335);
and U1908 (N_1908,N_420,N_367);
or U1909 (N_1909,N_705,N_457);
nand U1910 (N_1910,N_676,N_471);
xnor U1911 (N_1911,N_909,N_259);
or U1912 (N_1912,N_492,N_822);
and U1913 (N_1913,N_530,N_837);
xor U1914 (N_1914,N_374,N_620);
nand U1915 (N_1915,N_572,N_694);
xnor U1916 (N_1916,N_763,N_411);
nor U1917 (N_1917,N_954,N_72);
nand U1918 (N_1918,N_426,N_259);
nor U1919 (N_1919,N_416,N_968);
and U1920 (N_1920,N_609,N_605);
or U1921 (N_1921,N_834,N_533);
and U1922 (N_1922,N_918,N_513);
nor U1923 (N_1923,N_933,N_189);
or U1924 (N_1924,N_869,N_204);
xor U1925 (N_1925,N_763,N_309);
and U1926 (N_1926,N_107,N_931);
nand U1927 (N_1927,N_220,N_450);
nand U1928 (N_1928,N_891,N_226);
or U1929 (N_1929,N_922,N_514);
or U1930 (N_1930,N_704,N_827);
nor U1931 (N_1931,N_43,N_414);
nand U1932 (N_1932,N_47,N_842);
nand U1933 (N_1933,N_97,N_672);
and U1934 (N_1934,N_483,N_253);
and U1935 (N_1935,N_153,N_389);
xor U1936 (N_1936,N_178,N_25);
or U1937 (N_1937,N_49,N_187);
and U1938 (N_1938,N_875,N_273);
and U1939 (N_1939,N_801,N_769);
xor U1940 (N_1940,N_927,N_106);
xor U1941 (N_1941,N_670,N_591);
nand U1942 (N_1942,N_571,N_231);
nor U1943 (N_1943,N_262,N_420);
and U1944 (N_1944,N_90,N_590);
nor U1945 (N_1945,N_658,N_49);
and U1946 (N_1946,N_178,N_9);
and U1947 (N_1947,N_662,N_940);
nor U1948 (N_1948,N_928,N_286);
xnor U1949 (N_1949,N_427,N_714);
and U1950 (N_1950,N_459,N_103);
nand U1951 (N_1951,N_758,N_331);
or U1952 (N_1952,N_914,N_139);
nor U1953 (N_1953,N_889,N_419);
nand U1954 (N_1954,N_755,N_22);
and U1955 (N_1955,N_826,N_558);
nor U1956 (N_1956,N_321,N_523);
and U1957 (N_1957,N_641,N_16);
or U1958 (N_1958,N_785,N_991);
nor U1959 (N_1959,N_651,N_334);
xor U1960 (N_1960,N_312,N_474);
nand U1961 (N_1961,N_764,N_551);
and U1962 (N_1962,N_41,N_197);
nand U1963 (N_1963,N_65,N_966);
nor U1964 (N_1964,N_941,N_22);
or U1965 (N_1965,N_524,N_655);
nor U1966 (N_1966,N_92,N_209);
nor U1967 (N_1967,N_86,N_363);
or U1968 (N_1968,N_537,N_749);
nor U1969 (N_1969,N_738,N_983);
or U1970 (N_1970,N_815,N_942);
xnor U1971 (N_1971,N_187,N_545);
xor U1972 (N_1972,N_512,N_813);
nor U1973 (N_1973,N_813,N_71);
xor U1974 (N_1974,N_914,N_506);
xnor U1975 (N_1975,N_413,N_434);
or U1976 (N_1976,N_89,N_76);
or U1977 (N_1977,N_120,N_603);
and U1978 (N_1978,N_852,N_221);
or U1979 (N_1979,N_591,N_247);
nand U1980 (N_1980,N_370,N_432);
xnor U1981 (N_1981,N_324,N_419);
and U1982 (N_1982,N_970,N_459);
or U1983 (N_1983,N_243,N_166);
and U1984 (N_1984,N_181,N_244);
nand U1985 (N_1985,N_315,N_21);
xnor U1986 (N_1986,N_635,N_419);
nor U1987 (N_1987,N_59,N_332);
or U1988 (N_1988,N_721,N_732);
nor U1989 (N_1989,N_810,N_816);
nor U1990 (N_1990,N_314,N_247);
nor U1991 (N_1991,N_756,N_874);
nand U1992 (N_1992,N_336,N_299);
nand U1993 (N_1993,N_193,N_201);
and U1994 (N_1994,N_103,N_82);
xnor U1995 (N_1995,N_705,N_747);
nor U1996 (N_1996,N_165,N_574);
and U1997 (N_1997,N_31,N_903);
or U1998 (N_1998,N_502,N_680);
and U1999 (N_1999,N_610,N_333);
or U2000 (N_2000,N_1135,N_1654);
nand U2001 (N_2001,N_1564,N_1958);
or U2002 (N_2002,N_1801,N_1287);
or U2003 (N_2003,N_1110,N_1972);
and U2004 (N_2004,N_1744,N_1204);
nor U2005 (N_2005,N_1427,N_1263);
xor U2006 (N_2006,N_1589,N_1656);
xor U2007 (N_2007,N_1239,N_1151);
and U2008 (N_2008,N_1673,N_1786);
or U2009 (N_2009,N_1219,N_1713);
nor U2010 (N_2010,N_1806,N_1399);
xor U2011 (N_2011,N_1864,N_1906);
nand U2012 (N_2012,N_1561,N_1061);
nor U2013 (N_2013,N_1192,N_1167);
nor U2014 (N_2014,N_1512,N_1523);
nand U2015 (N_2015,N_1752,N_1207);
and U2016 (N_2016,N_1105,N_1186);
nor U2017 (N_2017,N_1180,N_1229);
nor U2018 (N_2018,N_1118,N_1054);
nand U2019 (N_2019,N_1353,N_1246);
or U2020 (N_2020,N_1015,N_1435);
nand U2021 (N_2021,N_1819,N_1632);
nor U2022 (N_2022,N_1603,N_1761);
and U2023 (N_2023,N_1617,N_1874);
or U2024 (N_2024,N_1507,N_1657);
or U2025 (N_2025,N_1292,N_1362);
or U2026 (N_2026,N_1371,N_1441);
or U2027 (N_2027,N_1164,N_1606);
nor U2028 (N_2028,N_1058,N_1517);
or U2029 (N_2029,N_1974,N_1121);
or U2030 (N_2030,N_1176,N_1250);
or U2031 (N_2031,N_1496,N_1079);
nand U2032 (N_2032,N_1500,N_1854);
nor U2033 (N_2033,N_1950,N_1882);
xnor U2034 (N_2034,N_1501,N_1962);
nand U2035 (N_2035,N_1634,N_1067);
nor U2036 (N_2036,N_1818,N_1934);
xnor U2037 (N_2037,N_1579,N_1807);
or U2038 (N_2038,N_1072,N_1382);
and U2039 (N_2039,N_1442,N_1374);
nand U2040 (N_2040,N_1877,N_1297);
nor U2041 (N_2041,N_1799,N_1554);
and U2042 (N_2042,N_1392,N_1381);
or U2043 (N_2043,N_1059,N_1691);
and U2044 (N_2044,N_1948,N_1965);
xnor U2045 (N_2045,N_1081,N_1481);
and U2046 (N_2046,N_1770,N_1754);
nand U2047 (N_2047,N_1134,N_1094);
xnor U2048 (N_2048,N_1391,N_1790);
nand U2049 (N_2049,N_1393,N_1581);
and U2050 (N_2050,N_1111,N_1420);
or U2051 (N_2051,N_1217,N_1194);
or U2052 (N_2052,N_1064,N_1910);
nor U2053 (N_2053,N_1650,N_1060);
or U2054 (N_2054,N_1339,N_1991);
xnor U2055 (N_2055,N_1244,N_1596);
nor U2056 (N_2056,N_1970,N_1921);
nor U2057 (N_2057,N_1548,N_1719);
nor U2058 (N_2058,N_1023,N_1705);
nand U2059 (N_2059,N_1325,N_1289);
nand U2060 (N_2060,N_1933,N_1089);
xor U2061 (N_2061,N_1628,N_1115);
nor U2062 (N_2062,N_1326,N_1275);
and U2063 (N_2063,N_1995,N_1421);
nor U2064 (N_2064,N_1723,N_1710);
nand U2065 (N_2065,N_1791,N_1891);
xor U2066 (N_2066,N_1739,N_1988);
and U2067 (N_2067,N_1711,N_1964);
nand U2068 (N_2068,N_1935,N_1919);
xor U2069 (N_2069,N_1528,N_1549);
nand U2070 (N_2070,N_1671,N_1722);
nand U2071 (N_2071,N_1133,N_1778);
and U2072 (N_2072,N_1859,N_1458);
xnor U2073 (N_2073,N_1439,N_1084);
xnor U2074 (N_2074,N_1471,N_1021);
xnor U2075 (N_2075,N_1216,N_1300);
or U2076 (N_2076,N_1355,N_1234);
nand U2077 (N_2077,N_1759,N_1994);
xor U2078 (N_2078,N_1815,N_1411);
nand U2079 (N_2079,N_1301,N_1526);
xnor U2080 (N_2080,N_1652,N_1210);
xnor U2081 (N_2081,N_1363,N_1558);
nand U2082 (N_2082,N_1259,N_1197);
xnor U2083 (N_2083,N_1459,N_1572);
or U2084 (N_2084,N_1655,N_1712);
and U2085 (N_2085,N_1651,N_1847);
or U2086 (N_2086,N_1456,N_1677);
or U2087 (N_2087,N_1174,N_1211);
nand U2088 (N_2088,N_1044,N_1403);
xnor U2089 (N_2089,N_1117,N_1334);
and U2090 (N_2090,N_1205,N_1062);
or U2091 (N_2091,N_1667,N_1880);
and U2092 (N_2092,N_1405,N_1227);
nor U2093 (N_2093,N_1980,N_1073);
nand U2094 (N_2094,N_1502,N_1514);
xnor U2095 (N_2095,N_1622,N_1727);
and U2096 (N_2096,N_1413,N_1758);
and U2097 (N_2097,N_1398,N_1510);
nor U2098 (N_2098,N_1269,N_1230);
nand U2099 (N_2099,N_1123,N_1085);
nor U2100 (N_2100,N_1542,N_1930);
xnor U2101 (N_2101,N_1175,N_1020);
or U2102 (N_2102,N_1714,N_1258);
and U2103 (N_2103,N_1647,N_1237);
nor U2104 (N_2104,N_1843,N_1530);
or U2105 (N_2105,N_1503,N_1648);
nand U2106 (N_2106,N_1899,N_1741);
or U2107 (N_2107,N_1277,N_1763);
xor U2108 (N_2108,N_1742,N_1241);
xor U2109 (N_2109,N_1975,N_1698);
and U2110 (N_2110,N_1331,N_1373);
nor U2111 (N_2111,N_1346,N_1866);
and U2112 (N_2112,N_1139,N_1488);
nand U2113 (N_2113,N_1011,N_1700);
nor U2114 (N_2114,N_1840,N_1137);
nand U2115 (N_2115,N_1850,N_1593);
or U2116 (N_2116,N_1003,N_1206);
and U2117 (N_2117,N_1920,N_1482);
or U2118 (N_2118,N_1889,N_1896);
or U2119 (N_2119,N_1341,N_1315);
nand U2120 (N_2120,N_1328,N_1783);
and U2121 (N_2121,N_1417,N_1963);
and U2122 (N_2122,N_1120,N_1016);
or U2123 (N_2123,N_1423,N_1360);
nor U2124 (N_2124,N_1922,N_1702);
nand U2125 (N_2125,N_1693,N_1412);
nand U2126 (N_2126,N_1279,N_1369);
xor U2127 (N_2127,N_1836,N_1352);
xnor U2128 (N_2128,N_1822,N_1943);
and U2129 (N_2129,N_1150,N_1418);
and U2130 (N_2130,N_1157,N_1303);
or U2131 (N_2131,N_1096,N_1795);
xnor U2132 (N_2132,N_1956,N_1440);
and U2133 (N_2133,N_1706,N_1235);
and U2134 (N_2134,N_1366,N_1156);
nand U2135 (N_2135,N_1479,N_1898);
or U2136 (N_2136,N_1116,N_1051);
nand U2137 (N_2137,N_1878,N_1871);
nor U2138 (N_2138,N_1766,N_1903);
xnor U2139 (N_2139,N_1979,N_1254);
and U2140 (N_2140,N_1132,N_1001);
and U2141 (N_2141,N_1681,N_1597);
nor U2142 (N_2142,N_1356,N_1213);
nand U2143 (N_2143,N_1773,N_1911);
xor U2144 (N_2144,N_1637,N_1200);
nand U2145 (N_2145,N_1358,N_1469);
nand U2146 (N_2146,N_1624,N_1686);
nand U2147 (N_2147,N_1784,N_1747);
nand U2148 (N_2148,N_1406,N_1097);
nor U2149 (N_2149,N_1344,N_1868);
or U2150 (N_2150,N_1971,N_1128);
nor U2151 (N_2151,N_1779,N_1689);
or U2152 (N_2152,N_1875,N_1426);
and U2153 (N_2153,N_1893,N_1857);
and U2154 (N_2154,N_1154,N_1886);
nor U2155 (N_2155,N_1050,N_1290);
and U2156 (N_2156,N_1944,N_1809);
or U2157 (N_2157,N_1811,N_1319);
nor U2158 (N_2158,N_1661,N_1342);
or U2159 (N_2159,N_1890,N_1845);
xnor U2160 (N_2160,N_1224,N_1915);
and U2161 (N_2161,N_1453,N_1794);
or U2162 (N_2162,N_1080,N_1546);
xor U2163 (N_2163,N_1796,N_1335);
or U2164 (N_2164,N_1019,N_1566);
or U2165 (N_2165,N_1800,N_1639);
and U2166 (N_2166,N_1031,N_1165);
xor U2167 (N_2167,N_1422,N_1372);
or U2168 (N_2168,N_1040,N_1643);
xnor U2169 (N_2169,N_1627,N_1273);
nor U2170 (N_2170,N_1102,N_1900);
or U2171 (N_2171,N_1489,N_1272);
nand U2172 (N_2172,N_1131,N_1522);
or U2173 (N_2173,N_1613,N_1513);
nand U2174 (N_2174,N_1155,N_1070);
and U2175 (N_2175,N_1692,N_1136);
and U2176 (N_2176,N_1295,N_1484);
xnor U2177 (N_2177,N_1798,N_1788);
nand U2178 (N_2178,N_1872,N_1029);
nand U2179 (N_2179,N_1166,N_1856);
nand U2180 (N_2180,N_1262,N_1498);
or U2181 (N_2181,N_1386,N_1032);
xnor U2182 (N_2182,N_1475,N_1521);
nor U2183 (N_2183,N_1495,N_1443);
and U2184 (N_2184,N_1619,N_1179);
and U2185 (N_2185,N_1104,N_1033);
and U2186 (N_2186,N_1220,N_1483);
and U2187 (N_2187,N_1183,N_1867);
xor U2188 (N_2188,N_1126,N_1537);
and U2189 (N_2189,N_1846,N_1336);
nand U2190 (N_2190,N_1370,N_1214);
xor U2191 (N_2191,N_1480,N_1068);
and U2192 (N_2192,N_1887,N_1114);
and U2193 (N_2193,N_1583,N_1129);
nand U2194 (N_2194,N_1720,N_1284);
xor U2195 (N_2195,N_1680,N_1063);
or U2196 (N_2196,N_1828,N_1257);
or U2197 (N_2197,N_1379,N_1309);
and U2198 (N_2198,N_1749,N_1924);
and U2199 (N_2199,N_1009,N_1873);
or U2200 (N_2200,N_1242,N_1598);
nor U2201 (N_2201,N_1993,N_1573);
or U2202 (N_2202,N_1715,N_1238);
nand U2203 (N_2203,N_1738,N_1999);
xnor U2204 (N_2204,N_1494,N_1519);
nand U2205 (N_2205,N_1380,N_1000);
and U2206 (N_2206,N_1223,N_1960);
and U2207 (N_2207,N_1983,N_1076);
nor U2208 (N_2208,N_1041,N_1550);
nor U2209 (N_2209,N_1330,N_1493);
nor U2210 (N_2210,N_1644,N_1557);
or U2211 (N_2211,N_1853,N_1106);
xnor U2212 (N_2212,N_1143,N_1416);
or U2213 (N_2213,N_1474,N_1078);
and U2214 (N_2214,N_1045,N_1551);
nor U2215 (N_2215,N_1168,N_1082);
nand U2216 (N_2216,N_1574,N_1347);
and U2217 (N_2217,N_1532,N_1035);
or U2218 (N_2218,N_1695,N_1193);
nand U2219 (N_2219,N_1071,N_1961);
xor U2220 (N_2220,N_1225,N_1232);
nor U2221 (N_2221,N_1535,N_1043);
and U2222 (N_2222,N_1954,N_1101);
or U2223 (N_2223,N_1833,N_1343);
nor U2224 (N_2224,N_1669,N_1236);
nand U2225 (N_2225,N_1696,N_1320);
and U2226 (N_2226,N_1536,N_1146);
nand U2227 (N_2227,N_1685,N_1614);
or U2228 (N_2228,N_1985,N_1264);
or U2229 (N_2229,N_1345,N_1162);
nand U2230 (N_2230,N_1946,N_1865);
xor U2231 (N_2231,N_1305,N_1444);
nand U2232 (N_2232,N_1547,N_1732);
nor U2233 (N_2233,N_1780,N_1490);
nor U2234 (N_2234,N_1879,N_1316);
xnor U2235 (N_2235,N_1725,N_1083);
and U2236 (N_2236,N_1861,N_1375);
or U2237 (N_2237,N_1728,N_1226);
or U2238 (N_2238,N_1916,N_1195);
xnor U2239 (N_2239,N_1088,N_1701);
nor U2240 (N_2240,N_1945,N_1631);
or U2241 (N_2241,N_1383,N_1976);
and U2242 (N_2242,N_1539,N_1604);
xor U2243 (N_2243,N_1929,N_1559);
nor U2244 (N_2244,N_1670,N_1449);
xor U2245 (N_2245,N_1048,N_1317);
or U2246 (N_2246,N_1308,N_1580);
or U2247 (N_2247,N_1772,N_1602);
or U2248 (N_2248,N_1529,N_1830);
nor U2249 (N_2249,N_1428,N_1684);
and U2250 (N_2250,N_1322,N_1311);
nand U2251 (N_2251,N_1672,N_1595);
or U2252 (N_2252,N_1454,N_1895);
or U2253 (N_2253,N_1432,N_1737);
or U2254 (N_2254,N_1208,N_1568);
and U2255 (N_2255,N_1491,N_1577);
and U2256 (N_2256,N_1851,N_1473);
nand U2257 (N_2257,N_1268,N_1966);
or U2258 (N_2258,N_1987,N_1608);
nor U2259 (N_2259,N_1802,N_1171);
xnor U2260 (N_2260,N_1074,N_1407);
and U2261 (N_2261,N_1265,N_1858);
and U2262 (N_2262,N_1090,N_1760);
xnor U2263 (N_2263,N_1683,N_1576);
nor U2264 (N_2264,N_1108,N_1447);
nand U2265 (N_2265,N_1302,N_1626);
nand U2266 (N_2266,N_1461,N_1615);
or U2267 (N_2267,N_1247,N_1282);
xor U2268 (N_2268,N_1429,N_1455);
or U2269 (N_2269,N_1823,N_1756);
and U2270 (N_2270,N_1928,N_1173);
or U2271 (N_2271,N_1694,N_1560);
nand U2272 (N_2272,N_1927,N_1863);
or U2273 (N_2273,N_1037,N_1792);
nor U2274 (N_2274,N_1401,N_1951);
xor U2275 (N_2275,N_1952,N_1007);
or U2276 (N_2276,N_1034,N_1027);
and U2277 (N_2277,N_1431,N_1520);
and U2278 (N_2278,N_1485,N_1942);
xnor U2279 (N_2279,N_1046,N_1189);
xnor U2280 (N_2280,N_1797,N_1022);
or U2281 (N_2281,N_1486,N_1757);
xor U2282 (N_2282,N_1251,N_1787);
xor U2283 (N_2283,N_1184,N_1645);
or U2284 (N_2284,N_1607,N_1190);
xor U2285 (N_2285,N_1909,N_1629);
and U2286 (N_2286,N_1552,N_1842);
and U2287 (N_2287,N_1625,N_1803);
xnor U2288 (N_2288,N_1069,N_1782);
xnor U2289 (N_2289,N_1582,N_1450);
and U2290 (N_2290,N_1812,N_1771);
xnor U2291 (N_2291,N_1017,N_1077);
or U2292 (N_2292,N_1215,N_1814);
and U2293 (N_2293,N_1394,N_1018);
nor U2294 (N_2294,N_1904,N_1902);
nand U2295 (N_2295,N_1404,N_1623);
and U2296 (N_2296,N_1735,N_1775);
nor U2297 (N_2297,N_1565,N_1437);
or U2298 (N_2298,N_1182,N_1294);
nand U2299 (N_2299,N_1389,N_1938);
nor U2300 (N_2300,N_1518,N_1152);
nand U2301 (N_2301,N_1410,N_1233);
or U2302 (N_2302,N_1914,N_1989);
xnor U2303 (N_2303,N_1107,N_1053);
nor U2304 (N_2304,N_1688,N_1533);
and U2305 (N_2305,N_1468,N_1313);
nand U2306 (N_2306,N_1387,N_1704);
nand U2307 (N_2307,N_1271,N_1436);
nor U2308 (N_2308,N_1203,N_1820);
or U2309 (N_2309,N_1438,N_1885);
or U2310 (N_2310,N_1364,N_1159);
or U2311 (N_2311,N_1025,N_1524);
or U2312 (N_2312,N_1913,N_1841);
xor U2313 (N_2313,N_1030,N_1630);
and U2314 (N_2314,N_1968,N_1746);
nor U2315 (N_2315,N_1912,N_1460);
nor U2316 (N_2316,N_1977,N_1119);
nand U2317 (N_2317,N_1222,N_1147);
nor U2318 (N_2318,N_1354,N_1620);
nor U2319 (N_2319,N_1047,N_1141);
nand U2320 (N_2320,N_1296,N_1953);
and U2321 (N_2321,N_1026,N_1751);
nand U2322 (N_2322,N_1897,N_1709);
and U2323 (N_2323,N_1361,N_1452);
nand U2324 (N_2324,N_1299,N_1451);
xnor U2325 (N_2325,N_1824,N_1445);
or U2326 (N_2326,N_1066,N_1270);
or U2327 (N_2327,N_1492,N_1286);
nor U2328 (N_2328,N_1351,N_1767);
nor U2329 (N_2329,N_1570,N_1649);
nand U2330 (N_2330,N_1855,N_1612);
nand U2331 (N_2331,N_1641,N_1196);
and U2332 (N_2332,N_1837,N_1562);
xor U2333 (N_2333,N_1553,N_1396);
or U2334 (N_2334,N_1969,N_1973);
and U2335 (N_2335,N_1957,N_1726);
or U2336 (N_2336,N_1789,N_1388);
and U2337 (N_2337,N_1594,N_1668);
or U2338 (N_2338,N_1285,N_1338);
or U2339 (N_2339,N_1584,N_1740);
or U2340 (N_2340,N_1831,N_1697);
nor U2341 (N_2341,N_1708,N_1377);
and U2342 (N_2342,N_1905,N_1663);
and U2343 (N_2343,N_1736,N_1984);
and U2344 (N_2344,N_1243,N_1327);
nand U2345 (N_2345,N_1092,N_1038);
and U2346 (N_2346,N_1130,N_1724);
nor U2347 (N_2347,N_1636,N_1433);
nor U2348 (N_2348,N_1590,N_1609);
or U2349 (N_2349,N_1218,N_1172);
nor U2350 (N_2350,N_1091,N_1281);
or U2351 (N_2351,N_1348,N_1690);
nor U2352 (N_2352,N_1476,N_1753);
nand U2353 (N_2353,N_1918,N_1013);
nor U2354 (N_2354,N_1505,N_1506);
nor U2355 (N_2355,N_1653,N_1252);
xor U2356 (N_2356,N_1256,N_1306);
xor U2357 (N_2357,N_1199,N_1852);
nand U2358 (N_2358,N_1087,N_1959);
nor U2359 (N_2359,N_1099,N_1333);
nand U2360 (N_2360,N_1276,N_1848);
and U2361 (N_2361,N_1642,N_1042);
and U2362 (N_2362,N_1178,N_1810);
and U2363 (N_2363,N_1587,N_1312);
xnor U2364 (N_2364,N_1621,N_1240);
nand U2365 (N_2365,N_1310,N_1384);
nor U2366 (N_2366,N_1996,N_1075);
nor U2367 (N_2367,N_1745,N_1158);
nand U2368 (N_2368,N_1527,N_1734);
and U2369 (N_2369,N_1478,N_1678);
nor U2370 (N_2370,N_1939,N_1253);
nand U2371 (N_2371,N_1635,N_1400);
nand U2372 (N_2372,N_1986,N_1765);
xor U2373 (N_2373,N_1997,N_1408);
or U2374 (N_2374,N_1395,N_1588);
or U2375 (N_2375,N_1161,N_1769);
nand U2376 (N_2376,N_1699,N_1004);
and U2377 (N_2377,N_1463,N_1298);
xor U2378 (N_2378,N_1002,N_1397);
nor U2379 (N_2379,N_1936,N_1144);
and U2380 (N_2380,N_1659,N_1640);
or U2381 (N_2381,N_1511,N_1926);
or U2382 (N_2382,N_1605,N_1777);
and U2383 (N_2383,N_1616,N_1876);
xor U2384 (N_2384,N_1563,N_1827);
xor U2385 (N_2385,N_1181,N_1884);
or U2386 (N_2386,N_1457,N_1764);
or U2387 (N_2387,N_1293,N_1274);
nor U2388 (N_2388,N_1228,N_1731);
and U2389 (N_2389,N_1055,N_1266);
or U2390 (N_2390,N_1005,N_1679);
nor U2391 (N_2391,N_1487,N_1221);
xnor U2392 (N_2392,N_1260,N_1967);
and U2393 (N_2393,N_1169,N_1349);
nor U2394 (N_2394,N_1600,N_1095);
or U2395 (N_2395,N_1212,N_1675);
xor U2396 (N_2396,N_1860,N_1755);
nand U2397 (N_2397,N_1267,N_1314);
or U2398 (N_2398,N_1955,N_1321);
nand U2399 (N_2399,N_1534,N_1231);
or U2400 (N_2400,N_1662,N_1940);
xor U2401 (N_2401,N_1012,N_1825);
nand U2402 (N_2402,N_1717,N_1065);
xor U2403 (N_2403,N_1470,N_1785);
xnor U2404 (N_2404,N_1467,N_1545);
or U2405 (N_2405,N_1531,N_1666);
nor U2406 (N_2406,N_1153,N_1359);
nor U2407 (N_2407,N_1056,N_1908);
nor U2408 (N_2408,N_1163,N_1508);
nand U2409 (N_2409,N_1881,N_1291);
nand U2410 (N_2410,N_1733,N_1808);
or U2411 (N_2411,N_1122,N_1776);
nand U2412 (N_2412,N_1086,N_1931);
or U2413 (N_2413,N_1592,N_1569);
nand U2414 (N_2414,N_1555,N_1992);
nor U2415 (N_2415,N_1743,N_1378);
nand U2416 (N_2416,N_1100,N_1591);
or U2417 (N_2417,N_1329,N_1368);
nor U2418 (N_2418,N_1504,N_1138);
and U2419 (N_2419,N_1805,N_1028);
and U2420 (N_2420,N_1248,N_1127);
xnor U2421 (N_2421,N_1280,N_1424);
xnor U2422 (N_2422,N_1525,N_1601);
nand U2423 (N_2423,N_1829,N_1448);
and U2424 (N_2424,N_1112,N_1198);
nor U2425 (N_2425,N_1124,N_1781);
and U2426 (N_2426,N_1892,N_1839);
and U2427 (N_2427,N_1148,N_1870);
nand U2428 (N_2428,N_1098,N_1010);
nor U2429 (N_2429,N_1888,N_1170);
xor U2430 (N_2430,N_1718,N_1835);
nor U2431 (N_2431,N_1611,N_1515);
or U2432 (N_2432,N_1462,N_1149);
or U2433 (N_2433,N_1419,N_1937);
or U2434 (N_2434,N_1177,N_1567);
nand U2435 (N_2435,N_1125,N_1323);
or U2436 (N_2436,N_1288,N_1466);
or U2437 (N_2437,N_1499,N_1385);
and U2438 (N_2438,N_1768,N_1707);
nand U2439 (N_2439,N_1014,N_1660);
nor U2440 (N_2440,N_1390,N_1367);
or U2441 (N_2441,N_1049,N_1923);
and U2442 (N_2442,N_1140,N_1730);
and U2443 (N_2443,N_1191,N_1729);
nand U2444 (N_2444,N_1665,N_1202);
or U2445 (N_2445,N_1516,N_1633);
and U2446 (N_2446,N_1185,N_1307);
nand U2447 (N_2447,N_1543,N_1610);
xnor U2448 (N_2448,N_1894,N_1978);
and U2449 (N_2449,N_1990,N_1465);
or U2450 (N_2450,N_1556,N_1674);
nor U2451 (N_2451,N_1816,N_1245);
and U2452 (N_2452,N_1332,N_1188);
and U2453 (N_2453,N_1917,N_1599);
nor U2454 (N_2454,N_1357,N_1703);
nand U2455 (N_2455,N_1261,N_1255);
or U2456 (N_2456,N_1834,N_1142);
nand U2457 (N_2457,N_1434,N_1981);
nor U2458 (N_2458,N_1844,N_1340);
nand U2459 (N_2459,N_1676,N_1425);
nor U2460 (N_2460,N_1402,N_1793);
and U2461 (N_2461,N_1052,N_1932);
nor U2462 (N_2462,N_1571,N_1409);
nand U2463 (N_2463,N_1509,N_1658);
nor U2464 (N_2464,N_1804,N_1249);
or U2465 (N_2465,N_1578,N_1838);
xnor U2466 (N_2466,N_1585,N_1664);
or U2467 (N_2467,N_1925,N_1716);
or U2468 (N_2468,N_1883,N_1721);
or U2469 (N_2469,N_1283,N_1774);
xnor U2470 (N_2470,N_1575,N_1145);
or U2471 (N_2471,N_1093,N_1541);
nor U2472 (N_2472,N_1949,N_1901);
xnor U2473 (N_2473,N_1618,N_1103);
or U2474 (N_2474,N_1039,N_1862);
nor U2475 (N_2475,N_1430,N_1324);
nor U2476 (N_2476,N_1036,N_1941);
or U2477 (N_2477,N_1376,N_1209);
xor U2478 (N_2478,N_1646,N_1472);
or U2479 (N_2479,N_1538,N_1817);
nor U2480 (N_2480,N_1982,N_1446);
nand U2481 (N_2481,N_1008,N_1497);
nor U2482 (N_2482,N_1414,N_1947);
nand U2483 (N_2483,N_1849,N_1907);
xor U2484 (N_2484,N_1832,N_1109);
and U2485 (N_2485,N_1337,N_1826);
or U2486 (N_2486,N_1160,N_1304);
and U2487 (N_2487,N_1687,N_1113);
or U2488 (N_2488,N_1024,N_1821);
or U2489 (N_2489,N_1006,N_1365);
and U2490 (N_2490,N_1540,N_1813);
xor U2491 (N_2491,N_1869,N_1748);
and U2492 (N_2492,N_1318,N_1682);
and U2493 (N_2493,N_1477,N_1998);
nor U2494 (N_2494,N_1187,N_1638);
and U2495 (N_2495,N_1350,N_1278);
xnor U2496 (N_2496,N_1057,N_1586);
nand U2497 (N_2497,N_1464,N_1201);
nor U2498 (N_2498,N_1415,N_1750);
and U2499 (N_2499,N_1762,N_1544);
nand U2500 (N_2500,N_1508,N_1284);
and U2501 (N_2501,N_1258,N_1958);
and U2502 (N_2502,N_1697,N_1155);
xor U2503 (N_2503,N_1179,N_1441);
or U2504 (N_2504,N_1644,N_1521);
xor U2505 (N_2505,N_1244,N_1959);
nand U2506 (N_2506,N_1528,N_1067);
xor U2507 (N_2507,N_1356,N_1584);
or U2508 (N_2508,N_1168,N_1970);
xnor U2509 (N_2509,N_1361,N_1500);
nor U2510 (N_2510,N_1870,N_1415);
xor U2511 (N_2511,N_1048,N_1585);
and U2512 (N_2512,N_1264,N_1505);
xnor U2513 (N_2513,N_1216,N_1038);
and U2514 (N_2514,N_1394,N_1890);
and U2515 (N_2515,N_1576,N_1285);
xnor U2516 (N_2516,N_1875,N_1753);
or U2517 (N_2517,N_1083,N_1775);
nor U2518 (N_2518,N_1336,N_1063);
or U2519 (N_2519,N_1096,N_1128);
xor U2520 (N_2520,N_1822,N_1416);
or U2521 (N_2521,N_1018,N_1329);
nand U2522 (N_2522,N_1993,N_1746);
and U2523 (N_2523,N_1245,N_1056);
or U2524 (N_2524,N_1184,N_1192);
nor U2525 (N_2525,N_1879,N_1103);
nor U2526 (N_2526,N_1805,N_1978);
and U2527 (N_2527,N_1840,N_1522);
nor U2528 (N_2528,N_1944,N_1876);
nor U2529 (N_2529,N_1237,N_1437);
xnor U2530 (N_2530,N_1462,N_1376);
or U2531 (N_2531,N_1805,N_1076);
or U2532 (N_2532,N_1113,N_1801);
nor U2533 (N_2533,N_1036,N_1087);
nand U2534 (N_2534,N_1635,N_1343);
nor U2535 (N_2535,N_1121,N_1538);
xnor U2536 (N_2536,N_1148,N_1213);
xnor U2537 (N_2537,N_1214,N_1152);
nand U2538 (N_2538,N_1721,N_1058);
or U2539 (N_2539,N_1759,N_1402);
nand U2540 (N_2540,N_1238,N_1610);
and U2541 (N_2541,N_1782,N_1171);
nand U2542 (N_2542,N_1726,N_1250);
nand U2543 (N_2543,N_1158,N_1133);
nand U2544 (N_2544,N_1285,N_1845);
or U2545 (N_2545,N_1622,N_1841);
nand U2546 (N_2546,N_1507,N_1318);
xnor U2547 (N_2547,N_1927,N_1114);
xnor U2548 (N_2548,N_1956,N_1589);
and U2549 (N_2549,N_1469,N_1271);
xor U2550 (N_2550,N_1542,N_1777);
xnor U2551 (N_2551,N_1577,N_1875);
xnor U2552 (N_2552,N_1644,N_1524);
and U2553 (N_2553,N_1771,N_1940);
or U2554 (N_2554,N_1248,N_1607);
or U2555 (N_2555,N_1458,N_1614);
nand U2556 (N_2556,N_1994,N_1692);
nand U2557 (N_2557,N_1533,N_1901);
and U2558 (N_2558,N_1839,N_1345);
and U2559 (N_2559,N_1683,N_1852);
xnor U2560 (N_2560,N_1931,N_1106);
and U2561 (N_2561,N_1262,N_1359);
nor U2562 (N_2562,N_1533,N_1192);
and U2563 (N_2563,N_1646,N_1510);
and U2564 (N_2564,N_1947,N_1504);
nand U2565 (N_2565,N_1696,N_1526);
nand U2566 (N_2566,N_1530,N_1947);
or U2567 (N_2567,N_1826,N_1109);
nand U2568 (N_2568,N_1579,N_1801);
nand U2569 (N_2569,N_1188,N_1141);
or U2570 (N_2570,N_1506,N_1708);
xor U2571 (N_2571,N_1668,N_1278);
nand U2572 (N_2572,N_1560,N_1566);
xnor U2573 (N_2573,N_1445,N_1943);
xor U2574 (N_2574,N_1173,N_1895);
nand U2575 (N_2575,N_1647,N_1374);
nand U2576 (N_2576,N_1336,N_1738);
or U2577 (N_2577,N_1652,N_1712);
xnor U2578 (N_2578,N_1127,N_1357);
and U2579 (N_2579,N_1997,N_1736);
xnor U2580 (N_2580,N_1549,N_1771);
nand U2581 (N_2581,N_1578,N_1694);
xnor U2582 (N_2582,N_1525,N_1475);
xnor U2583 (N_2583,N_1754,N_1831);
and U2584 (N_2584,N_1759,N_1163);
or U2585 (N_2585,N_1257,N_1559);
or U2586 (N_2586,N_1604,N_1834);
xor U2587 (N_2587,N_1563,N_1154);
or U2588 (N_2588,N_1421,N_1200);
and U2589 (N_2589,N_1114,N_1316);
nand U2590 (N_2590,N_1277,N_1129);
or U2591 (N_2591,N_1609,N_1673);
nand U2592 (N_2592,N_1345,N_1474);
xnor U2593 (N_2593,N_1449,N_1509);
or U2594 (N_2594,N_1215,N_1693);
nand U2595 (N_2595,N_1391,N_1469);
nand U2596 (N_2596,N_1550,N_1062);
nand U2597 (N_2597,N_1121,N_1497);
and U2598 (N_2598,N_1735,N_1623);
nor U2599 (N_2599,N_1096,N_1616);
xor U2600 (N_2600,N_1041,N_1797);
xor U2601 (N_2601,N_1781,N_1153);
nand U2602 (N_2602,N_1878,N_1748);
xor U2603 (N_2603,N_1373,N_1771);
nor U2604 (N_2604,N_1416,N_1828);
or U2605 (N_2605,N_1514,N_1655);
and U2606 (N_2606,N_1194,N_1115);
nand U2607 (N_2607,N_1236,N_1277);
xor U2608 (N_2608,N_1134,N_1273);
xor U2609 (N_2609,N_1818,N_1504);
xnor U2610 (N_2610,N_1008,N_1033);
nand U2611 (N_2611,N_1356,N_1183);
nand U2612 (N_2612,N_1607,N_1820);
xor U2613 (N_2613,N_1972,N_1852);
xor U2614 (N_2614,N_1093,N_1107);
nor U2615 (N_2615,N_1833,N_1615);
nor U2616 (N_2616,N_1068,N_1779);
and U2617 (N_2617,N_1377,N_1307);
or U2618 (N_2618,N_1658,N_1133);
nand U2619 (N_2619,N_1356,N_1555);
xnor U2620 (N_2620,N_1696,N_1747);
nor U2621 (N_2621,N_1636,N_1964);
xor U2622 (N_2622,N_1997,N_1516);
and U2623 (N_2623,N_1209,N_1228);
and U2624 (N_2624,N_1012,N_1325);
and U2625 (N_2625,N_1738,N_1178);
nor U2626 (N_2626,N_1952,N_1144);
or U2627 (N_2627,N_1038,N_1174);
nor U2628 (N_2628,N_1797,N_1857);
nand U2629 (N_2629,N_1128,N_1339);
nor U2630 (N_2630,N_1589,N_1945);
xnor U2631 (N_2631,N_1090,N_1993);
nand U2632 (N_2632,N_1190,N_1519);
or U2633 (N_2633,N_1482,N_1851);
and U2634 (N_2634,N_1193,N_1716);
and U2635 (N_2635,N_1716,N_1759);
nor U2636 (N_2636,N_1536,N_1303);
xor U2637 (N_2637,N_1399,N_1785);
xor U2638 (N_2638,N_1285,N_1376);
xnor U2639 (N_2639,N_1638,N_1886);
xor U2640 (N_2640,N_1794,N_1789);
nor U2641 (N_2641,N_1578,N_1554);
and U2642 (N_2642,N_1179,N_1830);
and U2643 (N_2643,N_1574,N_1114);
and U2644 (N_2644,N_1350,N_1318);
or U2645 (N_2645,N_1724,N_1955);
xnor U2646 (N_2646,N_1840,N_1193);
and U2647 (N_2647,N_1184,N_1468);
nand U2648 (N_2648,N_1201,N_1609);
nor U2649 (N_2649,N_1791,N_1261);
nor U2650 (N_2650,N_1926,N_1915);
xor U2651 (N_2651,N_1363,N_1496);
nand U2652 (N_2652,N_1915,N_1213);
and U2653 (N_2653,N_1841,N_1249);
nor U2654 (N_2654,N_1198,N_1412);
or U2655 (N_2655,N_1317,N_1766);
xor U2656 (N_2656,N_1951,N_1406);
or U2657 (N_2657,N_1687,N_1812);
or U2658 (N_2658,N_1523,N_1186);
or U2659 (N_2659,N_1499,N_1889);
or U2660 (N_2660,N_1105,N_1682);
nor U2661 (N_2661,N_1094,N_1123);
xor U2662 (N_2662,N_1597,N_1055);
nor U2663 (N_2663,N_1134,N_1613);
xor U2664 (N_2664,N_1710,N_1106);
or U2665 (N_2665,N_1936,N_1596);
nand U2666 (N_2666,N_1653,N_1606);
and U2667 (N_2667,N_1467,N_1407);
nor U2668 (N_2668,N_1928,N_1519);
nand U2669 (N_2669,N_1195,N_1235);
nand U2670 (N_2670,N_1003,N_1954);
xor U2671 (N_2671,N_1806,N_1339);
xnor U2672 (N_2672,N_1955,N_1213);
nor U2673 (N_2673,N_1542,N_1861);
or U2674 (N_2674,N_1985,N_1344);
or U2675 (N_2675,N_1955,N_1102);
nand U2676 (N_2676,N_1362,N_1159);
nor U2677 (N_2677,N_1612,N_1978);
xor U2678 (N_2678,N_1828,N_1982);
xor U2679 (N_2679,N_1297,N_1547);
nor U2680 (N_2680,N_1832,N_1464);
or U2681 (N_2681,N_1024,N_1678);
and U2682 (N_2682,N_1220,N_1217);
nand U2683 (N_2683,N_1049,N_1828);
or U2684 (N_2684,N_1434,N_1485);
or U2685 (N_2685,N_1592,N_1765);
or U2686 (N_2686,N_1803,N_1922);
nor U2687 (N_2687,N_1073,N_1512);
and U2688 (N_2688,N_1702,N_1307);
xnor U2689 (N_2689,N_1678,N_1260);
or U2690 (N_2690,N_1181,N_1930);
xor U2691 (N_2691,N_1610,N_1993);
nand U2692 (N_2692,N_1506,N_1729);
xor U2693 (N_2693,N_1329,N_1809);
and U2694 (N_2694,N_1482,N_1721);
nand U2695 (N_2695,N_1381,N_1738);
or U2696 (N_2696,N_1177,N_1367);
xnor U2697 (N_2697,N_1678,N_1520);
nor U2698 (N_2698,N_1778,N_1420);
nand U2699 (N_2699,N_1832,N_1306);
nand U2700 (N_2700,N_1695,N_1778);
xnor U2701 (N_2701,N_1635,N_1437);
nand U2702 (N_2702,N_1059,N_1072);
and U2703 (N_2703,N_1068,N_1491);
and U2704 (N_2704,N_1801,N_1026);
xor U2705 (N_2705,N_1581,N_1253);
or U2706 (N_2706,N_1898,N_1407);
nand U2707 (N_2707,N_1964,N_1735);
nor U2708 (N_2708,N_1280,N_1785);
xor U2709 (N_2709,N_1657,N_1951);
xor U2710 (N_2710,N_1315,N_1435);
and U2711 (N_2711,N_1288,N_1735);
xor U2712 (N_2712,N_1071,N_1753);
nand U2713 (N_2713,N_1398,N_1192);
xnor U2714 (N_2714,N_1387,N_1728);
or U2715 (N_2715,N_1992,N_1453);
and U2716 (N_2716,N_1900,N_1254);
nand U2717 (N_2717,N_1302,N_1891);
or U2718 (N_2718,N_1031,N_1727);
nand U2719 (N_2719,N_1707,N_1333);
xor U2720 (N_2720,N_1741,N_1206);
xnor U2721 (N_2721,N_1975,N_1346);
nor U2722 (N_2722,N_1824,N_1357);
or U2723 (N_2723,N_1241,N_1137);
nor U2724 (N_2724,N_1532,N_1368);
nor U2725 (N_2725,N_1543,N_1595);
xor U2726 (N_2726,N_1235,N_1530);
nor U2727 (N_2727,N_1487,N_1622);
xor U2728 (N_2728,N_1659,N_1996);
or U2729 (N_2729,N_1726,N_1097);
nand U2730 (N_2730,N_1958,N_1705);
or U2731 (N_2731,N_1031,N_1935);
nand U2732 (N_2732,N_1974,N_1004);
or U2733 (N_2733,N_1136,N_1685);
nor U2734 (N_2734,N_1703,N_1143);
nor U2735 (N_2735,N_1026,N_1694);
nor U2736 (N_2736,N_1779,N_1635);
nor U2737 (N_2737,N_1275,N_1027);
and U2738 (N_2738,N_1732,N_1756);
xnor U2739 (N_2739,N_1271,N_1813);
nor U2740 (N_2740,N_1268,N_1550);
and U2741 (N_2741,N_1540,N_1947);
nor U2742 (N_2742,N_1842,N_1863);
nand U2743 (N_2743,N_1980,N_1666);
nor U2744 (N_2744,N_1336,N_1601);
and U2745 (N_2745,N_1305,N_1085);
nor U2746 (N_2746,N_1710,N_1325);
nand U2747 (N_2747,N_1435,N_1334);
nor U2748 (N_2748,N_1584,N_1367);
nand U2749 (N_2749,N_1333,N_1137);
and U2750 (N_2750,N_1072,N_1602);
nand U2751 (N_2751,N_1864,N_1595);
or U2752 (N_2752,N_1049,N_1792);
or U2753 (N_2753,N_1917,N_1489);
or U2754 (N_2754,N_1486,N_1193);
xor U2755 (N_2755,N_1499,N_1987);
or U2756 (N_2756,N_1138,N_1688);
nor U2757 (N_2757,N_1906,N_1966);
xnor U2758 (N_2758,N_1995,N_1574);
or U2759 (N_2759,N_1451,N_1195);
xnor U2760 (N_2760,N_1825,N_1793);
nand U2761 (N_2761,N_1508,N_1077);
xnor U2762 (N_2762,N_1021,N_1199);
nor U2763 (N_2763,N_1936,N_1276);
nor U2764 (N_2764,N_1145,N_1218);
or U2765 (N_2765,N_1751,N_1282);
nor U2766 (N_2766,N_1469,N_1678);
nor U2767 (N_2767,N_1575,N_1982);
xor U2768 (N_2768,N_1161,N_1376);
and U2769 (N_2769,N_1925,N_1988);
nand U2770 (N_2770,N_1274,N_1359);
nand U2771 (N_2771,N_1874,N_1179);
xnor U2772 (N_2772,N_1860,N_1579);
xor U2773 (N_2773,N_1546,N_1376);
and U2774 (N_2774,N_1155,N_1755);
and U2775 (N_2775,N_1708,N_1833);
nand U2776 (N_2776,N_1669,N_1514);
nand U2777 (N_2777,N_1113,N_1913);
and U2778 (N_2778,N_1448,N_1431);
nor U2779 (N_2779,N_1304,N_1219);
or U2780 (N_2780,N_1504,N_1604);
xor U2781 (N_2781,N_1973,N_1374);
xor U2782 (N_2782,N_1379,N_1530);
or U2783 (N_2783,N_1223,N_1837);
xnor U2784 (N_2784,N_1653,N_1418);
xnor U2785 (N_2785,N_1016,N_1009);
nand U2786 (N_2786,N_1520,N_1049);
or U2787 (N_2787,N_1524,N_1388);
and U2788 (N_2788,N_1722,N_1788);
nor U2789 (N_2789,N_1265,N_1956);
nor U2790 (N_2790,N_1083,N_1483);
nor U2791 (N_2791,N_1454,N_1066);
and U2792 (N_2792,N_1875,N_1537);
or U2793 (N_2793,N_1574,N_1928);
or U2794 (N_2794,N_1547,N_1985);
xor U2795 (N_2795,N_1963,N_1551);
nand U2796 (N_2796,N_1353,N_1267);
and U2797 (N_2797,N_1688,N_1571);
or U2798 (N_2798,N_1402,N_1480);
or U2799 (N_2799,N_1314,N_1970);
and U2800 (N_2800,N_1917,N_1421);
nor U2801 (N_2801,N_1251,N_1285);
nand U2802 (N_2802,N_1462,N_1345);
and U2803 (N_2803,N_1631,N_1312);
nor U2804 (N_2804,N_1803,N_1759);
nor U2805 (N_2805,N_1933,N_1439);
nand U2806 (N_2806,N_1726,N_1022);
nand U2807 (N_2807,N_1258,N_1399);
xnor U2808 (N_2808,N_1894,N_1043);
and U2809 (N_2809,N_1017,N_1718);
nor U2810 (N_2810,N_1823,N_1377);
and U2811 (N_2811,N_1866,N_1843);
or U2812 (N_2812,N_1698,N_1880);
nand U2813 (N_2813,N_1741,N_1543);
xnor U2814 (N_2814,N_1361,N_1082);
or U2815 (N_2815,N_1728,N_1373);
nor U2816 (N_2816,N_1117,N_1262);
nand U2817 (N_2817,N_1188,N_1984);
or U2818 (N_2818,N_1970,N_1996);
or U2819 (N_2819,N_1004,N_1525);
nand U2820 (N_2820,N_1342,N_1481);
or U2821 (N_2821,N_1224,N_1002);
xnor U2822 (N_2822,N_1277,N_1211);
xnor U2823 (N_2823,N_1704,N_1086);
nor U2824 (N_2824,N_1022,N_1288);
nor U2825 (N_2825,N_1969,N_1165);
xor U2826 (N_2826,N_1446,N_1832);
nand U2827 (N_2827,N_1319,N_1949);
nor U2828 (N_2828,N_1979,N_1499);
nand U2829 (N_2829,N_1163,N_1088);
nor U2830 (N_2830,N_1785,N_1543);
nand U2831 (N_2831,N_1044,N_1086);
and U2832 (N_2832,N_1613,N_1506);
nand U2833 (N_2833,N_1842,N_1383);
nor U2834 (N_2834,N_1218,N_1354);
and U2835 (N_2835,N_1941,N_1325);
nand U2836 (N_2836,N_1353,N_1364);
and U2837 (N_2837,N_1653,N_1700);
and U2838 (N_2838,N_1895,N_1306);
and U2839 (N_2839,N_1168,N_1818);
nor U2840 (N_2840,N_1106,N_1659);
xor U2841 (N_2841,N_1283,N_1066);
xor U2842 (N_2842,N_1736,N_1389);
and U2843 (N_2843,N_1557,N_1852);
and U2844 (N_2844,N_1767,N_1382);
nor U2845 (N_2845,N_1830,N_1608);
nor U2846 (N_2846,N_1881,N_1089);
or U2847 (N_2847,N_1707,N_1673);
nor U2848 (N_2848,N_1111,N_1201);
or U2849 (N_2849,N_1733,N_1873);
xnor U2850 (N_2850,N_1147,N_1250);
and U2851 (N_2851,N_1877,N_1622);
and U2852 (N_2852,N_1910,N_1076);
nor U2853 (N_2853,N_1204,N_1132);
or U2854 (N_2854,N_1846,N_1883);
xnor U2855 (N_2855,N_1459,N_1275);
and U2856 (N_2856,N_1396,N_1828);
xnor U2857 (N_2857,N_1248,N_1505);
xnor U2858 (N_2858,N_1870,N_1986);
nand U2859 (N_2859,N_1028,N_1178);
xnor U2860 (N_2860,N_1871,N_1708);
xor U2861 (N_2861,N_1421,N_1588);
or U2862 (N_2862,N_1978,N_1974);
nand U2863 (N_2863,N_1778,N_1360);
or U2864 (N_2864,N_1239,N_1267);
or U2865 (N_2865,N_1516,N_1811);
nor U2866 (N_2866,N_1299,N_1594);
nor U2867 (N_2867,N_1988,N_1725);
nor U2868 (N_2868,N_1591,N_1086);
and U2869 (N_2869,N_1421,N_1462);
or U2870 (N_2870,N_1078,N_1081);
nor U2871 (N_2871,N_1942,N_1189);
nand U2872 (N_2872,N_1446,N_1853);
and U2873 (N_2873,N_1471,N_1394);
nor U2874 (N_2874,N_1716,N_1179);
nand U2875 (N_2875,N_1780,N_1125);
xnor U2876 (N_2876,N_1244,N_1550);
nor U2877 (N_2877,N_1942,N_1401);
nor U2878 (N_2878,N_1691,N_1792);
and U2879 (N_2879,N_1977,N_1449);
or U2880 (N_2880,N_1833,N_1057);
and U2881 (N_2881,N_1487,N_1963);
xnor U2882 (N_2882,N_1290,N_1419);
xnor U2883 (N_2883,N_1775,N_1434);
and U2884 (N_2884,N_1346,N_1414);
nor U2885 (N_2885,N_1220,N_1571);
xnor U2886 (N_2886,N_1905,N_1119);
xor U2887 (N_2887,N_1511,N_1887);
nand U2888 (N_2888,N_1056,N_1648);
nand U2889 (N_2889,N_1143,N_1193);
or U2890 (N_2890,N_1648,N_1250);
and U2891 (N_2891,N_1099,N_1410);
xor U2892 (N_2892,N_1925,N_1484);
or U2893 (N_2893,N_1196,N_1710);
xnor U2894 (N_2894,N_1893,N_1368);
nor U2895 (N_2895,N_1816,N_1806);
nor U2896 (N_2896,N_1105,N_1657);
nand U2897 (N_2897,N_1511,N_1378);
nand U2898 (N_2898,N_1018,N_1475);
or U2899 (N_2899,N_1242,N_1425);
and U2900 (N_2900,N_1375,N_1516);
or U2901 (N_2901,N_1852,N_1942);
or U2902 (N_2902,N_1536,N_1817);
and U2903 (N_2903,N_1343,N_1333);
or U2904 (N_2904,N_1196,N_1025);
nor U2905 (N_2905,N_1248,N_1174);
nor U2906 (N_2906,N_1257,N_1934);
and U2907 (N_2907,N_1836,N_1869);
xor U2908 (N_2908,N_1150,N_1926);
or U2909 (N_2909,N_1469,N_1882);
nor U2910 (N_2910,N_1642,N_1608);
xnor U2911 (N_2911,N_1927,N_1542);
xnor U2912 (N_2912,N_1185,N_1722);
and U2913 (N_2913,N_1434,N_1695);
nand U2914 (N_2914,N_1057,N_1389);
xor U2915 (N_2915,N_1738,N_1723);
and U2916 (N_2916,N_1130,N_1809);
or U2917 (N_2917,N_1096,N_1408);
xor U2918 (N_2918,N_1898,N_1797);
and U2919 (N_2919,N_1043,N_1048);
xnor U2920 (N_2920,N_1133,N_1378);
and U2921 (N_2921,N_1013,N_1360);
nand U2922 (N_2922,N_1995,N_1657);
nor U2923 (N_2923,N_1809,N_1589);
and U2924 (N_2924,N_1220,N_1849);
or U2925 (N_2925,N_1729,N_1915);
or U2926 (N_2926,N_1728,N_1565);
and U2927 (N_2927,N_1056,N_1820);
nand U2928 (N_2928,N_1639,N_1372);
or U2929 (N_2929,N_1771,N_1057);
or U2930 (N_2930,N_1420,N_1201);
and U2931 (N_2931,N_1452,N_1588);
nor U2932 (N_2932,N_1745,N_1277);
xor U2933 (N_2933,N_1599,N_1027);
or U2934 (N_2934,N_1821,N_1306);
xnor U2935 (N_2935,N_1738,N_1472);
or U2936 (N_2936,N_1986,N_1251);
xnor U2937 (N_2937,N_1651,N_1354);
xor U2938 (N_2938,N_1046,N_1515);
or U2939 (N_2939,N_1164,N_1973);
xnor U2940 (N_2940,N_1968,N_1118);
or U2941 (N_2941,N_1759,N_1971);
and U2942 (N_2942,N_1141,N_1747);
nand U2943 (N_2943,N_1742,N_1061);
or U2944 (N_2944,N_1787,N_1269);
nor U2945 (N_2945,N_1842,N_1760);
xnor U2946 (N_2946,N_1452,N_1597);
nor U2947 (N_2947,N_1971,N_1890);
xnor U2948 (N_2948,N_1573,N_1225);
nor U2949 (N_2949,N_1365,N_1112);
xor U2950 (N_2950,N_1451,N_1438);
or U2951 (N_2951,N_1385,N_1094);
xor U2952 (N_2952,N_1701,N_1017);
or U2953 (N_2953,N_1248,N_1126);
nand U2954 (N_2954,N_1029,N_1960);
and U2955 (N_2955,N_1153,N_1966);
nand U2956 (N_2956,N_1660,N_1398);
or U2957 (N_2957,N_1317,N_1110);
nand U2958 (N_2958,N_1781,N_1107);
or U2959 (N_2959,N_1512,N_1996);
nand U2960 (N_2960,N_1516,N_1152);
nor U2961 (N_2961,N_1454,N_1225);
nor U2962 (N_2962,N_1115,N_1811);
nor U2963 (N_2963,N_1226,N_1988);
and U2964 (N_2964,N_1832,N_1859);
and U2965 (N_2965,N_1400,N_1962);
or U2966 (N_2966,N_1042,N_1537);
nand U2967 (N_2967,N_1726,N_1802);
nand U2968 (N_2968,N_1608,N_1708);
nor U2969 (N_2969,N_1669,N_1192);
nand U2970 (N_2970,N_1027,N_1367);
or U2971 (N_2971,N_1230,N_1579);
and U2972 (N_2972,N_1744,N_1953);
nand U2973 (N_2973,N_1219,N_1261);
xnor U2974 (N_2974,N_1670,N_1719);
and U2975 (N_2975,N_1522,N_1874);
and U2976 (N_2976,N_1595,N_1219);
xnor U2977 (N_2977,N_1883,N_1241);
and U2978 (N_2978,N_1783,N_1387);
nor U2979 (N_2979,N_1050,N_1503);
nand U2980 (N_2980,N_1176,N_1815);
or U2981 (N_2981,N_1931,N_1729);
or U2982 (N_2982,N_1795,N_1695);
and U2983 (N_2983,N_1346,N_1908);
nand U2984 (N_2984,N_1589,N_1709);
or U2985 (N_2985,N_1930,N_1658);
xnor U2986 (N_2986,N_1157,N_1721);
nand U2987 (N_2987,N_1271,N_1969);
nand U2988 (N_2988,N_1735,N_1069);
or U2989 (N_2989,N_1078,N_1086);
or U2990 (N_2990,N_1008,N_1233);
or U2991 (N_2991,N_1099,N_1002);
and U2992 (N_2992,N_1059,N_1794);
nor U2993 (N_2993,N_1902,N_1033);
nor U2994 (N_2994,N_1044,N_1548);
or U2995 (N_2995,N_1956,N_1856);
xnor U2996 (N_2996,N_1204,N_1320);
nor U2997 (N_2997,N_1444,N_1725);
nand U2998 (N_2998,N_1192,N_1732);
or U2999 (N_2999,N_1421,N_1870);
and U3000 (N_3000,N_2245,N_2412);
xor U3001 (N_3001,N_2901,N_2104);
or U3002 (N_3002,N_2920,N_2409);
or U3003 (N_3003,N_2532,N_2498);
and U3004 (N_3004,N_2921,N_2310);
and U3005 (N_3005,N_2088,N_2678);
and U3006 (N_3006,N_2876,N_2798);
xor U3007 (N_3007,N_2361,N_2894);
nor U3008 (N_3008,N_2270,N_2283);
and U3009 (N_3009,N_2148,N_2114);
xor U3010 (N_3010,N_2181,N_2644);
nor U3011 (N_3011,N_2708,N_2555);
and U3012 (N_3012,N_2426,N_2237);
or U3013 (N_3013,N_2354,N_2761);
xor U3014 (N_3014,N_2500,N_2360);
xor U3015 (N_3015,N_2024,N_2556);
and U3016 (N_3016,N_2186,N_2472);
or U3017 (N_3017,N_2868,N_2036);
nor U3018 (N_3018,N_2201,N_2030);
and U3019 (N_3019,N_2497,N_2552);
nand U3020 (N_3020,N_2390,N_2255);
or U3021 (N_3021,N_2162,N_2840);
and U3022 (N_3022,N_2548,N_2022);
and U3023 (N_3023,N_2690,N_2624);
xnor U3024 (N_3024,N_2281,N_2356);
or U3025 (N_3025,N_2913,N_2608);
and U3026 (N_3026,N_2466,N_2735);
nor U3027 (N_3027,N_2067,N_2371);
xnor U3028 (N_3028,N_2776,N_2630);
nor U3029 (N_3029,N_2530,N_2531);
or U3030 (N_3030,N_2886,N_2347);
and U3031 (N_3031,N_2192,N_2247);
and U3032 (N_3032,N_2625,N_2597);
or U3033 (N_3033,N_2895,N_2955);
and U3034 (N_3034,N_2916,N_2286);
nand U3035 (N_3035,N_2642,N_2570);
or U3036 (N_3036,N_2438,N_2001);
nand U3037 (N_3037,N_2284,N_2378);
and U3038 (N_3038,N_2587,N_2646);
nor U3039 (N_3039,N_2989,N_2662);
nor U3040 (N_3040,N_2871,N_2524);
and U3041 (N_3041,N_2990,N_2723);
or U3042 (N_3042,N_2206,N_2097);
nor U3043 (N_3043,N_2892,N_2002);
or U3044 (N_3044,N_2471,N_2401);
and U3045 (N_3045,N_2359,N_2197);
nor U3046 (N_3046,N_2134,N_2758);
nor U3047 (N_3047,N_2170,N_2838);
nor U3048 (N_3048,N_2963,N_2043);
or U3049 (N_3049,N_2818,N_2275);
and U3050 (N_3050,N_2020,N_2804);
or U3051 (N_3051,N_2261,N_2098);
and U3052 (N_3052,N_2559,N_2504);
or U3053 (N_3053,N_2138,N_2700);
nor U3054 (N_3054,N_2883,N_2828);
and U3055 (N_3055,N_2567,N_2307);
xnor U3056 (N_3056,N_2054,N_2077);
xnor U3057 (N_3057,N_2660,N_2793);
nand U3058 (N_3058,N_2364,N_2156);
nor U3059 (N_3059,N_2533,N_2739);
nand U3060 (N_3060,N_2899,N_2317);
nand U3061 (N_3061,N_2745,N_2953);
or U3062 (N_3062,N_2773,N_2659);
xnor U3063 (N_3063,N_2262,N_2824);
and U3064 (N_3064,N_2334,N_2976);
or U3065 (N_3065,N_2414,N_2175);
xnor U3066 (N_3066,N_2765,N_2004);
and U3067 (N_3067,N_2127,N_2720);
nand U3068 (N_3068,N_2211,N_2740);
and U3069 (N_3069,N_2044,N_2606);
xor U3070 (N_3070,N_2130,N_2468);
or U3071 (N_3071,N_2943,N_2609);
nand U3072 (N_3072,N_2223,N_2415);
nand U3073 (N_3073,N_2975,N_2995);
xor U3074 (N_3074,N_2259,N_2189);
and U3075 (N_3075,N_2785,N_2406);
xnor U3076 (N_3076,N_2357,N_2389);
nand U3077 (N_3077,N_2458,N_2183);
nand U3078 (N_3078,N_2509,N_2935);
or U3079 (N_3079,N_2198,N_2946);
and U3080 (N_3080,N_2711,N_2638);
xor U3081 (N_3081,N_2507,N_2431);
nand U3082 (N_3082,N_2305,N_2381);
xnor U3083 (N_3083,N_2515,N_2537);
and U3084 (N_3084,N_2382,N_2521);
and U3085 (N_3085,N_2578,N_2163);
xnor U3086 (N_3086,N_2568,N_2397);
xor U3087 (N_3087,N_2264,N_2141);
or U3088 (N_3088,N_2376,N_2082);
nor U3089 (N_3089,N_2948,N_2404);
nor U3090 (N_3090,N_2228,N_2734);
nand U3091 (N_3091,N_2332,N_2658);
nand U3092 (N_3092,N_2058,N_2151);
nand U3093 (N_3093,N_2103,N_2577);
or U3094 (N_3094,N_2794,N_2726);
nand U3095 (N_3095,N_2834,N_2819);
xor U3096 (N_3096,N_2591,N_2462);
xnor U3097 (N_3097,N_2128,N_2959);
nand U3098 (N_3098,N_2105,N_2657);
xor U3099 (N_3099,N_2028,N_2408);
and U3100 (N_3100,N_2905,N_2047);
and U3101 (N_3101,N_2949,N_2633);
nor U3102 (N_3102,N_2122,N_2550);
nor U3103 (N_3103,N_2096,N_2790);
xnor U3104 (N_3104,N_2212,N_2979);
xor U3105 (N_3105,N_2852,N_2987);
or U3106 (N_3106,N_2450,N_2825);
and U3107 (N_3107,N_2807,N_2801);
nand U3108 (N_3108,N_2250,N_2144);
or U3109 (N_3109,N_2427,N_2200);
or U3110 (N_3110,N_2847,N_2319);
and U3111 (N_3111,N_2117,N_2488);
nor U3112 (N_3112,N_2111,N_2984);
nor U3113 (N_3113,N_2226,N_2266);
nand U3114 (N_3114,N_2210,N_2900);
or U3115 (N_3115,N_2499,N_2049);
or U3116 (N_3116,N_2338,N_2874);
xnor U3117 (N_3117,N_2831,N_2444);
and U3118 (N_3118,N_2733,N_2214);
nand U3119 (N_3119,N_2322,N_2491);
xnor U3120 (N_3120,N_2229,N_2246);
and U3121 (N_3121,N_2309,N_2551);
xnor U3122 (N_3122,N_2716,N_2039);
nand U3123 (N_3123,N_2118,N_2083);
or U3124 (N_3124,N_2437,N_2586);
nand U3125 (N_3125,N_2289,N_2355);
or U3126 (N_3126,N_2321,N_2326);
or U3127 (N_3127,N_2749,N_2903);
or U3128 (N_3128,N_2506,N_2493);
xnor U3129 (N_3129,N_2610,N_2421);
nand U3130 (N_3130,N_2405,N_2031);
or U3131 (N_3131,N_2486,N_2854);
or U3132 (N_3132,N_2782,N_2299);
nor U3133 (N_3133,N_2033,N_2712);
nor U3134 (N_3134,N_2452,N_2669);
nand U3135 (N_3135,N_2812,N_2000);
nor U3136 (N_3136,N_2403,N_2861);
nand U3137 (N_3137,N_2285,N_2072);
or U3138 (N_3138,N_2554,N_2387);
xnor U3139 (N_3139,N_2652,N_2196);
nor U3140 (N_3140,N_2126,N_2243);
and U3141 (N_3141,N_2702,N_2553);
or U3142 (N_3142,N_2827,N_2124);
or U3143 (N_3143,N_2327,N_2947);
xnor U3144 (N_3144,N_2062,N_2683);
xor U3145 (N_3145,N_2675,N_2475);
and U3146 (N_3146,N_2057,N_2641);
or U3147 (N_3147,N_2867,N_2316);
nor U3148 (N_3148,N_2590,N_2153);
xor U3149 (N_3149,N_2454,N_2649);
and U3150 (N_3150,N_2188,N_2460);
nor U3151 (N_3151,N_2816,N_2983);
nor U3152 (N_3152,N_2593,N_2168);
nand U3153 (N_3153,N_2686,N_2908);
nor U3154 (N_3154,N_2269,N_2166);
nor U3155 (N_3155,N_2887,N_2388);
or U3156 (N_3156,N_2737,N_2417);
and U3157 (N_3157,N_2048,N_2003);
and U3158 (N_3158,N_2121,N_2050);
nand U3159 (N_3159,N_2687,N_2012);
or U3160 (N_3160,N_2394,N_2337);
or U3161 (N_3161,N_2306,N_2843);
or U3162 (N_3162,N_2923,N_2482);
nand U3163 (N_3163,N_2607,N_2191);
nor U3164 (N_3164,N_2025,N_2557);
and U3165 (N_3165,N_2177,N_2396);
nor U3166 (N_3166,N_2015,N_2046);
nor U3167 (N_3167,N_2994,N_2848);
nand U3168 (N_3168,N_2034,N_2215);
nand U3169 (N_3169,N_2313,N_2194);
and U3170 (N_3170,N_2767,N_2370);
or U3171 (N_3171,N_2724,N_2845);
nand U3172 (N_3172,N_2013,N_2742);
and U3173 (N_3173,N_2407,N_2418);
nor U3174 (N_3174,N_2679,N_2068);
nand U3175 (N_3175,N_2330,N_2677);
nor U3176 (N_3176,N_2703,N_2091);
nor U3177 (N_3177,N_2231,N_2187);
xor U3178 (N_3178,N_2879,N_2732);
or U3179 (N_3179,N_2650,N_2511);
and U3180 (N_3180,N_2293,N_2563);
and U3181 (N_3181,N_2489,N_2547);
nor U3182 (N_3182,N_2478,N_2341);
or U3183 (N_3183,N_2169,N_2008);
nand U3184 (N_3184,N_2235,N_2143);
or U3185 (N_3185,N_2435,N_2997);
xnor U3186 (N_3186,N_2622,N_2932);
xnor U3187 (N_3187,N_2907,N_2584);
and U3188 (N_3188,N_2171,N_2353);
nand U3189 (N_3189,N_2743,N_2654);
nand U3190 (N_3190,N_2569,N_2797);
and U3191 (N_3191,N_2398,N_2695);
nand U3192 (N_3192,N_2224,N_2830);
nand U3193 (N_3193,N_2157,N_2674);
nor U3194 (N_3194,N_2236,N_2914);
nand U3195 (N_3195,N_2910,N_2693);
nand U3196 (N_3196,N_2463,N_2855);
nand U3197 (N_3197,N_2277,N_2872);
and U3198 (N_3198,N_2996,N_2069);
or U3199 (N_3199,N_2960,N_2333);
xnor U3200 (N_3200,N_2342,N_2882);
nor U3201 (N_3201,N_2931,N_2912);
nand U3202 (N_3202,N_2026,N_2680);
nand U3203 (N_3203,N_2070,N_2779);
or U3204 (N_3204,N_2549,N_2795);
xor U3205 (N_3205,N_2629,N_2086);
or U3206 (N_3206,N_2271,N_2813);
nand U3207 (N_3207,N_2564,N_2526);
nand U3208 (N_3208,N_2073,N_2560);
and U3209 (N_3209,N_2494,N_2799);
or U3210 (N_3210,N_2623,N_2320);
or U3211 (N_3211,N_2393,N_2451);
nor U3212 (N_3212,N_2880,N_2926);
nor U3213 (N_3213,N_2640,N_2936);
and U3214 (N_3214,N_2752,N_2656);
and U3215 (N_3215,N_2081,N_2736);
and U3216 (N_3216,N_2185,N_2889);
xnor U3217 (N_3217,N_2545,N_2216);
and U3218 (N_3218,N_2572,N_2826);
and U3219 (N_3219,N_2273,N_2856);
or U3220 (N_3220,N_2915,N_2479);
or U3221 (N_3221,N_2676,N_2006);
nand U3222 (N_3222,N_2257,N_2769);
xnor U3223 (N_3223,N_2512,N_2846);
or U3224 (N_3224,N_2328,N_2116);
nor U3225 (N_3225,N_2137,N_2029);
or U3226 (N_3226,N_2136,N_2434);
xnor U3227 (N_3227,N_2282,N_2694);
nor U3228 (N_3228,N_2222,N_2146);
and U3229 (N_3229,N_2254,N_2822);
and U3230 (N_3230,N_2350,N_2420);
nor U3231 (N_3231,N_2904,N_2585);
or U3232 (N_3232,N_2869,N_2325);
and U3233 (N_3233,N_2505,N_2052);
xnor U3234 (N_3234,N_2973,N_2476);
xnor U3235 (N_3235,N_2648,N_2783);
and U3236 (N_3236,N_2875,N_2707);
or U3237 (N_3237,N_2244,N_2358);
and U3238 (N_3238,N_2748,N_2429);
and U3239 (N_3239,N_2919,N_2534);
and U3240 (N_3240,N_2367,N_2614);
and U3241 (N_3241,N_2714,N_2589);
nand U3242 (N_3242,N_2579,N_2220);
nand U3243 (N_3243,N_2575,N_2823);
or U3244 (N_3244,N_2411,N_2730);
or U3245 (N_3245,N_2193,N_2635);
nor U3246 (N_3246,N_2670,N_2968);
nor U3247 (N_3247,N_2501,N_2777);
nand U3248 (N_3248,N_2351,N_2906);
or U3249 (N_3249,N_2965,N_2808);
nand U3250 (N_3250,N_2858,N_2841);
or U3251 (N_3251,N_2149,N_2303);
nand U3252 (N_3252,N_2032,N_2786);
nand U3253 (N_3253,N_2095,N_2014);
xor U3254 (N_3254,N_2422,N_2576);
nand U3255 (N_3255,N_2859,N_2380);
xor U3256 (N_3256,N_2815,N_2842);
and U3257 (N_3257,N_2469,N_2386);
and U3258 (N_3258,N_2789,N_2696);
and U3259 (N_3259,N_2538,N_2862);
xor U3260 (N_3260,N_2952,N_2035);
xnor U3261 (N_3261,N_2300,N_2115);
and U3262 (N_3262,N_2131,N_2304);
nor U3263 (N_3263,N_2203,N_2721);
xor U3264 (N_3264,N_2092,N_2150);
nand U3265 (N_3265,N_2084,N_2474);
or U3266 (N_3266,N_2268,N_2988);
and U3267 (N_3267,N_2541,N_2964);
nand U3268 (N_3268,N_2909,N_2839);
nor U3269 (N_3269,N_2562,N_2977);
and U3270 (N_3270,N_2287,N_2017);
and U3271 (N_3271,N_2957,N_2771);
and U3272 (N_3272,N_2911,N_2218);
nand U3273 (N_3273,N_2877,N_2011);
nor U3274 (N_3274,N_2445,N_2395);
xor U3275 (N_3275,N_2850,N_2249);
or U3276 (N_3276,N_2374,N_2490);
xor U3277 (N_3277,N_2836,N_2179);
and U3278 (N_3278,N_2992,N_2543);
and U3279 (N_3279,N_2164,N_2616);
or U3280 (N_3280,N_2159,N_2621);
and U3281 (N_3281,N_2123,N_2937);
or U3282 (N_3282,N_2385,N_2205);
xnor U3283 (N_3283,N_2125,N_2969);
nor U3284 (N_3284,N_2108,N_2517);
nor U3285 (N_3285,N_2612,N_2689);
or U3286 (N_3286,N_2535,N_2768);
or U3287 (N_3287,N_2542,N_2637);
xnor U3288 (N_3288,N_2204,N_2160);
and U3289 (N_3289,N_2558,N_2685);
xnor U3290 (N_3290,N_2738,N_2665);
nand U3291 (N_3291,N_2308,N_2312);
nand U3292 (N_3292,N_2573,N_2470);
xnor U3293 (N_3293,N_2448,N_2713);
or U3294 (N_3294,N_2784,N_2232);
xor U3295 (N_3295,N_2428,N_2966);
nor U3296 (N_3296,N_2722,N_2605);
nor U3297 (N_3297,N_2844,N_2918);
nand U3298 (N_3298,N_2864,N_2967);
and U3299 (N_3299,N_2230,N_2775);
nand U3300 (N_3300,N_2778,N_2618);
nor U3301 (N_3301,N_2750,N_2147);
and U3302 (N_3302,N_2898,N_2688);
xnor U3303 (N_3303,N_2941,N_2709);
nor U3304 (N_3304,N_2759,N_2480);
nand U3305 (N_3305,N_2094,N_2885);
or U3306 (N_3306,N_2484,N_2581);
nand U3307 (N_3307,N_2583,N_2888);
nand U3308 (N_3308,N_2391,N_2152);
or U3309 (N_3309,N_2087,N_2684);
or U3310 (N_3310,N_2772,N_2805);
nor U3311 (N_3311,N_2878,N_2917);
or U3312 (N_3312,N_2272,N_2719);
nor U3313 (N_3313,N_2315,N_2369);
nand U3314 (N_3314,N_2064,N_2061);
xnor U3315 (N_3315,N_2329,N_2705);
or U3316 (N_3316,N_2349,N_2529);
or U3317 (N_3317,N_2751,N_2718);
or U3318 (N_3318,N_2290,N_2076);
or U3319 (N_3319,N_2042,N_2433);
and U3320 (N_3320,N_2806,N_2296);
or U3321 (N_3321,N_2485,N_2717);
nand U3322 (N_3322,N_2741,N_2527);
nand U3323 (N_3323,N_2971,N_2110);
nor U3324 (N_3324,N_2671,N_2368);
xnor U3325 (N_3325,N_2851,N_2982);
and U3326 (N_3326,N_2167,N_2101);
and U3327 (N_3327,N_2755,N_2628);
or U3328 (N_3328,N_2710,N_2574);
and U3329 (N_3329,N_2063,N_2227);
xor U3330 (N_3330,N_2829,N_2986);
nand U3331 (N_3331,N_2544,N_2756);
or U3332 (N_3332,N_2725,N_2016);
nor U3333 (N_3333,N_2774,N_2155);
xor U3334 (N_3334,N_2757,N_2467);
nor U3335 (N_3335,N_2265,N_2496);
nor U3336 (N_3336,N_2252,N_2005);
or U3337 (N_3337,N_2100,N_2263);
nand U3338 (N_3338,N_2495,N_2803);
xor U3339 (N_3339,N_2985,N_2318);
or U3340 (N_3340,N_2199,N_2940);
and U3341 (N_3341,N_2344,N_2373);
nor U3342 (N_3342,N_2492,N_2365);
and U3343 (N_3343,N_2727,N_2375);
nand U3344 (N_3344,N_2040,N_2643);
nor U3345 (N_3345,N_2145,N_2972);
xor U3346 (N_3346,N_2787,N_2481);
nand U3347 (N_3347,N_2546,N_2837);
or U3348 (N_3348,N_2113,N_2863);
nor U3349 (N_3349,N_2881,N_2276);
nand U3350 (N_3350,N_2253,N_2956);
xor U3351 (N_3351,N_2619,N_2540);
nor U3352 (N_3352,N_2413,N_2377);
nor U3353 (N_3353,N_2580,N_2241);
nor U3354 (N_3354,N_2041,N_2811);
and U3355 (N_3355,N_2536,N_2184);
or U3356 (N_3356,N_2518,N_2446);
or U3357 (N_3357,N_2208,N_2279);
or U3358 (N_3358,N_2461,N_2933);
nand U3359 (N_3359,N_2440,N_2425);
or U3360 (N_3360,N_2256,N_2085);
or U3361 (N_3361,N_2664,N_2698);
nor U3362 (N_3362,N_2788,N_2833);
xnor U3363 (N_3363,N_2172,N_2951);
xor U3364 (N_3364,N_2860,N_2853);
or U3365 (N_3365,N_2372,N_2617);
and U3366 (N_3366,N_2673,N_2870);
xnor U3367 (N_3367,N_2423,N_2234);
xnor U3368 (N_3368,N_2345,N_2764);
or U3369 (N_3369,N_2217,N_2891);
xnor U3370 (N_3370,N_2945,N_2323);
xnor U3371 (N_3371,N_2502,N_2240);
xnor U3372 (N_3372,N_2007,N_2704);
xnor U3373 (N_3373,N_2582,N_2884);
nor U3374 (N_3374,N_2455,N_2636);
and U3375 (N_3375,N_2102,N_2295);
and U3376 (N_3376,N_2651,N_2439);
nand U3377 (N_3377,N_2219,N_2896);
nand U3378 (N_3378,N_2119,N_2419);
xnor U3379 (N_3379,N_2416,N_2950);
or U3380 (N_3380,N_2667,N_2139);
xor U3381 (N_3381,N_2280,N_2065);
nand U3382 (N_3382,N_2010,N_2561);
and U3383 (N_3383,N_2701,N_2897);
and U3384 (N_3384,N_2746,N_2078);
nor U3385 (N_3385,N_2075,N_2165);
xnor U3386 (N_3386,N_2132,N_2744);
xnor U3387 (N_3387,N_2929,N_2106);
xnor U3388 (N_3388,N_2056,N_2107);
xnor U3389 (N_3389,N_2592,N_2343);
and U3390 (N_3390,N_2457,N_2465);
nor U3391 (N_3391,N_2691,N_2443);
xnor U3392 (N_3392,N_2954,N_2729);
or U3393 (N_3393,N_2611,N_2161);
nand U3394 (N_3394,N_2780,N_2902);
or U3395 (N_3395,N_2302,N_2631);
xor U3396 (N_3396,N_2728,N_2348);
and U3397 (N_3397,N_2962,N_2278);
nor U3398 (N_3398,N_2666,N_2857);
nand U3399 (N_3399,N_2970,N_2681);
or U3400 (N_3400,N_2653,N_2634);
xor U3401 (N_3401,N_2301,N_2292);
nand U3402 (N_3402,N_2080,N_2384);
and U3403 (N_3403,N_2339,N_2632);
nand U3404 (N_3404,N_2849,N_2363);
nand U3405 (N_3405,N_2928,N_2938);
nand U3406 (N_3406,N_2958,N_2503);
nand U3407 (N_3407,N_2978,N_2991);
nand U3408 (N_3408,N_2516,N_2508);
nand U3409 (N_3409,N_2238,N_2038);
nand U3410 (N_3410,N_2598,N_2379);
xor U3411 (N_3411,N_2594,N_2449);
xor U3412 (N_3412,N_2291,N_2324);
nor U3413 (N_3413,N_2974,N_2865);
and U3414 (N_3414,N_2090,N_2093);
or U3415 (N_3415,N_2763,N_2209);
and U3416 (N_3416,N_2051,N_2835);
nor U3417 (N_3417,N_2615,N_2009);
xnor U3418 (N_3418,N_2174,N_2176);
xnor U3419 (N_3419,N_2890,N_2873);
xnor U3420 (N_3420,N_2999,N_2821);
and U3421 (N_3421,N_2021,N_2190);
or U3422 (N_3422,N_2655,N_2074);
nand U3423 (N_3423,N_2747,N_2523);
nor U3424 (N_3424,N_2258,N_2588);
and U3425 (N_3425,N_2399,N_2473);
or U3426 (N_3426,N_2601,N_2400);
and U3427 (N_3427,N_2762,N_2464);
xor U3428 (N_3428,N_2340,N_2980);
xnor U3429 (N_3429,N_2487,N_2142);
nand U3430 (N_3430,N_2925,N_2483);
nand U3431 (N_3431,N_2510,N_2055);
or U3432 (N_3432,N_2602,N_2297);
nor U3433 (N_3433,N_2770,N_2298);
xor U3434 (N_3434,N_2129,N_2934);
nand U3435 (N_3435,N_2753,N_2809);
xor U3436 (N_3436,N_2766,N_2993);
and U3437 (N_3437,N_2893,N_2314);
xnor U3438 (N_3438,N_2346,N_2331);
nor U3439 (N_3439,N_2663,N_2832);
or U3440 (N_3440,N_2383,N_2430);
xnor U3441 (N_3441,N_2441,N_2814);
or U3442 (N_3442,N_2519,N_2410);
or U3443 (N_3443,N_2796,N_2335);
xor U3444 (N_3444,N_2366,N_2682);
nand U3445 (N_3445,N_2599,N_2715);
and U3446 (N_3446,N_2311,N_2336);
and U3447 (N_3447,N_2288,N_2791);
nor U3448 (N_3448,N_2672,N_2178);
or U3449 (N_3449,N_2233,N_2447);
nor U3450 (N_3450,N_2639,N_2154);
nor U3451 (N_3451,N_2267,N_2424);
and U3452 (N_3452,N_2539,N_2754);
and U3453 (N_3453,N_2456,N_2513);
nor U3454 (N_3454,N_2866,N_2692);
or U3455 (N_3455,N_2019,N_2525);
or U3456 (N_3456,N_2221,N_2800);
and U3457 (N_3457,N_2626,N_2362);
nor U3458 (N_3458,N_2998,N_2613);
and U3459 (N_3459,N_2195,N_2180);
and U3460 (N_3460,N_2571,N_2242);
nor U3461 (N_3461,N_2731,N_2079);
xnor U3462 (N_3462,N_2699,N_2436);
or U3463 (N_3463,N_2453,N_2045);
nor U3464 (N_3464,N_2627,N_2939);
xor U3465 (N_3465,N_2661,N_2432);
nor U3466 (N_3466,N_2528,N_2158);
nor U3467 (N_3467,N_2930,N_2566);
and U3468 (N_3468,N_2792,N_2260);
or U3469 (N_3469,N_2202,N_2645);
nand U3470 (N_3470,N_2668,N_2520);
nor U3471 (N_3471,N_2459,N_2402);
or U3472 (N_3472,N_2239,N_2173);
nand U3473 (N_3473,N_2053,N_2182);
or U3474 (N_3474,N_2820,N_2251);
nand U3475 (N_3475,N_2135,N_2140);
nor U3476 (N_3476,N_2112,N_2477);
and U3477 (N_3477,N_2647,N_2213);
xor U3478 (N_3478,N_2944,N_2817);
and U3479 (N_3479,N_2089,N_2810);
or U3480 (N_3480,N_2059,N_2109);
xnor U3481 (N_3481,N_2802,N_2120);
nor U3482 (N_3482,N_2225,N_2274);
nand U3483 (N_3483,N_2922,N_2927);
xor U3484 (N_3484,N_2133,N_2924);
or U3485 (N_3485,N_2596,N_2352);
and U3486 (N_3486,N_2781,N_2604);
and U3487 (N_3487,N_2942,N_2442);
nor U3488 (N_3488,N_2706,N_2294);
nand U3489 (N_3489,N_2023,N_2981);
and U3490 (N_3490,N_2697,N_2760);
xor U3491 (N_3491,N_2099,N_2600);
nand U3492 (N_3492,N_2071,N_2066);
or U3493 (N_3493,N_2514,N_2595);
or U3494 (N_3494,N_2027,N_2392);
nand U3495 (N_3495,N_2522,N_2037);
xnor U3496 (N_3496,N_2018,N_2961);
or U3497 (N_3497,N_2060,N_2565);
or U3498 (N_3498,N_2207,N_2603);
nand U3499 (N_3499,N_2248,N_2620);
or U3500 (N_3500,N_2927,N_2925);
and U3501 (N_3501,N_2386,N_2392);
and U3502 (N_3502,N_2645,N_2289);
or U3503 (N_3503,N_2492,N_2277);
nand U3504 (N_3504,N_2415,N_2370);
and U3505 (N_3505,N_2569,N_2852);
and U3506 (N_3506,N_2183,N_2631);
nor U3507 (N_3507,N_2455,N_2496);
or U3508 (N_3508,N_2889,N_2457);
nand U3509 (N_3509,N_2970,N_2553);
or U3510 (N_3510,N_2741,N_2720);
nand U3511 (N_3511,N_2540,N_2030);
nand U3512 (N_3512,N_2090,N_2215);
nor U3513 (N_3513,N_2235,N_2955);
xnor U3514 (N_3514,N_2534,N_2330);
or U3515 (N_3515,N_2908,N_2082);
nand U3516 (N_3516,N_2689,N_2742);
nand U3517 (N_3517,N_2158,N_2035);
nand U3518 (N_3518,N_2141,N_2299);
xnor U3519 (N_3519,N_2815,N_2798);
nor U3520 (N_3520,N_2558,N_2011);
and U3521 (N_3521,N_2511,N_2182);
nand U3522 (N_3522,N_2755,N_2804);
xor U3523 (N_3523,N_2967,N_2849);
and U3524 (N_3524,N_2795,N_2214);
nand U3525 (N_3525,N_2488,N_2121);
and U3526 (N_3526,N_2015,N_2255);
nand U3527 (N_3527,N_2511,N_2750);
nor U3528 (N_3528,N_2886,N_2759);
or U3529 (N_3529,N_2882,N_2506);
or U3530 (N_3530,N_2020,N_2490);
xnor U3531 (N_3531,N_2504,N_2052);
and U3532 (N_3532,N_2997,N_2410);
xnor U3533 (N_3533,N_2821,N_2305);
nor U3534 (N_3534,N_2572,N_2847);
nand U3535 (N_3535,N_2348,N_2316);
xnor U3536 (N_3536,N_2240,N_2610);
nand U3537 (N_3537,N_2475,N_2269);
nand U3538 (N_3538,N_2425,N_2487);
nor U3539 (N_3539,N_2102,N_2800);
or U3540 (N_3540,N_2773,N_2784);
or U3541 (N_3541,N_2253,N_2734);
nand U3542 (N_3542,N_2778,N_2218);
xnor U3543 (N_3543,N_2076,N_2742);
nand U3544 (N_3544,N_2603,N_2018);
nand U3545 (N_3545,N_2063,N_2288);
xnor U3546 (N_3546,N_2190,N_2026);
nor U3547 (N_3547,N_2173,N_2054);
xnor U3548 (N_3548,N_2415,N_2166);
xnor U3549 (N_3549,N_2066,N_2137);
nor U3550 (N_3550,N_2285,N_2415);
nor U3551 (N_3551,N_2087,N_2949);
or U3552 (N_3552,N_2335,N_2185);
nor U3553 (N_3553,N_2978,N_2461);
nor U3554 (N_3554,N_2701,N_2322);
nand U3555 (N_3555,N_2573,N_2166);
nor U3556 (N_3556,N_2080,N_2566);
nand U3557 (N_3557,N_2334,N_2855);
nor U3558 (N_3558,N_2336,N_2676);
xnor U3559 (N_3559,N_2828,N_2351);
nand U3560 (N_3560,N_2180,N_2148);
nand U3561 (N_3561,N_2169,N_2934);
or U3562 (N_3562,N_2054,N_2102);
or U3563 (N_3563,N_2398,N_2468);
and U3564 (N_3564,N_2345,N_2651);
or U3565 (N_3565,N_2824,N_2342);
or U3566 (N_3566,N_2462,N_2753);
nor U3567 (N_3567,N_2219,N_2611);
nand U3568 (N_3568,N_2600,N_2068);
and U3569 (N_3569,N_2356,N_2062);
xor U3570 (N_3570,N_2231,N_2047);
nand U3571 (N_3571,N_2412,N_2188);
or U3572 (N_3572,N_2336,N_2270);
and U3573 (N_3573,N_2001,N_2079);
xor U3574 (N_3574,N_2557,N_2875);
nand U3575 (N_3575,N_2474,N_2118);
and U3576 (N_3576,N_2368,N_2933);
nand U3577 (N_3577,N_2000,N_2808);
nand U3578 (N_3578,N_2446,N_2698);
nand U3579 (N_3579,N_2850,N_2784);
nand U3580 (N_3580,N_2827,N_2315);
nand U3581 (N_3581,N_2209,N_2992);
nand U3582 (N_3582,N_2864,N_2296);
or U3583 (N_3583,N_2176,N_2812);
xor U3584 (N_3584,N_2666,N_2226);
xnor U3585 (N_3585,N_2899,N_2696);
or U3586 (N_3586,N_2810,N_2490);
and U3587 (N_3587,N_2993,N_2612);
and U3588 (N_3588,N_2807,N_2421);
or U3589 (N_3589,N_2616,N_2609);
and U3590 (N_3590,N_2679,N_2933);
nor U3591 (N_3591,N_2198,N_2621);
and U3592 (N_3592,N_2571,N_2788);
nor U3593 (N_3593,N_2390,N_2112);
xnor U3594 (N_3594,N_2261,N_2605);
or U3595 (N_3595,N_2627,N_2668);
nor U3596 (N_3596,N_2984,N_2940);
nand U3597 (N_3597,N_2512,N_2583);
or U3598 (N_3598,N_2122,N_2630);
nor U3599 (N_3599,N_2358,N_2575);
xor U3600 (N_3600,N_2845,N_2960);
nor U3601 (N_3601,N_2614,N_2702);
xor U3602 (N_3602,N_2528,N_2955);
nand U3603 (N_3603,N_2313,N_2046);
or U3604 (N_3604,N_2713,N_2667);
or U3605 (N_3605,N_2633,N_2840);
and U3606 (N_3606,N_2209,N_2482);
xor U3607 (N_3607,N_2166,N_2221);
and U3608 (N_3608,N_2005,N_2873);
nor U3609 (N_3609,N_2535,N_2433);
and U3610 (N_3610,N_2536,N_2549);
nor U3611 (N_3611,N_2976,N_2799);
or U3612 (N_3612,N_2716,N_2178);
or U3613 (N_3613,N_2017,N_2137);
nand U3614 (N_3614,N_2417,N_2171);
nor U3615 (N_3615,N_2239,N_2105);
or U3616 (N_3616,N_2125,N_2633);
and U3617 (N_3617,N_2665,N_2945);
and U3618 (N_3618,N_2327,N_2716);
nand U3619 (N_3619,N_2504,N_2014);
or U3620 (N_3620,N_2558,N_2128);
xor U3621 (N_3621,N_2733,N_2997);
and U3622 (N_3622,N_2412,N_2796);
or U3623 (N_3623,N_2841,N_2994);
xor U3624 (N_3624,N_2963,N_2066);
and U3625 (N_3625,N_2780,N_2175);
or U3626 (N_3626,N_2300,N_2466);
and U3627 (N_3627,N_2614,N_2111);
nor U3628 (N_3628,N_2362,N_2059);
xnor U3629 (N_3629,N_2645,N_2859);
or U3630 (N_3630,N_2519,N_2722);
or U3631 (N_3631,N_2978,N_2837);
or U3632 (N_3632,N_2777,N_2721);
or U3633 (N_3633,N_2042,N_2798);
and U3634 (N_3634,N_2363,N_2379);
or U3635 (N_3635,N_2020,N_2777);
nand U3636 (N_3636,N_2891,N_2585);
or U3637 (N_3637,N_2191,N_2042);
and U3638 (N_3638,N_2761,N_2982);
nor U3639 (N_3639,N_2119,N_2952);
nor U3640 (N_3640,N_2202,N_2017);
or U3641 (N_3641,N_2355,N_2027);
nand U3642 (N_3642,N_2151,N_2979);
and U3643 (N_3643,N_2803,N_2689);
nand U3644 (N_3644,N_2310,N_2046);
nand U3645 (N_3645,N_2936,N_2561);
nor U3646 (N_3646,N_2717,N_2529);
nand U3647 (N_3647,N_2763,N_2251);
nand U3648 (N_3648,N_2428,N_2653);
xnor U3649 (N_3649,N_2618,N_2027);
and U3650 (N_3650,N_2713,N_2571);
and U3651 (N_3651,N_2065,N_2326);
or U3652 (N_3652,N_2922,N_2797);
and U3653 (N_3653,N_2546,N_2913);
nor U3654 (N_3654,N_2896,N_2513);
and U3655 (N_3655,N_2220,N_2674);
or U3656 (N_3656,N_2693,N_2138);
and U3657 (N_3657,N_2872,N_2685);
nand U3658 (N_3658,N_2471,N_2160);
nand U3659 (N_3659,N_2967,N_2018);
or U3660 (N_3660,N_2030,N_2951);
and U3661 (N_3661,N_2693,N_2267);
and U3662 (N_3662,N_2080,N_2203);
nand U3663 (N_3663,N_2170,N_2043);
nor U3664 (N_3664,N_2154,N_2459);
or U3665 (N_3665,N_2723,N_2057);
or U3666 (N_3666,N_2195,N_2584);
nor U3667 (N_3667,N_2604,N_2865);
or U3668 (N_3668,N_2563,N_2444);
nand U3669 (N_3669,N_2307,N_2869);
and U3670 (N_3670,N_2375,N_2857);
nand U3671 (N_3671,N_2193,N_2874);
nor U3672 (N_3672,N_2797,N_2232);
and U3673 (N_3673,N_2259,N_2051);
and U3674 (N_3674,N_2546,N_2181);
xor U3675 (N_3675,N_2559,N_2940);
or U3676 (N_3676,N_2262,N_2859);
nor U3677 (N_3677,N_2291,N_2754);
and U3678 (N_3678,N_2474,N_2501);
or U3679 (N_3679,N_2782,N_2043);
nand U3680 (N_3680,N_2115,N_2698);
and U3681 (N_3681,N_2426,N_2441);
nand U3682 (N_3682,N_2027,N_2194);
or U3683 (N_3683,N_2680,N_2614);
nand U3684 (N_3684,N_2298,N_2939);
nor U3685 (N_3685,N_2615,N_2567);
nand U3686 (N_3686,N_2911,N_2020);
and U3687 (N_3687,N_2771,N_2900);
xor U3688 (N_3688,N_2260,N_2113);
nand U3689 (N_3689,N_2427,N_2791);
or U3690 (N_3690,N_2591,N_2312);
or U3691 (N_3691,N_2263,N_2257);
or U3692 (N_3692,N_2740,N_2622);
and U3693 (N_3693,N_2595,N_2211);
and U3694 (N_3694,N_2542,N_2459);
and U3695 (N_3695,N_2061,N_2809);
and U3696 (N_3696,N_2695,N_2677);
xnor U3697 (N_3697,N_2843,N_2344);
xnor U3698 (N_3698,N_2866,N_2719);
and U3699 (N_3699,N_2782,N_2275);
xnor U3700 (N_3700,N_2566,N_2595);
nand U3701 (N_3701,N_2186,N_2380);
nand U3702 (N_3702,N_2936,N_2985);
xor U3703 (N_3703,N_2402,N_2513);
nor U3704 (N_3704,N_2634,N_2208);
nor U3705 (N_3705,N_2271,N_2408);
nand U3706 (N_3706,N_2091,N_2152);
nor U3707 (N_3707,N_2422,N_2827);
and U3708 (N_3708,N_2388,N_2180);
and U3709 (N_3709,N_2778,N_2372);
nand U3710 (N_3710,N_2682,N_2179);
nor U3711 (N_3711,N_2228,N_2434);
and U3712 (N_3712,N_2106,N_2463);
or U3713 (N_3713,N_2584,N_2841);
xnor U3714 (N_3714,N_2317,N_2693);
nand U3715 (N_3715,N_2060,N_2441);
nand U3716 (N_3716,N_2452,N_2855);
or U3717 (N_3717,N_2820,N_2022);
and U3718 (N_3718,N_2145,N_2530);
and U3719 (N_3719,N_2499,N_2751);
and U3720 (N_3720,N_2686,N_2550);
and U3721 (N_3721,N_2422,N_2858);
nand U3722 (N_3722,N_2110,N_2144);
or U3723 (N_3723,N_2011,N_2918);
nand U3724 (N_3724,N_2776,N_2309);
and U3725 (N_3725,N_2654,N_2799);
and U3726 (N_3726,N_2514,N_2268);
nand U3727 (N_3727,N_2028,N_2249);
or U3728 (N_3728,N_2714,N_2669);
nor U3729 (N_3729,N_2386,N_2175);
or U3730 (N_3730,N_2733,N_2054);
and U3731 (N_3731,N_2180,N_2654);
xnor U3732 (N_3732,N_2888,N_2390);
nand U3733 (N_3733,N_2552,N_2532);
nand U3734 (N_3734,N_2688,N_2133);
or U3735 (N_3735,N_2059,N_2067);
or U3736 (N_3736,N_2999,N_2151);
nor U3737 (N_3737,N_2781,N_2270);
xor U3738 (N_3738,N_2529,N_2388);
and U3739 (N_3739,N_2483,N_2805);
or U3740 (N_3740,N_2382,N_2168);
and U3741 (N_3741,N_2382,N_2477);
xnor U3742 (N_3742,N_2252,N_2853);
nand U3743 (N_3743,N_2566,N_2097);
or U3744 (N_3744,N_2113,N_2892);
or U3745 (N_3745,N_2222,N_2071);
and U3746 (N_3746,N_2289,N_2800);
xnor U3747 (N_3747,N_2352,N_2400);
or U3748 (N_3748,N_2791,N_2324);
nand U3749 (N_3749,N_2463,N_2372);
nand U3750 (N_3750,N_2457,N_2105);
and U3751 (N_3751,N_2143,N_2806);
xor U3752 (N_3752,N_2779,N_2654);
nand U3753 (N_3753,N_2527,N_2772);
or U3754 (N_3754,N_2777,N_2079);
nor U3755 (N_3755,N_2963,N_2669);
nor U3756 (N_3756,N_2245,N_2004);
nor U3757 (N_3757,N_2407,N_2986);
nand U3758 (N_3758,N_2510,N_2490);
and U3759 (N_3759,N_2592,N_2462);
nor U3760 (N_3760,N_2547,N_2957);
nand U3761 (N_3761,N_2288,N_2793);
nand U3762 (N_3762,N_2171,N_2016);
or U3763 (N_3763,N_2411,N_2143);
and U3764 (N_3764,N_2704,N_2782);
xnor U3765 (N_3765,N_2350,N_2741);
nand U3766 (N_3766,N_2186,N_2939);
xnor U3767 (N_3767,N_2056,N_2804);
xor U3768 (N_3768,N_2780,N_2949);
or U3769 (N_3769,N_2660,N_2028);
or U3770 (N_3770,N_2203,N_2979);
and U3771 (N_3771,N_2014,N_2426);
nor U3772 (N_3772,N_2343,N_2460);
and U3773 (N_3773,N_2316,N_2043);
nor U3774 (N_3774,N_2005,N_2001);
and U3775 (N_3775,N_2275,N_2061);
and U3776 (N_3776,N_2372,N_2084);
nor U3777 (N_3777,N_2375,N_2453);
xnor U3778 (N_3778,N_2274,N_2376);
xnor U3779 (N_3779,N_2517,N_2138);
nor U3780 (N_3780,N_2725,N_2088);
xnor U3781 (N_3781,N_2899,N_2848);
nand U3782 (N_3782,N_2413,N_2627);
xnor U3783 (N_3783,N_2416,N_2885);
or U3784 (N_3784,N_2543,N_2123);
or U3785 (N_3785,N_2358,N_2713);
or U3786 (N_3786,N_2788,N_2083);
or U3787 (N_3787,N_2498,N_2608);
and U3788 (N_3788,N_2596,N_2740);
and U3789 (N_3789,N_2405,N_2733);
or U3790 (N_3790,N_2444,N_2248);
and U3791 (N_3791,N_2854,N_2736);
nor U3792 (N_3792,N_2678,N_2377);
nand U3793 (N_3793,N_2058,N_2057);
or U3794 (N_3794,N_2044,N_2211);
or U3795 (N_3795,N_2620,N_2622);
nor U3796 (N_3796,N_2141,N_2251);
and U3797 (N_3797,N_2228,N_2985);
nor U3798 (N_3798,N_2967,N_2321);
and U3799 (N_3799,N_2978,N_2774);
or U3800 (N_3800,N_2827,N_2183);
or U3801 (N_3801,N_2567,N_2582);
nand U3802 (N_3802,N_2809,N_2275);
nor U3803 (N_3803,N_2163,N_2779);
and U3804 (N_3804,N_2824,N_2591);
or U3805 (N_3805,N_2660,N_2689);
nor U3806 (N_3806,N_2413,N_2113);
or U3807 (N_3807,N_2253,N_2060);
nor U3808 (N_3808,N_2088,N_2080);
nand U3809 (N_3809,N_2106,N_2205);
xor U3810 (N_3810,N_2599,N_2488);
and U3811 (N_3811,N_2580,N_2868);
or U3812 (N_3812,N_2067,N_2494);
nand U3813 (N_3813,N_2550,N_2235);
nand U3814 (N_3814,N_2257,N_2756);
xor U3815 (N_3815,N_2810,N_2412);
or U3816 (N_3816,N_2378,N_2388);
xor U3817 (N_3817,N_2953,N_2074);
or U3818 (N_3818,N_2543,N_2090);
nand U3819 (N_3819,N_2782,N_2760);
nand U3820 (N_3820,N_2667,N_2132);
or U3821 (N_3821,N_2869,N_2924);
xnor U3822 (N_3822,N_2776,N_2123);
nand U3823 (N_3823,N_2938,N_2314);
and U3824 (N_3824,N_2520,N_2727);
nor U3825 (N_3825,N_2520,N_2839);
nor U3826 (N_3826,N_2283,N_2406);
xor U3827 (N_3827,N_2312,N_2188);
xor U3828 (N_3828,N_2132,N_2100);
and U3829 (N_3829,N_2020,N_2818);
nor U3830 (N_3830,N_2401,N_2961);
and U3831 (N_3831,N_2401,N_2088);
or U3832 (N_3832,N_2008,N_2846);
nor U3833 (N_3833,N_2835,N_2767);
or U3834 (N_3834,N_2698,N_2706);
nor U3835 (N_3835,N_2024,N_2858);
nand U3836 (N_3836,N_2264,N_2714);
xor U3837 (N_3837,N_2819,N_2382);
nand U3838 (N_3838,N_2112,N_2867);
or U3839 (N_3839,N_2479,N_2993);
xnor U3840 (N_3840,N_2082,N_2451);
or U3841 (N_3841,N_2465,N_2462);
and U3842 (N_3842,N_2074,N_2772);
nor U3843 (N_3843,N_2181,N_2579);
nor U3844 (N_3844,N_2945,N_2834);
xnor U3845 (N_3845,N_2753,N_2057);
xnor U3846 (N_3846,N_2873,N_2533);
xnor U3847 (N_3847,N_2589,N_2306);
and U3848 (N_3848,N_2578,N_2065);
nand U3849 (N_3849,N_2652,N_2628);
xor U3850 (N_3850,N_2377,N_2823);
nand U3851 (N_3851,N_2118,N_2374);
xnor U3852 (N_3852,N_2373,N_2222);
xnor U3853 (N_3853,N_2220,N_2639);
and U3854 (N_3854,N_2100,N_2360);
nor U3855 (N_3855,N_2876,N_2671);
nor U3856 (N_3856,N_2664,N_2179);
and U3857 (N_3857,N_2462,N_2654);
or U3858 (N_3858,N_2503,N_2699);
nor U3859 (N_3859,N_2736,N_2698);
nand U3860 (N_3860,N_2364,N_2446);
nor U3861 (N_3861,N_2769,N_2125);
or U3862 (N_3862,N_2844,N_2949);
or U3863 (N_3863,N_2938,N_2137);
and U3864 (N_3864,N_2359,N_2214);
and U3865 (N_3865,N_2466,N_2548);
and U3866 (N_3866,N_2504,N_2831);
xnor U3867 (N_3867,N_2319,N_2510);
nor U3868 (N_3868,N_2089,N_2902);
nand U3869 (N_3869,N_2900,N_2371);
and U3870 (N_3870,N_2478,N_2870);
nand U3871 (N_3871,N_2351,N_2676);
nor U3872 (N_3872,N_2136,N_2460);
nand U3873 (N_3873,N_2369,N_2686);
nand U3874 (N_3874,N_2570,N_2163);
nor U3875 (N_3875,N_2094,N_2824);
nand U3876 (N_3876,N_2375,N_2222);
and U3877 (N_3877,N_2305,N_2774);
nand U3878 (N_3878,N_2012,N_2753);
and U3879 (N_3879,N_2631,N_2462);
xor U3880 (N_3880,N_2462,N_2138);
or U3881 (N_3881,N_2453,N_2470);
nand U3882 (N_3882,N_2883,N_2202);
and U3883 (N_3883,N_2050,N_2739);
or U3884 (N_3884,N_2143,N_2944);
nor U3885 (N_3885,N_2063,N_2499);
and U3886 (N_3886,N_2770,N_2756);
nand U3887 (N_3887,N_2782,N_2473);
nor U3888 (N_3888,N_2498,N_2422);
nand U3889 (N_3889,N_2105,N_2525);
nor U3890 (N_3890,N_2487,N_2835);
xor U3891 (N_3891,N_2439,N_2967);
or U3892 (N_3892,N_2654,N_2777);
xor U3893 (N_3893,N_2326,N_2854);
xor U3894 (N_3894,N_2467,N_2172);
nor U3895 (N_3895,N_2861,N_2899);
nand U3896 (N_3896,N_2411,N_2300);
nor U3897 (N_3897,N_2077,N_2758);
nand U3898 (N_3898,N_2033,N_2740);
and U3899 (N_3899,N_2800,N_2566);
xor U3900 (N_3900,N_2768,N_2881);
and U3901 (N_3901,N_2575,N_2911);
nand U3902 (N_3902,N_2276,N_2407);
xor U3903 (N_3903,N_2307,N_2826);
nor U3904 (N_3904,N_2245,N_2633);
or U3905 (N_3905,N_2447,N_2031);
xor U3906 (N_3906,N_2080,N_2563);
or U3907 (N_3907,N_2260,N_2551);
or U3908 (N_3908,N_2747,N_2671);
nand U3909 (N_3909,N_2033,N_2710);
and U3910 (N_3910,N_2930,N_2638);
and U3911 (N_3911,N_2423,N_2769);
nand U3912 (N_3912,N_2352,N_2241);
nand U3913 (N_3913,N_2118,N_2012);
nand U3914 (N_3914,N_2293,N_2811);
and U3915 (N_3915,N_2295,N_2442);
nor U3916 (N_3916,N_2657,N_2518);
or U3917 (N_3917,N_2767,N_2058);
nand U3918 (N_3918,N_2298,N_2088);
or U3919 (N_3919,N_2663,N_2503);
xor U3920 (N_3920,N_2941,N_2638);
or U3921 (N_3921,N_2238,N_2588);
nor U3922 (N_3922,N_2917,N_2744);
nand U3923 (N_3923,N_2150,N_2057);
or U3924 (N_3924,N_2613,N_2073);
xor U3925 (N_3925,N_2379,N_2139);
xor U3926 (N_3926,N_2788,N_2036);
and U3927 (N_3927,N_2698,N_2382);
and U3928 (N_3928,N_2449,N_2649);
xnor U3929 (N_3929,N_2179,N_2714);
nor U3930 (N_3930,N_2180,N_2920);
xnor U3931 (N_3931,N_2075,N_2918);
or U3932 (N_3932,N_2459,N_2000);
nand U3933 (N_3933,N_2223,N_2212);
and U3934 (N_3934,N_2981,N_2409);
or U3935 (N_3935,N_2597,N_2944);
nand U3936 (N_3936,N_2897,N_2919);
xnor U3937 (N_3937,N_2423,N_2483);
and U3938 (N_3938,N_2273,N_2464);
nand U3939 (N_3939,N_2197,N_2532);
xnor U3940 (N_3940,N_2240,N_2010);
nor U3941 (N_3941,N_2502,N_2048);
xnor U3942 (N_3942,N_2511,N_2284);
nand U3943 (N_3943,N_2858,N_2485);
nor U3944 (N_3944,N_2492,N_2530);
nor U3945 (N_3945,N_2267,N_2378);
or U3946 (N_3946,N_2993,N_2650);
xnor U3947 (N_3947,N_2339,N_2873);
or U3948 (N_3948,N_2007,N_2459);
or U3949 (N_3949,N_2673,N_2539);
or U3950 (N_3950,N_2330,N_2910);
nand U3951 (N_3951,N_2603,N_2893);
nor U3952 (N_3952,N_2403,N_2738);
xor U3953 (N_3953,N_2608,N_2900);
and U3954 (N_3954,N_2821,N_2022);
or U3955 (N_3955,N_2760,N_2134);
or U3956 (N_3956,N_2008,N_2603);
nor U3957 (N_3957,N_2068,N_2290);
nor U3958 (N_3958,N_2896,N_2920);
nand U3959 (N_3959,N_2070,N_2891);
or U3960 (N_3960,N_2894,N_2410);
nor U3961 (N_3961,N_2051,N_2789);
nor U3962 (N_3962,N_2910,N_2067);
nand U3963 (N_3963,N_2020,N_2738);
nand U3964 (N_3964,N_2752,N_2467);
nand U3965 (N_3965,N_2207,N_2548);
or U3966 (N_3966,N_2711,N_2519);
nand U3967 (N_3967,N_2176,N_2894);
and U3968 (N_3968,N_2159,N_2436);
nor U3969 (N_3969,N_2342,N_2748);
and U3970 (N_3970,N_2967,N_2893);
xnor U3971 (N_3971,N_2332,N_2385);
nand U3972 (N_3972,N_2254,N_2729);
or U3973 (N_3973,N_2664,N_2902);
and U3974 (N_3974,N_2693,N_2178);
nand U3975 (N_3975,N_2705,N_2214);
and U3976 (N_3976,N_2169,N_2819);
nor U3977 (N_3977,N_2960,N_2998);
and U3978 (N_3978,N_2024,N_2971);
xnor U3979 (N_3979,N_2759,N_2580);
nor U3980 (N_3980,N_2779,N_2922);
nand U3981 (N_3981,N_2676,N_2440);
xor U3982 (N_3982,N_2736,N_2241);
xnor U3983 (N_3983,N_2959,N_2332);
or U3984 (N_3984,N_2155,N_2836);
nor U3985 (N_3985,N_2890,N_2500);
xnor U3986 (N_3986,N_2373,N_2821);
nand U3987 (N_3987,N_2990,N_2363);
nor U3988 (N_3988,N_2821,N_2601);
and U3989 (N_3989,N_2172,N_2005);
nor U3990 (N_3990,N_2446,N_2921);
and U3991 (N_3991,N_2248,N_2898);
nor U3992 (N_3992,N_2708,N_2329);
xor U3993 (N_3993,N_2469,N_2859);
xnor U3994 (N_3994,N_2781,N_2399);
nand U3995 (N_3995,N_2901,N_2006);
xor U3996 (N_3996,N_2289,N_2682);
xor U3997 (N_3997,N_2521,N_2682);
nand U3998 (N_3998,N_2208,N_2784);
xor U3999 (N_3999,N_2651,N_2557);
or U4000 (N_4000,N_3736,N_3624);
nor U4001 (N_4001,N_3269,N_3220);
or U4002 (N_4002,N_3536,N_3291);
or U4003 (N_4003,N_3766,N_3925);
xor U4004 (N_4004,N_3200,N_3371);
and U4005 (N_4005,N_3175,N_3859);
or U4006 (N_4006,N_3367,N_3613);
xor U4007 (N_4007,N_3442,N_3877);
and U4008 (N_4008,N_3718,N_3706);
xor U4009 (N_4009,N_3878,N_3399);
xor U4010 (N_4010,N_3654,N_3092);
or U4011 (N_4011,N_3252,N_3330);
or U4012 (N_4012,N_3166,N_3471);
nand U4013 (N_4013,N_3457,N_3641);
or U4014 (N_4014,N_3658,N_3637);
or U4015 (N_4015,N_3625,N_3904);
xnor U4016 (N_4016,N_3124,N_3229);
and U4017 (N_4017,N_3563,N_3807);
xnor U4018 (N_4018,N_3104,N_3984);
nor U4019 (N_4019,N_3545,N_3996);
nand U4020 (N_4020,N_3325,N_3599);
nor U4021 (N_4021,N_3887,N_3661);
or U4022 (N_4022,N_3967,N_3748);
nand U4023 (N_4023,N_3455,N_3403);
nor U4024 (N_4024,N_3711,N_3090);
xnor U4025 (N_4025,N_3049,N_3460);
or U4026 (N_4026,N_3633,N_3309);
or U4027 (N_4027,N_3667,N_3324);
or U4028 (N_4028,N_3136,N_3606);
or U4029 (N_4029,N_3825,N_3260);
nor U4030 (N_4030,N_3640,N_3814);
nor U4031 (N_4031,N_3816,N_3131);
and U4032 (N_4032,N_3621,N_3076);
xnor U4033 (N_4033,N_3946,N_3972);
nand U4034 (N_4034,N_3557,N_3231);
or U4035 (N_4035,N_3158,N_3970);
or U4036 (N_4036,N_3117,N_3644);
and U4037 (N_4037,N_3304,N_3138);
or U4038 (N_4038,N_3156,N_3547);
nor U4039 (N_4039,N_3401,N_3430);
or U4040 (N_4040,N_3947,N_3216);
and U4041 (N_4041,N_3580,N_3219);
and U4042 (N_4042,N_3337,N_3012);
xnor U4043 (N_4043,N_3931,N_3313);
xor U4044 (N_4044,N_3670,N_3833);
or U4045 (N_4045,N_3129,N_3505);
xor U4046 (N_4046,N_3973,N_3541);
xor U4047 (N_4047,N_3763,N_3623);
and U4048 (N_4048,N_3488,N_3635);
xor U4049 (N_4049,N_3015,N_3379);
nand U4050 (N_4050,N_3747,N_3162);
and U4051 (N_4051,N_3444,N_3465);
and U4052 (N_4052,N_3616,N_3643);
and U4053 (N_4053,N_3966,N_3802);
nor U4054 (N_4054,N_3798,N_3038);
nand U4055 (N_4055,N_3204,N_3426);
and U4056 (N_4056,N_3489,N_3879);
xnor U4057 (N_4057,N_3305,N_3612);
nor U4058 (N_4058,N_3757,N_3390);
nor U4059 (N_4059,N_3171,N_3868);
nor U4060 (N_4060,N_3112,N_3097);
and U4061 (N_4061,N_3762,N_3480);
xor U4062 (N_4062,N_3750,N_3163);
nand U4063 (N_4063,N_3466,N_3327);
nand U4064 (N_4064,N_3197,N_3082);
xor U4065 (N_4065,N_3537,N_3407);
and U4066 (N_4066,N_3133,N_3837);
and U4067 (N_4067,N_3772,N_3653);
and U4068 (N_4068,N_3053,N_3534);
and U4069 (N_4069,N_3700,N_3451);
xor U4070 (N_4070,N_3041,N_3533);
nand U4071 (N_4071,N_3923,N_3965);
and U4072 (N_4072,N_3227,N_3188);
nand U4073 (N_4073,N_3068,N_3607);
and U4074 (N_4074,N_3208,N_3276);
or U4075 (N_4075,N_3456,N_3414);
or U4076 (N_4076,N_3765,N_3713);
or U4077 (N_4077,N_3908,N_3777);
or U4078 (N_4078,N_3902,N_3919);
xnor U4079 (N_4079,N_3566,N_3727);
nand U4080 (N_4080,N_3067,N_3388);
and U4081 (N_4081,N_3650,N_3177);
or U4082 (N_4082,N_3195,N_3864);
and U4083 (N_4083,N_3699,N_3936);
xor U4084 (N_4084,N_3853,N_3093);
xor U4085 (N_4085,N_3478,N_3933);
xnor U4086 (N_4086,N_3334,N_3132);
nor U4087 (N_4087,N_3168,N_3590);
nor U4088 (N_4088,N_3027,N_3759);
nor U4089 (N_4089,N_3964,N_3627);
or U4090 (N_4090,N_3499,N_3732);
nor U4091 (N_4091,N_3078,N_3110);
nand U4092 (N_4092,N_3503,N_3292);
and U4093 (N_4093,N_3020,N_3105);
xnor U4094 (N_4094,N_3091,N_3826);
and U4095 (N_4095,N_3248,N_3823);
nor U4096 (N_4096,N_3400,N_3870);
nor U4097 (N_4097,N_3126,N_3761);
nor U4098 (N_4098,N_3062,N_3692);
nand U4099 (N_4099,N_3585,N_3361);
xnor U4100 (N_4100,N_3818,N_3949);
xnor U4101 (N_4101,N_3072,N_3472);
or U4102 (N_4102,N_3782,N_3137);
xor U4103 (N_4103,N_3708,N_3452);
nor U4104 (N_4104,N_3234,N_3264);
nand U4105 (N_4105,N_3036,N_3016);
nand U4106 (N_4106,N_3912,N_3787);
or U4107 (N_4107,N_3855,N_3061);
and U4108 (N_4108,N_3988,N_3368);
xor U4109 (N_4109,N_3120,N_3443);
xor U4110 (N_4110,N_3628,N_3075);
or U4111 (N_4111,N_3063,N_3495);
and U4112 (N_4112,N_3695,N_3603);
xor U4113 (N_4113,N_3697,N_3139);
and U4114 (N_4114,N_3882,N_3180);
or U4115 (N_4115,N_3303,N_3381);
or U4116 (N_4116,N_3207,N_3858);
nand U4117 (N_4117,N_3885,N_3588);
xnor U4118 (N_4118,N_3906,N_3098);
nor U4119 (N_4119,N_3159,N_3809);
and U4120 (N_4120,N_3555,N_3119);
and U4121 (N_4121,N_3290,N_3827);
nand U4122 (N_4122,N_3203,N_3352);
or U4123 (N_4123,N_3284,N_3948);
nor U4124 (N_4124,N_3316,N_3311);
and U4125 (N_4125,N_3006,N_3573);
xnor U4126 (N_4126,N_3420,N_3348);
nand U4127 (N_4127,N_3942,N_3866);
or U4128 (N_4128,N_3172,N_3510);
or U4129 (N_4129,N_3415,N_3295);
or U4130 (N_4130,N_3645,N_3889);
xor U4131 (N_4131,N_3312,N_3920);
nand U4132 (N_4132,N_3385,N_3358);
or U4133 (N_4133,N_3751,N_3449);
or U4134 (N_4134,N_3417,N_3184);
nand U4135 (N_4135,N_3294,N_3373);
nor U4136 (N_4136,N_3520,N_3301);
nand U4137 (N_4137,N_3134,N_3846);
nand U4138 (N_4138,N_3812,N_3228);
nand U4139 (N_4139,N_3940,N_3867);
nor U4140 (N_4140,N_3008,N_3490);
nand U4141 (N_4141,N_3926,N_3950);
or U4142 (N_4142,N_3094,N_3079);
or U4143 (N_4143,N_3578,N_3596);
nand U4144 (N_4144,N_3768,N_3000);
and U4145 (N_4145,N_3125,N_3341);
nor U4146 (N_4146,N_3386,N_3688);
nor U4147 (N_4147,N_3349,N_3754);
and U4148 (N_4148,N_3152,N_3551);
and U4149 (N_4149,N_3525,N_3854);
xor U4150 (N_4150,N_3107,N_3687);
or U4151 (N_4151,N_3981,N_3055);
nor U4152 (N_4152,N_3543,N_3485);
or U4153 (N_4153,N_3675,N_3800);
nand U4154 (N_4154,N_3085,N_3153);
or U4155 (N_4155,N_3225,N_3214);
nor U4156 (N_4156,N_3583,N_3288);
xnor U4157 (N_4157,N_3123,N_3318);
nor U4158 (N_4158,N_3860,N_3427);
or U4159 (N_4159,N_3416,N_3619);
nand U4160 (N_4160,N_3391,N_3895);
or U4161 (N_4161,N_3626,N_3888);
nand U4162 (N_4162,N_3293,N_3951);
xor U4163 (N_4163,N_3073,N_3458);
or U4164 (N_4164,N_3893,N_3486);
nor U4165 (N_4165,N_3238,N_3968);
nor U4166 (N_4166,N_3210,N_3002);
or U4167 (N_4167,N_3795,N_3561);
or U4168 (N_4168,N_3007,N_3307);
xnor U4169 (N_4169,N_3857,N_3283);
and U4170 (N_4170,N_3542,N_3767);
and U4171 (N_4171,N_3956,N_3605);
or U4172 (N_4172,N_3315,N_3657);
nor U4173 (N_4173,N_3514,N_3473);
or U4174 (N_4174,N_3775,N_3230);
and U4175 (N_4175,N_3587,N_3193);
nand U4176 (N_4176,N_3817,N_3360);
xor U4177 (N_4177,N_3672,N_3863);
xnor U4178 (N_4178,N_3102,N_3844);
nand U4179 (N_4179,N_3080,N_3211);
nand U4180 (N_4180,N_3709,N_3176);
and U4181 (N_4181,N_3577,N_3916);
nor U4182 (N_4182,N_3955,N_3004);
xor U4183 (N_4183,N_3862,N_3900);
xor U4184 (N_4184,N_3268,N_3232);
xnor U4185 (N_4185,N_3333,N_3244);
nand U4186 (N_4186,N_3069,N_3574);
nor U4187 (N_4187,N_3467,N_3716);
or U4188 (N_4188,N_3929,N_3508);
and U4189 (N_4189,N_3776,N_3087);
nand U4190 (N_4190,N_3247,N_3841);
xor U4191 (N_4191,N_3065,N_3831);
nand U4192 (N_4192,N_3764,N_3796);
nor U4193 (N_4193,N_3834,N_3589);
nand U4194 (N_4194,N_3610,N_3824);
or U4195 (N_4195,N_3187,N_3734);
nand U4196 (N_4196,N_3608,N_3310);
nor U4197 (N_4197,N_3298,N_3382);
nor U4198 (N_4198,N_3192,N_3639);
nor U4199 (N_4199,N_3261,N_3050);
and U4200 (N_4200,N_3045,N_3369);
or U4201 (N_4201,N_3468,N_3164);
and U4202 (N_4202,N_3898,N_3506);
and U4203 (N_4203,N_3969,N_3836);
nor U4204 (N_4204,N_3003,N_3629);
nor U4205 (N_4205,N_3032,N_3332);
nor U4206 (N_4206,N_3928,N_3521);
nand U4207 (N_4207,N_3081,N_3832);
or U4208 (N_4208,N_3493,N_3070);
nor U4209 (N_4209,N_3255,N_3202);
nor U4210 (N_4210,N_3249,N_3851);
and U4211 (N_4211,N_3986,N_3174);
nor U4212 (N_4212,N_3389,N_3372);
or U4213 (N_4213,N_3892,N_3236);
and U4214 (N_4214,N_3609,N_3270);
and U4215 (N_4215,N_3896,N_3448);
xor U4216 (N_4216,N_3218,N_3095);
nand U4217 (N_4217,N_3275,N_3453);
or U4218 (N_4218,N_3905,N_3022);
and U4219 (N_4219,N_3978,N_3285);
nand U4220 (N_4220,N_3845,N_3663);
and U4221 (N_4221,N_3582,N_3314);
and U4222 (N_4222,N_3549,N_3034);
xor U4223 (N_4223,N_3819,N_3057);
xnor U4224 (N_4224,N_3722,N_3331);
and U4225 (N_4225,N_3773,N_3861);
xnor U4226 (N_4226,N_3167,N_3839);
and U4227 (N_4227,N_3662,N_3890);
nand U4228 (N_4228,N_3149,N_3952);
or U4229 (N_4229,N_3556,N_3869);
xor U4230 (N_4230,N_3380,N_3976);
or U4231 (N_4231,N_3366,N_3299);
or U4232 (N_4232,N_3684,N_3704);
nand U4233 (N_4233,N_3350,N_3901);
xnor U4234 (N_4234,N_3475,N_3516);
and U4235 (N_4235,N_3852,N_3423);
or U4236 (N_4236,N_3393,N_3023);
xor U4237 (N_4237,N_3042,N_3962);
or U4238 (N_4238,N_3118,N_3433);
nand U4239 (N_4239,N_3226,N_3686);
xor U4240 (N_4240,N_3850,N_3335);
or U4241 (N_4241,N_3454,N_3529);
nand U4242 (N_4242,N_3685,N_3224);
and U4243 (N_4243,N_3028,N_3146);
nand U4244 (N_4244,N_3463,N_3733);
xnor U4245 (N_4245,N_3794,N_3838);
nand U4246 (N_4246,N_3037,N_3142);
nor U4247 (N_4247,N_3347,N_3266);
xor U4248 (N_4248,N_3482,N_3046);
and U4249 (N_4249,N_3274,N_3021);
xor U4250 (N_4250,N_3205,N_3954);
and U4251 (N_4251,N_3786,N_3918);
nand U4252 (N_4252,N_3494,N_3558);
or U4253 (N_4253,N_3982,N_3326);
nor U4254 (N_4254,N_3060,N_3096);
nand U4255 (N_4255,N_3913,N_3848);
xor U4256 (N_4256,N_3774,N_3646);
nor U4257 (N_4257,N_3677,N_3497);
or U4258 (N_4258,N_3921,N_3797);
or U4259 (N_4259,N_3805,N_3469);
and U4260 (N_4260,N_3029,N_3512);
nand U4261 (N_4261,N_3447,N_3601);
and U4262 (N_4262,N_3281,N_3539);
nand U4263 (N_4263,N_3030,N_3553);
xnor U4264 (N_4264,N_3048,N_3242);
nand U4265 (N_4265,N_3930,N_3530);
or U4266 (N_4266,N_3792,N_3598);
nor U4267 (N_4267,N_3944,N_3572);
and U4268 (N_4268,N_3217,N_3741);
xor U4269 (N_4269,N_3701,N_3440);
nor U4270 (N_4270,N_3277,N_3101);
nand U4271 (N_4271,N_3199,N_3883);
or U4272 (N_4272,N_3418,N_3527);
xnor U4273 (N_4273,N_3979,N_3263);
or U4274 (N_4274,N_3943,N_3279);
and U4275 (N_4275,N_3363,N_3945);
nand U4276 (N_4276,N_3740,N_3338);
and U4277 (N_4277,N_3784,N_3487);
or U4278 (N_4278,N_3491,N_3344);
and U4279 (N_4279,N_3297,N_3559);
xnor U4280 (N_4280,N_3398,N_3963);
and U4281 (N_4281,N_3799,N_3513);
nand U4282 (N_4282,N_3239,N_3903);
nand U4283 (N_4283,N_3779,N_3043);
xnor U4284 (N_4284,N_3265,N_3755);
and U4285 (N_4285,N_3111,N_3376);
xnor U4286 (N_4286,N_3121,N_3240);
xor U4287 (N_4287,N_3113,N_3743);
nor U4288 (N_4288,N_3682,N_3492);
nand U4289 (N_4289,N_3698,N_3346);
nand U4290 (N_4290,N_3907,N_3752);
nand U4291 (N_4291,N_3001,N_3911);
and U4292 (N_4292,N_3569,N_3144);
nor U4293 (N_4293,N_3383,N_3074);
or U4294 (N_4294,N_3614,N_3647);
xnor U4295 (N_4295,N_3822,N_3392);
nand U4296 (N_4296,N_3151,N_3434);
nand U4297 (N_4297,N_3351,N_3884);
xnor U4298 (N_4298,N_3189,N_3169);
and U4299 (N_4299,N_3897,N_3504);
nor U4300 (N_4300,N_3511,N_3375);
nand U4301 (N_4301,N_3507,N_3993);
xnor U4302 (N_4302,N_3329,N_3992);
and U4303 (N_4303,N_3665,N_3760);
xnor U4304 (N_4304,N_3995,N_3524);
nand U4305 (N_4305,N_3813,N_3746);
xnor U4306 (N_4306,N_3703,N_3025);
nor U4307 (N_4307,N_3742,N_3077);
xor U4308 (N_4308,N_3196,N_3179);
nor U4309 (N_4309,N_3306,N_3540);
and U4310 (N_4310,N_3791,N_3481);
xor U4311 (N_4311,N_3636,N_3106);
xor U4312 (N_4312,N_3615,N_3744);
xor U4313 (N_4313,N_3165,N_3222);
xor U4314 (N_4314,N_3419,N_3425);
nor U4315 (N_4315,N_3758,N_3509);
xor U4316 (N_4316,N_3690,N_3886);
nand U4317 (N_4317,N_3446,N_3632);
or U4318 (N_4318,N_3915,N_3876);
and U4319 (N_4319,N_3496,N_3059);
or U4320 (N_4320,N_3459,N_3723);
nor U4321 (N_4321,N_3031,N_3770);
or U4322 (N_4322,N_3961,N_3788);
nor U4323 (N_4323,N_3287,N_3241);
xor U4324 (N_4324,N_3396,N_3296);
xor U4325 (N_4325,N_3778,N_3130);
nand U4326 (N_4326,N_3565,N_3408);
and U4327 (N_4327,N_3983,N_3600);
nor U4328 (N_4328,N_3939,N_3450);
xnor U4329 (N_4329,N_3397,N_3273);
and U4330 (N_4330,N_3535,N_3847);
nor U4331 (N_4331,N_3980,N_3157);
nand U4332 (N_4332,N_3771,N_3322);
and U4333 (N_4333,N_3990,N_3522);
or U4334 (N_4334,N_3532,N_3689);
xor U4335 (N_4335,N_3694,N_3810);
nor U4336 (N_4336,N_3411,N_3568);
nand U4337 (N_4337,N_3808,N_3934);
nor U4338 (N_4338,N_3362,N_3567);
nor U4339 (N_4339,N_3710,N_3724);
xor U4340 (N_4340,N_3340,N_3725);
nor U4341 (N_4341,N_3317,N_3445);
and U4342 (N_4342,N_3715,N_3365);
nand U4343 (N_4343,N_3215,N_3576);
and U4344 (N_4344,N_3103,N_3738);
and U4345 (N_4345,N_3829,N_3147);
nand U4346 (N_4346,N_3739,N_3213);
nor U4347 (N_4347,N_3406,N_3395);
nor U4348 (N_4348,N_3441,N_3865);
nand U4349 (N_4349,N_3424,N_3871);
nor U4350 (N_4350,N_3470,N_3717);
xor U4351 (N_4351,N_3932,N_3570);
xnor U4352 (N_4352,N_3035,N_3251);
nand U4353 (N_4353,N_3575,N_3019);
nand U4354 (N_4354,N_3977,N_3518);
xnor U4355 (N_4355,N_3243,N_3611);
and U4356 (N_4356,N_3856,N_3116);
or U4357 (N_4357,N_3083,N_3975);
nand U4358 (N_4358,N_3122,N_3789);
nand U4359 (N_4359,N_3523,N_3250);
or U4360 (N_4360,N_3462,N_3483);
nor U4361 (N_4361,N_3874,N_3289);
xor U4362 (N_4362,N_3562,N_3412);
or U4363 (N_4363,N_3182,N_3484);
nor U4364 (N_4364,N_3413,N_3544);
xnor U4365 (N_4365,N_3880,N_3186);
nand U4366 (N_4366,N_3959,N_3498);
or U4367 (N_4367,N_3140,N_3378);
or U4368 (N_4368,N_3256,N_3278);
or U4369 (N_4369,N_3849,N_3707);
nor U4370 (N_4370,N_3464,N_3356);
and U4371 (N_4371,N_3668,N_3602);
nor U4372 (N_4372,N_3924,N_3502);
nor U4373 (N_4373,N_3353,N_3245);
or U4374 (N_4374,N_3084,N_3649);
or U4375 (N_4375,N_3128,N_3676);
xnor U4376 (N_4376,N_3592,N_3013);
and U4377 (N_4377,N_3927,N_3679);
nand U4378 (N_4378,N_3937,N_3875);
xnor U4379 (N_4379,N_3803,N_3246);
and U4380 (N_4380,N_3634,N_3815);
and U4381 (N_4381,N_3891,N_3622);
nand U4382 (N_4382,N_3579,N_3731);
nand U4383 (N_4383,N_3595,N_3233);
and U4384 (N_4384,N_3737,N_3018);
or U4385 (N_4385,N_3089,N_3552);
and U4386 (N_4386,N_3474,N_3958);
nand U4387 (N_4387,N_3678,N_3631);
nor U4388 (N_4388,N_3410,N_3801);
xnor U4389 (N_4389,N_3127,N_3476);
xnor U4390 (N_4390,N_3047,N_3781);
or U4391 (N_4391,N_3394,N_3143);
xor U4392 (N_4392,N_3058,N_3145);
nand U4393 (N_4393,N_3953,N_3756);
xor U4394 (N_4394,N_3014,N_3115);
nor U4395 (N_4395,N_3237,N_3033);
and U4396 (N_4396,N_3554,N_3660);
xor U4397 (N_4397,N_3223,N_3987);
nand U4398 (N_4398,N_3017,N_3336);
and U4399 (N_4399,N_3693,N_3384);
and U4400 (N_4400,N_3721,N_3370);
or U4401 (N_4401,N_3141,N_3749);
or U4402 (N_4402,N_3745,N_3461);
and U4403 (N_4403,N_3178,N_3160);
nand U4404 (N_4404,N_3064,N_3286);
nand U4405 (N_4405,N_3071,N_3840);
nand U4406 (N_4406,N_3364,N_3714);
and U4407 (N_4407,N_3664,N_3005);
or U4408 (N_4408,N_3438,N_3374);
and U4409 (N_4409,N_3343,N_3705);
and U4410 (N_4410,N_3319,N_3339);
and U4411 (N_4411,N_3806,N_3258);
xor U4412 (N_4412,N_3994,N_3431);
nor U4413 (N_4413,N_3730,N_3320);
or U4414 (N_4414,N_3999,N_3571);
xnor U4415 (N_4415,N_3357,N_3272);
nor U4416 (N_4416,N_3648,N_3100);
or U4417 (N_4417,N_3914,N_3282);
nor U4418 (N_4418,N_3432,N_3835);
xnor U4419 (N_4419,N_3935,N_3584);
nand U4420 (N_4420,N_3010,N_3894);
nand U4421 (N_4421,N_3719,N_3594);
nor U4422 (N_4422,N_3674,N_3617);
and U4423 (N_4423,N_3479,N_3769);
xor U4424 (N_4424,N_3656,N_3154);
nor U4425 (N_4425,N_3604,N_3780);
xor U4426 (N_4426,N_3652,N_3428);
nand U4427 (N_4427,N_3941,N_3683);
and U4428 (N_4428,N_3436,N_3024);
xor U4429 (N_4429,N_3011,N_3974);
nand U4430 (N_4430,N_3531,N_3191);
and U4431 (N_4431,N_3659,N_3728);
nand U4432 (N_4432,N_3729,N_3546);
nand U4433 (N_4433,N_3354,N_3785);
nor U4434 (N_4434,N_3691,N_3564);
and U4435 (N_4435,N_3429,N_3560);
xnor U4436 (N_4436,N_3991,N_3206);
nand U4437 (N_4437,N_3302,N_3387);
or U4438 (N_4438,N_3922,N_3828);
or U4439 (N_4439,N_3597,N_3783);
nand U4440 (N_4440,N_3026,N_3342);
and U4441 (N_4441,N_3066,N_3811);
and U4442 (N_4442,N_3404,N_3702);
and U4443 (N_4443,N_3235,N_3793);
or U4444 (N_4444,N_3439,N_3435);
or U4445 (N_4445,N_3681,N_3170);
nand U4446 (N_4446,N_3148,N_3402);
or U4447 (N_4447,N_3843,N_3842);
or U4448 (N_4448,N_3985,N_3044);
and U4449 (N_4449,N_3328,N_3620);
nand U4450 (N_4450,N_3056,N_3548);
or U4451 (N_4451,N_3183,N_3881);
nand U4452 (N_4452,N_3185,N_3262);
xor U4453 (N_4453,N_3910,N_3212);
nor U4454 (N_4454,N_3039,N_3150);
nor U4455 (N_4455,N_3308,N_3666);
or U4456 (N_4456,N_3528,N_3155);
or U4457 (N_4457,N_3593,N_3517);
nand U4458 (N_4458,N_3655,N_3321);
and U4459 (N_4459,N_3437,N_3550);
nand U4460 (N_4460,N_3267,N_3086);
xor U4461 (N_4461,N_3960,N_3052);
nor U4462 (N_4462,N_3581,N_3271);
xor U4463 (N_4463,N_3114,N_3917);
xor U4464 (N_4464,N_3345,N_3009);
xor U4465 (N_4465,N_3359,N_3198);
xor U4466 (N_4466,N_3753,N_3519);
nor U4467 (N_4467,N_3651,N_3194);
nor U4468 (N_4468,N_3804,N_3051);
or U4469 (N_4469,N_3161,N_3501);
nand U4470 (N_4470,N_3712,N_3221);
nand U4471 (N_4471,N_3173,N_3873);
and U4472 (N_4472,N_3630,N_3790);
or U4473 (N_4473,N_3673,N_3254);
nor U4474 (N_4474,N_3377,N_3591);
xor U4475 (N_4475,N_3209,N_3201);
and U4476 (N_4476,N_3642,N_3671);
and U4477 (N_4477,N_3421,N_3253);
xor U4478 (N_4478,N_3820,N_3526);
nand U4479 (N_4479,N_3355,N_3538);
nand U4480 (N_4480,N_3971,N_3821);
xor U4481 (N_4481,N_3181,N_3586);
xnor U4482 (N_4482,N_3109,N_3938);
and U4483 (N_4483,N_3909,N_3257);
and U4484 (N_4484,N_3088,N_3720);
and U4485 (N_4485,N_3997,N_3618);
or U4486 (N_4486,N_3696,N_3135);
xor U4487 (N_4487,N_3099,N_3872);
or U4488 (N_4488,N_3108,N_3280);
nand U4489 (N_4489,N_3957,N_3054);
nand U4490 (N_4490,N_3040,N_3409);
and U4491 (N_4491,N_3323,N_3680);
nor U4492 (N_4492,N_3989,N_3190);
and U4493 (N_4493,N_3899,N_3259);
or U4494 (N_4494,N_3735,N_3300);
or U4495 (N_4495,N_3726,N_3422);
xnor U4496 (N_4496,N_3405,N_3500);
and U4497 (N_4497,N_3669,N_3515);
nor U4498 (N_4498,N_3830,N_3998);
xor U4499 (N_4499,N_3477,N_3638);
nor U4500 (N_4500,N_3652,N_3681);
nand U4501 (N_4501,N_3860,N_3758);
or U4502 (N_4502,N_3741,N_3935);
nand U4503 (N_4503,N_3349,N_3416);
nor U4504 (N_4504,N_3899,N_3792);
or U4505 (N_4505,N_3697,N_3082);
nand U4506 (N_4506,N_3916,N_3284);
and U4507 (N_4507,N_3477,N_3835);
and U4508 (N_4508,N_3593,N_3198);
nor U4509 (N_4509,N_3364,N_3265);
and U4510 (N_4510,N_3767,N_3827);
nor U4511 (N_4511,N_3123,N_3976);
and U4512 (N_4512,N_3406,N_3002);
nor U4513 (N_4513,N_3979,N_3939);
or U4514 (N_4514,N_3552,N_3865);
or U4515 (N_4515,N_3669,N_3917);
nand U4516 (N_4516,N_3156,N_3502);
nand U4517 (N_4517,N_3967,N_3877);
xor U4518 (N_4518,N_3260,N_3933);
nor U4519 (N_4519,N_3606,N_3396);
xnor U4520 (N_4520,N_3905,N_3336);
and U4521 (N_4521,N_3634,N_3095);
and U4522 (N_4522,N_3031,N_3664);
or U4523 (N_4523,N_3267,N_3871);
or U4524 (N_4524,N_3231,N_3351);
and U4525 (N_4525,N_3723,N_3926);
and U4526 (N_4526,N_3012,N_3608);
nand U4527 (N_4527,N_3764,N_3855);
xnor U4528 (N_4528,N_3884,N_3625);
and U4529 (N_4529,N_3240,N_3905);
xor U4530 (N_4530,N_3648,N_3599);
nor U4531 (N_4531,N_3959,N_3243);
and U4532 (N_4532,N_3479,N_3816);
and U4533 (N_4533,N_3831,N_3215);
nor U4534 (N_4534,N_3840,N_3247);
nand U4535 (N_4535,N_3713,N_3414);
or U4536 (N_4536,N_3899,N_3132);
or U4537 (N_4537,N_3258,N_3073);
and U4538 (N_4538,N_3240,N_3442);
or U4539 (N_4539,N_3725,N_3064);
and U4540 (N_4540,N_3790,N_3874);
xnor U4541 (N_4541,N_3814,N_3534);
or U4542 (N_4542,N_3221,N_3361);
nor U4543 (N_4543,N_3129,N_3923);
or U4544 (N_4544,N_3488,N_3975);
nand U4545 (N_4545,N_3248,N_3608);
or U4546 (N_4546,N_3197,N_3440);
nor U4547 (N_4547,N_3002,N_3274);
and U4548 (N_4548,N_3977,N_3871);
xor U4549 (N_4549,N_3081,N_3148);
and U4550 (N_4550,N_3225,N_3688);
or U4551 (N_4551,N_3041,N_3261);
or U4552 (N_4552,N_3222,N_3042);
nand U4553 (N_4553,N_3412,N_3991);
nand U4554 (N_4554,N_3119,N_3462);
nand U4555 (N_4555,N_3137,N_3157);
nor U4556 (N_4556,N_3617,N_3910);
or U4557 (N_4557,N_3263,N_3864);
and U4558 (N_4558,N_3205,N_3881);
xor U4559 (N_4559,N_3337,N_3193);
xor U4560 (N_4560,N_3922,N_3723);
nand U4561 (N_4561,N_3384,N_3627);
xor U4562 (N_4562,N_3813,N_3395);
nor U4563 (N_4563,N_3358,N_3080);
nor U4564 (N_4564,N_3634,N_3390);
nand U4565 (N_4565,N_3252,N_3671);
xor U4566 (N_4566,N_3405,N_3545);
and U4567 (N_4567,N_3198,N_3314);
nor U4568 (N_4568,N_3698,N_3638);
and U4569 (N_4569,N_3785,N_3922);
and U4570 (N_4570,N_3759,N_3392);
and U4571 (N_4571,N_3969,N_3367);
and U4572 (N_4572,N_3071,N_3765);
xnor U4573 (N_4573,N_3306,N_3966);
nor U4574 (N_4574,N_3552,N_3152);
nand U4575 (N_4575,N_3340,N_3370);
xor U4576 (N_4576,N_3535,N_3956);
xor U4577 (N_4577,N_3670,N_3640);
nor U4578 (N_4578,N_3732,N_3899);
xnor U4579 (N_4579,N_3219,N_3780);
or U4580 (N_4580,N_3701,N_3064);
and U4581 (N_4581,N_3117,N_3418);
or U4582 (N_4582,N_3390,N_3326);
and U4583 (N_4583,N_3945,N_3456);
xnor U4584 (N_4584,N_3475,N_3217);
and U4585 (N_4585,N_3181,N_3304);
and U4586 (N_4586,N_3063,N_3416);
nor U4587 (N_4587,N_3252,N_3120);
nor U4588 (N_4588,N_3281,N_3639);
or U4589 (N_4589,N_3465,N_3675);
xor U4590 (N_4590,N_3109,N_3032);
xnor U4591 (N_4591,N_3411,N_3606);
nand U4592 (N_4592,N_3733,N_3359);
nor U4593 (N_4593,N_3584,N_3992);
or U4594 (N_4594,N_3686,N_3377);
xnor U4595 (N_4595,N_3840,N_3181);
or U4596 (N_4596,N_3069,N_3033);
xor U4597 (N_4597,N_3629,N_3242);
nand U4598 (N_4598,N_3242,N_3279);
nor U4599 (N_4599,N_3534,N_3392);
and U4600 (N_4600,N_3698,N_3538);
xnor U4601 (N_4601,N_3476,N_3417);
nor U4602 (N_4602,N_3170,N_3713);
xnor U4603 (N_4603,N_3309,N_3781);
or U4604 (N_4604,N_3269,N_3333);
xnor U4605 (N_4605,N_3418,N_3983);
and U4606 (N_4606,N_3516,N_3959);
and U4607 (N_4607,N_3761,N_3845);
nor U4608 (N_4608,N_3005,N_3522);
or U4609 (N_4609,N_3168,N_3767);
nand U4610 (N_4610,N_3308,N_3884);
xor U4611 (N_4611,N_3082,N_3260);
nand U4612 (N_4612,N_3530,N_3236);
and U4613 (N_4613,N_3411,N_3945);
or U4614 (N_4614,N_3576,N_3489);
xor U4615 (N_4615,N_3579,N_3614);
nand U4616 (N_4616,N_3668,N_3185);
or U4617 (N_4617,N_3569,N_3030);
xor U4618 (N_4618,N_3457,N_3420);
xnor U4619 (N_4619,N_3245,N_3205);
or U4620 (N_4620,N_3360,N_3322);
and U4621 (N_4621,N_3451,N_3744);
nor U4622 (N_4622,N_3684,N_3450);
and U4623 (N_4623,N_3604,N_3921);
nor U4624 (N_4624,N_3263,N_3240);
nand U4625 (N_4625,N_3463,N_3415);
nand U4626 (N_4626,N_3062,N_3480);
and U4627 (N_4627,N_3292,N_3374);
nor U4628 (N_4628,N_3425,N_3103);
and U4629 (N_4629,N_3069,N_3438);
or U4630 (N_4630,N_3314,N_3488);
nand U4631 (N_4631,N_3639,N_3165);
nand U4632 (N_4632,N_3892,N_3362);
xor U4633 (N_4633,N_3074,N_3862);
xnor U4634 (N_4634,N_3360,N_3884);
nor U4635 (N_4635,N_3009,N_3833);
xnor U4636 (N_4636,N_3701,N_3096);
xor U4637 (N_4637,N_3398,N_3318);
xnor U4638 (N_4638,N_3969,N_3789);
and U4639 (N_4639,N_3439,N_3064);
nand U4640 (N_4640,N_3051,N_3495);
and U4641 (N_4641,N_3739,N_3127);
nand U4642 (N_4642,N_3096,N_3619);
nor U4643 (N_4643,N_3683,N_3280);
xnor U4644 (N_4644,N_3713,N_3605);
xnor U4645 (N_4645,N_3881,N_3500);
xnor U4646 (N_4646,N_3855,N_3562);
and U4647 (N_4647,N_3216,N_3346);
xor U4648 (N_4648,N_3822,N_3848);
xor U4649 (N_4649,N_3040,N_3533);
and U4650 (N_4650,N_3253,N_3219);
xor U4651 (N_4651,N_3801,N_3224);
nor U4652 (N_4652,N_3066,N_3439);
or U4653 (N_4653,N_3879,N_3137);
xnor U4654 (N_4654,N_3045,N_3560);
or U4655 (N_4655,N_3213,N_3772);
nand U4656 (N_4656,N_3549,N_3272);
and U4657 (N_4657,N_3171,N_3639);
nand U4658 (N_4658,N_3040,N_3286);
or U4659 (N_4659,N_3161,N_3469);
nand U4660 (N_4660,N_3382,N_3497);
and U4661 (N_4661,N_3635,N_3001);
nor U4662 (N_4662,N_3773,N_3383);
nand U4663 (N_4663,N_3847,N_3578);
xor U4664 (N_4664,N_3401,N_3897);
nor U4665 (N_4665,N_3138,N_3201);
nor U4666 (N_4666,N_3345,N_3830);
xor U4667 (N_4667,N_3298,N_3561);
nand U4668 (N_4668,N_3933,N_3340);
or U4669 (N_4669,N_3900,N_3419);
nor U4670 (N_4670,N_3279,N_3726);
xnor U4671 (N_4671,N_3500,N_3089);
nand U4672 (N_4672,N_3383,N_3299);
xor U4673 (N_4673,N_3487,N_3133);
or U4674 (N_4674,N_3775,N_3251);
nor U4675 (N_4675,N_3751,N_3073);
and U4676 (N_4676,N_3472,N_3081);
xor U4677 (N_4677,N_3056,N_3070);
nand U4678 (N_4678,N_3681,N_3256);
and U4679 (N_4679,N_3505,N_3570);
and U4680 (N_4680,N_3046,N_3807);
nor U4681 (N_4681,N_3248,N_3717);
nand U4682 (N_4682,N_3859,N_3065);
nand U4683 (N_4683,N_3321,N_3714);
nand U4684 (N_4684,N_3571,N_3016);
or U4685 (N_4685,N_3170,N_3450);
and U4686 (N_4686,N_3876,N_3651);
xnor U4687 (N_4687,N_3815,N_3880);
xnor U4688 (N_4688,N_3669,N_3113);
and U4689 (N_4689,N_3858,N_3494);
nand U4690 (N_4690,N_3325,N_3484);
and U4691 (N_4691,N_3506,N_3955);
xnor U4692 (N_4692,N_3004,N_3079);
nand U4693 (N_4693,N_3472,N_3728);
or U4694 (N_4694,N_3226,N_3708);
nor U4695 (N_4695,N_3415,N_3640);
nand U4696 (N_4696,N_3293,N_3153);
or U4697 (N_4697,N_3651,N_3245);
xor U4698 (N_4698,N_3365,N_3661);
xor U4699 (N_4699,N_3708,N_3963);
xor U4700 (N_4700,N_3257,N_3036);
xor U4701 (N_4701,N_3669,N_3534);
and U4702 (N_4702,N_3943,N_3869);
nor U4703 (N_4703,N_3657,N_3691);
xnor U4704 (N_4704,N_3558,N_3730);
nand U4705 (N_4705,N_3190,N_3228);
or U4706 (N_4706,N_3359,N_3965);
or U4707 (N_4707,N_3128,N_3673);
nand U4708 (N_4708,N_3880,N_3837);
xnor U4709 (N_4709,N_3072,N_3134);
and U4710 (N_4710,N_3111,N_3959);
nor U4711 (N_4711,N_3565,N_3566);
and U4712 (N_4712,N_3264,N_3670);
nor U4713 (N_4713,N_3421,N_3891);
and U4714 (N_4714,N_3954,N_3862);
and U4715 (N_4715,N_3134,N_3551);
and U4716 (N_4716,N_3125,N_3637);
xor U4717 (N_4717,N_3738,N_3772);
nor U4718 (N_4718,N_3167,N_3423);
or U4719 (N_4719,N_3529,N_3007);
nand U4720 (N_4720,N_3783,N_3212);
and U4721 (N_4721,N_3663,N_3780);
and U4722 (N_4722,N_3379,N_3154);
and U4723 (N_4723,N_3941,N_3998);
nor U4724 (N_4724,N_3809,N_3978);
nand U4725 (N_4725,N_3940,N_3560);
or U4726 (N_4726,N_3508,N_3026);
xor U4727 (N_4727,N_3708,N_3308);
or U4728 (N_4728,N_3976,N_3825);
xor U4729 (N_4729,N_3346,N_3498);
xor U4730 (N_4730,N_3295,N_3981);
or U4731 (N_4731,N_3829,N_3660);
or U4732 (N_4732,N_3676,N_3207);
and U4733 (N_4733,N_3590,N_3238);
xnor U4734 (N_4734,N_3107,N_3225);
and U4735 (N_4735,N_3795,N_3374);
nand U4736 (N_4736,N_3998,N_3269);
nor U4737 (N_4737,N_3834,N_3647);
xnor U4738 (N_4738,N_3678,N_3400);
and U4739 (N_4739,N_3310,N_3759);
nand U4740 (N_4740,N_3392,N_3068);
and U4741 (N_4741,N_3264,N_3915);
nor U4742 (N_4742,N_3949,N_3331);
nand U4743 (N_4743,N_3556,N_3929);
or U4744 (N_4744,N_3875,N_3158);
xor U4745 (N_4745,N_3771,N_3890);
or U4746 (N_4746,N_3689,N_3490);
nor U4747 (N_4747,N_3553,N_3589);
xor U4748 (N_4748,N_3334,N_3583);
nand U4749 (N_4749,N_3087,N_3414);
nor U4750 (N_4750,N_3466,N_3356);
or U4751 (N_4751,N_3285,N_3386);
nor U4752 (N_4752,N_3284,N_3911);
nor U4753 (N_4753,N_3236,N_3599);
nand U4754 (N_4754,N_3518,N_3689);
nand U4755 (N_4755,N_3050,N_3444);
and U4756 (N_4756,N_3537,N_3711);
nor U4757 (N_4757,N_3111,N_3656);
xnor U4758 (N_4758,N_3991,N_3375);
and U4759 (N_4759,N_3525,N_3004);
nor U4760 (N_4760,N_3145,N_3358);
nor U4761 (N_4761,N_3033,N_3367);
and U4762 (N_4762,N_3437,N_3778);
xor U4763 (N_4763,N_3178,N_3356);
and U4764 (N_4764,N_3653,N_3841);
nor U4765 (N_4765,N_3506,N_3356);
nor U4766 (N_4766,N_3444,N_3775);
or U4767 (N_4767,N_3203,N_3538);
nor U4768 (N_4768,N_3259,N_3764);
and U4769 (N_4769,N_3479,N_3623);
xor U4770 (N_4770,N_3920,N_3051);
nor U4771 (N_4771,N_3363,N_3973);
or U4772 (N_4772,N_3616,N_3954);
nor U4773 (N_4773,N_3612,N_3694);
nand U4774 (N_4774,N_3852,N_3052);
nor U4775 (N_4775,N_3179,N_3297);
nor U4776 (N_4776,N_3791,N_3564);
xor U4777 (N_4777,N_3723,N_3181);
and U4778 (N_4778,N_3489,N_3325);
nand U4779 (N_4779,N_3567,N_3159);
or U4780 (N_4780,N_3578,N_3500);
nand U4781 (N_4781,N_3887,N_3979);
nor U4782 (N_4782,N_3813,N_3330);
nor U4783 (N_4783,N_3617,N_3366);
or U4784 (N_4784,N_3613,N_3283);
xor U4785 (N_4785,N_3711,N_3936);
and U4786 (N_4786,N_3030,N_3911);
or U4787 (N_4787,N_3917,N_3481);
and U4788 (N_4788,N_3859,N_3107);
xor U4789 (N_4789,N_3588,N_3330);
nand U4790 (N_4790,N_3893,N_3202);
or U4791 (N_4791,N_3921,N_3375);
or U4792 (N_4792,N_3061,N_3196);
xnor U4793 (N_4793,N_3013,N_3358);
nor U4794 (N_4794,N_3213,N_3468);
and U4795 (N_4795,N_3323,N_3785);
or U4796 (N_4796,N_3335,N_3938);
and U4797 (N_4797,N_3462,N_3737);
and U4798 (N_4798,N_3074,N_3412);
and U4799 (N_4799,N_3022,N_3964);
and U4800 (N_4800,N_3224,N_3175);
and U4801 (N_4801,N_3911,N_3472);
and U4802 (N_4802,N_3447,N_3675);
nand U4803 (N_4803,N_3316,N_3115);
or U4804 (N_4804,N_3741,N_3989);
or U4805 (N_4805,N_3953,N_3044);
or U4806 (N_4806,N_3166,N_3500);
xor U4807 (N_4807,N_3886,N_3590);
and U4808 (N_4808,N_3428,N_3233);
nand U4809 (N_4809,N_3827,N_3125);
nor U4810 (N_4810,N_3989,N_3732);
nand U4811 (N_4811,N_3401,N_3894);
or U4812 (N_4812,N_3247,N_3956);
nand U4813 (N_4813,N_3591,N_3358);
or U4814 (N_4814,N_3597,N_3382);
nor U4815 (N_4815,N_3995,N_3692);
or U4816 (N_4816,N_3459,N_3249);
or U4817 (N_4817,N_3875,N_3891);
nor U4818 (N_4818,N_3127,N_3384);
xor U4819 (N_4819,N_3286,N_3784);
nand U4820 (N_4820,N_3292,N_3069);
nand U4821 (N_4821,N_3963,N_3284);
nor U4822 (N_4822,N_3496,N_3263);
xor U4823 (N_4823,N_3428,N_3025);
or U4824 (N_4824,N_3991,N_3282);
nor U4825 (N_4825,N_3733,N_3123);
or U4826 (N_4826,N_3972,N_3004);
or U4827 (N_4827,N_3838,N_3783);
and U4828 (N_4828,N_3008,N_3062);
and U4829 (N_4829,N_3957,N_3824);
or U4830 (N_4830,N_3261,N_3202);
nand U4831 (N_4831,N_3491,N_3236);
or U4832 (N_4832,N_3846,N_3307);
and U4833 (N_4833,N_3711,N_3968);
nor U4834 (N_4834,N_3377,N_3019);
xor U4835 (N_4835,N_3361,N_3331);
nand U4836 (N_4836,N_3043,N_3517);
or U4837 (N_4837,N_3773,N_3778);
xor U4838 (N_4838,N_3565,N_3656);
or U4839 (N_4839,N_3366,N_3806);
nand U4840 (N_4840,N_3436,N_3168);
and U4841 (N_4841,N_3029,N_3941);
nand U4842 (N_4842,N_3261,N_3721);
nand U4843 (N_4843,N_3369,N_3804);
nand U4844 (N_4844,N_3432,N_3109);
xor U4845 (N_4845,N_3576,N_3342);
xnor U4846 (N_4846,N_3598,N_3799);
nand U4847 (N_4847,N_3220,N_3243);
and U4848 (N_4848,N_3670,N_3154);
nor U4849 (N_4849,N_3616,N_3944);
nand U4850 (N_4850,N_3745,N_3993);
nand U4851 (N_4851,N_3807,N_3164);
and U4852 (N_4852,N_3163,N_3730);
nor U4853 (N_4853,N_3224,N_3566);
xnor U4854 (N_4854,N_3860,N_3673);
xnor U4855 (N_4855,N_3891,N_3537);
nand U4856 (N_4856,N_3295,N_3386);
and U4857 (N_4857,N_3805,N_3571);
xor U4858 (N_4858,N_3762,N_3564);
and U4859 (N_4859,N_3421,N_3047);
nand U4860 (N_4860,N_3916,N_3275);
nor U4861 (N_4861,N_3100,N_3828);
and U4862 (N_4862,N_3134,N_3014);
and U4863 (N_4863,N_3796,N_3157);
or U4864 (N_4864,N_3847,N_3692);
xor U4865 (N_4865,N_3588,N_3268);
nand U4866 (N_4866,N_3678,N_3188);
nor U4867 (N_4867,N_3045,N_3471);
nor U4868 (N_4868,N_3719,N_3290);
or U4869 (N_4869,N_3999,N_3415);
xnor U4870 (N_4870,N_3682,N_3874);
or U4871 (N_4871,N_3724,N_3955);
or U4872 (N_4872,N_3840,N_3046);
or U4873 (N_4873,N_3555,N_3403);
nand U4874 (N_4874,N_3920,N_3903);
xor U4875 (N_4875,N_3632,N_3013);
and U4876 (N_4876,N_3409,N_3319);
xnor U4877 (N_4877,N_3232,N_3736);
nor U4878 (N_4878,N_3155,N_3870);
nand U4879 (N_4879,N_3979,N_3999);
and U4880 (N_4880,N_3363,N_3836);
and U4881 (N_4881,N_3157,N_3724);
and U4882 (N_4882,N_3279,N_3618);
or U4883 (N_4883,N_3277,N_3547);
xnor U4884 (N_4884,N_3501,N_3655);
and U4885 (N_4885,N_3344,N_3183);
xor U4886 (N_4886,N_3779,N_3755);
nand U4887 (N_4887,N_3737,N_3187);
xor U4888 (N_4888,N_3477,N_3259);
nand U4889 (N_4889,N_3350,N_3542);
nor U4890 (N_4890,N_3221,N_3904);
nor U4891 (N_4891,N_3331,N_3509);
or U4892 (N_4892,N_3292,N_3482);
nand U4893 (N_4893,N_3625,N_3310);
or U4894 (N_4894,N_3187,N_3822);
and U4895 (N_4895,N_3001,N_3049);
xor U4896 (N_4896,N_3355,N_3141);
xor U4897 (N_4897,N_3897,N_3475);
and U4898 (N_4898,N_3295,N_3911);
or U4899 (N_4899,N_3915,N_3974);
nor U4900 (N_4900,N_3119,N_3305);
xor U4901 (N_4901,N_3109,N_3589);
nor U4902 (N_4902,N_3613,N_3662);
xnor U4903 (N_4903,N_3547,N_3180);
and U4904 (N_4904,N_3089,N_3562);
nand U4905 (N_4905,N_3126,N_3259);
nand U4906 (N_4906,N_3952,N_3621);
xnor U4907 (N_4907,N_3792,N_3061);
nand U4908 (N_4908,N_3248,N_3189);
xor U4909 (N_4909,N_3498,N_3641);
xor U4910 (N_4910,N_3867,N_3241);
nor U4911 (N_4911,N_3388,N_3246);
or U4912 (N_4912,N_3570,N_3884);
and U4913 (N_4913,N_3098,N_3072);
nand U4914 (N_4914,N_3657,N_3293);
and U4915 (N_4915,N_3669,N_3617);
or U4916 (N_4916,N_3065,N_3708);
nor U4917 (N_4917,N_3513,N_3740);
xnor U4918 (N_4918,N_3711,N_3469);
xnor U4919 (N_4919,N_3861,N_3158);
or U4920 (N_4920,N_3354,N_3860);
and U4921 (N_4921,N_3801,N_3701);
or U4922 (N_4922,N_3259,N_3359);
or U4923 (N_4923,N_3555,N_3998);
or U4924 (N_4924,N_3565,N_3741);
nor U4925 (N_4925,N_3019,N_3847);
nand U4926 (N_4926,N_3807,N_3223);
and U4927 (N_4927,N_3692,N_3967);
or U4928 (N_4928,N_3986,N_3948);
nor U4929 (N_4929,N_3552,N_3088);
or U4930 (N_4930,N_3640,N_3560);
and U4931 (N_4931,N_3333,N_3883);
xor U4932 (N_4932,N_3251,N_3708);
and U4933 (N_4933,N_3711,N_3712);
nor U4934 (N_4934,N_3197,N_3000);
and U4935 (N_4935,N_3438,N_3389);
nand U4936 (N_4936,N_3457,N_3403);
nand U4937 (N_4937,N_3422,N_3064);
or U4938 (N_4938,N_3483,N_3688);
nand U4939 (N_4939,N_3732,N_3992);
nand U4940 (N_4940,N_3347,N_3471);
xnor U4941 (N_4941,N_3722,N_3059);
xor U4942 (N_4942,N_3862,N_3026);
and U4943 (N_4943,N_3972,N_3305);
xor U4944 (N_4944,N_3121,N_3653);
nor U4945 (N_4945,N_3589,N_3681);
xnor U4946 (N_4946,N_3174,N_3947);
xnor U4947 (N_4947,N_3834,N_3013);
xnor U4948 (N_4948,N_3239,N_3342);
nor U4949 (N_4949,N_3582,N_3256);
nor U4950 (N_4950,N_3216,N_3224);
nand U4951 (N_4951,N_3383,N_3508);
xor U4952 (N_4952,N_3716,N_3091);
nand U4953 (N_4953,N_3922,N_3370);
and U4954 (N_4954,N_3638,N_3586);
nand U4955 (N_4955,N_3035,N_3187);
nor U4956 (N_4956,N_3998,N_3038);
nand U4957 (N_4957,N_3332,N_3711);
xnor U4958 (N_4958,N_3881,N_3970);
nand U4959 (N_4959,N_3519,N_3624);
and U4960 (N_4960,N_3941,N_3024);
nand U4961 (N_4961,N_3323,N_3755);
nand U4962 (N_4962,N_3632,N_3656);
nor U4963 (N_4963,N_3957,N_3844);
nor U4964 (N_4964,N_3534,N_3609);
or U4965 (N_4965,N_3706,N_3185);
and U4966 (N_4966,N_3377,N_3127);
or U4967 (N_4967,N_3682,N_3653);
nor U4968 (N_4968,N_3934,N_3702);
xor U4969 (N_4969,N_3435,N_3855);
and U4970 (N_4970,N_3794,N_3955);
or U4971 (N_4971,N_3720,N_3923);
nor U4972 (N_4972,N_3331,N_3470);
nand U4973 (N_4973,N_3703,N_3224);
xor U4974 (N_4974,N_3610,N_3442);
xnor U4975 (N_4975,N_3597,N_3983);
or U4976 (N_4976,N_3076,N_3833);
nand U4977 (N_4977,N_3090,N_3835);
xnor U4978 (N_4978,N_3127,N_3314);
and U4979 (N_4979,N_3887,N_3022);
nor U4980 (N_4980,N_3783,N_3087);
or U4981 (N_4981,N_3415,N_3933);
nand U4982 (N_4982,N_3567,N_3186);
nand U4983 (N_4983,N_3211,N_3893);
nand U4984 (N_4984,N_3833,N_3139);
nor U4985 (N_4985,N_3969,N_3349);
or U4986 (N_4986,N_3434,N_3803);
nand U4987 (N_4987,N_3747,N_3968);
and U4988 (N_4988,N_3110,N_3910);
nand U4989 (N_4989,N_3080,N_3981);
nand U4990 (N_4990,N_3602,N_3598);
xor U4991 (N_4991,N_3272,N_3553);
xnor U4992 (N_4992,N_3745,N_3727);
and U4993 (N_4993,N_3628,N_3744);
xor U4994 (N_4994,N_3216,N_3761);
and U4995 (N_4995,N_3952,N_3080);
nor U4996 (N_4996,N_3019,N_3425);
nor U4997 (N_4997,N_3765,N_3804);
nor U4998 (N_4998,N_3198,N_3439);
and U4999 (N_4999,N_3855,N_3867);
or U5000 (N_5000,N_4912,N_4642);
xor U5001 (N_5001,N_4921,N_4805);
nand U5002 (N_5002,N_4398,N_4858);
nor U5003 (N_5003,N_4677,N_4511);
and U5004 (N_5004,N_4877,N_4565);
nand U5005 (N_5005,N_4338,N_4980);
and U5006 (N_5006,N_4420,N_4992);
xor U5007 (N_5007,N_4947,N_4527);
xor U5008 (N_5008,N_4055,N_4209);
xnor U5009 (N_5009,N_4036,N_4530);
or U5010 (N_5010,N_4926,N_4697);
nand U5011 (N_5011,N_4984,N_4014);
nand U5012 (N_5012,N_4415,N_4216);
and U5013 (N_5013,N_4798,N_4396);
xnor U5014 (N_5014,N_4377,N_4583);
xnor U5015 (N_5015,N_4199,N_4414);
or U5016 (N_5016,N_4599,N_4273);
or U5017 (N_5017,N_4234,N_4624);
nand U5018 (N_5018,N_4088,N_4572);
nor U5019 (N_5019,N_4295,N_4245);
or U5020 (N_5020,N_4728,N_4436);
nor U5021 (N_5021,N_4140,N_4372);
and U5022 (N_5022,N_4821,N_4491);
and U5023 (N_5023,N_4861,N_4819);
and U5024 (N_5024,N_4863,N_4483);
xnor U5025 (N_5025,N_4945,N_4767);
xor U5026 (N_5026,N_4561,N_4291);
or U5027 (N_5027,N_4710,N_4651);
nor U5028 (N_5028,N_4343,N_4161);
or U5029 (N_5029,N_4658,N_4669);
nor U5030 (N_5030,N_4843,N_4429);
nor U5031 (N_5031,N_4461,N_4387);
xor U5032 (N_5032,N_4688,N_4875);
nand U5033 (N_5033,N_4185,N_4846);
nand U5034 (N_5034,N_4737,N_4938);
nand U5035 (N_5035,N_4001,N_4519);
nand U5036 (N_5036,N_4477,N_4862);
nand U5037 (N_5037,N_4891,N_4366);
or U5038 (N_5038,N_4487,N_4760);
and U5039 (N_5039,N_4340,N_4730);
nand U5040 (N_5040,N_4474,N_4052);
nor U5041 (N_5041,N_4000,N_4750);
nor U5042 (N_5042,N_4460,N_4198);
or U5043 (N_5043,N_4820,N_4557);
and U5044 (N_5044,N_4870,N_4871);
nand U5045 (N_5045,N_4632,N_4224);
nor U5046 (N_5046,N_4687,N_4242);
and U5047 (N_5047,N_4418,N_4584);
nand U5048 (N_5048,N_4588,N_4543);
nor U5049 (N_5049,N_4319,N_4446);
nand U5050 (N_5050,N_4904,N_4153);
and U5051 (N_5051,N_4453,N_4038);
nor U5052 (N_5052,N_4508,N_4142);
and U5053 (N_5053,N_4410,N_4131);
and U5054 (N_5054,N_4620,N_4365);
xnor U5055 (N_5055,N_4797,N_4422);
nand U5056 (N_5056,N_4942,N_4794);
nor U5057 (N_5057,N_4850,N_4785);
and U5058 (N_5058,N_4804,N_4423);
and U5059 (N_5059,N_4200,N_4178);
or U5060 (N_5060,N_4930,N_4212);
nand U5061 (N_5061,N_4815,N_4704);
xnor U5062 (N_5062,N_4556,N_4791);
xor U5063 (N_5063,N_4262,N_4759);
nor U5064 (N_5064,N_4893,N_4496);
xor U5065 (N_5065,N_4364,N_4276);
nor U5066 (N_5066,N_4322,N_4480);
nor U5067 (N_5067,N_4093,N_4272);
or U5068 (N_5068,N_4520,N_4268);
nor U5069 (N_5069,N_4486,N_4296);
and U5070 (N_5070,N_4681,N_4678);
and U5071 (N_5071,N_4576,N_4983);
xor U5072 (N_5072,N_4439,N_4581);
and U5073 (N_5073,N_4179,N_4533);
xor U5074 (N_5074,N_4702,N_4978);
nor U5075 (N_5075,N_4154,N_4176);
nor U5076 (N_5076,N_4167,N_4975);
nand U5077 (N_5077,N_4267,N_4368);
and U5078 (N_5078,N_4585,N_4650);
nor U5079 (N_5079,N_4700,N_4493);
or U5080 (N_5080,N_4362,N_4716);
and U5081 (N_5081,N_4484,N_4866);
or U5082 (N_5082,N_4551,N_4749);
nor U5083 (N_5083,N_4416,N_4577);
nand U5084 (N_5084,N_4600,N_4696);
xnor U5085 (N_5085,N_4878,N_4417);
xnor U5086 (N_5086,N_4253,N_4649);
xnor U5087 (N_5087,N_4127,N_4129);
nand U5088 (N_5088,N_4977,N_4671);
nor U5089 (N_5089,N_4160,N_4255);
nand U5090 (N_5090,N_4189,N_4770);
xor U5091 (N_5091,N_4099,N_4067);
nand U5092 (N_5092,N_4044,N_4316);
nand U5093 (N_5093,N_4685,N_4727);
or U5094 (N_5094,N_4072,N_4703);
xor U5095 (N_5095,N_4633,N_4996);
nand U5096 (N_5096,N_4636,N_4569);
and U5097 (N_5097,N_4249,N_4523);
or U5098 (N_5098,N_4333,N_4943);
nand U5099 (N_5099,N_4999,N_4317);
xor U5100 (N_5100,N_4337,N_4313);
or U5101 (N_5101,N_4449,N_4196);
nand U5102 (N_5102,N_4789,N_4330);
or U5103 (N_5103,N_4083,N_4327);
xor U5104 (N_5104,N_4995,N_4358);
nor U5105 (N_5105,N_4973,N_4673);
xnor U5106 (N_5106,N_4241,N_4121);
nor U5107 (N_5107,N_4307,N_4957);
nor U5108 (N_5108,N_4353,N_4321);
nand U5109 (N_5109,N_4469,N_4745);
xor U5110 (N_5110,N_4345,N_4932);
nand U5111 (N_5111,N_4318,N_4148);
nor U5112 (N_5112,N_4645,N_4492);
and U5113 (N_5113,N_4908,N_4568);
nand U5114 (N_5114,N_4868,N_4187);
nand U5115 (N_5115,N_4689,N_4521);
xor U5116 (N_5116,N_4788,N_4763);
and U5117 (N_5117,N_4007,N_4331);
or U5118 (N_5118,N_4990,N_4674);
nand U5119 (N_5119,N_4857,N_4481);
nand U5120 (N_5120,N_4409,N_4698);
xor U5121 (N_5121,N_4352,N_4374);
nand U5122 (N_5122,N_4434,N_4931);
nand U5123 (N_5123,N_4030,N_4540);
nor U5124 (N_5124,N_4529,N_4679);
xnor U5125 (N_5125,N_4611,N_4715);
and U5126 (N_5126,N_4801,N_4652);
or U5127 (N_5127,N_4748,N_4133);
xnor U5128 (N_5128,N_4190,N_4013);
or U5129 (N_5129,N_4656,N_4287);
or U5130 (N_5130,N_4304,N_4100);
xor U5131 (N_5131,N_4281,N_4472);
or U5132 (N_5132,N_4828,N_4888);
xor U5133 (N_5133,N_4752,N_4940);
and U5134 (N_5134,N_4717,N_4170);
or U5135 (N_5135,N_4003,N_4357);
xor U5136 (N_5136,N_4388,N_4617);
and U5137 (N_5137,N_4810,N_4336);
nand U5138 (N_5138,N_4049,N_4243);
xor U5139 (N_5139,N_4927,N_4751);
nor U5140 (N_5140,N_4504,N_4407);
xnor U5141 (N_5141,N_4068,N_4714);
nand U5142 (N_5142,N_4740,N_4334);
or U5143 (N_5143,N_4676,N_4690);
xnor U5144 (N_5144,N_4818,N_4342);
nand U5145 (N_5145,N_4854,N_4265);
or U5146 (N_5146,N_4614,N_4762);
xnor U5147 (N_5147,N_4787,N_4571);
nand U5148 (N_5148,N_4310,N_4256);
and U5149 (N_5149,N_4860,N_4553);
and U5150 (N_5150,N_4430,N_4563);
and U5151 (N_5151,N_4378,N_4077);
nor U5152 (N_5152,N_4792,N_4950);
or U5153 (N_5153,N_4254,N_4096);
and U5154 (N_5154,N_4666,N_4827);
xor U5155 (N_5155,N_4668,N_4183);
nor U5156 (N_5156,N_4916,N_4811);
and U5157 (N_5157,N_4482,N_4227);
xnor U5158 (N_5158,N_4694,N_4974);
xor U5159 (N_5159,N_4203,N_4963);
or U5160 (N_5160,N_4528,N_4896);
or U5161 (N_5161,N_4367,N_4117);
and U5162 (N_5162,N_4552,N_4193);
nor U5163 (N_5163,N_4402,N_4479);
or U5164 (N_5164,N_4900,N_4173);
xnor U5165 (N_5165,N_4073,N_4107);
nand U5166 (N_5166,N_4080,N_4181);
xnor U5167 (N_5167,N_4314,N_4286);
or U5168 (N_5168,N_4873,N_4741);
and U5169 (N_5169,N_4166,N_4123);
and U5170 (N_5170,N_4831,N_4005);
nand U5171 (N_5171,N_4675,N_4596);
xor U5172 (N_5172,N_4539,N_4512);
nand U5173 (N_5173,N_4084,N_4053);
nand U5174 (N_5174,N_4898,N_4555);
nand U5175 (N_5175,N_4793,N_4376);
nor U5176 (N_5176,N_4274,N_4293);
and U5177 (N_5177,N_4011,N_4969);
and U5178 (N_5178,N_4644,N_4817);
and U5179 (N_5179,N_4610,N_4665);
xor U5180 (N_5180,N_4634,N_4455);
and U5181 (N_5181,N_4731,N_4693);
or U5182 (N_5182,N_4948,N_4278);
nor U5183 (N_5183,N_4116,N_4894);
xnor U5184 (N_5184,N_4701,N_4802);
xor U5185 (N_5185,N_4606,N_4790);
nor U5186 (N_5186,N_4803,N_4746);
or U5187 (N_5187,N_4724,N_4708);
and U5188 (N_5188,N_4747,N_4421);
or U5189 (N_5189,N_4324,N_4152);
nand U5190 (N_5190,N_4282,N_4922);
nand U5191 (N_5191,N_4607,N_4426);
and U5192 (N_5192,N_4468,N_4550);
nor U5193 (N_5193,N_4734,N_4413);
nand U5194 (N_5194,N_4777,N_4385);
and U5195 (N_5195,N_4782,N_4059);
or U5196 (N_5196,N_4027,N_4126);
and U5197 (N_5197,N_4609,N_4438);
nand U5198 (N_5198,N_4039,N_4350);
or U5199 (N_5199,N_4876,N_4020);
and U5200 (N_5200,N_4910,N_4134);
xnor U5201 (N_5201,N_4051,N_4213);
and U5202 (N_5202,N_4018,N_4769);
or U5203 (N_5203,N_4047,N_4269);
nor U5204 (N_5204,N_4458,N_4886);
nor U5205 (N_5205,N_4756,N_4298);
and U5206 (N_5206,N_4391,N_4294);
nand U5207 (N_5207,N_4229,N_4641);
or U5208 (N_5208,N_4643,N_4952);
and U5209 (N_5209,N_4814,N_4498);
nand U5210 (N_5210,N_4667,N_4002);
nor U5211 (N_5211,N_4879,N_4139);
and U5212 (N_5212,N_4598,N_4622);
nor U5213 (N_5213,N_4538,N_4202);
and U5214 (N_5214,N_4911,N_4816);
and U5215 (N_5215,N_4869,N_4435);
nor U5216 (N_5216,N_4949,N_4408);
and U5217 (N_5217,N_4120,N_4541);
nand U5218 (N_5218,N_4411,N_4381);
or U5219 (N_5219,N_4574,N_4718);
nand U5220 (N_5220,N_4783,N_4774);
or U5221 (N_5221,N_4115,N_4210);
or U5222 (N_5222,N_4288,N_4355);
or U5223 (N_5223,N_4230,N_4799);
nor U5224 (N_5224,N_4883,N_4069);
nor U5225 (N_5225,N_4686,N_4145);
nor U5226 (N_5226,N_4284,N_4394);
and U5227 (N_5227,N_4976,N_4061);
and U5228 (N_5228,N_4987,N_4156);
nor U5229 (N_5229,N_4165,N_4988);
xor U5230 (N_5230,N_4063,N_4035);
nor U5231 (N_5231,N_4755,N_4285);
or U5232 (N_5232,N_4251,N_4591);
xor U5233 (N_5233,N_4711,N_4619);
and U5234 (N_5234,N_4595,N_4844);
xnor U5235 (N_5235,N_4300,N_4305);
and U5236 (N_5236,N_4211,N_4761);
nor U5237 (N_5237,N_4989,N_4302);
or U5238 (N_5238,N_4829,N_4909);
or U5239 (N_5239,N_4220,N_4043);
nand U5240 (N_5240,N_4872,N_4264);
xor U5241 (N_5241,N_4114,N_4029);
nor U5242 (N_5242,N_4386,N_4847);
or U5243 (N_5243,N_4851,N_4075);
and U5244 (N_5244,N_4464,N_4985);
and U5245 (N_5245,N_4659,N_4205);
xor U5246 (N_5246,N_4354,N_4328);
nor U5247 (N_5247,N_4695,N_4040);
and U5248 (N_5248,N_4625,N_4979);
xnor U5249 (N_5249,N_4079,N_4935);
or U5250 (N_5250,N_4548,N_4822);
and U5251 (N_5251,N_4524,N_4841);
or U5252 (N_5252,N_4473,N_4054);
nor U5253 (N_5253,N_4986,N_4899);
nor U5254 (N_5254,N_4968,N_4476);
or U5255 (N_5255,N_4019,N_4110);
nor U5256 (N_5256,N_4004,N_4800);
and U5257 (N_5257,N_4323,N_4532);
or U5258 (N_5258,N_4138,N_4758);
xor U5259 (N_5259,N_4779,N_4171);
and U5260 (N_5260,N_4629,N_4006);
xnor U5261 (N_5261,N_4235,N_4885);
nand U5262 (N_5262,N_4301,N_4683);
nand U5263 (N_5263,N_4808,N_4903);
nand U5264 (N_5264,N_4918,N_4144);
xnor U5265 (N_5265,N_4733,N_4954);
and U5266 (N_5266,N_4082,N_4008);
xnor U5267 (N_5267,N_4346,N_4297);
or U5268 (N_5268,N_4309,N_4959);
xor U5269 (N_5269,N_4720,N_4849);
or U5270 (N_5270,N_4608,N_4425);
or U5271 (N_5271,N_4776,N_4128);
or U5272 (N_5272,N_4118,N_4451);
nor U5273 (N_5273,N_4603,N_4231);
nor U5274 (N_5274,N_4654,N_4501);
or U5275 (N_5275,N_4403,N_4105);
nand U5276 (N_5276,N_4500,N_4208);
and U5277 (N_5277,N_4824,N_4907);
and U5278 (N_5278,N_4856,N_4375);
or U5279 (N_5279,N_4605,N_4631);
or U5280 (N_5280,N_4852,N_4646);
and U5281 (N_5281,N_4807,N_4855);
and U5282 (N_5282,N_4955,N_4754);
xor U5283 (N_5283,N_4141,N_4835);
or U5284 (N_5284,N_4806,N_4657);
and U5285 (N_5285,N_4325,N_4025);
and U5286 (N_5286,N_4450,N_4085);
and U5287 (N_5287,N_4428,N_4045);
and U5288 (N_5288,N_4191,N_4292);
nand U5289 (N_5289,N_4956,N_4401);
nand U5290 (N_5290,N_4764,N_4465);
and U5291 (N_5291,N_4757,N_4503);
nand U5292 (N_5292,N_4567,N_4326);
or U5293 (N_5293,N_4914,N_4137);
xor U5294 (N_5294,N_4444,N_4440);
nand U5295 (N_5295,N_4640,N_4157);
or U5296 (N_5296,N_4470,N_4339);
and U5297 (N_5297,N_4923,N_4537);
nor U5298 (N_5298,N_4261,N_4149);
and U5299 (N_5299,N_4399,N_4159);
and U5300 (N_5300,N_4119,N_4536);
or U5301 (N_5301,N_4997,N_4594);
or U5302 (N_5302,N_4602,N_4880);
nand U5303 (N_5303,N_4023,N_4525);
and U5304 (N_5304,N_4928,N_4825);
xnor U5305 (N_5305,N_4832,N_4601);
nor U5306 (N_5306,N_4478,N_4662);
nor U5307 (N_5307,N_4887,N_4104);
or U5308 (N_5308,N_4592,N_4065);
and U5309 (N_5309,N_4913,N_4382);
or U5310 (N_5310,N_4351,N_4076);
or U5311 (N_5311,N_4545,N_4034);
xor U5312 (N_5312,N_4012,N_4897);
and U5313 (N_5313,N_4106,N_4534);
xor U5314 (N_5314,N_4933,N_4682);
xor U5315 (N_5315,N_4448,N_4299);
nor U5316 (N_5316,N_4623,N_4041);
xnor U5317 (N_5317,N_4130,N_4225);
and U5318 (N_5318,N_4062,N_4312);
nand U5319 (N_5319,N_4016,N_4499);
nor U5320 (N_5320,N_4960,N_4612);
nor U5321 (N_5321,N_4266,N_4833);
or U5322 (N_5322,N_4217,N_4834);
or U5323 (N_5323,N_4823,N_4573);
and U5324 (N_5324,N_4586,N_4842);
nand U5325 (N_5325,N_4672,N_4735);
or U5326 (N_5326,N_4188,N_4197);
nor U5327 (N_5327,N_4162,N_4837);
nor U5328 (N_5328,N_4836,N_4447);
or U5329 (N_5329,N_4158,N_4958);
nand U5330 (N_5330,N_4587,N_4889);
nor U5331 (N_5331,N_4826,N_4260);
nand U5332 (N_5332,N_4713,N_4699);
or U5333 (N_5333,N_4582,N_4795);
and U5334 (N_5334,N_4946,N_4929);
nor U5335 (N_5335,N_4580,N_4456);
nor U5336 (N_5336,N_4086,N_4445);
xor U5337 (N_5337,N_4575,N_4400);
or U5338 (N_5338,N_4739,N_4919);
and U5339 (N_5339,N_4172,N_4057);
and U5340 (N_5340,N_4744,N_4966);
xnor U5341 (N_5341,N_4169,N_4736);
or U5342 (N_5342,N_4902,N_4369);
nor U5343 (N_5343,N_4432,N_4991);
and U5344 (N_5344,N_4442,N_4066);
and U5345 (N_5345,N_4882,N_4344);
nand U5346 (N_5346,N_4661,N_4743);
and U5347 (N_5347,N_4604,N_4962);
nor U5348 (N_5348,N_4627,N_4441);
and U5349 (N_5349,N_4768,N_4554);
nor U5350 (N_5350,N_4853,N_4124);
and U5351 (N_5351,N_4163,N_4089);
or U5352 (N_5352,N_4164,N_4111);
xor U5353 (N_5353,N_4509,N_4092);
or U5354 (N_5354,N_4395,N_4071);
xor U5355 (N_5355,N_4237,N_4356);
xor U5356 (N_5356,N_4615,N_4784);
xor U5357 (N_5357,N_4182,N_4635);
nor U5358 (N_5358,N_4037,N_4967);
and U5359 (N_5359,N_4459,N_4306);
nand U5360 (N_5360,N_4335,N_4070);
and U5361 (N_5361,N_4452,N_4361);
or U5362 (N_5362,N_4772,N_4616);
nor U5363 (N_5363,N_4901,N_4705);
or U5364 (N_5364,N_4363,N_4613);
xor U5365 (N_5365,N_4431,N_4250);
or U5366 (N_5366,N_4812,N_4517);
xnor U5367 (N_5367,N_4223,N_4427);
nand U5368 (N_5368,N_4457,N_4544);
xor U5369 (N_5369,N_4280,N_4934);
and U5370 (N_5370,N_4936,N_4707);
xnor U5371 (N_5371,N_4648,N_4547);
or U5372 (N_5372,N_4031,N_4488);
nand U5373 (N_5373,N_4097,N_4247);
nor U5374 (N_5374,N_4526,N_4522);
and U5375 (N_5375,N_4147,N_4502);
and U5376 (N_5376,N_4135,N_4384);
and U5377 (N_5377,N_4865,N_4397);
nor U5378 (N_5378,N_4766,N_4151);
nor U5379 (N_5379,N_4143,N_4925);
or U5380 (N_5380,N_4495,N_4246);
and U5381 (N_5381,N_4513,N_4965);
and U5382 (N_5382,N_4579,N_4680);
nand U5383 (N_5383,N_4022,N_4215);
and U5384 (N_5384,N_4518,N_4094);
nand U5385 (N_5385,N_4275,N_4564);
and U5386 (N_5386,N_4125,N_4311);
or U5387 (N_5387,N_4028,N_4892);
and U5388 (N_5388,N_4542,N_4347);
and U5389 (N_5389,N_4753,N_4507);
xnor U5390 (N_5390,N_4691,N_4098);
xor U5391 (N_5391,N_4081,N_4271);
xor U5392 (N_5392,N_4221,N_4175);
or U5393 (N_5393,N_4108,N_4653);
and U5394 (N_5394,N_4087,N_4964);
or U5395 (N_5395,N_4320,N_4315);
and U5396 (N_5396,N_4578,N_4258);
and U5397 (N_5397,N_4109,N_4308);
xnor U5398 (N_5398,N_4618,N_4796);
nor U5399 (N_5399,N_4206,N_4722);
nand U5400 (N_5400,N_4859,N_4558);
nor U5401 (N_5401,N_4146,N_4048);
nand U5402 (N_5402,N_4924,N_4360);
nand U5403 (N_5403,N_4379,N_4380);
or U5404 (N_5404,N_4485,N_4510);
or U5405 (N_5405,N_4684,N_4463);
nor U5406 (N_5406,N_4971,N_4848);
and U5407 (N_5407,N_4091,N_4839);
or U5408 (N_5408,N_4090,N_4570);
and U5409 (N_5409,N_4709,N_4214);
or U5410 (N_5410,N_4303,N_4289);
nand U5411 (N_5411,N_4953,N_4721);
nor U5412 (N_5412,N_4155,N_4590);
nand U5413 (N_5413,N_4466,N_4462);
or U5414 (N_5414,N_4655,N_4639);
nor U5415 (N_5415,N_4890,N_4490);
nand U5416 (N_5416,N_4494,N_4630);
and U5417 (N_5417,N_4113,N_4729);
xor U5418 (N_5418,N_4244,N_4102);
and U5419 (N_5419,N_4670,N_4589);
nand U5420 (N_5420,N_4663,N_4845);
nor U5421 (N_5421,N_4078,N_4238);
xor U5422 (N_5422,N_4248,N_4279);
nor U5423 (N_5423,N_4471,N_4026);
and U5424 (N_5424,N_4184,N_4412);
nand U5425 (N_5425,N_4236,N_4941);
or U5426 (N_5426,N_4726,N_4060);
nor U5427 (N_5427,N_4021,N_4419);
xor U5428 (N_5428,N_4180,N_4867);
xor U5429 (N_5429,N_4993,N_4549);
nand U5430 (N_5430,N_4218,N_4033);
nor U5431 (N_5431,N_4010,N_4383);
or U5432 (N_5432,N_4195,N_4597);
xnor U5433 (N_5433,N_4228,N_4283);
nand U5434 (N_5434,N_4136,N_4024);
or U5435 (N_5435,N_4719,N_4951);
or U5436 (N_5436,N_4895,N_4424);
and U5437 (N_5437,N_4112,N_4204);
xnor U5438 (N_5438,N_4738,N_4660);
and U5439 (N_5439,N_4042,N_4546);
and U5440 (N_5440,N_4277,N_4535);
nor U5441 (N_5441,N_4467,N_4192);
or U5442 (N_5442,N_4207,N_4349);
and U5443 (N_5443,N_4329,N_4593);
nand U5444 (N_5444,N_4103,N_4150);
and U5445 (N_5445,N_4405,N_4560);
and U5446 (N_5446,N_4074,N_4982);
nor U5447 (N_5447,N_4712,N_4222);
or U5448 (N_5448,N_4773,N_4515);
xor U5449 (N_5449,N_4168,N_4058);
xnor U5450 (N_5450,N_4257,N_4219);
xnor U5451 (N_5451,N_4725,N_4692);
xor U5452 (N_5452,N_4626,N_4373);
xnor U5453 (N_5453,N_4433,N_4566);
nand U5454 (N_5454,N_4706,N_4270);
or U5455 (N_5455,N_4562,N_4406);
or U5456 (N_5456,N_4186,N_4475);
xnor U5457 (N_5457,N_4132,N_4830);
nor U5458 (N_5458,N_4838,N_4348);
nor U5459 (N_5459,N_4101,N_4778);
xor U5460 (N_5460,N_4122,N_4290);
xnor U5461 (N_5461,N_4009,N_4917);
nand U5462 (N_5462,N_4786,N_4232);
and U5463 (N_5463,N_4723,N_4638);
xnor U5464 (N_5464,N_4840,N_4392);
xor U5465 (N_5465,N_4939,N_4906);
nor U5466 (N_5466,N_4174,N_4514);
nor U5467 (N_5467,N_4516,N_4981);
xnor U5468 (N_5468,N_4252,N_4177);
nor U5469 (N_5469,N_4017,N_4371);
nor U5470 (N_5470,N_4095,N_4732);
xnor U5471 (N_5471,N_4937,N_4233);
or U5472 (N_5472,N_4201,N_4032);
xor U5473 (N_5473,N_4332,N_4437);
nand U5474 (N_5474,N_4226,N_4813);
and U5475 (N_5475,N_4046,N_4064);
or U5476 (N_5476,N_4390,N_4915);
xnor U5477 (N_5477,N_4972,N_4370);
nand U5478 (N_5478,N_4781,N_4240);
nand U5479 (N_5479,N_4389,N_4393);
nor U5480 (N_5480,N_4443,N_4359);
nor U5481 (N_5481,N_4497,N_4531);
or U5482 (N_5482,N_4621,N_4015);
or U5483 (N_5483,N_4961,N_4994);
nand U5484 (N_5484,N_4259,N_4647);
and U5485 (N_5485,N_4864,N_4905);
xor U5486 (N_5486,N_4944,N_4881);
nand U5487 (N_5487,N_4775,N_4809);
xor U5488 (N_5488,N_4263,N_4505);
and U5489 (N_5489,N_4998,N_4771);
and U5490 (N_5490,N_4920,N_4884);
nor U5491 (N_5491,N_4664,N_4194);
and U5492 (N_5492,N_4742,N_4874);
or U5493 (N_5493,N_4404,N_4780);
nand U5494 (N_5494,N_4050,N_4506);
or U5495 (N_5495,N_4489,N_4239);
and U5496 (N_5496,N_4341,N_4454);
or U5497 (N_5497,N_4765,N_4637);
xnor U5498 (N_5498,N_4970,N_4056);
nor U5499 (N_5499,N_4559,N_4628);
nand U5500 (N_5500,N_4802,N_4150);
or U5501 (N_5501,N_4286,N_4074);
xor U5502 (N_5502,N_4151,N_4754);
nor U5503 (N_5503,N_4073,N_4357);
nor U5504 (N_5504,N_4423,N_4887);
nand U5505 (N_5505,N_4195,N_4039);
or U5506 (N_5506,N_4631,N_4269);
or U5507 (N_5507,N_4152,N_4500);
and U5508 (N_5508,N_4871,N_4578);
xnor U5509 (N_5509,N_4736,N_4345);
xor U5510 (N_5510,N_4329,N_4412);
xnor U5511 (N_5511,N_4975,N_4728);
and U5512 (N_5512,N_4528,N_4147);
nand U5513 (N_5513,N_4890,N_4943);
nor U5514 (N_5514,N_4740,N_4971);
nor U5515 (N_5515,N_4580,N_4077);
and U5516 (N_5516,N_4318,N_4733);
or U5517 (N_5517,N_4979,N_4797);
and U5518 (N_5518,N_4996,N_4050);
nor U5519 (N_5519,N_4337,N_4186);
nor U5520 (N_5520,N_4668,N_4578);
and U5521 (N_5521,N_4428,N_4152);
nand U5522 (N_5522,N_4875,N_4867);
and U5523 (N_5523,N_4948,N_4765);
xor U5524 (N_5524,N_4367,N_4001);
or U5525 (N_5525,N_4795,N_4241);
and U5526 (N_5526,N_4209,N_4579);
xnor U5527 (N_5527,N_4999,N_4020);
nor U5528 (N_5528,N_4805,N_4627);
nor U5529 (N_5529,N_4337,N_4112);
nor U5530 (N_5530,N_4718,N_4646);
nor U5531 (N_5531,N_4852,N_4097);
or U5532 (N_5532,N_4024,N_4547);
nand U5533 (N_5533,N_4257,N_4388);
or U5534 (N_5534,N_4850,N_4554);
xor U5535 (N_5535,N_4912,N_4425);
nand U5536 (N_5536,N_4064,N_4293);
nand U5537 (N_5537,N_4322,N_4988);
nor U5538 (N_5538,N_4019,N_4705);
nand U5539 (N_5539,N_4525,N_4832);
xor U5540 (N_5540,N_4970,N_4739);
xor U5541 (N_5541,N_4502,N_4242);
nand U5542 (N_5542,N_4714,N_4803);
or U5543 (N_5543,N_4213,N_4948);
and U5544 (N_5544,N_4200,N_4931);
and U5545 (N_5545,N_4766,N_4453);
or U5546 (N_5546,N_4371,N_4478);
and U5547 (N_5547,N_4811,N_4005);
xnor U5548 (N_5548,N_4217,N_4548);
and U5549 (N_5549,N_4675,N_4699);
or U5550 (N_5550,N_4005,N_4543);
or U5551 (N_5551,N_4218,N_4339);
nor U5552 (N_5552,N_4150,N_4006);
nor U5553 (N_5553,N_4230,N_4713);
or U5554 (N_5554,N_4688,N_4852);
nand U5555 (N_5555,N_4745,N_4725);
nand U5556 (N_5556,N_4991,N_4332);
nor U5557 (N_5557,N_4187,N_4198);
and U5558 (N_5558,N_4948,N_4727);
nor U5559 (N_5559,N_4872,N_4283);
nand U5560 (N_5560,N_4926,N_4032);
and U5561 (N_5561,N_4466,N_4959);
nand U5562 (N_5562,N_4649,N_4413);
and U5563 (N_5563,N_4599,N_4142);
or U5564 (N_5564,N_4090,N_4550);
nand U5565 (N_5565,N_4146,N_4210);
and U5566 (N_5566,N_4567,N_4572);
nor U5567 (N_5567,N_4248,N_4985);
nor U5568 (N_5568,N_4401,N_4689);
nand U5569 (N_5569,N_4283,N_4002);
xnor U5570 (N_5570,N_4668,N_4551);
or U5571 (N_5571,N_4548,N_4986);
nand U5572 (N_5572,N_4320,N_4960);
or U5573 (N_5573,N_4974,N_4415);
xor U5574 (N_5574,N_4160,N_4072);
and U5575 (N_5575,N_4771,N_4478);
or U5576 (N_5576,N_4195,N_4467);
nand U5577 (N_5577,N_4600,N_4483);
or U5578 (N_5578,N_4300,N_4685);
and U5579 (N_5579,N_4569,N_4994);
xor U5580 (N_5580,N_4837,N_4758);
or U5581 (N_5581,N_4709,N_4682);
xor U5582 (N_5582,N_4802,N_4798);
nand U5583 (N_5583,N_4699,N_4671);
or U5584 (N_5584,N_4189,N_4085);
nor U5585 (N_5585,N_4148,N_4472);
nand U5586 (N_5586,N_4739,N_4046);
nand U5587 (N_5587,N_4531,N_4988);
nor U5588 (N_5588,N_4780,N_4037);
and U5589 (N_5589,N_4070,N_4973);
or U5590 (N_5590,N_4387,N_4497);
xor U5591 (N_5591,N_4492,N_4834);
xor U5592 (N_5592,N_4939,N_4916);
xor U5593 (N_5593,N_4307,N_4960);
xnor U5594 (N_5594,N_4755,N_4364);
or U5595 (N_5595,N_4647,N_4246);
or U5596 (N_5596,N_4145,N_4150);
xnor U5597 (N_5597,N_4724,N_4390);
and U5598 (N_5598,N_4950,N_4653);
nand U5599 (N_5599,N_4528,N_4156);
nor U5600 (N_5600,N_4867,N_4090);
and U5601 (N_5601,N_4937,N_4445);
or U5602 (N_5602,N_4624,N_4283);
or U5603 (N_5603,N_4057,N_4329);
and U5604 (N_5604,N_4151,N_4601);
or U5605 (N_5605,N_4566,N_4936);
or U5606 (N_5606,N_4565,N_4330);
xor U5607 (N_5607,N_4572,N_4194);
nor U5608 (N_5608,N_4643,N_4358);
nor U5609 (N_5609,N_4998,N_4140);
nand U5610 (N_5610,N_4567,N_4846);
and U5611 (N_5611,N_4964,N_4177);
xnor U5612 (N_5612,N_4383,N_4552);
or U5613 (N_5613,N_4347,N_4027);
and U5614 (N_5614,N_4682,N_4225);
and U5615 (N_5615,N_4961,N_4199);
nand U5616 (N_5616,N_4585,N_4548);
nor U5617 (N_5617,N_4920,N_4576);
or U5618 (N_5618,N_4585,N_4021);
nand U5619 (N_5619,N_4908,N_4302);
and U5620 (N_5620,N_4248,N_4203);
nor U5621 (N_5621,N_4879,N_4162);
and U5622 (N_5622,N_4673,N_4805);
nor U5623 (N_5623,N_4956,N_4810);
and U5624 (N_5624,N_4251,N_4817);
and U5625 (N_5625,N_4874,N_4563);
and U5626 (N_5626,N_4845,N_4184);
and U5627 (N_5627,N_4054,N_4800);
nor U5628 (N_5628,N_4780,N_4059);
or U5629 (N_5629,N_4653,N_4791);
nand U5630 (N_5630,N_4860,N_4109);
and U5631 (N_5631,N_4703,N_4230);
and U5632 (N_5632,N_4726,N_4374);
nand U5633 (N_5633,N_4110,N_4004);
xor U5634 (N_5634,N_4965,N_4087);
and U5635 (N_5635,N_4327,N_4713);
xor U5636 (N_5636,N_4260,N_4958);
xnor U5637 (N_5637,N_4943,N_4285);
or U5638 (N_5638,N_4671,N_4419);
and U5639 (N_5639,N_4174,N_4236);
nor U5640 (N_5640,N_4600,N_4757);
nor U5641 (N_5641,N_4997,N_4893);
xnor U5642 (N_5642,N_4693,N_4205);
nor U5643 (N_5643,N_4431,N_4761);
nor U5644 (N_5644,N_4909,N_4974);
and U5645 (N_5645,N_4262,N_4956);
and U5646 (N_5646,N_4486,N_4403);
and U5647 (N_5647,N_4120,N_4330);
nor U5648 (N_5648,N_4255,N_4177);
and U5649 (N_5649,N_4844,N_4776);
and U5650 (N_5650,N_4155,N_4154);
and U5651 (N_5651,N_4083,N_4274);
xnor U5652 (N_5652,N_4919,N_4123);
or U5653 (N_5653,N_4611,N_4515);
and U5654 (N_5654,N_4017,N_4707);
xor U5655 (N_5655,N_4786,N_4399);
nand U5656 (N_5656,N_4343,N_4226);
xor U5657 (N_5657,N_4638,N_4481);
and U5658 (N_5658,N_4089,N_4414);
nand U5659 (N_5659,N_4144,N_4365);
nor U5660 (N_5660,N_4525,N_4467);
and U5661 (N_5661,N_4964,N_4218);
nand U5662 (N_5662,N_4545,N_4769);
nor U5663 (N_5663,N_4610,N_4674);
nand U5664 (N_5664,N_4704,N_4709);
and U5665 (N_5665,N_4187,N_4361);
and U5666 (N_5666,N_4181,N_4604);
and U5667 (N_5667,N_4662,N_4518);
and U5668 (N_5668,N_4280,N_4414);
or U5669 (N_5669,N_4752,N_4673);
and U5670 (N_5670,N_4543,N_4459);
and U5671 (N_5671,N_4796,N_4535);
nand U5672 (N_5672,N_4164,N_4711);
or U5673 (N_5673,N_4408,N_4880);
nor U5674 (N_5674,N_4787,N_4285);
and U5675 (N_5675,N_4554,N_4744);
nor U5676 (N_5676,N_4961,N_4469);
xnor U5677 (N_5677,N_4056,N_4317);
and U5678 (N_5678,N_4024,N_4669);
nor U5679 (N_5679,N_4593,N_4412);
xor U5680 (N_5680,N_4230,N_4217);
or U5681 (N_5681,N_4538,N_4920);
xor U5682 (N_5682,N_4666,N_4659);
or U5683 (N_5683,N_4541,N_4831);
nor U5684 (N_5684,N_4959,N_4176);
and U5685 (N_5685,N_4382,N_4102);
xnor U5686 (N_5686,N_4321,N_4102);
xnor U5687 (N_5687,N_4981,N_4221);
nand U5688 (N_5688,N_4709,N_4999);
nand U5689 (N_5689,N_4282,N_4364);
and U5690 (N_5690,N_4057,N_4804);
nand U5691 (N_5691,N_4779,N_4849);
nor U5692 (N_5692,N_4817,N_4052);
or U5693 (N_5693,N_4063,N_4242);
or U5694 (N_5694,N_4152,N_4739);
nor U5695 (N_5695,N_4688,N_4714);
nor U5696 (N_5696,N_4097,N_4181);
nor U5697 (N_5697,N_4472,N_4146);
nor U5698 (N_5698,N_4505,N_4360);
nor U5699 (N_5699,N_4984,N_4280);
nor U5700 (N_5700,N_4323,N_4632);
and U5701 (N_5701,N_4099,N_4990);
nor U5702 (N_5702,N_4936,N_4118);
or U5703 (N_5703,N_4453,N_4391);
nor U5704 (N_5704,N_4482,N_4611);
and U5705 (N_5705,N_4923,N_4922);
xor U5706 (N_5706,N_4174,N_4698);
nand U5707 (N_5707,N_4651,N_4090);
xnor U5708 (N_5708,N_4421,N_4636);
nor U5709 (N_5709,N_4083,N_4114);
nor U5710 (N_5710,N_4993,N_4126);
and U5711 (N_5711,N_4566,N_4608);
and U5712 (N_5712,N_4852,N_4342);
xnor U5713 (N_5713,N_4751,N_4370);
nand U5714 (N_5714,N_4595,N_4042);
nor U5715 (N_5715,N_4490,N_4735);
and U5716 (N_5716,N_4045,N_4653);
and U5717 (N_5717,N_4214,N_4079);
nor U5718 (N_5718,N_4834,N_4024);
or U5719 (N_5719,N_4430,N_4795);
and U5720 (N_5720,N_4067,N_4495);
and U5721 (N_5721,N_4933,N_4203);
nand U5722 (N_5722,N_4487,N_4966);
and U5723 (N_5723,N_4512,N_4882);
nor U5724 (N_5724,N_4729,N_4884);
xnor U5725 (N_5725,N_4526,N_4895);
and U5726 (N_5726,N_4163,N_4392);
and U5727 (N_5727,N_4142,N_4601);
xor U5728 (N_5728,N_4361,N_4023);
or U5729 (N_5729,N_4976,N_4469);
or U5730 (N_5730,N_4111,N_4388);
or U5731 (N_5731,N_4851,N_4267);
xnor U5732 (N_5732,N_4534,N_4609);
or U5733 (N_5733,N_4678,N_4531);
and U5734 (N_5734,N_4802,N_4403);
nand U5735 (N_5735,N_4868,N_4465);
nand U5736 (N_5736,N_4448,N_4732);
nand U5737 (N_5737,N_4594,N_4181);
nor U5738 (N_5738,N_4943,N_4852);
or U5739 (N_5739,N_4451,N_4470);
or U5740 (N_5740,N_4813,N_4802);
and U5741 (N_5741,N_4954,N_4049);
and U5742 (N_5742,N_4391,N_4671);
or U5743 (N_5743,N_4429,N_4935);
nand U5744 (N_5744,N_4791,N_4498);
nand U5745 (N_5745,N_4823,N_4141);
and U5746 (N_5746,N_4662,N_4470);
nor U5747 (N_5747,N_4476,N_4867);
nor U5748 (N_5748,N_4052,N_4778);
xnor U5749 (N_5749,N_4192,N_4074);
xnor U5750 (N_5750,N_4263,N_4089);
and U5751 (N_5751,N_4765,N_4479);
nor U5752 (N_5752,N_4266,N_4511);
and U5753 (N_5753,N_4998,N_4595);
and U5754 (N_5754,N_4803,N_4470);
or U5755 (N_5755,N_4821,N_4056);
nand U5756 (N_5756,N_4598,N_4118);
xor U5757 (N_5757,N_4138,N_4353);
and U5758 (N_5758,N_4868,N_4098);
and U5759 (N_5759,N_4921,N_4252);
or U5760 (N_5760,N_4943,N_4965);
and U5761 (N_5761,N_4327,N_4181);
xnor U5762 (N_5762,N_4830,N_4826);
or U5763 (N_5763,N_4518,N_4504);
nand U5764 (N_5764,N_4205,N_4128);
or U5765 (N_5765,N_4179,N_4824);
nor U5766 (N_5766,N_4293,N_4827);
xnor U5767 (N_5767,N_4164,N_4367);
and U5768 (N_5768,N_4626,N_4935);
xor U5769 (N_5769,N_4603,N_4861);
or U5770 (N_5770,N_4644,N_4552);
or U5771 (N_5771,N_4144,N_4005);
and U5772 (N_5772,N_4920,N_4648);
xor U5773 (N_5773,N_4114,N_4186);
or U5774 (N_5774,N_4789,N_4546);
nor U5775 (N_5775,N_4263,N_4684);
and U5776 (N_5776,N_4326,N_4719);
and U5777 (N_5777,N_4284,N_4624);
xor U5778 (N_5778,N_4003,N_4605);
xor U5779 (N_5779,N_4207,N_4851);
xnor U5780 (N_5780,N_4618,N_4254);
nor U5781 (N_5781,N_4502,N_4214);
or U5782 (N_5782,N_4270,N_4573);
xnor U5783 (N_5783,N_4906,N_4022);
and U5784 (N_5784,N_4603,N_4604);
and U5785 (N_5785,N_4661,N_4126);
or U5786 (N_5786,N_4222,N_4365);
or U5787 (N_5787,N_4204,N_4273);
xnor U5788 (N_5788,N_4875,N_4681);
and U5789 (N_5789,N_4647,N_4990);
and U5790 (N_5790,N_4385,N_4409);
nor U5791 (N_5791,N_4006,N_4028);
nand U5792 (N_5792,N_4400,N_4433);
nand U5793 (N_5793,N_4421,N_4837);
nor U5794 (N_5794,N_4056,N_4680);
or U5795 (N_5795,N_4289,N_4763);
nand U5796 (N_5796,N_4263,N_4974);
nand U5797 (N_5797,N_4931,N_4099);
nand U5798 (N_5798,N_4824,N_4910);
nor U5799 (N_5799,N_4327,N_4304);
nor U5800 (N_5800,N_4498,N_4743);
or U5801 (N_5801,N_4757,N_4894);
nor U5802 (N_5802,N_4785,N_4017);
xnor U5803 (N_5803,N_4781,N_4250);
xnor U5804 (N_5804,N_4293,N_4320);
xor U5805 (N_5805,N_4109,N_4737);
and U5806 (N_5806,N_4767,N_4660);
nand U5807 (N_5807,N_4086,N_4757);
nand U5808 (N_5808,N_4441,N_4637);
nor U5809 (N_5809,N_4451,N_4857);
or U5810 (N_5810,N_4647,N_4825);
nor U5811 (N_5811,N_4199,N_4843);
and U5812 (N_5812,N_4445,N_4056);
xnor U5813 (N_5813,N_4770,N_4031);
xor U5814 (N_5814,N_4403,N_4977);
or U5815 (N_5815,N_4874,N_4631);
nand U5816 (N_5816,N_4317,N_4226);
nand U5817 (N_5817,N_4165,N_4137);
nor U5818 (N_5818,N_4272,N_4581);
xnor U5819 (N_5819,N_4710,N_4656);
nor U5820 (N_5820,N_4305,N_4149);
and U5821 (N_5821,N_4631,N_4681);
nor U5822 (N_5822,N_4515,N_4047);
nor U5823 (N_5823,N_4337,N_4316);
or U5824 (N_5824,N_4198,N_4792);
xnor U5825 (N_5825,N_4467,N_4217);
nand U5826 (N_5826,N_4561,N_4107);
nand U5827 (N_5827,N_4828,N_4815);
and U5828 (N_5828,N_4875,N_4264);
or U5829 (N_5829,N_4847,N_4927);
or U5830 (N_5830,N_4286,N_4958);
nand U5831 (N_5831,N_4519,N_4453);
and U5832 (N_5832,N_4500,N_4874);
or U5833 (N_5833,N_4898,N_4151);
nor U5834 (N_5834,N_4004,N_4918);
xnor U5835 (N_5835,N_4032,N_4810);
and U5836 (N_5836,N_4226,N_4711);
nand U5837 (N_5837,N_4987,N_4526);
nor U5838 (N_5838,N_4317,N_4480);
and U5839 (N_5839,N_4548,N_4730);
or U5840 (N_5840,N_4703,N_4557);
xnor U5841 (N_5841,N_4435,N_4266);
nor U5842 (N_5842,N_4741,N_4830);
nand U5843 (N_5843,N_4711,N_4764);
or U5844 (N_5844,N_4845,N_4961);
and U5845 (N_5845,N_4331,N_4020);
and U5846 (N_5846,N_4015,N_4645);
and U5847 (N_5847,N_4124,N_4126);
nand U5848 (N_5848,N_4849,N_4422);
nand U5849 (N_5849,N_4151,N_4994);
nand U5850 (N_5850,N_4906,N_4393);
nand U5851 (N_5851,N_4276,N_4938);
or U5852 (N_5852,N_4783,N_4598);
xnor U5853 (N_5853,N_4470,N_4333);
nand U5854 (N_5854,N_4961,N_4736);
xor U5855 (N_5855,N_4120,N_4314);
xor U5856 (N_5856,N_4833,N_4034);
and U5857 (N_5857,N_4611,N_4984);
nand U5858 (N_5858,N_4374,N_4330);
xor U5859 (N_5859,N_4376,N_4034);
and U5860 (N_5860,N_4400,N_4309);
or U5861 (N_5861,N_4628,N_4683);
nor U5862 (N_5862,N_4658,N_4330);
nor U5863 (N_5863,N_4880,N_4419);
or U5864 (N_5864,N_4554,N_4969);
nor U5865 (N_5865,N_4725,N_4813);
and U5866 (N_5866,N_4576,N_4633);
nand U5867 (N_5867,N_4105,N_4029);
nor U5868 (N_5868,N_4186,N_4208);
or U5869 (N_5869,N_4646,N_4173);
and U5870 (N_5870,N_4548,N_4317);
or U5871 (N_5871,N_4472,N_4089);
nor U5872 (N_5872,N_4394,N_4067);
nor U5873 (N_5873,N_4914,N_4212);
nor U5874 (N_5874,N_4257,N_4073);
and U5875 (N_5875,N_4884,N_4604);
nand U5876 (N_5876,N_4101,N_4458);
and U5877 (N_5877,N_4688,N_4516);
xor U5878 (N_5878,N_4901,N_4200);
and U5879 (N_5879,N_4582,N_4189);
nor U5880 (N_5880,N_4092,N_4331);
nand U5881 (N_5881,N_4441,N_4965);
xor U5882 (N_5882,N_4672,N_4431);
nand U5883 (N_5883,N_4301,N_4712);
xnor U5884 (N_5884,N_4988,N_4670);
nor U5885 (N_5885,N_4305,N_4790);
or U5886 (N_5886,N_4011,N_4018);
and U5887 (N_5887,N_4166,N_4941);
nand U5888 (N_5888,N_4026,N_4152);
xor U5889 (N_5889,N_4874,N_4428);
xor U5890 (N_5890,N_4665,N_4327);
nand U5891 (N_5891,N_4575,N_4987);
or U5892 (N_5892,N_4222,N_4792);
nor U5893 (N_5893,N_4805,N_4043);
xnor U5894 (N_5894,N_4531,N_4903);
nand U5895 (N_5895,N_4788,N_4718);
xnor U5896 (N_5896,N_4725,N_4357);
nor U5897 (N_5897,N_4110,N_4206);
and U5898 (N_5898,N_4922,N_4700);
nand U5899 (N_5899,N_4638,N_4077);
and U5900 (N_5900,N_4845,N_4150);
nand U5901 (N_5901,N_4484,N_4895);
or U5902 (N_5902,N_4595,N_4646);
nor U5903 (N_5903,N_4630,N_4423);
nor U5904 (N_5904,N_4940,N_4290);
and U5905 (N_5905,N_4978,N_4159);
xor U5906 (N_5906,N_4330,N_4922);
xnor U5907 (N_5907,N_4017,N_4770);
or U5908 (N_5908,N_4828,N_4288);
and U5909 (N_5909,N_4912,N_4599);
nor U5910 (N_5910,N_4647,N_4837);
nand U5911 (N_5911,N_4740,N_4137);
xnor U5912 (N_5912,N_4665,N_4156);
nand U5913 (N_5913,N_4598,N_4062);
nand U5914 (N_5914,N_4515,N_4697);
and U5915 (N_5915,N_4268,N_4315);
nor U5916 (N_5916,N_4838,N_4777);
and U5917 (N_5917,N_4136,N_4491);
xnor U5918 (N_5918,N_4060,N_4099);
and U5919 (N_5919,N_4010,N_4716);
xnor U5920 (N_5920,N_4055,N_4563);
or U5921 (N_5921,N_4948,N_4695);
or U5922 (N_5922,N_4456,N_4719);
nor U5923 (N_5923,N_4564,N_4553);
or U5924 (N_5924,N_4576,N_4854);
xor U5925 (N_5925,N_4730,N_4554);
nor U5926 (N_5926,N_4875,N_4156);
xor U5927 (N_5927,N_4025,N_4665);
and U5928 (N_5928,N_4731,N_4026);
and U5929 (N_5929,N_4082,N_4386);
nor U5930 (N_5930,N_4129,N_4956);
and U5931 (N_5931,N_4621,N_4543);
xnor U5932 (N_5932,N_4871,N_4786);
nor U5933 (N_5933,N_4580,N_4987);
nor U5934 (N_5934,N_4989,N_4824);
or U5935 (N_5935,N_4724,N_4673);
nor U5936 (N_5936,N_4585,N_4341);
or U5937 (N_5937,N_4294,N_4932);
and U5938 (N_5938,N_4687,N_4284);
and U5939 (N_5939,N_4780,N_4057);
nor U5940 (N_5940,N_4538,N_4800);
nand U5941 (N_5941,N_4691,N_4176);
and U5942 (N_5942,N_4727,N_4594);
or U5943 (N_5943,N_4366,N_4684);
and U5944 (N_5944,N_4784,N_4225);
and U5945 (N_5945,N_4079,N_4774);
xor U5946 (N_5946,N_4993,N_4129);
and U5947 (N_5947,N_4864,N_4298);
or U5948 (N_5948,N_4999,N_4711);
nand U5949 (N_5949,N_4217,N_4945);
xnor U5950 (N_5950,N_4846,N_4120);
xor U5951 (N_5951,N_4379,N_4164);
nand U5952 (N_5952,N_4931,N_4177);
nor U5953 (N_5953,N_4654,N_4692);
and U5954 (N_5954,N_4937,N_4197);
xnor U5955 (N_5955,N_4788,N_4924);
xnor U5956 (N_5956,N_4436,N_4017);
and U5957 (N_5957,N_4899,N_4791);
nand U5958 (N_5958,N_4375,N_4324);
nor U5959 (N_5959,N_4545,N_4795);
xnor U5960 (N_5960,N_4397,N_4647);
nor U5961 (N_5961,N_4938,N_4768);
nand U5962 (N_5962,N_4685,N_4739);
and U5963 (N_5963,N_4588,N_4911);
nand U5964 (N_5964,N_4377,N_4353);
and U5965 (N_5965,N_4474,N_4122);
nand U5966 (N_5966,N_4734,N_4766);
or U5967 (N_5967,N_4623,N_4264);
xor U5968 (N_5968,N_4458,N_4806);
or U5969 (N_5969,N_4860,N_4898);
nor U5970 (N_5970,N_4646,N_4837);
or U5971 (N_5971,N_4279,N_4176);
xnor U5972 (N_5972,N_4558,N_4172);
nor U5973 (N_5973,N_4052,N_4591);
or U5974 (N_5974,N_4970,N_4652);
nand U5975 (N_5975,N_4406,N_4063);
nor U5976 (N_5976,N_4030,N_4856);
or U5977 (N_5977,N_4257,N_4185);
nand U5978 (N_5978,N_4214,N_4412);
xor U5979 (N_5979,N_4730,N_4351);
or U5980 (N_5980,N_4675,N_4943);
xnor U5981 (N_5981,N_4678,N_4372);
nor U5982 (N_5982,N_4698,N_4386);
or U5983 (N_5983,N_4266,N_4880);
or U5984 (N_5984,N_4663,N_4790);
nor U5985 (N_5985,N_4842,N_4654);
and U5986 (N_5986,N_4736,N_4743);
nand U5987 (N_5987,N_4632,N_4038);
xnor U5988 (N_5988,N_4403,N_4402);
or U5989 (N_5989,N_4042,N_4154);
xnor U5990 (N_5990,N_4385,N_4326);
nand U5991 (N_5991,N_4147,N_4737);
nor U5992 (N_5992,N_4407,N_4961);
nor U5993 (N_5993,N_4979,N_4132);
or U5994 (N_5994,N_4114,N_4604);
and U5995 (N_5995,N_4509,N_4477);
nand U5996 (N_5996,N_4641,N_4051);
nand U5997 (N_5997,N_4823,N_4186);
or U5998 (N_5998,N_4265,N_4896);
nand U5999 (N_5999,N_4997,N_4075);
or U6000 (N_6000,N_5839,N_5374);
nor U6001 (N_6001,N_5728,N_5335);
nand U6002 (N_6002,N_5521,N_5247);
nor U6003 (N_6003,N_5501,N_5371);
nand U6004 (N_6004,N_5519,N_5674);
xnor U6005 (N_6005,N_5838,N_5128);
and U6006 (N_6006,N_5716,N_5555);
and U6007 (N_6007,N_5605,N_5717);
or U6008 (N_6008,N_5432,N_5575);
and U6009 (N_6009,N_5206,N_5922);
nor U6010 (N_6010,N_5229,N_5100);
nand U6011 (N_6011,N_5185,N_5828);
xor U6012 (N_6012,N_5204,N_5987);
nor U6013 (N_6013,N_5344,N_5392);
xor U6014 (N_6014,N_5012,N_5773);
nor U6015 (N_6015,N_5403,N_5009);
nor U6016 (N_6016,N_5168,N_5934);
nor U6017 (N_6017,N_5439,N_5240);
nor U6018 (N_6018,N_5177,N_5492);
nor U6019 (N_6019,N_5119,N_5988);
nand U6020 (N_6020,N_5661,N_5946);
nor U6021 (N_6021,N_5338,N_5108);
xor U6022 (N_6022,N_5470,N_5103);
and U6023 (N_6023,N_5880,N_5513);
nand U6024 (N_6024,N_5604,N_5270);
nor U6025 (N_6025,N_5453,N_5027);
nand U6026 (N_6026,N_5502,N_5446);
xor U6027 (N_6027,N_5864,N_5423);
xnor U6028 (N_6028,N_5540,N_5074);
xor U6029 (N_6029,N_5539,N_5632);
nor U6030 (N_6030,N_5591,N_5789);
or U6031 (N_6031,N_5785,N_5564);
nand U6032 (N_6032,N_5391,N_5738);
and U6033 (N_6033,N_5452,N_5112);
and U6034 (N_6034,N_5703,N_5192);
or U6035 (N_6035,N_5816,N_5412);
or U6036 (N_6036,N_5277,N_5053);
or U6037 (N_6037,N_5924,N_5817);
and U6038 (N_6038,N_5249,N_5754);
and U6039 (N_6039,N_5551,N_5169);
nand U6040 (N_6040,N_5760,N_5520);
xnor U6041 (N_6041,N_5508,N_5862);
nor U6042 (N_6042,N_5748,N_5241);
or U6043 (N_6043,N_5689,N_5741);
and U6044 (N_6044,N_5342,N_5263);
nand U6045 (N_6045,N_5003,N_5623);
and U6046 (N_6046,N_5228,N_5015);
and U6047 (N_6047,N_5352,N_5466);
nor U6048 (N_6048,N_5616,N_5954);
xnor U6049 (N_6049,N_5156,N_5246);
nand U6050 (N_6050,N_5145,N_5745);
or U6051 (N_6051,N_5291,N_5375);
and U6052 (N_6052,N_5357,N_5804);
nand U6053 (N_6053,N_5698,N_5991);
nor U6054 (N_6054,N_5434,N_5359);
nor U6055 (N_6055,N_5642,N_5589);
nor U6056 (N_6056,N_5460,N_5626);
nand U6057 (N_6057,N_5771,N_5800);
or U6058 (N_6058,N_5684,N_5346);
nor U6059 (N_6059,N_5621,N_5503);
xnor U6060 (N_6060,N_5682,N_5461);
or U6061 (N_6061,N_5381,N_5367);
nand U6062 (N_6062,N_5992,N_5272);
and U6063 (N_6063,N_5582,N_5147);
nor U6064 (N_6064,N_5530,N_5193);
xor U6065 (N_6065,N_5975,N_5651);
nand U6066 (N_6066,N_5814,N_5780);
nor U6067 (N_6067,N_5219,N_5625);
nor U6068 (N_6068,N_5711,N_5123);
nand U6069 (N_6069,N_5061,N_5259);
xor U6070 (N_6070,N_5732,N_5400);
and U6071 (N_6071,N_5404,N_5945);
nand U6072 (N_6072,N_5634,N_5523);
nand U6073 (N_6073,N_5552,N_5686);
nor U6074 (N_6074,N_5383,N_5170);
or U6075 (N_6075,N_5538,N_5268);
or U6076 (N_6076,N_5652,N_5330);
xnor U6077 (N_6077,N_5547,N_5543);
and U6078 (N_6078,N_5448,N_5244);
or U6079 (N_6079,N_5571,N_5829);
xor U6080 (N_6080,N_5340,N_5037);
or U6081 (N_6081,N_5557,N_5970);
or U6082 (N_6082,N_5072,N_5677);
xor U6083 (N_6083,N_5705,N_5603);
nand U6084 (N_6084,N_5960,N_5004);
nand U6085 (N_6085,N_5872,N_5458);
nand U6086 (N_6086,N_5051,N_5886);
or U6087 (N_6087,N_5030,N_5865);
or U6088 (N_6088,N_5570,N_5143);
or U6089 (N_6089,N_5251,N_5349);
xnor U6090 (N_6090,N_5545,N_5629);
nor U6091 (N_6091,N_5462,N_5791);
xor U6092 (N_6092,N_5468,N_5581);
or U6093 (N_6093,N_5336,N_5179);
and U6094 (N_6094,N_5046,N_5925);
nand U6095 (N_6095,N_5469,N_5242);
and U6096 (N_6096,N_5306,N_5062);
nor U6097 (N_6097,N_5735,N_5361);
and U6098 (N_6098,N_5088,N_5111);
nor U6099 (N_6099,N_5844,N_5495);
nand U6100 (N_6100,N_5653,N_5096);
xor U6101 (N_6101,N_5859,N_5070);
nand U6102 (N_6102,N_5284,N_5086);
nand U6103 (N_6103,N_5410,N_5282);
or U6104 (N_6104,N_5224,N_5038);
xor U6105 (N_6105,N_5022,N_5006);
xnor U6106 (N_6106,N_5333,N_5456);
nand U6107 (N_6107,N_5736,N_5216);
or U6108 (N_6108,N_5138,N_5560);
and U6109 (N_6109,N_5080,N_5858);
nor U6110 (N_6110,N_5226,N_5969);
nand U6111 (N_6111,N_5812,N_5120);
nand U6112 (N_6112,N_5093,N_5370);
or U6113 (N_6113,N_5943,N_5963);
nand U6114 (N_6114,N_5889,N_5426);
nand U6115 (N_6115,N_5576,N_5134);
nand U6116 (N_6116,N_5932,N_5874);
or U6117 (N_6117,N_5266,N_5092);
nor U6118 (N_6118,N_5965,N_5673);
and U6119 (N_6119,N_5904,N_5506);
or U6120 (N_6120,N_5064,N_5161);
nor U6121 (N_6121,N_5881,N_5611);
nand U6122 (N_6122,N_5183,N_5042);
or U6123 (N_6123,N_5348,N_5471);
and U6124 (N_6124,N_5721,N_5231);
and U6125 (N_6125,N_5562,N_5706);
and U6126 (N_6126,N_5610,N_5021);
nor U6127 (N_6127,N_5052,N_5985);
xnor U6128 (N_6128,N_5907,N_5917);
nor U6129 (N_6129,N_5890,N_5267);
xnor U6130 (N_6130,N_5303,N_5747);
or U6131 (N_6131,N_5989,N_5305);
or U6132 (N_6132,N_5429,N_5050);
xnor U6133 (N_6133,N_5607,N_5472);
and U6134 (N_6134,N_5522,N_5587);
nand U6135 (N_6135,N_5619,N_5307);
xnor U6136 (N_6136,N_5422,N_5056);
xnor U6137 (N_6137,N_5221,N_5424);
nor U6138 (N_6138,N_5384,N_5572);
and U6139 (N_6139,N_5905,N_5405);
nor U6140 (N_6140,N_5313,N_5002);
nor U6141 (N_6141,N_5309,N_5290);
xor U6142 (N_6142,N_5347,N_5912);
xnor U6143 (N_6143,N_5039,N_5644);
or U6144 (N_6144,N_5801,N_5067);
nor U6145 (N_6145,N_5876,N_5579);
xnor U6146 (N_6146,N_5578,N_5394);
nor U6147 (N_6147,N_5133,N_5250);
nand U6148 (N_6148,N_5967,N_5700);
xnor U6149 (N_6149,N_5189,N_5531);
and U6150 (N_6150,N_5797,N_5628);
nand U6151 (N_6151,N_5483,N_5713);
nand U6152 (N_6152,N_5379,N_5929);
nor U6153 (N_6153,N_5655,N_5569);
xnor U6154 (N_6154,N_5016,N_5436);
nand U6155 (N_6155,N_5317,N_5826);
and U6156 (N_6156,N_5909,N_5663);
and U6157 (N_6157,N_5648,N_5151);
xor U6158 (N_6158,N_5285,N_5157);
nor U6159 (N_6159,N_5852,N_5781);
xnor U6160 (N_6160,N_5040,N_5709);
and U6161 (N_6161,N_5159,N_5464);
nand U6162 (N_6162,N_5597,N_5299);
nor U6163 (N_6163,N_5851,N_5428);
or U6164 (N_6164,N_5645,N_5194);
nor U6165 (N_6165,N_5029,N_5903);
nand U6166 (N_6166,N_5755,N_5289);
nor U6167 (N_6167,N_5271,N_5697);
and U6168 (N_6168,N_5142,N_5395);
nor U6169 (N_6169,N_5149,N_5594);
and U6170 (N_6170,N_5236,N_5459);
and U6171 (N_6171,N_5961,N_5841);
xor U6172 (N_6172,N_5227,N_5136);
xor U6173 (N_6173,N_5435,N_5447);
nand U6174 (N_6174,N_5898,N_5406);
or U6175 (N_6175,N_5319,N_5366);
nand U6176 (N_6176,N_5883,N_5863);
nand U6177 (N_6177,N_5043,N_5982);
or U6178 (N_6178,N_5553,N_5048);
nand U6179 (N_6179,N_5065,N_5014);
nand U6180 (N_6180,N_5234,N_5107);
nor U6181 (N_6181,N_5121,N_5639);
and U6182 (N_6182,N_5514,N_5778);
nor U6183 (N_6183,N_5273,N_5203);
nor U6184 (N_6184,N_5467,N_5260);
nand U6185 (N_6185,N_5110,N_5327);
nor U6186 (N_6186,N_5976,N_5197);
nor U6187 (N_6187,N_5116,N_5171);
or U6188 (N_6188,N_5115,N_5692);
nand U6189 (N_6189,N_5060,N_5643);
or U6190 (N_6190,N_5507,N_5441);
nor U6191 (N_6191,N_5640,N_5548);
xnor U6192 (N_6192,N_5683,N_5845);
and U6193 (N_6193,N_5081,N_5978);
and U6194 (N_6194,N_5550,N_5165);
and U6195 (N_6195,N_5637,N_5613);
nor U6196 (N_6196,N_5546,N_5215);
xor U6197 (N_6197,N_5007,N_5650);
xnor U6198 (N_6198,N_5902,N_5387);
and U6199 (N_6199,N_5223,N_5822);
nor U6200 (N_6200,N_5117,N_5010);
or U6201 (N_6201,N_5083,N_5385);
or U6202 (N_6202,N_5199,N_5210);
or U6203 (N_6203,N_5025,N_5090);
nor U6204 (N_6204,N_5811,N_5959);
nor U6205 (N_6205,N_5847,N_5914);
and U6206 (N_6206,N_5580,N_5186);
or U6207 (N_6207,N_5983,N_5911);
and U6208 (N_6208,N_5444,N_5054);
xor U6209 (N_6209,N_5751,N_5465);
nor U6210 (N_6210,N_5662,N_5823);
xor U6211 (N_6211,N_5971,N_5779);
nor U6212 (N_6212,N_5534,N_5887);
xor U6213 (N_6213,N_5647,N_5350);
and U6214 (N_6214,N_5879,N_5897);
and U6215 (N_6215,N_5868,N_5311);
or U6216 (N_6216,N_5380,N_5358);
nand U6217 (N_6217,N_5213,N_5125);
and U6218 (N_6218,N_5664,N_5118);
xnor U6219 (N_6219,N_5916,N_5794);
xor U6220 (N_6220,N_5918,N_5718);
nand U6221 (N_6221,N_5832,N_5588);
nor U6222 (N_6222,N_5517,N_5856);
nor U6223 (N_6223,N_5390,N_5807);
or U6224 (N_6224,N_5066,N_5793);
or U6225 (N_6225,N_5923,N_5265);
xnor U6226 (N_6226,N_5681,N_5888);
and U6227 (N_6227,N_5026,N_5529);
or U6228 (N_6228,N_5297,N_5719);
and U6229 (N_6229,N_5996,N_5646);
xnor U6230 (N_6230,N_5568,N_5850);
or U6231 (N_6231,N_5678,N_5953);
xor U6232 (N_6232,N_5321,N_5209);
xnor U6233 (N_6233,N_5618,N_5397);
xnor U6234 (N_6234,N_5825,N_5252);
or U6235 (N_6235,N_5827,N_5820);
xor U6236 (N_6236,N_5544,N_5173);
and U6237 (N_6237,N_5255,N_5964);
nor U6238 (N_6238,N_5137,N_5031);
and U6239 (N_6239,N_5094,N_5979);
or U6240 (N_6240,N_5896,N_5630);
and U6241 (N_6241,N_5217,N_5415);
nor U6242 (N_6242,N_5787,N_5360);
nand U6243 (N_6243,N_5248,N_5861);
nor U6244 (N_6244,N_5463,N_5739);
xnor U6245 (N_6245,N_5600,N_5287);
nor U6246 (N_6246,N_5308,N_5175);
or U6247 (N_6247,N_5477,N_5920);
and U6248 (N_6248,N_5598,N_5750);
nor U6249 (N_6249,N_5314,N_5944);
and U6250 (N_6250,N_5803,N_5906);
nand U6251 (N_6251,N_5230,N_5243);
xor U6252 (N_6252,N_5950,N_5032);
or U6253 (N_6253,N_5376,N_5238);
nand U6254 (N_6254,N_5127,N_5563);
or U6255 (N_6255,N_5328,N_5331);
or U6256 (N_6256,N_5068,N_5777);
or U6257 (N_6257,N_5524,N_5294);
or U6258 (N_6258,N_5035,N_5511);
xnor U6259 (N_6259,N_5955,N_5972);
or U6260 (N_6260,N_5427,N_5990);
and U6261 (N_6261,N_5486,N_5498);
xnor U6262 (N_6262,N_5783,N_5413);
and U6263 (N_6263,N_5023,N_5809);
xor U6264 (N_6264,N_5326,N_5490);
and U6265 (N_6265,N_5191,N_5658);
xor U6266 (N_6266,N_5373,N_5608);
xnor U6267 (N_6267,N_5730,N_5363);
nand U6268 (N_6268,N_5766,N_5420);
nor U6269 (N_6269,N_5208,N_5334);
nor U6270 (N_6270,N_5532,N_5196);
or U6271 (N_6271,N_5126,N_5612);
or U6272 (N_6272,N_5910,N_5615);
nor U6273 (N_6273,N_5058,N_5774);
nor U6274 (N_6274,N_5087,N_5940);
nand U6275 (N_6275,N_5680,N_5198);
xor U6276 (N_6276,N_5212,N_5095);
nand U6277 (N_6277,N_5356,N_5891);
nor U6278 (N_6278,N_5763,N_5768);
and U6279 (N_6279,N_5676,N_5915);
and U6280 (N_6280,N_5860,N_5409);
nand U6281 (N_6281,N_5160,N_5276);
nor U6282 (N_6282,N_5695,N_5622);
xor U6283 (N_6283,N_5892,N_5382);
and U6284 (N_6284,N_5211,N_5353);
nor U6285 (N_6285,N_5813,N_5187);
nor U6286 (N_6286,N_5304,N_5158);
and U6287 (N_6287,N_5737,N_5586);
and U6288 (N_6288,N_5873,N_5949);
nor U6289 (N_6289,N_5997,N_5899);
nor U6290 (N_6290,N_5928,N_5275);
or U6291 (N_6291,N_5926,N_5188);
and U6292 (N_6292,N_5152,N_5659);
or U6293 (N_6293,N_5765,N_5166);
and U6294 (N_6294,N_5253,N_5135);
nor U6295 (N_6295,N_5837,N_5407);
nor U6296 (N_6296,N_5063,N_5256);
nor U6297 (N_6297,N_5870,N_5489);
nor U6298 (N_6298,N_5146,N_5525);
nand U6299 (N_6299,N_5332,N_5573);
or U6300 (N_6300,N_5584,N_5672);
xor U6301 (N_6301,N_5627,N_5488);
or U6302 (N_6302,N_5098,N_5144);
or U6303 (N_6303,N_5590,N_5831);
or U6304 (N_6304,N_5685,N_5476);
or U6305 (N_6305,N_5984,N_5494);
and U6306 (N_6306,N_5077,N_5254);
nand U6307 (N_6307,N_5894,N_5565);
nand U6308 (N_6308,N_5082,N_5131);
xor U6309 (N_6309,N_5853,N_5105);
nand U6310 (N_6310,N_5951,N_5139);
xnor U6311 (N_6311,N_5641,N_5937);
nand U6312 (N_6312,N_5833,N_5399);
nand U6313 (N_6313,N_5509,N_5049);
nor U6314 (N_6314,N_5526,N_5393);
or U6315 (N_6315,N_5702,N_5893);
and U6316 (N_6316,N_5871,N_5099);
and U6317 (N_6317,N_5936,N_5729);
nand U6318 (N_6318,N_5636,N_5323);
xnor U6319 (N_6319,N_5414,N_5527);
nand U6320 (N_6320,N_5849,N_5295);
nor U6321 (N_6321,N_5819,N_5731);
xor U6322 (N_6322,N_5301,N_5101);
and U6323 (N_6323,N_5746,N_5124);
and U6324 (N_6324,N_5073,N_5756);
and U6325 (N_6325,N_5869,N_5624);
and U6326 (N_6326,N_5274,N_5069);
or U6327 (N_6327,N_5140,N_5279);
xor U6328 (N_6328,N_5362,N_5667);
or U6329 (N_6329,N_5947,N_5518);
nor U6330 (N_6330,N_5288,N_5762);
xor U6331 (N_6331,N_5995,N_5974);
nor U6332 (N_6332,N_5011,N_5802);
or U6333 (N_6333,N_5554,N_5114);
nor U6334 (N_6334,N_5402,N_5986);
xnor U6335 (N_6335,N_5113,N_5132);
or U6336 (N_6336,N_5337,N_5878);
nand U6337 (N_6337,N_5660,N_5154);
or U6338 (N_6338,N_5496,N_5968);
nor U6339 (N_6339,N_5535,N_5102);
xor U6340 (N_6340,N_5207,N_5078);
xnor U6341 (N_6341,N_5045,N_5312);
xnor U6342 (N_6342,N_5656,N_5497);
or U6343 (N_6343,N_5815,N_5364);
nand U6344 (N_6344,N_5389,N_5602);
nor U6345 (N_6345,N_5141,N_5239);
nand U6346 (N_6346,N_5867,N_5556);
nand U6347 (N_6347,N_5431,N_5806);
xor U6348 (N_6348,N_5699,N_5033);
nor U6349 (N_6349,N_5085,N_5036);
xor U6350 (N_6350,N_5281,N_5283);
or U6351 (N_6351,N_5694,N_5200);
nand U6352 (N_6352,N_5245,N_5202);
and U6353 (N_6353,N_5733,N_5830);
xor U6354 (N_6354,N_5262,N_5232);
nor U6355 (N_6355,N_5485,N_5019);
or U6356 (N_6356,N_5900,N_5322);
nand U6357 (N_6357,N_5084,N_5805);
nor U6358 (N_6358,N_5454,N_5930);
or U6359 (N_6359,N_5707,N_5079);
xor U6360 (N_6360,N_5109,N_5034);
or U6361 (N_6361,N_5927,N_5343);
or U6362 (N_6362,N_5320,N_5775);
and U6363 (N_6363,N_5148,N_5388);
and U6364 (N_6364,N_5679,N_5723);
or U6365 (N_6365,N_5687,N_5601);
or U6366 (N_6366,N_5566,N_5877);
nor U6367 (N_6367,N_5478,N_5761);
nand U6368 (N_6368,N_5994,N_5952);
and U6369 (N_6369,N_5155,N_5980);
and U6370 (N_6370,N_5318,N_5044);
nor U6371 (N_6371,N_5355,N_5693);
nand U6372 (N_6372,N_5854,N_5796);
xor U6373 (N_6373,N_5438,N_5298);
nand U6374 (N_6374,N_5425,N_5769);
nor U6375 (N_6375,N_5195,N_5302);
nand U6376 (N_6376,N_5835,N_5005);
and U6377 (N_6377,N_5178,N_5493);
nor U6378 (N_6378,N_5421,N_5419);
nor U6379 (N_6379,N_5474,N_5316);
xor U6380 (N_6380,N_5451,N_5799);
or U6381 (N_6381,N_5688,N_5840);
xnor U6382 (N_6382,N_5325,N_5515);
nand U6383 (N_6383,N_5162,N_5842);
and U6384 (N_6384,N_5999,N_5510);
nand U6385 (N_6385,N_5834,N_5205);
or U6386 (N_6386,N_5310,N_5558);
xnor U6387 (N_6387,N_5948,N_5734);
and U6388 (N_6388,N_5669,N_5956);
or U6389 (N_6389,N_5237,N_5973);
or U6390 (N_6390,N_5788,N_5752);
nor U6391 (N_6391,N_5938,N_5901);
and U6392 (N_6392,N_5417,N_5163);
nor U6393 (N_6393,N_5449,N_5633);
nand U6394 (N_6394,N_5599,N_5559);
or U6395 (N_6395,N_5638,N_5505);
xnor U6396 (N_6396,N_5795,N_5567);
nor U6397 (N_6397,N_5300,N_5767);
xor U6398 (N_6398,N_5919,N_5184);
and U6399 (N_6399,N_5941,N_5286);
xnor U6400 (N_6400,N_5670,N_5714);
or U6401 (N_6401,N_5671,N_5715);
or U6402 (N_6402,N_5440,N_5512);
and U6403 (N_6403,N_5942,N_5635);
nand U6404 (N_6404,N_5372,N_5710);
nand U6405 (N_6405,N_5430,N_5824);
nor U6406 (N_6406,N_5176,N_5939);
nor U6407 (N_6407,N_5201,N_5445);
nand U6408 (N_6408,N_5377,N_5408);
and U6409 (N_6409,N_5541,N_5214);
and U6410 (N_6410,N_5480,N_5172);
or U6411 (N_6411,N_5690,N_5720);
and U6412 (N_6412,N_5725,N_5962);
xor U6413 (N_6413,N_5174,N_5668);
and U6414 (N_6414,N_5479,N_5583);
and U6415 (N_6415,N_5542,N_5821);
xnor U6416 (N_6416,N_5933,N_5913);
nor U6417 (N_6417,N_5481,N_5341);
and U6418 (N_6418,N_5704,N_5908);
or U6419 (N_6419,N_5818,N_5504);
and U6420 (N_6420,N_5017,N_5810);
or U6421 (N_6421,N_5180,N_5666);
or U6422 (N_6422,N_5235,N_5516);
or U6423 (N_6423,N_5368,N_5722);
or U6424 (N_6424,N_5654,N_5499);
or U6425 (N_6425,N_5457,N_5596);
xor U6426 (N_6426,N_5164,N_5921);
and U6427 (N_6427,N_5958,N_5024);
nand U6428 (N_6428,N_5089,N_5866);
nand U6429 (N_6429,N_5757,N_5491);
and U6430 (N_6430,N_5484,N_5475);
or U6431 (N_6431,N_5365,N_5885);
nor U6432 (N_6432,N_5258,N_5712);
nor U6433 (N_6433,N_5315,N_5631);
nand U6434 (N_6434,N_5450,N_5018);
or U6435 (N_6435,N_5798,N_5122);
nand U6436 (N_6436,N_5665,N_5220);
nand U6437 (N_6437,N_5740,N_5264);
and U6438 (N_6438,N_5561,N_5500);
and U6439 (N_6439,N_5727,N_5549);
and U6440 (N_6440,N_5981,N_5386);
xor U6441 (N_6441,N_5790,N_5091);
nor U6442 (N_6442,N_5617,N_5620);
nor U6443 (N_6443,N_5396,N_5846);
or U6444 (N_6444,N_5593,N_5351);
xor U6445 (N_6445,N_5537,N_5574);
nand U6446 (N_6446,N_5577,N_5057);
nor U6447 (N_6447,N_5585,N_5041);
nor U6448 (N_6448,N_5296,N_5691);
nand U6449 (N_6449,N_5416,N_5028);
or U6450 (N_6450,N_5225,N_5772);
or U6451 (N_6451,N_5675,N_5008);
or U6452 (N_6452,N_5369,N_5753);
nand U6453 (N_6453,N_5153,N_5786);
xor U6454 (N_6454,N_5000,N_5257);
or U6455 (N_6455,N_5884,N_5233);
and U6456 (N_6456,N_5528,N_5398);
or U6457 (N_6457,N_5855,N_5150);
nand U6458 (N_6458,N_5020,N_5776);
xnor U6459 (N_6459,N_5657,N_5592);
nand U6460 (N_6460,N_5487,N_5378);
or U6461 (N_6461,N_5957,N_5455);
xor U6462 (N_6462,N_5055,N_5609);
and U6463 (N_6463,N_5433,N_5345);
and U6464 (N_6464,N_5536,N_5401);
nand U6465 (N_6465,N_5190,N_5649);
nor U6466 (N_6466,N_5758,N_5473);
or U6467 (N_6467,N_5895,N_5076);
or U6468 (N_6468,N_5280,N_5071);
nand U6469 (N_6469,N_5059,N_5104);
nor U6470 (N_6470,N_5770,N_5437);
or U6471 (N_6471,N_5696,N_5269);
xnor U6472 (N_6472,N_5966,N_5130);
nand U6473 (N_6473,N_5764,N_5792);
or U6474 (N_6474,N_5843,N_5726);
or U6475 (N_6475,N_5875,N_5743);
nor U6476 (N_6476,N_5977,N_5292);
or U6477 (N_6477,N_5808,N_5354);
and U6478 (N_6478,N_5075,N_5935);
nand U6479 (N_6479,N_5848,N_5329);
or U6480 (N_6480,N_5782,N_5167);
xnor U6481 (N_6481,N_5882,N_5181);
or U6482 (N_6482,N_5784,N_5261);
xor U6483 (N_6483,N_5047,N_5708);
xnor U6484 (N_6484,N_5931,N_5724);
nor U6485 (N_6485,N_5836,N_5533);
or U6486 (N_6486,N_5701,N_5759);
xnor U6487 (N_6487,N_5106,N_5097);
nand U6488 (N_6488,N_5482,N_5324);
xor U6489 (N_6489,N_5614,N_5182);
and U6490 (N_6490,N_5013,N_5749);
nand U6491 (N_6491,N_5606,N_5998);
or U6492 (N_6492,N_5339,N_5293);
nand U6493 (N_6493,N_5442,N_5411);
nand U6494 (N_6494,N_5443,N_5418);
or U6495 (N_6495,N_5595,N_5218);
nand U6496 (N_6496,N_5001,N_5744);
nor U6497 (N_6497,N_5222,N_5857);
nand U6498 (N_6498,N_5129,N_5278);
and U6499 (N_6499,N_5742,N_5993);
xor U6500 (N_6500,N_5093,N_5745);
nand U6501 (N_6501,N_5966,N_5572);
and U6502 (N_6502,N_5344,N_5437);
and U6503 (N_6503,N_5520,N_5976);
nor U6504 (N_6504,N_5764,N_5738);
or U6505 (N_6505,N_5769,N_5767);
nor U6506 (N_6506,N_5661,N_5779);
nor U6507 (N_6507,N_5125,N_5751);
xor U6508 (N_6508,N_5050,N_5481);
or U6509 (N_6509,N_5490,N_5470);
xor U6510 (N_6510,N_5001,N_5761);
nor U6511 (N_6511,N_5243,N_5051);
xnor U6512 (N_6512,N_5714,N_5885);
nor U6513 (N_6513,N_5336,N_5873);
nand U6514 (N_6514,N_5157,N_5101);
and U6515 (N_6515,N_5663,N_5694);
and U6516 (N_6516,N_5512,N_5781);
xnor U6517 (N_6517,N_5709,N_5032);
nor U6518 (N_6518,N_5385,N_5350);
xor U6519 (N_6519,N_5721,N_5175);
nand U6520 (N_6520,N_5612,N_5723);
nor U6521 (N_6521,N_5650,N_5126);
or U6522 (N_6522,N_5931,N_5469);
and U6523 (N_6523,N_5816,N_5854);
or U6524 (N_6524,N_5960,N_5384);
nand U6525 (N_6525,N_5804,N_5078);
nand U6526 (N_6526,N_5696,N_5462);
nand U6527 (N_6527,N_5915,N_5111);
nand U6528 (N_6528,N_5882,N_5076);
and U6529 (N_6529,N_5853,N_5511);
xnor U6530 (N_6530,N_5169,N_5084);
nor U6531 (N_6531,N_5719,N_5285);
nor U6532 (N_6532,N_5902,N_5250);
or U6533 (N_6533,N_5572,N_5834);
xor U6534 (N_6534,N_5905,N_5622);
xnor U6535 (N_6535,N_5856,N_5295);
and U6536 (N_6536,N_5700,N_5584);
and U6537 (N_6537,N_5143,N_5059);
nor U6538 (N_6538,N_5090,N_5866);
nor U6539 (N_6539,N_5480,N_5344);
xnor U6540 (N_6540,N_5157,N_5451);
xor U6541 (N_6541,N_5981,N_5345);
or U6542 (N_6542,N_5900,N_5004);
or U6543 (N_6543,N_5581,N_5559);
and U6544 (N_6544,N_5795,N_5529);
or U6545 (N_6545,N_5056,N_5142);
xor U6546 (N_6546,N_5600,N_5146);
nor U6547 (N_6547,N_5495,N_5255);
nand U6548 (N_6548,N_5107,N_5989);
xor U6549 (N_6549,N_5001,N_5462);
xnor U6550 (N_6550,N_5632,N_5113);
or U6551 (N_6551,N_5209,N_5694);
or U6552 (N_6552,N_5832,N_5998);
and U6553 (N_6553,N_5565,N_5294);
and U6554 (N_6554,N_5727,N_5635);
nor U6555 (N_6555,N_5837,N_5523);
and U6556 (N_6556,N_5388,N_5290);
xnor U6557 (N_6557,N_5926,N_5734);
and U6558 (N_6558,N_5663,N_5800);
nand U6559 (N_6559,N_5182,N_5056);
xnor U6560 (N_6560,N_5554,N_5699);
xnor U6561 (N_6561,N_5352,N_5149);
or U6562 (N_6562,N_5222,N_5781);
nor U6563 (N_6563,N_5901,N_5186);
or U6564 (N_6564,N_5683,N_5791);
nor U6565 (N_6565,N_5869,N_5831);
nor U6566 (N_6566,N_5718,N_5006);
xor U6567 (N_6567,N_5953,N_5033);
or U6568 (N_6568,N_5451,N_5556);
nor U6569 (N_6569,N_5013,N_5422);
and U6570 (N_6570,N_5787,N_5808);
and U6571 (N_6571,N_5273,N_5525);
nand U6572 (N_6572,N_5382,N_5463);
and U6573 (N_6573,N_5000,N_5636);
xnor U6574 (N_6574,N_5695,N_5780);
and U6575 (N_6575,N_5203,N_5771);
nand U6576 (N_6576,N_5303,N_5368);
xnor U6577 (N_6577,N_5026,N_5342);
nor U6578 (N_6578,N_5327,N_5331);
or U6579 (N_6579,N_5537,N_5508);
and U6580 (N_6580,N_5536,N_5412);
nor U6581 (N_6581,N_5429,N_5151);
xnor U6582 (N_6582,N_5007,N_5744);
xnor U6583 (N_6583,N_5088,N_5436);
or U6584 (N_6584,N_5486,N_5825);
nor U6585 (N_6585,N_5100,N_5395);
and U6586 (N_6586,N_5363,N_5009);
nor U6587 (N_6587,N_5486,N_5495);
xnor U6588 (N_6588,N_5432,N_5288);
nor U6589 (N_6589,N_5754,N_5405);
nand U6590 (N_6590,N_5118,N_5998);
and U6591 (N_6591,N_5641,N_5607);
nand U6592 (N_6592,N_5759,N_5079);
or U6593 (N_6593,N_5329,N_5330);
nand U6594 (N_6594,N_5314,N_5464);
nand U6595 (N_6595,N_5559,N_5230);
and U6596 (N_6596,N_5933,N_5675);
or U6597 (N_6597,N_5831,N_5947);
and U6598 (N_6598,N_5904,N_5795);
nand U6599 (N_6599,N_5553,N_5195);
nor U6600 (N_6600,N_5996,N_5187);
nor U6601 (N_6601,N_5624,N_5172);
nor U6602 (N_6602,N_5569,N_5374);
xor U6603 (N_6603,N_5170,N_5171);
or U6604 (N_6604,N_5281,N_5968);
nand U6605 (N_6605,N_5629,N_5559);
and U6606 (N_6606,N_5334,N_5302);
xor U6607 (N_6607,N_5696,N_5940);
or U6608 (N_6608,N_5204,N_5691);
or U6609 (N_6609,N_5698,N_5562);
and U6610 (N_6610,N_5940,N_5057);
nand U6611 (N_6611,N_5351,N_5953);
nand U6612 (N_6612,N_5473,N_5872);
or U6613 (N_6613,N_5792,N_5622);
and U6614 (N_6614,N_5045,N_5152);
nand U6615 (N_6615,N_5127,N_5411);
xnor U6616 (N_6616,N_5430,N_5570);
nor U6617 (N_6617,N_5106,N_5907);
or U6618 (N_6618,N_5743,N_5936);
nand U6619 (N_6619,N_5468,N_5117);
and U6620 (N_6620,N_5101,N_5349);
and U6621 (N_6621,N_5541,N_5075);
or U6622 (N_6622,N_5553,N_5365);
xnor U6623 (N_6623,N_5763,N_5849);
xnor U6624 (N_6624,N_5599,N_5294);
nor U6625 (N_6625,N_5920,N_5170);
and U6626 (N_6626,N_5495,N_5030);
nand U6627 (N_6627,N_5832,N_5084);
and U6628 (N_6628,N_5196,N_5378);
nand U6629 (N_6629,N_5146,N_5397);
or U6630 (N_6630,N_5563,N_5290);
nand U6631 (N_6631,N_5677,N_5733);
and U6632 (N_6632,N_5913,N_5428);
nor U6633 (N_6633,N_5867,N_5828);
nand U6634 (N_6634,N_5916,N_5750);
and U6635 (N_6635,N_5037,N_5531);
or U6636 (N_6636,N_5289,N_5331);
nor U6637 (N_6637,N_5726,N_5093);
nand U6638 (N_6638,N_5572,N_5683);
nand U6639 (N_6639,N_5829,N_5690);
nand U6640 (N_6640,N_5721,N_5555);
and U6641 (N_6641,N_5344,N_5246);
nor U6642 (N_6642,N_5518,N_5012);
or U6643 (N_6643,N_5183,N_5532);
xnor U6644 (N_6644,N_5817,N_5693);
nand U6645 (N_6645,N_5293,N_5375);
or U6646 (N_6646,N_5549,N_5320);
nand U6647 (N_6647,N_5504,N_5957);
nand U6648 (N_6648,N_5156,N_5692);
nand U6649 (N_6649,N_5985,N_5821);
and U6650 (N_6650,N_5382,N_5587);
or U6651 (N_6651,N_5952,N_5172);
nand U6652 (N_6652,N_5293,N_5385);
xor U6653 (N_6653,N_5746,N_5668);
xnor U6654 (N_6654,N_5128,N_5175);
nand U6655 (N_6655,N_5873,N_5422);
xor U6656 (N_6656,N_5551,N_5792);
or U6657 (N_6657,N_5039,N_5458);
nor U6658 (N_6658,N_5303,N_5107);
xor U6659 (N_6659,N_5702,N_5953);
nor U6660 (N_6660,N_5421,N_5788);
xor U6661 (N_6661,N_5971,N_5626);
nand U6662 (N_6662,N_5575,N_5381);
or U6663 (N_6663,N_5066,N_5992);
nor U6664 (N_6664,N_5126,N_5266);
nor U6665 (N_6665,N_5623,N_5969);
nor U6666 (N_6666,N_5295,N_5363);
or U6667 (N_6667,N_5691,N_5290);
or U6668 (N_6668,N_5274,N_5624);
and U6669 (N_6669,N_5308,N_5715);
or U6670 (N_6670,N_5837,N_5106);
or U6671 (N_6671,N_5060,N_5346);
and U6672 (N_6672,N_5055,N_5791);
and U6673 (N_6673,N_5687,N_5500);
or U6674 (N_6674,N_5382,N_5240);
nor U6675 (N_6675,N_5806,N_5101);
and U6676 (N_6676,N_5681,N_5243);
nor U6677 (N_6677,N_5071,N_5761);
or U6678 (N_6678,N_5428,N_5188);
and U6679 (N_6679,N_5266,N_5302);
nand U6680 (N_6680,N_5535,N_5889);
or U6681 (N_6681,N_5607,N_5086);
and U6682 (N_6682,N_5460,N_5027);
xnor U6683 (N_6683,N_5507,N_5791);
nand U6684 (N_6684,N_5733,N_5611);
nand U6685 (N_6685,N_5253,N_5145);
xor U6686 (N_6686,N_5399,N_5806);
or U6687 (N_6687,N_5501,N_5415);
and U6688 (N_6688,N_5292,N_5714);
nand U6689 (N_6689,N_5064,N_5348);
nand U6690 (N_6690,N_5127,N_5593);
xnor U6691 (N_6691,N_5343,N_5971);
xnor U6692 (N_6692,N_5093,N_5502);
nor U6693 (N_6693,N_5309,N_5243);
xor U6694 (N_6694,N_5772,N_5483);
nor U6695 (N_6695,N_5716,N_5547);
and U6696 (N_6696,N_5781,N_5390);
nor U6697 (N_6697,N_5979,N_5228);
nor U6698 (N_6698,N_5365,N_5112);
nor U6699 (N_6699,N_5788,N_5794);
and U6700 (N_6700,N_5190,N_5626);
nand U6701 (N_6701,N_5973,N_5748);
and U6702 (N_6702,N_5477,N_5210);
and U6703 (N_6703,N_5018,N_5012);
and U6704 (N_6704,N_5595,N_5121);
and U6705 (N_6705,N_5571,N_5083);
or U6706 (N_6706,N_5038,N_5996);
and U6707 (N_6707,N_5467,N_5305);
xor U6708 (N_6708,N_5363,N_5081);
or U6709 (N_6709,N_5756,N_5295);
nand U6710 (N_6710,N_5621,N_5695);
nor U6711 (N_6711,N_5745,N_5359);
and U6712 (N_6712,N_5529,N_5958);
and U6713 (N_6713,N_5155,N_5116);
nor U6714 (N_6714,N_5385,N_5253);
and U6715 (N_6715,N_5543,N_5625);
nand U6716 (N_6716,N_5680,N_5788);
nor U6717 (N_6717,N_5542,N_5985);
and U6718 (N_6718,N_5296,N_5545);
nand U6719 (N_6719,N_5818,N_5302);
or U6720 (N_6720,N_5729,N_5040);
and U6721 (N_6721,N_5160,N_5552);
and U6722 (N_6722,N_5686,N_5204);
or U6723 (N_6723,N_5632,N_5652);
and U6724 (N_6724,N_5220,N_5060);
or U6725 (N_6725,N_5184,N_5078);
nand U6726 (N_6726,N_5596,N_5714);
or U6727 (N_6727,N_5930,N_5256);
nor U6728 (N_6728,N_5825,N_5410);
or U6729 (N_6729,N_5352,N_5638);
or U6730 (N_6730,N_5499,N_5743);
xnor U6731 (N_6731,N_5463,N_5599);
xnor U6732 (N_6732,N_5258,N_5842);
and U6733 (N_6733,N_5507,N_5159);
xnor U6734 (N_6734,N_5024,N_5020);
nor U6735 (N_6735,N_5835,N_5532);
and U6736 (N_6736,N_5085,N_5960);
xor U6737 (N_6737,N_5710,N_5887);
and U6738 (N_6738,N_5133,N_5669);
or U6739 (N_6739,N_5304,N_5330);
xor U6740 (N_6740,N_5076,N_5086);
and U6741 (N_6741,N_5762,N_5305);
and U6742 (N_6742,N_5285,N_5615);
and U6743 (N_6743,N_5746,N_5529);
xor U6744 (N_6744,N_5246,N_5408);
nor U6745 (N_6745,N_5047,N_5678);
nor U6746 (N_6746,N_5162,N_5837);
nand U6747 (N_6747,N_5248,N_5237);
nor U6748 (N_6748,N_5496,N_5340);
xor U6749 (N_6749,N_5634,N_5528);
xor U6750 (N_6750,N_5103,N_5724);
nor U6751 (N_6751,N_5118,N_5425);
or U6752 (N_6752,N_5946,N_5637);
and U6753 (N_6753,N_5979,N_5348);
or U6754 (N_6754,N_5654,N_5509);
and U6755 (N_6755,N_5652,N_5198);
and U6756 (N_6756,N_5488,N_5685);
nor U6757 (N_6757,N_5205,N_5030);
nor U6758 (N_6758,N_5157,N_5417);
nand U6759 (N_6759,N_5853,N_5572);
and U6760 (N_6760,N_5474,N_5138);
and U6761 (N_6761,N_5379,N_5071);
nor U6762 (N_6762,N_5681,N_5870);
or U6763 (N_6763,N_5398,N_5913);
nor U6764 (N_6764,N_5605,N_5748);
xor U6765 (N_6765,N_5790,N_5541);
xnor U6766 (N_6766,N_5084,N_5326);
and U6767 (N_6767,N_5036,N_5860);
and U6768 (N_6768,N_5183,N_5483);
or U6769 (N_6769,N_5767,N_5412);
nand U6770 (N_6770,N_5747,N_5770);
xnor U6771 (N_6771,N_5402,N_5915);
nand U6772 (N_6772,N_5589,N_5421);
or U6773 (N_6773,N_5906,N_5215);
or U6774 (N_6774,N_5851,N_5378);
nor U6775 (N_6775,N_5279,N_5647);
or U6776 (N_6776,N_5961,N_5491);
xnor U6777 (N_6777,N_5381,N_5396);
nand U6778 (N_6778,N_5922,N_5771);
nor U6779 (N_6779,N_5041,N_5141);
or U6780 (N_6780,N_5832,N_5052);
and U6781 (N_6781,N_5418,N_5964);
xnor U6782 (N_6782,N_5104,N_5701);
nor U6783 (N_6783,N_5751,N_5519);
and U6784 (N_6784,N_5950,N_5491);
xnor U6785 (N_6785,N_5958,N_5472);
nor U6786 (N_6786,N_5293,N_5206);
or U6787 (N_6787,N_5241,N_5029);
nor U6788 (N_6788,N_5732,N_5795);
and U6789 (N_6789,N_5103,N_5079);
or U6790 (N_6790,N_5156,N_5041);
xor U6791 (N_6791,N_5933,N_5947);
xnor U6792 (N_6792,N_5549,N_5486);
nand U6793 (N_6793,N_5389,N_5055);
or U6794 (N_6794,N_5343,N_5152);
nand U6795 (N_6795,N_5134,N_5351);
or U6796 (N_6796,N_5767,N_5993);
nand U6797 (N_6797,N_5284,N_5330);
and U6798 (N_6798,N_5080,N_5099);
nand U6799 (N_6799,N_5586,N_5174);
or U6800 (N_6800,N_5194,N_5216);
or U6801 (N_6801,N_5702,N_5275);
and U6802 (N_6802,N_5212,N_5774);
nor U6803 (N_6803,N_5640,N_5869);
or U6804 (N_6804,N_5691,N_5520);
xnor U6805 (N_6805,N_5775,N_5358);
or U6806 (N_6806,N_5923,N_5397);
nand U6807 (N_6807,N_5621,N_5311);
nand U6808 (N_6808,N_5284,N_5212);
or U6809 (N_6809,N_5096,N_5648);
nor U6810 (N_6810,N_5480,N_5984);
nand U6811 (N_6811,N_5402,N_5916);
and U6812 (N_6812,N_5679,N_5269);
nor U6813 (N_6813,N_5106,N_5789);
nor U6814 (N_6814,N_5095,N_5747);
nor U6815 (N_6815,N_5554,N_5901);
nand U6816 (N_6816,N_5360,N_5290);
and U6817 (N_6817,N_5335,N_5690);
nor U6818 (N_6818,N_5962,N_5643);
nor U6819 (N_6819,N_5016,N_5395);
and U6820 (N_6820,N_5947,N_5585);
or U6821 (N_6821,N_5945,N_5247);
nor U6822 (N_6822,N_5846,N_5618);
nand U6823 (N_6823,N_5082,N_5150);
nor U6824 (N_6824,N_5979,N_5851);
nor U6825 (N_6825,N_5815,N_5784);
xnor U6826 (N_6826,N_5174,N_5166);
and U6827 (N_6827,N_5276,N_5659);
and U6828 (N_6828,N_5331,N_5089);
nand U6829 (N_6829,N_5640,N_5668);
xnor U6830 (N_6830,N_5712,N_5453);
xor U6831 (N_6831,N_5899,N_5261);
or U6832 (N_6832,N_5305,N_5667);
nand U6833 (N_6833,N_5999,N_5179);
nand U6834 (N_6834,N_5145,N_5307);
xor U6835 (N_6835,N_5634,N_5665);
and U6836 (N_6836,N_5831,N_5753);
and U6837 (N_6837,N_5434,N_5572);
nor U6838 (N_6838,N_5884,N_5761);
and U6839 (N_6839,N_5823,N_5565);
nand U6840 (N_6840,N_5716,N_5088);
or U6841 (N_6841,N_5830,N_5753);
nand U6842 (N_6842,N_5265,N_5488);
or U6843 (N_6843,N_5648,N_5856);
xor U6844 (N_6844,N_5636,N_5767);
nor U6845 (N_6845,N_5662,N_5582);
nand U6846 (N_6846,N_5110,N_5022);
nor U6847 (N_6847,N_5834,N_5357);
or U6848 (N_6848,N_5969,N_5410);
and U6849 (N_6849,N_5696,N_5420);
nor U6850 (N_6850,N_5349,N_5731);
and U6851 (N_6851,N_5908,N_5877);
xor U6852 (N_6852,N_5289,N_5524);
nand U6853 (N_6853,N_5092,N_5553);
nand U6854 (N_6854,N_5974,N_5398);
and U6855 (N_6855,N_5628,N_5424);
nand U6856 (N_6856,N_5654,N_5319);
or U6857 (N_6857,N_5644,N_5603);
or U6858 (N_6858,N_5906,N_5820);
and U6859 (N_6859,N_5040,N_5778);
xor U6860 (N_6860,N_5751,N_5429);
or U6861 (N_6861,N_5760,N_5979);
and U6862 (N_6862,N_5313,N_5054);
nor U6863 (N_6863,N_5695,N_5647);
xnor U6864 (N_6864,N_5949,N_5226);
nand U6865 (N_6865,N_5157,N_5791);
or U6866 (N_6866,N_5160,N_5038);
xor U6867 (N_6867,N_5778,N_5454);
nor U6868 (N_6868,N_5314,N_5879);
nor U6869 (N_6869,N_5766,N_5644);
and U6870 (N_6870,N_5699,N_5762);
nand U6871 (N_6871,N_5683,N_5856);
or U6872 (N_6872,N_5018,N_5679);
or U6873 (N_6873,N_5776,N_5262);
nand U6874 (N_6874,N_5938,N_5659);
and U6875 (N_6875,N_5972,N_5724);
or U6876 (N_6876,N_5770,N_5823);
and U6877 (N_6877,N_5661,N_5969);
or U6878 (N_6878,N_5364,N_5996);
and U6879 (N_6879,N_5062,N_5753);
or U6880 (N_6880,N_5418,N_5888);
xnor U6881 (N_6881,N_5220,N_5276);
or U6882 (N_6882,N_5058,N_5391);
nor U6883 (N_6883,N_5507,N_5122);
and U6884 (N_6884,N_5314,N_5818);
xnor U6885 (N_6885,N_5213,N_5277);
and U6886 (N_6886,N_5009,N_5666);
nand U6887 (N_6887,N_5781,N_5786);
and U6888 (N_6888,N_5786,N_5697);
nand U6889 (N_6889,N_5952,N_5701);
and U6890 (N_6890,N_5278,N_5205);
and U6891 (N_6891,N_5064,N_5171);
nand U6892 (N_6892,N_5779,N_5773);
xnor U6893 (N_6893,N_5937,N_5755);
nor U6894 (N_6894,N_5273,N_5957);
nor U6895 (N_6895,N_5816,N_5794);
and U6896 (N_6896,N_5579,N_5631);
xnor U6897 (N_6897,N_5653,N_5485);
nor U6898 (N_6898,N_5585,N_5811);
xnor U6899 (N_6899,N_5597,N_5124);
nor U6900 (N_6900,N_5180,N_5108);
or U6901 (N_6901,N_5586,N_5141);
xor U6902 (N_6902,N_5917,N_5515);
or U6903 (N_6903,N_5515,N_5343);
nor U6904 (N_6904,N_5570,N_5577);
nand U6905 (N_6905,N_5010,N_5194);
and U6906 (N_6906,N_5830,N_5373);
and U6907 (N_6907,N_5470,N_5746);
and U6908 (N_6908,N_5509,N_5095);
nor U6909 (N_6909,N_5619,N_5685);
or U6910 (N_6910,N_5210,N_5205);
nor U6911 (N_6911,N_5397,N_5601);
and U6912 (N_6912,N_5838,N_5802);
xor U6913 (N_6913,N_5664,N_5325);
xor U6914 (N_6914,N_5847,N_5906);
or U6915 (N_6915,N_5683,N_5385);
xor U6916 (N_6916,N_5678,N_5022);
or U6917 (N_6917,N_5809,N_5669);
nand U6918 (N_6918,N_5219,N_5643);
or U6919 (N_6919,N_5341,N_5589);
nand U6920 (N_6920,N_5573,N_5927);
nand U6921 (N_6921,N_5569,N_5369);
or U6922 (N_6922,N_5599,N_5234);
xnor U6923 (N_6923,N_5837,N_5604);
nor U6924 (N_6924,N_5769,N_5900);
nor U6925 (N_6925,N_5265,N_5900);
or U6926 (N_6926,N_5824,N_5259);
nor U6927 (N_6927,N_5671,N_5830);
xnor U6928 (N_6928,N_5625,N_5513);
and U6929 (N_6929,N_5067,N_5593);
nand U6930 (N_6930,N_5081,N_5393);
nand U6931 (N_6931,N_5143,N_5530);
xnor U6932 (N_6932,N_5027,N_5048);
nand U6933 (N_6933,N_5488,N_5774);
nand U6934 (N_6934,N_5547,N_5305);
nor U6935 (N_6935,N_5444,N_5047);
or U6936 (N_6936,N_5016,N_5739);
and U6937 (N_6937,N_5610,N_5717);
xor U6938 (N_6938,N_5790,N_5127);
and U6939 (N_6939,N_5529,N_5351);
or U6940 (N_6940,N_5986,N_5405);
nor U6941 (N_6941,N_5926,N_5523);
or U6942 (N_6942,N_5661,N_5457);
or U6943 (N_6943,N_5381,N_5659);
nor U6944 (N_6944,N_5567,N_5306);
and U6945 (N_6945,N_5173,N_5061);
nand U6946 (N_6946,N_5787,N_5784);
or U6947 (N_6947,N_5537,N_5470);
nand U6948 (N_6948,N_5975,N_5625);
and U6949 (N_6949,N_5663,N_5674);
and U6950 (N_6950,N_5492,N_5845);
nand U6951 (N_6951,N_5535,N_5504);
and U6952 (N_6952,N_5858,N_5712);
xor U6953 (N_6953,N_5258,N_5984);
nor U6954 (N_6954,N_5775,N_5065);
xnor U6955 (N_6955,N_5763,N_5876);
nor U6956 (N_6956,N_5833,N_5713);
nor U6957 (N_6957,N_5017,N_5574);
nand U6958 (N_6958,N_5579,N_5113);
and U6959 (N_6959,N_5381,N_5253);
xnor U6960 (N_6960,N_5529,N_5408);
and U6961 (N_6961,N_5119,N_5488);
and U6962 (N_6962,N_5764,N_5082);
xnor U6963 (N_6963,N_5485,N_5994);
xor U6964 (N_6964,N_5357,N_5345);
nand U6965 (N_6965,N_5750,N_5051);
and U6966 (N_6966,N_5121,N_5794);
and U6967 (N_6967,N_5733,N_5863);
or U6968 (N_6968,N_5433,N_5095);
nand U6969 (N_6969,N_5189,N_5315);
nand U6970 (N_6970,N_5396,N_5725);
or U6971 (N_6971,N_5873,N_5679);
and U6972 (N_6972,N_5900,N_5348);
nor U6973 (N_6973,N_5789,N_5583);
and U6974 (N_6974,N_5324,N_5240);
and U6975 (N_6975,N_5110,N_5042);
nand U6976 (N_6976,N_5028,N_5532);
or U6977 (N_6977,N_5890,N_5212);
xnor U6978 (N_6978,N_5373,N_5346);
nand U6979 (N_6979,N_5537,N_5512);
and U6980 (N_6980,N_5704,N_5423);
nor U6981 (N_6981,N_5537,N_5414);
xor U6982 (N_6982,N_5320,N_5400);
nand U6983 (N_6983,N_5287,N_5626);
xor U6984 (N_6984,N_5761,N_5208);
or U6985 (N_6985,N_5460,N_5386);
nor U6986 (N_6986,N_5696,N_5113);
nand U6987 (N_6987,N_5974,N_5273);
or U6988 (N_6988,N_5531,N_5034);
nor U6989 (N_6989,N_5341,N_5330);
or U6990 (N_6990,N_5778,N_5589);
and U6991 (N_6991,N_5978,N_5828);
nand U6992 (N_6992,N_5166,N_5097);
and U6993 (N_6993,N_5756,N_5635);
and U6994 (N_6994,N_5832,N_5529);
and U6995 (N_6995,N_5396,N_5806);
and U6996 (N_6996,N_5354,N_5646);
xnor U6997 (N_6997,N_5275,N_5601);
or U6998 (N_6998,N_5715,N_5599);
and U6999 (N_6999,N_5405,N_5672);
nor U7000 (N_7000,N_6720,N_6846);
or U7001 (N_7001,N_6913,N_6831);
nand U7002 (N_7002,N_6791,N_6361);
or U7003 (N_7003,N_6341,N_6350);
xnor U7004 (N_7004,N_6596,N_6251);
xor U7005 (N_7005,N_6542,N_6051);
and U7006 (N_7006,N_6351,N_6144);
and U7007 (N_7007,N_6332,N_6110);
nor U7008 (N_7008,N_6628,N_6207);
and U7009 (N_7009,N_6632,N_6359);
or U7010 (N_7010,N_6132,N_6022);
nand U7011 (N_7011,N_6787,N_6533);
or U7012 (N_7012,N_6122,N_6045);
or U7013 (N_7013,N_6824,N_6299);
nor U7014 (N_7014,N_6433,N_6007);
nor U7015 (N_7015,N_6293,N_6891);
nor U7016 (N_7016,N_6668,N_6038);
nand U7017 (N_7017,N_6130,N_6300);
or U7018 (N_7018,N_6924,N_6977);
or U7019 (N_7019,N_6642,N_6855);
nor U7020 (N_7020,N_6111,N_6645);
xnor U7021 (N_7021,N_6555,N_6626);
nor U7022 (N_7022,N_6428,N_6362);
and U7023 (N_7023,N_6700,N_6690);
xor U7024 (N_7024,N_6035,N_6616);
xnor U7025 (N_7025,N_6313,N_6658);
or U7026 (N_7026,N_6286,N_6452);
and U7027 (N_7027,N_6121,N_6274);
or U7028 (N_7028,N_6379,N_6602);
and U7029 (N_7029,N_6931,N_6517);
or U7030 (N_7030,N_6972,N_6674);
nand U7031 (N_7031,N_6442,N_6735);
xor U7032 (N_7032,N_6413,N_6613);
or U7033 (N_7033,N_6146,N_6763);
nor U7034 (N_7034,N_6211,N_6687);
and U7035 (N_7035,N_6507,N_6488);
and U7036 (N_7036,N_6443,N_6863);
nor U7037 (N_7037,N_6744,N_6354);
and U7038 (N_7038,N_6834,N_6388);
and U7039 (N_7039,N_6518,N_6582);
nor U7040 (N_7040,N_6089,N_6896);
and U7041 (N_7041,N_6468,N_6346);
and U7042 (N_7042,N_6136,N_6218);
or U7043 (N_7043,N_6194,N_6727);
or U7044 (N_7044,N_6106,N_6941);
or U7045 (N_7045,N_6323,N_6385);
xor U7046 (N_7046,N_6027,N_6798);
xor U7047 (N_7047,N_6775,N_6307);
nor U7048 (N_7048,N_6963,N_6394);
xnor U7049 (N_7049,N_6571,N_6656);
xor U7050 (N_7050,N_6589,N_6568);
and U7051 (N_7051,N_6813,N_6137);
or U7052 (N_7052,N_6092,N_6415);
nor U7053 (N_7053,N_6115,N_6508);
and U7054 (N_7054,N_6303,N_6636);
xnor U7055 (N_7055,N_6965,N_6856);
nor U7056 (N_7056,N_6746,N_6393);
or U7057 (N_7057,N_6012,N_6193);
xnor U7058 (N_7058,N_6473,N_6812);
and U7059 (N_7059,N_6779,N_6356);
xnor U7060 (N_7060,N_6527,N_6974);
nand U7061 (N_7061,N_6531,N_6205);
and U7062 (N_7062,N_6565,N_6061);
nor U7063 (N_7063,N_6734,N_6246);
or U7064 (N_7064,N_6139,N_6434);
nor U7065 (N_7065,N_6033,N_6869);
or U7066 (N_7066,N_6269,N_6681);
or U7067 (N_7067,N_6366,N_6789);
xnor U7068 (N_7068,N_6826,N_6900);
xor U7069 (N_7069,N_6496,N_6664);
nor U7070 (N_7070,N_6797,N_6920);
or U7071 (N_7071,N_6322,N_6657);
and U7072 (N_7072,N_6058,N_6255);
nor U7073 (N_7073,N_6243,N_6551);
and U7074 (N_7074,N_6843,N_6231);
nand U7075 (N_7075,N_6738,N_6444);
nor U7076 (N_7076,N_6942,N_6208);
nand U7077 (N_7077,N_6295,N_6037);
xor U7078 (N_7078,N_6561,N_6807);
nor U7079 (N_7079,N_6588,N_6436);
nand U7080 (N_7080,N_6701,N_6279);
xnor U7081 (N_7081,N_6695,N_6864);
or U7082 (N_7082,N_6074,N_6823);
or U7083 (N_7083,N_6161,N_6730);
or U7084 (N_7084,N_6320,N_6182);
nor U7085 (N_7085,N_6649,N_6513);
nor U7086 (N_7086,N_6405,N_6921);
or U7087 (N_7087,N_6721,N_6955);
and U7088 (N_7088,N_6326,N_6857);
and U7089 (N_7089,N_6710,N_6395);
and U7090 (N_7090,N_6104,N_6774);
and U7091 (N_7091,N_6248,N_6036);
and U7092 (N_7092,N_6160,N_6138);
nand U7093 (N_7093,N_6992,N_6062);
and U7094 (N_7094,N_6788,N_6277);
nand U7095 (N_7095,N_6926,N_6123);
and U7096 (N_7096,N_6708,N_6666);
or U7097 (N_7097,N_6672,N_6052);
and U7098 (N_7098,N_6151,N_6566);
and U7099 (N_7099,N_6185,N_6770);
and U7100 (N_7100,N_6732,N_6001);
nor U7101 (N_7101,N_6619,N_6796);
or U7102 (N_7102,N_6614,N_6576);
or U7103 (N_7103,N_6853,N_6098);
or U7104 (N_7104,N_6819,N_6705);
and U7105 (N_7105,N_6731,N_6166);
or U7106 (N_7106,N_6252,N_6986);
and U7107 (N_7107,N_6489,N_6239);
nor U7108 (N_7108,N_6564,N_6538);
nand U7109 (N_7109,N_6479,N_6431);
or U7110 (N_7110,N_6919,N_6486);
nand U7111 (N_7111,N_6552,N_6319);
xnor U7112 (N_7112,N_6686,N_6877);
nand U7113 (N_7113,N_6522,N_6673);
or U7114 (N_7114,N_6094,N_6450);
nand U7115 (N_7115,N_6832,N_6339);
xor U7116 (N_7116,N_6102,N_6932);
xor U7117 (N_7117,N_6321,N_6806);
nand U7118 (N_7118,N_6310,N_6155);
nor U7119 (N_7119,N_6056,N_6401);
and U7120 (N_7120,N_6594,N_6641);
or U7121 (N_7121,N_6271,N_6344);
nor U7122 (N_7122,N_6331,N_6739);
and U7123 (N_7123,N_6375,N_6737);
nand U7124 (N_7124,N_6383,N_6934);
nand U7125 (N_7125,N_6912,N_6541);
or U7126 (N_7126,N_6838,N_6276);
and U7127 (N_7127,N_6068,N_6667);
xor U7128 (N_7128,N_6624,N_6814);
nand U7129 (N_7129,N_6964,N_6048);
xor U7130 (N_7130,N_6962,N_6836);
nand U7131 (N_7131,N_6778,N_6606);
xnor U7132 (N_7132,N_6726,N_6790);
and U7133 (N_7133,N_6783,N_6281);
xnor U7134 (N_7134,N_6993,N_6935);
and U7135 (N_7135,N_6483,N_6029);
xor U7136 (N_7136,N_6879,N_6675);
xnor U7137 (N_7137,N_6335,N_6163);
xnor U7138 (N_7138,N_6860,N_6506);
nand U7139 (N_7139,N_6190,N_6915);
and U7140 (N_7140,N_6071,N_6124);
nand U7141 (N_7141,N_6010,N_6605);
or U7142 (N_7142,N_6352,N_6376);
xor U7143 (N_7143,N_6192,N_6426);
xnor U7144 (N_7144,N_6117,N_6861);
nand U7145 (N_7145,N_6928,N_6917);
or U7146 (N_7146,N_6006,N_6471);
nand U7147 (N_7147,N_6600,N_6020);
and U7148 (N_7148,N_6250,N_6463);
nor U7149 (N_7149,N_6460,N_6887);
xor U7150 (N_7150,N_6096,N_6355);
nor U7151 (N_7151,N_6911,N_6189);
nand U7152 (N_7152,N_6262,N_6294);
xor U7153 (N_7153,N_6125,N_6345);
or U7154 (N_7154,N_6475,N_6546);
and U7155 (N_7155,N_6736,N_6892);
or U7156 (N_7156,N_6100,N_6607);
and U7157 (N_7157,N_6521,N_6429);
nand U7158 (N_7158,N_6617,N_6549);
xor U7159 (N_7159,N_6631,N_6618);
nand U7160 (N_7160,N_6063,N_6023);
nand U7161 (N_7161,N_6268,N_6871);
and U7162 (N_7162,N_6229,N_6118);
nand U7163 (N_7163,N_6478,N_6536);
nor U7164 (N_7164,N_6044,N_6398);
nor U7165 (N_7165,N_6402,N_6186);
nand U7166 (N_7166,N_6773,N_6256);
nor U7167 (N_7167,N_6927,N_6752);
nand U7168 (N_7168,N_6729,N_6984);
nor U7169 (N_7169,N_6692,N_6119);
nor U7170 (N_7170,N_6457,N_6309);
or U7171 (N_7171,N_6922,N_6622);
nor U7172 (N_7172,N_6704,N_6698);
nand U7173 (N_7173,N_6408,N_6755);
nor U7174 (N_7174,N_6906,N_6373);
nor U7175 (N_7175,N_6584,N_6390);
nor U7176 (N_7176,N_6446,N_6711);
xnor U7177 (N_7177,N_6011,N_6867);
nor U7178 (N_7178,N_6502,N_6004);
nand U7179 (N_7179,N_6159,N_6199);
nor U7180 (N_7180,N_6213,N_6849);
nand U7181 (N_7181,N_6358,N_6973);
or U7182 (N_7182,N_6372,N_6179);
xnor U7183 (N_7183,N_6227,N_6216);
and U7184 (N_7184,N_6265,N_6670);
nand U7185 (N_7185,N_6273,N_6156);
and U7186 (N_7186,N_6215,N_6031);
or U7187 (N_7187,N_6623,N_6289);
and U7188 (N_7188,N_6655,N_6261);
and U7189 (N_7189,N_6423,N_6528);
or U7190 (N_7190,N_6235,N_6610);
nor U7191 (N_7191,N_6621,N_6537);
xor U7192 (N_7192,N_6590,N_6712);
or U7193 (N_7193,N_6377,N_6706);
or U7194 (N_7194,N_6923,N_6938);
nand U7195 (N_7195,N_6747,N_6237);
xor U7196 (N_7196,N_6439,N_6282);
xnor U7197 (N_7197,N_6585,N_6175);
nand U7198 (N_7198,N_6288,N_6693);
xor U7199 (N_7199,N_6456,N_6363);
and U7200 (N_7200,N_6386,N_6197);
nand U7201 (N_7201,N_6238,N_6753);
and U7202 (N_7202,N_6794,N_6868);
nor U7203 (N_7203,N_6709,N_6142);
nand U7204 (N_7204,N_6847,N_6421);
nor U7205 (N_7205,N_6153,N_6954);
and U7206 (N_7206,N_6441,N_6776);
nor U7207 (N_7207,N_6573,N_6080);
or U7208 (N_7208,N_6002,N_6490);
and U7209 (N_7209,N_6660,N_6095);
nand U7210 (N_7210,N_6497,N_6420);
nand U7211 (N_7211,N_6976,N_6487);
and U7212 (N_7212,N_6512,N_6263);
or U7213 (N_7213,N_6957,N_6172);
and U7214 (N_7214,N_6563,N_6760);
nand U7215 (N_7215,N_6154,N_6325);
nor U7216 (N_7216,N_6406,N_6226);
xor U7217 (N_7217,N_6220,N_6648);
xnor U7218 (N_7218,N_6018,N_6762);
or U7219 (N_7219,N_6644,N_6560);
nor U7220 (N_7220,N_6685,N_6067);
or U7221 (N_7221,N_6874,N_6543);
nand U7222 (N_7222,N_6757,N_6422);
nand U7223 (N_7223,N_6811,N_6480);
xnor U7224 (N_7224,N_6329,N_6075);
nand U7225 (N_7225,N_6839,N_6223);
xnor U7226 (N_7226,N_6054,N_6167);
nor U7227 (N_7227,N_6983,N_6411);
or U7228 (N_7228,N_6653,N_6597);
xnor U7229 (N_7229,N_6761,N_6691);
nor U7230 (N_7230,N_6131,N_6903);
and U7231 (N_7231,N_6472,N_6574);
nand U7232 (N_7232,N_6825,N_6244);
nand U7233 (N_7233,N_6754,N_6909);
xnor U7234 (N_7234,N_6516,N_6640);
nand U7235 (N_7235,N_6540,N_6716);
nor U7236 (N_7236,N_6076,N_6050);
nor U7237 (N_7237,N_6509,N_6599);
xnor U7238 (N_7238,N_6224,N_6534);
xor U7239 (N_7239,N_6206,N_6247);
or U7240 (N_7240,N_6859,N_6404);
or U7241 (N_7241,N_6786,N_6535);
or U7242 (N_7242,N_6127,N_6759);
xnor U7243 (N_7243,N_6116,N_6053);
nor U7244 (N_7244,N_6365,N_6870);
and U7245 (N_7245,N_6980,N_6128);
and U7246 (N_7246,N_6914,N_6875);
or U7247 (N_7247,N_6852,N_6481);
nor U7248 (N_7248,N_6635,N_6009);
nor U7249 (N_7249,N_6382,N_6399);
nor U7250 (N_7250,N_6975,N_6267);
nand U7251 (N_7251,N_6799,N_6049);
nor U7252 (N_7252,N_6659,N_6093);
nand U7253 (N_7253,N_6815,N_6445);
nor U7254 (N_7254,N_6895,N_6925);
nand U7255 (N_7255,N_6283,N_6069);
nor U7256 (N_7256,N_6270,N_6232);
nor U7257 (N_7257,N_6781,N_6995);
and U7258 (N_7258,N_6165,N_6043);
and U7259 (N_7259,N_6897,N_6634);
xnor U7260 (N_7260,N_6024,N_6055);
nand U7261 (N_7261,N_6264,N_6242);
or U7262 (N_7262,N_6530,N_6217);
or U7263 (N_7263,N_6148,N_6134);
or U7264 (N_7264,N_6407,N_6461);
and U7265 (N_7265,N_6866,N_6629);
or U7266 (N_7266,N_6403,N_6081);
and U7267 (N_7267,N_6397,N_6550);
nor U7268 (N_7268,N_6065,N_6090);
and U7269 (N_7269,N_6818,N_6898);
or U7270 (N_7270,N_6240,N_6097);
and U7271 (N_7271,N_6703,N_6143);
or U7272 (N_7272,N_6586,N_6643);
and U7273 (N_7273,N_6418,N_6800);
xnor U7274 (N_7274,N_6005,N_6661);
xor U7275 (N_7275,N_6201,N_6633);
nand U7276 (N_7276,N_6357,N_6713);
or U7277 (N_7277,N_6158,N_6078);
or U7278 (N_7278,N_6449,N_6476);
and U7279 (N_7279,N_6349,N_6946);
nor U7280 (N_7280,N_6990,N_6105);
xnor U7281 (N_7281,N_6525,N_6079);
nand U7282 (N_7282,N_6292,N_6082);
or U7283 (N_7283,N_6996,N_6682);
nor U7284 (N_7284,N_6066,N_6702);
or U7285 (N_7285,N_6647,N_6750);
xnor U7286 (N_7286,N_6455,N_6598);
xor U7287 (N_7287,N_6370,N_6652);
xnor U7288 (N_7288,N_6991,N_6611);
and U7289 (N_7289,N_6196,N_6278);
nor U7290 (N_7290,N_6440,N_6503);
or U7291 (N_7291,N_6529,N_6494);
nand U7292 (N_7292,N_6872,N_6854);
xor U7293 (N_7293,N_6195,N_6340);
xnor U7294 (N_7294,N_6748,N_6949);
and U7295 (N_7295,N_6830,N_6287);
nand U7296 (N_7296,N_6767,N_6181);
nor U7297 (N_7297,N_6336,N_6907);
or U7298 (N_7298,N_6378,N_6228);
or U7299 (N_7299,N_6184,N_6929);
or U7300 (N_7300,N_6677,N_6200);
nor U7301 (N_7301,N_6878,N_6368);
and U7302 (N_7302,N_6047,N_6459);
or U7303 (N_7303,N_6858,N_6221);
or U7304 (N_7304,N_6465,N_6432);
nand U7305 (N_7305,N_6948,N_6724);
nor U7306 (N_7306,N_6367,N_6464);
or U7307 (N_7307,N_6091,N_6389);
nand U7308 (N_7308,N_6936,N_6723);
and U7309 (N_7309,N_6451,N_6554);
nor U7310 (N_7310,N_6837,N_6639);
and U7311 (N_7311,N_6572,N_6141);
xnor U7312 (N_7312,N_6930,N_6944);
nor U7313 (N_7313,N_6176,N_6482);
nand U7314 (N_7314,N_6678,N_6337);
xor U7315 (N_7315,N_6808,N_6654);
nand U7316 (N_7316,N_6514,N_6501);
nand U7317 (N_7317,N_6524,N_6257);
nand U7318 (N_7318,N_6173,N_6174);
xor U7319 (N_7319,N_6202,N_6785);
and U7320 (N_7320,N_6844,N_6017);
or U7321 (N_7321,N_6343,N_6694);
xor U7322 (N_7322,N_6330,N_6827);
nand U7323 (N_7323,N_6328,N_6427);
and U7324 (N_7324,N_6725,N_6064);
nor U7325 (N_7325,N_6802,N_6316);
and U7326 (N_7326,N_6742,N_6684);
or U7327 (N_7327,N_6569,N_6591);
and U7328 (N_7328,N_6046,N_6608);
nand U7329 (N_7329,N_6880,N_6595);
or U7330 (N_7330,N_6437,N_6214);
xnor U7331 (N_7331,N_6493,N_6212);
nand U7332 (N_7332,N_6638,N_6249);
nand U7333 (N_7333,N_6109,N_6970);
xnor U7334 (N_7334,N_6696,N_6520);
xnor U7335 (N_7335,N_6780,N_6910);
and U7336 (N_7336,N_6665,N_6312);
nand U7337 (N_7337,N_6342,N_6414);
and U7338 (N_7338,N_6901,N_6768);
xnor U7339 (N_7339,N_6581,N_6885);
nand U7340 (N_7340,N_6371,N_6301);
or U7341 (N_7341,N_6219,N_6210);
and U7342 (N_7342,N_6557,N_6318);
xnor U7343 (N_7343,N_6679,N_6733);
nand U7344 (N_7344,N_6989,N_6162);
xnor U7345 (N_7345,N_6107,N_6556);
nand U7346 (N_7346,N_6865,N_6412);
xnor U7347 (N_7347,N_6689,N_6553);
or U7348 (N_7348,N_6032,N_6805);
or U7349 (N_7349,N_6766,N_6454);
or U7350 (N_7350,N_6756,N_6937);
and U7351 (N_7351,N_6578,N_6391);
or U7352 (N_7352,N_6236,N_6987);
and U7353 (N_7353,N_6149,N_6466);
nand U7354 (N_7354,N_6374,N_6315);
and U7355 (N_7355,N_6245,N_6302);
xnor U7356 (N_7356,N_6745,N_6952);
nand U7357 (N_7357,N_6950,N_6592);
nand U7358 (N_7358,N_6191,N_6177);
xnor U7359 (N_7359,N_6577,N_6504);
and U7360 (N_7360,N_6112,N_6458);
nor U7361 (N_7361,N_6353,N_6088);
nand U7362 (N_7362,N_6842,N_6751);
and U7363 (N_7363,N_6669,N_6904);
and U7364 (N_7364,N_6209,N_6147);
nand U7365 (N_7365,N_6547,N_6234);
and U7366 (N_7366,N_6334,N_6615);
and U7367 (N_7367,N_6500,N_6894);
nand U7368 (N_7368,N_6792,N_6025);
xor U7369 (N_7369,N_6609,N_6170);
xnor U7370 (N_7370,N_6728,N_6492);
nand U7371 (N_7371,N_6835,N_6961);
nor U7372 (N_7372,N_6416,N_6150);
nor U7373 (N_7373,N_6718,N_6722);
nand U7374 (N_7374,N_6967,N_6782);
nand U7375 (N_7375,N_6933,N_6801);
nand U7376 (N_7376,N_6129,N_6960);
xor U7377 (N_7377,N_6495,N_6381);
or U7378 (N_7378,N_6662,N_6485);
nor U7379 (N_7379,N_6308,N_6804);
nand U7380 (N_7380,N_6663,N_6275);
nor U7381 (N_7381,N_6491,N_6715);
xor U7382 (N_7382,N_6559,N_6544);
and U7383 (N_7383,N_6028,N_6510);
nand U7384 (N_7384,N_6650,N_6997);
or U7385 (N_7385,N_6523,N_6285);
and U7386 (N_7386,N_6126,N_6298);
nor U7387 (N_7387,N_6570,N_6364);
xnor U7388 (N_7388,N_6347,N_6099);
xnor U7389 (N_7389,N_6630,N_6998);
and U7390 (N_7390,N_6086,N_6016);
xnor U7391 (N_7391,N_6168,N_6306);
xor U7392 (N_7392,N_6180,N_6034);
or U7393 (N_7393,N_6575,N_6470);
xnor U7394 (N_7394,N_6916,N_6042);
and U7395 (N_7395,N_6140,N_6258);
and U7396 (N_7396,N_6430,N_6969);
nand U7397 (N_7397,N_6327,N_6966);
or U7398 (N_7398,N_6030,N_6646);
xnor U7399 (N_7399,N_6988,N_6956);
xnor U7400 (N_7400,N_6765,N_6676);
nor U7401 (N_7401,N_6828,N_6070);
nand U7402 (N_7402,N_6060,N_6338);
nor U7403 (N_7403,N_6881,N_6810);
nor U7404 (N_7404,N_6448,N_6526);
nor U7405 (N_7405,N_6417,N_6953);
xnor U7406 (N_7406,N_6821,N_6719);
and U7407 (N_7407,N_6820,N_6021);
nand U7408 (N_7408,N_6886,N_6968);
nand U7409 (N_7409,N_6157,N_6841);
nand U7410 (N_7410,N_6587,N_6171);
nand U7411 (N_7411,N_6848,N_6410);
nand U7412 (N_7412,N_6850,N_6462);
nor U7413 (N_7413,N_6084,N_6816);
xor U7414 (N_7414,N_6183,N_6583);
nor U7415 (N_7415,N_6749,N_6829);
nand U7416 (N_7416,N_6333,N_6519);
xor U7417 (N_7417,N_6499,N_6254);
xor U7418 (N_7418,N_6041,N_6073);
or U7419 (N_7419,N_6113,N_6101);
nand U7420 (N_7420,N_6851,N_6680);
nand U7421 (N_7421,N_6994,N_6057);
and U7422 (N_7422,N_6889,N_6688);
nor U7423 (N_7423,N_6873,N_6883);
xnor U7424 (N_7424,N_6999,N_6888);
and U7425 (N_7425,N_6884,N_6260);
and U7426 (N_7426,N_6943,N_6072);
or U7427 (N_7427,N_6438,N_6699);
or U7428 (N_7428,N_6822,N_6424);
nor U7429 (N_7429,N_6793,N_6671);
nor U7430 (N_7430,N_6620,N_6515);
and U7431 (N_7431,N_6697,N_6169);
nor U7432 (N_7432,N_6777,N_6707);
or U7433 (N_7433,N_6284,N_6324);
xor U7434 (N_7434,N_6133,N_6548);
xor U7435 (N_7435,N_6203,N_6593);
or U7436 (N_7436,N_6817,N_6120);
or U7437 (N_7437,N_6266,N_6369);
or U7438 (N_7438,N_6259,N_6425);
and U7439 (N_7439,N_6135,N_6803);
nand U7440 (N_7440,N_6795,N_6601);
xor U7441 (N_7441,N_6862,N_6114);
and U7442 (N_7442,N_6103,N_6603);
nor U7443 (N_7443,N_6380,N_6474);
nand U7444 (N_7444,N_6290,N_6178);
or U7445 (N_7445,N_6145,N_6304);
or U7446 (N_7446,N_6840,N_6769);
xor U7447 (N_7447,N_6469,N_6253);
or U7448 (N_7448,N_6740,N_6348);
and U7449 (N_7449,N_6511,N_6225);
nor U7450 (N_7450,N_6280,N_6291);
and U7451 (N_7451,N_6579,N_6958);
xor U7452 (N_7452,N_6562,N_6453);
nand U7453 (N_7453,N_6083,N_6008);
or U7454 (N_7454,N_6845,N_6040);
nand U7455 (N_7455,N_6940,N_6204);
nand U7456 (N_7456,N_6311,N_6771);
and U7457 (N_7457,N_6477,N_6059);
or U7458 (N_7458,N_6890,N_6939);
and U7459 (N_7459,N_6188,N_6314);
nand U7460 (N_7460,N_6683,N_6400);
nand U7461 (N_7461,N_6545,N_6532);
and U7462 (N_7462,N_6013,N_6003);
xor U7463 (N_7463,N_6435,N_6971);
nor U7464 (N_7464,N_6447,N_6498);
nor U7465 (N_7465,N_6714,N_6085);
nand U7466 (N_7466,N_6959,N_6882);
xnor U7467 (N_7467,N_6539,N_6272);
nand U7468 (N_7468,N_6741,N_6982);
nor U7469 (N_7469,N_6039,N_6077);
nor U7470 (N_7470,N_6360,N_6000);
or U7471 (N_7471,N_6876,N_6164);
nor U7472 (N_7472,N_6019,N_6384);
xnor U7473 (N_7473,N_6558,N_6580);
or U7474 (N_7474,N_6612,N_6743);
xnor U7475 (N_7475,N_6625,N_6409);
xnor U7476 (N_7476,N_6305,N_6981);
xnor U7477 (N_7477,N_6947,N_6978);
nand U7478 (N_7478,N_6604,N_6809);
and U7479 (N_7479,N_6152,N_6784);
xnor U7480 (N_7480,N_6758,N_6908);
nor U7481 (N_7481,N_6717,N_6764);
xnor U7482 (N_7482,N_6187,N_6396);
or U7483 (N_7483,N_6015,N_6979);
and U7484 (N_7484,N_6902,N_6297);
nor U7485 (N_7485,N_6985,N_6893);
xnor U7486 (N_7486,N_6087,N_6108);
nor U7487 (N_7487,N_6419,N_6296);
nand U7488 (N_7488,N_6918,N_6637);
nand U7489 (N_7489,N_6651,N_6233);
or U7490 (N_7490,N_6772,N_6198);
xor U7491 (N_7491,N_6026,N_6241);
and U7492 (N_7492,N_6230,N_6951);
nand U7493 (N_7493,N_6222,N_6899);
and U7494 (N_7494,N_6833,N_6317);
nand U7495 (N_7495,N_6905,N_6567);
nand U7496 (N_7496,N_6627,N_6467);
or U7497 (N_7497,N_6392,N_6945);
nor U7498 (N_7498,N_6484,N_6387);
and U7499 (N_7499,N_6505,N_6014);
or U7500 (N_7500,N_6668,N_6111);
nor U7501 (N_7501,N_6197,N_6794);
and U7502 (N_7502,N_6595,N_6128);
and U7503 (N_7503,N_6056,N_6005);
or U7504 (N_7504,N_6486,N_6656);
nand U7505 (N_7505,N_6829,N_6922);
and U7506 (N_7506,N_6963,N_6641);
and U7507 (N_7507,N_6167,N_6966);
and U7508 (N_7508,N_6176,N_6420);
nand U7509 (N_7509,N_6894,N_6890);
and U7510 (N_7510,N_6232,N_6848);
nand U7511 (N_7511,N_6460,N_6926);
or U7512 (N_7512,N_6012,N_6957);
xnor U7513 (N_7513,N_6250,N_6666);
xnor U7514 (N_7514,N_6150,N_6016);
nor U7515 (N_7515,N_6399,N_6200);
nor U7516 (N_7516,N_6330,N_6811);
and U7517 (N_7517,N_6330,N_6900);
xor U7518 (N_7518,N_6421,N_6947);
nor U7519 (N_7519,N_6066,N_6980);
nor U7520 (N_7520,N_6773,N_6407);
nand U7521 (N_7521,N_6856,N_6474);
or U7522 (N_7522,N_6305,N_6376);
nand U7523 (N_7523,N_6402,N_6888);
xnor U7524 (N_7524,N_6091,N_6848);
or U7525 (N_7525,N_6032,N_6218);
nor U7526 (N_7526,N_6797,N_6239);
and U7527 (N_7527,N_6360,N_6549);
nand U7528 (N_7528,N_6400,N_6990);
and U7529 (N_7529,N_6925,N_6585);
xnor U7530 (N_7530,N_6933,N_6414);
xor U7531 (N_7531,N_6186,N_6780);
and U7532 (N_7532,N_6795,N_6428);
and U7533 (N_7533,N_6586,N_6778);
or U7534 (N_7534,N_6972,N_6346);
and U7535 (N_7535,N_6987,N_6285);
or U7536 (N_7536,N_6303,N_6392);
nand U7537 (N_7537,N_6817,N_6705);
xnor U7538 (N_7538,N_6061,N_6015);
or U7539 (N_7539,N_6455,N_6737);
nand U7540 (N_7540,N_6196,N_6496);
nor U7541 (N_7541,N_6062,N_6659);
nor U7542 (N_7542,N_6272,N_6990);
nor U7543 (N_7543,N_6716,N_6379);
nor U7544 (N_7544,N_6913,N_6968);
and U7545 (N_7545,N_6224,N_6778);
or U7546 (N_7546,N_6312,N_6571);
and U7547 (N_7547,N_6579,N_6087);
or U7548 (N_7548,N_6212,N_6046);
nand U7549 (N_7549,N_6541,N_6127);
xnor U7550 (N_7550,N_6471,N_6510);
nand U7551 (N_7551,N_6145,N_6575);
or U7552 (N_7552,N_6428,N_6194);
xor U7553 (N_7553,N_6841,N_6183);
nor U7554 (N_7554,N_6651,N_6325);
nand U7555 (N_7555,N_6936,N_6482);
nor U7556 (N_7556,N_6431,N_6393);
xnor U7557 (N_7557,N_6492,N_6474);
or U7558 (N_7558,N_6741,N_6221);
and U7559 (N_7559,N_6793,N_6496);
nor U7560 (N_7560,N_6432,N_6466);
xnor U7561 (N_7561,N_6951,N_6404);
xnor U7562 (N_7562,N_6133,N_6420);
xor U7563 (N_7563,N_6914,N_6476);
or U7564 (N_7564,N_6901,N_6566);
nor U7565 (N_7565,N_6490,N_6421);
and U7566 (N_7566,N_6245,N_6103);
xor U7567 (N_7567,N_6570,N_6460);
xor U7568 (N_7568,N_6600,N_6628);
nand U7569 (N_7569,N_6035,N_6454);
xnor U7570 (N_7570,N_6786,N_6686);
nand U7571 (N_7571,N_6808,N_6294);
nand U7572 (N_7572,N_6139,N_6907);
nor U7573 (N_7573,N_6124,N_6306);
nand U7574 (N_7574,N_6698,N_6222);
xor U7575 (N_7575,N_6851,N_6235);
xnor U7576 (N_7576,N_6158,N_6096);
nand U7577 (N_7577,N_6527,N_6850);
and U7578 (N_7578,N_6058,N_6505);
or U7579 (N_7579,N_6572,N_6421);
nor U7580 (N_7580,N_6032,N_6894);
nor U7581 (N_7581,N_6981,N_6061);
or U7582 (N_7582,N_6787,N_6355);
nor U7583 (N_7583,N_6120,N_6523);
or U7584 (N_7584,N_6043,N_6871);
nor U7585 (N_7585,N_6591,N_6949);
nand U7586 (N_7586,N_6613,N_6564);
nor U7587 (N_7587,N_6852,N_6198);
nor U7588 (N_7588,N_6349,N_6922);
nor U7589 (N_7589,N_6925,N_6214);
or U7590 (N_7590,N_6318,N_6641);
nand U7591 (N_7591,N_6539,N_6746);
and U7592 (N_7592,N_6513,N_6111);
nand U7593 (N_7593,N_6394,N_6771);
or U7594 (N_7594,N_6425,N_6136);
and U7595 (N_7595,N_6045,N_6310);
nand U7596 (N_7596,N_6017,N_6327);
xor U7597 (N_7597,N_6027,N_6119);
nor U7598 (N_7598,N_6586,N_6974);
nand U7599 (N_7599,N_6398,N_6920);
and U7600 (N_7600,N_6086,N_6064);
or U7601 (N_7601,N_6948,N_6491);
and U7602 (N_7602,N_6872,N_6865);
nand U7603 (N_7603,N_6331,N_6559);
xor U7604 (N_7604,N_6596,N_6797);
xor U7605 (N_7605,N_6724,N_6733);
nand U7606 (N_7606,N_6357,N_6941);
and U7607 (N_7607,N_6104,N_6997);
and U7608 (N_7608,N_6843,N_6610);
nand U7609 (N_7609,N_6520,N_6416);
nand U7610 (N_7610,N_6967,N_6932);
xor U7611 (N_7611,N_6173,N_6320);
nor U7612 (N_7612,N_6760,N_6344);
and U7613 (N_7613,N_6660,N_6040);
nor U7614 (N_7614,N_6628,N_6921);
nand U7615 (N_7615,N_6395,N_6873);
and U7616 (N_7616,N_6635,N_6057);
xnor U7617 (N_7617,N_6797,N_6712);
nor U7618 (N_7618,N_6450,N_6825);
and U7619 (N_7619,N_6076,N_6795);
xnor U7620 (N_7620,N_6598,N_6860);
nor U7621 (N_7621,N_6171,N_6971);
and U7622 (N_7622,N_6673,N_6837);
nor U7623 (N_7623,N_6742,N_6169);
and U7624 (N_7624,N_6587,N_6134);
and U7625 (N_7625,N_6670,N_6047);
and U7626 (N_7626,N_6085,N_6000);
nor U7627 (N_7627,N_6198,N_6161);
nand U7628 (N_7628,N_6291,N_6066);
and U7629 (N_7629,N_6423,N_6956);
and U7630 (N_7630,N_6727,N_6020);
or U7631 (N_7631,N_6002,N_6403);
nor U7632 (N_7632,N_6550,N_6449);
or U7633 (N_7633,N_6612,N_6631);
or U7634 (N_7634,N_6777,N_6068);
and U7635 (N_7635,N_6349,N_6182);
nor U7636 (N_7636,N_6517,N_6224);
xnor U7637 (N_7637,N_6990,N_6570);
nand U7638 (N_7638,N_6199,N_6530);
nor U7639 (N_7639,N_6374,N_6443);
xnor U7640 (N_7640,N_6493,N_6204);
or U7641 (N_7641,N_6394,N_6477);
or U7642 (N_7642,N_6185,N_6664);
nand U7643 (N_7643,N_6471,N_6850);
and U7644 (N_7644,N_6589,N_6368);
or U7645 (N_7645,N_6386,N_6137);
and U7646 (N_7646,N_6892,N_6303);
xnor U7647 (N_7647,N_6049,N_6157);
and U7648 (N_7648,N_6700,N_6084);
nand U7649 (N_7649,N_6984,N_6588);
nand U7650 (N_7650,N_6571,N_6833);
nor U7651 (N_7651,N_6665,N_6846);
or U7652 (N_7652,N_6643,N_6613);
nor U7653 (N_7653,N_6761,N_6423);
or U7654 (N_7654,N_6517,N_6868);
xnor U7655 (N_7655,N_6794,N_6648);
nor U7656 (N_7656,N_6758,N_6999);
xnor U7657 (N_7657,N_6929,N_6933);
or U7658 (N_7658,N_6874,N_6408);
xor U7659 (N_7659,N_6936,N_6779);
nand U7660 (N_7660,N_6106,N_6984);
and U7661 (N_7661,N_6376,N_6225);
or U7662 (N_7662,N_6357,N_6642);
and U7663 (N_7663,N_6886,N_6787);
nand U7664 (N_7664,N_6074,N_6049);
xor U7665 (N_7665,N_6470,N_6280);
nand U7666 (N_7666,N_6844,N_6559);
or U7667 (N_7667,N_6489,N_6856);
xnor U7668 (N_7668,N_6117,N_6114);
or U7669 (N_7669,N_6648,N_6928);
and U7670 (N_7670,N_6899,N_6718);
and U7671 (N_7671,N_6517,N_6700);
nor U7672 (N_7672,N_6812,N_6715);
nand U7673 (N_7673,N_6478,N_6113);
xnor U7674 (N_7674,N_6773,N_6489);
and U7675 (N_7675,N_6859,N_6482);
or U7676 (N_7676,N_6832,N_6911);
xnor U7677 (N_7677,N_6950,N_6183);
and U7678 (N_7678,N_6205,N_6251);
nand U7679 (N_7679,N_6811,N_6665);
nand U7680 (N_7680,N_6930,N_6640);
or U7681 (N_7681,N_6505,N_6089);
xor U7682 (N_7682,N_6251,N_6419);
nor U7683 (N_7683,N_6518,N_6551);
xor U7684 (N_7684,N_6665,N_6676);
and U7685 (N_7685,N_6651,N_6400);
or U7686 (N_7686,N_6550,N_6952);
and U7687 (N_7687,N_6246,N_6876);
xor U7688 (N_7688,N_6511,N_6840);
or U7689 (N_7689,N_6880,N_6075);
or U7690 (N_7690,N_6587,N_6994);
nand U7691 (N_7691,N_6708,N_6816);
or U7692 (N_7692,N_6606,N_6542);
nand U7693 (N_7693,N_6632,N_6465);
and U7694 (N_7694,N_6119,N_6505);
and U7695 (N_7695,N_6953,N_6582);
nand U7696 (N_7696,N_6856,N_6720);
nor U7697 (N_7697,N_6654,N_6407);
nor U7698 (N_7698,N_6773,N_6565);
nor U7699 (N_7699,N_6231,N_6102);
or U7700 (N_7700,N_6015,N_6385);
and U7701 (N_7701,N_6407,N_6418);
or U7702 (N_7702,N_6885,N_6795);
nor U7703 (N_7703,N_6895,N_6547);
xor U7704 (N_7704,N_6697,N_6956);
nor U7705 (N_7705,N_6765,N_6857);
xor U7706 (N_7706,N_6636,N_6068);
or U7707 (N_7707,N_6160,N_6596);
and U7708 (N_7708,N_6202,N_6052);
nor U7709 (N_7709,N_6655,N_6441);
and U7710 (N_7710,N_6429,N_6399);
nor U7711 (N_7711,N_6386,N_6588);
nor U7712 (N_7712,N_6390,N_6030);
nor U7713 (N_7713,N_6829,N_6496);
or U7714 (N_7714,N_6737,N_6524);
or U7715 (N_7715,N_6382,N_6935);
xnor U7716 (N_7716,N_6280,N_6136);
xor U7717 (N_7717,N_6562,N_6768);
xnor U7718 (N_7718,N_6076,N_6208);
or U7719 (N_7719,N_6601,N_6405);
nand U7720 (N_7720,N_6606,N_6703);
or U7721 (N_7721,N_6742,N_6774);
and U7722 (N_7722,N_6057,N_6210);
xor U7723 (N_7723,N_6054,N_6567);
xnor U7724 (N_7724,N_6960,N_6953);
nand U7725 (N_7725,N_6971,N_6878);
nand U7726 (N_7726,N_6486,N_6304);
or U7727 (N_7727,N_6792,N_6920);
nand U7728 (N_7728,N_6854,N_6950);
nor U7729 (N_7729,N_6766,N_6511);
or U7730 (N_7730,N_6090,N_6441);
xor U7731 (N_7731,N_6314,N_6840);
xor U7732 (N_7732,N_6916,N_6068);
nor U7733 (N_7733,N_6329,N_6619);
xor U7734 (N_7734,N_6062,N_6801);
nand U7735 (N_7735,N_6987,N_6185);
or U7736 (N_7736,N_6324,N_6587);
and U7737 (N_7737,N_6412,N_6921);
or U7738 (N_7738,N_6429,N_6379);
and U7739 (N_7739,N_6874,N_6831);
and U7740 (N_7740,N_6375,N_6837);
nand U7741 (N_7741,N_6529,N_6993);
xnor U7742 (N_7742,N_6342,N_6805);
xnor U7743 (N_7743,N_6969,N_6957);
xnor U7744 (N_7744,N_6491,N_6008);
xor U7745 (N_7745,N_6978,N_6130);
xor U7746 (N_7746,N_6266,N_6598);
nor U7747 (N_7747,N_6205,N_6354);
nor U7748 (N_7748,N_6630,N_6442);
xnor U7749 (N_7749,N_6710,N_6200);
nor U7750 (N_7750,N_6049,N_6655);
or U7751 (N_7751,N_6362,N_6590);
nor U7752 (N_7752,N_6297,N_6478);
nor U7753 (N_7753,N_6490,N_6948);
or U7754 (N_7754,N_6989,N_6533);
xor U7755 (N_7755,N_6468,N_6428);
nand U7756 (N_7756,N_6986,N_6245);
and U7757 (N_7757,N_6633,N_6329);
nand U7758 (N_7758,N_6343,N_6137);
nor U7759 (N_7759,N_6833,N_6344);
and U7760 (N_7760,N_6920,N_6362);
nor U7761 (N_7761,N_6502,N_6946);
nor U7762 (N_7762,N_6531,N_6625);
nand U7763 (N_7763,N_6498,N_6493);
or U7764 (N_7764,N_6564,N_6737);
nor U7765 (N_7765,N_6102,N_6968);
xor U7766 (N_7766,N_6831,N_6384);
xor U7767 (N_7767,N_6971,N_6358);
nor U7768 (N_7768,N_6636,N_6402);
or U7769 (N_7769,N_6660,N_6168);
xor U7770 (N_7770,N_6995,N_6108);
nor U7771 (N_7771,N_6432,N_6544);
or U7772 (N_7772,N_6780,N_6816);
or U7773 (N_7773,N_6189,N_6526);
xor U7774 (N_7774,N_6413,N_6344);
and U7775 (N_7775,N_6071,N_6933);
and U7776 (N_7776,N_6668,N_6813);
nand U7777 (N_7777,N_6111,N_6103);
xnor U7778 (N_7778,N_6061,N_6035);
xnor U7779 (N_7779,N_6473,N_6943);
nand U7780 (N_7780,N_6634,N_6273);
nand U7781 (N_7781,N_6959,N_6220);
nor U7782 (N_7782,N_6220,N_6708);
and U7783 (N_7783,N_6047,N_6867);
xnor U7784 (N_7784,N_6895,N_6606);
xnor U7785 (N_7785,N_6008,N_6776);
nand U7786 (N_7786,N_6890,N_6108);
nor U7787 (N_7787,N_6138,N_6389);
nor U7788 (N_7788,N_6545,N_6718);
xnor U7789 (N_7789,N_6725,N_6516);
nor U7790 (N_7790,N_6257,N_6412);
or U7791 (N_7791,N_6198,N_6494);
xor U7792 (N_7792,N_6427,N_6846);
xnor U7793 (N_7793,N_6632,N_6449);
nor U7794 (N_7794,N_6627,N_6670);
or U7795 (N_7795,N_6431,N_6633);
xor U7796 (N_7796,N_6628,N_6002);
or U7797 (N_7797,N_6944,N_6675);
nand U7798 (N_7798,N_6755,N_6784);
and U7799 (N_7799,N_6946,N_6168);
nand U7800 (N_7800,N_6376,N_6280);
xnor U7801 (N_7801,N_6710,N_6732);
and U7802 (N_7802,N_6377,N_6659);
nor U7803 (N_7803,N_6984,N_6426);
nand U7804 (N_7804,N_6679,N_6128);
xnor U7805 (N_7805,N_6801,N_6085);
xnor U7806 (N_7806,N_6978,N_6779);
or U7807 (N_7807,N_6509,N_6847);
or U7808 (N_7808,N_6382,N_6719);
nand U7809 (N_7809,N_6251,N_6176);
nor U7810 (N_7810,N_6570,N_6040);
nand U7811 (N_7811,N_6140,N_6735);
nor U7812 (N_7812,N_6576,N_6321);
and U7813 (N_7813,N_6525,N_6278);
nor U7814 (N_7814,N_6882,N_6057);
and U7815 (N_7815,N_6622,N_6664);
or U7816 (N_7816,N_6535,N_6079);
or U7817 (N_7817,N_6692,N_6859);
or U7818 (N_7818,N_6585,N_6359);
nand U7819 (N_7819,N_6694,N_6793);
nand U7820 (N_7820,N_6078,N_6509);
nor U7821 (N_7821,N_6707,N_6494);
or U7822 (N_7822,N_6211,N_6561);
and U7823 (N_7823,N_6732,N_6922);
nor U7824 (N_7824,N_6365,N_6842);
nand U7825 (N_7825,N_6209,N_6087);
xor U7826 (N_7826,N_6391,N_6048);
or U7827 (N_7827,N_6425,N_6815);
or U7828 (N_7828,N_6740,N_6252);
and U7829 (N_7829,N_6968,N_6491);
and U7830 (N_7830,N_6356,N_6624);
nand U7831 (N_7831,N_6476,N_6875);
xnor U7832 (N_7832,N_6778,N_6117);
xor U7833 (N_7833,N_6464,N_6816);
and U7834 (N_7834,N_6330,N_6427);
and U7835 (N_7835,N_6225,N_6276);
or U7836 (N_7836,N_6357,N_6666);
nand U7837 (N_7837,N_6387,N_6630);
or U7838 (N_7838,N_6806,N_6062);
nor U7839 (N_7839,N_6611,N_6875);
xor U7840 (N_7840,N_6584,N_6261);
xnor U7841 (N_7841,N_6450,N_6521);
xor U7842 (N_7842,N_6890,N_6060);
nor U7843 (N_7843,N_6748,N_6738);
xor U7844 (N_7844,N_6021,N_6517);
nand U7845 (N_7845,N_6285,N_6379);
xnor U7846 (N_7846,N_6742,N_6156);
xnor U7847 (N_7847,N_6913,N_6496);
or U7848 (N_7848,N_6996,N_6984);
or U7849 (N_7849,N_6823,N_6995);
and U7850 (N_7850,N_6235,N_6745);
xnor U7851 (N_7851,N_6207,N_6668);
or U7852 (N_7852,N_6386,N_6370);
nand U7853 (N_7853,N_6887,N_6326);
or U7854 (N_7854,N_6683,N_6374);
nor U7855 (N_7855,N_6473,N_6666);
and U7856 (N_7856,N_6682,N_6397);
nor U7857 (N_7857,N_6592,N_6100);
xnor U7858 (N_7858,N_6836,N_6631);
and U7859 (N_7859,N_6277,N_6238);
or U7860 (N_7860,N_6245,N_6223);
and U7861 (N_7861,N_6960,N_6673);
nor U7862 (N_7862,N_6585,N_6864);
xor U7863 (N_7863,N_6316,N_6966);
and U7864 (N_7864,N_6776,N_6106);
xor U7865 (N_7865,N_6496,N_6819);
nor U7866 (N_7866,N_6396,N_6890);
nor U7867 (N_7867,N_6549,N_6766);
and U7868 (N_7868,N_6037,N_6594);
nor U7869 (N_7869,N_6938,N_6551);
nand U7870 (N_7870,N_6477,N_6312);
and U7871 (N_7871,N_6074,N_6335);
nand U7872 (N_7872,N_6331,N_6757);
and U7873 (N_7873,N_6915,N_6442);
xor U7874 (N_7874,N_6011,N_6876);
nor U7875 (N_7875,N_6224,N_6022);
nor U7876 (N_7876,N_6736,N_6061);
nand U7877 (N_7877,N_6026,N_6275);
xor U7878 (N_7878,N_6003,N_6350);
nor U7879 (N_7879,N_6878,N_6295);
nand U7880 (N_7880,N_6684,N_6930);
nor U7881 (N_7881,N_6886,N_6458);
and U7882 (N_7882,N_6988,N_6767);
and U7883 (N_7883,N_6000,N_6309);
nor U7884 (N_7884,N_6823,N_6482);
nand U7885 (N_7885,N_6817,N_6030);
nand U7886 (N_7886,N_6143,N_6126);
or U7887 (N_7887,N_6839,N_6104);
and U7888 (N_7888,N_6197,N_6656);
and U7889 (N_7889,N_6212,N_6482);
nand U7890 (N_7890,N_6684,N_6457);
nand U7891 (N_7891,N_6091,N_6511);
nor U7892 (N_7892,N_6006,N_6159);
and U7893 (N_7893,N_6142,N_6533);
xnor U7894 (N_7894,N_6989,N_6715);
nand U7895 (N_7895,N_6958,N_6897);
or U7896 (N_7896,N_6469,N_6278);
and U7897 (N_7897,N_6120,N_6263);
or U7898 (N_7898,N_6007,N_6659);
xnor U7899 (N_7899,N_6648,N_6545);
nand U7900 (N_7900,N_6506,N_6192);
xor U7901 (N_7901,N_6655,N_6728);
nand U7902 (N_7902,N_6386,N_6218);
xor U7903 (N_7903,N_6366,N_6871);
nand U7904 (N_7904,N_6043,N_6349);
and U7905 (N_7905,N_6830,N_6192);
nor U7906 (N_7906,N_6926,N_6246);
and U7907 (N_7907,N_6052,N_6824);
nor U7908 (N_7908,N_6114,N_6442);
and U7909 (N_7909,N_6703,N_6921);
and U7910 (N_7910,N_6942,N_6145);
xor U7911 (N_7911,N_6155,N_6032);
and U7912 (N_7912,N_6736,N_6237);
or U7913 (N_7913,N_6361,N_6449);
and U7914 (N_7914,N_6360,N_6443);
or U7915 (N_7915,N_6374,N_6996);
nor U7916 (N_7916,N_6387,N_6881);
nor U7917 (N_7917,N_6647,N_6397);
or U7918 (N_7918,N_6060,N_6009);
and U7919 (N_7919,N_6145,N_6820);
and U7920 (N_7920,N_6431,N_6541);
nand U7921 (N_7921,N_6205,N_6395);
nor U7922 (N_7922,N_6330,N_6102);
and U7923 (N_7923,N_6523,N_6829);
or U7924 (N_7924,N_6654,N_6553);
xnor U7925 (N_7925,N_6907,N_6492);
and U7926 (N_7926,N_6405,N_6330);
nor U7927 (N_7927,N_6953,N_6287);
xor U7928 (N_7928,N_6334,N_6515);
or U7929 (N_7929,N_6112,N_6888);
and U7930 (N_7930,N_6292,N_6890);
and U7931 (N_7931,N_6276,N_6642);
nor U7932 (N_7932,N_6590,N_6863);
nand U7933 (N_7933,N_6304,N_6565);
xnor U7934 (N_7934,N_6896,N_6337);
nand U7935 (N_7935,N_6027,N_6639);
or U7936 (N_7936,N_6174,N_6481);
and U7937 (N_7937,N_6206,N_6558);
xor U7938 (N_7938,N_6688,N_6200);
nand U7939 (N_7939,N_6707,N_6071);
nor U7940 (N_7940,N_6730,N_6775);
xnor U7941 (N_7941,N_6499,N_6705);
and U7942 (N_7942,N_6750,N_6806);
nor U7943 (N_7943,N_6789,N_6032);
nand U7944 (N_7944,N_6507,N_6119);
nor U7945 (N_7945,N_6325,N_6931);
or U7946 (N_7946,N_6910,N_6790);
and U7947 (N_7947,N_6774,N_6368);
nand U7948 (N_7948,N_6111,N_6206);
nor U7949 (N_7949,N_6820,N_6289);
or U7950 (N_7950,N_6926,N_6044);
and U7951 (N_7951,N_6619,N_6596);
xor U7952 (N_7952,N_6073,N_6233);
and U7953 (N_7953,N_6978,N_6376);
or U7954 (N_7954,N_6555,N_6489);
xor U7955 (N_7955,N_6061,N_6856);
and U7956 (N_7956,N_6697,N_6116);
or U7957 (N_7957,N_6654,N_6745);
nand U7958 (N_7958,N_6876,N_6147);
or U7959 (N_7959,N_6289,N_6612);
nand U7960 (N_7960,N_6565,N_6838);
xor U7961 (N_7961,N_6013,N_6696);
nand U7962 (N_7962,N_6282,N_6440);
nand U7963 (N_7963,N_6146,N_6545);
nor U7964 (N_7964,N_6507,N_6976);
xnor U7965 (N_7965,N_6411,N_6548);
or U7966 (N_7966,N_6822,N_6914);
xnor U7967 (N_7967,N_6772,N_6085);
nor U7968 (N_7968,N_6520,N_6111);
nor U7969 (N_7969,N_6470,N_6799);
nor U7970 (N_7970,N_6318,N_6949);
nor U7971 (N_7971,N_6215,N_6143);
and U7972 (N_7972,N_6899,N_6431);
nor U7973 (N_7973,N_6977,N_6288);
and U7974 (N_7974,N_6446,N_6303);
xnor U7975 (N_7975,N_6601,N_6349);
nor U7976 (N_7976,N_6374,N_6289);
xnor U7977 (N_7977,N_6433,N_6089);
nor U7978 (N_7978,N_6857,N_6705);
and U7979 (N_7979,N_6819,N_6117);
xor U7980 (N_7980,N_6956,N_6502);
nor U7981 (N_7981,N_6104,N_6038);
and U7982 (N_7982,N_6577,N_6057);
nor U7983 (N_7983,N_6830,N_6213);
xor U7984 (N_7984,N_6215,N_6048);
xnor U7985 (N_7985,N_6247,N_6696);
nand U7986 (N_7986,N_6621,N_6271);
nor U7987 (N_7987,N_6397,N_6857);
xnor U7988 (N_7988,N_6626,N_6147);
nor U7989 (N_7989,N_6502,N_6148);
nor U7990 (N_7990,N_6022,N_6129);
or U7991 (N_7991,N_6707,N_6642);
or U7992 (N_7992,N_6782,N_6175);
nand U7993 (N_7993,N_6429,N_6718);
xor U7994 (N_7994,N_6255,N_6290);
xor U7995 (N_7995,N_6942,N_6057);
and U7996 (N_7996,N_6258,N_6026);
and U7997 (N_7997,N_6364,N_6413);
nand U7998 (N_7998,N_6045,N_6723);
and U7999 (N_7999,N_6501,N_6818);
nor U8000 (N_8000,N_7904,N_7782);
or U8001 (N_8001,N_7452,N_7602);
or U8002 (N_8002,N_7775,N_7046);
xor U8003 (N_8003,N_7160,N_7663);
or U8004 (N_8004,N_7079,N_7637);
nand U8005 (N_8005,N_7983,N_7342);
xnor U8006 (N_8006,N_7657,N_7170);
xor U8007 (N_8007,N_7708,N_7744);
nand U8008 (N_8008,N_7013,N_7878);
or U8009 (N_8009,N_7634,N_7505);
nand U8010 (N_8010,N_7721,N_7416);
xor U8011 (N_8011,N_7591,N_7597);
or U8012 (N_8012,N_7988,N_7815);
and U8013 (N_8013,N_7444,N_7454);
and U8014 (N_8014,N_7670,N_7778);
and U8015 (N_8015,N_7433,N_7705);
nor U8016 (N_8016,N_7536,N_7964);
and U8017 (N_8017,N_7542,N_7723);
and U8018 (N_8018,N_7600,N_7659);
or U8019 (N_8019,N_7066,N_7768);
or U8020 (N_8020,N_7306,N_7661);
xnor U8021 (N_8021,N_7167,N_7840);
and U8022 (N_8022,N_7906,N_7489);
nand U8023 (N_8023,N_7493,N_7128);
nand U8024 (N_8024,N_7217,N_7293);
or U8025 (N_8025,N_7315,N_7126);
nor U8026 (N_8026,N_7621,N_7432);
nand U8027 (N_8027,N_7430,N_7387);
xnor U8028 (N_8028,N_7797,N_7015);
or U8029 (N_8029,N_7758,N_7463);
xnor U8030 (N_8030,N_7875,N_7051);
or U8031 (N_8031,N_7014,N_7521);
nor U8032 (N_8032,N_7762,N_7985);
xnor U8033 (N_8033,N_7265,N_7370);
nor U8034 (N_8034,N_7070,N_7226);
xnor U8035 (N_8035,N_7673,N_7156);
or U8036 (N_8036,N_7465,N_7199);
nor U8037 (N_8037,N_7526,N_7140);
nor U8038 (N_8038,N_7638,N_7543);
nand U8039 (N_8039,N_7149,N_7898);
nand U8040 (N_8040,N_7257,N_7854);
nor U8041 (N_8041,N_7755,N_7063);
xor U8042 (N_8042,N_7012,N_7656);
and U8043 (N_8043,N_7154,N_7296);
nand U8044 (N_8044,N_7279,N_7553);
or U8045 (N_8045,N_7089,N_7077);
nand U8046 (N_8046,N_7350,N_7415);
nor U8047 (N_8047,N_7820,N_7180);
xor U8048 (N_8048,N_7053,N_7589);
xnor U8049 (N_8049,N_7400,N_7485);
nand U8050 (N_8050,N_7232,N_7980);
xnor U8051 (N_8051,N_7410,N_7780);
nand U8052 (N_8052,N_7940,N_7733);
or U8053 (N_8053,N_7291,N_7698);
nand U8054 (N_8054,N_7675,N_7848);
nand U8055 (N_8055,N_7380,N_7484);
nor U8056 (N_8056,N_7990,N_7501);
or U8057 (N_8057,N_7408,N_7067);
and U8058 (N_8058,N_7435,N_7347);
nand U8059 (N_8059,N_7955,N_7532);
and U8060 (N_8060,N_7165,N_7795);
and U8061 (N_8061,N_7443,N_7606);
nor U8062 (N_8062,N_7006,N_7910);
xnor U8063 (N_8063,N_7935,N_7789);
nor U8064 (N_8064,N_7281,N_7139);
xor U8065 (N_8065,N_7561,N_7938);
or U8066 (N_8066,N_7831,N_7740);
nand U8067 (N_8067,N_7337,N_7665);
xnor U8068 (N_8068,N_7372,N_7141);
nor U8069 (N_8069,N_7897,N_7678);
or U8070 (N_8070,N_7256,N_7473);
xor U8071 (N_8071,N_7407,N_7556);
or U8072 (N_8072,N_7330,N_7274);
nand U8073 (N_8073,N_7168,N_7530);
and U8074 (N_8074,N_7539,N_7952);
and U8075 (N_8075,N_7286,N_7642);
xor U8076 (N_8076,N_7653,N_7502);
xor U8077 (N_8077,N_7321,N_7449);
and U8078 (N_8078,N_7022,N_7054);
nand U8079 (N_8079,N_7273,N_7162);
or U8080 (N_8080,N_7324,N_7929);
and U8081 (N_8081,N_7468,N_7576);
nand U8082 (N_8082,N_7475,N_7138);
nor U8083 (N_8083,N_7119,N_7424);
and U8084 (N_8084,N_7696,N_7428);
xor U8085 (N_8085,N_7945,N_7996);
nand U8086 (N_8086,N_7111,N_7537);
or U8087 (N_8087,N_7084,N_7693);
nor U8088 (N_8088,N_7800,N_7555);
xor U8089 (N_8089,N_7779,N_7335);
nor U8090 (N_8090,N_7214,N_7828);
and U8091 (N_8091,N_7161,N_7689);
nor U8092 (N_8092,N_7511,N_7982);
and U8093 (N_8093,N_7301,N_7426);
nor U8094 (N_8094,N_7813,N_7244);
or U8095 (N_8095,N_7453,N_7508);
nor U8096 (N_8096,N_7857,N_7056);
nor U8097 (N_8097,N_7130,N_7922);
nor U8098 (N_8098,N_7114,N_7303);
xor U8099 (N_8099,N_7242,N_7667);
or U8100 (N_8100,N_7967,N_7710);
xor U8101 (N_8101,N_7102,N_7345);
xor U8102 (N_8102,N_7429,N_7245);
or U8103 (N_8103,N_7065,N_7125);
xor U8104 (N_8104,N_7143,N_7490);
xor U8105 (N_8105,N_7000,N_7403);
nand U8106 (N_8106,N_7756,N_7282);
nand U8107 (N_8107,N_7839,N_7095);
and U8108 (N_8108,N_7654,N_7632);
and U8109 (N_8109,N_7367,N_7110);
nand U8110 (N_8110,N_7640,N_7185);
xor U8111 (N_8111,N_7129,N_7995);
xor U8112 (N_8112,N_7233,N_7725);
nand U8113 (N_8113,N_7458,N_7826);
xnor U8114 (N_8114,N_7099,N_7961);
nor U8115 (N_8115,N_7984,N_7237);
xor U8116 (N_8116,N_7767,N_7639);
xnor U8117 (N_8117,N_7451,N_7541);
xor U8118 (N_8118,N_7598,N_7506);
nand U8119 (N_8119,N_7374,N_7890);
or U8120 (N_8120,N_7920,N_7595);
nand U8121 (N_8121,N_7106,N_7219);
nand U8122 (N_8122,N_7847,N_7150);
nand U8123 (N_8123,N_7580,N_7072);
xor U8124 (N_8124,N_7781,N_7031);
nand U8125 (N_8125,N_7518,N_7575);
or U8126 (N_8126,N_7590,N_7799);
xor U8127 (N_8127,N_7169,N_7413);
nand U8128 (N_8128,N_7745,N_7849);
nand U8129 (N_8129,N_7047,N_7229);
nor U8130 (N_8130,N_7329,N_7866);
xnor U8131 (N_8131,N_7172,N_7123);
xor U8132 (N_8132,N_7001,N_7085);
or U8133 (N_8133,N_7810,N_7087);
nand U8134 (N_8134,N_7627,N_7397);
or U8135 (N_8135,N_7934,N_7236);
nand U8136 (N_8136,N_7535,N_7307);
or U8137 (N_8137,N_7609,N_7911);
nand U8138 (N_8138,N_7837,N_7592);
xor U8139 (N_8139,N_7208,N_7743);
xnor U8140 (N_8140,N_7914,N_7681);
or U8141 (N_8141,N_7533,N_7071);
nor U8142 (N_8142,N_7958,N_7183);
nand U8143 (N_8143,N_7297,N_7488);
nor U8144 (N_8144,N_7531,N_7896);
and U8145 (N_8145,N_7155,N_7951);
nor U8146 (N_8146,N_7855,N_7086);
or U8147 (N_8147,N_7747,N_7596);
nor U8148 (N_8148,N_7613,N_7157);
and U8149 (N_8149,N_7188,N_7997);
nor U8150 (N_8150,N_7300,N_7507);
and U8151 (N_8151,N_7749,N_7491);
xnor U8152 (N_8152,N_7908,N_7177);
or U8153 (N_8153,N_7729,N_7630);
or U8154 (N_8154,N_7970,N_7514);
nor U8155 (N_8155,N_7892,N_7614);
and U8156 (N_8156,N_7361,N_7028);
xnor U8157 (N_8157,N_7204,N_7651);
nand U8158 (N_8158,N_7247,N_7211);
xor U8159 (N_8159,N_7615,N_7624);
or U8160 (N_8160,N_7806,N_7702);
nand U8161 (N_8161,N_7176,N_7680);
nand U8162 (N_8162,N_7075,N_7009);
xnor U8163 (N_8163,N_7883,N_7133);
or U8164 (N_8164,N_7512,N_7704);
nor U8165 (N_8165,N_7016,N_7937);
xor U8166 (N_8166,N_7522,N_7406);
xor U8167 (N_8167,N_7579,N_7719);
xor U8168 (N_8168,N_7033,N_7690);
and U8169 (N_8169,N_7390,N_7159);
or U8170 (N_8170,N_7373,N_7998);
xnor U8171 (N_8171,N_7968,N_7442);
nor U8172 (N_8172,N_7635,N_7213);
xnor U8173 (N_8173,N_7646,N_7112);
xnor U8174 (N_8174,N_7860,N_7037);
nor U8175 (N_8175,N_7455,N_7326);
and U8176 (N_8176,N_7010,N_7986);
nor U8177 (N_8177,N_7474,N_7703);
and U8178 (N_8178,N_7513,N_7552);
xor U8179 (N_8179,N_7568,N_7164);
xnor U8180 (N_8180,N_7200,N_7540);
xnor U8181 (N_8181,N_7790,N_7885);
xor U8182 (N_8182,N_7915,N_7272);
or U8183 (N_8183,N_7956,N_7664);
xnor U8184 (N_8184,N_7499,N_7363);
or U8185 (N_8185,N_7946,N_7459);
and U8186 (N_8186,N_7832,N_7323);
and U8187 (N_8187,N_7973,N_7889);
xnor U8188 (N_8188,N_7369,N_7117);
xnor U8189 (N_8189,N_7251,N_7283);
or U8190 (N_8190,N_7030,N_7633);
xor U8191 (N_8191,N_7097,N_7305);
xnor U8192 (N_8192,N_7467,N_7868);
nand U8193 (N_8193,N_7757,N_7327);
xor U8194 (N_8194,N_7577,N_7405);
or U8195 (N_8195,N_7549,N_7909);
nor U8196 (N_8196,N_7829,N_7446);
or U8197 (N_8197,N_7817,N_7146);
xnor U8198 (N_8198,N_7811,N_7726);
nor U8199 (N_8199,N_7059,N_7179);
xor U8200 (N_8200,N_7375,N_7772);
nand U8201 (N_8201,N_7366,N_7730);
nor U8202 (N_8202,N_7560,N_7954);
nand U8203 (N_8203,N_7127,N_7944);
and U8204 (N_8204,N_7818,N_7497);
xor U8205 (N_8205,N_7346,N_7816);
nor U8206 (N_8206,N_7287,N_7103);
and U8207 (N_8207,N_7585,N_7975);
nor U8208 (N_8208,N_7671,N_7419);
nor U8209 (N_8209,N_7255,N_7234);
nand U8210 (N_8210,N_7333,N_7166);
nor U8211 (N_8211,N_7316,N_7082);
or U8212 (N_8212,N_7688,N_7069);
and U8213 (N_8213,N_7519,N_7581);
xnor U8214 (N_8214,N_7358,N_7094);
and U8215 (N_8215,N_7571,N_7684);
xnor U8216 (N_8216,N_7728,N_7224);
or U8217 (N_8217,N_7992,N_7202);
and U8218 (N_8218,N_7736,N_7605);
and U8219 (N_8219,N_7043,N_7073);
nor U8220 (N_8220,N_7100,N_7819);
and U8221 (N_8221,N_7979,N_7939);
and U8222 (N_8222,N_7331,N_7147);
or U8223 (N_8223,N_7978,N_7376);
xor U8224 (N_8224,N_7476,N_7221);
or U8225 (N_8225,N_7631,N_7360);
nor U8226 (N_8226,N_7804,N_7152);
or U8227 (N_8227,N_7520,N_7480);
or U8228 (N_8228,N_7824,N_7379);
xnor U8229 (N_8229,N_7076,N_7421);
nor U8230 (N_8230,N_7115,N_7777);
xor U8231 (N_8231,N_7096,N_7724);
and U8232 (N_8232,N_7737,N_7572);
or U8233 (N_8233,N_7351,N_7567);
nand U8234 (N_8234,N_7873,N_7439);
nand U8235 (N_8235,N_7108,N_7026);
nand U8236 (N_8236,N_7931,N_7151);
or U8237 (N_8237,N_7354,N_7864);
xor U8238 (N_8238,N_7548,N_7715);
and U8239 (N_8239,N_7275,N_7011);
nand U8240 (N_8240,N_7923,N_7083);
nor U8241 (N_8241,N_7999,N_7215);
and U8242 (N_8242,N_7713,N_7289);
nand U8243 (N_8243,N_7821,N_7398);
or U8244 (N_8244,N_7695,N_7960);
and U8245 (N_8245,N_7706,N_7765);
or U8246 (N_8246,N_7932,N_7271);
xor U8247 (N_8247,N_7278,N_7017);
nand U8248 (N_8248,N_7867,N_7963);
or U8249 (N_8249,N_7196,N_7791);
nor U8250 (N_8250,N_7163,N_7309);
xor U8251 (N_8251,N_7893,N_7976);
nor U8252 (N_8252,N_7807,N_7966);
nand U8253 (N_8253,N_7793,N_7220);
or U8254 (N_8254,N_7645,N_7238);
nor U8255 (N_8255,N_7647,N_7971);
and U8256 (N_8256,N_7525,N_7178);
xnor U8257 (N_8257,N_7641,N_7294);
and U8258 (N_8258,N_7034,N_7677);
xor U8259 (N_8259,N_7469,N_7871);
xnor U8260 (N_8260,N_7044,N_7668);
or U8261 (N_8261,N_7801,N_7352);
nand U8262 (N_8262,N_7392,N_7748);
and U8263 (N_8263,N_7718,N_7477);
nand U8264 (N_8264,N_7529,N_7322);
nand U8265 (N_8265,N_7662,N_7534);
xor U8266 (N_8266,N_7487,N_7672);
xnor U8267 (N_8267,N_7570,N_7741);
nand U8268 (N_8268,N_7882,N_7239);
nor U8269 (N_8269,N_7395,N_7830);
or U8270 (N_8270,N_7061,N_7792);
nand U8271 (N_8271,N_7833,N_7921);
xnor U8272 (N_8272,N_7563,N_7766);
or U8273 (N_8273,N_7040,N_7965);
or U8274 (N_8274,N_7422,N_7254);
nor U8275 (N_8275,N_7478,N_7803);
nor U8276 (N_8276,N_7863,N_7835);
nor U8277 (N_8277,N_7611,N_7423);
nor U8278 (N_8278,N_7240,N_7391);
and U8279 (N_8279,N_7124,N_7562);
or U8280 (N_8280,N_7717,N_7314);
nand U8281 (N_8281,N_7062,N_7158);
nand U8282 (N_8282,N_7699,N_7005);
xnor U8283 (N_8283,N_7144,N_7649);
or U8284 (N_8284,N_7586,N_7735);
xnor U8285 (N_8285,N_7685,N_7742);
nor U8286 (N_8286,N_7216,N_7796);
xor U8287 (N_8287,N_7994,N_7687);
or U8288 (N_8288,N_7510,N_7137);
nor U8289 (N_8289,N_7886,N_7905);
xor U8290 (N_8290,N_7859,N_7175);
nor U8291 (N_8291,N_7225,N_7784);
nand U8292 (N_8292,N_7470,N_7593);
nor U8293 (N_8293,N_7599,N_7738);
nand U8294 (N_8294,N_7991,N_7618);
or U8295 (N_8295,N_7527,N_7173);
and U8296 (N_8296,N_7045,N_7362);
xnor U8297 (N_8297,N_7720,N_7023);
or U8298 (N_8298,N_7104,N_7035);
xor U8299 (N_8299,N_7858,N_7107);
nor U8300 (N_8300,N_7620,N_7862);
nand U8301 (N_8301,N_7235,N_7381);
nor U8302 (N_8302,N_7121,N_7334);
nor U8303 (N_8303,N_7482,N_7223);
xnor U8304 (N_8304,N_7925,N_7136);
nor U8305 (N_8305,N_7093,N_7304);
xor U8306 (N_8306,N_7383,N_7365);
nand U8307 (N_8307,N_7834,N_7926);
nor U8308 (N_8308,N_7636,N_7650);
xor U8309 (N_8309,N_7288,N_7941);
xor U8310 (N_8310,N_7814,N_7626);
nor U8311 (N_8311,N_7879,N_7625);
nand U8312 (N_8312,N_7460,N_7686);
or U8313 (N_8313,N_7280,N_7264);
xor U8314 (N_8314,N_7852,N_7872);
nor U8315 (N_8315,N_7295,N_7588);
nand U8316 (N_8316,N_7524,N_7900);
xnor U8317 (N_8317,N_7569,N_7546);
xor U8318 (N_8318,N_7573,N_7957);
nand U8319 (N_8319,N_7888,N_7312);
or U8320 (N_8320,N_7697,N_7252);
xnor U8321 (N_8321,N_7655,N_7770);
nand U8322 (N_8322,N_7019,N_7064);
nor U8323 (N_8323,N_7574,N_7648);
or U8324 (N_8324,N_7763,N_7861);
nor U8325 (N_8325,N_7195,N_7565);
nor U8326 (N_8326,N_7382,N_7583);
xor U8327 (N_8327,N_7843,N_7148);
or U8328 (N_8328,N_7055,N_7846);
xnor U8329 (N_8329,N_7193,N_7068);
or U8330 (N_8330,N_7676,N_7943);
nand U8331 (N_8331,N_7538,N_7924);
xor U8332 (N_8332,N_7794,N_7558);
xor U8333 (N_8333,N_7285,N_7092);
and U8334 (N_8334,N_7771,N_7977);
xnor U8335 (N_8335,N_7427,N_7191);
nand U8336 (N_8336,N_7456,N_7187);
xnor U8337 (N_8337,N_7759,N_7388);
nand U8338 (N_8338,N_7825,N_7628);
and U8339 (N_8339,N_7972,N_7788);
xor U8340 (N_8340,N_7041,N_7623);
or U8341 (N_8341,N_7218,N_7343);
nor U8342 (N_8342,N_7750,N_7036);
xor U8343 (N_8343,N_7258,N_7503);
nor U8344 (N_8344,N_7716,N_7052);
xor U8345 (N_8345,N_7171,N_7617);
xnor U8346 (N_8346,N_7936,N_7584);
or U8347 (N_8347,N_7393,N_7032);
xnor U8348 (N_8348,N_7132,N_7042);
or U8349 (N_8349,N_7783,N_7808);
and U8350 (N_8350,N_7682,N_7269);
or U8351 (N_8351,N_7189,N_7604);
and U8352 (N_8352,N_7320,N_7660);
and U8353 (N_8353,N_7120,N_7057);
nor U8354 (N_8354,N_7739,N_7669);
nor U8355 (N_8355,N_7608,N_7544);
and U8356 (N_8356,N_7927,N_7643);
and U8357 (N_8357,N_7190,N_7754);
or U8358 (N_8358,N_7494,N_7338);
nor U8359 (N_8359,N_7298,N_7619);
and U8360 (N_8360,N_7845,N_7877);
xnor U8361 (N_8361,N_7098,N_7761);
or U8362 (N_8362,N_7805,N_7377);
or U8363 (N_8363,N_7116,N_7020);
xor U8364 (N_8364,N_7989,N_7891);
or U8365 (N_8365,N_7008,N_7776);
xnor U8366 (N_8366,N_7385,N_7746);
xor U8367 (N_8367,N_7384,N_7887);
nand U8368 (N_8368,N_7339,N_7142);
nand U8369 (N_8369,N_7587,N_7722);
xor U8370 (N_8370,N_7709,N_7050);
nand U8371 (N_8371,N_7090,N_7658);
and U8372 (N_8372,N_7049,N_7207);
nand U8373 (N_8373,N_7004,N_7901);
nand U8374 (N_8374,N_7263,N_7302);
xnor U8375 (N_8375,N_7058,N_7348);
or U8376 (N_8376,N_7311,N_7268);
or U8377 (N_8377,N_7876,N_7880);
xnor U8378 (N_8378,N_7394,N_7153);
xor U8379 (N_8379,N_7993,N_7332);
nand U8380 (N_8380,N_7024,N_7448);
or U8381 (N_8381,N_7974,N_7261);
xnor U8382 (N_8382,N_7039,N_7355);
xor U8383 (N_8383,N_7838,N_7959);
xnor U8384 (N_8384,N_7894,N_7317);
or U8385 (N_8385,N_7727,N_7319);
or U8386 (N_8386,N_7201,N_7559);
nand U8387 (N_8387,N_7438,N_7088);
or U8388 (N_8388,N_7582,N_7396);
nand U8389 (N_8389,N_7145,N_7248);
xor U8390 (N_8390,N_7437,N_7652);
xor U8391 (N_8391,N_7479,N_7205);
nor U8392 (N_8392,N_7349,N_7851);
xnor U8393 (N_8393,N_7341,N_7629);
or U8394 (N_8394,N_7025,N_7260);
nand U8395 (N_8395,N_7074,N_7773);
nand U8396 (N_8396,N_7947,N_7386);
xnor U8397 (N_8397,N_7492,N_7292);
and U8398 (N_8398,N_7197,N_7787);
or U8399 (N_8399,N_7812,N_7564);
xor U8400 (N_8400,N_7504,N_7495);
or U8401 (N_8401,N_7622,N_7753);
nand U8402 (N_8402,N_7987,N_7694);
xor U8403 (N_8403,N_7578,N_7371);
nor U8404 (N_8404,N_7357,N_7498);
and U8405 (N_8405,N_7554,N_7930);
xor U8406 (N_8406,N_7949,N_7368);
xnor U8407 (N_8407,N_7483,N_7404);
or U8408 (N_8408,N_7550,N_7230);
and U8409 (N_8409,N_7950,N_7557);
or U8410 (N_8410,N_7547,N_7203);
nor U8411 (N_8411,N_7184,N_7912);
nor U8412 (N_8412,N_7774,N_7091);
nand U8413 (N_8413,N_7299,N_7594);
xnor U8414 (N_8414,N_7222,N_7290);
and U8415 (N_8415,N_7276,N_7340);
xor U8416 (N_8416,N_7603,N_7711);
nor U8417 (N_8417,N_7842,N_7270);
or U8418 (N_8418,N_7029,N_7420);
xor U8419 (N_8419,N_7359,N_7691);
nand U8420 (N_8420,N_7122,N_7827);
xnor U8421 (N_8421,N_7409,N_7250);
nor U8422 (N_8422,N_7919,N_7021);
xor U8423 (N_8423,N_7003,N_7516);
nor U8424 (N_8424,N_7118,N_7325);
nand U8425 (N_8425,N_7198,N_7953);
nand U8426 (N_8426,N_7356,N_7701);
or U8427 (N_8427,N_7707,N_7809);
xnor U8428 (N_8428,N_7060,N_7402);
or U8429 (N_8429,N_7481,N_7227);
or U8430 (N_8430,N_7038,N_7607);
or U8431 (N_8431,N_7284,N_7486);
nand U8432 (N_8432,N_7318,N_7181);
nor U8433 (N_8433,N_7823,N_7109);
xor U8434 (N_8434,N_7007,N_7378);
nor U8435 (N_8435,N_7471,N_7853);
and U8436 (N_8436,N_7440,N_7445);
nor U8437 (N_8437,N_7266,N_7364);
and U8438 (N_8438,N_7277,N_7389);
nor U8439 (N_8439,N_7509,N_7464);
nor U8440 (N_8440,N_7884,N_7870);
xnor U8441 (N_8441,N_7948,N_7308);
and U8442 (N_8442,N_7844,N_7865);
nand U8443 (N_8443,N_7899,N_7895);
nand U8444 (N_8444,N_7210,N_7644);
and U8445 (N_8445,N_7785,N_7802);
nand U8446 (N_8446,N_7209,N_7135);
nand U8447 (N_8447,N_7523,N_7798);
or U8448 (N_8448,N_7353,N_7414);
nor U8449 (N_8449,N_7981,N_7683);
and U8450 (N_8450,N_7249,N_7466);
nor U8451 (N_8451,N_7856,N_7734);
or U8452 (N_8452,N_7764,N_7850);
and U8453 (N_8453,N_7447,N_7457);
and U8454 (N_8454,N_7048,N_7411);
nand U8455 (N_8455,N_7212,N_7874);
and U8456 (N_8456,N_7666,N_7336);
nor U8457 (N_8457,N_7610,N_7869);
xnor U8458 (N_8458,N_7328,N_7174);
nor U8459 (N_8459,N_7822,N_7918);
xnor U8460 (N_8460,N_7841,N_7472);
xor U8461 (N_8461,N_7902,N_7515);
xnor U8462 (N_8462,N_7916,N_7002);
and U8463 (N_8463,N_7425,N_7344);
nor U8464 (N_8464,N_7228,N_7679);
and U8465 (N_8465,N_7399,N_7969);
nand U8466 (N_8466,N_7246,N_7412);
and U8467 (N_8467,N_7241,N_7732);
or U8468 (N_8468,N_7113,N_7500);
or U8469 (N_8469,N_7461,N_7903);
xor U8470 (N_8470,N_7450,N_7313);
and U8471 (N_8471,N_7692,N_7192);
and U8472 (N_8472,N_7078,N_7913);
xor U8473 (N_8473,N_7101,N_7182);
nand U8474 (N_8474,N_7231,N_7712);
or U8475 (N_8475,N_7786,N_7517);
nor U8476 (N_8476,N_7496,N_7928);
and U8477 (N_8477,N_7417,N_7194);
nand U8478 (N_8478,N_7431,N_7080);
or U8479 (N_8479,N_7259,N_7206);
xor U8480 (N_8480,N_7836,N_7027);
and U8481 (N_8481,N_7434,N_7769);
nand U8482 (N_8482,N_7566,N_7545);
and U8483 (N_8483,N_7134,N_7714);
and U8484 (N_8484,N_7186,N_7942);
or U8485 (N_8485,N_7760,N_7700);
nand U8486 (N_8486,N_7441,N_7436);
xnor U8487 (N_8487,N_7243,N_7933);
or U8488 (N_8488,N_7616,N_7081);
xor U8489 (N_8489,N_7751,N_7131);
and U8490 (N_8490,N_7962,N_7907);
or U8491 (N_8491,N_7612,N_7267);
nand U8492 (N_8492,N_7674,N_7418);
and U8493 (N_8493,N_7105,N_7253);
or U8494 (N_8494,N_7528,N_7401);
or U8495 (N_8495,N_7881,N_7551);
nand U8496 (N_8496,N_7731,N_7752);
xnor U8497 (N_8497,N_7262,N_7601);
nand U8498 (N_8498,N_7462,N_7018);
and U8499 (N_8499,N_7310,N_7917);
and U8500 (N_8500,N_7177,N_7554);
or U8501 (N_8501,N_7323,N_7756);
and U8502 (N_8502,N_7650,N_7380);
xor U8503 (N_8503,N_7979,N_7978);
xnor U8504 (N_8504,N_7939,N_7829);
and U8505 (N_8505,N_7415,N_7904);
nor U8506 (N_8506,N_7297,N_7739);
xnor U8507 (N_8507,N_7831,N_7656);
xor U8508 (N_8508,N_7047,N_7409);
nand U8509 (N_8509,N_7902,N_7970);
xnor U8510 (N_8510,N_7389,N_7069);
or U8511 (N_8511,N_7172,N_7385);
nand U8512 (N_8512,N_7635,N_7827);
nor U8513 (N_8513,N_7133,N_7180);
and U8514 (N_8514,N_7513,N_7939);
nor U8515 (N_8515,N_7051,N_7686);
nor U8516 (N_8516,N_7452,N_7163);
or U8517 (N_8517,N_7611,N_7652);
nand U8518 (N_8518,N_7702,N_7644);
xor U8519 (N_8519,N_7893,N_7138);
xor U8520 (N_8520,N_7946,N_7108);
and U8521 (N_8521,N_7323,N_7672);
nor U8522 (N_8522,N_7428,N_7972);
or U8523 (N_8523,N_7244,N_7182);
and U8524 (N_8524,N_7335,N_7174);
nor U8525 (N_8525,N_7590,N_7812);
and U8526 (N_8526,N_7336,N_7748);
nand U8527 (N_8527,N_7614,N_7420);
and U8528 (N_8528,N_7565,N_7994);
xor U8529 (N_8529,N_7527,N_7299);
xor U8530 (N_8530,N_7338,N_7370);
and U8531 (N_8531,N_7850,N_7830);
nor U8532 (N_8532,N_7313,N_7360);
or U8533 (N_8533,N_7566,N_7524);
xnor U8534 (N_8534,N_7275,N_7133);
and U8535 (N_8535,N_7650,N_7935);
xor U8536 (N_8536,N_7345,N_7619);
nor U8537 (N_8537,N_7934,N_7227);
and U8538 (N_8538,N_7731,N_7200);
and U8539 (N_8539,N_7752,N_7944);
xnor U8540 (N_8540,N_7692,N_7200);
xor U8541 (N_8541,N_7235,N_7855);
nor U8542 (N_8542,N_7899,N_7469);
nand U8543 (N_8543,N_7876,N_7727);
xnor U8544 (N_8544,N_7559,N_7910);
nand U8545 (N_8545,N_7362,N_7264);
nand U8546 (N_8546,N_7057,N_7944);
nand U8547 (N_8547,N_7423,N_7266);
and U8548 (N_8548,N_7437,N_7610);
nor U8549 (N_8549,N_7137,N_7314);
or U8550 (N_8550,N_7028,N_7645);
and U8551 (N_8551,N_7331,N_7922);
nand U8552 (N_8552,N_7334,N_7194);
and U8553 (N_8553,N_7285,N_7181);
nand U8554 (N_8554,N_7054,N_7769);
and U8555 (N_8555,N_7794,N_7696);
xor U8556 (N_8556,N_7248,N_7328);
xnor U8557 (N_8557,N_7532,N_7541);
and U8558 (N_8558,N_7591,N_7078);
nor U8559 (N_8559,N_7509,N_7550);
nand U8560 (N_8560,N_7680,N_7840);
nand U8561 (N_8561,N_7231,N_7742);
xor U8562 (N_8562,N_7771,N_7437);
or U8563 (N_8563,N_7036,N_7501);
xnor U8564 (N_8564,N_7343,N_7146);
nand U8565 (N_8565,N_7841,N_7510);
nor U8566 (N_8566,N_7684,N_7059);
nand U8567 (N_8567,N_7607,N_7683);
xor U8568 (N_8568,N_7264,N_7177);
and U8569 (N_8569,N_7033,N_7982);
nand U8570 (N_8570,N_7246,N_7843);
xnor U8571 (N_8571,N_7673,N_7425);
or U8572 (N_8572,N_7885,N_7429);
xor U8573 (N_8573,N_7478,N_7980);
nand U8574 (N_8574,N_7012,N_7474);
or U8575 (N_8575,N_7598,N_7466);
nand U8576 (N_8576,N_7874,N_7272);
nor U8577 (N_8577,N_7265,N_7134);
or U8578 (N_8578,N_7637,N_7186);
or U8579 (N_8579,N_7491,N_7585);
nand U8580 (N_8580,N_7656,N_7607);
xnor U8581 (N_8581,N_7478,N_7971);
nand U8582 (N_8582,N_7654,N_7360);
or U8583 (N_8583,N_7401,N_7292);
xor U8584 (N_8584,N_7973,N_7500);
xor U8585 (N_8585,N_7726,N_7351);
and U8586 (N_8586,N_7674,N_7327);
xor U8587 (N_8587,N_7899,N_7945);
and U8588 (N_8588,N_7530,N_7251);
and U8589 (N_8589,N_7998,N_7297);
or U8590 (N_8590,N_7900,N_7746);
nand U8591 (N_8591,N_7992,N_7791);
and U8592 (N_8592,N_7949,N_7330);
nor U8593 (N_8593,N_7309,N_7951);
nor U8594 (N_8594,N_7024,N_7790);
nor U8595 (N_8595,N_7447,N_7188);
and U8596 (N_8596,N_7976,N_7104);
xor U8597 (N_8597,N_7012,N_7963);
nor U8598 (N_8598,N_7404,N_7615);
and U8599 (N_8599,N_7106,N_7099);
xor U8600 (N_8600,N_7476,N_7983);
nand U8601 (N_8601,N_7216,N_7810);
nand U8602 (N_8602,N_7993,N_7304);
nor U8603 (N_8603,N_7477,N_7390);
or U8604 (N_8604,N_7005,N_7332);
nand U8605 (N_8605,N_7694,N_7003);
nor U8606 (N_8606,N_7985,N_7458);
or U8607 (N_8607,N_7031,N_7628);
or U8608 (N_8608,N_7963,N_7457);
nand U8609 (N_8609,N_7738,N_7223);
and U8610 (N_8610,N_7757,N_7905);
nor U8611 (N_8611,N_7526,N_7549);
xnor U8612 (N_8612,N_7748,N_7333);
or U8613 (N_8613,N_7384,N_7368);
and U8614 (N_8614,N_7242,N_7137);
and U8615 (N_8615,N_7820,N_7325);
xnor U8616 (N_8616,N_7080,N_7945);
xnor U8617 (N_8617,N_7607,N_7994);
xnor U8618 (N_8618,N_7577,N_7784);
and U8619 (N_8619,N_7015,N_7055);
and U8620 (N_8620,N_7824,N_7893);
xor U8621 (N_8621,N_7014,N_7864);
nor U8622 (N_8622,N_7489,N_7305);
xor U8623 (N_8623,N_7205,N_7534);
xor U8624 (N_8624,N_7215,N_7079);
nor U8625 (N_8625,N_7379,N_7318);
nor U8626 (N_8626,N_7336,N_7156);
nand U8627 (N_8627,N_7605,N_7980);
and U8628 (N_8628,N_7332,N_7031);
nor U8629 (N_8629,N_7198,N_7712);
xnor U8630 (N_8630,N_7450,N_7691);
or U8631 (N_8631,N_7177,N_7304);
or U8632 (N_8632,N_7010,N_7418);
and U8633 (N_8633,N_7253,N_7334);
nand U8634 (N_8634,N_7219,N_7034);
xor U8635 (N_8635,N_7204,N_7590);
and U8636 (N_8636,N_7937,N_7780);
xor U8637 (N_8637,N_7439,N_7575);
xnor U8638 (N_8638,N_7294,N_7248);
xor U8639 (N_8639,N_7678,N_7853);
nor U8640 (N_8640,N_7016,N_7929);
nand U8641 (N_8641,N_7791,N_7443);
or U8642 (N_8642,N_7528,N_7052);
and U8643 (N_8643,N_7096,N_7381);
and U8644 (N_8644,N_7658,N_7765);
nor U8645 (N_8645,N_7417,N_7558);
nor U8646 (N_8646,N_7633,N_7561);
nand U8647 (N_8647,N_7858,N_7406);
or U8648 (N_8648,N_7033,N_7852);
nor U8649 (N_8649,N_7465,N_7285);
and U8650 (N_8650,N_7433,N_7871);
nand U8651 (N_8651,N_7402,N_7945);
xor U8652 (N_8652,N_7222,N_7322);
nand U8653 (N_8653,N_7413,N_7517);
nand U8654 (N_8654,N_7472,N_7421);
xor U8655 (N_8655,N_7597,N_7449);
xnor U8656 (N_8656,N_7865,N_7681);
nand U8657 (N_8657,N_7024,N_7854);
nand U8658 (N_8658,N_7917,N_7982);
nand U8659 (N_8659,N_7416,N_7543);
or U8660 (N_8660,N_7283,N_7239);
xnor U8661 (N_8661,N_7481,N_7029);
and U8662 (N_8662,N_7424,N_7836);
nand U8663 (N_8663,N_7770,N_7761);
or U8664 (N_8664,N_7306,N_7831);
nor U8665 (N_8665,N_7085,N_7098);
or U8666 (N_8666,N_7308,N_7359);
nand U8667 (N_8667,N_7602,N_7218);
and U8668 (N_8668,N_7077,N_7154);
nand U8669 (N_8669,N_7453,N_7126);
nand U8670 (N_8670,N_7126,N_7279);
nand U8671 (N_8671,N_7679,N_7717);
and U8672 (N_8672,N_7111,N_7381);
nand U8673 (N_8673,N_7385,N_7959);
or U8674 (N_8674,N_7195,N_7286);
nand U8675 (N_8675,N_7611,N_7563);
or U8676 (N_8676,N_7697,N_7442);
nand U8677 (N_8677,N_7957,N_7489);
or U8678 (N_8678,N_7144,N_7213);
and U8679 (N_8679,N_7085,N_7984);
nand U8680 (N_8680,N_7008,N_7001);
or U8681 (N_8681,N_7193,N_7835);
and U8682 (N_8682,N_7996,N_7345);
nor U8683 (N_8683,N_7733,N_7292);
and U8684 (N_8684,N_7659,N_7534);
or U8685 (N_8685,N_7617,N_7035);
and U8686 (N_8686,N_7794,N_7235);
or U8687 (N_8687,N_7658,N_7170);
nor U8688 (N_8688,N_7010,N_7851);
nand U8689 (N_8689,N_7795,N_7006);
or U8690 (N_8690,N_7040,N_7152);
nor U8691 (N_8691,N_7495,N_7997);
nand U8692 (N_8692,N_7850,N_7013);
or U8693 (N_8693,N_7049,N_7789);
nand U8694 (N_8694,N_7226,N_7507);
xnor U8695 (N_8695,N_7490,N_7252);
nor U8696 (N_8696,N_7808,N_7905);
xnor U8697 (N_8697,N_7471,N_7782);
or U8698 (N_8698,N_7023,N_7740);
xnor U8699 (N_8699,N_7357,N_7090);
nor U8700 (N_8700,N_7989,N_7631);
and U8701 (N_8701,N_7640,N_7472);
and U8702 (N_8702,N_7003,N_7904);
and U8703 (N_8703,N_7237,N_7404);
nand U8704 (N_8704,N_7881,N_7410);
or U8705 (N_8705,N_7601,N_7521);
and U8706 (N_8706,N_7296,N_7027);
nor U8707 (N_8707,N_7060,N_7536);
nor U8708 (N_8708,N_7264,N_7229);
or U8709 (N_8709,N_7332,N_7488);
and U8710 (N_8710,N_7260,N_7990);
or U8711 (N_8711,N_7235,N_7297);
or U8712 (N_8712,N_7120,N_7822);
and U8713 (N_8713,N_7547,N_7794);
xnor U8714 (N_8714,N_7019,N_7680);
xnor U8715 (N_8715,N_7537,N_7570);
xor U8716 (N_8716,N_7768,N_7296);
and U8717 (N_8717,N_7442,N_7517);
nand U8718 (N_8718,N_7081,N_7397);
nor U8719 (N_8719,N_7014,N_7659);
or U8720 (N_8720,N_7793,N_7646);
xnor U8721 (N_8721,N_7007,N_7300);
and U8722 (N_8722,N_7663,N_7569);
nor U8723 (N_8723,N_7078,N_7352);
nor U8724 (N_8724,N_7390,N_7196);
nand U8725 (N_8725,N_7718,N_7444);
or U8726 (N_8726,N_7574,N_7446);
or U8727 (N_8727,N_7576,N_7339);
nor U8728 (N_8728,N_7147,N_7765);
nand U8729 (N_8729,N_7302,N_7793);
and U8730 (N_8730,N_7187,N_7368);
nor U8731 (N_8731,N_7961,N_7169);
and U8732 (N_8732,N_7542,N_7861);
xor U8733 (N_8733,N_7371,N_7709);
nor U8734 (N_8734,N_7218,N_7295);
nor U8735 (N_8735,N_7545,N_7980);
and U8736 (N_8736,N_7186,N_7328);
nor U8737 (N_8737,N_7835,N_7768);
nor U8738 (N_8738,N_7510,N_7205);
or U8739 (N_8739,N_7312,N_7370);
or U8740 (N_8740,N_7646,N_7938);
or U8741 (N_8741,N_7483,N_7296);
nor U8742 (N_8742,N_7463,N_7309);
xor U8743 (N_8743,N_7531,N_7705);
xnor U8744 (N_8744,N_7418,N_7994);
xnor U8745 (N_8745,N_7380,N_7580);
xnor U8746 (N_8746,N_7397,N_7415);
xor U8747 (N_8747,N_7634,N_7029);
or U8748 (N_8748,N_7693,N_7879);
nand U8749 (N_8749,N_7942,N_7407);
and U8750 (N_8750,N_7880,N_7222);
xnor U8751 (N_8751,N_7328,N_7140);
or U8752 (N_8752,N_7164,N_7286);
and U8753 (N_8753,N_7100,N_7719);
nand U8754 (N_8754,N_7014,N_7556);
nor U8755 (N_8755,N_7200,N_7609);
xnor U8756 (N_8756,N_7061,N_7989);
or U8757 (N_8757,N_7474,N_7996);
xnor U8758 (N_8758,N_7060,N_7258);
nand U8759 (N_8759,N_7639,N_7880);
xnor U8760 (N_8760,N_7896,N_7161);
or U8761 (N_8761,N_7316,N_7249);
nand U8762 (N_8762,N_7906,N_7396);
and U8763 (N_8763,N_7119,N_7995);
nor U8764 (N_8764,N_7607,N_7110);
and U8765 (N_8765,N_7834,N_7554);
or U8766 (N_8766,N_7713,N_7595);
or U8767 (N_8767,N_7276,N_7115);
and U8768 (N_8768,N_7400,N_7668);
nor U8769 (N_8769,N_7347,N_7568);
or U8770 (N_8770,N_7218,N_7783);
and U8771 (N_8771,N_7985,N_7228);
or U8772 (N_8772,N_7495,N_7075);
nand U8773 (N_8773,N_7959,N_7639);
and U8774 (N_8774,N_7013,N_7106);
xor U8775 (N_8775,N_7286,N_7866);
xnor U8776 (N_8776,N_7182,N_7684);
xor U8777 (N_8777,N_7903,N_7637);
nor U8778 (N_8778,N_7160,N_7542);
xnor U8779 (N_8779,N_7426,N_7936);
nor U8780 (N_8780,N_7749,N_7310);
nand U8781 (N_8781,N_7898,N_7684);
nor U8782 (N_8782,N_7938,N_7011);
or U8783 (N_8783,N_7670,N_7135);
nor U8784 (N_8784,N_7193,N_7194);
xor U8785 (N_8785,N_7358,N_7834);
nand U8786 (N_8786,N_7085,N_7217);
nor U8787 (N_8787,N_7722,N_7376);
or U8788 (N_8788,N_7900,N_7564);
xor U8789 (N_8789,N_7479,N_7093);
nand U8790 (N_8790,N_7505,N_7638);
or U8791 (N_8791,N_7644,N_7663);
xor U8792 (N_8792,N_7246,N_7521);
nor U8793 (N_8793,N_7598,N_7451);
or U8794 (N_8794,N_7868,N_7230);
and U8795 (N_8795,N_7232,N_7659);
and U8796 (N_8796,N_7270,N_7347);
nand U8797 (N_8797,N_7591,N_7937);
and U8798 (N_8798,N_7091,N_7163);
nand U8799 (N_8799,N_7467,N_7582);
or U8800 (N_8800,N_7940,N_7100);
nor U8801 (N_8801,N_7465,N_7318);
or U8802 (N_8802,N_7971,N_7594);
or U8803 (N_8803,N_7455,N_7707);
and U8804 (N_8804,N_7602,N_7904);
nor U8805 (N_8805,N_7187,N_7601);
xnor U8806 (N_8806,N_7545,N_7409);
or U8807 (N_8807,N_7335,N_7371);
xor U8808 (N_8808,N_7629,N_7454);
and U8809 (N_8809,N_7579,N_7381);
xnor U8810 (N_8810,N_7788,N_7348);
or U8811 (N_8811,N_7348,N_7047);
nand U8812 (N_8812,N_7657,N_7599);
or U8813 (N_8813,N_7837,N_7218);
or U8814 (N_8814,N_7492,N_7055);
nand U8815 (N_8815,N_7059,N_7256);
or U8816 (N_8816,N_7927,N_7826);
and U8817 (N_8817,N_7567,N_7629);
or U8818 (N_8818,N_7341,N_7299);
and U8819 (N_8819,N_7684,N_7116);
xnor U8820 (N_8820,N_7425,N_7107);
xor U8821 (N_8821,N_7051,N_7345);
nand U8822 (N_8822,N_7901,N_7535);
xor U8823 (N_8823,N_7414,N_7123);
xnor U8824 (N_8824,N_7886,N_7373);
nor U8825 (N_8825,N_7100,N_7468);
and U8826 (N_8826,N_7742,N_7734);
nor U8827 (N_8827,N_7530,N_7173);
nor U8828 (N_8828,N_7956,N_7728);
and U8829 (N_8829,N_7922,N_7475);
nor U8830 (N_8830,N_7937,N_7296);
and U8831 (N_8831,N_7434,N_7721);
or U8832 (N_8832,N_7102,N_7256);
nand U8833 (N_8833,N_7268,N_7194);
or U8834 (N_8834,N_7755,N_7249);
or U8835 (N_8835,N_7819,N_7632);
nor U8836 (N_8836,N_7367,N_7629);
and U8837 (N_8837,N_7548,N_7337);
nor U8838 (N_8838,N_7074,N_7062);
nand U8839 (N_8839,N_7980,N_7786);
or U8840 (N_8840,N_7350,N_7738);
xor U8841 (N_8841,N_7527,N_7168);
nand U8842 (N_8842,N_7821,N_7474);
nor U8843 (N_8843,N_7365,N_7670);
and U8844 (N_8844,N_7892,N_7721);
nor U8845 (N_8845,N_7309,N_7593);
or U8846 (N_8846,N_7887,N_7444);
and U8847 (N_8847,N_7998,N_7008);
or U8848 (N_8848,N_7521,N_7668);
and U8849 (N_8849,N_7865,N_7626);
xor U8850 (N_8850,N_7159,N_7002);
nor U8851 (N_8851,N_7236,N_7392);
or U8852 (N_8852,N_7527,N_7829);
xnor U8853 (N_8853,N_7654,N_7775);
nor U8854 (N_8854,N_7428,N_7362);
or U8855 (N_8855,N_7355,N_7680);
xnor U8856 (N_8856,N_7969,N_7886);
or U8857 (N_8857,N_7167,N_7656);
and U8858 (N_8858,N_7378,N_7441);
nand U8859 (N_8859,N_7690,N_7389);
and U8860 (N_8860,N_7710,N_7392);
nor U8861 (N_8861,N_7113,N_7320);
and U8862 (N_8862,N_7246,N_7174);
xor U8863 (N_8863,N_7850,N_7224);
nand U8864 (N_8864,N_7996,N_7240);
or U8865 (N_8865,N_7528,N_7066);
nor U8866 (N_8866,N_7501,N_7055);
nand U8867 (N_8867,N_7031,N_7201);
or U8868 (N_8868,N_7956,N_7771);
nor U8869 (N_8869,N_7944,N_7082);
xnor U8870 (N_8870,N_7480,N_7238);
nand U8871 (N_8871,N_7664,N_7333);
xnor U8872 (N_8872,N_7858,N_7049);
nor U8873 (N_8873,N_7762,N_7019);
xor U8874 (N_8874,N_7614,N_7124);
nor U8875 (N_8875,N_7395,N_7178);
nand U8876 (N_8876,N_7730,N_7132);
and U8877 (N_8877,N_7250,N_7613);
and U8878 (N_8878,N_7046,N_7822);
and U8879 (N_8879,N_7861,N_7581);
xnor U8880 (N_8880,N_7593,N_7059);
and U8881 (N_8881,N_7376,N_7916);
or U8882 (N_8882,N_7519,N_7880);
xnor U8883 (N_8883,N_7029,N_7755);
and U8884 (N_8884,N_7466,N_7035);
or U8885 (N_8885,N_7241,N_7304);
or U8886 (N_8886,N_7505,N_7104);
and U8887 (N_8887,N_7548,N_7185);
nor U8888 (N_8888,N_7193,N_7926);
and U8889 (N_8889,N_7629,N_7472);
or U8890 (N_8890,N_7890,N_7818);
nand U8891 (N_8891,N_7572,N_7273);
nand U8892 (N_8892,N_7574,N_7357);
xor U8893 (N_8893,N_7291,N_7012);
nand U8894 (N_8894,N_7838,N_7260);
xnor U8895 (N_8895,N_7054,N_7923);
or U8896 (N_8896,N_7345,N_7071);
and U8897 (N_8897,N_7113,N_7971);
or U8898 (N_8898,N_7744,N_7838);
nor U8899 (N_8899,N_7636,N_7499);
nor U8900 (N_8900,N_7560,N_7359);
xnor U8901 (N_8901,N_7978,N_7136);
xnor U8902 (N_8902,N_7631,N_7107);
nor U8903 (N_8903,N_7353,N_7940);
nor U8904 (N_8904,N_7670,N_7817);
xor U8905 (N_8905,N_7760,N_7276);
or U8906 (N_8906,N_7286,N_7006);
nor U8907 (N_8907,N_7384,N_7208);
nor U8908 (N_8908,N_7532,N_7057);
xnor U8909 (N_8909,N_7144,N_7657);
nor U8910 (N_8910,N_7178,N_7500);
nor U8911 (N_8911,N_7480,N_7001);
nor U8912 (N_8912,N_7496,N_7165);
nor U8913 (N_8913,N_7413,N_7390);
nand U8914 (N_8914,N_7187,N_7864);
or U8915 (N_8915,N_7552,N_7784);
and U8916 (N_8916,N_7430,N_7786);
nand U8917 (N_8917,N_7630,N_7329);
nor U8918 (N_8918,N_7390,N_7068);
xnor U8919 (N_8919,N_7607,N_7945);
xnor U8920 (N_8920,N_7776,N_7344);
xnor U8921 (N_8921,N_7737,N_7722);
or U8922 (N_8922,N_7090,N_7363);
nand U8923 (N_8923,N_7455,N_7598);
nor U8924 (N_8924,N_7509,N_7243);
nor U8925 (N_8925,N_7976,N_7495);
and U8926 (N_8926,N_7028,N_7088);
and U8927 (N_8927,N_7828,N_7442);
nor U8928 (N_8928,N_7548,N_7215);
xor U8929 (N_8929,N_7799,N_7298);
and U8930 (N_8930,N_7595,N_7835);
and U8931 (N_8931,N_7031,N_7502);
nor U8932 (N_8932,N_7087,N_7992);
nor U8933 (N_8933,N_7225,N_7836);
or U8934 (N_8934,N_7994,N_7170);
and U8935 (N_8935,N_7328,N_7869);
xnor U8936 (N_8936,N_7418,N_7206);
or U8937 (N_8937,N_7961,N_7110);
nand U8938 (N_8938,N_7193,N_7315);
or U8939 (N_8939,N_7318,N_7614);
nor U8940 (N_8940,N_7375,N_7132);
or U8941 (N_8941,N_7655,N_7287);
and U8942 (N_8942,N_7173,N_7295);
nand U8943 (N_8943,N_7151,N_7328);
xnor U8944 (N_8944,N_7056,N_7515);
or U8945 (N_8945,N_7755,N_7506);
xor U8946 (N_8946,N_7887,N_7997);
or U8947 (N_8947,N_7783,N_7361);
and U8948 (N_8948,N_7971,N_7635);
and U8949 (N_8949,N_7964,N_7866);
nand U8950 (N_8950,N_7996,N_7833);
and U8951 (N_8951,N_7732,N_7090);
nand U8952 (N_8952,N_7537,N_7562);
or U8953 (N_8953,N_7152,N_7546);
nor U8954 (N_8954,N_7738,N_7250);
nand U8955 (N_8955,N_7168,N_7429);
xnor U8956 (N_8956,N_7596,N_7255);
nand U8957 (N_8957,N_7761,N_7586);
or U8958 (N_8958,N_7088,N_7842);
nand U8959 (N_8959,N_7887,N_7216);
or U8960 (N_8960,N_7034,N_7857);
and U8961 (N_8961,N_7780,N_7787);
and U8962 (N_8962,N_7593,N_7999);
nor U8963 (N_8963,N_7090,N_7281);
or U8964 (N_8964,N_7043,N_7455);
nor U8965 (N_8965,N_7492,N_7722);
xor U8966 (N_8966,N_7406,N_7603);
nor U8967 (N_8967,N_7780,N_7293);
or U8968 (N_8968,N_7380,N_7082);
nand U8969 (N_8969,N_7694,N_7307);
nor U8970 (N_8970,N_7811,N_7833);
nand U8971 (N_8971,N_7085,N_7306);
nand U8972 (N_8972,N_7418,N_7474);
nand U8973 (N_8973,N_7075,N_7062);
xor U8974 (N_8974,N_7659,N_7230);
and U8975 (N_8975,N_7702,N_7630);
xor U8976 (N_8976,N_7432,N_7473);
or U8977 (N_8977,N_7927,N_7120);
nand U8978 (N_8978,N_7258,N_7961);
or U8979 (N_8979,N_7022,N_7015);
and U8980 (N_8980,N_7506,N_7547);
and U8981 (N_8981,N_7955,N_7907);
xnor U8982 (N_8982,N_7197,N_7845);
and U8983 (N_8983,N_7375,N_7353);
xnor U8984 (N_8984,N_7289,N_7263);
nor U8985 (N_8985,N_7802,N_7560);
nor U8986 (N_8986,N_7078,N_7681);
or U8987 (N_8987,N_7686,N_7013);
nor U8988 (N_8988,N_7607,N_7713);
nor U8989 (N_8989,N_7085,N_7595);
nor U8990 (N_8990,N_7380,N_7184);
nor U8991 (N_8991,N_7418,N_7905);
xnor U8992 (N_8992,N_7902,N_7519);
xnor U8993 (N_8993,N_7759,N_7239);
or U8994 (N_8994,N_7180,N_7693);
and U8995 (N_8995,N_7331,N_7881);
or U8996 (N_8996,N_7764,N_7674);
and U8997 (N_8997,N_7395,N_7150);
nand U8998 (N_8998,N_7359,N_7088);
nor U8999 (N_8999,N_7030,N_7033);
and U9000 (N_9000,N_8839,N_8278);
nand U9001 (N_9001,N_8108,N_8378);
nand U9002 (N_9002,N_8700,N_8016);
and U9003 (N_9003,N_8810,N_8934);
nor U9004 (N_9004,N_8339,N_8431);
nand U9005 (N_9005,N_8753,N_8835);
nand U9006 (N_9006,N_8976,N_8920);
or U9007 (N_9007,N_8291,N_8873);
and U9008 (N_9008,N_8069,N_8484);
nand U9009 (N_9009,N_8355,N_8912);
or U9010 (N_9010,N_8034,N_8553);
and U9011 (N_9011,N_8226,N_8494);
nor U9012 (N_9012,N_8988,N_8817);
xnor U9013 (N_9013,N_8617,N_8423);
nand U9014 (N_9014,N_8891,N_8677);
or U9015 (N_9015,N_8369,N_8330);
and U9016 (N_9016,N_8635,N_8244);
nand U9017 (N_9017,N_8476,N_8075);
xnor U9018 (N_9018,N_8396,N_8883);
and U9019 (N_9019,N_8562,N_8032);
nand U9020 (N_9020,N_8812,N_8548);
or U9021 (N_9021,N_8798,N_8570);
nand U9022 (N_9022,N_8148,N_8914);
nor U9023 (N_9023,N_8434,N_8552);
and U9024 (N_9024,N_8213,N_8448);
nand U9025 (N_9025,N_8061,N_8158);
or U9026 (N_9026,N_8681,N_8357);
and U9027 (N_9027,N_8366,N_8654);
nor U9028 (N_9028,N_8403,N_8168);
xnor U9029 (N_9029,N_8749,N_8302);
and U9030 (N_9030,N_8325,N_8008);
xnor U9031 (N_9031,N_8203,N_8478);
and U9032 (N_9032,N_8876,N_8721);
or U9033 (N_9033,N_8050,N_8619);
nand U9034 (N_9034,N_8692,N_8204);
nand U9035 (N_9035,N_8684,N_8809);
nor U9036 (N_9036,N_8329,N_8400);
and U9037 (N_9037,N_8164,N_8121);
nor U9038 (N_9038,N_8287,N_8986);
or U9039 (N_9039,N_8348,N_8374);
xnor U9040 (N_9040,N_8547,N_8490);
xor U9041 (N_9041,N_8206,N_8615);
xnor U9042 (N_9042,N_8257,N_8272);
xnor U9043 (N_9043,N_8246,N_8450);
and U9044 (N_9044,N_8136,N_8077);
xnor U9045 (N_9045,N_8924,N_8189);
nor U9046 (N_9046,N_8200,N_8701);
nor U9047 (N_9047,N_8500,N_8998);
and U9048 (N_9048,N_8002,N_8483);
xnor U9049 (N_9049,N_8215,N_8183);
xnor U9050 (N_9050,N_8704,N_8543);
xor U9051 (N_9051,N_8087,N_8099);
and U9052 (N_9052,N_8740,N_8301);
nor U9053 (N_9053,N_8620,N_8387);
nand U9054 (N_9054,N_8937,N_8537);
nand U9055 (N_9055,N_8637,N_8385);
xor U9056 (N_9056,N_8129,N_8482);
xor U9057 (N_9057,N_8974,N_8877);
nand U9058 (N_9058,N_8182,N_8344);
nor U9059 (N_9059,N_8970,N_8541);
and U9060 (N_9060,N_8673,N_8456);
or U9061 (N_9061,N_8640,N_8699);
nand U9062 (N_9062,N_8493,N_8993);
and U9063 (N_9063,N_8091,N_8955);
nand U9064 (N_9064,N_8885,N_8795);
or U9065 (N_9065,N_8328,N_8017);
nand U9066 (N_9066,N_8720,N_8205);
nor U9067 (N_9067,N_8777,N_8459);
and U9068 (N_9068,N_8978,N_8686);
or U9069 (N_9069,N_8851,N_8815);
nor U9070 (N_9070,N_8828,N_8783);
or U9071 (N_9071,N_8001,N_8600);
nor U9072 (N_9072,N_8953,N_8659);
nor U9073 (N_9073,N_8706,N_8950);
nand U9074 (N_9074,N_8649,N_8167);
and U9075 (N_9075,N_8288,N_8729);
and U9076 (N_9076,N_8404,N_8438);
and U9077 (N_9077,N_8264,N_8405);
xnor U9078 (N_9078,N_8137,N_8664);
or U9079 (N_9079,N_8718,N_8286);
nand U9080 (N_9080,N_8020,N_8259);
or U9081 (N_9081,N_8837,N_8894);
nor U9082 (N_9082,N_8299,N_8643);
nor U9083 (N_9083,N_8453,N_8878);
xor U9084 (N_9084,N_8064,N_8967);
or U9085 (N_9085,N_8298,N_8157);
or U9086 (N_9086,N_8665,N_8505);
or U9087 (N_9087,N_8152,N_8680);
and U9088 (N_9088,N_8055,N_8309);
nand U9089 (N_9089,N_8965,N_8430);
nor U9090 (N_9090,N_8504,N_8793);
and U9091 (N_9091,N_8112,N_8223);
xor U9092 (N_9092,N_8388,N_8393);
or U9093 (N_9093,N_8280,N_8954);
nor U9094 (N_9094,N_8492,N_8766);
and U9095 (N_9095,N_8927,N_8778);
and U9096 (N_9096,N_8065,N_8319);
nand U9097 (N_9097,N_8524,N_8980);
or U9098 (N_9098,N_8243,N_8256);
xor U9099 (N_9099,N_8224,N_8119);
and U9100 (N_9100,N_8781,N_8907);
xnor U9101 (N_9101,N_8134,N_8426);
nor U9102 (N_9102,N_8195,N_8479);
nand U9103 (N_9103,N_8441,N_8916);
or U9104 (N_9104,N_8846,N_8807);
nand U9105 (N_9105,N_8058,N_8520);
or U9106 (N_9106,N_8031,N_8439);
nor U9107 (N_9107,N_8565,N_8586);
or U9108 (N_9108,N_8053,N_8521);
or U9109 (N_9109,N_8944,N_8481);
nor U9110 (N_9110,N_8592,N_8155);
nand U9111 (N_9111,N_8171,N_8669);
and U9112 (N_9112,N_8964,N_8271);
nor U9113 (N_9113,N_8282,N_8227);
or U9114 (N_9114,N_8502,N_8668);
or U9115 (N_9115,N_8116,N_8297);
xor U9116 (N_9116,N_8792,N_8544);
nand U9117 (N_9117,N_8130,N_8776);
nand U9118 (N_9118,N_8220,N_8103);
nor U9119 (N_9119,N_8047,N_8782);
xnor U9120 (N_9120,N_8219,N_8834);
and U9121 (N_9121,N_8917,N_8187);
or U9122 (N_9122,N_8341,N_8760);
xnor U9123 (N_9123,N_8429,N_8896);
or U9124 (N_9124,N_8336,N_8392);
and U9125 (N_9125,N_8176,N_8702);
nor U9126 (N_9126,N_8101,N_8254);
nor U9127 (N_9127,N_8790,N_8806);
or U9128 (N_9128,N_8146,N_8651);
nand U9129 (N_9129,N_8634,N_8987);
or U9130 (N_9130,N_8276,N_8554);
nand U9131 (N_9131,N_8049,N_8273);
or U9132 (N_9132,N_8144,N_8506);
and U9133 (N_9133,N_8150,N_8905);
nand U9134 (N_9134,N_8390,N_8169);
nand U9135 (N_9135,N_8024,N_8952);
or U9136 (N_9136,N_8908,N_8292);
nor U9137 (N_9137,N_8915,N_8051);
nor U9138 (N_9138,N_8451,N_8567);
nor U9139 (N_9139,N_8335,N_8501);
nand U9140 (N_9140,N_8229,N_8910);
xnor U9141 (N_9141,N_8421,N_8946);
nor U9142 (N_9142,N_8580,N_8962);
xnor U9143 (N_9143,N_8076,N_8402);
nand U9144 (N_9144,N_8349,N_8661);
nor U9145 (N_9145,N_8599,N_8646);
or U9146 (N_9146,N_8270,N_8004);
and U9147 (N_9147,N_8853,N_8179);
xor U9148 (N_9148,N_8687,N_8125);
or U9149 (N_9149,N_8576,N_8797);
and U9150 (N_9150,N_8117,N_8975);
or U9151 (N_9151,N_8671,N_8041);
nor U9152 (N_9152,N_8039,N_8327);
and U9153 (N_9153,N_8631,N_8585);
nor U9154 (N_9154,N_8695,N_8983);
or U9155 (N_9155,N_8762,N_8021);
or U9156 (N_9156,N_8942,N_8571);
xnor U9157 (N_9157,N_8512,N_8735);
xnor U9158 (N_9158,N_8488,N_8437);
nor U9159 (N_9159,N_8497,N_8086);
nor U9160 (N_9160,N_8089,N_8650);
nor U9161 (N_9161,N_8898,N_8399);
and U9162 (N_9162,N_8526,N_8078);
xor U9163 (N_9163,N_8621,N_8084);
or U9164 (N_9164,N_8030,N_8676);
or U9165 (N_9165,N_8864,N_8132);
and U9166 (N_9166,N_8638,N_8295);
nor U9167 (N_9167,N_8139,N_8574);
xnor U9168 (N_9168,N_8813,N_8048);
nor U9169 (N_9169,N_8845,N_8252);
and U9170 (N_9170,N_8192,N_8353);
xnor U9171 (N_9171,N_8727,N_8231);
or U9172 (N_9172,N_8308,N_8066);
or U9173 (N_9173,N_8623,N_8761);
or U9174 (N_9174,N_8391,N_8507);
nand U9175 (N_9175,N_8377,N_8029);
xor U9176 (N_9176,N_8829,N_8575);
nand U9177 (N_9177,N_8928,N_8546);
or U9178 (N_9178,N_8734,N_8703);
and U9179 (N_9179,N_8542,N_8859);
and U9180 (N_9180,N_8079,N_8123);
xnor U9181 (N_9181,N_8773,N_8332);
nor U9182 (N_9182,N_8359,N_8250);
and U9183 (N_9183,N_8268,N_8865);
and U9184 (N_9184,N_8923,N_8630);
nor U9185 (N_9185,N_8613,N_8995);
xnor U9186 (N_9186,N_8214,N_8682);
nor U9187 (N_9187,N_8265,N_8019);
xnor U9188 (N_9188,N_8808,N_8312);
and U9189 (N_9189,N_8406,N_8491);
xor U9190 (N_9190,N_8833,N_8610);
nand U9191 (N_9191,N_8140,N_8445);
and U9192 (N_9192,N_8342,N_8315);
nand U9193 (N_9193,N_8305,N_8105);
nand U9194 (N_9194,N_8338,N_8283);
or U9195 (N_9195,N_8296,N_8948);
or U9196 (N_9196,N_8056,N_8147);
and U9197 (N_9197,N_8424,N_8841);
and U9198 (N_9198,N_8323,N_8408);
and U9199 (N_9199,N_8872,N_8667);
nor U9200 (N_9200,N_8550,N_8011);
xnor U9201 (N_9201,N_8616,N_8557);
nor U9202 (N_9202,N_8417,N_8759);
xor U9203 (N_9203,N_8080,N_8895);
and U9204 (N_9204,N_8464,N_8867);
or U9205 (N_9205,N_8940,N_8629);
or U9206 (N_9206,N_8201,N_8584);
xnor U9207 (N_9207,N_8444,N_8248);
and U9208 (N_9208,N_8870,N_8320);
or U9209 (N_9209,N_8156,N_8627);
nand U9210 (N_9210,N_8715,N_8579);
nor U9211 (N_9211,N_8925,N_8757);
and U9212 (N_9212,N_8842,N_8868);
and U9213 (N_9213,N_8655,N_8674);
and U9214 (N_9214,N_8966,N_8693);
and U9215 (N_9215,N_8522,N_8281);
nor U9216 (N_9216,N_8538,N_8689);
or U9217 (N_9217,N_8931,N_8433);
or U9218 (N_9218,N_8819,N_8143);
nand U9219 (N_9219,N_8455,N_8710);
nand U9220 (N_9220,N_8595,N_8858);
nor U9221 (N_9221,N_8606,N_8266);
nor U9222 (N_9222,N_8892,N_8487);
and U9223 (N_9223,N_8515,N_8277);
xor U9224 (N_9224,N_8862,N_8785);
or U9225 (N_9225,N_8059,N_8111);
and U9226 (N_9226,N_8025,N_8672);
xor U9227 (N_9227,N_8717,N_8383);
or U9228 (N_9228,N_8696,N_8409);
nand U9229 (N_9229,N_8151,N_8899);
nand U9230 (N_9230,N_8871,N_8678);
and U9231 (N_9231,N_8849,N_8318);
nand U9232 (N_9232,N_8745,N_8234);
and U9233 (N_9233,N_8770,N_8193);
and U9234 (N_9234,N_8255,N_8648);
nor U9235 (N_9235,N_8074,N_8470);
xor U9236 (N_9236,N_8207,N_8890);
nor U9237 (N_9237,N_8474,N_8794);
and U9238 (N_9238,N_8957,N_8831);
nand U9239 (N_9239,N_8596,N_8855);
xor U9240 (N_9240,N_8211,N_8949);
or U9241 (N_9241,N_8670,N_8549);
nor U9242 (N_9242,N_8560,N_8352);
or U9243 (N_9243,N_8713,N_8376);
and U9244 (N_9244,N_8977,N_8569);
nand U9245 (N_9245,N_8178,N_8698);
xnor U9246 (N_9246,N_8919,N_8442);
nand U9247 (N_9247,N_8251,N_8503);
nor U9248 (N_9248,N_8893,N_8612);
nand U9249 (N_9249,N_8748,N_8690);
and U9250 (N_9250,N_8465,N_8856);
nor U9251 (N_9251,N_8943,N_8093);
and U9252 (N_9252,N_8758,N_8714);
nor U9253 (N_9253,N_8558,N_8389);
xnor U9254 (N_9254,N_8816,N_8477);
xor U9255 (N_9255,N_8365,N_8906);
or U9256 (N_9256,N_8197,N_8420);
or U9257 (N_9257,N_8581,N_8126);
nor U9258 (N_9258,N_8607,N_8113);
nand U9259 (N_9259,N_8992,N_8485);
or U9260 (N_9260,N_8830,N_8994);
nand U9261 (N_9261,N_8947,N_8982);
nor U9262 (N_9262,N_8469,N_8343);
and U9263 (N_9263,N_8901,N_8052);
nor U9264 (N_9264,N_8471,N_8632);
nand U9265 (N_9265,N_8744,N_8658);
nand U9266 (N_9266,N_8368,N_8751);
nor U9267 (N_9267,N_8708,N_8881);
nor U9268 (N_9268,N_8609,N_8060);
and U9269 (N_9269,N_8131,N_8394);
and U9270 (N_9270,N_8645,N_8597);
or U9271 (N_9271,N_8561,N_8054);
nor U9272 (N_9272,N_8922,N_8889);
or U9273 (N_9273,N_8539,N_8691);
nand U9274 (N_9274,N_8840,N_8913);
xnor U9275 (N_9275,N_8027,N_8769);
nand U9276 (N_9276,N_8968,N_8209);
and U9277 (N_9277,N_8733,N_8354);
or U9278 (N_9278,N_8598,N_8294);
xor U9279 (N_9279,N_8334,N_8918);
or U9280 (N_9280,N_8989,N_8238);
or U9281 (N_9281,N_8044,N_8832);
nor U9282 (N_9282,N_8743,N_8114);
xnor U9283 (N_9283,N_8719,N_8236);
or U9284 (N_9284,N_8162,N_8884);
and U9285 (N_9285,N_8432,N_8072);
nor U9286 (N_9286,N_8083,N_8014);
and U9287 (N_9287,N_8173,N_8124);
xnor U9288 (N_9288,N_8346,N_8530);
and U9289 (N_9289,N_8331,N_8958);
and U9290 (N_9290,N_8764,N_8533);
or U9291 (N_9291,N_8921,N_8767);
and U9292 (N_9292,N_8232,N_8133);
xor U9293 (N_9293,N_8208,N_8363);
xor U9294 (N_9294,N_8003,N_8730);
or U9295 (N_9295,N_8191,N_8628);
nor U9296 (N_9296,N_8563,N_8780);
nor U9297 (N_9297,N_8517,N_8033);
xnor U9298 (N_9298,N_8886,N_8768);
nor U9299 (N_9299,N_8181,N_8447);
and U9300 (N_9300,N_8847,N_8367);
nor U9301 (N_9301,N_8882,N_8073);
nor U9302 (N_9302,N_8971,N_8731);
or U9303 (N_9303,N_8887,N_8275);
xor U9304 (N_9304,N_8245,N_8801);
or U9305 (N_9305,N_8358,N_8775);
and U9306 (N_9306,N_8472,N_8235);
nor U9307 (N_9307,N_8258,N_8351);
xor U9308 (N_9308,N_8446,N_8568);
or U9309 (N_9309,N_8460,N_8821);
nand U9310 (N_9310,N_8666,N_8216);
nand U9311 (N_9311,N_8196,N_8737);
nor U9312 (N_9312,N_8165,N_8185);
and U9313 (N_9313,N_8804,N_8362);
nor U9314 (N_9314,N_8006,N_8023);
or U9315 (N_9315,N_8642,N_8791);
or U9316 (N_9316,N_8239,N_8267);
and U9317 (N_9317,N_8888,N_8373);
nor U9318 (N_9318,N_8796,N_8375);
xor U9319 (N_9319,N_8822,N_8956);
and U9320 (N_9320,N_8153,N_8532);
and U9321 (N_9321,N_8866,N_8711);
nor U9322 (N_9322,N_8127,N_8653);
and U9323 (N_9323,N_8799,N_8556);
or U9324 (N_9324,N_8736,N_8848);
and U9325 (N_9325,N_8138,N_8763);
nand U9326 (N_9326,N_8037,N_8863);
or U9327 (N_9327,N_8395,N_8588);
nor U9328 (N_9328,N_8860,N_8589);
or U9329 (N_9329,N_8109,N_8462);
xnor U9330 (N_9330,N_8739,N_8260);
xor U9331 (N_9331,N_8973,N_8159);
or U9332 (N_9332,N_8959,N_8716);
nor U9333 (N_9333,N_8062,N_8725);
and U9334 (N_9334,N_8009,N_8564);
nand U9335 (N_9335,N_8529,N_8466);
and U9336 (N_9336,N_8741,N_8583);
and U9337 (N_9337,N_8118,N_8765);
nor U9338 (N_9338,N_8262,N_8379);
or U9339 (N_9339,N_8941,N_8573);
nor U9340 (N_9340,N_8679,N_8932);
xnor U9341 (N_9341,N_8662,N_8401);
and U9342 (N_9342,N_8422,N_8135);
nor U9343 (N_9343,N_8082,N_8000);
xor U9344 (N_9344,N_8608,N_8427);
nor U9345 (N_9345,N_8461,N_8779);
and U9346 (N_9346,N_8789,N_8416);
nor U9347 (N_9347,N_8322,N_8188);
nand U9348 (N_9348,N_8516,N_8418);
nor U9349 (N_9349,N_8480,N_8514);
nand U9350 (N_9350,N_8811,N_8685);
or U9351 (N_9351,N_8939,N_8688);
nand U9352 (N_9352,N_8326,N_8614);
nor U9353 (N_9353,N_8874,N_8705);
or U9354 (N_9354,N_8194,N_8467);
or U9355 (N_9355,N_8384,N_8045);
nand U9356 (N_9356,N_8038,N_8641);
nor U9357 (N_9357,N_8750,N_8593);
and U9358 (N_9358,N_8802,N_8128);
or U9359 (N_9359,N_8694,N_8435);
or U9360 (N_9360,N_8857,N_8306);
xor U9361 (N_9361,N_8106,N_8774);
nor U9362 (N_9362,N_8601,N_8100);
nand U9363 (N_9363,N_8028,N_8879);
or U9364 (N_9364,N_8228,N_8827);
and U9365 (N_9365,N_8177,N_8566);
nand U9366 (N_9366,N_8425,N_8709);
nand U9367 (N_9367,N_8356,N_8578);
nor U9368 (N_9368,N_8436,N_8284);
nor U9369 (N_9369,N_8935,N_8249);
or U9370 (N_9370,N_8861,N_8602);
and U9371 (N_9371,N_8788,N_8911);
and U9372 (N_9372,N_8321,N_8198);
or U9373 (N_9373,N_8551,N_8996);
nand U9374 (N_9374,N_8412,N_8222);
and U9375 (N_9375,N_8904,N_8046);
and U9376 (N_9376,N_8337,N_8347);
xnor U9377 (N_9377,N_8285,N_8314);
nor U9378 (N_9378,N_8772,N_8969);
nand U9379 (N_9379,N_8818,N_8005);
and U9380 (N_9380,N_8850,N_8217);
nor U9381 (N_9381,N_8035,N_8724);
or U9382 (N_9382,N_8534,N_8929);
nand U9383 (N_9383,N_8622,N_8316);
or U9384 (N_9384,N_8202,N_8398);
nor U9385 (N_9385,N_8712,N_8022);
xor U9386 (N_9386,N_8519,N_8094);
nand U9387 (N_9387,N_8577,N_8869);
nor U9388 (N_9388,N_8897,N_8951);
nand U9389 (N_9389,N_8572,N_8333);
and U9390 (N_9390,N_8149,N_8122);
nand U9391 (N_9391,N_8241,N_8722);
xnor U9392 (N_9392,N_8990,N_8909);
or U9393 (N_9393,N_8513,N_8945);
or U9394 (N_9394,N_8210,N_8242);
or U9395 (N_9395,N_8902,N_8499);
nor U9396 (N_9396,N_8199,N_8269);
or U9397 (N_9397,N_8747,N_8936);
nand U9398 (N_9398,N_8440,N_8095);
or U9399 (N_9399,N_8836,N_8647);
and U9400 (N_9400,N_8605,N_8536);
nand U9401 (N_9401,N_8311,N_8361);
and U9402 (N_9402,N_8040,N_8457);
xnor U9403 (N_9403,N_8754,N_8324);
xnor U9404 (N_9404,N_8010,N_8085);
nor U9405 (N_9405,N_8397,N_8142);
nand U9406 (N_9406,N_8371,N_8372);
nand U9407 (N_9407,N_8510,N_8237);
and U9408 (N_9408,N_8824,N_8926);
nand U9409 (N_9409,N_8340,N_8261);
xor U9410 (N_9410,N_8820,N_8413);
and U9411 (N_9411,N_8317,N_8407);
and U9412 (N_9412,N_8525,N_8012);
or U9413 (N_9413,N_8068,N_8107);
and U9414 (N_9414,N_8495,N_8604);
nor U9415 (N_9415,N_8636,N_8771);
or U9416 (N_9416,N_8972,N_8212);
xnor U9417 (N_9417,N_8380,N_8611);
nor U9418 (N_9418,N_8752,N_8071);
xnor U9419 (N_9419,N_8307,N_8170);
or U9420 (N_9420,N_8723,N_8096);
xnor U9421 (N_9421,N_8999,N_8290);
nand U9422 (N_9422,N_8843,N_8279);
nand U9423 (N_9423,N_8555,N_8683);
xor U9424 (N_9424,N_8697,N_8088);
nand U9425 (N_9425,N_8304,N_8825);
and U9426 (N_9426,N_8414,N_8468);
and U9427 (N_9427,N_8300,N_8043);
xor U9428 (N_9428,N_8545,N_8496);
xnor U9429 (N_9429,N_8154,N_8590);
or U9430 (N_9430,N_8540,N_8742);
or U9431 (N_9431,N_8410,N_8900);
and U9432 (N_9432,N_8784,N_8063);
or U9433 (N_9433,N_8233,N_8067);
nor U9434 (N_9434,N_8018,N_8070);
xor U9435 (N_9435,N_8104,N_8523);
or U9436 (N_9436,N_8419,N_8186);
or U9437 (N_9437,N_8180,N_8814);
nor U9438 (N_9438,N_8528,N_8381);
nand U9439 (N_9439,N_8452,N_8527);
and U9440 (N_9440,N_8221,N_8428);
and U9441 (N_9441,N_8458,N_8175);
xnor U9442 (N_9442,N_8618,N_8145);
nor U9443 (N_9443,N_8633,N_8184);
nand U9444 (N_9444,N_8755,N_8225);
nand U9445 (N_9445,N_8559,N_8303);
xor U9446 (N_9446,N_8042,N_8036);
xor U9447 (N_9447,N_8026,N_8738);
nand U9448 (N_9448,N_8443,N_8930);
xor U9449 (N_9449,N_8786,N_8838);
nand U9450 (N_9450,N_8253,N_8880);
xnor U9451 (N_9451,N_8092,N_8531);
nor U9452 (N_9452,N_8293,N_8350);
xnor U9453 (N_9453,N_8963,N_8933);
nor U9454 (N_9454,N_8102,N_8449);
xor U9455 (N_9455,N_8263,N_8475);
nor U9456 (N_9456,N_8463,N_8746);
nand U9457 (N_9457,N_8370,N_8174);
or U9458 (N_9458,N_8938,N_8875);
nor U9459 (N_9459,N_8639,N_8160);
or U9460 (N_9460,N_8007,N_8508);
nor U9461 (N_9461,N_8756,N_8852);
nand U9462 (N_9462,N_8663,N_8726);
nor U9463 (N_9463,N_8509,N_8115);
and U9464 (N_9464,N_8675,N_8015);
or U9465 (N_9465,N_8518,N_8535);
or U9466 (N_9466,N_8454,N_8844);
and U9467 (N_9467,N_8090,N_8411);
nor U9468 (N_9468,N_8984,N_8486);
nor U9469 (N_9469,N_8057,N_8013);
or U9470 (N_9470,N_8240,N_8707);
nor U9471 (N_9471,N_8644,N_8854);
nor U9472 (N_9472,N_8289,N_8313);
and U9473 (N_9473,N_8603,N_8591);
nand U9474 (N_9474,N_8489,N_8805);
or U9475 (N_9475,N_8310,N_8511);
or U9476 (N_9476,N_8190,N_8415);
nand U9477 (N_9477,N_8382,N_8141);
and U9478 (N_9478,N_8803,N_8961);
and U9479 (N_9479,N_8652,N_8728);
nor U9480 (N_9480,N_8594,N_8360);
nand U9481 (N_9481,N_8991,N_8473);
nand U9482 (N_9482,N_8624,N_8979);
or U9483 (N_9483,N_8161,N_8985);
nor U9484 (N_9484,N_8787,N_8386);
or U9485 (N_9485,N_8120,N_8247);
and U9486 (N_9486,N_8997,N_8903);
or U9487 (N_9487,N_8587,N_8218);
xnor U9488 (N_9488,N_8626,N_8166);
xor U9489 (N_9489,N_8826,N_8660);
and U9490 (N_9490,N_8172,N_8656);
xnor U9491 (N_9491,N_8800,N_8498);
or U9492 (N_9492,N_8960,N_8823);
and U9493 (N_9493,N_8110,N_8163);
or U9494 (N_9494,N_8364,N_8098);
xor U9495 (N_9495,N_8981,N_8345);
nand U9496 (N_9496,N_8657,N_8582);
and U9497 (N_9497,N_8625,N_8274);
xnor U9498 (N_9498,N_8732,N_8230);
nand U9499 (N_9499,N_8097,N_8081);
nor U9500 (N_9500,N_8010,N_8562);
and U9501 (N_9501,N_8945,N_8178);
and U9502 (N_9502,N_8786,N_8636);
and U9503 (N_9503,N_8704,N_8203);
or U9504 (N_9504,N_8070,N_8051);
xor U9505 (N_9505,N_8365,N_8523);
or U9506 (N_9506,N_8529,N_8123);
and U9507 (N_9507,N_8360,N_8200);
and U9508 (N_9508,N_8946,N_8529);
or U9509 (N_9509,N_8202,N_8067);
nand U9510 (N_9510,N_8985,N_8129);
or U9511 (N_9511,N_8243,N_8673);
nand U9512 (N_9512,N_8260,N_8099);
xor U9513 (N_9513,N_8253,N_8151);
nor U9514 (N_9514,N_8239,N_8623);
xor U9515 (N_9515,N_8455,N_8243);
nand U9516 (N_9516,N_8978,N_8386);
or U9517 (N_9517,N_8736,N_8961);
or U9518 (N_9518,N_8519,N_8724);
xor U9519 (N_9519,N_8012,N_8885);
and U9520 (N_9520,N_8140,N_8340);
nand U9521 (N_9521,N_8368,N_8062);
or U9522 (N_9522,N_8488,N_8022);
and U9523 (N_9523,N_8279,N_8293);
nand U9524 (N_9524,N_8153,N_8418);
xnor U9525 (N_9525,N_8898,N_8645);
and U9526 (N_9526,N_8814,N_8156);
or U9527 (N_9527,N_8815,N_8086);
and U9528 (N_9528,N_8506,N_8744);
nor U9529 (N_9529,N_8486,N_8944);
nand U9530 (N_9530,N_8476,N_8156);
xor U9531 (N_9531,N_8097,N_8911);
xor U9532 (N_9532,N_8890,N_8994);
xnor U9533 (N_9533,N_8789,N_8162);
or U9534 (N_9534,N_8286,N_8843);
xnor U9535 (N_9535,N_8139,N_8150);
or U9536 (N_9536,N_8093,N_8226);
nor U9537 (N_9537,N_8057,N_8350);
nor U9538 (N_9538,N_8348,N_8804);
and U9539 (N_9539,N_8540,N_8026);
xor U9540 (N_9540,N_8263,N_8467);
and U9541 (N_9541,N_8581,N_8827);
nand U9542 (N_9542,N_8084,N_8775);
or U9543 (N_9543,N_8766,N_8840);
xnor U9544 (N_9544,N_8455,N_8245);
xnor U9545 (N_9545,N_8699,N_8060);
nor U9546 (N_9546,N_8232,N_8113);
and U9547 (N_9547,N_8302,N_8745);
nor U9548 (N_9548,N_8830,N_8767);
or U9549 (N_9549,N_8626,N_8627);
or U9550 (N_9550,N_8870,N_8433);
or U9551 (N_9551,N_8494,N_8146);
xor U9552 (N_9552,N_8394,N_8313);
or U9553 (N_9553,N_8056,N_8817);
nor U9554 (N_9554,N_8661,N_8740);
xnor U9555 (N_9555,N_8098,N_8055);
or U9556 (N_9556,N_8649,N_8130);
xnor U9557 (N_9557,N_8628,N_8433);
and U9558 (N_9558,N_8197,N_8317);
or U9559 (N_9559,N_8225,N_8702);
or U9560 (N_9560,N_8758,N_8009);
and U9561 (N_9561,N_8773,N_8798);
or U9562 (N_9562,N_8814,N_8705);
or U9563 (N_9563,N_8248,N_8068);
and U9564 (N_9564,N_8545,N_8572);
nand U9565 (N_9565,N_8092,N_8394);
nand U9566 (N_9566,N_8256,N_8876);
nand U9567 (N_9567,N_8872,N_8976);
and U9568 (N_9568,N_8916,N_8986);
and U9569 (N_9569,N_8832,N_8073);
nor U9570 (N_9570,N_8737,N_8608);
xor U9571 (N_9571,N_8525,N_8741);
or U9572 (N_9572,N_8628,N_8441);
xor U9573 (N_9573,N_8586,N_8754);
nor U9574 (N_9574,N_8532,N_8067);
and U9575 (N_9575,N_8856,N_8187);
and U9576 (N_9576,N_8213,N_8429);
nand U9577 (N_9577,N_8627,N_8630);
nor U9578 (N_9578,N_8061,N_8280);
nand U9579 (N_9579,N_8767,N_8095);
nor U9580 (N_9580,N_8862,N_8137);
nand U9581 (N_9581,N_8894,N_8542);
and U9582 (N_9582,N_8842,N_8543);
nand U9583 (N_9583,N_8775,N_8333);
xnor U9584 (N_9584,N_8064,N_8005);
xor U9585 (N_9585,N_8218,N_8075);
and U9586 (N_9586,N_8238,N_8097);
and U9587 (N_9587,N_8379,N_8877);
nand U9588 (N_9588,N_8084,N_8509);
xor U9589 (N_9589,N_8614,N_8152);
and U9590 (N_9590,N_8632,N_8622);
nand U9591 (N_9591,N_8914,N_8353);
nand U9592 (N_9592,N_8022,N_8930);
and U9593 (N_9593,N_8745,N_8458);
nor U9594 (N_9594,N_8418,N_8287);
or U9595 (N_9595,N_8296,N_8955);
nand U9596 (N_9596,N_8706,N_8433);
or U9597 (N_9597,N_8274,N_8263);
nand U9598 (N_9598,N_8264,N_8703);
and U9599 (N_9599,N_8338,N_8622);
nand U9600 (N_9600,N_8978,N_8085);
xor U9601 (N_9601,N_8398,N_8449);
and U9602 (N_9602,N_8224,N_8859);
or U9603 (N_9603,N_8288,N_8308);
and U9604 (N_9604,N_8524,N_8020);
nand U9605 (N_9605,N_8027,N_8508);
xor U9606 (N_9606,N_8214,N_8312);
or U9607 (N_9607,N_8201,N_8436);
or U9608 (N_9608,N_8008,N_8169);
nand U9609 (N_9609,N_8800,N_8450);
or U9610 (N_9610,N_8937,N_8568);
or U9611 (N_9611,N_8362,N_8825);
or U9612 (N_9612,N_8147,N_8625);
nand U9613 (N_9613,N_8964,N_8403);
nand U9614 (N_9614,N_8351,N_8003);
nand U9615 (N_9615,N_8051,N_8773);
or U9616 (N_9616,N_8489,N_8352);
nand U9617 (N_9617,N_8895,N_8327);
nor U9618 (N_9618,N_8938,N_8708);
xor U9619 (N_9619,N_8346,N_8069);
nand U9620 (N_9620,N_8724,N_8228);
and U9621 (N_9621,N_8016,N_8125);
and U9622 (N_9622,N_8909,N_8285);
nor U9623 (N_9623,N_8373,N_8609);
and U9624 (N_9624,N_8340,N_8002);
nand U9625 (N_9625,N_8515,N_8560);
nand U9626 (N_9626,N_8309,N_8831);
xnor U9627 (N_9627,N_8602,N_8679);
nand U9628 (N_9628,N_8387,N_8966);
nor U9629 (N_9629,N_8192,N_8693);
and U9630 (N_9630,N_8038,N_8893);
xor U9631 (N_9631,N_8293,N_8949);
nand U9632 (N_9632,N_8795,N_8856);
nand U9633 (N_9633,N_8105,N_8194);
or U9634 (N_9634,N_8152,N_8716);
nand U9635 (N_9635,N_8810,N_8023);
nand U9636 (N_9636,N_8894,N_8093);
xnor U9637 (N_9637,N_8762,N_8411);
nand U9638 (N_9638,N_8306,N_8492);
nor U9639 (N_9639,N_8385,N_8247);
and U9640 (N_9640,N_8771,N_8668);
or U9641 (N_9641,N_8926,N_8533);
nand U9642 (N_9642,N_8162,N_8853);
and U9643 (N_9643,N_8978,N_8602);
nor U9644 (N_9644,N_8962,N_8988);
nor U9645 (N_9645,N_8660,N_8988);
nand U9646 (N_9646,N_8360,N_8344);
and U9647 (N_9647,N_8027,N_8354);
nor U9648 (N_9648,N_8589,N_8873);
and U9649 (N_9649,N_8102,N_8584);
nand U9650 (N_9650,N_8192,N_8315);
and U9651 (N_9651,N_8867,N_8537);
nand U9652 (N_9652,N_8253,N_8369);
nand U9653 (N_9653,N_8427,N_8794);
nand U9654 (N_9654,N_8402,N_8380);
and U9655 (N_9655,N_8416,N_8446);
nor U9656 (N_9656,N_8971,N_8306);
nand U9657 (N_9657,N_8107,N_8461);
and U9658 (N_9658,N_8979,N_8193);
nor U9659 (N_9659,N_8300,N_8149);
and U9660 (N_9660,N_8754,N_8573);
nor U9661 (N_9661,N_8920,N_8108);
or U9662 (N_9662,N_8473,N_8387);
nand U9663 (N_9663,N_8845,N_8704);
and U9664 (N_9664,N_8100,N_8462);
or U9665 (N_9665,N_8825,N_8706);
and U9666 (N_9666,N_8981,N_8375);
nand U9667 (N_9667,N_8295,N_8956);
and U9668 (N_9668,N_8456,N_8547);
nand U9669 (N_9669,N_8563,N_8700);
nor U9670 (N_9670,N_8887,N_8077);
and U9671 (N_9671,N_8304,N_8007);
xor U9672 (N_9672,N_8172,N_8893);
or U9673 (N_9673,N_8664,N_8689);
xnor U9674 (N_9674,N_8217,N_8609);
and U9675 (N_9675,N_8854,N_8516);
or U9676 (N_9676,N_8877,N_8619);
nor U9677 (N_9677,N_8954,N_8225);
nor U9678 (N_9678,N_8821,N_8383);
nand U9679 (N_9679,N_8619,N_8696);
and U9680 (N_9680,N_8179,N_8451);
nand U9681 (N_9681,N_8675,N_8458);
or U9682 (N_9682,N_8243,N_8797);
nand U9683 (N_9683,N_8018,N_8617);
xor U9684 (N_9684,N_8791,N_8924);
nand U9685 (N_9685,N_8397,N_8027);
or U9686 (N_9686,N_8686,N_8238);
and U9687 (N_9687,N_8913,N_8545);
and U9688 (N_9688,N_8430,N_8397);
or U9689 (N_9689,N_8575,N_8526);
xor U9690 (N_9690,N_8211,N_8042);
or U9691 (N_9691,N_8805,N_8486);
or U9692 (N_9692,N_8424,N_8565);
nand U9693 (N_9693,N_8868,N_8711);
xnor U9694 (N_9694,N_8022,N_8315);
or U9695 (N_9695,N_8424,N_8908);
and U9696 (N_9696,N_8682,N_8867);
nand U9697 (N_9697,N_8005,N_8493);
nand U9698 (N_9698,N_8852,N_8277);
nand U9699 (N_9699,N_8958,N_8658);
and U9700 (N_9700,N_8352,N_8984);
or U9701 (N_9701,N_8129,N_8026);
or U9702 (N_9702,N_8537,N_8607);
and U9703 (N_9703,N_8178,N_8399);
nand U9704 (N_9704,N_8848,N_8950);
and U9705 (N_9705,N_8275,N_8560);
nand U9706 (N_9706,N_8569,N_8463);
or U9707 (N_9707,N_8288,N_8405);
or U9708 (N_9708,N_8367,N_8188);
nand U9709 (N_9709,N_8058,N_8268);
and U9710 (N_9710,N_8513,N_8392);
nor U9711 (N_9711,N_8924,N_8191);
or U9712 (N_9712,N_8861,N_8332);
xor U9713 (N_9713,N_8868,N_8624);
nand U9714 (N_9714,N_8320,N_8603);
nand U9715 (N_9715,N_8815,N_8482);
and U9716 (N_9716,N_8654,N_8286);
or U9717 (N_9717,N_8675,N_8797);
nand U9718 (N_9718,N_8959,N_8288);
nand U9719 (N_9719,N_8364,N_8958);
and U9720 (N_9720,N_8393,N_8426);
and U9721 (N_9721,N_8030,N_8940);
xor U9722 (N_9722,N_8093,N_8806);
or U9723 (N_9723,N_8337,N_8116);
nor U9724 (N_9724,N_8568,N_8914);
nor U9725 (N_9725,N_8530,N_8737);
and U9726 (N_9726,N_8709,N_8666);
nor U9727 (N_9727,N_8509,N_8812);
and U9728 (N_9728,N_8987,N_8843);
xor U9729 (N_9729,N_8718,N_8892);
nor U9730 (N_9730,N_8149,N_8677);
nand U9731 (N_9731,N_8090,N_8452);
nand U9732 (N_9732,N_8376,N_8022);
or U9733 (N_9733,N_8617,N_8439);
nor U9734 (N_9734,N_8173,N_8759);
or U9735 (N_9735,N_8064,N_8671);
xnor U9736 (N_9736,N_8128,N_8740);
nor U9737 (N_9737,N_8943,N_8170);
nand U9738 (N_9738,N_8791,N_8913);
nor U9739 (N_9739,N_8391,N_8488);
nor U9740 (N_9740,N_8108,N_8285);
or U9741 (N_9741,N_8132,N_8728);
and U9742 (N_9742,N_8009,N_8400);
nor U9743 (N_9743,N_8061,N_8261);
nand U9744 (N_9744,N_8276,N_8471);
nor U9745 (N_9745,N_8450,N_8468);
or U9746 (N_9746,N_8145,N_8831);
and U9747 (N_9747,N_8812,N_8852);
nand U9748 (N_9748,N_8645,N_8218);
or U9749 (N_9749,N_8129,N_8276);
or U9750 (N_9750,N_8769,N_8958);
and U9751 (N_9751,N_8647,N_8790);
nand U9752 (N_9752,N_8340,N_8252);
or U9753 (N_9753,N_8608,N_8061);
xor U9754 (N_9754,N_8144,N_8462);
nand U9755 (N_9755,N_8014,N_8611);
nand U9756 (N_9756,N_8199,N_8356);
nand U9757 (N_9757,N_8532,N_8483);
or U9758 (N_9758,N_8850,N_8509);
or U9759 (N_9759,N_8397,N_8133);
nand U9760 (N_9760,N_8161,N_8527);
nor U9761 (N_9761,N_8963,N_8681);
or U9762 (N_9762,N_8257,N_8735);
nor U9763 (N_9763,N_8207,N_8551);
nor U9764 (N_9764,N_8741,N_8265);
or U9765 (N_9765,N_8204,N_8982);
and U9766 (N_9766,N_8254,N_8804);
nand U9767 (N_9767,N_8062,N_8619);
xnor U9768 (N_9768,N_8222,N_8614);
and U9769 (N_9769,N_8364,N_8378);
nor U9770 (N_9770,N_8704,N_8607);
nand U9771 (N_9771,N_8405,N_8676);
nor U9772 (N_9772,N_8107,N_8444);
or U9773 (N_9773,N_8186,N_8437);
xor U9774 (N_9774,N_8475,N_8721);
nand U9775 (N_9775,N_8426,N_8852);
nor U9776 (N_9776,N_8394,N_8287);
and U9777 (N_9777,N_8649,N_8584);
and U9778 (N_9778,N_8378,N_8390);
nand U9779 (N_9779,N_8054,N_8344);
xnor U9780 (N_9780,N_8760,N_8653);
xor U9781 (N_9781,N_8716,N_8585);
nor U9782 (N_9782,N_8327,N_8907);
xor U9783 (N_9783,N_8034,N_8548);
nand U9784 (N_9784,N_8797,N_8558);
or U9785 (N_9785,N_8502,N_8410);
and U9786 (N_9786,N_8650,N_8945);
or U9787 (N_9787,N_8790,N_8234);
and U9788 (N_9788,N_8553,N_8446);
or U9789 (N_9789,N_8225,N_8864);
or U9790 (N_9790,N_8712,N_8986);
nor U9791 (N_9791,N_8056,N_8317);
nor U9792 (N_9792,N_8696,N_8971);
nand U9793 (N_9793,N_8840,N_8616);
and U9794 (N_9794,N_8731,N_8350);
or U9795 (N_9795,N_8160,N_8034);
nand U9796 (N_9796,N_8123,N_8823);
nor U9797 (N_9797,N_8714,N_8740);
nor U9798 (N_9798,N_8208,N_8711);
xnor U9799 (N_9799,N_8025,N_8093);
xnor U9800 (N_9800,N_8178,N_8507);
and U9801 (N_9801,N_8306,N_8933);
nand U9802 (N_9802,N_8210,N_8113);
and U9803 (N_9803,N_8959,N_8014);
xnor U9804 (N_9804,N_8929,N_8790);
or U9805 (N_9805,N_8951,N_8722);
and U9806 (N_9806,N_8731,N_8571);
nand U9807 (N_9807,N_8418,N_8564);
and U9808 (N_9808,N_8474,N_8037);
nor U9809 (N_9809,N_8819,N_8274);
nand U9810 (N_9810,N_8172,N_8951);
or U9811 (N_9811,N_8246,N_8949);
xor U9812 (N_9812,N_8310,N_8756);
and U9813 (N_9813,N_8255,N_8043);
nor U9814 (N_9814,N_8680,N_8846);
nor U9815 (N_9815,N_8405,N_8878);
nand U9816 (N_9816,N_8794,N_8320);
and U9817 (N_9817,N_8144,N_8577);
nand U9818 (N_9818,N_8615,N_8291);
xnor U9819 (N_9819,N_8412,N_8409);
xnor U9820 (N_9820,N_8105,N_8829);
or U9821 (N_9821,N_8314,N_8466);
and U9822 (N_9822,N_8013,N_8700);
xnor U9823 (N_9823,N_8265,N_8484);
and U9824 (N_9824,N_8077,N_8284);
and U9825 (N_9825,N_8864,N_8193);
nor U9826 (N_9826,N_8459,N_8039);
nand U9827 (N_9827,N_8727,N_8707);
nand U9828 (N_9828,N_8508,N_8398);
or U9829 (N_9829,N_8270,N_8477);
nand U9830 (N_9830,N_8091,N_8206);
nand U9831 (N_9831,N_8226,N_8658);
nor U9832 (N_9832,N_8465,N_8537);
or U9833 (N_9833,N_8411,N_8871);
nand U9834 (N_9834,N_8292,N_8632);
nor U9835 (N_9835,N_8143,N_8188);
and U9836 (N_9836,N_8736,N_8458);
or U9837 (N_9837,N_8199,N_8369);
nor U9838 (N_9838,N_8154,N_8355);
nor U9839 (N_9839,N_8184,N_8397);
nand U9840 (N_9840,N_8954,N_8601);
or U9841 (N_9841,N_8835,N_8728);
or U9842 (N_9842,N_8028,N_8691);
xnor U9843 (N_9843,N_8947,N_8907);
and U9844 (N_9844,N_8080,N_8584);
and U9845 (N_9845,N_8634,N_8035);
nor U9846 (N_9846,N_8705,N_8880);
nand U9847 (N_9847,N_8718,N_8130);
or U9848 (N_9848,N_8924,N_8628);
nand U9849 (N_9849,N_8645,N_8567);
and U9850 (N_9850,N_8313,N_8391);
nand U9851 (N_9851,N_8668,N_8293);
nand U9852 (N_9852,N_8205,N_8655);
or U9853 (N_9853,N_8307,N_8379);
and U9854 (N_9854,N_8758,N_8271);
xor U9855 (N_9855,N_8106,N_8054);
nand U9856 (N_9856,N_8036,N_8744);
xor U9857 (N_9857,N_8675,N_8308);
or U9858 (N_9858,N_8430,N_8536);
xor U9859 (N_9859,N_8880,N_8782);
xnor U9860 (N_9860,N_8400,N_8854);
and U9861 (N_9861,N_8595,N_8780);
nand U9862 (N_9862,N_8758,N_8625);
xor U9863 (N_9863,N_8786,N_8260);
nand U9864 (N_9864,N_8734,N_8896);
nor U9865 (N_9865,N_8597,N_8283);
xor U9866 (N_9866,N_8397,N_8749);
and U9867 (N_9867,N_8135,N_8278);
and U9868 (N_9868,N_8628,N_8634);
nand U9869 (N_9869,N_8161,N_8422);
nor U9870 (N_9870,N_8640,N_8396);
and U9871 (N_9871,N_8735,N_8824);
nand U9872 (N_9872,N_8689,N_8872);
or U9873 (N_9873,N_8773,N_8121);
and U9874 (N_9874,N_8115,N_8396);
and U9875 (N_9875,N_8319,N_8295);
or U9876 (N_9876,N_8032,N_8919);
nand U9877 (N_9877,N_8315,N_8840);
and U9878 (N_9878,N_8321,N_8579);
nor U9879 (N_9879,N_8708,N_8962);
and U9880 (N_9880,N_8851,N_8483);
xor U9881 (N_9881,N_8902,N_8971);
and U9882 (N_9882,N_8576,N_8046);
and U9883 (N_9883,N_8317,N_8241);
and U9884 (N_9884,N_8186,N_8027);
nor U9885 (N_9885,N_8227,N_8719);
or U9886 (N_9886,N_8876,N_8323);
xnor U9887 (N_9887,N_8174,N_8104);
and U9888 (N_9888,N_8846,N_8785);
and U9889 (N_9889,N_8037,N_8249);
xor U9890 (N_9890,N_8106,N_8919);
nor U9891 (N_9891,N_8309,N_8615);
xnor U9892 (N_9892,N_8057,N_8110);
nand U9893 (N_9893,N_8563,N_8653);
and U9894 (N_9894,N_8826,N_8638);
xnor U9895 (N_9895,N_8749,N_8210);
nor U9896 (N_9896,N_8500,N_8607);
xnor U9897 (N_9897,N_8751,N_8891);
xor U9898 (N_9898,N_8236,N_8974);
nand U9899 (N_9899,N_8288,N_8116);
or U9900 (N_9900,N_8918,N_8857);
or U9901 (N_9901,N_8791,N_8170);
xor U9902 (N_9902,N_8869,N_8003);
nor U9903 (N_9903,N_8316,N_8460);
nor U9904 (N_9904,N_8057,N_8816);
and U9905 (N_9905,N_8911,N_8044);
nand U9906 (N_9906,N_8519,N_8383);
xor U9907 (N_9907,N_8517,N_8760);
nor U9908 (N_9908,N_8658,N_8799);
nand U9909 (N_9909,N_8614,N_8726);
or U9910 (N_9910,N_8045,N_8164);
xor U9911 (N_9911,N_8127,N_8783);
and U9912 (N_9912,N_8646,N_8605);
xor U9913 (N_9913,N_8240,N_8346);
nor U9914 (N_9914,N_8578,N_8378);
or U9915 (N_9915,N_8613,N_8279);
or U9916 (N_9916,N_8310,N_8982);
xnor U9917 (N_9917,N_8193,N_8957);
or U9918 (N_9918,N_8919,N_8321);
nor U9919 (N_9919,N_8043,N_8247);
xor U9920 (N_9920,N_8539,N_8292);
nand U9921 (N_9921,N_8976,N_8074);
xor U9922 (N_9922,N_8286,N_8478);
and U9923 (N_9923,N_8389,N_8463);
xnor U9924 (N_9924,N_8033,N_8739);
nor U9925 (N_9925,N_8697,N_8083);
nor U9926 (N_9926,N_8489,N_8633);
or U9927 (N_9927,N_8629,N_8464);
or U9928 (N_9928,N_8391,N_8806);
or U9929 (N_9929,N_8952,N_8513);
xnor U9930 (N_9930,N_8129,N_8184);
and U9931 (N_9931,N_8638,N_8900);
nand U9932 (N_9932,N_8275,N_8265);
xor U9933 (N_9933,N_8391,N_8239);
xor U9934 (N_9934,N_8742,N_8296);
nand U9935 (N_9935,N_8188,N_8085);
nor U9936 (N_9936,N_8857,N_8597);
and U9937 (N_9937,N_8206,N_8763);
nand U9938 (N_9938,N_8281,N_8862);
xnor U9939 (N_9939,N_8989,N_8744);
xor U9940 (N_9940,N_8585,N_8581);
nand U9941 (N_9941,N_8028,N_8334);
or U9942 (N_9942,N_8921,N_8484);
or U9943 (N_9943,N_8009,N_8042);
xnor U9944 (N_9944,N_8875,N_8426);
nand U9945 (N_9945,N_8129,N_8530);
nor U9946 (N_9946,N_8989,N_8966);
nor U9947 (N_9947,N_8777,N_8394);
xor U9948 (N_9948,N_8480,N_8407);
nor U9949 (N_9949,N_8891,N_8270);
xor U9950 (N_9950,N_8569,N_8716);
nor U9951 (N_9951,N_8181,N_8467);
xor U9952 (N_9952,N_8684,N_8047);
nor U9953 (N_9953,N_8960,N_8984);
nor U9954 (N_9954,N_8699,N_8341);
and U9955 (N_9955,N_8312,N_8572);
xnor U9956 (N_9956,N_8646,N_8296);
nand U9957 (N_9957,N_8231,N_8272);
and U9958 (N_9958,N_8884,N_8307);
and U9959 (N_9959,N_8806,N_8282);
nor U9960 (N_9960,N_8138,N_8506);
and U9961 (N_9961,N_8591,N_8989);
and U9962 (N_9962,N_8282,N_8074);
and U9963 (N_9963,N_8727,N_8295);
and U9964 (N_9964,N_8657,N_8396);
nand U9965 (N_9965,N_8932,N_8962);
xor U9966 (N_9966,N_8780,N_8321);
and U9967 (N_9967,N_8682,N_8075);
xnor U9968 (N_9968,N_8926,N_8736);
nor U9969 (N_9969,N_8363,N_8169);
nand U9970 (N_9970,N_8612,N_8749);
nand U9971 (N_9971,N_8442,N_8780);
or U9972 (N_9972,N_8467,N_8611);
or U9973 (N_9973,N_8770,N_8329);
nand U9974 (N_9974,N_8619,N_8335);
nand U9975 (N_9975,N_8997,N_8614);
nor U9976 (N_9976,N_8000,N_8644);
or U9977 (N_9977,N_8930,N_8867);
and U9978 (N_9978,N_8306,N_8534);
or U9979 (N_9979,N_8680,N_8236);
xor U9980 (N_9980,N_8515,N_8202);
and U9981 (N_9981,N_8675,N_8755);
nand U9982 (N_9982,N_8410,N_8544);
xor U9983 (N_9983,N_8951,N_8335);
and U9984 (N_9984,N_8858,N_8472);
nor U9985 (N_9985,N_8307,N_8449);
nor U9986 (N_9986,N_8970,N_8458);
nor U9987 (N_9987,N_8050,N_8080);
nand U9988 (N_9988,N_8137,N_8200);
xnor U9989 (N_9989,N_8833,N_8810);
and U9990 (N_9990,N_8001,N_8910);
nor U9991 (N_9991,N_8576,N_8385);
nand U9992 (N_9992,N_8698,N_8994);
or U9993 (N_9993,N_8217,N_8245);
or U9994 (N_9994,N_8764,N_8899);
and U9995 (N_9995,N_8096,N_8646);
or U9996 (N_9996,N_8168,N_8404);
nand U9997 (N_9997,N_8518,N_8571);
nand U9998 (N_9998,N_8244,N_8463);
and U9999 (N_9999,N_8148,N_8502);
and U10000 (N_10000,N_9989,N_9720);
nor U10001 (N_10001,N_9201,N_9859);
nor U10002 (N_10002,N_9271,N_9539);
xor U10003 (N_10003,N_9204,N_9956);
nor U10004 (N_10004,N_9895,N_9420);
nand U10005 (N_10005,N_9086,N_9979);
nand U10006 (N_10006,N_9572,N_9862);
nand U10007 (N_10007,N_9334,N_9181);
nor U10008 (N_10008,N_9673,N_9132);
or U10009 (N_10009,N_9723,N_9958);
nor U10010 (N_10010,N_9412,N_9037);
xor U10011 (N_10011,N_9076,N_9292);
and U10012 (N_10012,N_9478,N_9495);
and U10013 (N_10013,N_9087,N_9146);
or U10014 (N_10014,N_9456,N_9735);
nor U10015 (N_10015,N_9343,N_9206);
nor U10016 (N_10016,N_9545,N_9325);
nand U10017 (N_10017,N_9254,N_9019);
and U10018 (N_10018,N_9971,N_9195);
or U10019 (N_10019,N_9494,N_9133);
and U10020 (N_10020,N_9027,N_9586);
nor U10021 (N_10021,N_9554,N_9661);
xnor U10022 (N_10022,N_9308,N_9916);
or U10023 (N_10023,N_9966,N_9319);
or U10024 (N_10024,N_9251,N_9237);
nand U10025 (N_10025,N_9876,N_9769);
nand U10026 (N_10026,N_9563,N_9279);
or U10027 (N_10027,N_9333,N_9025);
nand U10028 (N_10028,N_9622,N_9527);
and U10029 (N_10029,N_9134,N_9096);
or U10030 (N_10030,N_9187,N_9659);
nand U10031 (N_10031,N_9328,N_9843);
nand U10032 (N_10032,N_9380,N_9479);
or U10033 (N_10033,N_9561,N_9414);
and U10034 (N_10034,N_9141,N_9755);
nor U10035 (N_10035,N_9189,N_9826);
or U10036 (N_10036,N_9510,N_9612);
or U10037 (N_10037,N_9126,N_9063);
or U10038 (N_10038,N_9581,N_9831);
xnor U10039 (N_10039,N_9176,N_9579);
xnor U10040 (N_10040,N_9807,N_9764);
and U10041 (N_10041,N_9531,N_9792);
and U10042 (N_10042,N_9459,N_9587);
and U10043 (N_10043,N_9706,N_9908);
or U10044 (N_10044,N_9691,N_9144);
or U10045 (N_10045,N_9703,N_9613);
nor U10046 (N_10046,N_9508,N_9896);
and U10047 (N_10047,N_9178,N_9986);
nor U10048 (N_10048,N_9315,N_9159);
or U10049 (N_10049,N_9066,N_9633);
or U10050 (N_10050,N_9616,N_9120);
or U10051 (N_10051,N_9227,N_9145);
or U10052 (N_10052,N_9244,N_9467);
nand U10053 (N_10053,N_9926,N_9048);
xor U10054 (N_10054,N_9996,N_9083);
or U10055 (N_10055,N_9636,N_9101);
and U10056 (N_10056,N_9378,N_9737);
or U10057 (N_10057,N_9656,N_9443);
or U10058 (N_10058,N_9482,N_9270);
and U10059 (N_10059,N_9236,N_9310);
and U10060 (N_10060,N_9867,N_9839);
nand U10061 (N_10061,N_9719,N_9652);
and U10062 (N_10062,N_9232,N_9252);
and U10063 (N_10063,N_9742,N_9336);
xor U10064 (N_10064,N_9074,N_9782);
xor U10065 (N_10065,N_9611,N_9157);
xor U10066 (N_10066,N_9212,N_9199);
xor U10067 (N_10067,N_9142,N_9355);
or U10068 (N_10068,N_9722,N_9487);
nand U10069 (N_10069,N_9866,N_9920);
xnor U10070 (N_10070,N_9569,N_9477);
or U10071 (N_10071,N_9436,N_9033);
nand U10072 (N_10072,N_9677,N_9179);
or U10073 (N_10073,N_9624,N_9379);
xor U10074 (N_10074,N_9814,N_9103);
or U10075 (N_10075,N_9757,N_9762);
xnor U10076 (N_10076,N_9369,N_9701);
nand U10077 (N_10077,N_9752,N_9630);
nor U10078 (N_10078,N_9205,N_9714);
xnor U10079 (N_10079,N_9941,N_9562);
or U10080 (N_10080,N_9055,N_9286);
nor U10081 (N_10081,N_9389,N_9273);
xnor U10082 (N_10082,N_9517,N_9220);
nand U10083 (N_10083,N_9301,N_9243);
or U10084 (N_10084,N_9793,N_9054);
xnor U10085 (N_10085,N_9638,N_9897);
and U10086 (N_10086,N_9987,N_9363);
nor U10087 (N_10087,N_9289,N_9288);
and U10088 (N_10088,N_9760,N_9915);
and U10089 (N_10089,N_9365,N_9553);
xnor U10090 (N_10090,N_9679,N_9795);
or U10091 (N_10091,N_9909,N_9395);
and U10092 (N_10092,N_9257,N_9598);
and U10093 (N_10093,N_9667,N_9682);
nand U10094 (N_10094,N_9607,N_9291);
nor U10095 (N_10095,N_9448,N_9700);
or U10096 (N_10096,N_9344,N_9689);
nor U10097 (N_10097,N_9164,N_9560);
and U10098 (N_10098,N_9617,N_9771);
and U10099 (N_10099,N_9676,N_9842);
and U10100 (N_10100,N_9584,N_9687);
nor U10101 (N_10101,N_9422,N_9558);
nor U10102 (N_10102,N_9810,N_9768);
xor U10103 (N_10103,N_9637,N_9042);
and U10104 (N_10104,N_9609,N_9396);
and U10105 (N_10105,N_9634,N_9465);
nor U10106 (N_10106,N_9215,N_9258);
and U10107 (N_10107,N_9317,N_9829);
and U10108 (N_10108,N_9845,N_9648);
and U10109 (N_10109,N_9715,N_9969);
xnor U10110 (N_10110,N_9809,N_9529);
and U10111 (N_10111,N_9833,N_9654);
or U10112 (N_10112,N_9307,N_9946);
nand U10113 (N_10113,N_9403,N_9177);
or U10114 (N_10114,N_9248,N_9528);
or U10115 (N_10115,N_9321,N_9192);
nor U10116 (N_10116,N_9435,N_9658);
nor U10117 (N_10117,N_9547,N_9089);
xnor U10118 (N_10118,N_9770,N_9670);
or U10119 (N_10119,N_9975,N_9018);
nand U10120 (N_10120,N_9822,N_9499);
nand U10121 (N_10121,N_9062,N_9049);
or U10122 (N_10122,N_9841,N_9534);
nor U10123 (N_10123,N_9047,N_9107);
nor U10124 (N_10124,N_9774,N_9784);
nand U10125 (N_10125,N_9260,N_9031);
or U10126 (N_10126,N_9228,N_9098);
xor U10127 (N_10127,N_9549,N_9580);
or U10128 (N_10128,N_9441,N_9513);
or U10129 (N_10129,N_9022,N_9068);
or U10130 (N_10130,N_9827,N_9651);
or U10131 (N_10131,N_9813,N_9754);
or U10132 (N_10132,N_9102,N_9388);
and U10133 (N_10133,N_9836,N_9474);
xor U10134 (N_10134,N_9300,N_9129);
or U10135 (N_10135,N_9058,N_9850);
or U10136 (N_10136,N_9413,N_9469);
and U10137 (N_10137,N_9451,N_9263);
or U10138 (N_10138,N_9311,N_9932);
and U10139 (N_10139,N_9644,N_9811);
nand U10140 (N_10140,N_9353,N_9578);
nor U10141 (N_10141,N_9835,N_9590);
xor U10142 (N_10142,N_9997,N_9697);
and U10143 (N_10143,N_9340,N_9583);
or U10144 (N_10144,N_9978,N_9012);
or U10145 (N_10145,N_9500,N_9172);
or U10146 (N_10146,N_9858,N_9818);
and U10147 (N_10147,N_9766,N_9071);
and U10148 (N_10148,N_9429,N_9238);
and U10149 (N_10149,N_9819,N_9825);
nor U10150 (N_10150,N_9577,N_9543);
nand U10151 (N_10151,N_9116,N_9548);
nand U10152 (N_10152,N_9602,N_9625);
and U10153 (N_10153,N_9444,N_9026);
xor U10154 (N_10154,N_9015,N_9377);
nand U10155 (N_10155,N_9555,N_9806);
xor U10156 (N_10156,N_9475,N_9029);
nand U10157 (N_10157,N_9724,N_9837);
and U10158 (N_10158,N_9155,N_9610);
nor U10159 (N_10159,N_9461,N_9044);
and U10160 (N_10160,N_9373,N_9733);
nand U10161 (N_10161,N_9203,N_9851);
nand U10162 (N_10162,N_9940,N_9118);
nor U10163 (N_10163,N_9886,N_9032);
and U10164 (N_10164,N_9955,N_9171);
xor U10165 (N_10165,N_9211,N_9681);
nand U10166 (N_10166,N_9174,N_9471);
and U10167 (N_10167,N_9405,N_9943);
nand U10168 (N_10168,N_9949,N_9326);
nand U10169 (N_10169,N_9481,N_9374);
or U10170 (N_10170,N_9226,N_9900);
and U10171 (N_10171,N_9341,N_9386);
nand U10172 (N_10172,N_9387,N_9162);
nor U10173 (N_10173,N_9596,N_9184);
xor U10174 (N_10174,N_9599,N_9158);
nand U10175 (N_10175,N_9967,N_9566);
or U10176 (N_10176,N_9834,N_9092);
nor U10177 (N_10177,N_9650,N_9128);
nand U10178 (N_10178,N_9692,N_9445);
xnor U10179 (N_10179,N_9284,N_9964);
nand U10180 (N_10180,N_9193,N_9780);
nand U10181 (N_10181,N_9017,N_9295);
nor U10182 (N_10182,N_9143,N_9030);
or U10183 (N_10183,N_9261,N_9385);
xor U10184 (N_10184,N_9246,N_9139);
nand U10185 (N_10185,N_9889,N_9484);
and U10186 (N_10186,N_9117,N_9269);
or U10187 (N_10187,N_9789,N_9803);
or U10188 (N_10188,N_9530,N_9537);
or U10189 (N_10189,N_9954,N_9135);
nor U10190 (N_10190,N_9446,N_9067);
xnor U10191 (N_10191,N_9253,N_9983);
and U10192 (N_10192,N_9888,N_9398);
xnor U10193 (N_10193,N_9400,N_9699);
or U10194 (N_10194,N_9472,N_9170);
nand U10195 (N_10195,N_9546,N_9277);
and U10196 (N_10196,N_9797,N_9005);
nor U10197 (N_10197,N_9702,N_9427);
nand U10198 (N_10198,N_9191,N_9007);
xor U10199 (N_10199,N_9927,N_9993);
nand U10200 (N_10200,N_9592,N_9351);
nor U10201 (N_10201,N_9753,N_9108);
nor U10202 (N_10202,N_9939,N_9914);
xnor U10203 (N_10203,N_9938,N_9731);
and U10204 (N_10204,N_9864,N_9505);
and U10205 (N_10205,N_9815,N_9669);
xnor U10206 (N_10206,N_9423,N_9274);
xor U10207 (N_10207,N_9588,N_9210);
xnor U10208 (N_10208,N_9382,N_9984);
xor U10209 (N_10209,N_9272,N_9114);
or U10210 (N_10210,N_9163,N_9557);
nand U10211 (N_10211,N_9934,N_9194);
nor U10212 (N_10212,N_9875,N_9235);
nand U10213 (N_10213,N_9614,N_9840);
or U10214 (N_10214,N_9173,N_9240);
nand U10215 (N_10215,N_9416,N_9544);
or U10216 (N_10216,N_9898,N_9570);
nand U10217 (N_10217,N_9437,N_9974);
nor U10218 (N_10218,N_9830,N_9259);
xnor U10219 (N_10219,N_9621,N_9631);
xor U10220 (N_10220,N_9094,N_9600);
or U10221 (N_10221,N_9462,N_9642);
and U10222 (N_10222,N_9090,N_9904);
nand U10223 (N_10223,N_9404,N_9485);
or U10224 (N_10224,N_9454,N_9911);
nand U10225 (N_10225,N_9838,N_9804);
nor U10226 (N_10226,N_9294,N_9216);
xnor U10227 (N_10227,N_9628,N_9359);
nor U10228 (N_10228,N_9305,N_9748);
and U10229 (N_10229,N_9758,N_9347);
xnor U10230 (N_10230,N_9053,N_9698);
nor U10231 (N_10231,N_9736,N_9696);
and U10232 (N_10232,N_9933,N_9313);
and U10233 (N_10233,N_9085,N_9980);
nand U10234 (N_10234,N_9734,N_9917);
nor U10235 (N_10235,N_9705,N_9879);
and U10236 (N_10236,N_9104,N_9945);
nor U10237 (N_10237,N_9779,N_9937);
or U10238 (N_10238,N_9823,N_9364);
or U10239 (N_10239,N_9410,N_9419);
and U10240 (N_10240,N_9952,N_9013);
nor U10241 (N_10241,N_9618,N_9957);
or U10242 (N_10242,N_9641,N_9185);
and U10243 (N_10243,N_9525,N_9501);
and U10244 (N_10244,N_9418,N_9121);
and U10245 (N_10245,N_9573,N_9947);
xor U10246 (N_10246,N_9093,N_9368);
nand U10247 (N_10247,N_9111,N_9148);
nor U10248 (N_10248,N_9992,N_9564);
nand U10249 (N_10249,N_9283,N_9848);
or U10250 (N_10250,N_9538,N_9002);
nor U10251 (N_10251,N_9685,N_9824);
and U10252 (N_10252,N_9084,N_9421);
xor U10253 (N_10253,N_9516,N_9524);
and U10254 (N_10254,N_9514,N_9710);
and U10255 (N_10255,N_9518,N_9653);
or U10256 (N_10256,N_9693,N_9629);
or U10257 (N_10257,N_9891,N_9690);
xnor U10258 (N_10258,N_9728,N_9304);
nand U10259 (N_10259,N_9360,N_9276);
or U10260 (N_10260,N_9765,N_9894);
nand U10261 (N_10261,N_9990,N_9161);
nor U10262 (N_10262,N_9038,N_9605);
and U10263 (N_10263,N_9646,N_9202);
nand U10264 (N_10264,N_9097,N_9490);
or U10265 (N_10265,N_9739,N_9493);
xnor U10266 (N_10266,N_9239,N_9250);
nand U10267 (N_10267,N_9371,N_9079);
nor U10268 (N_10268,N_9275,N_9738);
nand U10269 (N_10269,N_9040,N_9781);
xnor U10270 (N_10270,N_9535,N_9854);
nor U10271 (N_10271,N_9608,N_9151);
and U10272 (N_10272,N_9794,N_9775);
nand U10273 (N_10273,N_9010,N_9391);
and U10274 (N_10274,N_9601,N_9893);
nand U10275 (N_10275,N_9743,N_9455);
or U10276 (N_10276,N_9401,N_9298);
nand U10277 (N_10277,N_9623,N_9082);
and U10278 (N_10278,N_9870,N_9167);
nor U10279 (N_10279,N_9282,N_9376);
or U10280 (N_10280,N_9496,N_9683);
xor U10281 (N_10281,N_9776,N_9965);
nor U10282 (N_10282,N_9995,N_9973);
or U10283 (N_10283,N_9209,N_9878);
nor U10284 (N_10284,N_9483,N_9571);
xnor U10285 (N_10285,N_9046,N_9532);
or U10286 (N_10286,N_9664,N_9309);
and U10287 (N_10287,N_9928,N_9817);
nand U10288 (N_10288,N_9709,N_9004);
and U10289 (N_10289,N_9882,N_9657);
or U10290 (N_10290,N_9712,N_9799);
and U10291 (N_10291,N_9241,N_9064);
nor U10292 (N_10292,N_9988,N_9660);
xnor U10293 (N_10293,N_9783,N_9217);
nor U10294 (N_10294,N_9856,N_9585);
xnor U10295 (N_10295,N_9907,N_9632);
nor U10296 (N_10296,N_9113,N_9680);
nor U10297 (N_10297,N_9065,N_9931);
nand U10298 (N_10298,N_9218,N_9798);
nand U10299 (N_10299,N_9960,N_9922);
xnor U10300 (N_10300,N_9968,N_9077);
or U10301 (N_10301,N_9402,N_9725);
nor U10302 (N_10302,N_9392,N_9778);
nand U10303 (N_10303,N_9749,N_9727);
or U10304 (N_10304,N_9338,N_9078);
or U10305 (N_10305,N_9221,N_9999);
and U10306 (N_10306,N_9721,N_9497);
or U10307 (N_10307,N_9520,N_9375);
xnor U10308 (N_10308,N_9884,N_9635);
nor U10309 (N_10309,N_9816,N_9464);
xor U10310 (N_10310,N_9846,N_9873);
nor U10311 (N_10311,N_9384,N_9383);
xnor U10312 (N_10312,N_9515,N_9675);
nor U10313 (N_10313,N_9639,N_9109);
and U10314 (N_10314,N_9166,N_9045);
xnor U10315 (N_10315,N_9708,N_9498);
nand U10316 (N_10316,N_9293,N_9339);
and U10317 (N_10317,N_9844,N_9224);
or U10318 (N_10318,N_9352,N_9821);
nand U10319 (N_10319,N_9565,N_9009);
nor U10320 (N_10320,N_9320,N_9615);
or U10321 (N_10321,N_9910,N_9381);
nand U10322 (N_10322,N_9869,N_9024);
nand U10323 (N_10323,N_9741,N_9440);
xnor U10324 (N_10324,N_9759,N_9367);
nor U10325 (N_10325,N_9672,N_9242);
xnor U10326 (N_10326,N_9099,N_9366);
nor U10327 (N_10327,N_9688,N_9589);
and U10328 (N_10328,N_9245,N_9439);
and U10329 (N_10329,N_9329,N_9332);
nor U10330 (N_10330,N_9393,N_9732);
nor U10331 (N_10331,N_9105,N_9591);
xnor U10332 (N_10332,N_9785,N_9188);
nor U10333 (N_10333,N_9767,N_9021);
nor U10334 (N_10334,N_9963,N_9847);
xor U10335 (N_10335,N_9213,N_9711);
xnor U10336 (N_10336,N_9521,N_9372);
nand U10337 (N_10337,N_9713,N_9020);
and U10338 (N_10338,N_9407,N_9674);
or U10339 (N_10339,N_9786,N_9137);
nor U10340 (N_10340,N_9503,N_9507);
and U10341 (N_10341,N_9504,N_9057);
and U10342 (N_10342,N_9290,N_9885);
nand U10343 (N_10343,N_9169,N_9417);
and U10344 (N_10344,N_9492,N_9265);
nor U10345 (N_10345,N_9060,N_9249);
or U10346 (N_10346,N_9299,N_9935);
or U10347 (N_10347,N_9744,N_9604);
xor U10348 (N_10348,N_9871,N_9136);
or U10349 (N_10349,N_9576,N_9750);
and U10350 (N_10350,N_9686,N_9175);
nor U10351 (N_10351,N_9695,N_9281);
or U10352 (N_10352,N_9800,N_9346);
or U10353 (N_10353,N_9944,N_9468);
xnor U10354 (N_10354,N_9302,N_9930);
nor U10355 (N_10355,N_9627,N_9805);
nor U10356 (N_10356,N_9912,N_9594);
or U10357 (N_10357,N_9409,N_9522);
nand U10358 (N_10358,N_9287,N_9154);
xnor U10359 (N_10359,N_9153,N_9665);
or U10360 (N_10360,N_9394,N_9466);
xnor U10361 (N_10361,N_9540,N_9948);
xor U10362 (N_10362,N_9460,N_9168);
nand U10363 (N_10363,N_9533,N_9354);
xor U10364 (N_10364,N_9881,N_9165);
nand U10365 (N_10365,N_9953,N_9088);
nand U10366 (N_10366,N_9863,N_9214);
and U10367 (N_10367,N_9223,N_9905);
nand U10368 (N_10368,N_9509,N_9595);
or U10369 (N_10369,N_9337,N_9458);
and U10370 (N_10370,N_9684,N_9014);
nor U10371 (N_10371,N_9853,N_9619);
or U10372 (N_10372,N_9432,N_9425);
and U10373 (N_10373,N_9463,N_9450);
and U10374 (N_10374,N_9150,N_9050);
and U10375 (N_10375,N_9131,N_9929);
nand U10376 (N_10376,N_9647,N_9707);
and U10377 (N_10377,N_9230,N_9872);
nand U10378 (N_10378,N_9790,N_9551);
nor U10379 (N_10379,N_9156,N_9991);
nor U10380 (N_10380,N_9011,N_9470);
and U10381 (N_10381,N_9716,N_9397);
nand U10382 (N_10382,N_9312,N_9149);
xnor U10383 (N_10383,N_9812,N_9874);
nor U10384 (N_10384,N_9262,N_9491);
nand U10385 (N_10385,N_9222,N_9314);
xor U10386 (N_10386,N_9303,N_9138);
xor U10387 (N_10387,N_9852,N_9036);
or U10388 (N_10388,N_9075,N_9962);
xnor U10389 (N_10389,N_9606,N_9070);
or U10390 (N_10390,N_9919,N_9977);
or U10391 (N_10391,N_9903,N_9358);
and U10392 (N_10392,N_9219,N_9772);
or U10393 (N_10393,N_9523,N_9480);
xor U10394 (N_10394,N_9072,N_9902);
or U10395 (N_10395,N_9730,N_9649);
or U10396 (N_10396,N_9296,N_9006);
xor U10397 (N_10397,N_9003,N_9008);
nor U10398 (N_10398,N_9457,N_9620);
xor U10399 (N_10399,N_9655,N_9438);
or U10400 (N_10400,N_9849,N_9023);
and U10401 (N_10401,N_9428,N_9122);
or U10402 (N_10402,N_9115,N_9453);
or U10403 (N_10403,N_9147,N_9473);
or U10404 (N_10404,N_9626,N_9411);
nor U10405 (N_10405,N_9593,N_9119);
nor U10406 (N_10406,N_9541,N_9056);
and U10407 (N_10407,N_9556,N_9645);
or U10408 (N_10408,N_9582,N_9180);
and U10409 (N_10409,N_9890,N_9802);
or U10410 (N_10410,N_9127,N_9511);
nand U10411 (N_10411,N_9860,N_9322);
nand U10412 (N_10412,N_9704,N_9868);
xor U10413 (N_10413,N_9324,N_9921);
and U10414 (N_10414,N_9406,N_9415);
or U10415 (N_10415,N_9452,N_9865);
and U10416 (N_10416,N_9348,N_9125);
xor U10417 (N_10417,N_9801,N_9526);
nand U10418 (N_10418,N_9362,N_9390);
nand U10419 (N_10419,N_9186,N_9536);
and U10420 (N_10420,N_9773,N_9791);
xor U10421 (N_10421,N_9820,N_9855);
nor U10422 (N_10422,N_9502,N_9316);
or U10423 (N_10423,N_9361,N_9640);
xnor U10424 (N_10424,N_9357,N_9198);
and U10425 (N_10425,N_9208,N_9512);
xnor U10426 (N_10426,N_9597,N_9740);
nor U10427 (N_10427,N_9080,N_9035);
or U10428 (N_10428,N_9430,N_9777);
or U10429 (N_10429,N_9255,N_9519);
and U10430 (N_10430,N_9488,N_9747);
nor U10431 (N_10431,N_9370,N_9233);
and U10432 (N_10432,N_9106,N_9892);
nor U10433 (N_10433,N_9746,N_9123);
or U10434 (N_10434,N_9000,N_9350);
nor U10435 (N_10435,N_9559,N_9756);
or U10436 (N_10436,N_9323,N_9981);
xor U10437 (N_10437,N_9994,N_9745);
nand U10438 (N_10438,N_9061,N_9972);
xor U10439 (N_10439,N_9160,N_9726);
or U10440 (N_10440,N_9506,N_9998);
xor U10441 (N_10441,N_9331,N_9399);
nor U10442 (N_10442,N_9280,N_9913);
and U10443 (N_10443,N_9936,N_9923);
xnor U10444 (N_10444,N_9486,N_9051);
nand U10445 (N_10445,N_9069,N_9426);
and U10446 (N_10446,N_9552,N_9318);
or U10447 (N_10447,N_9433,N_9717);
xnor U10448 (N_10448,N_9883,N_9662);
xor U10449 (N_10449,N_9231,N_9666);
nor U10450 (N_10450,N_9196,N_9942);
nand U10451 (N_10451,N_9130,N_9285);
and U10452 (N_10452,N_9190,N_9918);
nor U10453 (N_10453,N_9110,N_9267);
and U10454 (N_10454,N_9542,N_9976);
nand U10455 (N_10455,N_9330,N_9112);
nor U10456 (N_10456,N_9229,N_9345);
xnor U10457 (N_10457,N_9266,N_9729);
or U10458 (N_10458,N_9268,N_9901);
or U10459 (N_10459,N_9671,N_9041);
and U10460 (N_10460,N_9906,N_9574);
or U10461 (N_10461,N_9476,N_9264);
nand U10462 (N_10462,N_9924,N_9751);
or U10463 (N_10463,N_9028,N_9124);
nand U10464 (N_10464,N_9039,N_9349);
or U10465 (N_10465,N_9073,N_9887);
nand U10466 (N_10466,N_9408,N_9550);
and U10467 (N_10467,N_9761,N_9763);
xor U10468 (N_10468,N_9234,N_9925);
or U10469 (N_10469,N_9183,N_9016);
nand U10470 (N_10470,N_9052,N_9297);
xnor U10471 (N_10471,N_9356,N_9034);
nor U10472 (N_10472,N_9663,N_9951);
xnor U10473 (N_10473,N_9095,N_9950);
xor U10474 (N_10474,N_9828,N_9059);
nor U10475 (N_10475,N_9335,N_9643);
xor U10476 (N_10476,N_9197,N_9899);
nor U10477 (N_10477,N_9140,N_9152);
nor U10478 (N_10478,N_9668,N_9001);
xor U10479 (N_10479,N_9256,N_9787);
nand U10480 (N_10480,N_9718,N_9877);
nand U10481 (N_10481,N_9694,N_9424);
nand U10482 (N_10482,N_9788,N_9567);
nand U10483 (N_10483,N_9225,N_9327);
and U10484 (N_10484,N_9880,N_9603);
and U10485 (N_10485,N_9489,N_9278);
and U10486 (N_10486,N_9449,N_9857);
nand U10487 (N_10487,N_9575,N_9434);
nand U10488 (N_10488,N_9796,N_9442);
and U10489 (N_10489,N_9182,N_9568);
and U10490 (N_10490,N_9091,N_9678);
and U10491 (N_10491,N_9342,N_9043);
and U10492 (N_10492,N_9861,N_9985);
and U10493 (N_10493,N_9970,N_9447);
nor U10494 (N_10494,N_9431,N_9247);
nor U10495 (N_10495,N_9200,N_9100);
nor U10496 (N_10496,N_9959,N_9306);
xnor U10497 (N_10497,N_9961,N_9982);
nand U10498 (N_10498,N_9081,N_9207);
or U10499 (N_10499,N_9832,N_9808);
or U10500 (N_10500,N_9803,N_9563);
or U10501 (N_10501,N_9264,N_9854);
xnor U10502 (N_10502,N_9535,N_9383);
nor U10503 (N_10503,N_9140,N_9510);
or U10504 (N_10504,N_9131,N_9029);
or U10505 (N_10505,N_9798,N_9944);
and U10506 (N_10506,N_9616,N_9649);
nand U10507 (N_10507,N_9184,N_9137);
and U10508 (N_10508,N_9170,N_9135);
nor U10509 (N_10509,N_9981,N_9773);
xor U10510 (N_10510,N_9202,N_9919);
nand U10511 (N_10511,N_9270,N_9808);
and U10512 (N_10512,N_9199,N_9961);
and U10513 (N_10513,N_9629,N_9107);
nor U10514 (N_10514,N_9294,N_9154);
xor U10515 (N_10515,N_9647,N_9178);
and U10516 (N_10516,N_9721,N_9078);
xnor U10517 (N_10517,N_9789,N_9097);
and U10518 (N_10518,N_9114,N_9674);
nor U10519 (N_10519,N_9348,N_9445);
and U10520 (N_10520,N_9846,N_9578);
xor U10521 (N_10521,N_9689,N_9525);
xnor U10522 (N_10522,N_9867,N_9868);
nor U10523 (N_10523,N_9235,N_9217);
nand U10524 (N_10524,N_9891,N_9817);
nand U10525 (N_10525,N_9352,N_9273);
xor U10526 (N_10526,N_9444,N_9708);
nor U10527 (N_10527,N_9956,N_9958);
nand U10528 (N_10528,N_9937,N_9166);
nor U10529 (N_10529,N_9229,N_9040);
or U10530 (N_10530,N_9423,N_9713);
or U10531 (N_10531,N_9884,N_9414);
or U10532 (N_10532,N_9272,N_9678);
nor U10533 (N_10533,N_9608,N_9861);
nor U10534 (N_10534,N_9477,N_9391);
or U10535 (N_10535,N_9427,N_9271);
nand U10536 (N_10536,N_9411,N_9281);
and U10537 (N_10537,N_9073,N_9757);
nor U10538 (N_10538,N_9674,N_9131);
and U10539 (N_10539,N_9123,N_9352);
nor U10540 (N_10540,N_9205,N_9093);
nor U10541 (N_10541,N_9219,N_9189);
or U10542 (N_10542,N_9758,N_9774);
and U10543 (N_10543,N_9850,N_9353);
nand U10544 (N_10544,N_9820,N_9977);
nand U10545 (N_10545,N_9992,N_9493);
and U10546 (N_10546,N_9765,N_9804);
xnor U10547 (N_10547,N_9163,N_9055);
nor U10548 (N_10548,N_9267,N_9870);
nand U10549 (N_10549,N_9927,N_9876);
nand U10550 (N_10550,N_9959,N_9054);
nor U10551 (N_10551,N_9466,N_9200);
and U10552 (N_10552,N_9094,N_9684);
nor U10553 (N_10553,N_9887,N_9024);
nor U10554 (N_10554,N_9581,N_9412);
and U10555 (N_10555,N_9078,N_9155);
and U10556 (N_10556,N_9010,N_9358);
and U10557 (N_10557,N_9346,N_9103);
or U10558 (N_10558,N_9070,N_9211);
nor U10559 (N_10559,N_9060,N_9610);
nand U10560 (N_10560,N_9357,N_9640);
or U10561 (N_10561,N_9418,N_9305);
nand U10562 (N_10562,N_9829,N_9144);
and U10563 (N_10563,N_9470,N_9501);
xnor U10564 (N_10564,N_9842,N_9435);
xnor U10565 (N_10565,N_9624,N_9931);
nor U10566 (N_10566,N_9344,N_9125);
nand U10567 (N_10567,N_9997,N_9198);
and U10568 (N_10568,N_9158,N_9890);
xor U10569 (N_10569,N_9810,N_9694);
nand U10570 (N_10570,N_9580,N_9665);
or U10571 (N_10571,N_9687,N_9946);
xor U10572 (N_10572,N_9603,N_9953);
nor U10573 (N_10573,N_9716,N_9010);
and U10574 (N_10574,N_9317,N_9318);
xor U10575 (N_10575,N_9038,N_9753);
xor U10576 (N_10576,N_9238,N_9850);
and U10577 (N_10577,N_9707,N_9761);
or U10578 (N_10578,N_9007,N_9491);
or U10579 (N_10579,N_9078,N_9257);
xor U10580 (N_10580,N_9757,N_9517);
nor U10581 (N_10581,N_9963,N_9406);
nor U10582 (N_10582,N_9755,N_9968);
xor U10583 (N_10583,N_9227,N_9620);
xor U10584 (N_10584,N_9805,N_9578);
xor U10585 (N_10585,N_9162,N_9453);
xnor U10586 (N_10586,N_9851,N_9717);
and U10587 (N_10587,N_9228,N_9511);
nand U10588 (N_10588,N_9457,N_9335);
xor U10589 (N_10589,N_9195,N_9288);
nand U10590 (N_10590,N_9938,N_9614);
nand U10591 (N_10591,N_9095,N_9511);
or U10592 (N_10592,N_9967,N_9443);
or U10593 (N_10593,N_9664,N_9938);
or U10594 (N_10594,N_9877,N_9358);
and U10595 (N_10595,N_9116,N_9673);
nand U10596 (N_10596,N_9859,N_9094);
and U10597 (N_10597,N_9952,N_9883);
xnor U10598 (N_10598,N_9404,N_9158);
and U10599 (N_10599,N_9128,N_9645);
nand U10600 (N_10600,N_9626,N_9824);
nand U10601 (N_10601,N_9519,N_9041);
nor U10602 (N_10602,N_9360,N_9878);
xor U10603 (N_10603,N_9166,N_9155);
or U10604 (N_10604,N_9192,N_9129);
or U10605 (N_10605,N_9792,N_9867);
nand U10606 (N_10606,N_9582,N_9978);
and U10607 (N_10607,N_9942,N_9289);
or U10608 (N_10608,N_9896,N_9094);
or U10609 (N_10609,N_9720,N_9689);
nand U10610 (N_10610,N_9293,N_9808);
nor U10611 (N_10611,N_9966,N_9362);
xnor U10612 (N_10612,N_9945,N_9690);
nor U10613 (N_10613,N_9583,N_9088);
or U10614 (N_10614,N_9631,N_9243);
and U10615 (N_10615,N_9873,N_9831);
or U10616 (N_10616,N_9829,N_9593);
xor U10617 (N_10617,N_9496,N_9615);
and U10618 (N_10618,N_9424,N_9344);
or U10619 (N_10619,N_9819,N_9370);
nand U10620 (N_10620,N_9047,N_9661);
xnor U10621 (N_10621,N_9513,N_9717);
or U10622 (N_10622,N_9922,N_9850);
or U10623 (N_10623,N_9405,N_9438);
and U10624 (N_10624,N_9245,N_9672);
or U10625 (N_10625,N_9610,N_9190);
nand U10626 (N_10626,N_9067,N_9265);
xnor U10627 (N_10627,N_9232,N_9202);
nand U10628 (N_10628,N_9220,N_9856);
or U10629 (N_10629,N_9537,N_9061);
nor U10630 (N_10630,N_9308,N_9603);
or U10631 (N_10631,N_9961,N_9593);
and U10632 (N_10632,N_9907,N_9273);
or U10633 (N_10633,N_9061,N_9072);
nor U10634 (N_10634,N_9179,N_9980);
nand U10635 (N_10635,N_9784,N_9926);
xnor U10636 (N_10636,N_9771,N_9826);
xnor U10637 (N_10637,N_9845,N_9321);
nand U10638 (N_10638,N_9004,N_9268);
or U10639 (N_10639,N_9245,N_9348);
and U10640 (N_10640,N_9298,N_9139);
nand U10641 (N_10641,N_9960,N_9472);
xnor U10642 (N_10642,N_9084,N_9781);
nor U10643 (N_10643,N_9810,N_9281);
and U10644 (N_10644,N_9253,N_9002);
nor U10645 (N_10645,N_9723,N_9461);
xor U10646 (N_10646,N_9243,N_9727);
nand U10647 (N_10647,N_9113,N_9116);
xnor U10648 (N_10648,N_9393,N_9745);
xor U10649 (N_10649,N_9963,N_9619);
nand U10650 (N_10650,N_9903,N_9471);
nand U10651 (N_10651,N_9581,N_9891);
or U10652 (N_10652,N_9401,N_9468);
xnor U10653 (N_10653,N_9795,N_9271);
or U10654 (N_10654,N_9546,N_9335);
nor U10655 (N_10655,N_9191,N_9942);
nor U10656 (N_10656,N_9256,N_9364);
nor U10657 (N_10657,N_9717,N_9533);
xnor U10658 (N_10658,N_9350,N_9418);
nand U10659 (N_10659,N_9254,N_9102);
xor U10660 (N_10660,N_9355,N_9494);
nand U10661 (N_10661,N_9027,N_9175);
or U10662 (N_10662,N_9568,N_9129);
or U10663 (N_10663,N_9083,N_9296);
nor U10664 (N_10664,N_9416,N_9258);
xnor U10665 (N_10665,N_9715,N_9423);
xnor U10666 (N_10666,N_9291,N_9878);
and U10667 (N_10667,N_9561,N_9480);
xnor U10668 (N_10668,N_9550,N_9222);
nor U10669 (N_10669,N_9577,N_9558);
or U10670 (N_10670,N_9405,N_9255);
or U10671 (N_10671,N_9943,N_9679);
xnor U10672 (N_10672,N_9021,N_9575);
nor U10673 (N_10673,N_9715,N_9328);
or U10674 (N_10674,N_9647,N_9595);
or U10675 (N_10675,N_9448,N_9452);
or U10676 (N_10676,N_9486,N_9505);
nand U10677 (N_10677,N_9213,N_9710);
nor U10678 (N_10678,N_9095,N_9208);
or U10679 (N_10679,N_9161,N_9553);
xnor U10680 (N_10680,N_9247,N_9494);
or U10681 (N_10681,N_9588,N_9885);
xor U10682 (N_10682,N_9939,N_9324);
xor U10683 (N_10683,N_9409,N_9915);
nor U10684 (N_10684,N_9765,N_9006);
and U10685 (N_10685,N_9604,N_9678);
xor U10686 (N_10686,N_9132,N_9225);
nor U10687 (N_10687,N_9195,N_9941);
xnor U10688 (N_10688,N_9653,N_9596);
and U10689 (N_10689,N_9544,N_9935);
nor U10690 (N_10690,N_9645,N_9639);
and U10691 (N_10691,N_9047,N_9917);
and U10692 (N_10692,N_9266,N_9144);
and U10693 (N_10693,N_9587,N_9844);
nand U10694 (N_10694,N_9237,N_9258);
or U10695 (N_10695,N_9187,N_9376);
and U10696 (N_10696,N_9726,N_9563);
xor U10697 (N_10697,N_9039,N_9255);
and U10698 (N_10698,N_9048,N_9976);
nor U10699 (N_10699,N_9547,N_9541);
and U10700 (N_10700,N_9879,N_9553);
xnor U10701 (N_10701,N_9645,N_9259);
nand U10702 (N_10702,N_9307,N_9698);
nor U10703 (N_10703,N_9868,N_9048);
nand U10704 (N_10704,N_9139,N_9452);
and U10705 (N_10705,N_9363,N_9821);
and U10706 (N_10706,N_9396,N_9006);
nor U10707 (N_10707,N_9823,N_9782);
xor U10708 (N_10708,N_9523,N_9784);
xnor U10709 (N_10709,N_9189,N_9728);
nand U10710 (N_10710,N_9265,N_9707);
nor U10711 (N_10711,N_9684,N_9627);
and U10712 (N_10712,N_9119,N_9622);
nand U10713 (N_10713,N_9568,N_9817);
or U10714 (N_10714,N_9566,N_9344);
and U10715 (N_10715,N_9652,N_9940);
nor U10716 (N_10716,N_9311,N_9039);
xnor U10717 (N_10717,N_9794,N_9415);
or U10718 (N_10718,N_9668,N_9302);
and U10719 (N_10719,N_9785,N_9044);
or U10720 (N_10720,N_9456,N_9717);
nor U10721 (N_10721,N_9061,N_9727);
nand U10722 (N_10722,N_9571,N_9213);
nand U10723 (N_10723,N_9721,N_9310);
and U10724 (N_10724,N_9633,N_9328);
nand U10725 (N_10725,N_9797,N_9882);
or U10726 (N_10726,N_9342,N_9301);
xnor U10727 (N_10727,N_9068,N_9968);
and U10728 (N_10728,N_9896,N_9086);
nor U10729 (N_10729,N_9307,N_9996);
xor U10730 (N_10730,N_9683,N_9625);
or U10731 (N_10731,N_9325,N_9125);
xor U10732 (N_10732,N_9955,N_9760);
or U10733 (N_10733,N_9793,N_9623);
nor U10734 (N_10734,N_9395,N_9885);
xor U10735 (N_10735,N_9490,N_9268);
nor U10736 (N_10736,N_9941,N_9732);
xor U10737 (N_10737,N_9906,N_9592);
or U10738 (N_10738,N_9832,N_9091);
or U10739 (N_10739,N_9008,N_9147);
or U10740 (N_10740,N_9303,N_9892);
xnor U10741 (N_10741,N_9017,N_9387);
nor U10742 (N_10742,N_9755,N_9904);
or U10743 (N_10743,N_9471,N_9115);
xnor U10744 (N_10744,N_9509,N_9037);
nor U10745 (N_10745,N_9564,N_9285);
xor U10746 (N_10746,N_9144,N_9455);
nand U10747 (N_10747,N_9235,N_9055);
xnor U10748 (N_10748,N_9343,N_9389);
or U10749 (N_10749,N_9175,N_9993);
nand U10750 (N_10750,N_9601,N_9163);
and U10751 (N_10751,N_9864,N_9580);
nor U10752 (N_10752,N_9573,N_9759);
xor U10753 (N_10753,N_9373,N_9928);
or U10754 (N_10754,N_9633,N_9063);
nand U10755 (N_10755,N_9244,N_9451);
nor U10756 (N_10756,N_9870,N_9441);
nand U10757 (N_10757,N_9847,N_9421);
or U10758 (N_10758,N_9797,N_9455);
xnor U10759 (N_10759,N_9168,N_9286);
nand U10760 (N_10760,N_9245,N_9772);
and U10761 (N_10761,N_9504,N_9999);
nor U10762 (N_10762,N_9491,N_9446);
or U10763 (N_10763,N_9292,N_9471);
nand U10764 (N_10764,N_9393,N_9881);
nor U10765 (N_10765,N_9545,N_9073);
and U10766 (N_10766,N_9003,N_9512);
nor U10767 (N_10767,N_9409,N_9837);
and U10768 (N_10768,N_9653,N_9423);
xnor U10769 (N_10769,N_9012,N_9538);
and U10770 (N_10770,N_9047,N_9702);
nor U10771 (N_10771,N_9448,N_9558);
and U10772 (N_10772,N_9328,N_9695);
or U10773 (N_10773,N_9045,N_9057);
and U10774 (N_10774,N_9149,N_9783);
or U10775 (N_10775,N_9775,N_9052);
nor U10776 (N_10776,N_9829,N_9197);
or U10777 (N_10777,N_9747,N_9410);
and U10778 (N_10778,N_9549,N_9782);
nand U10779 (N_10779,N_9777,N_9382);
and U10780 (N_10780,N_9657,N_9946);
xor U10781 (N_10781,N_9694,N_9350);
and U10782 (N_10782,N_9820,N_9569);
xor U10783 (N_10783,N_9197,N_9427);
and U10784 (N_10784,N_9058,N_9680);
nand U10785 (N_10785,N_9434,N_9964);
xor U10786 (N_10786,N_9464,N_9498);
nand U10787 (N_10787,N_9827,N_9015);
nor U10788 (N_10788,N_9960,N_9658);
or U10789 (N_10789,N_9022,N_9221);
or U10790 (N_10790,N_9644,N_9819);
or U10791 (N_10791,N_9245,N_9576);
or U10792 (N_10792,N_9194,N_9007);
nand U10793 (N_10793,N_9196,N_9130);
nor U10794 (N_10794,N_9082,N_9165);
nand U10795 (N_10795,N_9385,N_9044);
nor U10796 (N_10796,N_9790,N_9896);
nor U10797 (N_10797,N_9175,N_9695);
xor U10798 (N_10798,N_9355,N_9336);
xor U10799 (N_10799,N_9532,N_9877);
or U10800 (N_10800,N_9602,N_9914);
and U10801 (N_10801,N_9194,N_9293);
xnor U10802 (N_10802,N_9564,N_9085);
nor U10803 (N_10803,N_9904,N_9265);
nor U10804 (N_10804,N_9556,N_9049);
nand U10805 (N_10805,N_9032,N_9598);
xnor U10806 (N_10806,N_9996,N_9402);
nor U10807 (N_10807,N_9141,N_9327);
or U10808 (N_10808,N_9163,N_9427);
nor U10809 (N_10809,N_9706,N_9254);
nor U10810 (N_10810,N_9218,N_9339);
nor U10811 (N_10811,N_9916,N_9880);
xnor U10812 (N_10812,N_9623,N_9878);
xnor U10813 (N_10813,N_9983,N_9495);
xnor U10814 (N_10814,N_9255,N_9909);
nand U10815 (N_10815,N_9656,N_9364);
nor U10816 (N_10816,N_9241,N_9343);
or U10817 (N_10817,N_9281,N_9549);
nor U10818 (N_10818,N_9050,N_9966);
and U10819 (N_10819,N_9025,N_9335);
and U10820 (N_10820,N_9491,N_9131);
nand U10821 (N_10821,N_9635,N_9707);
or U10822 (N_10822,N_9983,N_9329);
and U10823 (N_10823,N_9821,N_9947);
or U10824 (N_10824,N_9838,N_9591);
and U10825 (N_10825,N_9261,N_9705);
nand U10826 (N_10826,N_9918,N_9792);
nand U10827 (N_10827,N_9996,N_9769);
and U10828 (N_10828,N_9826,N_9992);
xor U10829 (N_10829,N_9045,N_9994);
nand U10830 (N_10830,N_9410,N_9776);
xor U10831 (N_10831,N_9999,N_9418);
nand U10832 (N_10832,N_9931,N_9706);
and U10833 (N_10833,N_9303,N_9409);
and U10834 (N_10834,N_9637,N_9234);
xnor U10835 (N_10835,N_9920,N_9325);
nor U10836 (N_10836,N_9180,N_9177);
nand U10837 (N_10837,N_9073,N_9250);
and U10838 (N_10838,N_9242,N_9686);
and U10839 (N_10839,N_9765,N_9486);
xor U10840 (N_10840,N_9412,N_9178);
nand U10841 (N_10841,N_9207,N_9058);
or U10842 (N_10842,N_9520,N_9386);
nor U10843 (N_10843,N_9090,N_9775);
and U10844 (N_10844,N_9772,N_9883);
and U10845 (N_10845,N_9614,N_9338);
and U10846 (N_10846,N_9483,N_9531);
or U10847 (N_10847,N_9100,N_9460);
and U10848 (N_10848,N_9058,N_9203);
or U10849 (N_10849,N_9711,N_9845);
xor U10850 (N_10850,N_9286,N_9021);
nand U10851 (N_10851,N_9637,N_9130);
nand U10852 (N_10852,N_9693,N_9134);
or U10853 (N_10853,N_9877,N_9884);
xor U10854 (N_10854,N_9927,N_9976);
nor U10855 (N_10855,N_9458,N_9534);
nand U10856 (N_10856,N_9338,N_9804);
nor U10857 (N_10857,N_9150,N_9611);
or U10858 (N_10858,N_9102,N_9051);
and U10859 (N_10859,N_9166,N_9868);
or U10860 (N_10860,N_9599,N_9654);
and U10861 (N_10861,N_9738,N_9069);
nand U10862 (N_10862,N_9204,N_9580);
nand U10863 (N_10863,N_9255,N_9330);
nor U10864 (N_10864,N_9371,N_9578);
or U10865 (N_10865,N_9702,N_9123);
xnor U10866 (N_10866,N_9977,N_9199);
xor U10867 (N_10867,N_9749,N_9338);
xor U10868 (N_10868,N_9372,N_9135);
nand U10869 (N_10869,N_9380,N_9325);
and U10870 (N_10870,N_9991,N_9861);
and U10871 (N_10871,N_9213,N_9224);
or U10872 (N_10872,N_9642,N_9613);
xor U10873 (N_10873,N_9106,N_9400);
nand U10874 (N_10874,N_9867,N_9159);
nor U10875 (N_10875,N_9659,N_9031);
xnor U10876 (N_10876,N_9194,N_9988);
xnor U10877 (N_10877,N_9066,N_9272);
or U10878 (N_10878,N_9664,N_9835);
or U10879 (N_10879,N_9602,N_9399);
xor U10880 (N_10880,N_9596,N_9072);
and U10881 (N_10881,N_9663,N_9302);
xnor U10882 (N_10882,N_9952,N_9244);
nor U10883 (N_10883,N_9981,N_9261);
or U10884 (N_10884,N_9026,N_9343);
nor U10885 (N_10885,N_9936,N_9819);
nand U10886 (N_10886,N_9513,N_9372);
xnor U10887 (N_10887,N_9787,N_9891);
or U10888 (N_10888,N_9397,N_9439);
or U10889 (N_10889,N_9471,N_9937);
nor U10890 (N_10890,N_9189,N_9645);
or U10891 (N_10891,N_9880,N_9795);
or U10892 (N_10892,N_9441,N_9995);
xnor U10893 (N_10893,N_9569,N_9122);
nand U10894 (N_10894,N_9249,N_9691);
nand U10895 (N_10895,N_9708,N_9763);
nand U10896 (N_10896,N_9590,N_9080);
or U10897 (N_10897,N_9241,N_9611);
nand U10898 (N_10898,N_9384,N_9789);
nor U10899 (N_10899,N_9887,N_9335);
and U10900 (N_10900,N_9442,N_9516);
xor U10901 (N_10901,N_9231,N_9786);
and U10902 (N_10902,N_9145,N_9836);
xnor U10903 (N_10903,N_9244,N_9727);
nand U10904 (N_10904,N_9577,N_9481);
nor U10905 (N_10905,N_9796,N_9261);
xnor U10906 (N_10906,N_9971,N_9463);
xor U10907 (N_10907,N_9402,N_9767);
nor U10908 (N_10908,N_9039,N_9027);
xor U10909 (N_10909,N_9775,N_9957);
xor U10910 (N_10910,N_9766,N_9367);
nand U10911 (N_10911,N_9459,N_9807);
nand U10912 (N_10912,N_9742,N_9618);
nand U10913 (N_10913,N_9138,N_9707);
nand U10914 (N_10914,N_9417,N_9717);
nand U10915 (N_10915,N_9545,N_9542);
or U10916 (N_10916,N_9230,N_9433);
nor U10917 (N_10917,N_9014,N_9201);
or U10918 (N_10918,N_9591,N_9304);
nor U10919 (N_10919,N_9837,N_9070);
or U10920 (N_10920,N_9941,N_9730);
or U10921 (N_10921,N_9548,N_9610);
or U10922 (N_10922,N_9423,N_9316);
and U10923 (N_10923,N_9261,N_9158);
xor U10924 (N_10924,N_9502,N_9909);
nand U10925 (N_10925,N_9488,N_9190);
xor U10926 (N_10926,N_9980,N_9302);
and U10927 (N_10927,N_9408,N_9897);
xnor U10928 (N_10928,N_9381,N_9011);
xnor U10929 (N_10929,N_9388,N_9686);
and U10930 (N_10930,N_9880,N_9977);
or U10931 (N_10931,N_9449,N_9886);
nand U10932 (N_10932,N_9557,N_9055);
and U10933 (N_10933,N_9431,N_9573);
and U10934 (N_10934,N_9129,N_9411);
and U10935 (N_10935,N_9830,N_9848);
or U10936 (N_10936,N_9495,N_9746);
or U10937 (N_10937,N_9374,N_9858);
nand U10938 (N_10938,N_9526,N_9669);
nor U10939 (N_10939,N_9065,N_9455);
nand U10940 (N_10940,N_9660,N_9006);
or U10941 (N_10941,N_9162,N_9015);
xor U10942 (N_10942,N_9746,N_9992);
xnor U10943 (N_10943,N_9442,N_9934);
nand U10944 (N_10944,N_9847,N_9959);
xor U10945 (N_10945,N_9342,N_9308);
nor U10946 (N_10946,N_9678,N_9118);
or U10947 (N_10947,N_9516,N_9147);
nor U10948 (N_10948,N_9854,N_9842);
and U10949 (N_10949,N_9150,N_9994);
nand U10950 (N_10950,N_9964,N_9752);
nor U10951 (N_10951,N_9373,N_9477);
and U10952 (N_10952,N_9326,N_9559);
and U10953 (N_10953,N_9907,N_9287);
and U10954 (N_10954,N_9233,N_9152);
and U10955 (N_10955,N_9023,N_9396);
nand U10956 (N_10956,N_9224,N_9935);
nand U10957 (N_10957,N_9900,N_9395);
nor U10958 (N_10958,N_9428,N_9061);
xnor U10959 (N_10959,N_9010,N_9873);
and U10960 (N_10960,N_9376,N_9736);
nand U10961 (N_10961,N_9806,N_9230);
nand U10962 (N_10962,N_9904,N_9155);
and U10963 (N_10963,N_9544,N_9859);
or U10964 (N_10964,N_9921,N_9749);
and U10965 (N_10965,N_9025,N_9121);
nand U10966 (N_10966,N_9804,N_9794);
nor U10967 (N_10967,N_9200,N_9859);
xor U10968 (N_10968,N_9817,N_9554);
and U10969 (N_10969,N_9706,N_9806);
or U10970 (N_10970,N_9730,N_9179);
nor U10971 (N_10971,N_9879,N_9984);
nor U10972 (N_10972,N_9975,N_9925);
xor U10973 (N_10973,N_9276,N_9416);
nor U10974 (N_10974,N_9969,N_9622);
nor U10975 (N_10975,N_9531,N_9830);
nor U10976 (N_10976,N_9683,N_9520);
xnor U10977 (N_10977,N_9824,N_9934);
nor U10978 (N_10978,N_9637,N_9499);
and U10979 (N_10979,N_9865,N_9048);
and U10980 (N_10980,N_9288,N_9511);
nor U10981 (N_10981,N_9930,N_9910);
nand U10982 (N_10982,N_9635,N_9396);
and U10983 (N_10983,N_9859,N_9027);
nand U10984 (N_10984,N_9140,N_9595);
nor U10985 (N_10985,N_9021,N_9880);
nor U10986 (N_10986,N_9623,N_9277);
and U10987 (N_10987,N_9250,N_9467);
xnor U10988 (N_10988,N_9194,N_9548);
or U10989 (N_10989,N_9116,N_9287);
or U10990 (N_10990,N_9198,N_9906);
nor U10991 (N_10991,N_9303,N_9500);
nand U10992 (N_10992,N_9683,N_9606);
nand U10993 (N_10993,N_9622,N_9284);
nand U10994 (N_10994,N_9851,N_9761);
nand U10995 (N_10995,N_9652,N_9214);
xnor U10996 (N_10996,N_9017,N_9244);
and U10997 (N_10997,N_9925,N_9645);
xnor U10998 (N_10998,N_9604,N_9987);
or U10999 (N_10999,N_9695,N_9965);
nor U11000 (N_11000,N_10686,N_10161);
or U11001 (N_11001,N_10751,N_10454);
nand U11002 (N_11002,N_10027,N_10959);
nor U11003 (N_11003,N_10905,N_10312);
xnor U11004 (N_11004,N_10259,N_10449);
or U11005 (N_11005,N_10094,N_10292);
nor U11006 (N_11006,N_10574,N_10783);
nand U11007 (N_11007,N_10323,N_10355);
nand U11008 (N_11008,N_10950,N_10277);
nor U11009 (N_11009,N_10412,N_10171);
xnor U11010 (N_11010,N_10251,N_10321);
xnor U11011 (N_11011,N_10472,N_10169);
xnor U11012 (N_11012,N_10765,N_10213);
and U11013 (N_11013,N_10249,N_10502);
nor U11014 (N_11014,N_10416,N_10481);
nor U11015 (N_11015,N_10828,N_10096);
or U11016 (N_11016,N_10946,N_10392);
xnor U11017 (N_11017,N_10922,N_10128);
or U11018 (N_11018,N_10967,N_10314);
xor U11019 (N_11019,N_10555,N_10699);
nor U11020 (N_11020,N_10630,N_10237);
or U11021 (N_11021,N_10855,N_10977);
and U11022 (N_11022,N_10224,N_10667);
xor U11023 (N_11023,N_10427,N_10365);
xnor U11024 (N_11024,N_10152,N_10095);
or U11025 (N_11025,N_10285,N_10430);
nor U11026 (N_11026,N_10076,N_10371);
or U11027 (N_11027,N_10401,N_10448);
or U11028 (N_11028,N_10850,N_10810);
nand U11029 (N_11029,N_10269,N_10694);
xnor U11030 (N_11030,N_10796,N_10549);
xnor U11031 (N_11031,N_10640,N_10522);
nand U11032 (N_11032,N_10623,N_10725);
nor U11033 (N_11033,N_10331,N_10439);
or U11034 (N_11034,N_10511,N_10866);
and U11035 (N_11035,N_10088,N_10507);
nand U11036 (N_11036,N_10784,N_10927);
nand U11037 (N_11037,N_10330,N_10366);
xor U11038 (N_11038,N_10650,N_10772);
xnor U11039 (N_11039,N_10433,N_10553);
xnor U11040 (N_11040,N_10638,N_10230);
and U11041 (N_11041,N_10232,N_10024);
nand U11042 (N_11042,N_10973,N_10681);
nor U11043 (N_11043,N_10202,N_10917);
or U11044 (N_11044,N_10865,N_10939);
nor U11045 (N_11045,N_10443,N_10659);
and U11046 (N_11046,N_10656,N_10087);
xnor U11047 (N_11047,N_10792,N_10918);
nor U11048 (N_11048,N_10505,N_10933);
nand U11049 (N_11049,N_10453,N_10451);
xor U11050 (N_11050,N_10531,N_10113);
nor U11051 (N_11051,N_10352,N_10697);
xnor U11052 (N_11052,N_10123,N_10708);
and U11053 (N_11053,N_10423,N_10390);
or U11054 (N_11054,N_10016,N_10499);
xnor U11055 (N_11055,N_10740,N_10308);
xnor U11056 (N_11056,N_10821,N_10122);
nand U11057 (N_11057,N_10081,N_10090);
and U11058 (N_11058,N_10182,N_10856);
and U11059 (N_11059,N_10183,N_10537);
nor U11060 (N_11060,N_10389,N_10737);
or U11061 (N_11061,N_10750,N_10085);
and U11062 (N_11062,N_10009,N_10884);
xnor U11063 (N_11063,N_10260,N_10711);
or U11064 (N_11064,N_10653,N_10347);
or U11065 (N_11065,N_10872,N_10188);
nand U11066 (N_11066,N_10108,N_10763);
nor U11067 (N_11067,N_10860,N_10280);
nor U11068 (N_11068,N_10376,N_10851);
and U11069 (N_11069,N_10688,N_10603);
xor U11070 (N_11070,N_10215,N_10078);
or U11071 (N_11071,N_10031,N_10503);
nand U11072 (N_11072,N_10227,N_10310);
nand U11073 (N_11073,N_10972,N_10039);
nand U11074 (N_11074,N_10834,N_10521);
xnor U11075 (N_11075,N_10781,N_10332);
xnor U11076 (N_11076,N_10391,N_10173);
or U11077 (N_11077,N_10168,N_10929);
xor U11078 (N_11078,N_10944,N_10646);
nor U11079 (N_11079,N_10621,N_10988);
nand U11080 (N_11080,N_10995,N_10999);
or U11081 (N_11081,N_10844,N_10106);
or U11082 (N_11082,N_10518,N_10836);
or U11083 (N_11083,N_10490,N_10265);
nand U11084 (N_11084,N_10703,N_10261);
xor U11085 (N_11085,N_10738,N_10165);
nand U11086 (N_11086,N_10786,N_10317);
xnor U11087 (N_11087,N_10466,N_10824);
nor U11088 (N_11088,N_10220,N_10222);
or U11089 (N_11089,N_10561,N_10931);
nor U11090 (N_11090,N_10357,N_10368);
or U11091 (N_11091,N_10002,N_10342);
nand U11092 (N_11092,N_10256,N_10761);
nand U11093 (N_11093,N_10373,N_10397);
nor U11094 (N_11094,N_10780,N_10969);
and U11095 (N_11095,N_10057,N_10691);
xnor U11096 (N_11096,N_10870,N_10877);
xnor U11097 (N_11097,N_10146,N_10890);
xor U11098 (N_11098,N_10483,N_10971);
xnor U11099 (N_11099,N_10255,N_10897);
xnor U11100 (N_11100,N_10825,N_10904);
nor U11101 (N_11101,N_10558,N_10712);
and U11102 (N_11102,N_10046,N_10941);
or U11103 (N_11103,N_10579,N_10315);
or U11104 (N_11104,N_10385,N_10990);
xnor U11105 (N_11105,N_10976,N_10678);
nor U11106 (N_11106,N_10666,N_10673);
nor U11107 (N_11107,N_10982,N_10636);
nor U11108 (N_11108,N_10428,N_10798);
nand U11109 (N_11109,N_10609,N_10879);
nor U11110 (N_11110,N_10114,N_10829);
and U11111 (N_11111,N_10911,N_10670);
xor U11112 (N_11112,N_10231,N_10745);
nand U11113 (N_11113,N_10706,N_10271);
or U11114 (N_11114,N_10162,N_10773);
and U11115 (N_11115,N_10077,N_10595);
or U11116 (N_11116,N_10845,N_10369);
or U11117 (N_11117,N_10891,N_10937);
nor U11118 (N_11118,N_10318,N_10302);
nand U11119 (N_11119,N_10372,N_10004);
nor U11120 (N_11120,N_10075,N_10446);
or U11121 (N_11121,N_10926,N_10934);
xor U11122 (N_11122,N_10042,N_10746);
and U11123 (N_11123,N_10203,N_10334);
xnor U11124 (N_11124,N_10730,N_10327);
nand U11125 (N_11125,N_10665,N_10105);
or U11126 (N_11126,N_10777,N_10395);
and U11127 (N_11127,N_10386,N_10525);
or U11128 (N_11128,N_10023,N_10361);
nand U11129 (N_11129,N_10047,N_10238);
nand U11130 (N_11130,N_10402,N_10497);
or U11131 (N_11131,N_10135,N_10298);
and U11132 (N_11132,N_10727,N_10808);
nor U11133 (N_11133,N_10104,N_10282);
xor U11134 (N_11134,N_10894,N_10160);
or U11135 (N_11135,N_10262,N_10247);
nor U11136 (N_11136,N_10229,N_10089);
xnor U11137 (N_11137,N_10025,N_10830);
and U11138 (N_11138,N_10593,N_10818);
nand U11139 (N_11139,N_10017,N_10809);
nand U11140 (N_11140,N_10696,N_10311);
xnor U11141 (N_11141,N_10217,N_10572);
nand U11142 (N_11142,N_10354,N_10543);
nand U11143 (N_11143,N_10793,N_10072);
or U11144 (N_11144,N_10148,N_10337);
nand U11145 (N_11145,N_10540,N_10677);
nor U11146 (N_11146,N_10283,N_10137);
or U11147 (N_11147,N_10329,N_10859);
or U11148 (N_11148,N_10952,N_10120);
nor U11149 (N_11149,N_10007,N_10649);
nor U11150 (N_11150,N_10582,N_10043);
nor U11151 (N_11151,N_10820,N_10356);
xnor U11152 (N_11152,N_10468,N_10698);
xor U11153 (N_11153,N_10536,N_10167);
nand U11154 (N_11154,N_10841,N_10550);
nand U11155 (N_11155,N_10274,N_10441);
and U11156 (N_11156,N_10320,N_10436);
nor U11157 (N_11157,N_10486,N_10571);
nand U11158 (N_11158,N_10112,N_10534);
or U11159 (N_11159,N_10058,N_10524);
nand U11160 (N_11160,N_10339,N_10151);
or U11161 (N_11161,N_10467,N_10252);
nor U11162 (N_11162,N_10364,N_10930);
and U11163 (N_11163,N_10049,N_10626);
and U11164 (N_11164,N_10111,N_10200);
nor U11165 (N_11165,N_10858,N_10407);
xnor U11166 (N_11166,N_10597,N_10544);
or U11167 (N_11167,N_10133,N_10216);
and U11168 (N_11168,N_10605,N_10063);
or U11169 (N_11169,N_10770,N_10463);
or U11170 (N_11170,N_10294,N_10790);
xnor U11171 (N_11171,N_10878,N_10797);
xor U11172 (N_11172,N_10760,N_10629);
and U11173 (N_11173,N_10241,N_10375);
or U11174 (N_11174,N_10726,N_10799);
xnor U11175 (N_11175,N_10715,N_10492);
xor U11176 (N_11176,N_10559,N_10618);
or U11177 (N_11177,N_10353,N_10705);
nand U11178 (N_11178,N_10403,N_10343);
and U11179 (N_11179,N_10288,N_10289);
nor U11180 (N_11180,N_10800,N_10811);
or U11181 (N_11181,N_10854,N_10936);
and U11182 (N_11182,N_10663,N_10557);
and U11183 (N_11183,N_10145,N_10538);
and U11184 (N_11184,N_10056,N_10303);
nand U11185 (N_11185,N_10370,N_10156);
nand U11186 (N_11186,N_10583,N_10073);
and U11187 (N_11187,N_10869,N_10138);
or U11188 (N_11188,N_10379,N_10533);
and U11189 (N_11189,N_10005,N_10189);
or U11190 (N_11190,N_10886,N_10669);
nor U11191 (N_11191,N_10101,N_10489);
and U11192 (N_11192,N_10822,N_10498);
and U11193 (N_11193,N_10209,N_10421);
nand U11194 (N_11194,N_10129,N_10126);
nor U11195 (N_11195,N_10325,N_10187);
xor U11196 (N_11196,N_10565,N_10932);
nand U11197 (N_11197,N_10040,N_10580);
xnor U11198 (N_11198,N_10476,N_10617);
nor U11199 (N_11199,N_10083,N_10912);
or U11200 (N_11200,N_10170,N_10814);
nor U11201 (N_11201,N_10720,N_10608);
nand U11202 (N_11202,N_10889,N_10921);
and U11203 (N_11203,N_10632,N_10000);
nand U11204 (N_11204,N_10084,N_10431);
nand U11205 (N_11205,N_10465,N_10450);
nand U11206 (N_11206,N_10457,N_10097);
and U11207 (N_11207,N_10299,N_10198);
nor U11208 (N_11208,N_10517,N_10835);
and U11209 (N_11209,N_10975,N_10414);
or U11210 (N_11210,N_10634,N_10838);
or U11211 (N_11211,N_10943,N_10333);
nand U11212 (N_11212,N_10248,N_10053);
xor U11213 (N_11213,N_10034,N_10791);
xor U11214 (N_11214,N_10140,N_10909);
and U11215 (N_11215,N_10473,N_10803);
or U11216 (N_11216,N_10281,N_10991);
nor U11217 (N_11217,N_10279,N_10885);
or U11218 (N_11218,N_10242,N_10736);
or U11219 (N_11219,N_10071,N_10254);
xnor U11220 (N_11220,N_10601,N_10585);
nor U11221 (N_11221,N_10127,N_10445);
and U11222 (N_11222,N_10819,N_10309);
nand U11223 (N_11223,N_10052,N_10551);
nand U11224 (N_11224,N_10876,N_10197);
nand U11225 (N_11225,N_10506,N_10576);
xor U11226 (N_11226,N_10328,N_10606);
and U11227 (N_11227,N_10484,N_10050);
nor U11228 (N_11228,N_10635,N_10253);
xor U11229 (N_11229,N_10074,N_10477);
nor U11230 (N_11230,N_10616,N_10861);
nor U11231 (N_11231,N_10258,N_10619);
and U11232 (N_11232,N_10532,N_10970);
nor U11233 (N_11233,N_10948,N_10704);
nor U11234 (N_11234,N_10748,N_10631);
and U11235 (N_11235,N_10048,N_10304);
xnor U11236 (N_11236,N_10776,N_10037);
xnor U11237 (N_11237,N_10622,N_10755);
xor U11238 (N_11238,N_10575,N_10853);
xor U11239 (N_11239,N_10464,N_10657);
and U11240 (N_11240,N_10324,N_10979);
nor U11241 (N_11241,N_10022,N_10707);
and U11242 (N_11242,N_10724,N_10749);
or U11243 (N_11243,N_10660,N_10150);
and U11244 (N_11244,N_10459,N_10722);
xor U11245 (N_11245,N_10219,N_10272);
nor U11246 (N_11246,N_10296,N_10510);
nor U11247 (N_11247,N_10384,N_10983);
or U11248 (N_11248,N_10257,N_10569);
and U11249 (N_11249,N_10006,N_10419);
nand U11250 (N_11250,N_10080,N_10482);
nand U11251 (N_11251,N_10341,N_10003);
and U11252 (N_11252,N_10462,N_10475);
and U11253 (N_11253,N_10455,N_10587);
and U11254 (N_11254,N_10951,N_10030);
xor U11255 (N_11255,N_10900,N_10035);
nand U11256 (N_11256,N_10306,N_10994);
or U11257 (N_11257,N_10898,N_10149);
and U11258 (N_11258,N_10675,N_10029);
xor U11259 (N_11259,N_10644,N_10286);
nor U11260 (N_11260,N_10680,N_10935);
nor U11261 (N_11261,N_10420,N_10195);
nand U11262 (N_11262,N_10692,N_10599);
xnor U11263 (N_11263,N_10846,N_10903);
nand U11264 (N_11264,N_10815,N_10297);
nor U11265 (N_11265,N_10588,N_10516);
nor U11266 (N_11266,N_10539,N_10514);
nand U11267 (N_11267,N_10409,N_10584);
nor U11268 (N_11268,N_10611,N_10562);
nand U11269 (N_11269,N_10914,N_10968);
or U11270 (N_11270,N_10501,N_10461);
and U11271 (N_11271,N_10958,N_10774);
and U11272 (N_11272,N_10275,N_10250);
nor U11273 (N_11273,N_10847,N_10782);
nand U11274 (N_11274,N_10739,N_10945);
or U11275 (N_11275,N_10100,N_10179);
nor U11276 (N_11276,N_10731,N_10924);
nand U11277 (N_11277,N_10523,N_10652);
nor U11278 (N_11278,N_10741,N_10319);
xnor U11279 (N_11279,N_10639,N_10415);
nand U11280 (N_11280,N_10118,N_10488);
and U11281 (N_11281,N_10529,N_10018);
nand U11282 (N_11282,N_10066,N_10805);
xnor U11283 (N_11283,N_10228,N_10381);
xor U11284 (N_11284,N_10452,N_10664);
nand U11285 (N_11285,N_10615,N_10789);
nand U11286 (N_11286,N_10567,N_10210);
and U11287 (N_11287,N_10961,N_10028);
nand U11288 (N_11288,N_10642,N_10020);
or U11289 (N_11289,N_10326,N_10713);
nand U11290 (N_11290,N_10719,N_10019);
nor U11291 (N_11291,N_10848,N_10244);
nor U11292 (N_11292,N_10172,N_10413);
and U11293 (N_11293,N_10117,N_10671);
and U11294 (N_11294,N_10987,N_10676);
and U11295 (N_11295,N_10940,N_10766);
nor U11296 (N_11296,N_10079,N_10693);
nor U11297 (N_11297,N_10193,N_10344);
nand U11298 (N_11298,N_10164,N_10012);
or U11299 (N_11299,N_10554,N_10794);
or U11300 (N_11300,N_10065,N_10602);
and U11301 (N_11301,N_10956,N_10440);
or U11302 (N_11302,N_10163,N_10823);
xnor U11303 (N_11303,N_10542,N_10775);
nand U11304 (N_11304,N_10610,N_10054);
nand U11305 (N_11305,N_10873,N_10273);
xor U11306 (N_11306,N_10573,N_10062);
xor U11307 (N_11307,N_10175,N_10181);
nor U11308 (N_11308,N_10996,N_10812);
xnor U11309 (N_11309,N_10925,N_10570);
or U11310 (N_11310,N_10221,N_10989);
nand U11311 (N_11311,N_10068,N_10684);
nor U11312 (N_11312,N_10378,N_10960);
or U11313 (N_11313,N_10234,N_10059);
xor U11314 (N_11314,N_10702,N_10211);
nor U11315 (N_11315,N_10756,N_10155);
xnor U11316 (N_11316,N_10778,N_10284);
and U11317 (N_11317,N_10493,N_10655);
xor U11318 (N_11318,N_10432,N_10633);
nor U11319 (N_11319,N_10986,N_10208);
or U11320 (N_11320,N_10394,N_10266);
nor U11321 (N_11321,N_10586,N_10612);
nand U11322 (N_11322,N_10293,N_10103);
nand U11323 (N_11323,N_10426,N_10758);
xor U11324 (N_11324,N_10001,N_10067);
and U11325 (N_11325,N_10604,N_10546);
nand U11326 (N_11326,N_10144,N_10863);
nor U11327 (N_11327,N_10226,N_10654);
or U11328 (N_11328,N_10192,N_10185);
or U11329 (N_11329,N_10893,N_10743);
and U11330 (N_11330,N_10700,N_10607);
nand U11331 (N_11331,N_10816,N_10628);
nand U11332 (N_11332,N_10833,N_10316);
and U11333 (N_11333,N_10041,N_10881);
xor U11334 (N_11334,N_10624,N_10469);
or U11335 (N_11335,N_10504,N_10136);
xor U11336 (N_11336,N_10913,N_10398);
xor U11337 (N_11337,N_10674,N_10668);
nand U11338 (N_11338,N_10458,N_10560);
or U11339 (N_11339,N_10070,N_10487);
nand U11340 (N_11340,N_10752,N_10620);
nor U11341 (N_11341,N_10839,N_10648);
nor U11342 (N_11342,N_10011,N_10055);
and U11343 (N_11343,N_10245,N_10278);
and U11344 (N_11344,N_10207,N_10957);
xnor U11345 (N_11345,N_10268,N_10928);
xor U11346 (N_11346,N_10240,N_10125);
and U11347 (N_11347,N_10036,N_10683);
xor U11348 (N_11348,N_10910,N_10474);
xnor U11349 (N_11349,N_10092,N_10199);
nand U11350 (N_11350,N_10290,N_10444);
or U11351 (N_11351,N_10134,N_10747);
or U11352 (N_11352,N_10981,N_10902);
nand U11353 (N_11353,N_10919,N_10166);
nor U11354 (N_11354,N_10807,N_10093);
or U11355 (N_11355,N_10153,N_10535);
xnor U11356 (N_11356,N_10955,N_10500);
or U11357 (N_11357,N_10154,N_10887);
or U11358 (N_11358,N_10788,N_10382);
nor U11359 (N_11359,N_10225,N_10592);
or U11360 (N_11360,N_10978,N_10346);
nand U11361 (N_11361,N_10119,N_10520);
and U11362 (N_11362,N_10641,N_10026);
or U11363 (N_11363,N_10374,N_10060);
nand U11364 (N_11364,N_10132,N_10235);
and U11365 (N_11365,N_10843,N_10116);
and U11366 (N_11366,N_10051,N_10980);
and U11367 (N_11367,N_10985,N_10710);
nor U11368 (N_11368,N_10578,N_10141);
or U11369 (N_11369,N_10061,N_10380);
and U11370 (N_11370,N_10107,N_10239);
and U11371 (N_11371,N_10735,N_10264);
nor U11372 (N_11372,N_10625,N_10840);
and U11373 (N_11373,N_10435,N_10864);
nor U11374 (N_11374,N_10753,N_10637);
or U11375 (N_11375,N_10340,N_10779);
nand U11376 (N_11376,N_10813,N_10831);
nand U11377 (N_11377,N_10837,N_10658);
or U11378 (N_11378,N_10404,N_10672);
nand U11379 (N_11379,N_10447,N_10733);
nand U11380 (N_11380,N_10530,N_10301);
nor U11381 (N_11381,N_10548,N_10920);
or U11382 (N_11382,N_10515,N_10563);
and U11383 (N_11383,N_10509,N_10045);
and U11384 (N_11384,N_10410,N_10716);
xnor U11385 (N_11385,N_10405,N_10687);
or U11386 (N_11386,N_10177,N_10362);
xor U11387 (N_11387,N_10868,N_10589);
nand U11388 (N_11388,N_10098,N_10964);
and U11389 (N_11389,N_10817,N_10754);
nand U11390 (N_11390,N_10614,N_10010);
nor U11391 (N_11391,N_10896,N_10787);
xor U11392 (N_11392,N_10335,N_10471);
nor U11393 (N_11393,N_10295,N_10246);
and U11394 (N_11394,N_10723,N_10947);
or U11395 (N_11395,N_10709,N_10827);
nand U11396 (N_11396,N_10021,N_10400);
or U11397 (N_11397,N_10243,N_10867);
xnor U11398 (N_11398,N_10801,N_10849);
nand U11399 (N_11399,N_10233,N_10842);
nor U11400 (N_11400,N_10008,N_10032);
or U11401 (N_11401,N_10857,N_10962);
nor U11402 (N_11402,N_10434,N_10963);
and U11403 (N_11403,N_10157,N_10287);
or U11404 (N_11404,N_10349,N_10742);
nand U11405 (N_11405,N_10178,N_10204);
nand U11406 (N_11406,N_10862,N_10044);
xor U11407 (N_11407,N_10442,N_10527);
nor U11408 (N_11408,N_10966,N_10767);
nor U11409 (N_11409,N_10528,N_10802);
xnor U11410 (N_11410,N_10734,N_10594);
or U11411 (N_11411,N_10267,N_10908);
and U11412 (N_11412,N_10313,N_10184);
nor U11413 (N_11413,N_10015,N_10429);
and U11414 (N_11414,N_10645,N_10759);
nor U11415 (N_11415,N_10883,N_10345);
xor U11416 (N_11416,N_10744,N_10764);
xor U11417 (N_11417,N_10115,N_10984);
nor U11418 (N_11418,N_10437,N_10880);
xor U11419 (N_11419,N_10411,N_10965);
and U11420 (N_11420,N_10142,N_10300);
nor U11421 (N_11421,N_10033,N_10769);
and U11422 (N_11422,N_10064,N_10383);
xor U11423 (N_11423,N_10013,N_10091);
nand U11424 (N_11424,N_10263,N_10218);
nor U11425 (N_11425,N_10307,N_10591);
nor U11426 (N_11426,N_10627,N_10494);
and U11427 (N_11427,N_10552,N_10069);
and U11428 (N_11428,N_10363,N_10360);
and U11429 (N_11429,N_10491,N_10086);
and U11430 (N_11430,N_10212,N_10690);
xor U11431 (N_11431,N_10901,N_10875);
or U11432 (N_11432,N_10393,N_10131);
or U11433 (N_11433,N_10270,N_10682);
xnor U11434 (N_11434,N_10895,N_10495);
or U11435 (N_11435,N_10547,N_10613);
xnor U11436 (N_11436,N_10806,N_10186);
xor U11437 (N_11437,N_10038,N_10470);
xnor U11438 (N_11438,N_10479,N_10406);
xnor U11439 (N_11439,N_10997,N_10662);
nor U11440 (N_11440,N_10729,N_10350);
nor U11441 (N_11441,N_10721,N_10305);
or U11442 (N_11442,N_10367,N_10771);
or U11443 (N_11443,N_10992,N_10916);
xor U11444 (N_11444,N_10892,N_10942);
or U11445 (N_11445,N_10581,N_10418);
nand U11446 (N_11446,N_10201,N_10695);
or U11447 (N_11447,N_10110,N_10545);
or U11448 (N_11448,N_10564,N_10882);
or U11449 (N_11449,N_10899,N_10496);
and U11450 (N_11450,N_10647,N_10577);
and U11451 (N_11451,N_10102,N_10590);
nand U11452 (N_11452,N_10762,N_10661);
or U11453 (N_11453,N_10456,N_10679);
or U11454 (N_11454,N_10714,N_10954);
and U11455 (N_11455,N_10396,N_10974);
or U11456 (N_11456,N_10358,N_10014);
nand U11457 (N_11457,N_10147,N_10214);
nand U11458 (N_11458,N_10139,N_10526);
xnor U11459 (N_11459,N_10351,N_10852);
nor U11460 (N_11460,N_10832,N_10176);
and U11461 (N_11461,N_10399,N_10508);
nor U11462 (N_11462,N_10408,N_10417);
nand U11463 (N_11463,N_10438,N_10568);
or U11464 (N_11464,N_10387,N_10651);
nand U11465 (N_11465,N_10124,N_10512);
and U11466 (N_11466,N_10159,N_10757);
xnor U11467 (N_11467,N_10206,N_10938);
and U11468 (N_11468,N_10099,N_10596);
and U11469 (N_11469,N_10888,N_10717);
or U11470 (N_11470,N_10205,N_10194);
nor U11471 (N_11471,N_10953,N_10190);
nand U11472 (N_11472,N_10480,N_10513);
nor U11473 (N_11473,N_10998,N_10424);
xnor U11474 (N_11474,N_10804,N_10130);
nor U11475 (N_11475,N_10768,N_10348);
xor U11476 (N_11476,N_10795,N_10422);
or U11477 (N_11477,N_10600,N_10425);
or U11478 (N_11478,N_10915,N_10377);
nand U11479 (N_11479,N_10728,N_10907);
and U11480 (N_11480,N_10718,N_10541);
xnor U11481 (N_11481,N_10732,N_10121);
or U11482 (N_11482,N_10291,N_10874);
or U11483 (N_11483,N_10336,N_10460);
xor U11484 (N_11484,N_10485,N_10993);
nand U11485 (N_11485,N_10519,N_10826);
xor U11486 (N_11486,N_10598,N_10388);
nor U11487 (N_11487,N_10643,N_10180);
nor U11488 (N_11488,N_10685,N_10871);
and U11489 (N_11489,N_10906,N_10338);
and U11490 (N_11490,N_10082,N_10109);
and U11491 (N_11491,N_10785,N_10158);
and U11492 (N_11492,N_10949,N_10322);
nor U11493 (N_11493,N_10359,N_10143);
xor U11494 (N_11494,N_10478,N_10689);
nand U11495 (N_11495,N_10701,N_10223);
nand U11496 (N_11496,N_10923,N_10236);
nand U11497 (N_11497,N_10276,N_10196);
and U11498 (N_11498,N_10191,N_10174);
nor U11499 (N_11499,N_10566,N_10556);
nand U11500 (N_11500,N_10783,N_10073);
nor U11501 (N_11501,N_10279,N_10847);
or U11502 (N_11502,N_10899,N_10584);
nor U11503 (N_11503,N_10573,N_10428);
nand U11504 (N_11504,N_10852,N_10977);
xnor U11505 (N_11505,N_10199,N_10322);
xnor U11506 (N_11506,N_10331,N_10907);
and U11507 (N_11507,N_10723,N_10280);
nand U11508 (N_11508,N_10555,N_10218);
nand U11509 (N_11509,N_10916,N_10763);
and U11510 (N_11510,N_10066,N_10576);
xnor U11511 (N_11511,N_10459,N_10392);
and U11512 (N_11512,N_10959,N_10262);
nand U11513 (N_11513,N_10820,N_10193);
and U11514 (N_11514,N_10203,N_10683);
and U11515 (N_11515,N_10852,N_10243);
nand U11516 (N_11516,N_10302,N_10232);
nand U11517 (N_11517,N_10481,N_10151);
nand U11518 (N_11518,N_10247,N_10588);
or U11519 (N_11519,N_10817,N_10039);
nand U11520 (N_11520,N_10296,N_10546);
nor U11521 (N_11521,N_10062,N_10463);
xor U11522 (N_11522,N_10549,N_10325);
nand U11523 (N_11523,N_10302,N_10354);
or U11524 (N_11524,N_10298,N_10678);
xnor U11525 (N_11525,N_10216,N_10252);
and U11526 (N_11526,N_10112,N_10269);
nor U11527 (N_11527,N_10572,N_10949);
or U11528 (N_11528,N_10132,N_10642);
nand U11529 (N_11529,N_10107,N_10324);
xor U11530 (N_11530,N_10004,N_10007);
and U11531 (N_11531,N_10679,N_10516);
or U11532 (N_11532,N_10946,N_10748);
nand U11533 (N_11533,N_10973,N_10974);
and U11534 (N_11534,N_10033,N_10558);
nand U11535 (N_11535,N_10489,N_10743);
xnor U11536 (N_11536,N_10213,N_10824);
nand U11537 (N_11537,N_10008,N_10685);
and U11538 (N_11538,N_10972,N_10806);
nand U11539 (N_11539,N_10730,N_10624);
xnor U11540 (N_11540,N_10458,N_10478);
nor U11541 (N_11541,N_10522,N_10491);
or U11542 (N_11542,N_10320,N_10164);
or U11543 (N_11543,N_10575,N_10049);
xnor U11544 (N_11544,N_10080,N_10906);
nor U11545 (N_11545,N_10155,N_10119);
and U11546 (N_11546,N_10637,N_10845);
or U11547 (N_11547,N_10687,N_10256);
nor U11548 (N_11548,N_10340,N_10567);
nor U11549 (N_11549,N_10114,N_10519);
nor U11550 (N_11550,N_10966,N_10296);
and U11551 (N_11551,N_10423,N_10714);
nor U11552 (N_11552,N_10812,N_10751);
or U11553 (N_11553,N_10242,N_10376);
or U11554 (N_11554,N_10968,N_10829);
and U11555 (N_11555,N_10081,N_10684);
and U11556 (N_11556,N_10161,N_10677);
xor U11557 (N_11557,N_10455,N_10766);
nand U11558 (N_11558,N_10257,N_10901);
xnor U11559 (N_11559,N_10520,N_10270);
or U11560 (N_11560,N_10759,N_10004);
and U11561 (N_11561,N_10535,N_10435);
nand U11562 (N_11562,N_10367,N_10680);
nor U11563 (N_11563,N_10678,N_10517);
nand U11564 (N_11564,N_10649,N_10643);
xnor U11565 (N_11565,N_10892,N_10422);
and U11566 (N_11566,N_10618,N_10205);
xor U11567 (N_11567,N_10921,N_10446);
or U11568 (N_11568,N_10130,N_10138);
nor U11569 (N_11569,N_10482,N_10367);
nor U11570 (N_11570,N_10449,N_10050);
nand U11571 (N_11571,N_10799,N_10462);
nand U11572 (N_11572,N_10525,N_10470);
nor U11573 (N_11573,N_10405,N_10364);
and U11574 (N_11574,N_10740,N_10759);
nand U11575 (N_11575,N_10753,N_10957);
and U11576 (N_11576,N_10633,N_10473);
or U11577 (N_11577,N_10410,N_10618);
nand U11578 (N_11578,N_10287,N_10048);
nor U11579 (N_11579,N_10661,N_10812);
and U11580 (N_11580,N_10025,N_10044);
and U11581 (N_11581,N_10803,N_10891);
nor U11582 (N_11582,N_10151,N_10300);
nand U11583 (N_11583,N_10859,N_10846);
xnor U11584 (N_11584,N_10399,N_10941);
or U11585 (N_11585,N_10817,N_10894);
or U11586 (N_11586,N_10424,N_10765);
and U11587 (N_11587,N_10211,N_10474);
nand U11588 (N_11588,N_10496,N_10670);
nand U11589 (N_11589,N_10982,N_10203);
and U11590 (N_11590,N_10932,N_10322);
and U11591 (N_11591,N_10999,N_10638);
and U11592 (N_11592,N_10721,N_10968);
and U11593 (N_11593,N_10136,N_10823);
nand U11594 (N_11594,N_10624,N_10755);
nor U11595 (N_11595,N_10614,N_10377);
or U11596 (N_11596,N_10969,N_10267);
nor U11597 (N_11597,N_10725,N_10127);
or U11598 (N_11598,N_10832,N_10455);
or U11599 (N_11599,N_10967,N_10826);
and U11600 (N_11600,N_10778,N_10266);
xor U11601 (N_11601,N_10110,N_10507);
nand U11602 (N_11602,N_10682,N_10112);
and U11603 (N_11603,N_10268,N_10743);
and U11604 (N_11604,N_10914,N_10646);
nand U11605 (N_11605,N_10824,N_10349);
nor U11606 (N_11606,N_10037,N_10703);
xor U11607 (N_11607,N_10194,N_10214);
xnor U11608 (N_11608,N_10494,N_10689);
and U11609 (N_11609,N_10630,N_10341);
and U11610 (N_11610,N_10007,N_10661);
nor U11611 (N_11611,N_10348,N_10073);
nor U11612 (N_11612,N_10831,N_10285);
or U11613 (N_11613,N_10110,N_10995);
and U11614 (N_11614,N_10371,N_10177);
xor U11615 (N_11615,N_10041,N_10966);
xor U11616 (N_11616,N_10616,N_10952);
nor U11617 (N_11617,N_10301,N_10516);
xor U11618 (N_11618,N_10859,N_10084);
xnor U11619 (N_11619,N_10761,N_10335);
xnor U11620 (N_11620,N_10123,N_10514);
and U11621 (N_11621,N_10420,N_10082);
nand U11622 (N_11622,N_10700,N_10938);
or U11623 (N_11623,N_10992,N_10528);
nor U11624 (N_11624,N_10657,N_10130);
and U11625 (N_11625,N_10236,N_10780);
nand U11626 (N_11626,N_10159,N_10042);
xor U11627 (N_11627,N_10478,N_10065);
and U11628 (N_11628,N_10363,N_10593);
nor U11629 (N_11629,N_10749,N_10349);
nand U11630 (N_11630,N_10433,N_10740);
and U11631 (N_11631,N_10660,N_10464);
nand U11632 (N_11632,N_10812,N_10701);
nor U11633 (N_11633,N_10520,N_10724);
xor U11634 (N_11634,N_10678,N_10253);
xor U11635 (N_11635,N_10081,N_10837);
or U11636 (N_11636,N_10738,N_10653);
nand U11637 (N_11637,N_10414,N_10504);
or U11638 (N_11638,N_10079,N_10454);
nand U11639 (N_11639,N_10117,N_10687);
nand U11640 (N_11640,N_10915,N_10014);
nor U11641 (N_11641,N_10665,N_10926);
nor U11642 (N_11642,N_10238,N_10780);
nand U11643 (N_11643,N_10598,N_10098);
nand U11644 (N_11644,N_10284,N_10425);
nand U11645 (N_11645,N_10736,N_10300);
and U11646 (N_11646,N_10057,N_10324);
xnor U11647 (N_11647,N_10632,N_10385);
xor U11648 (N_11648,N_10923,N_10815);
or U11649 (N_11649,N_10144,N_10986);
xnor U11650 (N_11650,N_10456,N_10101);
or U11651 (N_11651,N_10104,N_10322);
nor U11652 (N_11652,N_10253,N_10213);
or U11653 (N_11653,N_10427,N_10163);
nor U11654 (N_11654,N_10920,N_10491);
nor U11655 (N_11655,N_10437,N_10769);
nor U11656 (N_11656,N_10224,N_10874);
nand U11657 (N_11657,N_10499,N_10886);
xor U11658 (N_11658,N_10182,N_10220);
nand U11659 (N_11659,N_10560,N_10408);
nand U11660 (N_11660,N_10450,N_10677);
xor U11661 (N_11661,N_10145,N_10259);
nand U11662 (N_11662,N_10863,N_10906);
and U11663 (N_11663,N_10292,N_10280);
nand U11664 (N_11664,N_10359,N_10543);
nor U11665 (N_11665,N_10664,N_10888);
and U11666 (N_11666,N_10346,N_10436);
nand U11667 (N_11667,N_10974,N_10320);
nor U11668 (N_11668,N_10081,N_10142);
or U11669 (N_11669,N_10587,N_10685);
nor U11670 (N_11670,N_10467,N_10889);
xnor U11671 (N_11671,N_10726,N_10161);
or U11672 (N_11672,N_10611,N_10860);
nor U11673 (N_11673,N_10011,N_10881);
xnor U11674 (N_11674,N_10141,N_10072);
nor U11675 (N_11675,N_10381,N_10321);
nor U11676 (N_11676,N_10096,N_10083);
and U11677 (N_11677,N_10403,N_10333);
nor U11678 (N_11678,N_10675,N_10224);
xnor U11679 (N_11679,N_10607,N_10539);
and U11680 (N_11680,N_10777,N_10521);
nand U11681 (N_11681,N_10529,N_10186);
xnor U11682 (N_11682,N_10458,N_10803);
nor U11683 (N_11683,N_10509,N_10947);
nor U11684 (N_11684,N_10532,N_10412);
nor U11685 (N_11685,N_10609,N_10784);
xnor U11686 (N_11686,N_10329,N_10759);
xor U11687 (N_11687,N_10369,N_10029);
nand U11688 (N_11688,N_10163,N_10936);
or U11689 (N_11689,N_10723,N_10920);
and U11690 (N_11690,N_10642,N_10921);
or U11691 (N_11691,N_10068,N_10950);
nand U11692 (N_11692,N_10149,N_10481);
or U11693 (N_11693,N_10626,N_10434);
and U11694 (N_11694,N_10490,N_10879);
nor U11695 (N_11695,N_10197,N_10283);
or U11696 (N_11696,N_10393,N_10694);
and U11697 (N_11697,N_10855,N_10118);
or U11698 (N_11698,N_10909,N_10521);
xnor U11699 (N_11699,N_10908,N_10618);
and U11700 (N_11700,N_10422,N_10692);
and U11701 (N_11701,N_10186,N_10542);
nor U11702 (N_11702,N_10282,N_10789);
nand U11703 (N_11703,N_10445,N_10373);
xnor U11704 (N_11704,N_10031,N_10366);
nand U11705 (N_11705,N_10746,N_10462);
and U11706 (N_11706,N_10206,N_10823);
xnor U11707 (N_11707,N_10218,N_10996);
and U11708 (N_11708,N_10161,N_10273);
nor U11709 (N_11709,N_10234,N_10478);
xor U11710 (N_11710,N_10989,N_10981);
or U11711 (N_11711,N_10504,N_10359);
nand U11712 (N_11712,N_10740,N_10300);
xnor U11713 (N_11713,N_10661,N_10599);
nor U11714 (N_11714,N_10532,N_10801);
and U11715 (N_11715,N_10206,N_10200);
nor U11716 (N_11716,N_10334,N_10738);
and U11717 (N_11717,N_10917,N_10985);
nand U11718 (N_11718,N_10497,N_10651);
or U11719 (N_11719,N_10812,N_10190);
and U11720 (N_11720,N_10971,N_10500);
nand U11721 (N_11721,N_10929,N_10356);
and U11722 (N_11722,N_10559,N_10225);
or U11723 (N_11723,N_10093,N_10403);
and U11724 (N_11724,N_10074,N_10144);
and U11725 (N_11725,N_10924,N_10852);
nor U11726 (N_11726,N_10400,N_10827);
and U11727 (N_11727,N_10423,N_10183);
and U11728 (N_11728,N_10535,N_10983);
nand U11729 (N_11729,N_10947,N_10074);
nor U11730 (N_11730,N_10338,N_10067);
or U11731 (N_11731,N_10416,N_10489);
and U11732 (N_11732,N_10328,N_10850);
nand U11733 (N_11733,N_10295,N_10553);
or U11734 (N_11734,N_10940,N_10225);
xor U11735 (N_11735,N_10135,N_10822);
xnor U11736 (N_11736,N_10551,N_10995);
xnor U11737 (N_11737,N_10330,N_10111);
nor U11738 (N_11738,N_10554,N_10999);
xnor U11739 (N_11739,N_10362,N_10735);
nor U11740 (N_11740,N_10359,N_10162);
and U11741 (N_11741,N_10778,N_10469);
or U11742 (N_11742,N_10405,N_10052);
xnor U11743 (N_11743,N_10273,N_10440);
and U11744 (N_11744,N_10245,N_10613);
nand U11745 (N_11745,N_10795,N_10529);
nor U11746 (N_11746,N_10802,N_10074);
or U11747 (N_11747,N_10663,N_10709);
nand U11748 (N_11748,N_10198,N_10955);
or U11749 (N_11749,N_10336,N_10111);
nand U11750 (N_11750,N_10275,N_10349);
nand U11751 (N_11751,N_10671,N_10205);
nor U11752 (N_11752,N_10410,N_10310);
nor U11753 (N_11753,N_10265,N_10360);
and U11754 (N_11754,N_10927,N_10118);
nor U11755 (N_11755,N_10364,N_10735);
xnor U11756 (N_11756,N_10417,N_10111);
and U11757 (N_11757,N_10416,N_10761);
or U11758 (N_11758,N_10120,N_10459);
xnor U11759 (N_11759,N_10470,N_10307);
and U11760 (N_11760,N_10290,N_10050);
and U11761 (N_11761,N_10763,N_10180);
or U11762 (N_11762,N_10597,N_10422);
and U11763 (N_11763,N_10756,N_10644);
or U11764 (N_11764,N_10960,N_10124);
nand U11765 (N_11765,N_10027,N_10792);
nor U11766 (N_11766,N_10516,N_10272);
nor U11767 (N_11767,N_10720,N_10361);
and U11768 (N_11768,N_10305,N_10424);
xnor U11769 (N_11769,N_10328,N_10454);
or U11770 (N_11770,N_10761,N_10466);
nand U11771 (N_11771,N_10464,N_10313);
nand U11772 (N_11772,N_10567,N_10004);
and U11773 (N_11773,N_10928,N_10788);
nand U11774 (N_11774,N_10005,N_10957);
or U11775 (N_11775,N_10106,N_10184);
nand U11776 (N_11776,N_10091,N_10134);
xor U11777 (N_11777,N_10422,N_10050);
xor U11778 (N_11778,N_10841,N_10884);
or U11779 (N_11779,N_10046,N_10723);
xnor U11780 (N_11780,N_10298,N_10797);
or U11781 (N_11781,N_10049,N_10988);
nand U11782 (N_11782,N_10046,N_10287);
xnor U11783 (N_11783,N_10235,N_10794);
nand U11784 (N_11784,N_10228,N_10636);
nor U11785 (N_11785,N_10750,N_10034);
or U11786 (N_11786,N_10897,N_10770);
and U11787 (N_11787,N_10710,N_10633);
and U11788 (N_11788,N_10896,N_10376);
nor U11789 (N_11789,N_10842,N_10249);
nand U11790 (N_11790,N_10524,N_10640);
or U11791 (N_11791,N_10191,N_10860);
and U11792 (N_11792,N_10684,N_10962);
nor U11793 (N_11793,N_10797,N_10581);
or U11794 (N_11794,N_10008,N_10040);
and U11795 (N_11795,N_10026,N_10112);
nand U11796 (N_11796,N_10137,N_10325);
or U11797 (N_11797,N_10331,N_10276);
xnor U11798 (N_11798,N_10264,N_10311);
nor U11799 (N_11799,N_10468,N_10833);
nor U11800 (N_11800,N_10427,N_10210);
nand U11801 (N_11801,N_10828,N_10180);
and U11802 (N_11802,N_10295,N_10203);
and U11803 (N_11803,N_10540,N_10554);
nand U11804 (N_11804,N_10015,N_10273);
nor U11805 (N_11805,N_10408,N_10562);
or U11806 (N_11806,N_10015,N_10660);
nand U11807 (N_11807,N_10652,N_10734);
nand U11808 (N_11808,N_10396,N_10243);
or U11809 (N_11809,N_10986,N_10239);
nor U11810 (N_11810,N_10182,N_10258);
nand U11811 (N_11811,N_10957,N_10865);
nor U11812 (N_11812,N_10269,N_10441);
nor U11813 (N_11813,N_10178,N_10127);
and U11814 (N_11814,N_10897,N_10051);
xnor U11815 (N_11815,N_10400,N_10287);
nand U11816 (N_11816,N_10159,N_10033);
nand U11817 (N_11817,N_10562,N_10763);
or U11818 (N_11818,N_10263,N_10709);
or U11819 (N_11819,N_10919,N_10501);
and U11820 (N_11820,N_10313,N_10690);
nor U11821 (N_11821,N_10700,N_10609);
xor U11822 (N_11822,N_10485,N_10339);
and U11823 (N_11823,N_10900,N_10487);
nor U11824 (N_11824,N_10371,N_10432);
xor U11825 (N_11825,N_10235,N_10886);
xnor U11826 (N_11826,N_10131,N_10402);
or U11827 (N_11827,N_10087,N_10349);
nand U11828 (N_11828,N_10868,N_10937);
nand U11829 (N_11829,N_10917,N_10374);
or U11830 (N_11830,N_10575,N_10398);
nand U11831 (N_11831,N_10351,N_10095);
xnor U11832 (N_11832,N_10312,N_10505);
xor U11833 (N_11833,N_10340,N_10668);
nand U11834 (N_11834,N_10322,N_10158);
xor U11835 (N_11835,N_10694,N_10572);
nand U11836 (N_11836,N_10485,N_10841);
and U11837 (N_11837,N_10515,N_10050);
xnor U11838 (N_11838,N_10733,N_10315);
nand U11839 (N_11839,N_10080,N_10018);
and U11840 (N_11840,N_10905,N_10372);
xor U11841 (N_11841,N_10665,N_10877);
nand U11842 (N_11842,N_10473,N_10920);
nor U11843 (N_11843,N_10166,N_10769);
xor U11844 (N_11844,N_10056,N_10286);
or U11845 (N_11845,N_10911,N_10086);
nand U11846 (N_11846,N_10626,N_10549);
xnor U11847 (N_11847,N_10938,N_10846);
and U11848 (N_11848,N_10622,N_10627);
or U11849 (N_11849,N_10119,N_10875);
and U11850 (N_11850,N_10754,N_10814);
xnor U11851 (N_11851,N_10793,N_10649);
nor U11852 (N_11852,N_10510,N_10647);
nor U11853 (N_11853,N_10781,N_10287);
and U11854 (N_11854,N_10649,N_10025);
nor U11855 (N_11855,N_10417,N_10502);
and U11856 (N_11856,N_10580,N_10379);
or U11857 (N_11857,N_10548,N_10424);
xnor U11858 (N_11858,N_10935,N_10209);
or U11859 (N_11859,N_10945,N_10601);
xnor U11860 (N_11860,N_10897,N_10217);
and U11861 (N_11861,N_10404,N_10538);
or U11862 (N_11862,N_10282,N_10568);
nand U11863 (N_11863,N_10692,N_10965);
nand U11864 (N_11864,N_10236,N_10674);
nand U11865 (N_11865,N_10565,N_10003);
nand U11866 (N_11866,N_10566,N_10849);
nor U11867 (N_11867,N_10482,N_10683);
or U11868 (N_11868,N_10297,N_10446);
and U11869 (N_11869,N_10612,N_10775);
xor U11870 (N_11870,N_10505,N_10699);
or U11871 (N_11871,N_10738,N_10186);
xnor U11872 (N_11872,N_10677,N_10511);
xnor U11873 (N_11873,N_10157,N_10689);
nor U11874 (N_11874,N_10285,N_10010);
and U11875 (N_11875,N_10650,N_10544);
nand U11876 (N_11876,N_10482,N_10939);
or U11877 (N_11877,N_10518,N_10691);
or U11878 (N_11878,N_10536,N_10348);
nor U11879 (N_11879,N_10338,N_10665);
xor U11880 (N_11880,N_10927,N_10936);
nor U11881 (N_11881,N_10396,N_10982);
nor U11882 (N_11882,N_10999,N_10400);
nor U11883 (N_11883,N_10736,N_10403);
and U11884 (N_11884,N_10460,N_10203);
nor U11885 (N_11885,N_10188,N_10642);
xnor U11886 (N_11886,N_10481,N_10827);
nand U11887 (N_11887,N_10842,N_10648);
nand U11888 (N_11888,N_10103,N_10096);
or U11889 (N_11889,N_10995,N_10118);
nor U11890 (N_11890,N_10792,N_10983);
or U11891 (N_11891,N_10471,N_10872);
nand U11892 (N_11892,N_10782,N_10509);
nand U11893 (N_11893,N_10640,N_10471);
nor U11894 (N_11894,N_10636,N_10704);
or U11895 (N_11895,N_10368,N_10635);
nand U11896 (N_11896,N_10002,N_10709);
or U11897 (N_11897,N_10697,N_10376);
nand U11898 (N_11898,N_10869,N_10151);
and U11899 (N_11899,N_10361,N_10448);
or U11900 (N_11900,N_10105,N_10985);
nor U11901 (N_11901,N_10858,N_10746);
and U11902 (N_11902,N_10391,N_10509);
nor U11903 (N_11903,N_10048,N_10585);
or U11904 (N_11904,N_10018,N_10638);
or U11905 (N_11905,N_10392,N_10331);
or U11906 (N_11906,N_10606,N_10187);
or U11907 (N_11907,N_10141,N_10836);
xnor U11908 (N_11908,N_10828,N_10450);
nor U11909 (N_11909,N_10582,N_10807);
or U11910 (N_11910,N_10372,N_10839);
and U11911 (N_11911,N_10089,N_10065);
nand U11912 (N_11912,N_10032,N_10735);
and U11913 (N_11913,N_10175,N_10854);
nand U11914 (N_11914,N_10672,N_10798);
nor U11915 (N_11915,N_10098,N_10441);
or U11916 (N_11916,N_10850,N_10999);
xnor U11917 (N_11917,N_10010,N_10233);
xor U11918 (N_11918,N_10153,N_10126);
or U11919 (N_11919,N_10458,N_10159);
xor U11920 (N_11920,N_10135,N_10588);
or U11921 (N_11921,N_10911,N_10448);
and U11922 (N_11922,N_10369,N_10795);
and U11923 (N_11923,N_10230,N_10408);
nand U11924 (N_11924,N_10529,N_10969);
and U11925 (N_11925,N_10122,N_10442);
or U11926 (N_11926,N_10036,N_10448);
nor U11927 (N_11927,N_10123,N_10827);
and U11928 (N_11928,N_10401,N_10671);
nor U11929 (N_11929,N_10166,N_10246);
xor U11930 (N_11930,N_10303,N_10218);
xor U11931 (N_11931,N_10702,N_10713);
or U11932 (N_11932,N_10842,N_10269);
xnor U11933 (N_11933,N_10358,N_10781);
or U11934 (N_11934,N_10471,N_10304);
or U11935 (N_11935,N_10470,N_10680);
nand U11936 (N_11936,N_10706,N_10999);
nor U11937 (N_11937,N_10605,N_10964);
xnor U11938 (N_11938,N_10633,N_10645);
and U11939 (N_11939,N_10181,N_10596);
or U11940 (N_11940,N_10292,N_10093);
and U11941 (N_11941,N_10388,N_10393);
nand U11942 (N_11942,N_10639,N_10297);
or U11943 (N_11943,N_10367,N_10017);
xor U11944 (N_11944,N_10422,N_10903);
and U11945 (N_11945,N_10348,N_10241);
xnor U11946 (N_11946,N_10864,N_10677);
nor U11947 (N_11947,N_10194,N_10804);
or U11948 (N_11948,N_10319,N_10018);
nor U11949 (N_11949,N_10848,N_10087);
nand U11950 (N_11950,N_10970,N_10429);
and U11951 (N_11951,N_10058,N_10452);
or U11952 (N_11952,N_10291,N_10162);
and U11953 (N_11953,N_10800,N_10698);
nand U11954 (N_11954,N_10422,N_10636);
nor U11955 (N_11955,N_10364,N_10361);
nand U11956 (N_11956,N_10135,N_10887);
and U11957 (N_11957,N_10722,N_10026);
nor U11958 (N_11958,N_10612,N_10579);
xnor U11959 (N_11959,N_10267,N_10120);
xor U11960 (N_11960,N_10730,N_10895);
or U11961 (N_11961,N_10829,N_10179);
nor U11962 (N_11962,N_10646,N_10751);
nand U11963 (N_11963,N_10264,N_10580);
xnor U11964 (N_11964,N_10805,N_10361);
and U11965 (N_11965,N_10449,N_10552);
nand U11966 (N_11966,N_10128,N_10689);
xnor U11967 (N_11967,N_10127,N_10275);
nor U11968 (N_11968,N_10140,N_10503);
nor U11969 (N_11969,N_10397,N_10370);
and U11970 (N_11970,N_10800,N_10307);
xor U11971 (N_11971,N_10138,N_10915);
and U11972 (N_11972,N_10270,N_10742);
and U11973 (N_11973,N_10662,N_10317);
nand U11974 (N_11974,N_10521,N_10644);
nand U11975 (N_11975,N_10225,N_10161);
or U11976 (N_11976,N_10826,N_10098);
nand U11977 (N_11977,N_10796,N_10054);
or U11978 (N_11978,N_10079,N_10739);
or U11979 (N_11979,N_10986,N_10459);
and U11980 (N_11980,N_10601,N_10555);
or U11981 (N_11981,N_10594,N_10466);
xor U11982 (N_11982,N_10721,N_10058);
nor U11983 (N_11983,N_10796,N_10922);
and U11984 (N_11984,N_10212,N_10948);
xor U11985 (N_11985,N_10996,N_10806);
nand U11986 (N_11986,N_10940,N_10700);
nor U11987 (N_11987,N_10308,N_10635);
nor U11988 (N_11988,N_10630,N_10058);
and U11989 (N_11989,N_10391,N_10988);
nand U11990 (N_11990,N_10135,N_10900);
xnor U11991 (N_11991,N_10948,N_10069);
and U11992 (N_11992,N_10024,N_10318);
xnor U11993 (N_11993,N_10710,N_10771);
or U11994 (N_11994,N_10713,N_10320);
xnor U11995 (N_11995,N_10824,N_10857);
nand U11996 (N_11996,N_10752,N_10779);
or U11997 (N_11997,N_10786,N_10114);
or U11998 (N_11998,N_10016,N_10347);
nand U11999 (N_11999,N_10135,N_10363);
nand U12000 (N_12000,N_11467,N_11203);
nand U12001 (N_12001,N_11630,N_11275);
or U12002 (N_12002,N_11712,N_11673);
and U12003 (N_12003,N_11551,N_11047);
nor U12004 (N_12004,N_11483,N_11652);
nor U12005 (N_12005,N_11296,N_11651);
and U12006 (N_12006,N_11852,N_11675);
nor U12007 (N_12007,N_11092,N_11858);
and U12008 (N_12008,N_11680,N_11164);
and U12009 (N_12009,N_11685,N_11141);
nand U12010 (N_12010,N_11476,N_11072);
nor U12011 (N_12011,N_11801,N_11109);
xnor U12012 (N_12012,N_11155,N_11174);
xnor U12013 (N_12013,N_11175,N_11715);
or U12014 (N_12014,N_11495,N_11977);
xor U12015 (N_12015,N_11487,N_11748);
xnor U12016 (N_12016,N_11116,N_11714);
and U12017 (N_12017,N_11118,N_11128);
xor U12018 (N_12018,N_11833,N_11081);
nor U12019 (N_12019,N_11716,N_11181);
and U12020 (N_12020,N_11364,N_11247);
nand U12021 (N_12021,N_11202,N_11733);
or U12022 (N_12022,N_11307,N_11271);
and U12023 (N_12023,N_11731,N_11260);
nand U12024 (N_12024,N_11370,N_11310);
or U12025 (N_12025,N_11200,N_11432);
xor U12026 (N_12026,N_11624,N_11626);
nand U12027 (N_12027,N_11071,N_11008);
nor U12028 (N_12028,N_11914,N_11779);
xnor U12029 (N_12029,N_11736,N_11573);
or U12030 (N_12030,N_11864,N_11887);
or U12031 (N_12031,N_11287,N_11598);
nor U12032 (N_12032,N_11967,N_11760);
nor U12033 (N_12033,N_11208,N_11187);
nand U12034 (N_12034,N_11042,N_11322);
xor U12035 (N_12035,N_11439,N_11683);
or U12036 (N_12036,N_11284,N_11509);
nor U12037 (N_12037,N_11461,N_11125);
nor U12038 (N_12038,N_11418,N_11923);
and U12039 (N_12039,N_11829,N_11752);
nand U12040 (N_12040,N_11941,N_11514);
or U12041 (N_12041,N_11412,N_11453);
or U12042 (N_12042,N_11798,N_11448);
xor U12043 (N_12043,N_11191,N_11520);
and U12044 (N_12044,N_11304,N_11906);
and U12045 (N_12045,N_11216,N_11342);
nand U12046 (N_12046,N_11353,N_11654);
and U12047 (N_12047,N_11761,N_11366);
nand U12048 (N_12048,N_11783,N_11215);
nor U12049 (N_12049,N_11728,N_11511);
or U12050 (N_12050,N_11534,N_11268);
and U12051 (N_12051,N_11340,N_11985);
nand U12052 (N_12052,N_11740,N_11237);
xor U12053 (N_12053,N_11111,N_11017);
xnor U12054 (N_12054,N_11006,N_11501);
nor U12055 (N_12055,N_11754,N_11455);
nor U12056 (N_12056,N_11359,N_11242);
nand U12057 (N_12057,N_11180,N_11007);
nor U12058 (N_12058,N_11688,N_11171);
or U12059 (N_12059,N_11670,N_11085);
and U12060 (N_12060,N_11606,N_11818);
or U12061 (N_12061,N_11096,N_11751);
nand U12062 (N_12062,N_11568,N_11547);
xor U12063 (N_12063,N_11472,N_11037);
and U12064 (N_12064,N_11621,N_11192);
and U12065 (N_12065,N_11756,N_11479);
nor U12066 (N_12066,N_11417,N_11392);
nand U12067 (N_12067,N_11556,N_11857);
or U12068 (N_12068,N_11622,N_11320);
nor U12069 (N_12069,N_11146,N_11594);
and U12070 (N_12070,N_11947,N_11734);
and U12071 (N_12071,N_11302,N_11213);
nor U12072 (N_12072,N_11648,N_11710);
xor U12073 (N_12073,N_11542,N_11350);
or U12074 (N_12074,N_11363,N_11639);
nand U12075 (N_12075,N_11659,N_11936);
nand U12076 (N_12076,N_11229,N_11299);
xor U12077 (N_12077,N_11014,N_11574);
or U12078 (N_12078,N_11442,N_11387);
xor U12079 (N_12079,N_11196,N_11951);
nor U12080 (N_12080,N_11324,N_11904);
or U12081 (N_12081,N_11823,N_11845);
xor U12082 (N_12082,N_11793,N_11438);
or U12083 (N_12083,N_11078,N_11348);
nand U12084 (N_12084,N_11620,N_11462);
and U12085 (N_12085,N_11226,N_11609);
and U12086 (N_12086,N_11984,N_11671);
and U12087 (N_12087,N_11494,N_11976);
and U12088 (N_12088,N_11170,N_11650);
xnor U12089 (N_12089,N_11532,N_11486);
xor U12090 (N_12090,N_11381,N_11787);
nand U12091 (N_12091,N_11571,N_11988);
xor U12092 (N_12092,N_11935,N_11682);
and U12093 (N_12093,N_11747,N_11335);
nand U12094 (N_12094,N_11137,N_11429);
xor U12095 (N_12095,N_11896,N_11909);
nor U12096 (N_12096,N_11293,N_11173);
nor U12097 (N_12097,N_11944,N_11323);
xnor U12098 (N_12098,N_11261,N_11677);
or U12099 (N_12099,N_11450,N_11510);
or U12100 (N_12100,N_11378,N_11055);
or U12101 (N_12101,N_11603,N_11145);
xnor U12102 (N_12102,N_11653,N_11668);
xnor U12103 (N_12103,N_11953,N_11874);
nand U12104 (N_12104,N_11778,N_11218);
xnor U12105 (N_12105,N_11054,N_11934);
nor U12106 (N_12106,N_11662,N_11924);
or U12107 (N_12107,N_11182,N_11178);
nor U12108 (N_12108,N_11545,N_11357);
nand U12109 (N_12109,N_11552,N_11913);
and U12110 (N_12110,N_11836,N_11349);
xor U12111 (N_12111,N_11385,N_11640);
and U12112 (N_12112,N_11837,N_11217);
or U12113 (N_12113,N_11308,N_11029);
and U12114 (N_12114,N_11251,N_11372);
and U12115 (N_12115,N_11133,N_11883);
nand U12116 (N_12116,N_11138,N_11537);
and U12117 (N_12117,N_11591,N_11456);
and U12118 (N_12118,N_11679,N_11123);
nor U12119 (N_12119,N_11828,N_11023);
or U12120 (N_12120,N_11341,N_11958);
nor U12121 (N_12121,N_11800,N_11035);
and U12122 (N_12122,N_11223,N_11488);
nand U12123 (N_12123,N_11559,N_11315);
or U12124 (N_12124,N_11420,N_11356);
and U12125 (N_12125,N_11068,N_11497);
xnor U12126 (N_12126,N_11295,N_11666);
xnor U12127 (N_12127,N_11755,N_11794);
nand U12128 (N_12128,N_11692,N_11777);
xor U12129 (N_12129,N_11886,N_11233);
nand U12130 (N_12130,N_11469,N_11615);
and U12131 (N_12131,N_11930,N_11767);
and U12132 (N_12132,N_11262,N_11028);
nand U12133 (N_12133,N_11563,N_11291);
nand U12134 (N_12134,N_11012,N_11610);
and U12135 (N_12135,N_11239,N_11691);
nand U12136 (N_12136,N_11409,N_11865);
nor U12137 (N_12137,N_11139,N_11795);
nand U12138 (N_12138,N_11707,N_11144);
nor U12139 (N_12139,N_11234,N_11780);
nor U12140 (N_12140,N_11204,N_11797);
or U12141 (N_12141,N_11721,N_11278);
nand U12142 (N_12142,N_11269,N_11088);
and U12143 (N_12143,N_11541,N_11148);
xor U12144 (N_12144,N_11980,N_11880);
nand U12145 (N_12145,N_11523,N_11910);
nor U12146 (N_12146,N_11916,N_11709);
nor U12147 (N_12147,N_11879,N_11881);
nor U12148 (N_12148,N_11533,N_11219);
nor U12149 (N_12149,N_11562,N_11264);
nand U12150 (N_12150,N_11373,N_11664);
or U12151 (N_12151,N_11990,N_11112);
nand U12152 (N_12152,N_11513,N_11386);
or U12153 (N_12153,N_11946,N_11190);
nor U12154 (N_12154,N_11343,N_11838);
or U12155 (N_12155,N_11013,N_11784);
nand U12156 (N_12156,N_11531,N_11704);
nor U12157 (N_12157,N_11843,N_11831);
and U12158 (N_12158,N_11389,N_11991);
nand U12159 (N_12159,N_11592,N_11207);
nand U12160 (N_12160,N_11079,N_11926);
or U12161 (N_12161,N_11451,N_11711);
xnor U12162 (N_12162,N_11873,N_11806);
xnor U12163 (N_12163,N_11056,N_11086);
nor U12164 (N_12164,N_11119,N_11500);
xor U12165 (N_12165,N_11863,N_11333);
nor U12166 (N_12166,N_11397,N_11866);
or U12167 (N_12167,N_11026,N_11222);
nand U12168 (N_12168,N_11994,N_11297);
or U12169 (N_12169,N_11940,N_11582);
and U12170 (N_12170,N_11195,N_11974);
nor U12171 (N_12171,N_11318,N_11376);
nand U12172 (N_12172,N_11063,N_11430);
nand U12173 (N_12173,N_11903,N_11665);
nand U12174 (N_12174,N_11585,N_11498);
or U12175 (N_12175,N_11782,N_11027);
xor U12176 (N_12176,N_11150,N_11809);
or U12177 (N_12177,N_11314,N_11775);
xnor U12178 (N_12178,N_11834,N_11978);
nand U12179 (N_12179,N_11311,N_11546);
or U12180 (N_12180,N_11550,N_11766);
nor U12181 (N_12181,N_11328,N_11928);
xor U12182 (N_12182,N_11720,N_11177);
nor U12183 (N_12183,N_11435,N_11996);
and U12184 (N_12184,N_11205,N_11243);
nand U12185 (N_12185,N_11095,N_11949);
or U12186 (N_12186,N_11558,N_11601);
and U12187 (N_12187,N_11898,N_11176);
nor U12188 (N_12188,N_11030,N_11750);
xnor U12189 (N_12189,N_11628,N_11280);
nor U12190 (N_12190,N_11010,N_11312);
xor U12191 (N_12191,N_11194,N_11584);
and U12192 (N_12192,N_11566,N_11244);
and U12193 (N_12193,N_11768,N_11152);
nand U12194 (N_12194,N_11839,N_11238);
or U12195 (N_12195,N_11301,N_11437);
nand U12196 (N_12196,N_11365,N_11266);
or U12197 (N_12197,N_11443,N_11022);
nand U12198 (N_12198,N_11273,N_11169);
nor U12199 (N_12199,N_11396,N_11950);
nor U12200 (N_12200,N_11764,N_11143);
xor U12201 (N_12201,N_11334,N_11127);
nor U12202 (N_12202,N_11745,N_11188);
nand U12203 (N_12203,N_11856,N_11762);
or U12204 (N_12204,N_11306,N_11292);
and U12205 (N_12205,N_11832,N_11231);
nand U12206 (N_12206,N_11769,N_11894);
nand U12207 (N_12207,N_11093,N_11912);
nor U12208 (N_12208,N_11586,N_11371);
nand U12209 (N_12209,N_11632,N_11960);
nor U12210 (N_12210,N_11588,N_11465);
xor U12211 (N_12211,N_11637,N_11475);
or U12212 (N_12212,N_11059,N_11607);
and U12213 (N_12213,N_11701,N_11581);
nand U12214 (N_12214,N_11104,N_11230);
nand U12215 (N_12215,N_11629,N_11744);
nand U12216 (N_12216,N_11590,N_11694);
xnor U12217 (N_12217,N_11004,N_11957);
xnor U12218 (N_12218,N_11115,N_11616);
or U12219 (N_12219,N_11689,N_11519);
nand U12220 (N_12220,N_11065,N_11993);
or U12221 (N_12221,N_11792,N_11868);
and U12222 (N_12222,N_11623,N_11159);
xnor U12223 (N_12223,N_11053,N_11454);
nand U12224 (N_12224,N_11384,N_11331);
or U12225 (N_12225,N_11048,N_11725);
nor U12226 (N_12226,N_11436,N_11038);
nand U12227 (N_12227,N_11773,N_11419);
xnor U12228 (N_12228,N_11102,N_11021);
and U12229 (N_12229,N_11132,N_11433);
or U12230 (N_12230,N_11851,N_11485);
and U12231 (N_12231,N_11527,N_11032);
nand U12232 (N_12232,N_11530,N_11423);
nor U12233 (N_12233,N_11379,N_11228);
nand U12234 (N_12234,N_11872,N_11739);
nor U12235 (N_12235,N_11303,N_11221);
or U12236 (N_12236,N_11158,N_11000);
xnor U12237 (N_12237,N_11841,N_11339);
nand U12238 (N_12238,N_11827,N_11713);
or U12239 (N_12239,N_11406,N_11478);
nor U12240 (N_12240,N_11763,N_11110);
and U12241 (N_12241,N_11270,N_11258);
xnor U12242 (N_12242,N_11512,N_11041);
nor U12243 (N_12243,N_11708,N_11161);
nand U12244 (N_12244,N_11289,N_11625);
xnor U12245 (N_12245,N_11998,N_11189);
xor U12246 (N_12246,N_11253,N_11122);
xnor U12247 (N_12247,N_11759,N_11252);
nand U12248 (N_12248,N_11888,N_11987);
or U12249 (N_12249,N_11964,N_11791);
nor U12250 (N_12250,N_11460,N_11403);
or U12251 (N_12251,N_11254,N_11599);
nor U12252 (N_12252,N_11248,N_11565);
and U12253 (N_12253,N_11210,N_11447);
nor U12254 (N_12254,N_11540,N_11617);
nor U12255 (N_12255,N_11724,N_11415);
and U12256 (N_12256,N_11660,N_11405);
nand U12257 (N_12257,N_11272,N_11702);
or U12258 (N_12258,N_11193,N_11646);
nand U12259 (N_12259,N_11877,N_11698);
nor U12260 (N_12260,N_11643,N_11062);
or U12261 (N_12261,N_11893,N_11050);
nor U12262 (N_12262,N_11089,N_11388);
xor U12263 (N_12263,N_11185,N_11165);
and U12264 (N_12264,N_11596,N_11965);
and U12265 (N_12265,N_11332,N_11224);
or U12266 (N_12266,N_11686,N_11718);
nor U12267 (N_12267,N_11570,N_11464);
and U12268 (N_12268,N_11220,N_11235);
and U12269 (N_12269,N_11799,N_11250);
nor U12270 (N_12270,N_11847,N_11211);
or U12271 (N_12271,N_11362,N_11920);
and U12272 (N_12272,N_11066,N_11700);
or U12273 (N_12273,N_11099,N_11649);
nor U12274 (N_12274,N_11168,N_11561);
xnor U12275 (N_12275,N_11058,N_11618);
or U12276 (N_12276,N_11608,N_11882);
or U12277 (N_12277,N_11410,N_11466);
and U12278 (N_12278,N_11867,N_11457);
nand U12279 (N_12279,N_11166,N_11094);
or U12280 (N_12280,N_11862,N_11149);
nand U12281 (N_12281,N_11087,N_11674);
xnor U12282 (N_12282,N_11484,N_11667);
nand U12283 (N_12283,N_11826,N_11080);
and U12284 (N_12284,N_11070,N_11549);
or U12285 (N_12285,N_11730,N_11286);
and U12286 (N_12286,N_11493,N_11846);
nand U12287 (N_12287,N_11699,N_11595);
or U12288 (N_12288,N_11597,N_11274);
nor U12289 (N_12289,N_11481,N_11232);
nor U12290 (N_12290,N_11140,N_11426);
nor U12291 (N_12291,N_11113,N_11580);
nand U12292 (N_12292,N_11383,N_11503);
xnor U12293 (N_12293,N_11516,N_11647);
xor U12294 (N_12294,N_11645,N_11449);
nand U12295 (N_12295,N_11979,N_11124);
or U12296 (N_12296,N_11589,N_11298);
nor U12297 (N_12297,N_11183,N_11121);
or U12298 (N_12298,N_11933,N_11108);
xor U12299 (N_12299,N_11130,N_11074);
nand U12300 (N_12300,N_11458,N_11075);
nand U12301 (N_12301,N_11288,N_11101);
nor U12302 (N_12302,N_11840,N_11817);
nand U12303 (N_12303,N_11908,N_11199);
nor U12304 (N_12304,N_11490,N_11945);
and U12305 (N_12305,N_11536,N_11576);
or U12306 (N_12306,N_11690,N_11395);
nor U12307 (N_12307,N_11198,N_11502);
and U12308 (N_12308,N_11696,N_11695);
nor U12309 (N_12309,N_11360,N_11572);
and U12310 (N_12310,N_11434,N_11678);
nor U12311 (N_12311,N_11895,N_11738);
xor U12312 (N_12312,N_11876,N_11635);
and U12313 (N_12313,N_11100,N_11508);
and U12314 (N_12314,N_11861,N_11788);
nor U12315 (N_12315,N_11741,N_11614);
or U12316 (N_12316,N_11044,N_11179);
nor U12317 (N_12317,N_11361,N_11020);
nand U12318 (N_12318,N_11970,N_11236);
nor U12319 (N_12319,N_11517,N_11019);
and U12320 (N_12320,N_11687,N_11822);
nor U12321 (N_12321,N_11672,N_11153);
nor U12322 (N_12322,N_11459,N_11470);
or U12323 (N_12323,N_11040,N_11742);
nand U12324 (N_12324,N_11214,N_11844);
or U12325 (N_12325,N_11555,N_11544);
xor U12326 (N_12326,N_11636,N_11084);
and U12327 (N_12327,N_11316,N_11212);
nand U12328 (N_12328,N_11382,N_11619);
and U12329 (N_12329,N_11956,N_11963);
and U12330 (N_12330,N_11681,N_11375);
xor U12331 (N_12331,N_11521,N_11989);
nand U12332 (N_12332,N_11142,N_11612);
nand U12333 (N_12333,N_11564,N_11962);
nand U12334 (N_12334,N_11515,N_11758);
and U12335 (N_12335,N_11390,N_11676);
and U12336 (N_12336,N_11727,N_11154);
nor U12337 (N_12337,N_11401,N_11391);
xnor U12338 (N_12338,N_11206,N_11034);
xnor U12339 (N_12339,N_11067,N_11524);
nand U12340 (N_12340,N_11285,N_11107);
or U12341 (N_12341,N_11404,N_11669);
or U12342 (N_12342,N_11411,N_11538);
and U12343 (N_12343,N_11813,N_11528);
xor U12344 (N_12344,N_11553,N_11703);
xnor U12345 (N_12345,N_11255,N_11186);
nor U12346 (N_12346,N_11400,N_11352);
and U12347 (N_12347,N_11684,N_11518);
and U12348 (N_12348,N_11560,N_11380);
or U12349 (N_12349,N_11942,N_11283);
or U12350 (N_12350,N_11575,N_11753);
or U12351 (N_12351,N_11927,N_11117);
or U12352 (N_12352,N_11808,N_11824);
and U12353 (N_12353,N_11329,N_11917);
and U12354 (N_12354,N_11016,N_11735);
nor U12355 (N_12355,N_11441,N_11644);
nand U12356 (N_12356,N_11911,N_11162);
or U12357 (N_12357,N_11638,N_11491);
nor U12358 (N_12358,N_11983,N_11024);
xor U12359 (N_12359,N_11240,N_11003);
or U12360 (N_12360,N_11507,N_11245);
and U12361 (N_12361,N_11358,N_11971);
or U12362 (N_12362,N_11046,N_11605);
xor U12363 (N_12363,N_11120,N_11959);
xor U12364 (N_12364,N_11445,N_11830);
nor U12365 (N_12365,N_11772,N_11408);
and U12366 (N_12366,N_11633,N_11265);
and U12367 (N_12367,N_11083,N_11069);
nand U12368 (N_12368,N_11746,N_11557);
nand U12369 (N_12369,N_11480,N_11554);
nand U12370 (N_12370,N_11136,N_11925);
nor U12371 (N_12371,N_11197,N_11002);
and U12372 (N_12372,N_11351,N_11090);
nand U12373 (N_12373,N_11025,N_11897);
and U12374 (N_12374,N_11249,N_11870);
and U12375 (N_12375,N_11398,N_11871);
or U12376 (N_12376,N_11001,N_11992);
xor U12377 (N_12377,N_11076,N_11593);
and U12378 (N_12378,N_11820,N_11835);
and U12379 (N_12379,N_11786,N_11889);
or U12380 (N_12380,N_11103,N_11627);
or U12381 (N_12381,N_11539,N_11869);
xnor U12382 (N_12382,N_11961,N_11267);
or U12383 (N_12383,N_11948,N_11496);
and U12384 (N_12384,N_11354,N_11878);
or U12385 (N_12385,N_11172,N_11804);
nor U12386 (N_12386,N_11812,N_11317);
or U12387 (N_12387,N_11663,N_11693);
or U12388 (N_12388,N_11902,N_11567);
nand U12389 (N_12389,N_11770,N_11729);
and U12390 (N_12390,N_11452,N_11431);
nand U12391 (N_12391,N_11717,N_11129);
nor U12392 (N_12392,N_11548,N_11057);
nor U12393 (N_12393,N_11135,N_11427);
nand U12394 (N_12394,N_11757,N_11325);
or U12395 (N_12395,N_11337,N_11091);
or U12396 (N_12396,N_11504,N_11468);
nor U12397 (N_12397,N_11973,N_11931);
and U12398 (N_12398,N_11814,N_11526);
nor U12399 (N_12399,N_11241,N_11256);
nand U12400 (N_12400,N_11907,N_11492);
xor U12401 (N_12401,N_11184,N_11899);
nand U12402 (N_12402,N_11807,N_11369);
nand U12403 (N_12403,N_11901,N_11986);
nand U12404 (N_12404,N_11743,N_11005);
or U12405 (N_12405,N_11097,N_11975);
nand U12406 (N_12406,N_11114,N_11969);
nor U12407 (N_12407,N_11859,N_11854);
and U12408 (N_12408,N_11377,N_11082);
xnor U12409 (N_12409,N_11011,N_11631);
nand U12410 (N_12410,N_11522,N_11578);
nand U12411 (N_12411,N_11884,N_11577);
or U12412 (N_12412,N_11073,N_11816);
xnor U12413 (N_12413,N_11105,N_11471);
nand U12414 (N_12414,N_11656,N_11393);
nor U12415 (N_12415,N_11848,N_11602);
and U12416 (N_12416,N_11326,N_11587);
xor U12417 (N_12417,N_11892,N_11855);
or U12418 (N_12418,N_11313,N_11529);
nor U12419 (N_12419,N_11600,N_11999);
nand U12420 (N_12420,N_11319,N_11802);
and U12421 (N_12421,N_11955,N_11446);
xnor U12422 (N_12422,N_11771,N_11276);
or U12423 (N_12423,N_11049,N_11658);
or U12424 (N_12424,N_11282,N_11579);
and U12425 (N_12425,N_11064,N_11416);
nor U12426 (N_12426,N_11425,N_11163);
or U12427 (N_12427,N_11277,N_11294);
nand U12428 (N_12428,N_11891,N_11009);
nor U12429 (N_12429,N_11613,N_11422);
nand U12430 (N_12430,N_11705,N_11167);
and U12431 (N_12431,N_11052,N_11657);
xnor U12432 (N_12432,N_11106,N_11345);
nor U12433 (N_12433,N_11407,N_11305);
xnor U12434 (N_12434,N_11413,N_11932);
and U12435 (N_12435,N_11722,N_11031);
xor U12436 (N_12436,N_11825,N_11790);
or U12437 (N_12437,N_11723,N_11444);
nor U12438 (N_12438,N_11061,N_11915);
xnor U12439 (N_12439,N_11749,N_11367);
nand U12440 (N_12440,N_11972,N_11368);
nand U12441 (N_12441,N_11810,N_11732);
or U12442 (N_12442,N_11330,N_11919);
nand U12443 (N_12443,N_11160,N_11796);
and U12444 (N_12444,N_11850,N_11506);
xnor U12445 (N_12445,N_11815,N_11227);
or U12446 (N_12446,N_11875,N_11921);
nand U12447 (N_12447,N_11505,N_11535);
and U12448 (N_12448,N_11399,N_11300);
xnor U12449 (N_12449,N_11463,N_11655);
nor U12450 (N_12450,N_11344,N_11134);
or U12451 (N_12451,N_11860,N_11604);
nor U12452 (N_12452,N_11355,N_11929);
xor U12453 (N_12453,N_11943,N_11719);
and U12454 (N_12454,N_11785,N_11428);
or U12455 (N_12455,N_11279,N_11938);
nor U12456 (N_12456,N_11905,N_11885);
nand U12457 (N_12457,N_11821,N_11209);
xor U12458 (N_12458,N_11737,N_11151);
nor U12459 (N_12459,N_11954,N_11338);
or U12460 (N_12460,N_11997,N_11394);
or U12461 (N_12461,N_11033,N_11257);
or U12462 (N_12462,N_11321,N_11374);
nor U12463 (N_12463,N_11849,N_11474);
nand U12464 (N_12464,N_11347,N_11131);
xor U12465 (N_12465,N_11890,N_11853);
and U12466 (N_12466,N_11477,N_11968);
or U12467 (N_12467,N_11842,N_11661);
xnor U12468 (N_12468,N_11803,N_11765);
nor U12469 (N_12469,N_11290,N_11499);
nand U12470 (N_12470,N_11819,N_11157);
nor U12471 (N_12471,N_11201,N_11952);
or U12472 (N_12472,N_11077,N_11811);
nor U12473 (N_12473,N_11036,N_11018);
or U12474 (N_12474,N_11045,N_11634);
and U12475 (N_12475,N_11776,N_11147);
nand U12476 (N_12476,N_11440,N_11642);
and U12477 (N_12477,N_11583,N_11336);
nand U12478 (N_12478,N_11939,N_11569);
xor U12479 (N_12479,N_11489,N_11346);
xnor U12480 (N_12480,N_11697,N_11641);
and U12481 (N_12481,N_11706,N_11473);
and U12482 (N_12482,N_11281,N_11543);
nand U12483 (N_12483,N_11043,N_11726);
nand U12484 (N_12484,N_11937,N_11126);
and U12485 (N_12485,N_11982,N_11327);
nand U12486 (N_12486,N_11015,N_11263);
nor U12487 (N_12487,N_11611,N_11482);
nor U12488 (N_12488,N_11922,N_11225);
or U12489 (N_12489,N_11414,N_11981);
nand U12490 (N_12490,N_11918,N_11060);
xnor U12491 (N_12491,N_11774,N_11781);
or U12492 (N_12492,N_11424,N_11098);
nand U12493 (N_12493,N_11966,N_11309);
or U12494 (N_12494,N_11246,N_11039);
xnor U12495 (N_12495,N_11259,N_11421);
or U12496 (N_12496,N_11789,N_11900);
nand U12497 (N_12497,N_11525,N_11156);
xor U12498 (N_12498,N_11995,N_11402);
nor U12499 (N_12499,N_11805,N_11051);
or U12500 (N_12500,N_11134,N_11331);
nand U12501 (N_12501,N_11268,N_11630);
or U12502 (N_12502,N_11440,N_11802);
nor U12503 (N_12503,N_11976,N_11863);
and U12504 (N_12504,N_11543,N_11473);
nor U12505 (N_12505,N_11801,N_11212);
and U12506 (N_12506,N_11555,N_11857);
nand U12507 (N_12507,N_11038,N_11173);
or U12508 (N_12508,N_11922,N_11621);
nor U12509 (N_12509,N_11341,N_11039);
and U12510 (N_12510,N_11443,N_11603);
and U12511 (N_12511,N_11175,N_11631);
nor U12512 (N_12512,N_11796,N_11719);
xnor U12513 (N_12513,N_11024,N_11446);
nor U12514 (N_12514,N_11251,N_11906);
and U12515 (N_12515,N_11216,N_11657);
nand U12516 (N_12516,N_11709,N_11585);
or U12517 (N_12517,N_11320,N_11620);
nand U12518 (N_12518,N_11468,N_11136);
nand U12519 (N_12519,N_11719,N_11465);
or U12520 (N_12520,N_11275,N_11359);
and U12521 (N_12521,N_11223,N_11071);
or U12522 (N_12522,N_11848,N_11020);
or U12523 (N_12523,N_11995,N_11875);
xor U12524 (N_12524,N_11367,N_11764);
xnor U12525 (N_12525,N_11284,N_11500);
nand U12526 (N_12526,N_11559,N_11367);
nor U12527 (N_12527,N_11284,N_11277);
nor U12528 (N_12528,N_11193,N_11087);
xnor U12529 (N_12529,N_11103,N_11415);
or U12530 (N_12530,N_11924,N_11457);
or U12531 (N_12531,N_11423,N_11896);
nand U12532 (N_12532,N_11845,N_11630);
xor U12533 (N_12533,N_11959,N_11547);
nand U12534 (N_12534,N_11391,N_11792);
nor U12535 (N_12535,N_11570,N_11237);
or U12536 (N_12536,N_11472,N_11044);
nand U12537 (N_12537,N_11874,N_11872);
nand U12538 (N_12538,N_11382,N_11844);
xnor U12539 (N_12539,N_11627,N_11580);
nand U12540 (N_12540,N_11405,N_11860);
or U12541 (N_12541,N_11888,N_11170);
and U12542 (N_12542,N_11325,N_11300);
nor U12543 (N_12543,N_11474,N_11688);
xor U12544 (N_12544,N_11616,N_11043);
or U12545 (N_12545,N_11776,N_11884);
or U12546 (N_12546,N_11972,N_11435);
and U12547 (N_12547,N_11915,N_11347);
or U12548 (N_12548,N_11518,N_11552);
xor U12549 (N_12549,N_11016,N_11661);
nor U12550 (N_12550,N_11427,N_11081);
nor U12551 (N_12551,N_11570,N_11198);
nand U12552 (N_12552,N_11245,N_11631);
nand U12553 (N_12553,N_11661,N_11024);
or U12554 (N_12554,N_11513,N_11002);
xnor U12555 (N_12555,N_11185,N_11425);
nand U12556 (N_12556,N_11588,N_11739);
and U12557 (N_12557,N_11010,N_11819);
nor U12558 (N_12558,N_11586,N_11805);
and U12559 (N_12559,N_11568,N_11744);
nor U12560 (N_12560,N_11376,N_11179);
or U12561 (N_12561,N_11360,N_11597);
and U12562 (N_12562,N_11272,N_11635);
and U12563 (N_12563,N_11883,N_11439);
nor U12564 (N_12564,N_11660,N_11945);
xor U12565 (N_12565,N_11779,N_11131);
or U12566 (N_12566,N_11134,N_11068);
nand U12567 (N_12567,N_11680,N_11991);
xor U12568 (N_12568,N_11278,N_11362);
or U12569 (N_12569,N_11323,N_11096);
nor U12570 (N_12570,N_11873,N_11756);
or U12571 (N_12571,N_11898,N_11661);
xnor U12572 (N_12572,N_11113,N_11427);
nand U12573 (N_12573,N_11863,N_11679);
nand U12574 (N_12574,N_11341,N_11456);
nand U12575 (N_12575,N_11036,N_11010);
xor U12576 (N_12576,N_11600,N_11835);
or U12577 (N_12577,N_11515,N_11076);
nor U12578 (N_12578,N_11771,N_11706);
or U12579 (N_12579,N_11122,N_11184);
nor U12580 (N_12580,N_11086,N_11516);
or U12581 (N_12581,N_11902,N_11683);
or U12582 (N_12582,N_11661,N_11771);
nor U12583 (N_12583,N_11250,N_11083);
and U12584 (N_12584,N_11196,N_11609);
xnor U12585 (N_12585,N_11597,N_11323);
or U12586 (N_12586,N_11345,N_11142);
xnor U12587 (N_12587,N_11070,N_11452);
xor U12588 (N_12588,N_11965,N_11589);
xor U12589 (N_12589,N_11698,N_11468);
and U12590 (N_12590,N_11784,N_11466);
and U12591 (N_12591,N_11212,N_11903);
and U12592 (N_12592,N_11536,N_11930);
nand U12593 (N_12593,N_11933,N_11750);
and U12594 (N_12594,N_11494,N_11818);
and U12595 (N_12595,N_11940,N_11576);
nor U12596 (N_12596,N_11277,N_11795);
nor U12597 (N_12597,N_11264,N_11854);
nand U12598 (N_12598,N_11687,N_11680);
nor U12599 (N_12599,N_11380,N_11925);
and U12600 (N_12600,N_11172,N_11926);
xor U12601 (N_12601,N_11655,N_11929);
nor U12602 (N_12602,N_11597,N_11398);
and U12603 (N_12603,N_11835,N_11710);
xor U12604 (N_12604,N_11207,N_11840);
xnor U12605 (N_12605,N_11360,N_11994);
or U12606 (N_12606,N_11253,N_11309);
or U12607 (N_12607,N_11311,N_11898);
nor U12608 (N_12608,N_11343,N_11279);
nor U12609 (N_12609,N_11509,N_11080);
xnor U12610 (N_12610,N_11613,N_11450);
xor U12611 (N_12611,N_11943,N_11703);
nor U12612 (N_12612,N_11390,N_11494);
nor U12613 (N_12613,N_11532,N_11598);
nand U12614 (N_12614,N_11499,N_11317);
nor U12615 (N_12615,N_11946,N_11780);
nor U12616 (N_12616,N_11440,N_11158);
or U12617 (N_12617,N_11770,N_11934);
or U12618 (N_12618,N_11259,N_11764);
xor U12619 (N_12619,N_11662,N_11160);
and U12620 (N_12620,N_11088,N_11749);
or U12621 (N_12621,N_11567,N_11991);
and U12622 (N_12622,N_11992,N_11923);
nor U12623 (N_12623,N_11761,N_11062);
nor U12624 (N_12624,N_11880,N_11448);
nor U12625 (N_12625,N_11610,N_11604);
or U12626 (N_12626,N_11060,N_11234);
nor U12627 (N_12627,N_11034,N_11894);
nand U12628 (N_12628,N_11510,N_11218);
and U12629 (N_12629,N_11913,N_11632);
xor U12630 (N_12630,N_11216,N_11513);
nor U12631 (N_12631,N_11102,N_11776);
xnor U12632 (N_12632,N_11136,N_11838);
nor U12633 (N_12633,N_11844,N_11532);
nor U12634 (N_12634,N_11838,N_11596);
or U12635 (N_12635,N_11419,N_11410);
and U12636 (N_12636,N_11409,N_11203);
nand U12637 (N_12637,N_11003,N_11878);
nor U12638 (N_12638,N_11448,N_11688);
and U12639 (N_12639,N_11704,N_11989);
or U12640 (N_12640,N_11538,N_11877);
and U12641 (N_12641,N_11835,N_11434);
xnor U12642 (N_12642,N_11099,N_11194);
or U12643 (N_12643,N_11028,N_11811);
nand U12644 (N_12644,N_11376,N_11146);
nor U12645 (N_12645,N_11366,N_11238);
xor U12646 (N_12646,N_11475,N_11691);
xor U12647 (N_12647,N_11731,N_11650);
or U12648 (N_12648,N_11537,N_11838);
or U12649 (N_12649,N_11242,N_11537);
nand U12650 (N_12650,N_11254,N_11660);
nor U12651 (N_12651,N_11309,N_11002);
nand U12652 (N_12652,N_11211,N_11951);
nand U12653 (N_12653,N_11019,N_11882);
nand U12654 (N_12654,N_11576,N_11283);
xor U12655 (N_12655,N_11752,N_11590);
and U12656 (N_12656,N_11665,N_11933);
and U12657 (N_12657,N_11280,N_11851);
or U12658 (N_12658,N_11407,N_11835);
or U12659 (N_12659,N_11009,N_11717);
nand U12660 (N_12660,N_11934,N_11652);
or U12661 (N_12661,N_11339,N_11241);
nor U12662 (N_12662,N_11641,N_11025);
xnor U12663 (N_12663,N_11569,N_11202);
or U12664 (N_12664,N_11531,N_11543);
or U12665 (N_12665,N_11069,N_11609);
nand U12666 (N_12666,N_11187,N_11778);
nor U12667 (N_12667,N_11985,N_11565);
nand U12668 (N_12668,N_11361,N_11575);
and U12669 (N_12669,N_11023,N_11408);
and U12670 (N_12670,N_11852,N_11791);
xnor U12671 (N_12671,N_11367,N_11351);
or U12672 (N_12672,N_11437,N_11279);
and U12673 (N_12673,N_11294,N_11233);
nand U12674 (N_12674,N_11118,N_11502);
xnor U12675 (N_12675,N_11649,N_11361);
nor U12676 (N_12676,N_11749,N_11747);
xor U12677 (N_12677,N_11650,N_11020);
nand U12678 (N_12678,N_11656,N_11599);
nand U12679 (N_12679,N_11326,N_11561);
and U12680 (N_12680,N_11549,N_11888);
xor U12681 (N_12681,N_11003,N_11285);
and U12682 (N_12682,N_11821,N_11797);
xor U12683 (N_12683,N_11454,N_11556);
xor U12684 (N_12684,N_11997,N_11823);
or U12685 (N_12685,N_11081,N_11640);
or U12686 (N_12686,N_11946,N_11733);
or U12687 (N_12687,N_11392,N_11423);
nand U12688 (N_12688,N_11245,N_11189);
or U12689 (N_12689,N_11949,N_11633);
nand U12690 (N_12690,N_11170,N_11610);
or U12691 (N_12691,N_11266,N_11788);
or U12692 (N_12692,N_11049,N_11126);
and U12693 (N_12693,N_11236,N_11115);
nand U12694 (N_12694,N_11844,N_11691);
or U12695 (N_12695,N_11985,N_11428);
and U12696 (N_12696,N_11780,N_11595);
xor U12697 (N_12697,N_11482,N_11551);
and U12698 (N_12698,N_11746,N_11880);
or U12699 (N_12699,N_11110,N_11706);
nor U12700 (N_12700,N_11153,N_11965);
and U12701 (N_12701,N_11881,N_11590);
nor U12702 (N_12702,N_11269,N_11464);
or U12703 (N_12703,N_11816,N_11568);
xnor U12704 (N_12704,N_11655,N_11337);
nand U12705 (N_12705,N_11829,N_11453);
nor U12706 (N_12706,N_11721,N_11299);
or U12707 (N_12707,N_11285,N_11728);
or U12708 (N_12708,N_11932,N_11358);
nand U12709 (N_12709,N_11590,N_11737);
nor U12710 (N_12710,N_11617,N_11221);
xnor U12711 (N_12711,N_11216,N_11705);
and U12712 (N_12712,N_11760,N_11345);
xor U12713 (N_12713,N_11100,N_11808);
nor U12714 (N_12714,N_11253,N_11456);
nor U12715 (N_12715,N_11978,N_11396);
xor U12716 (N_12716,N_11233,N_11941);
and U12717 (N_12717,N_11857,N_11013);
nand U12718 (N_12718,N_11801,N_11138);
or U12719 (N_12719,N_11834,N_11531);
xor U12720 (N_12720,N_11884,N_11692);
and U12721 (N_12721,N_11642,N_11183);
or U12722 (N_12722,N_11955,N_11732);
or U12723 (N_12723,N_11677,N_11898);
xnor U12724 (N_12724,N_11786,N_11955);
or U12725 (N_12725,N_11976,N_11818);
and U12726 (N_12726,N_11280,N_11696);
xnor U12727 (N_12727,N_11147,N_11991);
nand U12728 (N_12728,N_11770,N_11692);
and U12729 (N_12729,N_11820,N_11729);
nor U12730 (N_12730,N_11126,N_11273);
or U12731 (N_12731,N_11635,N_11878);
xnor U12732 (N_12732,N_11878,N_11423);
xor U12733 (N_12733,N_11129,N_11130);
nand U12734 (N_12734,N_11380,N_11583);
and U12735 (N_12735,N_11150,N_11337);
nor U12736 (N_12736,N_11717,N_11944);
or U12737 (N_12737,N_11871,N_11142);
nand U12738 (N_12738,N_11223,N_11897);
nor U12739 (N_12739,N_11231,N_11729);
and U12740 (N_12740,N_11146,N_11481);
and U12741 (N_12741,N_11516,N_11865);
nand U12742 (N_12742,N_11441,N_11527);
xnor U12743 (N_12743,N_11236,N_11136);
nor U12744 (N_12744,N_11574,N_11096);
and U12745 (N_12745,N_11258,N_11562);
nor U12746 (N_12746,N_11040,N_11825);
and U12747 (N_12747,N_11306,N_11555);
and U12748 (N_12748,N_11368,N_11655);
or U12749 (N_12749,N_11886,N_11179);
or U12750 (N_12750,N_11183,N_11475);
nor U12751 (N_12751,N_11390,N_11721);
nor U12752 (N_12752,N_11908,N_11656);
xnor U12753 (N_12753,N_11108,N_11243);
and U12754 (N_12754,N_11061,N_11966);
nor U12755 (N_12755,N_11702,N_11124);
nand U12756 (N_12756,N_11109,N_11229);
or U12757 (N_12757,N_11636,N_11206);
or U12758 (N_12758,N_11034,N_11075);
or U12759 (N_12759,N_11697,N_11346);
xnor U12760 (N_12760,N_11872,N_11940);
or U12761 (N_12761,N_11225,N_11837);
nand U12762 (N_12762,N_11276,N_11358);
nor U12763 (N_12763,N_11828,N_11386);
nand U12764 (N_12764,N_11198,N_11558);
nor U12765 (N_12765,N_11646,N_11989);
and U12766 (N_12766,N_11642,N_11816);
and U12767 (N_12767,N_11537,N_11818);
or U12768 (N_12768,N_11632,N_11927);
and U12769 (N_12769,N_11119,N_11560);
nand U12770 (N_12770,N_11399,N_11892);
and U12771 (N_12771,N_11272,N_11931);
nor U12772 (N_12772,N_11393,N_11578);
or U12773 (N_12773,N_11579,N_11695);
or U12774 (N_12774,N_11249,N_11854);
or U12775 (N_12775,N_11009,N_11292);
or U12776 (N_12776,N_11909,N_11748);
xnor U12777 (N_12777,N_11297,N_11975);
and U12778 (N_12778,N_11269,N_11992);
or U12779 (N_12779,N_11939,N_11472);
xnor U12780 (N_12780,N_11562,N_11447);
or U12781 (N_12781,N_11499,N_11110);
xor U12782 (N_12782,N_11063,N_11036);
nand U12783 (N_12783,N_11740,N_11737);
nor U12784 (N_12784,N_11551,N_11360);
nor U12785 (N_12785,N_11381,N_11240);
nand U12786 (N_12786,N_11455,N_11123);
nor U12787 (N_12787,N_11773,N_11080);
and U12788 (N_12788,N_11728,N_11630);
nor U12789 (N_12789,N_11867,N_11632);
nand U12790 (N_12790,N_11972,N_11321);
xnor U12791 (N_12791,N_11692,N_11744);
nand U12792 (N_12792,N_11556,N_11049);
or U12793 (N_12793,N_11793,N_11432);
or U12794 (N_12794,N_11768,N_11161);
nor U12795 (N_12795,N_11073,N_11310);
and U12796 (N_12796,N_11687,N_11580);
or U12797 (N_12797,N_11568,N_11114);
xor U12798 (N_12798,N_11606,N_11811);
nor U12799 (N_12799,N_11414,N_11087);
or U12800 (N_12800,N_11706,N_11820);
nand U12801 (N_12801,N_11939,N_11113);
and U12802 (N_12802,N_11639,N_11924);
nor U12803 (N_12803,N_11838,N_11211);
or U12804 (N_12804,N_11390,N_11162);
nor U12805 (N_12805,N_11768,N_11120);
nand U12806 (N_12806,N_11243,N_11492);
xnor U12807 (N_12807,N_11876,N_11610);
and U12808 (N_12808,N_11700,N_11184);
or U12809 (N_12809,N_11353,N_11825);
and U12810 (N_12810,N_11062,N_11621);
xor U12811 (N_12811,N_11405,N_11145);
nand U12812 (N_12812,N_11896,N_11566);
nand U12813 (N_12813,N_11683,N_11574);
nand U12814 (N_12814,N_11601,N_11069);
or U12815 (N_12815,N_11330,N_11466);
xnor U12816 (N_12816,N_11638,N_11586);
or U12817 (N_12817,N_11809,N_11578);
nand U12818 (N_12818,N_11083,N_11256);
nor U12819 (N_12819,N_11796,N_11505);
and U12820 (N_12820,N_11634,N_11942);
nand U12821 (N_12821,N_11049,N_11776);
or U12822 (N_12822,N_11058,N_11965);
or U12823 (N_12823,N_11863,N_11958);
or U12824 (N_12824,N_11656,N_11910);
nand U12825 (N_12825,N_11657,N_11243);
xor U12826 (N_12826,N_11155,N_11312);
xor U12827 (N_12827,N_11307,N_11544);
xor U12828 (N_12828,N_11527,N_11387);
or U12829 (N_12829,N_11277,N_11765);
and U12830 (N_12830,N_11514,N_11949);
and U12831 (N_12831,N_11845,N_11968);
xnor U12832 (N_12832,N_11033,N_11104);
or U12833 (N_12833,N_11146,N_11172);
nand U12834 (N_12834,N_11321,N_11024);
and U12835 (N_12835,N_11880,N_11671);
and U12836 (N_12836,N_11061,N_11273);
and U12837 (N_12837,N_11353,N_11576);
xor U12838 (N_12838,N_11763,N_11762);
nor U12839 (N_12839,N_11352,N_11107);
or U12840 (N_12840,N_11603,N_11504);
xnor U12841 (N_12841,N_11599,N_11905);
xnor U12842 (N_12842,N_11673,N_11567);
nand U12843 (N_12843,N_11387,N_11893);
nor U12844 (N_12844,N_11643,N_11702);
xor U12845 (N_12845,N_11996,N_11616);
nand U12846 (N_12846,N_11257,N_11857);
and U12847 (N_12847,N_11346,N_11396);
and U12848 (N_12848,N_11864,N_11853);
nor U12849 (N_12849,N_11531,N_11340);
or U12850 (N_12850,N_11125,N_11922);
xnor U12851 (N_12851,N_11504,N_11781);
nor U12852 (N_12852,N_11110,N_11122);
nand U12853 (N_12853,N_11613,N_11608);
nand U12854 (N_12854,N_11599,N_11416);
and U12855 (N_12855,N_11899,N_11008);
nor U12856 (N_12856,N_11875,N_11766);
nand U12857 (N_12857,N_11847,N_11481);
and U12858 (N_12858,N_11616,N_11546);
nor U12859 (N_12859,N_11095,N_11189);
xor U12860 (N_12860,N_11421,N_11508);
nor U12861 (N_12861,N_11783,N_11398);
and U12862 (N_12862,N_11008,N_11269);
nand U12863 (N_12863,N_11241,N_11213);
or U12864 (N_12864,N_11867,N_11866);
or U12865 (N_12865,N_11292,N_11416);
and U12866 (N_12866,N_11380,N_11493);
nor U12867 (N_12867,N_11852,N_11506);
nand U12868 (N_12868,N_11798,N_11325);
and U12869 (N_12869,N_11240,N_11962);
nor U12870 (N_12870,N_11827,N_11452);
or U12871 (N_12871,N_11629,N_11636);
nand U12872 (N_12872,N_11338,N_11533);
or U12873 (N_12873,N_11341,N_11069);
or U12874 (N_12874,N_11337,N_11008);
nand U12875 (N_12875,N_11524,N_11992);
and U12876 (N_12876,N_11369,N_11393);
and U12877 (N_12877,N_11023,N_11963);
nand U12878 (N_12878,N_11717,N_11123);
and U12879 (N_12879,N_11509,N_11038);
or U12880 (N_12880,N_11216,N_11763);
nand U12881 (N_12881,N_11498,N_11126);
nand U12882 (N_12882,N_11825,N_11700);
nand U12883 (N_12883,N_11878,N_11078);
xor U12884 (N_12884,N_11713,N_11611);
and U12885 (N_12885,N_11855,N_11085);
or U12886 (N_12886,N_11000,N_11694);
xnor U12887 (N_12887,N_11406,N_11767);
nand U12888 (N_12888,N_11846,N_11489);
or U12889 (N_12889,N_11927,N_11111);
nor U12890 (N_12890,N_11541,N_11322);
and U12891 (N_12891,N_11313,N_11175);
or U12892 (N_12892,N_11720,N_11963);
nor U12893 (N_12893,N_11567,N_11260);
or U12894 (N_12894,N_11996,N_11774);
xnor U12895 (N_12895,N_11004,N_11365);
nor U12896 (N_12896,N_11061,N_11976);
or U12897 (N_12897,N_11376,N_11894);
nand U12898 (N_12898,N_11100,N_11569);
and U12899 (N_12899,N_11810,N_11617);
and U12900 (N_12900,N_11390,N_11952);
nand U12901 (N_12901,N_11823,N_11924);
nand U12902 (N_12902,N_11976,N_11201);
nand U12903 (N_12903,N_11867,N_11147);
xor U12904 (N_12904,N_11935,N_11176);
or U12905 (N_12905,N_11997,N_11323);
xor U12906 (N_12906,N_11274,N_11725);
and U12907 (N_12907,N_11945,N_11871);
and U12908 (N_12908,N_11899,N_11697);
xor U12909 (N_12909,N_11290,N_11172);
nor U12910 (N_12910,N_11780,N_11285);
nor U12911 (N_12911,N_11933,N_11037);
or U12912 (N_12912,N_11632,N_11658);
nand U12913 (N_12913,N_11162,N_11487);
nor U12914 (N_12914,N_11502,N_11888);
xor U12915 (N_12915,N_11891,N_11699);
or U12916 (N_12916,N_11039,N_11370);
and U12917 (N_12917,N_11719,N_11614);
or U12918 (N_12918,N_11186,N_11114);
xor U12919 (N_12919,N_11376,N_11747);
nand U12920 (N_12920,N_11683,N_11425);
or U12921 (N_12921,N_11660,N_11869);
nor U12922 (N_12922,N_11556,N_11552);
and U12923 (N_12923,N_11582,N_11357);
and U12924 (N_12924,N_11717,N_11208);
or U12925 (N_12925,N_11367,N_11095);
nand U12926 (N_12926,N_11371,N_11567);
nor U12927 (N_12927,N_11879,N_11489);
nand U12928 (N_12928,N_11347,N_11693);
or U12929 (N_12929,N_11744,N_11289);
and U12930 (N_12930,N_11992,N_11888);
nor U12931 (N_12931,N_11613,N_11776);
xnor U12932 (N_12932,N_11361,N_11817);
nor U12933 (N_12933,N_11199,N_11390);
xnor U12934 (N_12934,N_11538,N_11370);
or U12935 (N_12935,N_11879,N_11320);
or U12936 (N_12936,N_11777,N_11696);
or U12937 (N_12937,N_11915,N_11018);
xor U12938 (N_12938,N_11019,N_11094);
nor U12939 (N_12939,N_11773,N_11967);
nand U12940 (N_12940,N_11721,N_11755);
or U12941 (N_12941,N_11636,N_11545);
and U12942 (N_12942,N_11178,N_11502);
nand U12943 (N_12943,N_11686,N_11800);
nor U12944 (N_12944,N_11536,N_11471);
xnor U12945 (N_12945,N_11874,N_11840);
nor U12946 (N_12946,N_11274,N_11017);
nor U12947 (N_12947,N_11440,N_11558);
nand U12948 (N_12948,N_11013,N_11174);
and U12949 (N_12949,N_11310,N_11487);
and U12950 (N_12950,N_11844,N_11047);
and U12951 (N_12951,N_11538,N_11023);
nand U12952 (N_12952,N_11828,N_11054);
or U12953 (N_12953,N_11856,N_11209);
nor U12954 (N_12954,N_11672,N_11147);
nand U12955 (N_12955,N_11963,N_11107);
nor U12956 (N_12956,N_11435,N_11948);
and U12957 (N_12957,N_11233,N_11821);
xor U12958 (N_12958,N_11621,N_11756);
nand U12959 (N_12959,N_11592,N_11025);
or U12960 (N_12960,N_11088,N_11031);
nor U12961 (N_12961,N_11284,N_11565);
nor U12962 (N_12962,N_11089,N_11600);
nor U12963 (N_12963,N_11354,N_11241);
xnor U12964 (N_12964,N_11403,N_11220);
nand U12965 (N_12965,N_11533,N_11060);
xor U12966 (N_12966,N_11894,N_11446);
or U12967 (N_12967,N_11770,N_11980);
xnor U12968 (N_12968,N_11128,N_11139);
nor U12969 (N_12969,N_11191,N_11528);
xor U12970 (N_12970,N_11493,N_11010);
nand U12971 (N_12971,N_11351,N_11278);
xor U12972 (N_12972,N_11906,N_11689);
or U12973 (N_12973,N_11761,N_11145);
nand U12974 (N_12974,N_11509,N_11616);
and U12975 (N_12975,N_11810,N_11296);
and U12976 (N_12976,N_11332,N_11060);
nand U12977 (N_12977,N_11304,N_11670);
nor U12978 (N_12978,N_11609,N_11232);
and U12979 (N_12979,N_11394,N_11840);
nor U12980 (N_12980,N_11635,N_11912);
nand U12981 (N_12981,N_11391,N_11640);
nand U12982 (N_12982,N_11674,N_11280);
or U12983 (N_12983,N_11224,N_11564);
nor U12984 (N_12984,N_11143,N_11820);
xor U12985 (N_12985,N_11416,N_11452);
xnor U12986 (N_12986,N_11230,N_11233);
xnor U12987 (N_12987,N_11019,N_11137);
xor U12988 (N_12988,N_11795,N_11784);
and U12989 (N_12989,N_11698,N_11228);
nand U12990 (N_12990,N_11044,N_11467);
xor U12991 (N_12991,N_11640,N_11624);
or U12992 (N_12992,N_11542,N_11257);
nand U12993 (N_12993,N_11016,N_11127);
and U12994 (N_12994,N_11030,N_11483);
or U12995 (N_12995,N_11557,N_11630);
nor U12996 (N_12996,N_11471,N_11237);
or U12997 (N_12997,N_11859,N_11720);
nor U12998 (N_12998,N_11083,N_11562);
and U12999 (N_12999,N_11443,N_11308);
or U13000 (N_13000,N_12635,N_12552);
xnor U13001 (N_13001,N_12451,N_12544);
and U13002 (N_13002,N_12940,N_12172);
nor U13003 (N_13003,N_12641,N_12714);
nand U13004 (N_13004,N_12941,N_12442);
or U13005 (N_13005,N_12511,N_12217);
and U13006 (N_13006,N_12730,N_12043);
nor U13007 (N_13007,N_12454,N_12231);
and U13008 (N_13008,N_12058,N_12411);
or U13009 (N_13009,N_12117,N_12556);
nor U13010 (N_13010,N_12616,N_12580);
nor U13011 (N_13011,N_12783,N_12044);
or U13012 (N_13012,N_12956,N_12663);
nor U13013 (N_13013,N_12294,N_12260);
or U13014 (N_13014,N_12180,N_12393);
and U13015 (N_13015,N_12850,N_12004);
nor U13016 (N_13016,N_12990,N_12258);
and U13017 (N_13017,N_12877,N_12789);
nand U13018 (N_13018,N_12277,N_12984);
or U13019 (N_13019,N_12848,N_12605);
nor U13020 (N_13020,N_12832,N_12950);
nand U13021 (N_13021,N_12200,N_12517);
xor U13022 (N_13022,N_12664,N_12072);
and U13023 (N_13023,N_12887,N_12251);
xnor U13024 (N_13024,N_12570,N_12904);
xnor U13025 (N_13025,N_12286,N_12746);
nand U13026 (N_13026,N_12619,N_12938);
and U13027 (N_13027,N_12086,N_12640);
nor U13028 (N_13028,N_12159,N_12001);
nor U13029 (N_13029,N_12092,N_12825);
and U13030 (N_13030,N_12573,N_12842);
or U13031 (N_13031,N_12829,N_12281);
nand U13032 (N_13032,N_12499,N_12890);
or U13033 (N_13033,N_12710,N_12244);
or U13034 (N_13034,N_12724,N_12997);
or U13035 (N_13035,N_12612,N_12388);
and U13036 (N_13036,N_12684,N_12571);
xnor U13037 (N_13037,N_12741,N_12514);
or U13038 (N_13038,N_12838,N_12207);
nand U13039 (N_13039,N_12740,N_12161);
and U13040 (N_13040,N_12321,N_12192);
or U13041 (N_13041,N_12360,N_12869);
nor U13042 (N_13042,N_12666,N_12711);
or U13043 (N_13043,N_12494,N_12876);
nand U13044 (N_13044,N_12445,N_12343);
or U13045 (N_13045,N_12491,N_12558);
xor U13046 (N_13046,N_12975,N_12475);
or U13047 (N_13047,N_12766,N_12361);
nand U13048 (N_13048,N_12249,N_12079);
or U13049 (N_13049,N_12198,N_12121);
or U13050 (N_13050,N_12218,N_12708);
nand U13051 (N_13051,N_12132,N_12398);
and U13052 (N_13052,N_12028,N_12248);
xnor U13053 (N_13053,N_12501,N_12851);
xnor U13054 (N_13054,N_12670,N_12531);
xnor U13055 (N_13055,N_12939,N_12165);
nor U13056 (N_13056,N_12889,N_12691);
xnor U13057 (N_13057,N_12459,N_12503);
nor U13058 (N_13058,N_12130,N_12137);
nor U13059 (N_13059,N_12696,N_12625);
nor U13060 (N_13060,N_12768,N_12389);
nor U13061 (N_13061,N_12003,N_12386);
or U13062 (N_13062,N_12632,N_12201);
nand U13063 (N_13063,N_12481,N_12733);
nand U13064 (N_13064,N_12845,N_12861);
xor U13065 (N_13065,N_12098,N_12992);
or U13066 (N_13066,N_12588,N_12559);
nor U13067 (N_13067,N_12524,N_12016);
nor U13068 (N_13068,N_12506,N_12094);
nor U13069 (N_13069,N_12444,N_12053);
nand U13070 (N_13070,N_12858,N_12119);
or U13071 (N_13071,N_12408,N_12808);
nor U13072 (N_13072,N_12685,N_12855);
nand U13073 (N_13073,N_12193,N_12278);
xor U13074 (N_13074,N_12776,N_12608);
or U13075 (N_13075,N_12817,N_12572);
and U13076 (N_13076,N_12465,N_12493);
or U13077 (N_13077,N_12377,N_12896);
or U13078 (N_13078,N_12324,N_12177);
or U13079 (N_13079,N_12692,N_12759);
and U13080 (N_13080,N_12924,N_12968);
nor U13081 (N_13081,N_12074,N_12203);
xnor U13082 (N_13082,N_12242,N_12148);
nor U13083 (N_13083,N_12773,N_12282);
or U13084 (N_13084,N_12097,N_12757);
nor U13085 (N_13085,N_12788,N_12857);
or U13086 (N_13086,N_12652,N_12885);
and U13087 (N_13087,N_12843,N_12801);
nor U13088 (N_13088,N_12113,N_12932);
nand U13089 (N_13089,N_12315,N_12156);
xor U13090 (N_13090,N_12256,N_12686);
and U13091 (N_13091,N_12219,N_12308);
and U13092 (N_13092,N_12124,N_12337);
or U13093 (N_13093,N_12657,N_12577);
or U13094 (N_13094,N_12383,N_12178);
nor U13095 (N_13095,N_12373,N_12918);
nor U13096 (N_13096,N_12955,N_12886);
nand U13097 (N_13097,N_12152,N_12881);
and U13098 (N_13098,N_12407,N_12909);
nand U13099 (N_13099,N_12934,N_12205);
nand U13100 (N_13100,N_12923,N_12257);
or U13101 (N_13101,N_12457,N_12913);
and U13102 (N_13102,N_12742,N_12611);
or U13103 (N_13103,N_12674,N_12723);
xor U13104 (N_13104,N_12069,N_12979);
or U13105 (N_13105,N_12266,N_12374);
and U13106 (N_13106,N_12008,N_12694);
and U13107 (N_13107,N_12787,N_12122);
and U13108 (N_13108,N_12535,N_12705);
xor U13109 (N_13109,N_12301,N_12187);
or U13110 (N_13110,N_12778,N_12196);
xor U13111 (N_13111,N_12617,N_12025);
or U13112 (N_13112,N_12066,N_12300);
xor U13113 (N_13113,N_12158,N_12164);
nand U13114 (N_13114,N_12143,N_12819);
or U13115 (N_13115,N_12675,N_12009);
and U13116 (N_13116,N_12946,N_12472);
nor U13117 (N_13117,N_12628,N_12983);
nand U13118 (N_13118,N_12905,N_12450);
or U13119 (N_13119,N_12206,N_12210);
xor U13120 (N_13120,N_12888,N_12765);
xor U13121 (N_13121,N_12812,N_12860);
or U13122 (N_13122,N_12650,N_12126);
nand U13123 (N_13123,N_12963,N_12809);
nor U13124 (N_13124,N_12703,N_12077);
and U13125 (N_13125,N_12613,N_12800);
or U13126 (N_13126,N_12797,N_12129);
nand U13127 (N_13127,N_12565,N_12316);
nor U13128 (N_13128,N_12065,N_12590);
xnor U13129 (N_13129,N_12828,N_12977);
or U13130 (N_13130,N_12562,N_12397);
nor U13131 (N_13131,N_12404,N_12189);
or U13132 (N_13132,N_12067,N_12157);
nand U13133 (N_13133,N_12777,N_12339);
or U13134 (N_13134,N_12171,N_12792);
or U13135 (N_13135,N_12167,N_12998);
or U13136 (N_13136,N_12994,N_12479);
and U13137 (N_13137,N_12959,N_12023);
xnor U13138 (N_13138,N_12409,N_12183);
and U13139 (N_13139,N_12031,N_12774);
xnor U13140 (N_13140,N_12868,N_12995);
xor U13141 (N_13141,N_12991,N_12330);
nor U13142 (N_13142,N_12226,N_12292);
or U13143 (N_13143,N_12006,N_12485);
nand U13144 (N_13144,N_12721,N_12542);
or U13145 (N_13145,N_12458,N_12594);
or U13146 (N_13146,N_12970,N_12665);
or U13147 (N_13147,N_12089,N_12533);
nor U13148 (N_13148,N_12856,N_12754);
nand U13149 (N_13149,N_12854,N_12228);
nand U13150 (N_13150,N_12747,N_12264);
and U13151 (N_13151,N_12350,N_12356);
nor U13152 (N_13152,N_12021,N_12568);
xor U13153 (N_13153,N_12927,N_12470);
and U13154 (N_13154,N_12914,N_12035);
or U13155 (N_13155,N_12654,N_12578);
and U13156 (N_13156,N_12631,N_12247);
xnor U13157 (N_13157,N_12414,N_12907);
or U13158 (N_13158,N_12478,N_12463);
nand U13159 (N_13159,N_12596,N_12287);
or U13160 (N_13160,N_12996,N_12466);
xor U13161 (N_13161,N_12497,N_12492);
nor U13162 (N_13162,N_12880,N_12081);
xor U13163 (N_13163,N_12438,N_12637);
nand U13164 (N_13164,N_12191,N_12620);
or U13165 (N_13165,N_12636,N_12624);
and U13166 (N_13166,N_12986,N_12239);
and U13167 (N_13167,N_12050,N_12500);
or U13168 (N_13168,N_12720,N_12405);
and U13169 (N_13169,N_12769,N_12736);
xor U13170 (N_13170,N_12756,N_12135);
xnor U13171 (N_13171,N_12427,N_12846);
xnor U13172 (N_13172,N_12690,N_12583);
xor U13173 (N_13173,N_12253,N_12026);
or U13174 (N_13174,N_12839,N_12213);
and U13175 (N_13175,N_12722,N_12238);
or U13176 (N_13176,N_12311,N_12919);
and U13177 (N_13177,N_12668,N_12310);
or U13178 (N_13178,N_12468,N_12548);
nand U13179 (N_13179,N_12883,N_12731);
nor U13180 (N_13180,N_12547,N_12318);
xnor U13181 (N_13181,N_12585,N_12614);
xor U13182 (N_13182,N_12279,N_12399);
nand U13183 (N_13183,N_12847,N_12280);
nor U13184 (N_13184,N_12662,N_12948);
and U13185 (N_13185,N_12709,N_12477);
xnor U13186 (N_13186,N_12194,N_12530);
and U13187 (N_13187,N_12334,N_12420);
or U13188 (N_13188,N_12095,N_12153);
nand U13189 (N_13189,N_12402,N_12988);
nor U13190 (N_13190,N_12949,N_12967);
nor U13191 (N_13191,N_12704,N_12894);
nor U13192 (N_13192,N_12853,N_12743);
or U13193 (N_13193,N_12621,N_12212);
or U13194 (N_13194,N_12943,N_12116);
xor U13195 (N_13195,N_12322,N_12529);
or U13196 (N_13196,N_12702,N_12453);
and U13197 (N_13197,N_12040,N_12519);
nand U13198 (N_13198,N_12082,N_12048);
nor U13199 (N_13199,N_12767,N_12929);
and U13200 (N_13200,N_12293,N_12326);
or U13201 (N_13201,N_12681,N_12697);
nand U13202 (N_13202,N_12110,N_12298);
and U13203 (N_13203,N_12452,N_12312);
and U13204 (N_13204,N_12348,N_12999);
and U13205 (N_13205,N_12794,N_12749);
xor U13206 (N_13206,N_12252,N_12953);
nand U13207 (N_13207,N_12243,N_12971);
or U13208 (N_13208,N_12168,N_12276);
nor U13209 (N_13209,N_12160,N_12391);
nand U13210 (N_13210,N_12601,N_12735);
nor U13211 (N_13211,N_12528,N_12197);
nand U13212 (N_13212,N_12345,N_12807);
or U13213 (N_13213,N_12969,N_12917);
xnor U13214 (N_13214,N_12595,N_12421);
or U13215 (N_13215,N_12879,N_12430);
and U13216 (N_13216,N_12209,N_12344);
nor U13217 (N_13217,N_12314,N_12323);
nand U13218 (N_13218,N_12693,N_12683);
xor U13219 (N_13219,N_12549,N_12974);
nor U13220 (N_13220,N_12810,N_12866);
and U13221 (N_13221,N_12151,N_12052);
xor U13222 (N_13222,N_12096,N_12423);
xnor U13223 (N_13223,N_12329,N_12865);
xnor U13224 (N_13224,N_12891,N_12062);
nor U13225 (N_13225,N_12815,N_12071);
xnor U13226 (N_13226,N_12426,N_12726);
xor U13227 (N_13227,N_12455,N_12575);
or U13228 (N_13228,N_12139,N_12336);
nand U13229 (N_13229,N_12782,N_12643);
xor U13230 (N_13230,N_12718,N_12429);
nand U13231 (N_13231,N_12957,N_12555);
xor U13232 (N_13232,N_12406,N_12060);
or U13233 (N_13233,N_12149,N_12593);
nor U13234 (N_13234,N_12673,N_12771);
nand U13235 (N_13235,N_12250,N_12005);
nor U13236 (N_13236,N_12523,N_12014);
or U13237 (N_13237,N_12597,N_12371);
and U13238 (N_13238,N_12753,N_12010);
nand U13239 (N_13239,N_12878,N_12816);
nor U13240 (N_13240,N_12365,N_12521);
nand U13241 (N_13241,N_12190,N_12037);
nand U13242 (N_13242,N_12036,N_12283);
xor U13243 (N_13243,N_12304,N_12772);
or U13244 (N_13244,N_12054,N_12138);
xnor U13245 (N_13245,N_12083,N_12925);
nand U13246 (N_13246,N_12342,N_12688);
nand U13247 (N_13247,N_12012,N_12546);
nor U13248 (N_13248,N_12906,N_12443);
or U13249 (N_13249,N_12607,N_12978);
nand U13250 (N_13250,N_12958,N_12638);
nor U13251 (N_13251,N_12592,N_12539);
nor U13252 (N_13252,N_12394,N_12553);
nor U13253 (N_13253,N_12030,N_12056);
or U13254 (N_13254,N_12897,N_12428);
nand U13255 (N_13255,N_12352,N_12609);
and U13256 (N_13256,N_12512,N_12385);
xnor U13257 (N_13257,N_12677,N_12667);
or U13258 (N_13258,N_12813,N_12358);
and U13259 (N_13259,N_12090,N_12114);
nor U13260 (N_13260,N_12915,N_12413);
nand U13261 (N_13261,N_12013,N_12111);
or U13262 (N_13262,N_12554,N_12615);
nor U13263 (N_13263,N_12259,N_12381);
nor U13264 (N_13264,N_12488,N_12751);
xnor U13265 (N_13265,N_12989,N_12687);
or U13266 (N_13266,N_12502,N_12039);
nand U13267 (N_13267,N_12712,N_12019);
nor U13268 (N_13268,N_12713,N_12951);
and U13269 (N_13269,N_12962,N_12793);
xnor U13270 (N_13270,N_12170,N_12265);
and U13271 (N_13271,N_12034,N_12051);
nand U13272 (N_13272,N_12223,N_12824);
nor U13273 (N_13273,N_12835,N_12372);
nand U13274 (N_13274,N_12105,N_12145);
xnor U13275 (N_13275,N_12920,N_12942);
and U13276 (N_13276,N_12763,N_12327);
nand U13277 (N_13277,N_12269,N_12826);
nand U13278 (N_13278,N_12790,N_12563);
xnor U13279 (N_13279,N_12230,N_12805);
or U13280 (N_13280,N_12061,N_12150);
nor U13281 (N_13281,N_12146,N_12000);
xor U13282 (N_13282,N_12384,N_12425);
nor U13283 (N_13283,N_12284,N_12290);
or U13284 (N_13284,N_12263,N_12707);
or U13285 (N_13285,N_12830,N_12833);
nor U13286 (N_13286,N_12415,N_12627);
nor U13287 (N_13287,N_12701,N_12873);
xor U13288 (N_13288,N_12820,N_12537);
or U13289 (N_13289,N_12618,N_12085);
and U13290 (N_13290,N_12821,N_12002);
and U13291 (N_13291,N_12202,N_12435);
and U13292 (N_13292,N_12540,N_12748);
nor U13293 (N_13293,N_12863,N_12375);
and U13294 (N_13294,N_12018,N_12649);
and U13295 (N_13295,N_12109,N_12022);
nor U13296 (N_13296,N_12581,N_12987);
nand U13297 (N_13297,N_12755,N_12952);
xnor U13298 (N_13298,N_12606,N_12155);
or U13299 (N_13299,N_12678,N_12447);
and U13300 (N_13300,N_12660,N_12574);
nand U13301 (N_13301,N_12717,N_12604);
xnor U13302 (N_13302,N_12104,N_12779);
or U13303 (N_13303,N_12550,N_12525);
and U13304 (N_13304,N_12127,N_12680);
or U13305 (N_13305,N_12262,N_12236);
nand U13306 (N_13306,N_12134,N_12945);
nand U13307 (N_13307,N_12834,N_12305);
xnor U13308 (N_13308,N_12204,N_12538);
and U13309 (N_13309,N_12319,N_12128);
or U13310 (N_13310,N_12070,N_12564);
nand U13311 (N_13311,N_12392,N_12719);
nor U13312 (N_13312,N_12275,N_12029);
or U13313 (N_13313,N_12299,N_12584);
and U13314 (N_13314,N_12123,N_12598);
xnor U13315 (N_13315,N_12799,N_12007);
nor U13316 (N_13316,N_12669,N_12785);
xnor U13317 (N_13317,N_12446,N_12274);
or U13318 (N_13318,N_12981,N_12099);
nor U13319 (N_13319,N_12115,N_12295);
xor U13320 (N_13320,N_12032,N_12432);
nor U13321 (N_13321,N_12483,N_12656);
and U13322 (N_13322,N_12973,N_12395);
or U13323 (N_13323,N_12333,N_12179);
or U13324 (N_13324,N_12645,N_12520);
xnor U13325 (N_13325,N_12341,N_12623);
and U13326 (N_13326,N_12527,N_12534);
or U13327 (N_13327,N_12133,N_12362);
xnor U13328 (N_13328,N_12101,N_12335);
nor U13329 (N_13329,N_12806,N_12142);
nand U13330 (N_13330,N_12770,N_12396);
and U13331 (N_13331,N_12068,N_12734);
nand U13332 (N_13332,N_12510,N_12017);
xnor U13333 (N_13333,N_12364,N_12390);
nor U13334 (N_13334,N_12307,N_12867);
and U13335 (N_13335,N_12268,N_12216);
nor U13336 (N_13336,N_12490,N_12715);
nor U13337 (N_13337,N_12504,N_12175);
nor U13338 (N_13338,N_12208,N_12267);
and U13339 (N_13339,N_12120,N_12173);
and U13340 (N_13340,N_12761,N_12661);
nand U13341 (N_13341,N_12582,N_12439);
nor U13342 (N_13342,N_12784,N_12679);
nand U13343 (N_13343,N_12441,N_12639);
and U13344 (N_13344,N_12976,N_12078);
and U13345 (N_13345,N_12515,N_12671);
nand U13346 (N_13346,N_12728,N_12370);
nor U13347 (N_13347,N_12634,N_12232);
nor U13348 (N_13348,N_12184,N_12185);
and U13349 (N_13349,N_12112,N_12507);
or U13350 (N_13350,N_12526,N_12599);
xor U13351 (N_13351,N_12169,N_12076);
nor U13352 (N_13352,N_12804,N_12935);
or U13353 (N_13353,N_12075,N_12795);
and U13354 (N_13354,N_12476,N_12353);
and U13355 (N_13355,N_12576,N_12303);
and U13356 (N_13356,N_12147,N_12727);
nand U13357 (N_13357,N_12367,N_12561);
or U13358 (N_13358,N_12162,N_12874);
and U13359 (N_13359,N_12750,N_12055);
or U13360 (N_13360,N_12700,N_12895);
nand U13361 (N_13361,N_12254,N_12498);
nor U13362 (N_13362,N_12982,N_12921);
nor U13363 (N_13363,N_12802,N_12359);
nor U13364 (N_13364,N_12296,N_12933);
and U13365 (N_13365,N_12985,N_12195);
nand U13366 (N_13366,N_12046,N_12516);
nand U13367 (N_13367,N_12419,N_12460);
or U13368 (N_13368,N_12912,N_12648);
nand U13369 (N_13369,N_12602,N_12655);
nor U13370 (N_13370,N_12380,N_12928);
nand U13371 (N_13371,N_12798,N_12182);
xnor U13372 (N_13372,N_12831,N_12433);
nand U13373 (N_13373,N_12418,N_12107);
and U13374 (N_13374,N_12560,N_12474);
xnor U13375 (N_13375,N_12461,N_12225);
nor U13376 (N_13376,N_12786,N_12059);
and U13377 (N_13377,N_12698,N_12566);
and U13378 (N_13378,N_12401,N_12870);
nor U13379 (N_13379,N_12108,N_12424);
or U13380 (N_13380,N_12467,N_12422);
nor U13381 (N_13381,N_12541,N_12930);
xnor U13382 (N_13382,N_12289,N_12522);
nor U13383 (N_13383,N_12382,N_12448);
and U13384 (N_13384,N_12496,N_12369);
xnor U13385 (N_13385,N_12049,N_12355);
nor U13386 (N_13386,N_12993,N_12557);
nor U13387 (N_13387,N_12317,N_12245);
nor U13388 (N_13388,N_12551,N_12106);
xnor U13389 (N_13389,N_12543,N_12237);
xor U13390 (N_13390,N_12509,N_12093);
or U13391 (N_13391,N_12659,N_12403);
xor U13392 (N_13392,N_12901,N_12964);
xor U13393 (N_13393,N_12349,N_12822);
nand U13394 (N_13394,N_12633,N_12291);
or U13395 (N_13395,N_12469,N_12297);
nor U13396 (N_13396,N_12224,N_12732);
xnor U13397 (N_13397,N_12545,N_12306);
or U13398 (N_13398,N_12695,N_12589);
and U13399 (N_13399,N_12682,N_12063);
and U13400 (N_13400,N_12760,N_12347);
and U13401 (N_13401,N_12091,N_12449);
or U13402 (N_13402,N_12725,N_12440);
and U13403 (N_13403,N_12980,N_12651);
and U13404 (N_13404,N_12908,N_12136);
nor U13405 (N_13405,N_12144,N_12222);
nor U13406 (N_13406,N_12629,N_12603);
nand U13407 (N_13407,N_12015,N_12569);
and U13408 (N_13408,N_12893,N_12271);
nor U13409 (N_13409,N_12505,N_12346);
and U13410 (N_13410,N_12781,N_12220);
xor U13411 (N_13411,N_12176,N_12309);
nor U13412 (N_13412,N_12495,N_12737);
nand U13413 (N_13413,N_12610,N_12689);
xnor U13414 (N_13414,N_12064,N_12872);
xor U13415 (N_13415,N_12814,N_12328);
nor U13416 (N_13416,N_12859,N_12456);
nor U13417 (N_13417,N_12903,N_12902);
and U13418 (N_13418,N_12486,N_12073);
or U13419 (N_13419,N_12188,N_12215);
or U13420 (N_13420,N_12379,N_12823);
xnor U13421 (N_13421,N_12011,N_12482);
or U13422 (N_13422,N_12140,N_12892);
or U13423 (N_13423,N_12199,N_12387);
and U13424 (N_13424,N_12100,N_12841);
xnor U13425 (N_13425,N_12818,N_12332);
nand U13426 (N_13426,N_12780,N_12057);
and U13427 (N_13427,N_12272,N_12622);
or U13428 (N_13428,N_12084,N_12261);
nor U13429 (N_13429,N_12255,N_12027);
nand U13430 (N_13430,N_12313,N_12240);
and U13431 (N_13431,N_12118,N_12235);
xnor U13432 (N_13432,N_12811,N_12875);
and U13433 (N_13433,N_12431,N_12926);
or U13434 (N_13434,N_12900,N_12088);
xnor U13435 (N_13435,N_12410,N_12416);
nor U13436 (N_13436,N_12487,N_12864);
and U13437 (N_13437,N_12320,N_12473);
nand U13438 (N_13438,N_12745,N_12163);
and U13439 (N_13439,N_12366,N_12174);
or U13440 (N_13440,N_12400,N_12672);
or U13441 (N_13441,N_12849,N_12211);
nor U13442 (N_13442,N_12270,N_12233);
xor U13443 (N_13443,N_12434,N_12234);
xor U13444 (N_13444,N_12508,N_12363);
nand U13445 (N_13445,N_12947,N_12033);
nand U13446 (N_13446,N_12045,N_12436);
nand U13447 (N_13447,N_12647,N_12102);
or U13448 (N_13448,N_12351,N_12041);
nor U13449 (N_13449,N_12716,N_12325);
nor U13450 (N_13450,N_12462,N_12331);
or U13451 (N_13451,N_12518,N_12916);
nor U13452 (N_13452,N_12739,N_12844);
or U13453 (N_13453,N_12644,N_12437);
or U13454 (N_13454,N_12181,N_12471);
or U13455 (N_13455,N_12020,N_12862);
or U13456 (N_13456,N_12340,N_12417);
nand U13457 (N_13457,N_12357,N_12131);
nand U13458 (N_13458,N_12042,N_12412);
and U13459 (N_13459,N_12944,N_12954);
xnor U13460 (N_13460,N_12931,N_12758);
xnor U13461 (N_13461,N_12729,N_12038);
or U13462 (N_13462,N_12464,N_12764);
or U13463 (N_13463,N_12586,N_12837);
and U13464 (N_13464,N_12836,N_12827);
or U13465 (N_13465,N_12630,N_12536);
nand U13466 (N_13466,N_12936,N_12699);
and U13467 (N_13467,N_12882,N_12840);
nand U13468 (N_13468,N_12080,N_12658);
xor U13469 (N_13469,N_12884,N_12960);
and U13470 (N_13470,N_12229,N_12646);
nor U13471 (N_13471,N_12484,N_12273);
xor U13472 (N_13472,N_12378,N_12899);
and U13473 (N_13473,N_12087,N_12965);
nor U13474 (N_13474,N_12752,N_12966);
nor U13475 (N_13475,N_12368,N_12354);
nor U13476 (N_13476,N_12600,N_12898);
xnor U13477 (N_13477,N_12513,N_12922);
xnor U13478 (N_13478,N_12911,N_12762);
and U13479 (N_13479,N_12796,N_12489);
nor U13480 (N_13480,N_12376,N_12937);
xor U13481 (N_13481,N_12338,N_12567);
xnor U13482 (N_13482,N_12738,N_12302);
nor U13483 (N_13483,N_12642,N_12024);
nand U13484 (N_13484,N_12246,N_12803);
and U13485 (N_13485,N_12591,N_12214);
and U13486 (N_13486,N_12141,N_12972);
nand U13487 (N_13487,N_12186,N_12775);
nand U13488 (N_13488,N_12103,N_12241);
and U13489 (N_13489,N_12791,N_12047);
xor U13490 (N_13490,N_12587,N_12221);
nor U13491 (N_13491,N_12288,N_12227);
xor U13492 (N_13492,N_12154,N_12125);
and U13493 (N_13493,N_12744,N_12961);
or U13494 (N_13494,N_12910,N_12579);
or U13495 (N_13495,N_12532,N_12676);
nand U13496 (N_13496,N_12166,N_12653);
or U13497 (N_13497,N_12480,N_12871);
xor U13498 (N_13498,N_12852,N_12285);
nor U13499 (N_13499,N_12626,N_12706);
nand U13500 (N_13500,N_12336,N_12207);
nand U13501 (N_13501,N_12594,N_12643);
nor U13502 (N_13502,N_12894,N_12264);
nand U13503 (N_13503,N_12303,N_12082);
or U13504 (N_13504,N_12663,N_12091);
and U13505 (N_13505,N_12581,N_12656);
nor U13506 (N_13506,N_12780,N_12838);
nor U13507 (N_13507,N_12542,N_12733);
nand U13508 (N_13508,N_12580,N_12863);
or U13509 (N_13509,N_12818,N_12117);
and U13510 (N_13510,N_12539,N_12525);
xor U13511 (N_13511,N_12993,N_12947);
nand U13512 (N_13512,N_12106,N_12148);
nor U13513 (N_13513,N_12429,N_12410);
nand U13514 (N_13514,N_12241,N_12601);
nand U13515 (N_13515,N_12066,N_12950);
nand U13516 (N_13516,N_12952,N_12672);
nor U13517 (N_13517,N_12457,N_12551);
nor U13518 (N_13518,N_12870,N_12210);
or U13519 (N_13519,N_12512,N_12685);
nand U13520 (N_13520,N_12300,N_12732);
and U13521 (N_13521,N_12374,N_12768);
and U13522 (N_13522,N_12438,N_12897);
nor U13523 (N_13523,N_12824,N_12615);
xor U13524 (N_13524,N_12600,N_12554);
and U13525 (N_13525,N_12223,N_12422);
xnor U13526 (N_13526,N_12348,N_12544);
xor U13527 (N_13527,N_12461,N_12628);
nand U13528 (N_13528,N_12393,N_12846);
xnor U13529 (N_13529,N_12925,N_12033);
nor U13530 (N_13530,N_12889,N_12801);
nand U13531 (N_13531,N_12450,N_12029);
and U13532 (N_13532,N_12670,N_12706);
or U13533 (N_13533,N_12127,N_12504);
or U13534 (N_13534,N_12973,N_12058);
nor U13535 (N_13535,N_12145,N_12362);
and U13536 (N_13536,N_12404,N_12346);
nand U13537 (N_13537,N_12618,N_12398);
nand U13538 (N_13538,N_12435,N_12495);
xnor U13539 (N_13539,N_12476,N_12551);
and U13540 (N_13540,N_12980,N_12217);
or U13541 (N_13541,N_12641,N_12440);
or U13542 (N_13542,N_12745,N_12336);
nand U13543 (N_13543,N_12733,N_12201);
and U13544 (N_13544,N_12903,N_12895);
or U13545 (N_13545,N_12139,N_12355);
and U13546 (N_13546,N_12692,N_12286);
or U13547 (N_13547,N_12771,N_12146);
or U13548 (N_13548,N_12608,N_12311);
nor U13549 (N_13549,N_12216,N_12112);
and U13550 (N_13550,N_12469,N_12474);
or U13551 (N_13551,N_12807,N_12276);
nand U13552 (N_13552,N_12903,N_12241);
nand U13553 (N_13553,N_12258,N_12665);
xor U13554 (N_13554,N_12883,N_12980);
or U13555 (N_13555,N_12950,N_12618);
xor U13556 (N_13556,N_12017,N_12189);
nand U13557 (N_13557,N_12937,N_12962);
nand U13558 (N_13558,N_12965,N_12720);
xnor U13559 (N_13559,N_12040,N_12714);
and U13560 (N_13560,N_12669,N_12118);
and U13561 (N_13561,N_12250,N_12661);
nand U13562 (N_13562,N_12154,N_12972);
nand U13563 (N_13563,N_12191,N_12728);
nor U13564 (N_13564,N_12207,N_12384);
or U13565 (N_13565,N_12579,N_12529);
nor U13566 (N_13566,N_12310,N_12467);
and U13567 (N_13567,N_12544,N_12909);
or U13568 (N_13568,N_12647,N_12756);
nor U13569 (N_13569,N_12821,N_12705);
and U13570 (N_13570,N_12222,N_12428);
xnor U13571 (N_13571,N_12621,N_12784);
or U13572 (N_13572,N_12968,N_12301);
nor U13573 (N_13573,N_12633,N_12823);
nor U13574 (N_13574,N_12941,N_12661);
or U13575 (N_13575,N_12950,N_12814);
and U13576 (N_13576,N_12140,N_12213);
and U13577 (N_13577,N_12682,N_12851);
nor U13578 (N_13578,N_12878,N_12849);
or U13579 (N_13579,N_12468,N_12074);
or U13580 (N_13580,N_12347,N_12264);
nor U13581 (N_13581,N_12860,N_12434);
and U13582 (N_13582,N_12442,N_12076);
nor U13583 (N_13583,N_12106,N_12241);
or U13584 (N_13584,N_12701,N_12656);
or U13585 (N_13585,N_12614,N_12845);
or U13586 (N_13586,N_12363,N_12010);
xnor U13587 (N_13587,N_12843,N_12870);
xnor U13588 (N_13588,N_12457,N_12317);
xnor U13589 (N_13589,N_12463,N_12602);
and U13590 (N_13590,N_12685,N_12304);
nor U13591 (N_13591,N_12346,N_12977);
xor U13592 (N_13592,N_12219,N_12467);
nor U13593 (N_13593,N_12568,N_12163);
nand U13594 (N_13594,N_12706,N_12068);
and U13595 (N_13595,N_12705,N_12269);
or U13596 (N_13596,N_12825,N_12025);
nor U13597 (N_13597,N_12187,N_12275);
or U13598 (N_13598,N_12662,N_12927);
nand U13599 (N_13599,N_12599,N_12717);
xor U13600 (N_13600,N_12581,N_12354);
and U13601 (N_13601,N_12280,N_12145);
nand U13602 (N_13602,N_12393,N_12570);
or U13603 (N_13603,N_12824,N_12716);
or U13604 (N_13604,N_12527,N_12656);
nand U13605 (N_13605,N_12697,N_12433);
nor U13606 (N_13606,N_12822,N_12175);
xnor U13607 (N_13607,N_12513,N_12772);
and U13608 (N_13608,N_12842,N_12097);
and U13609 (N_13609,N_12170,N_12809);
xor U13610 (N_13610,N_12391,N_12485);
or U13611 (N_13611,N_12916,N_12567);
xor U13612 (N_13612,N_12276,N_12783);
nand U13613 (N_13613,N_12501,N_12567);
or U13614 (N_13614,N_12085,N_12197);
and U13615 (N_13615,N_12657,N_12204);
or U13616 (N_13616,N_12154,N_12047);
xnor U13617 (N_13617,N_12491,N_12174);
xnor U13618 (N_13618,N_12521,N_12001);
nand U13619 (N_13619,N_12691,N_12141);
or U13620 (N_13620,N_12139,N_12553);
and U13621 (N_13621,N_12205,N_12662);
nor U13622 (N_13622,N_12480,N_12178);
xor U13623 (N_13623,N_12700,N_12996);
nor U13624 (N_13624,N_12205,N_12830);
or U13625 (N_13625,N_12977,N_12095);
nand U13626 (N_13626,N_12025,N_12501);
nand U13627 (N_13627,N_12317,N_12424);
nand U13628 (N_13628,N_12780,N_12295);
and U13629 (N_13629,N_12106,N_12515);
or U13630 (N_13630,N_12366,N_12790);
xnor U13631 (N_13631,N_12066,N_12170);
nand U13632 (N_13632,N_12031,N_12132);
or U13633 (N_13633,N_12550,N_12206);
and U13634 (N_13634,N_12519,N_12500);
or U13635 (N_13635,N_12634,N_12863);
nand U13636 (N_13636,N_12837,N_12526);
nor U13637 (N_13637,N_12536,N_12620);
nor U13638 (N_13638,N_12977,N_12581);
or U13639 (N_13639,N_12542,N_12992);
nor U13640 (N_13640,N_12391,N_12948);
xor U13641 (N_13641,N_12777,N_12095);
and U13642 (N_13642,N_12275,N_12039);
nor U13643 (N_13643,N_12587,N_12785);
nor U13644 (N_13644,N_12161,N_12827);
nor U13645 (N_13645,N_12748,N_12769);
nor U13646 (N_13646,N_12290,N_12878);
nor U13647 (N_13647,N_12356,N_12065);
and U13648 (N_13648,N_12240,N_12886);
nor U13649 (N_13649,N_12915,N_12383);
and U13650 (N_13650,N_12601,N_12701);
and U13651 (N_13651,N_12024,N_12508);
or U13652 (N_13652,N_12896,N_12234);
nand U13653 (N_13653,N_12574,N_12263);
and U13654 (N_13654,N_12427,N_12880);
and U13655 (N_13655,N_12474,N_12310);
xnor U13656 (N_13656,N_12631,N_12260);
nor U13657 (N_13657,N_12551,N_12728);
and U13658 (N_13658,N_12312,N_12711);
nand U13659 (N_13659,N_12918,N_12170);
and U13660 (N_13660,N_12174,N_12868);
nand U13661 (N_13661,N_12836,N_12365);
and U13662 (N_13662,N_12641,N_12889);
xnor U13663 (N_13663,N_12092,N_12004);
nand U13664 (N_13664,N_12307,N_12798);
and U13665 (N_13665,N_12228,N_12445);
nand U13666 (N_13666,N_12670,N_12732);
or U13667 (N_13667,N_12231,N_12485);
or U13668 (N_13668,N_12215,N_12368);
xor U13669 (N_13669,N_12873,N_12397);
nor U13670 (N_13670,N_12703,N_12920);
nor U13671 (N_13671,N_12461,N_12458);
and U13672 (N_13672,N_12707,N_12814);
xor U13673 (N_13673,N_12291,N_12287);
nand U13674 (N_13674,N_12430,N_12415);
nand U13675 (N_13675,N_12284,N_12336);
nor U13676 (N_13676,N_12156,N_12221);
nor U13677 (N_13677,N_12752,N_12516);
and U13678 (N_13678,N_12709,N_12612);
and U13679 (N_13679,N_12451,N_12683);
or U13680 (N_13680,N_12299,N_12853);
nand U13681 (N_13681,N_12773,N_12867);
and U13682 (N_13682,N_12901,N_12302);
nor U13683 (N_13683,N_12068,N_12069);
or U13684 (N_13684,N_12088,N_12292);
nand U13685 (N_13685,N_12391,N_12557);
nor U13686 (N_13686,N_12696,N_12447);
nor U13687 (N_13687,N_12224,N_12534);
nand U13688 (N_13688,N_12128,N_12284);
nand U13689 (N_13689,N_12991,N_12829);
xnor U13690 (N_13690,N_12248,N_12111);
xnor U13691 (N_13691,N_12897,N_12284);
nand U13692 (N_13692,N_12484,N_12735);
xor U13693 (N_13693,N_12007,N_12157);
xnor U13694 (N_13694,N_12457,N_12640);
or U13695 (N_13695,N_12893,N_12277);
xnor U13696 (N_13696,N_12283,N_12185);
or U13697 (N_13697,N_12205,N_12988);
or U13698 (N_13698,N_12378,N_12598);
nand U13699 (N_13699,N_12727,N_12529);
or U13700 (N_13700,N_12606,N_12075);
nand U13701 (N_13701,N_12651,N_12187);
and U13702 (N_13702,N_12605,N_12667);
and U13703 (N_13703,N_12043,N_12032);
nand U13704 (N_13704,N_12107,N_12714);
or U13705 (N_13705,N_12171,N_12681);
or U13706 (N_13706,N_12783,N_12675);
or U13707 (N_13707,N_12457,N_12132);
nor U13708 (N_13708,N_12829,N_12261);
and U13709 (N_13709,N_12163,N_12682);
nor U13710 (N_13710,N_12462,N_12352);
xor U13711 (N_13711,N_12675,N_12296);
or U13712 (N_13712,N_12912,N_12504);
or U13713 (N_13713,N_12464,N_12783);
and U13714 (N_13714,N_12405,N_12589);
xnor U13715 (N_13715,N_12938,N_12517);
nor U13716 (N_13716,N_12649,N_12212);
and U13717 (N_13717,N_12929,N_12224);
or U13718 (N_13718,N_12161,N_12067);
nand U13719 (N_13719,N_12874,N_12305);
nor U13720 (N_13720,N_12698,N_12089);
and U13721 (N_13721,N_12304,N_12956);
or U13722 (N_13722,N_12377,N_12384);
or U13723 (N_13723,N_12060,N_12942);
and U13724 (N_13724,N_12890,N_12152);
nand U13725 (N_13725,N_12453,N_12128);
or U13726 (N_13726,N_12223,N_12075);
nand U13727 (N_13727,N_12736,N_12069);
nand U13728 (N_13728,N_12327,N_12002);
nand U13729 (N_13729,N_12438,N_12851);
or U13730 (N_13730,N_12096,N_12931);
nor U13731 (N_13731,N_12500,N_12752);
nor U13732 (N_13732,N_12345,N_12556);
nor U13733 (N_13733,N_12743,N_12182);
nor U13734 (N_13734,N_12644,N_12471);
or U13735 (N_13735,N_12139,N_12985);
nand U13736 (N_13736,N_12281,N_12180);
nand U13737 (N_13737,N_12341,N_12040);
xnor U13738 (N_13738,N_12340,N_12347);
and U13739 (N_13739,N_12264,N_12616);
nor U13740 (N_13740,N_12042,N_12325);
nor U13741 (N_13741,N_12833,N_12590);
nand U13742 (N_13742,N_12781,N_12493);
nand U13743 (N_13743,N_12242,N_12321);
xor U13744 (N_13744,N_12673,N_12295);
nand U13745 (N_13745,N_12870,N_12262);
xor U13746 (N_13746,N_12815,N_12554);
nor U13747 (N_13747,N_12041,N_12583);
xnor U13748 (N_13748,N_12114,N_12942);
or U13749 (N_13749,N_12635,N_12106);
and U13750 (N_13750,N_12321,N_12964);
or U13751 (N_13751,N_12085,N_12425);
xnor U13752 (N_13752,N_12222,N_12830);
nand U13753 (N_13753,N_12399,N_12689);
or U13754 (N_13754,N_12129,N_12096);
xor U13755 (N_13755,N_12817,N_12803);
or U13756 (N_13756,N_12969,N_12299);
nor U13757 (N_13757,N_12870,N_12827);
nor U13758 (N_13758,N_12227,N_12037);
nor U13759 (N_13759,N_12664,N_12831);
xnor U13760 (N_13760,N_12215,N_12941);
and U13761 (N_13761,N_12150,N_12906);
xnor U13762 (N_13762,N_12947,N_12749);
or U13763 (N_13763,N_12945,N_12489);
or U13764 (N_13764,N_12343,N_12612);
or U13765 (N_13765,N_12086,N_12435);
nor U13766 (N_13766,N_12834,N_12243);
and U13767 (N_13767,N_12183,N_12164);
nand U13768 (N_13768,N_12277,N_12711);
or U13769 (N_13769,N_12686,N_12040);
nand U13770 (N_13770,N_12529,N_12849);
nand U13771 (N_13771,N_12204,N_12404);
xor U13772 (N_13772,N_12079,N_12510);
and U13773 (N_13773,N_12161,N_12352);
nand U13774 (N_13774,N_12349,N_12803);
or U13775 (N_13775,N_12495,N_12674);
or U13776 (N_13776,N_12125,N_12269);
or U13777 (N_13777,N_12687,N_12779);
nor U13778 (N_13778,N_12951,N_12529);
and U13779 (N_13779,N_12149,N_12789);
or U13780 (N_13780,N_12743,N_12204);
nor U13781 (N_13781,N_12401,N_12550);
nor U13782 (N_13782,N_12251,N_12702);
xor U13783 (N_13783,N_12803,N_12464);
xnor U13784 (N_13784,N_12056,N_12415);
xor U13785 (N_13785,N_12657,N_12757);
nor U13786 (N_13786,N_12697,N_12872);
nand U13787 (N_13787,N_12969,N_12133);
and U13788 (N_13788,N_12467,N_12843);
xor U13789 (N_13789,N_12105,N_12359);
xnor U13790 (N_13790,N_12907,N_12458);
or U13791 (N_13791,N_12861,N_12225);
and U13792 (N_13792,N_12476,N_12793);
and U13793 (N_13793,N_12147,N_12100);
nor U13794 (N_13794,N_12989,N_12666);
nor U13795 (N_13795,N_12453,N_12580);
xnor U13796 (N_13796,N_12327,N_12004);
or U13797 (N_13797,N_12376,N_12690);
xor U13798 (N_13798,N_12467,N_12804);
nand U13799 (N_13799,N_12429,N_12206);
xnor U13800 (N_13800,N_12518,N_12907);
nand U13801 (N_13801,N_12934,N_12167);
nor U13802 (N_13802,N_12289,N_12388);
or U13803 (N_13803,N_12143,N_12368);
or U13804 (N_13804,N_12549,N_12687);
or U13805 (N_13805,N_12380,N_12995);
or U13806 (N_13806,N_12753,N_12136);
xor U13807 (N_13807,N_12427,N_12082);
nand U13808 (N_13808,N_12516,N_12059);
or U13809 (N_13809,N_12489,N_12532);
or U13810 (N_13810,N_12960,N_12977);
nor U13811 (N_13811,N_12450,N_12955);
nor U13812 (N_13812,N_12361,N_12075);
nand U13813 (N_13813,N_12689,N_12528);
nand U13814 (N_13814,N_12096,N_12473);
and U13815 (N_13815,N_12378,N_12307);
and U13816 (N_13816,N_12425,N_12120);
or U13817 (N_13817,N_12458,N_12766);
nor U13818 (N_13818,N_12401,N_12572);
and U13819 (N_13819,N_12498,N_12748);
and U13820 (N_13820,N_12991,N_12758);
and U13821 (N_13821,N_12433,N_12175);
or U13822 (N_13822,N_12392,N_12367);
and U13823 (N_13823,N_12320,N_12635);
or U13824 (N_13824,N_12662,N_12321);
and U13825 (N_13825,N_12854,N_12495);
nor U13826 (N_13826,N_12583,N_12375);
and U13827 (N_13827,N_12223,N_12387);
nand U13828 (N_13828,N_12440,N_12881);
or U13829 (N_13829,N_12377,N_12717);
xor U13830 (N_13830,N_12390,N_12208);
nand U13831 (N_13831,N_12122,N_12248);
and U13832 (N_13832,N_12666,N_12003);
or U13833 (N_13833,N_12496,N_12046);
nand U13834 (N_13834,N_12255,N_12522);
and U13835 (N_13835,N_12734,N_12852);
and U13836 (N_13836,N_12847,N_12732);
xnor U13837 (N_13837,N_12751,N_12219);
or U13838 (N_13838,N_12668,N_12047);
nand U13839 (N_13839,N_12634,N_12213);
nand U13840 (N_13840,N_12375,N_12511);
xor U13841 (N_13841,N_12392,N_12755);
nor U13842 (N_13842,N_12297,N_12531);
xor U13843 (N_13843,N_12362,N_12661);
or U13844 (N_13844,N_12717,N_12041);
or U13845 (N_13845,N_12170,N_12542);
nand U13846 (N_13846,N_12466,N_12037);
nand U13847 (N_13847,N_12911,N_12443);
and U13848 (N_13848,N_12692,N_12117);
and U13849 (N_13849,N_12585,N_12112);
nor U13850 (N_13850,N_12502,N_12585);
or U13851 (N_13851,N_12017,N_12119);
nor U13852 (N_13852,N_12269,N_12846);
or U13853 (N_13853,N_12790,N_12150);
nand U13854 (N_13854,N_12811,N_12490);
nor U13855 (N_13855,N_12364,N_12702);
nand U13856 (N_13856,N_12940,N_12480);
nand U13857 (N_13857,N_12559,N_12131);
xor U13858 (N_13858,N_12639,N_12736);
and U13859 (N_13859,N_12029,N_12080);
and U13860 (N_13860,N_12864,N_12827);
nor U13861 (N_13861,N_12194,N_12381);
or U13862 (N_13862,N_12321,N_12061);
nor U13863 (N_13863,N_12623,N_12904);
nand U13864 (N_13864,N_12371,N_12134);
nand U13865 (N_13865,N_12715,N_12191);
and U13866 (N_13866,N_12754,N_12052);
nand U13867 (N_13867,N_12102,N_12151);
xnor U13868 (N_13868,N_12308,N_12482);
and U13869 (N_13869,N_12435,N_12563);
nand U13870 (N_13870,N_12741,N_12996);
or U13871 (N_13871,N_12470,N_12037);
xnor U13872 (N_13872,N_12580,N_12488);
or U13873 (N_13873,N_12643,N_12813);
xnor U13874 (N_13874,N_12104,N_12484);
nand U13875 (N_13875,N_12101,N_12546);
nand U13876 (N_13876,N_12976,N_12846);
xor U13877 (N_13877,N_12743,N_12096);
or U13878 (N_13878,N_12862,N_12402);
nand U13879 (N_13879,N_12066,N_12738);
xnor U13880 (N_13880,N_12812,N_12006);
xor U13881 (N_13881,N_12559,N_12777);
and U13882 (N_13882,N_12728,N_12762);
xor U13883 (N_13883,N_12098,N_12240);
xnor U13884 (N_13884,N_12667,N_12898);
or U13885 (N_13885,N_12645,N_12430);
xor U13886 (N_13886,N_12156,N_12121);
xnor U13887 (N_13887,N_12977,N_12670);
nand U13888 (N_13888,N_12982,N_12457);
nand U13889 (N_13889,N_12931,N_12940);
and U13890 (N_13890,N_12878,N_12799);
nand U13891 (N_13891,N_12169,N_12155);
xor U13892 (N_13892,N_12345,N_12056);
or U13893 (N_13893,N_12566,N_12689);
nand U13894 (N_13894,N_12901,N_12096);
nand U13895 (N_13895,N_12468,N_12414);
nor U13896 (N_13896,N_12486,N_12005);
and U13897 (N_13897,N_12292,N_12825);
or U13898 (N_13898,N_12016,N_12775);
and U13899 (N_13899,N_12054,N_12815);
nor U13900 (N_13900,N_12229,N_12636);
nor U13901 (N_13901,N_12727,N_12687);
nand U13902 (N_13902,N_12984,N_12654);
or U13903 (N_13903,N_12765,N_12253);
nor U13904 (N_13904,N_12769,N_12604);
xnor U13905 (N_13905,N_12471,N_12797);
nand U13906 (N_13906,N_12954,N_12432);
xnor U13907 (N_13907,N_12046,N_12359);
xnor U13908 (N_13908,N_12751,N_12871);
nor U13909 (N_13909,N_12294,N_12132);
and U13910 (N_13910,N_12915,N_12328);
and U13911 (N_13911,N_12002,N_12981);
or U13912 (N_13912,N_12732,N_12931);
nor U13913 (N_13913,N_12132,N_12000);
or U13914 (N_13914,N_12748,N_12131);
nor U13915 (N_13915,N_12624,N_12716);
and U13916 (N_13916,N_12741,N_12217);
nand U13917 (N_13917,N_12854,N_12394);
or U13918 (N_13918,N_12520,N_12942);
nor U13919 (N_13919,N_12193,N_12972);
and U13920 (N_13920,N_12358,N_12779);
and U13921 (N_13921,N_12109,N_12529);
nand U13922 (N_13922,N_12665,N_12038);
nor U13923 (N_13923,N_12313,N_12707);
xor U13924 (N_13924,N_12587,N_12095);
xor U13925 (N_13925,N_12842,N_12550);
nor U13926 (N_13926,N_12475,N_12685);
nand U13927 (N_13927,N_12341,N_12694);
or U13928 (N_13928,N_12572,N_12735);
or U13929 (N_13929,N_12756,N_12855);
xnor U13930 (N_13930,N_12967,N_12471);
or U13931 (N_13931,N_12867,N_12019);
nand U13932 (N_13932,N_12510,N_12529);
or U13933 (N_13933,N_12490,N_12035);
or U13934 (N_13934,N_12339,N_12151);
nand U13935 (N_13935,N_12039,N_12949);
or U13936 (N_13936,N_12266,N_12021);
nor U13937 (N_13937,N_12561,N_12251);
or U13938 (N_13938,N_12166,N_12349);
and U13939 (N_13939,N_12131,N_12990);
and U13940 (N_13940,N_12027,N_12381);
xnor U13941 (N_13941,N_12175,N_12036);
or U13942 (N_13942,N_12340,N_12645);
or U13943 (N_13943,N_12431,N_12477);
nand U13944 (N_13944,N_12471,N_12113);
and U13945 (N_13945,N_12615,N_12355);
xnor U13946 (N_13946,N_12118,N_12786);
xor U13947 (N_13947,N_12910,N_12667);
or U13948 (N_13948,N_12289,N_12818);
and U13949 (N_13949,N_12852,N_12963);
xnor U13950 (N_13950,N_12464,N_12496);
and U13951 (N_13951,N_12277,N_12854);
nor U13952 (N_13952,N_12276,N_12235);
or U13953 (N_13953,N_12695,N_12160);
nor U13954 (N_13954,N_12548,N_12015);
or U13955 (N_13955,N_12249,N_12457);
and U13956 (N_13956,N_12429,N_12734);
nand U13957 (N_13957,N_12209,N_12695);
nor U13958 (N_13958,N_12317,N_12462);
and U13959 (N_13959,N_12027,N_12701);
and U13960 (N_13960,N_12300,N_12465);
and U13961 (N_13961,N_12261,N_12872);
nand U13962 (N_13962,N_12031,N_12040);
nor U13963 (N_13963,N_12262,N_12146);
nor U13964 (N_13964,N_12094,N_12836);
nor U13965 (N_13965,N_12946,N_12018);
and U13966 (N_13966,N_12978,N_12660);
xnor U13967 (N_13967,N_12120,N_12489);
xnor U13968 (N_13968,N_12353,N_12502);
nor U13969 (N_13969,N_12034,N_12618);
nand U13970 (N_13970,N_12419,N_12113);
nand U13971 (N_13971,N_12852,N_12443);
and U13972 (N_13972,N_12951,N_12543);
or U13973 (N_13973,N_12079,N_12937);
xor U13974 (N_13974,N_12887,N_12898);
nand U13975 (N_13975,N_12950,N_12704);
or U13976 (N_13976,N_12090,N_12531);
nor U13977 (N_13977,N_12516,N_12480);
or U13978 (N_13978,N_12617,N_12260);
or U13979 (N_13979,N_12791,N_12114);
and U13980 (N_13980,N_12814,N_12622);
nand U13981 (N_13981,N_12576,N_12359);
nand U13982 (N_13982,N_12948,N_12281);
and U13983 (N_13983,N_12219,N_12616);
or U13984 (N_13984,N_12140,N_12956);
xor U13985 (N_13985,N_12094,N_12948);
xor U13986 (N_13986,N_12895,N_12393);
nor U13987 (N_13987,N_12769,N_12199);
nor U13988 (N_13988,N_12510,N_12968);
nor U13989 (N_13989,N_12593,N_12673);
xor U13990 (N_13990,N_12139,N_12724);
and U13991 (N_13991,N_12099,N_12610);
xnor U13992 (N_13992,N_12223,N_12955);
and U13993 (N_13993,N_12509,N_12100);
and U13994 (N_13994,N_12166,N_12022);
or U13995 (N_13995,N_12411,N_12679);
xnor U13996 (N_13996,N_12359,N_12317);
nand U13997 (N_13997,N_12433,N_12011);
and U13998 (N_13998,N_12746,N_12227);
and U13999 (N_13999,N_12514,N_12543);
or U14000 (N_14000,N_13875,N_13640);
or U14001 (N_14001,N_13506,N_13386);
and U14002 (N_14002,N_13300,N_13568);
or U14003 (N_14003,N_13317,N_13566);
nand U14004 (N_14004,N_13809,N_13078);
and U14005 (N_14005,N_13426,N_13036);
xnor U14006 (N_14006,N_13969,N_13354);
nor U14007 (N_14007,N_13112,N_13655);
xnor U14008 (N_14008,N_13251,N_13684);
nor U14009 (N_14009,N_13819,N_13323);
xor U14010 (N_14010,N_13126,N_13547);
nor U14011 (N_14011,N_13401,N_13518);
xnor U14012 (N_14012,N_13352,N_13827);
and U14013 (N_14013,N_13254,N_13691);
or U14014 (N_14014,N_13835,N_13402);
and U14015 (N_14015,N_13424,N_13891);
and U14016 (N_14016,N_13140,N_13485);
nand U14017 (N_14017,N_13977,N_13326);
or U14018 (N_14018,N_13173,N_13293);
and U14019 (N_14019,N_13631,N_13760);
xnor U14020 (N_14020,N_13692,N_13549);
and U14021 (N_14021,N_13041,N_13296);
nor U14022 (N_14022,N_13004,N_13916);
nand U14023 (N_14023,N_13821,N_13860);
and U14024 (N_14024,N_13271,N_13218);
nand U14025 (N_14025,N_13629,N_13661);
nand U14026 (N_14026,N_13110,N_13325);
xnor U14027 (N_14027,N_13998,N_13953);
nand U14028 (N_14028,N_13214,N_13146);
nor U14029 (N_14029,N_13528,N_13715);
nand U14030 (N_14030,N_13718,N_13019);
or U14031 (N_14031,N_13383,N_13738);
nor U14032 (N_14032,N_13970,N_13888);
or U14033 (N_14033,N_13353,N_13656);
and U14034 (N_14034,N_13707,N_13674);
or U14035 (N_14035,N_13964,N_13184);
xor U14036 (N_14036,N_13454,N_13109);
nor U14037 (N_14037,N_13039,N_13289);
and U14038 (N_14038,N_13590,N_13924);
and U14039 (N_14039,N_13725,N_13706);
nor U14040 (N_14040,N_13759,N_13127);
and U14041 (N_14041,N_13796,N_13807);
or U14042 (N_14042,N_13076,N_13519);
xnor U14043 (N_14043,N_13018,N_13909);
or U14044 (N_14044,N_13766,N_13502);
and U14045 (N_14045,N_13174,N_13987);
nor U14046 (N_14046,N_13571,N_13726);
xor U14047 (N_14047,N_13358,N_13688);
nor U14048 (N_14048,N_13348,N_13583);
nand U14049 (N_14049,N_13852,N_13495);
xnor U14050 (N_14050,N_13037,N_13989);
nand U14051 (N_14051,N_13842,N_13187);
nand U14052 (N_14052,N_13949,N_13600);
xor U14053 (N_14053,N_13452,N_13260);
and U14054 (N_14054,N_13713,N_13031);
or U14055 (N_14055,N_13845,N_13231);
nor U14056 (N_14056,N_13520,N_13869);
and U14057 (N_14057,N_13151,N_13580);
and U14058 (N_14058,N_13034,N_13002);
or U14059 (N_14059,N_13768,N_13478);
xnor U14060 (N_14060,N_13683,N_13407);
xnor U14061 (N_14061,N_13360,N_13840);
nor U14062 (N_14062,N_13483,N_13010);
or U14063 (N_14063,N_13879,N_13915);
nor U14064 (N_14064,N_13367,N_13711);
or U14065 (N_14065,N_13570,N_13606);
nor U14066 (N_14066,N_13800,N_13277);
xor U14067 (N_14067,N_13224,N_13792);
and U14068 (N_14068,N_13922,N_13665);
and U14069 (N_14069,N_13333,N_13921);
nand U14070 (N_14070,N_13156,N_13124);
nor U14071 (N_14071,N_13132,N_13066);
and U14072 (N_14072,N_13329,N_13469);
or U14073 (N_14073,N_13742,N_13274);
or U14074 (N_14074,N_13737,N_13794);
nand U14075 (N_14075,N_13903,N_13539);
nand U14076 (N_14076,N_13458,N_13605);
and U14077 (N_14077,N_13746,N_13930);
nand U14078 (N_14078,N_13065,N_13636);
nor U14079 (N_14079,N_13475,N_13734);
nor U14080 (N_14080,N_13292,N_13052);
or U14081 (N_14081,N_13536,N_13121);
xor U14082 (N_14082,N_13464,N_13983);
nand U14083 (N_14083,N_13532,N_13428);
nand U14084 (N_14084,N_13462,N_13069);
and U14085 (N_14085,N_13979,N_13769);
xnor U14086 (N_14086,N_13240,N_13847);
and U14087 (N_14087,N_13612,N_13445);
nor U14088 (N_14088,N_13040,N_13350);
nand U14089 (N_14089,N_13543,N_13550);
nor U14090 (N_14090,N_13933,N_13148);
and U14091 (N_14091,N_13617,N_13061);
nand U14092 (N_14092,N_13524,N_13311);
xor U14093 (N_14093,N_13158,N_13681);
and U14094 (N_14094,N_13551,N_13493);
nor U14095 (N_14095,N_13102,N_13955);
nand U14096 (N_14096,N_13802,N_13907);
nor U14097 (N_14097,N_13843,N_13815);
or U14098 (N_14098,N_13745,N_13466);
xor U14099 (N_14099,N_13614,N_13851);
nand U14100 (N_14100,N_13133,N_13494);
and U14101 (N_14101,N_13778,N_13702);
nor U14102 (N_14102,N_13762,N_13561);
nand U14103 (N_14103,N_13413,N_13653);
xor U14104 (N_14104,N_13144,N_13408);
xnor U14105 (N_14105,N_13959,N_13649);
xor U14106 (N_14106,N_13098,N_13247);
nor U14107 (N_14107,N_13832,N_13659);
nand U14108 (N_14108,N_13563,N_13216);
nor U14109 (N_14109,N_13491,N_13730);
or U14110 (N_14110,N_13752,N_13935);
xor U14111 (N_14111,N_13203,N_13431);
nor U14112 (N_14112,N_13474,N_13880);
or U14113 (N_14113,N_13077,N_13128);
or U14114 (N_14114,N_13176,N_13196);
xnor U14115 (N_14115,N_13811,N_13269);
nand U14116 (N_14116,N_13117,N_13107);
or U14117 (N_14117,N_13535,N_13479);
xor U14118 (N_14118,N_13042,N_13958);
nand U14119 (N_14119,N_13836,N_13394);
and U14120 (N_14120,N_13744,N_13722);
nand U14121 (N_14121,N_13048,N_13508);
xnor U14122 (N_14122,N_13417,N_13850);
and U14123 (N_14123,N_13304,N_13434);
or U14124 (N_14124,N_13803,N_13418);
nand U14125 (N_14125,N_13438,N_13676);
nand U14126 (N_14126,N_13461,N_13511);
nand U14127 (N_14127,N_13223,N_13232);
and U14128 (N_14128,N_13498,N_13425);
nor U14129 (N_14129,N_13575,N_13279);
and U14130 (N_14130,N_13763,N_13094);
and U14131 (N_14131,N_13190,N_13748);
xor U14132 (N_14132,N_13113,N_13627);
nor U14133 (N_14133,N_13749,N_13030);
xnor U14134 (N_14134,N_13270,N_13639);
nor U14135 (N_14135,N_13451,N_13777);
and U14136 (N_14136,N_13839,N_13962);
and U14137 (N_14137,N_13599,N_13523);
nor U14138 (N_14138,N_13255,N_13765);
nor U14139 (N_14139,N_13952,N_13626);
nor U14140 (N_14140,N_13172,N_13741);
nor U14141 (N_14141,N_13757,N_13537);
and U14142 (N_14142,N_13586,N_13697);
or U14143 (N_14143,N_13507,N_13138);
nand U14144 (N_14144,N_13059,N_13185);
or U14145 (N_14145,N_13585,N_13758);
nand U14146 (N_14146,N_13897,N_13285);
and U14147 (N_14147,N_13849,N_13488);
nor U14148 (N_14148,N_13645,N_13772);
nand U14149 (N_14149,N_13261,N_13384);
or U14150 (N_14150,N_13305,N_13238);
and U14151 (N_14151,N_13122,N_13510);
or U14152 (N_14152,N_13457,N_13370);
xnor U14153 (N_14153,N_13801,N_13993);
nand U14154 (N_14154,N_13235,N_13552);
or U14155 (N_14155,N_13785,N_13893);
nand U14156 (N_14156,N_13100,N_13638);
and U14157 (N_14157,N_13447,N_13472);
nor U14158 (N_14158,N_13141,N_13275);
nand U14159 (N_14159,N_13966,N_13854);
xnor U14160 (N_14160,N_13167,N_13686);
nand U14161 (N_14161,N_13948,N_13346);
nor U14162 (N_14162,N_13415,N_13985);
xnor U14163 (N_14163,N_13594,N_13157);
xnor U14164 (N_14164,N_13946,N_13319);
nor U14165 (N_14165,N_13833,N_13504);
xnor U14166 (N_14166,N_13743,N_13540);
nand U14167 (N_14167,N_13406,N_13500);
nand U14168 (N_14168,N_13115,N_13327);
or U14169 (N_14169,N_13054,N_13541);
or U14170 (N_14170,N_13694,N_13544);
xor U14171 (N_14171,N_13391,N_13435);
xnor U14172 (N_14172,N_13429,N_13620);
or U14173 (N_14173,N_13817,N_13119);
or U14174 (N_14174,N_13186,N_13669);
xor U14175 (N_14175,N_13633,N_13227);
and U14176 (N_14176,N_13997,N_13120);
nor U14177 (N_14177,N_13682,N_13177);
nor U14178 (N_14178,N_13171,N_13963);
nor U14179 (N_14179,N_13108,N_13318);
nand U14180 (N_14180,N_13487,N_13846);
nor U14181 (N_14181,N_13822,N_13103);
or U14182 (N_14182,N_13191,N_13538);
xnor U14183 (N_14183,N_13058,N_13663);
and U14184 (N_14184,N_13899,N_13482);
nand U14185 (N_14185,N_13377,N_13204);
xor U14186 (N_14186,N_13215,N_13602);
and U14187 (N_14187,N_13404,N_13432);
nand U14188 (N_14188,N_13717,N_13219);
and U14189 (N_14189,N_13032,N_13211);
nand U14190 (N_14190,N_13939,N_13642);
and U14191 (N_14191,N_13818,N_13349);
nor U14192 (N_14192,N_13314,N_13316);
and U14193 (N_14193,N_13033,N_13603);
or U14194 (N_14194,N_13644,N_13099);
nand U14195 (N_14195,N_13199,N_13525);
nand U14196 (N_14196,N_13878,N_13558);
and U14197 (N_14197,N_13134,N_13994);
nand U14198 (N_14198,N_13755,N_13096);
nor U14199 (N_14199,N_13623,N_13727);
and U14200 (N_14200,N_13929,N_13797);
xor U14201 (N_14201,N_13947,N_13135);
nor U14202 (N_14202,N_13233,N_13616);
or U14203 (N_14203,N_13266,N_13877);
or U14204 (N_14204,N_13780,N_13201);
nor U14205 (N_14205,N_13637,N_13856);
nor U14206 (N_14206,N_13978,N_13322);
or U14207 (N_14207,N_13072,N_13608);
or U14208 (N_14208,N_13695,N_13971);
and U14209 (N_14209,N_13687,N_13373);
and U14210 (N_14210,N_13816,N_13272);
nand U14211 (N_14211,N_13043,N_13347);
and U14212 (N_14212,N_13728,N_13806);
nand U14213 (N_14213,N_13870,N_13101);
and U14214 (N_14214,N_13131,N_13601);
or U14215 (N_14215,N_13481,N_13624);
xor U14216 (N_14216,N_13844,N_13906);
or U14217 (N_14217,N_13175,N_13795);
xnor U14218 (N_14218,N_13060,N_13363);
or U14219 (N_14219,N_13496,N_13179);
or U14220 (N_14220,N_13701,N_13864);
nor U14221 (N_14221,N_13992,N_13268);
or U14222 (N_14222,N_13419,N_13973);
and U14223 (N_14223,N_13513,N_13613);
nor U14224 (N_14224,N_13609,N_13841);
nor U14225 (N_14225,N_13904,N_13335);
xor U14226 (N_14226,N_13673,N_13020);
xnor U14227 (N_14227,N_13618,N_13721);
and U14228 (N_14228,N_13622,N_13125);
nand U14229 (N_14229,N_13351,N_13340);
nand U14230 (N_14230,N_13160,N_13658);
nand U14231 (N_14231,N_13943,N_13517);
nor U14232 (N_14232,N_13490,N_13667);
and U14233 (N_14233,N_13996,N_13398);
nand U14234 (N_14234,N_13198,N_13244);
nand U14235 (N_14235,N_13375,N_13611);
or U14236 (N_14236,N_13450,N_13263);
nand U14237 (N_14237,N_13567,N_13063);
or U14238 (N_14238,N_13381,N_13881);
xor U14239 (N_14239,N_13650,N_13761);
nand U14240 (N_14240,N_13308,N_13501);
xor U14241 (N_14241,N_13423,N_13330);
xor U14242 (N_14242,N_13572,N_13055);
or U14243 (N_14243,N_13182,N_13430);
nor U14244 (N_14244,N_13831,N_13087);
and U14245 (N_14245,N_13968,N_13773);
xnor U14246 (N_14246,N_13596,N_13284);
xor U14247 (N_14247,N_13666,N_13183);
or U14248 (N_14248,N_13256,N_13014);
xnor U14249 (N_14249,N_13641,N_13678);
nor U14250 (N_14250,N_13889,N_13643);
xor U14251 (N_14251,N_13262,N_13465);
and U14252 (N_14252,N_13826,N_13712);
xor U14253 (N_14253,N_13385,N_13209);
nor U14254 (N_14254,N_13399,N_13439);
xnor U14255 (N_14255,N_13011,N_13788);
nor U14256 (N_14256,N_13280,N_13693);
nor U14257 (N_14257,N_13781,N_13576);
and U14258 (N_14258,N_13163,N_13876);
xnor U14259 (N_14259,N_13205,N_13793);
and U14260 (N_14260,N_13147,N_13872);
nand U14261 (N_14261,N_13267,N_13514);
and U14262 (N_14262,N_13775,N_13595);
or U14263 (N_14263,N_13926,N_13503);
nor U14264 (N_14264,N_13022,N_13392);
nand U14265 (N_14265,N_13965,N_13791);
or U14266 (N_14266,N_13364,N_13779);
xor U14267 (N_14267,N_13356,N_13867);
nand U14268 (N_14268,N_13288,N_13615);
xor U14269 (N_14269,N_13050,N_13564);
xnor U14270 (N_14270,N_13813,N_13950);
xor U14271 (N_14271,N_13286,N_13111);
xor U14272 (N_14272,N_13009,N_13515);
nor U14273 (N_14273,N_13278,N_13310);
xor U14274 (N_14274,N_13213,N_13938);
xnor U14275 (N_14275,N_13896,N_13253);
or U14276 (N_14276,N_13522,N_13104);
and U14277 (N_14277,N_13095,N_13449);
nor U14278 (N_14278,N_13142,N_13764);
and U14279 (N_14279,N_13632,N_13696);
nand U14280 (N_14280,N_13302,N_13028);
xnor U14281 (N_14281,N_13393,N_13007);
xor U14282 (N_14282,N_13116,N_13448);
nand U14283 (N_14283,N_13901,N_13143);
and U14284 (N_14284,N_13597,N_13008);
and U14285 (N_14285,N_13362,N_13823);
xnor U14286 (N_14286,N_13328,N_13804);
or U14287 (N_14287,N_13243,N_13898);
xor U14288 (N_14288,N_13130,N_13049);
xor U14289 (N_14289,N_13027,N_13887);
or U14290 (N_14290,N_13168,N_13917);
and U14291 (N_14291,N_13660,N_13756);
nand U14292 (N_14292,N_13086,N_13338);
nor U14293 (N_14293,N_13298,N_13732);
or U14294 (N_14294,N_13920,N_13936);
nand U14295 (N_14295,N_13589,N_13276);
xor U14296 (N_14296,N_13303,N_13222);
or U14297 (N_14297,N_13810,N_13798);
nor U14298 (N_14298,N_13092,N_13857);
or U14299 (N_14299,N_13341,N_13956);
nor U14300 (N_14300,N_13700,N_13170);
nand U14301 (N_14301,N_13237,N_13123);
nand U14302 (N_14302,N_13197,N_13584);
and U14303 (N_14303,N_13376,N_13421);
or U14304 (N_14304,N_13581,N_13925);
nor U14305 (N_14305,N_13006,N_13165);
or U14306 (N_14306,N_13015,N_13074);
and U14307 (N_14307,N_13531,N_13720);
and U14308 (N_14308,N_13651,N_13265);
and U14309 (N_14309,N_13212,N_13820);
xnor U14310 (N_14310,N_13509,N_13161);
xor U14311 (N_14311,N_13309,N_13331);
nand U14312 (N_14312,N_13709,N_13357);
xor U14313 (N_14313,N_13866,N_13229);
or U14314 (N_14314,N_13988,N_13467);
nor U14315 (N_14315,N_13405,N_13181);
xnor U14316 (N_14316,N_13868,N_13976);
xnor U14317 (N_14317,N_13067,N_13388);
and U14318 (N_14318,N_13912,N_13361);
nor U14319 (N_14319,N_13366,N_13118);
nand U14320 (N_14320,N_13081,N_13410);
xnor U14321 (N_14321,N_13089,N_13200);
or U14322 (N_14322,N_13740,N_13918);
and U14323 (N_14323,N_13064,N_13646);
nand U14324 (N_14324,N_13648,N_13654);
and U14325 (N_14325,N_13497,N_13705);
or U14326 (N_14326,N_13986,N_13412);
or U14327 (N_14327,N_13610,N_13320);
nand U14328 (N_14328,N_13071,N_13239);
or U14329 (N_14329,N_13657,N_13456);
nor U14330 (N_14330,N_13188,N_13056);
or U14331 (N_14331,N_13675,N_13591);
nor U14332 (N_14332,N_13739,N_13306);
xor U14333 (N_14333,N_13001,N_13771);
nor U14334 (N_14334,N_13137,N_13097);
xor U14335 (N_14335,N_13937,N_13026);
xor U14336 (N_14336,N_13044,N_13805);
nand U14337 (N_14337,N_13248,N_13960);
nor U14338 (N_14338,N_13105,N_13565);
or U14339 (N_14339,N_13075,N_13910);
and U14340 (N_14340,N_13312,N_13865);
and U14341 (N_14341,N_13652,N_13257);
nor U14342 (N_14342,N_13114,N_13139);
xor U14343 (N_14343,N_13382,N_13057);
nor U14344 (N_14344,N_13295,N_13714);
nor U14345 (N_14345,N_13884,N_13577);
xnor U14346 (N_14346,N_13273,N_13829);
xnor U14347 (N_14347,N_13991,N_13516);
nor U14348 (N_14348,N_13545,N_13945);
nor U14349 (N_14349,N_13371,N_13024);
or U14350 (N_14350,N_13226,N_13068);
nand U14351 (N_14351,N_13153,N_13940);
nor U14352 (N_14352,N_13194,N_13716);
or U14353 (N_14353,N_13557,N_13900);
xor U14354 (N_14354,N_13928,N_13149);
or U14355 (N_14355,N_13073,N_13374);
nor U14356 (N_14356,N_13974,N_13420);
xnor U14357 (N_14357,N_13954,N_13981);
nor U14358 (N_14358,N_13982,N_13178);
nor U14359 (N_14359,N_13051,N_13914);
nand U14360 (N_14360,N_13786,N_13664);
and U14361 (N_14361,N_13345,N_13192);
nor U14362 (N_14362,N_13812,N_13895);
nand U14363 (N_14363,N_13202,N_13790);
nor U14364 (N_14364,N_13588,N_13995);
xnor U14365 (N_14365,N_13972,N_13554);
and U14366 (N_14366,N_13294,N_13162);
xnor U14367 (N_14367,N_13246,N_13750);
or U14368 (N_14368,N_13206,N_13848);
nand U14369 (N_14369,N_13250,N_13000);
nor U14370 (N_14370,N_13855,N_13228);
xor U14371 (N_14371,N_13783,N_13070);
nand U14372 (N_14372,N_13249,N_13853);
nand U14373 (N_14373,N_13908,N_13677);
or U14374 (N_14374,N_13281,N_13578);
nor U14375 (N_14375,N_13241,N_13217);
or U14376 (N_14376,N_13913,N_13710);
or U14377 (N_14377,N_13290,N_13886);
nand U14378 (N_14378,N_13468,N_13210);
and U14379 (N_14379,N_13662,N_13332);
and U14380 (N_14380,N_13980,N_13619);
or U14381 (N_14381,N_13337,N_13164);
xnor U14382 (N_14382,N_13283,N_13021);
and U14383 (N_14383,N_13442,N_13441);
xnor U14384 (N_14384,N_13808,N_13091);
or U14385 (N_14385,N_13708,N_13324);
and U14386 (N_14386,N_13013,N_13136);
and U14387 (N_14387,N_13824,N_13368);
nand U14388 (N_14388,N_13892,N_13409);
nor U14389 (N_14389,N_13593,N_13344);
nor U14390 (N_14390,N_13023,N_13476);
xor U14391 (N_14391,N_13628,N_13470);
and U14392 (N_14392,N_13090,N_13967);
nand U14393 (N_14393,N_13934,N_13975);
and U14394 (N_14394,N_13512,N_13598);
and U14395 (N_14395,N_13321,N_13751);
nand U14396 (N_14396,N_13556,N_13574);
and U14397 (N_14397,N_13225,N_13258);
xor U14398 (N_14398,N_13990,N_13047);
nor U14399 (N_14399,N_13607,N_13416);
nand U14400 (N_14400,N_13703,N_13883);
nand U14401 (N_14401,N_13830,N_13873);
nand U14402 (N_14402,N_13236,N_13342);
nand U14403 (N_14403,N_13690,N_13754);
nor U14404 (N_14404,N_13984,N_13221);
nor U14405 (N_14405,N_13106,N_13301);
and U14406 (N_14406,N_13150,N_13154);
nor U14407 (N_14407,N_13486,N_13427);
and U14408 (N_14408,N_13460,N_13957);
or U14409 (N_14409,N_13894,N_13559);
nor U14410 (N_14410,N_13861,N_13230);
nand U14411 (N_14411,N_13369,N_13315);
nand U14412 (N_14412,N_13307,N_13814);
nor U14413 (N_14413,N_13379,N_13569);
or U14414 (N_14414,N_13529,N_13477);
or U14415 (N_14415,N_13169,N_13679);
nor U14416 (N_14416,N_13999,N_13489);
nor U14417 (N_14417,N_13025,N_13029);
and U14418 (N_14418,N_13471,N_13252);
and U14419 (N_14419,N_13621,N_13411);
xnor U14420 (N_14420,N_13723,N_13735);
or U14421 (N_14421,N_13724,N_13422);
and U14422 (N_14422,N_13733,N_13680);
and U14423 (N_14423,N_13685,N_13942);
or U14424 (N_14424,N_13582,N_13579);
or U14425 (N_14425,N_13573,N_13767);
xor U14426 (N_14426,N_13944,N_13088);
nand U14427 (N_14427,N_13635,N_13526);
nand U14428 (N_14428,N_13634,N_13927);
and U14429 (N_14429,N_13291,N_13670);
nand U14430 (N_14430,N_13195,N_13546);
nand U14431 (N_14431,N_13560,N_13587);
nand U14432 (N_14432,N_13951,N_13480);
nor U14433 (N_14433,N_13297,N_13264);
or U14434 (N_14434,N_13336,N_13389);
nor U14435 (N_14435,N_13542,N_13902);
or U14436 (N_14436,N_13919,N_13453);
or U14437 (N_14437,N_13863,N_13005);
nand U14438 (N_14438,N_13885,N_13862);
or U14439 (N_14439,N_13825,N_13380);
and U14440 (N_14440,N_13647,N_13530);
xnor U14441 (N_14441,N_13395,N_13129);
or U14442 (N_14442,N_13672,N_13443);
xnor U14443 (N_14443,N_13414,N_13671);
and U14444 (N_14444,N_13630,N_13729);
and U14445 (N_14445,N_13062,N_13365);
nor U14446 (N_14446,N_13625,N_13245);
xor U14447 (N_14447,N_13799,N_13874);
nor U14448 (N_14448,N_13704,N_13747);
nor U14449 (N_14449,N_13343,N_13553);
xor U14450 (N_14450,N_13046,N_13941);
xor U14451 (N_14451,N_13166,N_13932);
nand U14452 (N_14452,N_13961,N_13220);
xnor U14453 (N_14453,N_13834,N_13355);
nor U14454 (N_14454,N_13604,N_13189);
xnor U14455 (N_14455,N_13890,N_13828);
nand U14456 (N_14456,N_13459,N_13882);
or U14457 (N_14457,N_13378,N_13012);
or U14458 (N_14458,N_13242,N_13437);
or U14459 (N_14459,N_13079,N_13871);
xnor U14460 (N_14460,N_13774,N_13017);
or U14461 (N_14461,N_13440,N_13038);
nand U14462 (N_14462,N_13159,N_13155);
or U14463 (N_14463,N_13484,N_13396);
or U14464 (N_14464,N_13003,N_13776);
xor U14465 (N_14465,N_13787,N_13299);
or U14466 (N_14466,N_13193,N_13045);
xor U14467 (N_14467,N_13208,N_13084);
nor U14468 (N_14468,N_13145,N_13499);
nor U14469 (N_14469,N_13689,N_13400);
nor U14470 (N_14470,N_13282,N_13080);
nand U14471 (N_14471,N_13789,N_13397);
or U14472 (N_14472,N_13259,N_13313);
or U14473 (N_14473,N_13083,N_13455);
and U14474 (N_14474,N_13911,N_13463);
and U14475 (N_14475,N_13082,N_13180);
nand U14476 (N_14476,N_13207,N_13359);
and U14477 (N_14477,N_13562,N_13339);
and U14478 (N_14478,N_13782,N_13433);
or U14479 (N_14479,N_13521,N_13035);
and U14480 (N_14480,N_13699,N_13387);
nor U14481 (N_14481,N_13390,N_13592);
or U14482 (N_14482,N_13505,N_13436);
and U14483 (N_14483,N_13859,N_13152);
nand U14484 (N_14484,N_13731,N_13905);
nor U14485 (N_14485,N_13533,N_13093);
or U14486 (N_14486,N_13837,N_13923);
xnor U14487 (N_14487,N_13053,N_13736);
and U14488 (N_14488,N_13555,N_13719);
or U14489 (N_14489,N_13931,N_13534);
xor U14490 (N_14490,N_13838,N_13668);
nor U14491 (N_14491,N_13444,N_13784);
xor U14492 (N_14492,N_13527,N_13334);
and U14493 (N_14493,N_13492,N_13770);
or U14494 (N_14494,N_13016,N_13548);
nor U14495 (N_14495,N_13403,N_13446);
nor U14496 (N_14496,N_13473,N_13234);
xnor U14497 (N_14497,N_13287,N_13753);
xnor U14498 (N_14498,N_13858,N_13372);
nor U14499 (N_14499,N_13085,N_13698);
nand U14500 (N_14500,N_13659,N_13763);
and U14501 (N_14501,N_13805,N_13059);
and U14502 (N_14502,N_13640,N_13435);
or U14503 (N_14503,N_13388,N_13757);
xnor U14504 (N_14504,N_13056,N_13754);
nor U14505 (N_14505,N_13706,N_13718);
or U14506 (N_14506,N_13032,N_13633);
nor U14507 (N_14507,N_13136,N_13220);
nor U14508 (N_14508,N_13192,N_13823);
or U14509 (N_14509,N_13340,N_13330);
nand U14510 (N_14510,N_13415,N_13436);
or U14511 (N_14511,N_13682,N_13805);
xnor U14512 (N_14512,N_13344,N_13042);
and U14513 (N_14513,N_13673,N_13961);
nor U14514 (N_14514,N_13392,N_13841);
and U14515 (N_14515,N_13047,N_13541);
or U14516 (N_14516,N_13281,N_13293);
nand U14517 (N_14517,N_13676,N_13725);
nor U14518 (N_14518,N_13197,N_13779);
or U14519 (N_14519,N_13949,N_13391);
and U14520 (N_14520,N_13377,N_13118);
xor U14521 (N_14521,N_13602,N_13532);
nand U14522 (N_14522,N_13881,N_13427);
nand U14523 (N_14523,N_13779,N_13343);
xnor U14524 (N_14524,N_13679,N_13655);
xnor U14525 (N_14525,N_13739,N_13510);
xnor U14526 (N_14526,N_13038,N_13708);
nand U14527 (N_14527,N_13160,N_13065);
and U14528 (N_14528,N_13708,N_13525);
and U14529 (N_14529,N_13855,N_13802);
and U14530 (N_14530,N_13282,N_13591);
nor U14531 (N_14531,N_13332,N_13475);
or U14532 (N_14532,N_13612,N_13391);
or U14533 (N_14533,N_13882,N_13161);
and U14534 (N_14534,N_13920,N_13398);
or U14535 (N_14535,N_13466,N_13990);
and U14536 (N_14536,N_13228,N_13643);
nor U14537 (N_14537,N_13466,N_13924);
nand U14538 (N_14538,N_13628,N_13350);
xor U14539 (N_14539,N_13701,N_13726);
nor U14540 (N_14540,N_13807,N_13610);
nor U14541 (N_14541,N_13373,N_13329);
nand U14542 (N_14542,N_13540,N_13380);
nand U14543 (N_14543,N_13004,N_13226);
and U14544 (N_14544,N_13924,N_13887);
or U14545 (N_14545,N_13867,N_13620);
xnor U14546 (N_14546,N_13711,N_13239);
or U14547 (N_14547,N_13045,N_13226);
nand U14548 (N_14548,N_13744,N_13715);
nor U14549 (N_14549,N_13218,N_13972);
or U14550 (N_14550,N_13551,N_13778);
xor U14551 (N_14551,N_13813,N_13852);
xor U14552 (N_14552,N_13256,N_13249);
xor U14553 (N_14553,N_13503,N_13481);
nand U14554 (N_14554,N_13921,N_13545);
or U14555 (N_14555,N_13737,N_13073);
xnor U14556 (N_14556,N_13684,N_13396);
xor U14557 (N_14557,N_13185,N_13140);
nor U14558 (N_14558,N_13357,N_13822);
xnor U14559 (N_14559,N_13093,N_13806);
or U14560 (N_14560,N_13936,N_13493);
xnor U14561 (N_14561,N_13978,N_13790);
nand U14562 (N_14562,N_13339,N_13656);
xnor U14563 (N_14563,N_13733,N_13435);
or U14564 (N_14564,N_13477,N_13746);
or U14565 (N_14565,N_13614,N_13181);
and U14566 (N_14566,N_13037,N_13036);
and U14567 (N_14567,N_13488,N_13984);
and U14568 (N_14568,N_13747,N_13752);
or U14569 (N_14569,N_13039,N_13884);
nor U14570 (N_14570,N_13582,N_13704);
nor U14571 (N_14571,N_13089,N_13658);
and U14572 (N_14572,N_13775,N_13510);
or U14573 (N_14573,N_13038,N_13015);
nand U14574 (N_14574,N_13717,N_13341);
and U14575 (N_14575,N_13980,N_13972);
xor U14576 (N_14576,N_13244,N_13701);
and U14577 (N_14577,N_13151,N_13859);
and U14578 (N_14578,N_13104,N_13678);
nor U14579 (N_14579,N_13667,N_13375);
nand U14580 (N_14580,N_13015,N_13475);
and U14581 (N_14581,N_13312,N_13597);
xnor U14582 (N_14582,N_13674,N_13003);
xor U14583 (N_14583,N_13162,N_13575);
xor U14584 (N_14584,N_13585,N_13997);
or U14585 (N_14585,N_13971,N_13315);
or U14586 (N_14586,N_13613,N_13299);
nor U14587 (N_14587,N_13603,N_13599);
nand U14588 (N_14588,N_13294,N_13621);
and U14589 (N_14589,N_13695,N_13669);
and U14590 (N_14590,N_13817,N_13763);
or U14591 (N_14591,N_13874,N_13274);
and U14592 (N_14592,N_13365,N_13162);
nor U14593 (N_14593,N_13748,N_13069);
and U14594 (N_14594,N_13901,N_13375);
nand U14595 (N_14595,N_13836,N_13978);
or U14596 (N_14596,N_13570,N_13399);
xnor U14597 (N_14597,N_13532,N_13019);
and U14598 (N_14598,N_13354,N_13360);
nor U14599 (N_14599,N_13194,N_13037);
xnor U14600 (N_14600,N_13314,N_13479);
nand U14601 (N_14601,N_13791,N_13357);
nand U14602 (N_14602,N_13739,N_13775);
nor U14603 (N_14603,N_13610,N_13913);
nor U14604 (N_14604,N_13096,N_13943);
or U14605 (N_14605,N_13302,N_13875);
and U14606 (N_14606,N_13524,N_13306);
nor U14607 (N_14607,N_13318,N_13822);
nand U14608 (N_14608,N_13598,N_13354);
nor U14609 (N_14609,N_13437,N_13570);
nor U14610 (N_14610,N_13286,N_13332);
xnor U14611 (N_14611,N_13072,N_13039);
xnor U14612 (N_14612,N_13651,N_13487);
nor U14613 (N_14613,N_13007,N_13841);
and U14614 (N_14614,N_13454,N_13121);
and U14615 (N_14615,N_13916,N_13194);
xor U14616 (N_14616,N_13922,N_13972);
and U14617 (N_14617,N_13220,N_13854);
and U14618 (N_14618,N_13016,N_13059);
xor U14619 (N_14619,N_13014,N_13060);
xor U14620 (N_14620,N_13298,N_13323);
and U14621 (N_14621,N_13389,N_13114);
and U14622 (N_14622,N_13720,N_13833);
nand U14623 (N_14623,N_13816,N_13576);
xnor U14624 (N_14624,N_13413,N_13250);
or U14625 (N_14625,N_13219,N_13831);
xnor U14626 (N_14626,N_13157,N_13035);
xnor U14627 (N_14627,N_13466,N_13130);
nand U14628 (N_14628,N_13150,N_13604);
nor U14629 (N_14629,N_13867,N_13951);
nor U14630 (N_14630,N_13829,N_13077);
xnor U14631 (N_14631,N_13609,N_13718);
xnor U14632 (N_14632,N_13390,N_13759);
and U14633 (N_14633,N_13715,N_13493);
nor U14634 (N_14634,N_13499,N_13983);
nor U14635 (N_14635,N_13519,N_13326);
and U14636 (N_14636,N_13184,N_13342);
or U14637 (N_14637,N_13759,N_13997);
xor U14638 (N_14638,N_13484,N_13251);
nand U14639 (N_14639,N_13805,N_13596);
nand U14640 (N_14640,N_13951,N_13342);
or U14641 (N_14641,N_13083,N_13398);
or U14642 (N_14642,N_13550,N_13308);
nand U14643 (N_14643,N_13117,N_13618);
nor U14644 (N_14644,N_13496,N_13988);
or U14645 (N_14645,N_13740,N_13598);
or U14646 (N_14646,N_13925,N_13500);
xor U14647 (N_14647,N_13293,N_13772);
or U14648 (N_14648,N_13728,N_13505);
xor U14649 (N_14649,N_13042,N_13259);
nand U14650 (N_14650,N_13117,N_13943);
nand U14651 (N_14651,N_13178,N_13312);
nand U14652 (N_14652,N_13508,N_13909);
nand U14653 (N_14653,N_13586,N_13461);
xor U14654 (N_14654,N_13640,N_13788);
or U14655 (N_14655,N_13062,N_13711);
xor U14656 (N_14656,N_13041,N_13946);
and U14657 (N_14657,N_13474,N_13926);
or U14658 (N_14658,N_13235,N_13267);
nand U14659 (N_14659,N_13464,N_13817);
xnor U14660 (N_14660,N_13662,N_13903);
nand U14661 (N_14661,N_13955,N_13932);
nor U14662 (N_14662,N_13903,N_13404);
or U14663 (N_14663,N_13899,N_13832);
xor U14664 (N_14664,N_13640,N_13665);
nand U14665 (N_14665,N_13545,N_13497);
nor U14666 (N_14666,N_13751,N_13710);
nand U14667 (N_14667,N_13532,N_13272);
or U14668 (N_14668,N_13765,N_13226);
xnor U14669 (N_14669,N_13905,N_13736);
nand U14670 (N_14670,N_13508,N_13530);
nand U14671 (N_14671,N_13775,N_13138);
nand U14672 (N_14672,N_13286,N_13198);
or U14673 (N_14673,N_13487,N_13143);
nor U14674 (N_14674,N_13803,N_13965);
xnor U14675 (N_14675,N_13374,N_13868);
xor U14676 (N_14676,N_13025,N_13178);
and U14677 (N_14677,N_13708,N_13644);
or U14678 (N_14678,N_13937,N_13615);
nor U14679 (N_14679,N_13355,N_13098);
or U14680 (N_14680,N_13704,N_13864);
xnor U14681 (N_14681,N_13189,N_13987);
and U14682 (N_14682,N_13920,N_13742);
xnor U14683 (N_14683,N_13119,N_13282);
nor U14684 (N_14684,N_13697,N_13376);
xor U14685 (N_14685,N_13931,N_13367);
nor U14686 (N_14686,N_13681,N_13597);
xor U14687 (N_14687,N_13937,N_13929);
and U14688 (N_14688,N_13709,N_13291);
nand U14689 (N_14689,N_13001,N_13016);
and U14690 (N_14690,N_13783,N_13349);
xnor U14691 (N_14691,N_13070,N_13925);
xnor U14692 (N_14692,N_13107,N_13646);
or U14693 (N_14693,N_13523,N_13983);
and U14694 (N_14694,N_13379,N_13917);
or U14695 (N_14695,N_13295,N_13072);
nand U14696 (N_14696,N_13166,N_13457);
nor U14697 (N_14697,N_13053,N_13929);
and U14698 (N_14698,N_13350,N_13621);
or U14699 (N_14699,N_13965,N_13384);
or U14700 (N_14700,N_13175,N_13326);
nor U14701 (N_14701,N_13408,N_13589);
and U14702 (N_14702,N_13222,N_13694);
and U14703 (N_14703,N_13553,N_13504);
nand U14704 (N_14704,N_13487,N_13262);
nor U14705 (N_14705,N_13996,N_13069);
nand U14706 (N_14706,N_13961,N_13965);
nand U14707 (N_14707,N_13589,N_13955);
and U14708 (N_14708,N_13170,N_13593);
and U14709 (N_14709,N_13018,N_13821);
nor U14710 (N_14710,N_13064,N_13783);
and U14711 (N_14711,N_13285,N_13679);
nor U14712 (N_14712,N_13367,N_13280);
and U14713 (N_14713,N_13380,N_13393);
and U14714 (N_14714,N_13453,N_13602);
or U14715 (N_14715,N_13230,N_13212);
nor U14716 (N_14716,N_13027,N_13730);
or U14717 (N_14717,N_13905,N_13412);
and U14718 (N_14718,N_13473,N_13287);
xnor U14719 (N_14719,N_13013,N_13530);
nand U14720 (N_14720,N_13661,N_13582);
nor U14721 (N_14721,N_13053,N_13774);
and U14722 (N_14722,N_13890,N_13682);
nor U14723 (N_14723,N_13456,N_13945);
nand U14724 (N_14724,N_13268,N_13682);
xor U14725 (N_14725,N_13532,N_13283);
and U14726 (N_14726,N_13321,N_13252);
nor U14727 (N_14727,N_13133,N_13818);
xnor U14728 (N_14728,N_13354,N_13910);
or U14729 (N_14729,N_13641,N_13698);
xnor U14730 (N_14730,N_13777,N_13271);
nand U14731 (N_14731,N_13172,N_13629);
or U14732 (N_14732,N_13633,N_13843);
nand U14733 (N_14733,N_13418,N_13581);
and U14734 (N_14734,N_13918,N_13344);
or U14735 (N_14735,N_13062,N_13969);
xor U14736 (N_14736,N_13609,N_13571);
or U14737 (N_14737,N_13566,N_13802);
or U14738 (N_14738,N_13868,N_13019);
or U14739 (N_14739,N_13826,N_13050);
nor U14740 (N_14740,N_13645,N_13050);
nand U14741 (N_14741,N_13816,N_13036);
nand U14742 (N_14742,N_13090,N_13180);
or U14743 (N_14743,N_13822,N_13983);
or U14744 (N_14744,N_13252,N_13987);
or U14745 (N_14745,N_13084,N_13306);
nand U14746 (N_14746,N_13235,N_13027);
nor U14747 (N_14747,N_13992,N_13171);
nand U14748 (N_14748,N_13389,N_13264);
nand U14749 (N_14749,N_13221,N_13384);
nand U14750 (N_14750,N_13846,N_13281);
or U14751 (N_14751,N_13534,N_13735);
or U14752 (N_14752,N_13695,N_13694);
and U14753 (N_14753,N_13146,N_13221);
nor U14754 (N_14754,N_13441,N_13781);
and U14755 (N_14755,N_13278,N_13631);
nand U14756 (N_14756,N_13947,N_13941);
and U14757 (N_14757,N_13969,N_13272);
and U14758 (N_14758,N_13697,N_13201);
and U14759 (N_14759,N_13948,N_13447);
xor U14760 (N_14760,N_13934,N_13929);
nand U14761 (N_14761,N_13818,N_13319);
nand U14762 (N_14762,N_13176,N_13582);
and U14763 (N_14763,N_13750,N_13923);
xnor U14764 (N_14764,N_13511,N_13733);
nor U14765 (N_14765,N_13819,N_13636);
and U14766 (N_14766,N_13257,N_13173);
or U14767 (N_14767,N_13653,N_13664);
xnor U14768 (N_14768,N_13199,N_13264);
or U14769 (N_14769,N_13699,N_13287);
xor U14770 (N_14770,N_13046,N_13205);
nor U14771 (N_14771,N_13541,N_13521);
and U14772 (N_14772,N_13708,N_13174);
xnor U14773 (N_14773,N_13561,N_13929);
and U14774 (N_14774,N_13182,N_13853);
xnor U14775 (N_14775,N_13401,N_13620);
or U14776 (N_14776,N_13686,N_13456);
and U14777 (N_14777,N_13954,N_13940);
nand U14778 (N_14778,N_13832,N_13042);
or U14779 (N_14779,N_13941,N_13666);
and U14780 (N_14780,N_13857,N_13628);
and U14781 (N_14781,N_13533,N_13070);
and U14782 (N_14782,N_13579,N_13026);
xor U14783 (N_14783,N_13449,N_13006);
and U14784 (N_14784,N_13114,N_13796);
or U14785 (N_14785,N_13324,N_13287);
nand U14786 (N_14786,N_13294,N_13817);
nor U14787 (N_14787,N_13183,N_13497);
and U14788 (N_14788,N_13725,N_13088);
nand U14789 (N_14789,N_13595,N_13840);
xor U14790 (N_14790,N_13647,N_13944);
nand U14791 (N_14791,N_13410,N_13834);
nor U14792 (N_14792,N_13150,N_13936);
xor U14793 (N_14793,N_13924,N_13597);
nor U14794 (N_14794,N_13149,N_13001);
xnor U14795 (N_14795,N_13435,N_13499);
nand U14796 (N_14796,N_13321,N_13457);
xnor U14797 (N_14797,N_13007,N_13199);
and U14798 (N_14798,N_13029,N_13245);
and U14799 (N_14799,N_13194,N_13311);
and U14800 (N_14800,N_13706,N_13768);
nand U14801 (N_14801,N_13797,N_13759);
xor U14802 (N_14802,N_13094,N_13308);
nand U14803 (N_14803,N_13039,N_13980);
nand U14804 (N_14804,N_13044,N_13515);
xor U14805 (N_14805,N_13023,N_13329);
nor U14806 (N_14806,N_13243,N_13479);
and U14807 (N_14807,N_13721,N_13174);
and U14808 (N_14808,N_13592,N_13365);
or U14809 (N_14809,N_13570,N_13821);
and U14810 (N_14810,N_13476,N_13116);
and U14811 (N_14811,N_13442,N_13940);
and U14812 (N_14812,N_13772,N_13519);
nor U14813 (N_14813,N_13096,N_13229);
xnor U14814 (N_14814,N_13648,N_13899);
xnor U14815 (N_14815,N_13428,N_13356);
xor U14816 (N_14816,N_13028,N_13602);
xor U14817 (N_14817,N_13089,N_13353);
nor U14818 (N_14818,N_13643,N_13281);
xnor U14819 (N_14819,N_13417,N_13001);
and U14820 (N_14820,N_13140,N_13143);
nor U14821 (N_14821,N_13243,N_13022);
xnor U14822 (N_14822,N_13350,N_13860);
nor U14823 (N_14823,N_13212,N_13547);
xor U14824 (N_14824,N_13432,N_13445);
nor U14825 (N_14825,N_13744,N_13483);
nand U14826 (N_14826,N_13647,N_13780);
and U14827 (N_14827,N_13867,N_13412);
nand U14828 (N_14828,N_13433,N_13480);
nand U14829 (N_14829,N_13201,N_13604);
or U14830 (N_14830,N_13567,N_13749);
xor U14831 (N_14831,N_13312,N_13321);
nor U14832 (N_14832,N_13193,N_13186);
nor U14833 (N_14833,N_13252,N_13187);
or U14834 (N_14834,N_13926,N_13262);
nand U14835 (N_14835,N_13731,N_13535);
or U14836 (N_14836,N_13373,N_13527);
or U14837 (N_14837,N_13186,N_13778);
nor U14838 (N_14838,N_13609,N_13668);
and U14839 (N_14839,N_13202,N_13626);
xnor U14840 (N_14840,N_13128,N_13950);
and U14841 (N_14841,N_13136,N_13467);
xnor U14842 (N_14842,N_13232,N_13616);
nor U14843 (N_14843,N_13823,N_13675);
nand U14844 (N_14844,N_13049,N_13399);
nand U14845 (N_14845,N_13676,N_13031);
and U14846 (N_14846,N_13033,N_13739);
or U14847 (N_14847,N_13794,N_13516);
xor U14848 (N_14848,N_13409,N_13584);
xnor U14849 (N_14849,N_13160,N_13105);
and U14850 (N_14850,N_13893,N_13708);
and U14851 (N_14851,N_13663,N_13692);
nor U14852 (N_14852,N_13624,N_13897);
and U14853 (N_14853,N_13119,N_13726);
and U14854 (N_14854,N_13461,N_13708);
or U14855 (N_14855,N_13187,N_13742);
xor U14856 (N_14856,N_13177,N_13350);
or U14857 (N_14857,N_13070,N_13459);
or U14858 (N_14858,N_13666,N_13264);
nor U14859 (N_14859,N_13430,N_13248);
nor U14860 (N_14860,N_13305,N_13071);
and U14861 (N_14861,N_13707,N_13983);
or U14862 (N_14862,N_13495,N_13426);
nand U14863 (N_14863,N_13379,N_13404);
xor U14864 (N_14864,N_13639,N_13654);
xnor U14865 (N_14865,N_13431,N_13925);
or U14866 (N_14866,N_13436,N_13132);
and U14867 (N_14867,N_13541,N_13108);
xnor U14868 (N_14868,N_13148,N_13381);
nor U14869 (N_14869,N_13393,N_13869);
and U14870 (N_14870,N_13379,N_13766);
nand U14871 (N_14871,N_13186,N_13954);
xor U14872 (N_14872,N_13223,N_13876);
xnor U14873 (N_14873,N_13484,N_13912);
or U14874 (N_14874,N_13676,N_13808);
nor U14875 (N_14875,N_13196,N_13167);
nor U14876 (N_14876,N_13301,N_13851);
or U14877 (N_14877,N_13158,N_13917);
or U14878 (N_14878,N_13463,N_13306);
nor U14879 (N_14879,N_13394,N_13725);
or U14880 (N_14880,N_13614,N_13279);
nand U14881 (N_14881,N_13311,N_13322);
or U14882 (N_14882,N_13782,N_13232);
nor U14883 (N_14883,N_13756,N_13168);
nand U14884 (N_14884,N_13550,N_13362);
nor U14885 (N_14885,N_13660,N_13585);
nor U14886 (N_14886,N_13296,N_13774);
nor U14887 (N_14887,N_13764,N_13487);
or U14888 (N_14888,N_13867,N_13683);
and U14889 (N_14889,N_13142,N_13548);
or U14890 (N_14890,N_13339,N_13465);
or U14891 (N_14891,N_13518,N_13002);
nand U14892 (N_14892,N_13744,N_13909);
nor U14893 (N_14893,N_13448,N_13206);
or U14894 (N_14894,N_13878,N_13167);
or U14895 (N_14895,N_13092,N_13419);
and U14896 (N_14896,N_13973,N_13020);
nor U14897 (N_14897,N_13473,N_13771);
xor U14898 (N_14898,N_13907,N_13575);
nand U14899 (N_14899,N_13222,N_13241);
and U14900 (N_14900,N_13378,N_13649);
nand U14901 (N_14901,N_13972,N_13266);
or U14902 (N_14902,N_13651,N_13065);
nor U14903 (N_14903,N_13940,N_13794);
and U14904 (N_14904,N_13423,N_13919);
and U14905 (N_14905,N_13975,N_13355);
nor U14906 (N_14906,N_13873,N_13366);
nor U14907 (N_14907,N_13185,N_13188);
xnor U14908 (N_14908,N_13029,N_13649);
nand U14909 (N_14909,N_13367,N_13320);
and U14910 (N_14910,N_13335,N_13586);
xnor U14911 (N_14911,N_13511,N_13774);
and U14912 (N_14912,N_13093,N_13729);
xor U14913 (N_14913,N_13746,N_13885);
and U14914 (N_14914,N_13316,N_13021);
and U14915 (N_14915,N_13173,N_13096);
and U14916 (N_14916,N_13096,N_13775);
xnor U14917 (N_14917,N_13429,N_13380);
nand U14918 (N_14918,N_13161,N_13625);
nand U14919 (N_14919,N_13023,N_13461);
nor U14920 (N_14920,N_13735,N_13545);
nand U14921 (N_14921,N_13231,N_13836);
or U14922 (N_14922,N_13776,N_13335);
nor U14923 (N_14923,N_13671,N_13912);
and U14924 (N_14924,N_13217,N_13849);
xnor U14925 (N_14925,N_13005,N_13543);
nor U14926 (N_14926,N_13498,N_13476);
or U14927 (N_14927,N_13045,N_13841);
nor U14928 (N_14928,N_13357,N_13850);
nand U14929 (N_14929,N_13473,N_13725);
or U14930 (N_14930,N_13681,N_13737);
xnor U14931 (N_14931,N_13746,N_13431);
nand U14932 (N_14932,N_13744,N_13020);
xnor U14933 (N_14933,N_13135,N_13701);
nor U14934 (N_14934,N_13156,N_13937);
nand U14935 (N_14935,N_13105,N_13779);
xor U14936 (N_14936,N_13754,N_13871);
nand U14937 (N_14937,N_13395,N_13972);
xor U14938 (N_14938,N_13685,N_13983);
or U14939 (N_14939,N_13144,N_13583);
nor U14940 (N_14940,N_13876,N_13886);
or U14941 (N_14941,N_13294,N_13210);
and U14942 (N_14942,N_13306,N_13634);
nand U14943 (N_14943,N_13972,N_13164);
nand U14944 (N_14944,N_13888,N_13827);
or U14945 (N_14945,N_13006,N_13748);
or U14946 (N_14946,N_13661,N_13786);
nor U14947 (N_14947,N_13904,N_13214);
xnor U14948 (N_14948,N_13699,N_13962);
xnor U14949 (N_14949,N_13567,N_13100);
nand U14950 (N_14950,N_13542,N_13044);
and U14951 (N_14951,N_13214,N_13788);
and U14952 (N_14952,N_13321,N_13475);
or U14953 (N_14953,N_13961,N_13848);
and U14954 (N_14954,N_13955,N_13054);
and U14955 (N_14955,N_13480,N_13818);
nand U14956 (N_14956,N_13125,N_13569);
or U14957 (N_14957,N_13110,N_13960);
xnor U14958 (N_14958,N_13865,N_13145);
xnor U14959 (N_14959,N_13893,N_13310);
or U14960 (N_14960,N_13274,N_13088);
or U14961 (N_14961,N_13748,N_13618);
or U14962 (N_14962,N_13333,N_13347);
xor U14963 (N_14963,N_13006,N_13895);
and U14964 (N_14964,N_13486,N_13884);
nand U14965 (N_14965,N_13417,N_13754);
or U14966 (N_14966,N_13533,N_13104);
nor U14967 (N_14967,N_13922,N_13237);
and U14968 (N_14968,N_13246,N_13955);
xnor U14969 (N_14969,N_13810,N_13158);
and U14970 (N_14970,N_13155,N_13726);
nor U14971 (N_14971,N_13416,N_13508);
and U14972 (N_14972,N_13418,N_13059);
and U14973 (N_14973,N_13180,N_13681);
nor U14974 (N_14974,N_13666,N_13606);
or U14975 (N_14975,N_13686,N_13900);
or U14976 (N_14976,N_13564,N_13501);
nand U14977 (N_14977,N_13862,N_13483);
and U14978 (N_14978,N_13941,N_13982);
nor U14979 (N_14979,N_13868,N_13614);
nor U14980 (N_14980,N_13069,N_13962);
nor U14981 (N_14981,N_13120,N_13573);
nand U14982 (N_14982,N_13281,N_13799);
and U14983 (N_14983,N_13147,N_13516);
or U14984 (N_14984,N_13371,N_13119);
nand U14985 (N_14985,N_13294,N_13685);
nor U14986 (N_14986,N_13018,N_13572);
or U14987 (N_14987,N_13269,N_13124);
and U14988 (N_14988,N_13991,N_13866);
nand U14989 (N_14989,N_13740,N_13672);
or U14990 (N_14990,N_13520,N_13199);
or U14991 (N_14991,N_13198,N_13336);
nor U14992 (N_14992,N_13763,N_13905);
xor U14993 (N_14993,N_13659,N_13486);
or U14994 (N_14994,N_13768,N_13632);
nor U14995 (N_14995,N_13984,N_13355);
or U14996 (N_14996,N_13908,N_13957);
nor U14997 (N_14997,N_13385,N_13484);
xor U14998 (N_14998,N_13312,N_13696);
xnor U14999 (N_14999,N_13728,N_13211);
nand U15000 (N_15000,N_14652,N_14674);
and U15001 (N_15001,N_14713,N_14530);
and U15002 (N_15002,N_14274,N_14888);
nor U15003 (N_15003,N_14796,N_14664);
nand U15004 (N_15004,N_14181,N_14495);
nand U15005 (N_15005,N_14071,N_14716);
nor U15006 (N_15006,N_14051,N_14761);
nand U15007 (N_15007,N_14203,N_14421);
or U15008 (N_15008,N_14344,N_14848);
nand U15009 (N_15009,N_14657,N_14013);
nand U15010 (N_15010,N_14210,N_14041);
xnor U15011 (N_15011,N_14944,N_14454);
xnor U15012 (N_15012,N_14624,N_14538);
or U15013 (N_15013,N_14650,N_14149);
xor U15014 (N_15014,N_14705,N_14262);
nand U15015 (N_15015,N_14593,N_14570);
xor U15016 (N_15016,N_14609,N_14161);
xor U15017 (N_15017,N_14438,N_14197);
xor U15018 (N_15018,N_14244,N_14045);
nand U15019 (N_15019,N_14623,N_14924);
nand U15020 (N_15020,N_14837,N_14594);
xor U15021 (N_15021,N_14672,N_14114);
and U15022 (N_15022,N_14878,N_14376);
and U15023 (N_15023,N_14010,N_14330);
nand U15024 (N_15024,N_14760,N_14007);
nand U15025 (N_15025,N_14963,N_14622);
and U15026 (N_15026,N_14771,N_14112);
or U15027 (N_15027,N_14939,N_14946);
nor U15028 (N_15028,N_14332,N_14909);
and U15029 (N_15029,N_14659,N_14397);
and U15030 (N_15030,N_14847,N_14224);
nand U15031 (N_15031,N_14971,N_14882);
and U15032 (N_15032,N_14876,N_14074);
nor U15033 (N_15033,N_14829,N_14626);
and U15034 (N_15034,N_14868,N_14465);
nand U15035 (N_15035,N_14490,N_14961);
xnor U15036 (N_15036,N_14702,N_14700);
nor U15037 (N_15037,N_14663,N_14922);
or U15038 (N_15038,N_14335,N_14742);
or U15039 (N_15039,N_14388,N_14870);
nand U15040 (N_15040,N_14245,N_14549);
or U15041 (N_15041,N_14604,N_14461);
nand U15042 (N_15042,N_14865,N_14102);
and U15043 (N_15043,N_14562,N_14240);
or U15044 (N_15044,N_14903,N_14118);
and U15045 (N_15045,N_14757,N_14524);
or U15046 (N_15046,N_14030,N_14838);
and U15047 (N_15047,N_14543,N_14690);
xnor U15048 (N_15048,N_14751,N_14456);
or U15049 (N_15049,N_14853,N_14644);
xnor U15050 (N_15050,N_14960,N_14859);
nor U15051 (N_15051,N_14890,N_14046);
or U15052 (N_15052,N_14320,N_14239);
xnor U15053 (N_15053,N_14318,N_14028);
xnor U15054 (N_15054,N_14250,N_14762);
and U15055 (N_15055,N_14364,N_14616);
nand U15056 (N_15056,N_14347,N_14380);
nor U15057 (N_15057,N_14085,N_14297);
nand U15058 (N_15058,N_14133,N_14015);
nor U15059 (N_15059,N_14532,N_14775);
nand U15060 (N_15060,N_14576,N_14354);
nand U15061 (N_15061,N_14415,N_14135);
nand U15062 (N_15062,N_14111,N_14730);
and U15063 (N_15063,N_14810,N_14787);
or U15064 (N_15064,N_14029,N_14062);
xor U15065 (N_15065,N_14034,N_14639);
or U15066 (N_15066,N_14492,N_14993);
xnor U15067 (N_15067,N_14917,N_14405);
nand U15068 (N_15068,N_14166,N_14381);
and U15069 (N_15069,N_14324,N_14568);
or U15070 (N_15070,N_14601,N_14485);
or U15071 (N_15071,N_14989,N_14432);
nor U15072 (N_15072,N_14575,N_14143);
and U15073 (N_15073,N_14969,N_14247);
nor U15074 (N_15074,N_14186,N_14583);
and U15075 (N_15075,N_14764,N_14795);
and U15076 (N_15076,N_14752,N_14906);
xor U15077 (N_15077,N_14152,N_14833);
or U15078 (N_15078,N_14400,N_14175);
or U15079 (N_15079,N_14450,N_14280);
xnor U15080 (N_15080,N_14005,N_14695);
xor U15081 (N_15081,N_14926,N_14942);
and U15082 (N_15082,N_14130,N_14475);
or U15083 (N_15083,N_14464,N_14264);
and U15084 (N_15084,N_14208,N_14800);
nand U15085 (N_15085,N_14872,N_14086);
nor U15086 (N_15086,N_14978,N_14393);
xnor U15087 (N_15087,N_14653,N_14977);
nand U15088 (N_15088,N_14372,N_14692);
and U15089 (N_15089,N_14647,N_14371);
and U15090 (N_15090,N_14723,N_14610);
xor U15091 (N_15091,N_14706,N_14444);
nand U15092 (N_15092,N_14957,N_14841);
and U15093 (N_15093,N_14417,N_14083);
or U15094 (N_15094,N_14539,N_14769);
xnor U15095 (N_15095,N_14355,N_14056);
xor U15096 (N_15096,N_14548,N_14377);
and U15097 (N_15097,N_14325,N_14476);
nor U15098 (N_15098,N_14044,N_14763);
nor U15099 (N_15099,N_14555,N_14899);
xor U15100 (N_15100,N_14719,N_14814);
or U15101 (N_15101,N_14823,N_14357);
xor U15102 (N_15102,N_14003,N_14246);
and U15103 (N_15103,N_14714,N_14098);
xnor U15104 (N_15104,N_14067,N_14195);
xor U15105 (N_15105,N_14501,N_14423);
and U15106 (N_15106,N_14749,N_14808);
and U15107 (N_15107,N_14687,N_14361);
nand U15108 (N_15108,N_14852,N_14670);
nand U15109 (N_15109,N_14498,N_14304);
or U15110 (N_15110,N_14504,N_14923);
nor U15111 (N_15111,N_14669,N_14807);
and U15112 (N_15112,N_14054,N_14835);
nand U15113 (N_15113,N_14370,N_14039);
and U15114 (N_15114,N_14430,N_14140);
and U15115 (N_15115,N_14386,N_14907);
nand U15116 (N_15116,N_14571,N_14614);
or U15117 (N_15117,N_14011,N_14235);
or U15118 (N_15118,N_14937,N_14840);
nand U15119 (N_15119,N_14493,N_14455);
nand U15120 (N_15120,N_14665,N_14266);
and U15121 (N_15121,N_14980,N_14373);
or U15122 (N_15122,N_14612,N_14349);
nor U15123 (N_15123,N_14685,N_14411);
nand U15124 (N_15124,N_14126,N_14927);
and U15125 (N_15125,N_14179,N_14517);
or U15126 (N_15126,N_14252,N_14592);
and U15127 (N_15127,N_14103,N_14230);
xor U15128 (N_15128,N_14082,N_14748);
or U15129 (N_15129,N_14368,N_14962);
nor U15130 (N_15130,N_14484,N_14259);
and U15131 (N_15131,N_14299,N_14394);
and U15132 (N_15132,N_14613,N_14791);
or U15133 (N_15133,N_14422,N_14919);
nor U15134 (N_15134,N_14611,N_14064);
and U15135 (N_15135,N_14414,N_14910);
xor U15136 (N_15136,N_14273,N_14667);
or U15137 (N_15137,N_14597,N_14819);
xor U15138 (N_15138,N_14968,N_14319);
and U15139 (N_15139,N_14774,N_14228);
and U15140 (N_15140,N_14879,N_14912);
xor U15141 (N_15141,N_14416,N_14811);
nor U15142 (N_15142,N_14300,N_14173);
or U15143 (N_15143,N_14871,N_14633);
or U15144 (N_15144,N_14435,N_14383);
or U15145 (N_15145,N_14312,N_14269);
or U15146 (N_15146,N_14891,N_14309);
nand U15147 (N_15147,N_14251,N_14880);
nor U15148 (N_15148,N_14217,N_14518);
and U15149 (N_15149,N_14164,N_14732);
xor U15150 (N_15150,N_14204,N_14905);
nand U15151 (N_15151,N_14092,N_14385);
nand U15152 (N_15152,N_14487,N_14141);
and U15153 (N_15153,N_14467,N_14825);
and U15154 (N_15154,N_14231,N_14654);
and U15155 (N_15155,N_14897,N_14359);
xor U15156 (N_15156,N_14177,N_14873);
nand U15157 (N_15157,N_14241,N_14452);
nand U15158 (N_15158,N_14901,N_14027);
nor U15159 (N_15159,N_14268,N_14638);
or U15160 (N_15160,N_14012,N_14754);
and U15161 (N_15161,N_14463,N_14983);
or U15162 (N_15162,N_14060,N_14786);
xor U15163 (N_15163,N_14818,N_14689);
nor U15164 (N_15164,N_14079,N_14059);
or U15165 (N_15165,N_14733,N_14686);
and U15166 (N_15166,N_14780,N_14794);
nand U15167 (N_15167,N_14914,N_14600);
nor U15168 (N_15168,N_14488,N_14651);
nand U15169 (N_15169,N_14401,N_14860);
nand U15170 (N_15170,N_14147,N_14328);
or U15171 (N_15171,N_14781,N_14360);
nand U15172 (N_15172,N_14547,N_14916);
nor U15173 (N_15173,N_14929,N_14322);
and U15174 (N_15174,N_14342,N_14499);
xnor U15175 (N_15175,N_14420,N_14567);
nor U15176 (N_15176,N_14643,N_14132);
nand U15177 (N_15177,N_14122,N_14243);
xnor U15178 (N_15178,N_14680,N_14374);
xor U15179 (N_15179,N_14406,N_14995);
xnor U15180 (N_15180,N_14256,N_14874);
and U15181 (N_15181,N_14947,N_14174);
nand U15182 (N_15182,N_14974,N_14693);
nor U15183 (N_15183,N_14785,N_14998);
or U15184 (N_15184,N_14694,N_14001);
nor U15185 (N_15185,N_14207,N_14471);
xor U15186 (N_15186,N_14019,N_14316);
and U15187 (N_15187,N_14075,N_14821);
nor U15188 (N_15188,N_14788,N_14271);
nor U15189 (N_15189,N_14031,N_14088);
nor U15190 (N_15190,N_14527,N_14681);
and U15191 (N_15191,N_14768,N_14094);
and U15192 (N_15192,N_14709,N_14233);
and U15193 (N_15193,N_14218,N_14213);
nand U15194 (N_15194,N_14072,N_14267);
or U15195 (N_15195,N_14148,N_14817);
or U15196 (N_15196,N_14589,N_14893);
nand U15197 (N_15197,N_14525,N_14073);
xnor U15198 (N_15198,N_14286,N_14790);
nor U15199 (N_15199,N_14261,N_14341);
xnor U15200 (N_15200,N_14433,N_14199);
nand U15201 (N_15201,N_14100,N_14707);
xor U15202 (N_15202,N_14289,N_14620);
nand U15203 (N_15203,N_14295,N_14820);
nand U15204 (N_15204,N_14290,N_14497);
or U15205 (N_15205,N_14223,N_14982);
nand U15206 (N_15206,N_14541,N_14949);
or U15207 (N_15207,N_14187,N_14955);
nor U15208 (N_15208,N_14718,N_14281);
xor U15209 (N_15209,N_14509,N_14183);
and U15210 (N_15210,N_14738,N_14196);
or U15211 (N_15211,N_14249,N_14201);
nand U15212 (N_15212,N_14745,N_14991);
and U15213 (N_15213,N_14529,N_14336);
xor U15214 (N_15214,N_14607,N_14911);
or U15215 (N_15215,N_14999,N_14482);
or U15216 (N_15216,N_14194,N_14744);
and U15217 (N_15217,N_14737,N_14329);
or U15218 (N_15218,N_14120,N_14782);
nor U15219 (N_15219,N_14503,N_14163);
nand U15220 (N_15220,N_14678,N_14512);
or U15221 (N_15221,N_14367,N_14779);
xnor U15222 (N_15222,N_14629,N_14282);
and U15223 (N_15223,N_14353,N_14331);
or U15224 (N_15224,N_14699,N_14778);
xor U15225 (N_15225,N_14468,N_14026);
nor U15226 (N_15226,N_14717,N_14887);
xor U15227 (N_15227,N_14958,N_14598);
nand U15228 (N_15228,N_14439,N_14660);
nand U15229 (N_15229,N_14984,N_14996);
and U15230 (N_15230,N_14864,N_14496);
xnor U15231 (N_15231,N_14976,N_14154);
and U15232 (N_15232,N_14069,N_14954);
or U15233 (N_15233,N_14153,N_14544);
nor U15234 (N_15234,N_14540,N_14018);
nand U15235 (N_15235,N_14478,N_14459);
nor U15236 (N_15236,N_14824,N_14915);
nand U15237 (N_15237,N_14317,N_14508);
and U15238 (N_15238,N_14750,N_14193);
nand U15239 (N_15239,N_14580,N_14953);
and U15240 (N_15240,N_14124,N_14108);
or U15241 (N_15241,N_14125,N_14830);
or U15242 (N_15242,N_14588,N_14429);
and U15243 (N_15243,N_14158,N_14107);
xor U15244 (N_15244,N_14747,N_14628);
nor U15245 (N_15245,N_14849,N_14908);
or U15246 (N_15246,N_14520,N_14418);
or U15247 (N_15247,N_14936,N_14697);
nor U15248 (N_15248,N_14608,N_14565);
xnor U15249 (N_15249,N_14635,N_14987);
nor U15250 (N_15250,N_14146,N_14284);
nor U15251 (N_15251,N_14867,N_14586);
or U15252 (N_15252,N_14646,N_14425);
nor U15253 (N_15253,N_14673,N_14144);
nor U15254 (N_15254,N_14232,N_14602);
or U15255 (N_15255,N_14581,N_14077);
xnor U15256 (N_15256,N_14057,N_14428);
nor U15257 (N_15257,N_14945,N_14225);
nor U15258 (N_15258,N_14449,N_14850);
or U15259 (N_15259,N_14921,N_14988);
or U15260 (N_15260,N_14533,N_14831);
nor U15261 (N_15261,N_14469,N_14701);
and U15262 (N_15262,N_14630,N_14772);
nor U15263 (N_15263,N_14605,N_14137);
or U15264 (N_15264,N_14410,N_14311);
and U15265 (N_15265,N_14227,N_14753);
nor U15266 (N_15266,N_14739,N_14352);
nor U15267 (N_15267,N_14343,N_14515);
or U15268 (N_15268,N_14812,N_14229);
nor U15269 (N_15269,N_14260,N_14279);
nor U15270 (N_15270,N_14827,N_14389);
or U15271 (N_15271,N_14710,N_14139);
or U15272 (N_15272,N_14740,N_14104);
nor U15273 (N_15273,N_14448,N_14479);
and U15274 (N_15274,N_14301,N_14313);
nand U15275 (N_15275,N_14662,N_14185);
and U15276 (N_15276,N_14815,N_14641);
xnor U15277 (N_15277,N_14572,N_14399);
xnor U15278 (N_15278,N_14160,N_14097);
and U15279 (N_15279,N_14885,N_14065);
and U15280 (N_15280,N_14023,N_14728);
nand U15281 (N_15281,N_14558,N_14105);
nor U15282 (N_15282,N_14668,N_14883);
nor U15283 (N_15283,N_14191,N_14677);
nor U15284 (N_15284,N_14434,N_14315);
and U15285 (N_15285,N_14959,N_14258);
or U15286 (N_15286,N_14507,N_14894);
nand U15287 (N_15287,N_14306,N_14395);
xor U15288 (N_15288,N_14436,N_14783);
nor U15289 (N_15289,N_14789,N_14656);
and U15290 (N_15290,N_14390,N_14755);
and U15291 (N_15291,N_14648,N_14992);
xnor U15292 (N_15292,N_14291,N_14460);
and U15293 (N_15293,N_14123,N_14006);
or U15294 (N_15294,N_14895,N_14032);
xnor U15295 (N_15295,N_14595,N_14408);
or U15296 (N_15296,N_14806,N_14084);
nand U15297 (N_15297,N_14986,N_14138);
nand U15298 (N_15298,N_14283,N_14952);
xor U15299 (N_15299,N_14440,N_14720);
nor U15300 (N_15300,N_14024,N_14546);
nand U15301 (N_15301,N_14106,N_14658);
nor U15302 (N_15302,N_14159,N_14263);
xnor U15303 (N_15303,N_14900,N_14254);
nand U15304 (N_15304,N_14021,N_14404);
or U15305 (N_15305,N_14542,N_14803);
xnor U15306 (N_15306,N_14366,N_14171);
xnor U15307 (N_15307,N_14834,N_14938);
nor U15308 (N_15308,N_14169,N_14902);
or U15309 (N_15309,N_14134,N_14997);
or U15310 (N_15310,N_14222,N_14211);
or U15311 (N_15311,N_14127,N_14550);
xor U15312 (N_15312,N_14632,N_14564);
and U15313 (N_15313,N_14113,N_14898);
nand U15314 (N_15314,N_14047,N_14861);
xnor U15315 (N_15315,N_14877,N_14334);
nand U15316 (N_15316,N_14000,N_14676);
and U15317 (N_15317,N_14513,N_14407);
nor U15318 (N_15318,N_14008,N_14928);
nand U15319 (N_15319,N_14151,N_14930);
or U15320 (N_15320,N_14042,N_14270);
nor U15321 (N_15321,N_14866,N_14275);
nand U15322 (N_15322,N_14292,N_14688);
nor U15323 (N_15323,N_14721,N_14426);
or U15324 (N_15324,N_14666,N_14587);
xnor U15325 (N_15325,N_14698,N_14150);
xor U15326 (N_15326,N_14110,N_14813);
xor U15327 (N_15327,N_14458,N_14724);
and U15328 (N_15328,N_14531,N_14809);
nor U15329 (N_15329,N_14474,N_14981);
or U15330 (N_15330,N_14964,N_14337);
nand U15331 (N_15331,N_14486,N_14551);
xnor U15332 (N_15332,N_14087,N_14040);
nand U15333 (N_15333,N_14759,N_14766);
or U15334 (N_15334,N_14345,N_14875);
xnor U15335 (N_15335,N_14350,N_14131);
and U15336 (N_15336,N_14178,N_14055);
or U15337 (N_15337,N_14682,N_14384);
or U15338 (N_15338,N_14053,N_14726);
and U15339 (N_15339,N_14119,N_14574);
or U15340 (N_15340,N_14855,N_14773);
xor U15341 (N_15341,N_14093,N_14462);
nand U15342 (N_15342,N_14365,N_14437);
nor U15343 (N_15343,N_14424,N_14396);
and U15344 (N_15344,N_14128,N_14577);
xor U15345 (N_15345,N_14842,N_14172);
xnor U15346 (N_15346,N_14037,N_14526);
and U15347 (N_15347,N_14591,N_14226);
nand U15348 (N_15348,N_14886,N_14985);
xor U15349 (N_15349,N_14048,N_14277);
xor U15350 (N_15350,N_14216,N_14884);
and U15351 (N_15351,N_14606,N_14711);
or U15352 (N_15352,N_14704,N_14188);
or U15353 (N_15353,N_14634,N_14826);
or U15354 (N_15354,N_14238,N_14050);
nor U15355 (N_15355,N_14115,N_14802);
xor U15356 (N_15356,N_14070,N_14298);
or U15357 (N_15357,N_14722,N_14801);
and U15358 (N_15358,N_14180,N_14451);
nand U15359 (N_15359,N_14058,N_14409);
or U15360 (N_15360,N_14176,N_14036);
or U15361 (N_15361,N_14348,N_14412);
xor U15362 (N_15362,N_14950,N_14303);
nor U15363 (N_15363,N_14441,N_14913);
nor U15364 (N_15364,N_14637,N_14844);
xnor U15365 (N_15365,N_14038,N_14965);
or U15366 (N_15366,N_14285,N_14889);
nor U15367 (N_15367,N_14323,N_14379);
and U15368 (N_15368,N_14091,N_14655);
or U15369 (N_15369,N_14804,N_14170);
xnor U15370 (N_15370,N_14703,N_14559);
and U15371 (N_15371,N_14052,N_14453);
and U15372 (N_15372,N_14973,N_14473);
and U15373 (N_15373,N_14061,N_14477);
and U15374 (N_15374,N_14202,N_14743);
and U15375 (N_15375,N_14002,N_14142);
xnor U15376 (N_15376,N_14155,N_14967);
nand U15377 (N_15377,N_14502,N_14552);
and U15378 (N_15378,N_14931,N_14675);
xor U15379 (N_15379,N_14481,N_14470);
nor U15380 (N_15380,N_14579,N_14242);
or U15381 (N_15381,N_14727,N_14619);
nand U15382 (N_15382,N_14734,N_14767);
xor U15383 (N_15383,N_14234,N_14640);
or U15384 (N_15384,N_14362,N_14265);
nor U15385 (N_15385,N_14972,N_14198);
xor U15386 (N_15386,N_14480,N_14272);
or U15387 (N_15387,N_14095,N_14956);
xnor U15388 (N_15388,N_14190,N_14636);
or U15389 (N_15389,N_14136,N_14934);
nor U15390 (N_15390,N_14979,N_14340);
or U15391 (N_15391,N_14708,N_14212);
nand U15392 (N_15392,N_14712,N_14863);
xor U15393 (N_15393,N_14661,N_14096);
nor U15394 (N_15394,N_14975,N_14798);
xor U15395 (N_15395,N_14472,N_14221);
nand U15396 (N_15396,N_14278,N_14033);
xor U15397 (N_15397,N_14049,N_14896);
nor U15398 (N_15398,N_14584,N_14683);
nand U15399 (N_15399,N_14854,N_14741);
and U15400 (N_15400,N_14016,N_14206);
xnor U15401 (N_15401,N_14553,N_14326);
xor U15402 (N_15402,N_14725,N_14932);
or U15403 (N_15403,N_14145,N_14519);
nand U15404 (N_15404,N_14182,N_14398);
nor U15405 (N_15405,N_14603,N_14510);
xnor U15406 (N_15406,N_14736,N_14523);
or U15407 (N_15407,N_14522,N_14925);
xnor U15408 (N_15408,N_14904,N_14020);
xnor U15409 (N_15409,N_14856,N_14797);
xor U15410 (N_15410,N_14514,N_14715);
and U15411 (N_15411,N_14892,N_14220);
nand U15412 (N_15412,N_14684,N_14446);
and U15413 (N_15413,N_14382,N_14516);
nand U15414 (N_15414,N_14560,N_14729);
or U15415 (N_15415,N_14920,N_14255);
and U15416 (N_15416,N_14427,N_14731);
nor U15417 (N_15417,N_14535,N_14288);
nand U15418 (N_15418,N_14066,N_14165);
or U15419 (N_15419,N_14537,N_14287);
or U15420 (N_15420,N_14935,N_14117);
xnor U15421 (N_15421,N_14009,N_14735);
and U15422 (N_15422,N_14671,N_14157);
xnor U15423 (N_15423,N_14257,N_14184);
xnor U15424 (N_15424,N_14068,N_14792);
nor U15425 (N_15425,N_14746,N_14836);
and U15426 (N_15426,N_14858,N_14770);
and U15427 (N_15427,N_14491,N_14189);
and U15428 (N_15428,N_14839,N_14489);
or U15429 (N_15429,N_14599,N_14308);
nor U15430 (N_15430,N_14310,N_14391);
or U15431 (N_15431,N_14327,N_14442);
xor U15432 (N_15432,N_14582,N_14443);
nand U15433 (N_15433,N_14990,N_14200);
xor U15434 (N_15434,N_14305,N_14578);
xor U15435 (N_15435,N_14500,N_14799);
xor U15436 (N_15436,N_14642,N_14691);
nand U15437 (N_15437,N_14109,N_14294);
and U15438 (N_15438,N_14116,N_14918);
and U15439 (N_15439,N_14017,N_14078);
and U15440 (N_15440,N_14043,N_14941);
xor U15441 (N_15441,N_14022,N_14413);
or U15442 (N_15442,N_14561,N_14556);
and U15443 (N_15443,N_14756,N_14276);
or U15444 (N_15444,N_14994,N_14948);
nand U15445 (N_15445,N_14063,N_14805);
or U15446 (N_15446,N_14076,N_14090);
xnor U15447 (N_15447,N_14403,N_14346);
nor U15448 (N_15448,N_14793,N_14205);
and U15449 (N_15449,N_14156,N_14765);
xnor U15450 (N_15450,N_14832,N_14563);
nand U15451 (N_15451,N_14121,N_14828);
and U15452 (N_15452,N_14862,N_14339);
nand U15453 (N_15453,N_14679,N_14943);
and U15454 (N_15454,N_14356,N_14857);
nand U15455 (N_15455,N_14569,N_14025);
nor U15456 (N_15456,N_14696,N_14375);
nor U15457 (N_15457,N_14387,N_14521);
nor U15458 (N_15458,N_14253,N_14214);
nor U15459 (N_15459,N_14618,N_14966);
or U15460 (N_15460,N_14392,N_14004);
xnor U15461 (N_15461,N_14236,N_14099);
or U15462 (N_15462,N_14419,N_14296);
nor U15463 (N_15463,N_14585,N_14363);
nand U15464 (N_15464,N_14940,N_14843);
nand U15465 (N_15465,N_14447,N_14080);
nand U15466 (N_15466,N_14645,N_14162);
xnor U15467 (N_15467,N_14621,N_14557);
nand U15468 (N_15468,N_14483,N_14505);
or U15469 (N_15469,N_14192,N_14237);
xor U15470 (N_15470,N_14528,N_14615);
xor U15471 (N_15471,N_14378,N_14307);
nand U15472 (N_15472,N_14293,N_14369);
nand U15473 (N_15473,N_14554,N_14776);
or U15474 (N_15474,N_14573,N_14466);
or U15475 (N_15475,N_14351,N_14089);
and U15476 (N_15476,N_14219,N_14566);
nand U15477 (N_15477,N_14101,N_14402);
and U15478 (N_15478,N_14215,N_14777);
nand U15479 (N_15479,N_14822,N_14511);
and U15480 (N_15480,N_14445,N_14881);
xnor U15481 (N_15481,N_14970,N_14758);
and U15482 (N_15482,N_14816,N_14845);
and U15483 (N_15483,N_14333,N_14617);
xor U15484 (N_15484,N_14631,N_14129);
xor U15485 (N_15485,N_14851,N_14248);
and U15486 (N_15486,N_14506,N_14035);
or U15487 (N_15487,N_14869,N_14933);
or U15488 (N_15488,N_14846,N_14209);
and U15489 (N_15489,N_14457,N_14596);
nor U15490 (N_15490,N_14314,N_14494);
nand U15491 (N_15491,N_14534,N_14168);
or U15492 (N_15492,N_14302,N_14358);
nand U15493 (N_15493,N_14627,N_14167);
or U15494 (N_15494,N_14338,N_14649);
or U15495 (N_15495,N_14545,N_14431);
nand U15496 (N_15496,N_14014,N_14784);
nand U15497 (N_15497,N_14321,N_14536);
or U15498 (N_15498,N_14625,N_14951);
and U15499 (N_15499,N_14081,N_14590);
xor U15500 (N_15500,N_14080,N_14091);
xnor U15501 (N_15501,N_14482,N_14111);
xor U15502 (N_15502,N_14962,N_14642);
and U15503 (N_15503,N_14853,N_14429);
nand U15504 (N_15504,N_14101,N_14155);
and U15505 (N_15505,N_14188,N_14062);
or U15506 (N_15506,N_14522,N_14918);
or U15507 (N_15507,N_14521,N_14841);
and U15508 (N_15508,N_14828,N_14653);
nand U15509 (N_15509,N_14286,N_14492);
and U15510 (N_15510,N_14844,N_14019);
nand U15511 (N_15511,N_14048,N_14808);
nand U15512 (N_15512,N_14272,N_14777);
nand U15513 (N_15513,N_14612,N_14905);
nor U15514 (N_15514,N_14022,N_14377);
xor U15515 (N_15515,N_14828,N_14153);
nand U15516 (N_15516,N_14883,N_14525);
xnor U15517 (N_15517,N_14212,N_14133);
or U15518 (N_15518,N_14775,N_14226);
nand U15519 (N_15519,N_14427,N_14534);
nor U15520 (N_15520,N_14906,N_14078);
and U15521 (N_15521,N_14487,N_14976);
and U15522 (N_15522,N_14820,N_14572);
or U15523 (N_15523,N_14532,N_14438);
or U15524 (N_15524,N_14237,N_14827);
or U15525 (N_15525,N_14545,N_14211);
nor U15526 (N_15526,N_14876,N_14273);
and U15527 (N_15527,N_14815,N_14919);
nand U15528 (N_15528,N_14225,N_14422);
or U15529 (N_15529,N_14914,N_14976);
and U15530 (N_15530,N_14407,N_14308);
nand U15531 (N_15531,N_14205,N_14832);
nor U15532 (N_15532,N_14071,N_14839);
and U15533 (N_15533,N_14492,N_14774);
or U15534 (N_15534,N_14649,N_14946);
xnor U15535 (N_15535,N_14298,N_14419);
nand U15536 (N_15536,N_14263,N_14652);
nand U15537 (N_15537,N_14860,N_14962);
nand U15538 (N_15538,N_14375,N_14360);
xor U15539 (N_15539,N_14344,N_14091);
nor U15540 (N_15540,N_14396,N_14389);
and U15541 (N_15541,N_14400,N_14892);
or U15542 (N_15542,N_14084,N_14194);
xor U15543 (N_15543,N_14268,N_14728);
nand U15544 (N_15544,N_14493,N_14740);
nor U15545 (N_15545,N_14296,N_14565);
xnor U15546 (N_15546,N_14639,N_14755);
nand U15547 (N_15547,N_14992,N_14084);
nand U15548 (N_15548,N_14743,N_14629);
nand U15549 (N_15549,N_14624,N_14508);
nand U15550 (N_15550,N_14322,N_14964);
or U15551 (N_15551,N_14517,N_14047);
nor U15552 (N_15552,N_14842,N_14924);
and U15553 (N_15553,N_14166,N_14259);
xor U15554 (N_15554,N_14726,N_14603);
nor U15555 (N_15555,N_14004,N_14759);
or U15556 (N_15556,N_14895,N_14711);
nor U15557 (N_15557,N_14873,N_14386);
xnor U15558 (N_15558,N_14904,N_14849);
and U15559 (N_15559,N_14297,N_14971);
or U15560 (N_15560,N_14067,N_14037);
xor U15561 (N_15561,N_14061,N_14700);
and U15562 (N_15562,N_14465,N_14350);
xnor U15563 (N_15563,N_14561,N_14229);
and U15564 (N_15564,N_14137,N_14076);
nor U15565 (N_15565,N_14660,N_14885);
and U15566 (N_15566,N_14254,N_14890);
nor U15567 (N_15567,N_14494,N_14056);
or U15568 (N_15568,N_14736,N_14083);
nor U15569 (N_15569,N_14924,N_14558);
nand U15570 (N_15570,N_14301,N_14596);
and U15571 (N_15571,N_14367,N_14845);
nor U15572 (N_15572,N_14108,N_14504);
nor U15573 (N_15573,N_14150,N_14493);
or U15574 (N_15574,N_14541,N_14290);
or U15575 (N_15575,N_14817,N_14564);
nand U15576 (N_15576,N_14795,N_14747);
nor U15577 (N_15577,N_14858,N_14496);
nor U15578 (N_15578,N_14211,N_14072);
and U15579 (N_15579,N_14909,N_14710);
xor U15580 (N_15580,N_14705,N_14501);
nor U15581 (N_15581,N_14141,N_14563);
and U15582 (N_15582,N_14731,N_14317);
nor U15583 (N_15583,N_14976,N_14308);
xnor U15584 (N_15584,N_14672,N_14392);
nor U15585 (N_15585,N_14629,N_14156);
nor U15586 (N_15586,N_14352,N_14807);
nor U15587 (N_15587,N_14848,N_14601);
or U15588 (N_15588,N_14961,N_14581);
xor U15589 (N_15589,N_14561,N_14828);
nor U15590 (N_15590,N_14348,N_14227);
xnor U15591 (N_15591,N_14575,N_14739);
nand U15592 (N_15592,N_14387,N_14300);
nor U15593 (N_15593,N_14781,N_14595);
nand U15594 (N_15594,N_14708,N_14185);
nor U15595 (N_15595,N_14244,N_14933);
nand U15596 (N_15596,N_14208,N_14825);
and U15597 (N_15597,N_14064,N_14841);
nor U15598 (N_15598,N_14948,N_14969);
xnor U15599 (N_15599,N_14064,N_14284);
nand U15600 (N_15600,N_14697,N_14055);
xor U15601 (N_15601,N_14991,N_14035);
nor U15602 (N_15602,N_14201,N_14768);
xnor U15603 (N_15603,N_14282,N_14726);
xor U15604 (N_15604,N_14729,N_14481);
nor U15605 (N_15605,N_14047,N_14851);
xor U15606 (N_15606,N_14132,N_14746);
nor U15607 (N_15607,N_14650,N_14672);
nand U15608 (N_15608,N_14564,N_14681);
xnor U15609 (N_15609,N_14575,N_14256);
or U15610 (N_15610,N_14690,N_14880);
nor U15611 (N_15611,N_14486,N_14344);
xor U15612 (N_15612,N_14982,N_14172);
nor U15613 (N_15613,N_14501,N_14688);
and U15614 (N_15614,N_14396,N_14742);
and U15615 (N_15615,N_14260,N_14887);
nor U15616 (N_15616,N_14425,N_14699);
xor U15617 (N_15617,N_14153,N_14714);
and U15618 (N_15618,N_14187,N_14567);
and U15619 (N_15619,N_14516,N_14311);
or U15620 (N_15620,N_14014,N_14585);
xor U15621 (N_15621,N_14130,N_14965);
nand U15622 (N_15622,N_14001,N_14166);
nand U15623 (N_15623,N_14994,N_14951);
nor U15624 (N_15624,N_14721,N_14341);
nor U15625 (N_15625,N_14723,N_14375);
nor U15626 (N_15626,N_14717,N_14611);
and U15627 (N_15627,N_14721,N_14207);
or U15628 (N_15628,N_14030,N_14344);
nand U15629 (N_15629,N_14304,N_14976);
nand U15630 (N_15630,N_14491,N_14525);
nor U15631 (N_15631,N_14040,N_14845);
nor U15632 (N_15632,N_14571,N_14565);
nand U15633 (N_15633,N_14020,N_14869);
nand U15634 (N_15634,N_14640,N_14385);
nand U15635 (N_15635,N_14963,N_14497);
nor U15636 (N_15636,N_14068,N_14425);
or U15637 (N_15637,N_14973,N_14202);
and U15638 (N_15638,N_14833,N_14113);
nand U15639 (N_15639,N_14289,N_14078);
and U15640 (N_15640,N_14233,N_14653);
and U15641 (N_15641,N_14175,N_14872);
nand U15642 (N_15642,N_14908,N_14411);
or U15643 (N_15643,N_14095,N_14057);
and U15644 (N_15644,N_14296,N_14607);
xnor U15645 (N_15645,N_14303,N_14582);
nand U15646 (N_15646,N_14148,N_14558);
and U15647 (N_15647,N_14092,N_14289);
nor U15648 (N_15648,N_14112,N_14166);
xor U15649 (N_15649,N_14830,N_14391);
nand U15650 (N_15650,N_14221,N_14656);
nand U15651 (N_15651,N_14667,N_14712);
and U15652 (N_15652,N_14056,N_14270);
and U15653 (N_15653,N_14862,N_14643);
nand U15654 (N_15654,N_14575,N_14371);
nand U15655 (N_15655,N_14344,N_14929);
nor U15656 (N_15656,N_14104,N_14006);
xnor U15657 (N_15657,N_14758,N_14364);
xnor U15658 (N_15658,N_14869,N_14085);
or U15659 (N_15659,N_14642,N_14057);
or U15660 (N_15660,N_14461,N_14613);
nor U15661 (N_15661,N_14489,N_14186);
and U15662 (N_15662,N_14876,N_14194);
nor U15663 (N_15663,N_14800,N_14252);
or U15664 (N_15664,N_14026,N_14318);
nand U15665 (N_15665,N_14385,N_14205);
and U15666 (N_15666,N_14489,N_14886);
or U15667 (N_15667,N_14463,N_14854);
nand U15668 (N_15668,N_14681,N_14654);
nor U15669 (N_15669,N_14438,N_14831);
nand U15670 (N_15670,N_14346,N_14696);
nor U15671 (N_15671,N_14888,N_14342);
or U15672 (N_15672,N_14043,N_14361);
or U15673 (N_15673,N_14732,N_14192);
or U15674 (N_15674,N_14939,N_14812);
or U15675 (N_15675,N_14734,N_14472);
or U15676 (N_15676,N_14340,N_14070);
nand U15677 (N_15677,N_14121,N_14114);
or U15678 (N_15678,N_14098,N_14704);
and U15679 (N_15679,N_14301,N_14776);
nand U15680 (N_15680,N_14834,N_14205);
and U15681 (N_15681,N_14758,N_14630);
and U15682 (N_15682,N_14145,N_14582);
or U15683 (N_15683,N_14553,N_14857);
and U15684 (N_15684,N_14205,N_14083);
nand U15685 (N_15685,N_14483,N_14902);
nor U15686 (N_15686,N_14539,N_14540);
nand U15687 (N_15687,N_14471,N_14429);
and U15688 (N_15688,N_14438,N_14717);
xnor U15689 (N_15689,N_14434,N_14317);
and U15690 (N_15690,N_14400,N_14487);
nor U15691 (N_15691,N_14063,N_14032);
and U15692 (N_15692,N_14443,N_14054);
nand U15693 (N_15693,N_14833,N_14751);
nor U15694 (N_15694,N_14791,N_14324);
nor U15695 (N_15695,N_14924,N_14085);
nor U15696 (N_15696,N_14489,N_14470);
and U15697 (N_15697,N_14403,N_14702);
or U15698 (N_15698,N_14832,N_14062);
nor U15699 (N_15699,N_14784,N_14681);
nand U15700 (N_15700,N_14528,N_14420);
nor U15701 (N_15701,N_14625,N_14404);
and U15702 (N_15702,N_14022,N_14368);
nand U15703 (N_15703,N_14707,N_14061);
or U15704 (N_15704,N_14224,N_14998);
nor U15705 (N_15705,N_14096,N_14663);
xnor U15706 (N_15706,N_14257,N_14270);
or U15707 (N_15707,N_14396,N_14978);
and U15708 (N_15708,N_14434,N_14552);
or U15709 (N_15709,N_14884,N_14056);
nand U15710 (N_15710,N_14539,N_14497);
or U15711 (N_15711,N_14131,N_14590);
xnor U15712 (N_15712,N_14155,N_14457);
and U15713 (N_15713,N_14398,N_14647);
nor U15714 (N_15714,N_14734,N_14553);
and U15715 (N_15715,N_14356,N_14049);
or U15716 (N_15716,N_14398,N_14765);
xnor U15717 (N_15717,N_14826,N_14181);
xor U15718 (N_15718,N_14107,N_14091);
and U15719 (N_15719,N_14352,N_14852);
nand U15720 (N_15720,N_14113,N_14860);
xnor U15721 (N_15721,N_14406,N_14861);
and U15722 (N_15722,N_14301,N_14178);
or U15723 (N_15723,N_14824,N_14151);
nand U15724 (N_15724,N_14140,N_14730);
or U15725 (N_15725,N_14991,N_14836);
or U15726 (N_15726,N_14860,N_14686);
and U15727 (N_15727,N_14124,N_14819);
nor U15728 (N_15728,N_14223,N_14617);
nand U15729 (N_15729,N_14704,N_14461);
xor U15730 (N_15730,N_14521,N_14191);
nor U15731 (N_15731,N_14696,N_14304);
nor U15732 (N_15732,N_14883,N_14745);
nor U15733 (N_15733,N_14377,N_14536);
and U15734 (N_15734,N_14304,N_14570);
or U15735 (N_15735,N_14714,N_14341);
xor U15736 (N_15736,N_14442,N_14661);
xor U15737 (N_15737,N_14164,N_14994);
xnor U15738 (N_15738,N_14290,N_14082);
or U15739 (N_15739,N_14178,N_14490);
xnor U15740 (N_15740,N_14545,N_14240);
or U15741 (N_15741,N_14817,N_14442);
nand U15742 (N_15742,N_14472,N_14719);
and U15743 (N_15743,N_14366,N_14498);
or U15744 (N_15744,N_14877,N_14416);
nor U15745 (N_15745,N_14275,N_14612);
and U15746 (N_15746,N_14109,N_14629);
or U15747 (N_15747,N_14410,N_14685);
nor U15748 (N_15748,N_14961,N_14476);
or U15749 (N_15749,N_14022,N_14556);
nand U15750 (N_15750,N_14688,N_14168);
xor U15751 (N_15751,N_14839,N_14562);
xnor U15752 (N_15752,N_14269,N_14553);
or U15753 (N_15753,N_14009,N_14673);
nand U15754 (N_15754,N_14624,N_14382);
xor U15755 (N_15755,N_14183,N_14115);
nor U15756 (N_15756,N_14424,N_14380);
xor U15757 (N_15757,N_14020,N_14988);
nor U15758 (N_15758,N_14148,N_14656);
or U15759 (N_15759,N_14224,N_14170);
or U15760 (N_15760,N_14231,N_14979);
nor U15761 (N_15761,N_14823,N_14638);
xnor U15762 (N_15762,N_14805,N_14028);
xor U15763 (N_15763,N_14459,N_14479);
nor U15764 (N_15764,N_14875,N_14457);
xnor U15765 (N_15765,N_14684,N_14412);
and U15766 (N_15766,N_14836,N_14300);
and U15767 (N_15767,N_14412,N_14470);
or U15768 (N_15768,N_14572,N_14757);
nand U15769 (N_15769,N_14909,N_14713);
or U15770 (N_15770,N_14075,N_14618);
and U15771 (N_15771,N_14046,N_14648);
nand U15772 (N_15772,N_14254,N_14366);
xnor U15773 (N_15773,N_14859,N_14781);
or U15774 (N_15774,N_14337,N_14014);
nor U15775 (N_15775,N_14353,N_14374);
xnor U15776 (N_15776,N_14211,N_14349);
or U15777 (N_15777,N_14674,N_14291);
or U15778 (N_15778,N_14012,N_14653);
nand U15779 (N_15779,N_14594,N_14809);
or U15780 (N_15780,N_14352,N_14727);
nor U15781 (N_15781,N_14650,N_14091);
xor U15782 (N_15782,N_14797,N_14813);
xnor U15783 (N_15783,N_14179,N_14319);
and U15784 (N_15784,N_14231,N_14241);
or U15785 (N_15785,N_14697,N_14514);
or U15786 (N_15786,N_14292,N_14523);
or U15787 (N_15787,N_14578,N_14863);
and U15788 (N_15788,N_14364,N_14982);
and U15789 (N_15789,N_14400,N_14928);
nand U15790 (N_15790,N_14446,N_14257);
or U15791 (N_15791,N_14817,N_14958);
xor U15792 (N_15792,N_14415,N_14378);
nand U15793 (N_15793,N_14095,N_14536);
xor U15794 (N_15794,N_14313,N_14205);
nor U15795 (N_15795,N_14415,N_14514);
nand U15796 (N_15796,N_14606,N_14982);
xnor U15797 (N_15797,N_14891,N_14717);
or U15798 (N_15798,N_14989,N_14222);
or U15799 (N_15799,N_14122,N_14255);
and U15800 (N_15800,N_14326,N_14631);
xor U15801 (N_15801,N_14164,N_14390);
nor U15802 (N_15802,N_14668,N_14512);
nand U15803 (N_15803,N_14603,N_14192);
or U15804 (N_15804,N_14522,N_14492);
nand U15805 (N_15805,N_14908,N_14343);
nor U15806 (N_15806,N_14711,N_14589);
and U15807 (N_15807,N_14661,N_14684);
or U15808 (N_15808,N_14349,N_14279);
nand U15809 (N_15809,N_14043,N_14994);
nand U15810 (N_15810,N_14866,N_14471);
nand U15811 (N_15811,N_14742,N_14224);
and U15812 (N_15812,N_14849,N_14588);
xnor U15813 (N_15813,N_14304,N_14272);
nand U15814 (N_15814,N_14974,N_14426);
xnor U15815 (N_15815,N_14389,N_14752);
nand U15816 (N_15816,N_14000,N_14038);
nand U15817 (N_15817,N_14203,N_14835);
nand U15818 (N_15818,N_14086,N_14360);
and U15819 (N_15819,N_14671,N_14274);
nor U15820 (N_15820,N_14358,N_14125);
nand U15821 (N_15821,N_14445,N_14400);
xor U15822 (N_15822,N_14920,N_14107);
xnor U15823 (N_15823,N_14085,N_14488);
or U15824 (N_15824,N_14170,N_14483);
nand U15825 (N_15825,N_14052,N_14982);
nand U15826 (N_15826,N_14720,N_14171);
xor U15827 (N_15827,N_14685,N_14342);
and U15828 (N_15828,N_14284,N_14057);
xnor U15829 (N_15829,N_14476,N_14628);
and U15830 (N_15830,N_14386,N_14976);
xnor U15831 (N_15831,N_14154,N_14371);
nor U15832 (N_15832,N_14558,N_14098);
xor U15833 (N_15833,N_14401,N_14473);
nand U15834 (N_15834,N_14611,N_14885);
and U15835 (N_15835,N_14514,N_14952);
nor U15836 (N_15836,N_14191,N_14451);
nand U15837 (N_15837,N_14982,N_14010);
nor U15838 (N_15838,N_14740,N_14472);
xor U15839 (N_15839,N_14981,N_14100);
or U15840 (N_15840,N_14080,N_14345);
and U15841 (N_15841,N_14866,N_14459);
nor U15842 (N_15842,N_14661,N_14113);
nor U15843 (N_15843,N_14546,N_14153);
nor U15844 (N_15844,N_14899,N_14333);
xnor U15845 (N_15845,N_14176,N_14230);
and U15846 (N_15846,N_14724,N_14638);
nor U15847 (N_15847,N_14658,N_14082);
nor U15848 (N_15848,N_14052,N_14376);
nand U15849 (N_15849,N_14711,N_14293);
nand U15850 (N_15850,N_14301,N_14319);
nand U15851 (N_15851,N_14212,N_14357);
nand U15852 (N_15852,N_14988,N_14330);
xor U15853 (N_15853,N_14229,N_14329);
xor U15854 (N_15854,N_14940,N_14557);
or U15855 (N_15855,N_14065,N_14925);
nand U15856 (N_15856,N_14122,N_14660);
nor U15857 (N_15857,N_14500,N_14986);
and U15858 (N_15858,N_14078,N_14499);
or U15859 (N_15859,N_14082,N_14972);
nor U15860 (N_15860,N_14272,N_14734);
and U15861 (N_15861,N_14164,N_14257);
nor U15862 (N_15862,N_14651,N_14466);
nor U15863 (N_15863,N_14737,N_14425);
nor U15864 (N_15864,N_14512,N_14216);
or U15865 (N_15865,N_14636,N_14035);
xor U15866 (N_15866,N_14790,N_14941);
or U15867 (N_15867,N_14662,N_14152);
and U15868 (N_15868,N_14072,N_14371);
xor U15869 (N_15869,N_14159,N_14237);
or U15870 (N_15870,N_14574,N_14279);
xnor U15871 (N_15871,N_14596,N_14923);
xnor U15872 (N_15872,N_14432,N_14463);
and U15873 (N_15873,N_14043,N_14913);
and U15874 (N_15874,N_14513,N_14128);
nand U15875 (N_15875,N_14959,N_14564);
nor U15876 (N_15876,N_14159,N_14437);
nor U15877 (N_15877,N_14009,N_14261);
nor U15878 (N_15878,N_14227,N_14305);
and U15879 (N_15879,N_14683,N_14902);
nand U15880 (N_15880,N_14501,N_14245);
and U15881 (N_15881,N_14043,N_14479);
nor U15882 (N_15882,N_14021,N_14293);
xor U15883 (N_15883,N_14909,N_14724);
xor U15884 (N_15884,N_14056,N_14215);
xnor U15885 (N_15885,N_14117,N_14414);
nand U15886 (N_15886,N_14553,N_14710);
or U15887 (N_15887,N_14160,N_14064);
nand U15888 (N_15888,N_14180,N_14211);
or U15889 (N_15889,N_14846,N_14602);
nor U15890 (N_15890,N_14737,N_14866);
xnor U15891 (N_15891,N_14786,N_14453);
nor U15892 (N_15892,N_14134,N_14041);
nor U15893 (N_15893,N_14339,N_14593);
nand U15894 (N_15894,N_14019,N_14085);
nand U15895 (N_15895,N_14617,N_14587);
nand U15896 (N_15896,N_14446,N_14243);
xor U15897 (N_15897,N_14130,N_14611);
nand U15898 (N_15898,N_14944,N_14456);
nand U15899 (N_15899,N_14430,N_14295);
or U15900 (N_15900,N_14177,N_14710);
nand U15901 (N_15901,N_14732,N_14460);
xnor U15902 (N_15902,N_14899,N_14171);
xor U15903 (N_15903,N_14104,N_14914);
and U15904 (N_15904,N_14430,N_14225);
nand U15905 (N_15905,N_14828,N_14002);
nand U15906 (N_15906,N_14712,N_14235);
or U15907 (N_15907,N_14502,N_14065);
nand U15908 (N_15908,N_14569,N_14984);
nor U15909 (N_15909,N_14680,N_14828);
or U15910 (N_15910,N_14399,N_14383);
or U15911 (N_15911,N_14636,N_14880);
or U15912 (N_15912,N_14360,N_14097);
xor U15913 (N_15913,N_14753,N_14484);
nand U15914 (N_15914,N_14614,N_14711);
nand U15915 (N_15915,N_14417,N_14670);
nand U15916 (N_15916,N_14820,N_14234);
xor U15917 (N_15917,N_14609,N_14634);
nand U15918 (N_15918,N_14958,N_14265);
and U15919 (N_15919,N_14517,N_14862);
or U15920 (N_15920,N_14766,N_14339);
nand U15921 (N_15921,N_14854,N_14060);
xor U15922 (N_15922,N_14393,N_14352);
or U15923 (N_15923,N_14120,N_14283);
or U15924 (N_15924,N_14836,N_14664);
nor U15925 (N_15925,N_14576,N_14430);
or U15926 (N_15926,N_14937,N_14730);
nand U15927 (N_15927,N_14516,N_14137);
nor U15928 (N_15928,N_14816,N_14647);
and U15929 (N_15929,N_14384,N_14178);
and U15930 (N_15930,N_14009,N_14169);
xor U15931 (N_15931,N_14084,N_14614);
xor U15932 (N_15932,N_14662,N_14125);
nand U15933 (N_15933,N_14828,N_14444);
or U15934 (N_15934,N_14197,N_14166);
xnor U15935 (N_15935,N_14784,N_14812);
xnor U15936 (N_15936,N_14861,N_14749);
nor U15937 (N_15937,N_14727,N_14709);
and U15938 (N_15938,N_14623,N_14237);
or U15939 (N_15939,N_14590,N_14701);
and U15940 (N_15940,N_14500,N_14357);
or U15941 (N_15941,N_14530,N_14463);
nand U15942 (N_15942,N_14856,N_14022);
or U15943 (N_15943,N_14068,N_14326);
nand U15944 (N_15944,N_14899,N_14087);
nor U15945 (N_15945,N_14367,N_14353);
and U15946 (N_15946,N_14598,N_14345);
nor U15947 (N_15947,N_14325,N_14698);
or U15948 (N_15948,N_14421,N_14405);
or U15949 (N_15949,N_14109,N_14303);
nand U15950 (N_15950,N_14291,N_14435);
xor U15951 (N_15951,N_14784,N_14471);
nand U15952 (N_15952,N_14810,N_14980);
or U15953 (N_15953,N_14705,N_14620);
and U15954 (N_15954,N_14771,N_14181);
xor U15955 (N_15955,N_14500,N_14924);
nand U15956 (N_15956,N_14272,N_14371);
or U15957 (N_15957,N_14482,N_14095);
xor U15958 (N_15958,N_14299,N_14220);
nand U15959 (N_15959,N_14992,N_14037);
xnor U15960 (N_15960,N_14161,N_14392);
and U15961 (N_15961,N_14895,N_14827);
nor U15962 (N_15962,N_14795,N_14852);
xor U15963 (N_15963,N_14039,N_14454);
or U15964 (N_15964,N_14596,N_14920);
xnor U15965 (N_15965,N_14503,N_14147);
and U15966 (N_15966,N_14604,N_14984);
nor U15967 (N_15967,N_14662,N_14335);
nor U15968 (N_15968,N_14329,N_14869);
and U15969 (N_15969,N_14864,N_14685);
and U15970 (N_15970,N_14757,N_14662);
nor U15971 (N_15971,N_14072,N_14900);
xor U15972 (N_15972,N_14240,N_14942);
and U15973 (N_15973,N_14457,N_14686);
xor U15974 (N_15974,N_14627,N_14461);
xnor U15975 (N_15975,N_14596,N_14693);
xnor U15976 (N_15976,N_14792,N_14445);
or U15977 (N_15977,N_14017,N_14660);
xor U15978 (N_15978,N_14986,N_14338);
xnor U15979 (N_15979,N_14710,N_14196);
and U15980 (N_15980,N_14472,N_14386);
nor U15981 (N_15981,N_14139,N_14689);
or U15982 (N_15982,N_14511,N_14894);
nand U15983 (N_15983,N_14742,N_14390);
and U15984 (N_15984,N_14563,N_14987);
xor U15985 (N_15985,N_14533,N_14526);
nand U15986 (N_15986,N_14283,N_14105);
xnor U15987 (N_15987,N_14849,N_14162);
xor U15988 (N_15988,N_14895,N_14870);
nor U15989 (N_15989,N_14932,N_14766);
nor U15990 (N_15990,N_14143,N_14073);
nand U15991 (N_15991,N_14316,N_14203);
xor U15992 (N_15992,N_14732,N_14657);
nand U15993 (N_15993,N_14392,N_14786);
nand U15994 (N_15994,N_14766,N_14837);
nand U15995 (N_15995,N_14902,N_14850);
and U15996 (N_15996,N_14868,N_14130);
xnor U15997 (N_15997,N_14822,N_14594);
and U15998 (N_15998,N_14409,N_14093);
xnor U15999 (N_15999,N_14518,N_14278);
nor U16000 (N_16000,N_15334,N_15543);
or U16001 (N_16001,N_15705,N_15665);
nor U16002 (N_16002,N_15793,N_15650);
xor U16003 (N_16003,N_15963,N_15842);
nand U16004 (N_16004,N_15968,N_15727);
nor U16005 (N_16005,N_15876,N_15918);
or U16006 (N_16006,N_15508,N_15360);
xor U16007 (N_16007,N_15518,N_15662);
xnor U16008 (N_16008,N_15633,N_15310);
nand U16009 (N_16009,N_15696,N_15279);
nor U16010 (N_16010,N_15988,N_15252);
xnor U16011 (N_16011,N_15701,N_15156);
and U16012 (N_16012,N_15517,N_15493);
nor U16013 (N_16013,N_15086,N_15632);
xor U16014 (N_16014,N_15767,N_15284);
or U16015 (N_16015,N_15901,N_15207);
and U16016 (N_16016,N_15238,N_15681);
nor U16017 (N_16017,N_15406,N_15470);
or U16018 (N_16018,N_15249,N_15531);
xnor U16019 (N_16019,N_15673,N_15983);
nand U16020 (N_16020,N_15747,N_15574);
or U16021 (N_16021,N_15029,N_15514);
or U16022 (N_16022,N_15686,N_15698);
and U16023 (N_16023,N_15787,N_15516);
nand U16024 (N_16024,N_15886,N_15208);
and U16025 (N_16025,N_15078,N_15391);
nor U16026 (N_16026,N_15437,N_15889);
and U16027 (N_16027,N_15578,N_15049);
xnor U16028 (N_16028,N_15659,N_15134);
nand U16029 (N_16029,N_15151,N_15611);
nor U16030 (N_16030,N_15964,N_15711);
nor U16031 (N_16031,N_15240,N_15872);
nor U16032 (N_16032,N_15112,N_15800);
nor U16033 (N_16033,N_15625,N_15837);
and U16034 (N_16034,N_15716,N_15266);
and U16035 (N_16035,N_15098,N_15942);
nand U16036 (N_16036,N_15458,N_15172);
and U16037 (N_16037,N_15162,N_15168);
nand U16038 (N_16038,N_15413,N_15763);
and U16039 (N_16039,N_15989,N_15569);
xnor U16040 (N_16040,N_15728,N_15147);
xnor U16041 (N_16041,N_15575,N_15772);
or U16042 (N_16042,N_15548,N_15538);
xnor U16043 (N_16043,N_15265,N_15580);
or U16044 (N_16044,N_15074,N_15934);
nand U16045 (N_16045,N_15161,N_15140);
nor U16046 (N_16046,N_15606,N_15392);
xor U16047 (N_16047,N_15794,N_15670);
and U16048 (N_16048,N_15402,N_15327);
xnor U16049 (N_16049,N_15163,N_15072);
or U16050 (N_16050,N_15788,N_15521);
and U16051 (N_16051,N_15329,N_15979);
or U16052 (N_16052,N_15210,N_15453);
or U16053 (N_16053,N_15860,N_15125);
or U16054 (N_16054,N_15830,N_15454);
and U16055 (N_16055,N_15082,N_15067);
xor U16056 (N_16056,N_15897,N_15755);
or U16057 (N_16057,N_15032,N_15275);
nor U16058 (N_16058,N_15190,N_15272);
nand U16059 (N_16059,N_15894,N_15441);
nand U16060 (N_16060,N_15189,N_15631);
nor U16061 (N_16061,N_15022,N_15034);
xnor U16062 (N_16062,N_15654,N_15945);
nor U16063 (N_16063,N_15177,N_15375);
nand U16064 (N_16064,N_15510,N_15605);
or U16065 (N_16065,N_15976,N_15912);
nand U16066 (N_16066,N_15774,N_15960);
or U16067 (N_16067,N_15776,N_15498);
and U16068 (N_16068,N_15791,N_15121);
xor U16069 (N_16069,N_15176,N_15496);
xor U16070 (N_16070,N_15330,N_15201);
nand U16071 (N_16071,N_15640,N_15424);
and U16072 (N_16072,N_15314,N_15014);
or U16073 (N_16073,N_15018,N_15223);
and U16074 (N_16074,N_15095,N_15479);
and U16075 (N_16075,N_15855,N_15104);
or U16076 (N_16076,N_15846,N_15011);
nor U16077 (N_16077,N_15278,N_15205);
nand U16078 (N_16078,N_15925,N_15347);
nor U16079 (N_16079,N_15867,N_15806);
and U16080 (N_16080,N_15101,N_15396);
nand U16081 (N_16081,N_15380,N_15059);
or U16082 (N_16082,N_15142,N_15592);
nand U16083 (N_16083,N_15649,N_15468);
and U16084 (N_16084,N_15965,N_15568);
or U16085 (N_16085,N_15534,N_15039);
xnor U16086 (N_16086,N_15981,N_15612);
nor U16087 (N_16087,N_15823,N_15440);
nor U16088 (N_16088,N_15319,N_15218);
or U16089 (N_16089,N_15445,N_15955);
nand U16090 (N_16090,N_15923,N_15141);
or U16091 (N_16091,N_15819,N_15048);
xnor U16092 (N_16092,N_15024,N_15922);
and U16093 (N_16093,N_15017,N_15751);
or U16094 (N_16094,N_15801,N_15961);
nand U16095 (N_16095,N_15571,N_15224);
xnor U16096 (N_16096,N_15890,N_15164);
or U16097 (N_16097,N_15697,N_15308);
nand U16098 (N_16098,N_15583,N_15461);
nor U16099 (N_16099,N_15335,N_15732);
nand U16100 (N_16100,N_15115,N_15044);
and U16101 (N_16101,N_15301,N_15497);
nand U16102 (N_16102,N_15621,N_15685);
xor U16103 (N_16103,N_15462,N_15924);
xnor U16104 (N_16104,N_15825,N_15427);
xnor U16105 (N_16105,N_15630,N_15160);
xor U16106 (N_16106,N_15930,N_15434);
xor U16107 (N_16107,N_15904,N_15020);
nor U16108 (N_16108,N_15386,N_15645);
and U16109 (N_16109,N_15602,N_15744);
nand U16110 (N_16110,N_15834,N_15753);
nand U16111 (N_16111,N_15439,N_15704);
or U16112 (N_16112,N_15920,N_15417);
nand U16113 (N_16113,N_15500,N_15844);
nand U16114 (N_16114,N_15501,N_15393);
or U16115 (N_16115,N_15353,N_15264);
and U16116 (N_16116,N_15731,N_15700);
nand U16117 (N_16117,N_15259,N_15225);
nand U16118 (N_16118,N_15345,N_15430);
or U16119 (N_16119,N_15146,N_15053);
nand U16120 (N_16120,N_15560,N_15490);
and U16121 (N_16121,N_15581,N_15332);
or U16122 (N_16122,N_15084,N_15343);
and U16123 (N_16123,N_15505,N_15882);
or U16124 (N_16124,N_15478,N_15137);
or U16125 (N_16125,N_15364,N_15178);
xnor U16126 (N_16126,N_15619,N_15358);
nand U16127 (N_16127,N_15292,N_15277);
and U16128 (N_16128,N_15390,N_15276);
or U16129 (N_16129,N_15643,N_15641);
xnor U16130 (N_16130,N_15322,N_15451);
xnor U16131 (N_16131,N_15863,N_15384);
xor U16132 (N_16132,N_15241,N_15809);
nand U16133 (N_16133,N_15985,N_15947);
xor U16134 (N_16134,N_15399,N_15449);
nand U16135 (N_16135,N_15423,N_15750);
xnor U16136 (N_16136,N_15484,N_15573);
xor U16137 (N_16137,N_15622,N_15227);
xor U16138 (N_16138,N_15653,N_15799);
nand U16139 (N_16139,N_15236,N_15365);
or U16140 (N_16140,N_15344,N_15715);
nand U16141 (N_16141,N_15624,N_15895);
nand U16142 (N_16142,N_15303,N_15033);
and U16143 (N_16143,N_15457,N_15455);
or U16144 (N_16144,N_15688,N_15987);
nor U16145 (N_16145,N_15250,N_15133);
or U16146 (N_16146,N_15743,N_15467);
nand U16147 (N_16147,N_15061,N_15850);
or U16148 (N_16148,N_15937,N_15851);
and U16149 (N_16149,N_15542,N_15356);
nor U16150 (N_16150,N_15898,N_15587);
nand U16151 (N_16151,N_15056,N_15940);
nor U16152 (N_16152,N_15166,N_15181);
nor U16153 (N_16153,N_15369,N_15756);
nor U16154 (N_16154,N_15749,N_15055);
xnor U16155 (N_16155,N_15174,N_15674);
and U16156 (N_16156,N_15415,N_15013);
nor U16157 (N_16157,N_15476,N_15070);
nor U16158 (N_16158,N_15745,N_15324);
xor U16159 (N_16159,N_15376,N_15927);
nand U16160 (N_16160,N_15746,N_15248);
nor U16161 (N_16161,N_15970,N_15768);
xor U16162 (N_16162,N_15191,N_15807);
and U16163 (N_16163,N_15131,N_15342);
nor U16164 (N_16164,N_15975,N_15007);
nand U16165 (N_16165,N_15286,N_15599);
or U16166 (N_16166,N_15796,N_15389);
xor U16167 (N_16167,N_15471,N_15220);
nand U16168 (N_16168,N_15952,N_15526);
or U16169 (N_16169,N_15996,N_15068);
and U16170 (N_16170,N_15054,N_15312);
xnor U16171 (N_16171,N_15792,N_15184);
nand U16172 (N_16172,N_15817,N_15758);
nor U16173 (N_16173,N_15341,N_15910);
nand U16174 (N_16174,N_15089,N_15903);
nor U16175 (N_16175,N_15117,N_15735);
nand U16176 (N_16176,N_15403,N_15042);
xnor U16177 (N_16177,N_15243,N_15331);
nand U16178 (N_16178,N_15422,N_15601);
xnor U16179 (N_16179,N_15757,N_15107);
and U16180 (N_16180,N_15929,N_15660);
xor U16181 (N_16181,N_15198,N_15720);
nand U16182 (N_16182,N_15246,N_15684);
nor U16183 (N_16183,N_15325,N_15972);
nor U16184 (N_16184,N_15244,N_15433);
nand U16185 (N_16185,N_15815,N_15617);
nor U16186 (N_16186,N_15520,N_15169);
or U16187 (N_16187,N_15992,N_15754);
nor U16188 (N_16188,N_15443,N_15426);
nand U16189 (N_16189,N_15442,N_15299);
xnor U16190 (N_16190,N_15999,N_15762);
or U16191 (N_16191,N_15216,N_15719);
or U16192 (N_16192,N_15118,N_15721);
nor U16193 (N_16193,N_15969,N_15447);
nand U16194 (N_16194,N_15946,N_15629);
and U16195 (N_16195,N_15382,N_15843);
or U16196 (N_16196,N_15919,N_15820);
and U16197 (N_16197,N_15884,N_15984);
nor U16198 (N_16198,N_15866,N_15603);
nand U16199 (N_16199,N_15337,N_15388);
or U16200 (N_16200,N_15450,N_15371);
nand U16201 (N_16201,N_15222,N_15595);
nand U16202 (N_16202,N_15600,N_15586);
or U16203 (N_16203,N_15003,N_15075);
and U16204 (N_16204,N_15309,N_15857);
nand U16205 (N_16205,N_15714,N_15444);
xor U16206 (N_16206,N_15194,N_15057);
and U16207 (N_16207,N_15723,N_15880);
xnor U16208 (N_16208,N_15565,N_15536);
nor U16209 (N_16209,N_15040,N_15047);
xnor U16210 (N_16210,N_15703,N_15609);
and U16211 (N_16211,N_15827,N_15463);
or U16212 (N_16212,N_15563,N_15879);
nor U16213 (N_16213,N_15483,N_15247);
nor U16214 (N_16214,N_15544,N_15495);
nor U16215 (N_16215,N_15030,N_15859);
nand U16216 (N_16216,N_15352,N_15110);
or U16217 (N_16217,N_15338,N_15294);
nand U16218 (N_16218,N_15663,N_15209);
nor U16219 (N_16219,N_15366,N_15432);
nor U16220 (N_16220,N_15780,N_15111);
or U16221 (N_16221,N_15256,N_15974);
xor U16222 (N_16222,N_15533,N_15349);
or U16223 (N_16223,N_15537,N_15302);
or U16224 (N_16224,N_15893,N_15734);
or U16225 (N_16225,N_15865,N_15932);
and U16226 (N_16226,N_15885,N_15122);
nand U16227 (N_16227,N_15847,N_15124);
xnor U16228 (N_16228,N_15785,N_15775);
and U16229 (N_16229,N_15570,N_15050);
nand U16230 (N_16230,N_15858,N_15395);
and U16231 (N_16231,N_15318,N_15379);
or U16232 (N_16232,N_15182,N_15092);
or U16233 (N_16233,N_15438,N_15914);
nand U16234 (N_16234,N_15881,N_15411);
nor U16235 (N_16235,N_15550,N_15203);
xnor U16236 (N_16236,N_15096,N_15547);
nand U16237 (N_16237,N_15149,N_15835);
and U16238 (N_16238,N_15956,N_15966);
nor U16239 (N_16239,N_15480,N_15041);
or U16240 (N_16240,N_15724,N_15200);
and U16241 (N_16241,N_15921,N_15598);
nor U16242 (N_16242,N_15502,N_15973);
or U16243 (N_16243,N_15350,N_15492);
nand U16244 (N_16244,N_15414,N_15691);
or U16245 (N_16245,N_15957,N_15810);
and U16246 (N_16246,N_15839,N_15404);
nand U16247 (N_16247,N_15005,N_15226);
xor U16248 (N_16248,N_15473,N_15270);
or U16249 (N_16249,N_15094,N_15316);
nor U16250 (N_16250,N_15525,N_15362);
and U16251 (N_16251,N_15287,N_15738);
nor U16252 (N_16252,N_15069,N_15091);
nor U16253 (N_16253,N_15572,N_15513);
nor U16254 (N_16254,N_15900,N_15398);
or U16255 (N_16255,N_15180,N_15120);
and U16256 (N_16256,N_15229,N_15425);
and U16257 (N_16257,N_15764,N_15677);
nand U16258 (N_16258,N_15130,N_15113);
xnor U16259 (N_16259,N_15908,N_15737);
or U16260 (N_16260,N_15618,N_15295);
and U16261 (N_16261,N_15108,N_15448);
nand U16262 (N_16262,N_15642,N_15849);
nor U16263 (N_16263,N_15675,N_15887);
nand U16264 (N_16264,N_15173,N_15135);
nand U16265 (N_16265,N_15838,N_15896);
or U16266 (N_16266,N_15410,N_15816);
nand U16267 (N_16267,N_15077,N_15431);
nand U16268 (N_16268,N_15577,N_15071);
nor U16269 (N_16269,N_15596,N_15854);
nor U16270 (N_16270,N_15931,N_15915);
nand U16271 (N_16271,N_15759,N_15004);
nand U16272 (N_16272,N_15967,N_15260);
and U16273 (N_16273,N_15261,N_15676);
and U16274 (N_16274,N_15304,N_15652);
and U16275 (N_16275,N_15841,N_15954);
nor U16276 (N_16276,N_15891,N_15143);
xor U16277 (N_16277,N_15001,N_15980);
or U16278 (N_16278,N_15928,N_15373);
or U16279 (N_16279,N_15367,N_15636);
and U16280 (N_16280,N_15401,N_15482);
nor U16281 (N_16281,N_15281,N_15035);
and U16282 (N_16282,N_15293,N_15986);
nor U16283 (N_16283,N_15128,N_15043);
or U16284 (N_16284,N_15037,N_15469);
nand U16285 (N_16285,N_15845,N_15795);
xor U16286 (N_16286,N_15661,N_15824);
xor U16287 (N_16287,N_15193,N_15667);
and U16288 (N_16288,N_15736,N_15009);
or U16289 (N_16289,N_15188,N_15808);
xor U16290 (N_16290,N_15826,N_15320);
xor U16291 (N_16291,N_15564,N_15805);
or U16292 (N_16292,N_15405,N_15085);
or U16293 (N_16293,N_15199,N_15995);
xnor U16294 (N_16294,N_15524,N_15585);
xor U16295 (N_16295,N_15726,N_15027);
or U16296 (N_16296,N_15228,N_15594);
xor U16297 (N_16297,N_15202,N_15997);
nor U16298 (N_16298,N_15786,N_15706);
nand U16299 (N_16299,N_15710,N_15941);
xor U16300 (N_16300,N_15875,N_15582);
or U16301 (N_16301,N_15852,N_15475);
nand U16302 (N_16302,N_15740,N_15693);
and U16303 (N_16303,N_15217,N_15519);
nor U16304 (N_16304,N_15267,N_15456);
or U16305 (N_16305,N_15452,N_15771);
and U16306 (N_16306,N_15627,N_15487);
or U16307 (N_16307,N_15378,N_15080);
and U16308 (N_16308,N_15552,N_15822);
or U16309 (N_16309,N_15213,N_15678);
xor U16310 (N_16310,N_15953,N_15197);
nand U16311 (N_16311,N_15647,N_15639);
xor U16312 (N_16312,N_15076,N_15298);
and U16313 (N_16313,N_15832,N_15836);
nor U16314 (N_16314,N_15368,N_15351);
nor U16315 (N_16315,N_15421,N_15129);
or U16316 (N_16316,N_15576,N_15765);
and U16317 (N_16317,N_15917,N_15268);
nand U16318 (N_16318,N_15274,N_15789);
nor U16319 (N_16319,N_15944,N_15991);
nand U16320 (N_16320,N_15233,N_15263);
or U16321 (N_16321,N_15614,N_15902);
or U16322 (N_16322,N_15237,N_15503);
nor U16323 (N_16323,N_15257,N_15766);
nor U16324 (N_16324,N_15026,N_15702);
nor U16325 (N_16325,N_15515,N_15167);
nor U16326 (N_16326,N_15400,N_15540);
xor U16327 (N_16327,N_15725,N_15230);
and U16328 (N_16328,N_15769,N_15959);
or U16329 (N_16329,N_15152,N_15109);
or U16330 (N_16330,N_15713,N_15804);
xor U16331 (N_16331,N_15588,N_15803);
and U16332 (N_16332,N_15459,N_15848);
and U16333 (N_16333,N_15387,N_15802);
nor U16334 (N_16334,N_15127,N_15313);
xnor U16335 (N_16335,N_15783,N_15797);
nor U16336 (N_16336,N_15814,N_15148);
nor U16337 (N_16337,N_15994,N_15340);
xnor U16338 (N_16338,N_15555,N_15474);
nand U16339 (N_16339,N_15253,N_15878);
nor U16340 (N_16340,N_15255,N_15584);
nor U16341 (N_16341,N_15099,N_15262);
nor U16342 (N_16342,N_15407,N_15290);
and U16343 (N_16343,N_15635,N_15006);
and U16344 (N_16344,N_15179,N_15221);
and U16345 (N_16345,N_15656,N_15978);
nand U16346 (N_16346,N_15012,N_15778);
or U16347 (N_16347,N_15010,N_15593);
and U16348 (N_16348,N_15073,N_15155);
nor U16349 (N_16349,N_15561,N_15363);
and U16350 (N_16350,N_15307,N_15718);
and U16351 (N_16351,N_15465,N_15509);
or U16352 (N_16352,N_15938,N_15782);
nand U16353 (N_16353,N_15139,N_15219);
nor U16354 (N_16354,N_15297,N_15911);
nor U16355 (N_16355,N_15485,N_15062);
or U16356 (N_16356,N_15874,N_15045);
or U16357 (N_16357,N_15046,N_15739);
and U16358 (N_16358,N_15326,N_15689);
nand U16359 (N_16359,N_15385,N_15507);
and U16360 (N_16360,N_15321,N_15206);
nor U16361 (N_16361,N_15549,N_15254);
and U16362 (N_16362,N_15418,N_15813);
or U16363 (N_16363,N_15950,N_15899);
and U16364 (N_16364,N_15864,N_15812);
nand U16365 (N_16365,N_15192,N_15119);
and U16366 (N_16366,N_15913,N_15694);
nand U16367 (N_16367,N_15008,N_15021);
or U16368 (N_16368,N_15840,N_15195);
nand U16369 (N_16369,N_15370,N_15690);
nand U16370 (N_16370,N_15869,N_15993);
nand U16371 (N_16371,N_15185,N_15712);
nand U16372 (N_16372,N_15760,N_15905);
nand U16373 (N_16373,N_15512,N_15409);
xor U16374 (N_16374,N_15936,N_15752);
xor U16375 (N_16375,N_15877,N_15958);
or U16376 (N_16376,N_15394,N_15486);
or U16377 (N_16377,N_15528,N_15861);
nor U16378 (N_16378,N_15657,N_15285);
and U16379 (N_16379,N_15023,N_15669);
xnor U16380 (N_16380,N_15291,N_15031);
nor U16381 (N_16381,N_15907,N_15477);
xnor U16382 (N_16382,N_15655,N_15242);
and U16383 (N_16383,N_15136,N_15158);
and U16384 (N_16384,N_15666,N_15436);
xor U16385 (N_16385,N_15183,N_15412);
nand U16386 (N_16386,N_15589,N_15644);
or U16387 (N_16387,N_15093,N_15729);
and U16388 (N_16388,N_15977,N_15790);
nor U16389 (N_16389,N_15990,N_15620);
or U16390 (N_16390,N_15773,N_15638);
xnor U16391 (N_16391,N_15311,N_15679);
or U16392 (N_16392,N_15066,N_15888);
nor U16393 (N_16393,N_15523,N_15058);
or U16394 (N_16394,N_15153,N_15489);
nor U16395 (N_16395,N_15672,N_15871);
xor U16396 (N_16396,N_15002,N_15028);
nor U16397 (N_16397,N_15658,N_15355);
xor U16398 (N_16398,N_15777,N_15943);
nand U16399 (N_16399,N_15289,N_15591);
nor U16400 (N_16400,N_15154,N_15204);
or U16401 (N_16401,N_15408,N_15687);
xor U16402 (N_16402,N_15504,N_15811);
and U16403 (N_16403,N_15336,N_15545);
or U16404 (N_16404,N_15527,N_15597);
xnor U16405 (N_16405,N_15613,N_15138);
or U16406 (N_16406,N_15615,N_15211);
nor U16407 (N_16407,N_15870,N_15419);
and U16408 (N_16408,N_15779,N_15323);
and U16409 (N_16409,N_15081,N_15283);
or U16410 (N_16410,N_15126,N_15377);
nand U16411 (N_16411,N_15511,N_15951);
xor U16412 (N_16412,N_15541,N_15892);
and U16413 (N_16413,N_15818,N_15562);
nand U16414 (N_16414,N_15273,N_15962);
xnor U16415 (N_16415,N_15546,N_15051);
and U16416 (N_16416,N_15251,N_15935);
xor U16417 (N_16417,N_15717,N_15038);
and U16418 (N_16418,N_15535,N_15446);
nand U16419 (N_16419,N_15231,N_15579);
or U16420 (N_16420,N_15116,N_15671);
or U16421 (N_16421,N_15558,N_15175);
or U16422 (N_16422,N_15494,N_15102);
xnor U16423 (N_16423,N_15829,N_15648);
and U16424 (N_16424,N_15730,N_15556);
nor U16425 (N_16425,N_15114,N_15328);
nand U16426 (N_16426,N_15464,N_15604);
nand U16427 (N_16427,N_15566,N_15868);
nand U16428 (N_16428,N_15397,N_15488);
nor U16429 (N_16429,N_15144,N_15239);
and U16430 (N_16430,N_15105,N_15145);
or U16431 (N_16431,N_15460,N_15235);
nand U16432 (N_16432,N_15269,N_15709);
or U16433 (N_16433,N_15567,N_15909);
nor U16434 (N_16434,N_15616,N_15186);
nor U16435 (N_16435,N_15361,N_15828);
or U16436 (N_16436,N_15982,N_15491);
nand U16437 (N_16437,N_15060,N_15171);
nand U16438 (N_16438,N_15036,N_15998);
nand U16439 (N_16439,N_15083,N_15761);
and U16440 (N_16440,N_15472,N_15357);
xor U16441 (N_16441,N_15833,N_15087);
nand U16442 (N_16442,N_15097,N_15348);
or U16443 (N_16443,N_15466,N_15300);
or U16444 (N_16444,N_15831,N_15280);
nor U16445 (N_16445,N_15634,N_15853);
xnor U16446 (N_16446,N_15100,N_15150);
nor U16447 (N_16447,N_15532,N_15607);
nor U16448 (N_16448,N_15063,N_15079);
and U16449 (N_16449,N_15165,N_15015);
and U16450 (N_16450,N_15381,N_15234);
nor U16451 (N_16451,N_15682,N_15668);
or U16452 (N_16452,N_15019,N_15608);
and U16453 (N_16453,N_15196,N_15354);
xor U16454 (N_16454,N_15559,N_15692);
and U16455 (N_16455,N_15305,N_15064);
nor U16456 (N_16456,N_15680,N_15282);
xnor U16457 (N_16457,N_15626,N_15245);
nand U16458 (N_16458,N_15435,N_15339);
nand U16459 (N_16459,N_15383,N_15722);
and U16460 (N_16460,N_15333,N_15428);
nor U16461 (N_16461,N_15103,N_15939);
nor U16462 (N_16462,N_15215,N_15906);
and U16463 (N_16463,N_15016,N_15288);
and U16464 (N_16464,N_15933,N_15557);
nor U16465 (N_16465,N_15212,N_15232);
xor U16466 (N_16466,N_15551,N_15429);
or U16467 (N_16467,N_15916,N_15025);
and U16468 (N_16468,N_15157,N_15741);
nand U16469 (N_16469,N_15315,N_15522);
nand U16470 (N_16470,N_15862,N_15346);
or U16471 (N_16471,N_15530,N_15499);
and U16472 (N_16472,N_15372,N_15506);
xor U16473 (N_16473,N_15374,N_15317);
nand U16474 (N_16474,N_15416,N_15707);
xnor U16475 (N_16475,N_15481,N_15610);
nor U16476 (N_16476,N_15000,N_15539);
nor U16477 (N_16477,N_15748,N_15733);
and U16478 (N_16478,N_15065,N_15637);
or U16479 (N_16479,N_15359,N_15420);
nand U16480 (N_16480,N_15554,N_15664);
xnor U16481 (N_16481,N_15646,N_15090);
xnor U16482 (N_16482,N_15770,N_15781);
nor U16483 (N_16483,N_15873,N_15856);
xor U16484 (N_16484,N_15784,N_15699);
nor U16485 (N_16485,N_15553,N_15214);
and U16486 (N_16486,N_15926,N_15258);
xnor U16487 (N_16487,N_15052,N_15683);
nand U16488 (N_16488,N_15529,N_15623);
and U16489 (N_16489,N_15628,N_15106);
nor U16490 (N_16490,N_15590,N_15159);
and U16491 (N_16491,N_15949,N_15695);
nand U16492 (N_16492,N_15742,N_15798);
and U16493 (N_16493,N_15306,N_15088);
and U16494 (N_16494,N_15170,N_15271);
nor U16495 (N_16495,N_15132,N_15821);
xor U16496 (N_16496,N_15296,N_15948);
or U16497 (N_16497,N_15883,N_15971);
and U16498 (N_16498,N_15651,N_15708);
nand U16499 (N_16499,N_15187,N_15123);
or U16500 (N_16500,N_15531,N_15460);
or U16501 (N_16501,N_15346,N_15252);
and U16502 (N_16502,N_15514,N_15150);
or U16503 (N_16503,N_15526,N_15034);
xnor U16504 (N_16504,N_15722,N_15737);
and U16505 (N_16505,N_15795,N_15291);
nand U16506 (N_16506,N_15366,N_15641);
nand U16507 (N_16507,N_15367,N_15961);
nand U16508 (N_16508,N_15057,N_15162);
nor U16509 (N_16509,N_15963,N_15322);
and U16510 (N_16510,N_15304,N_15488);
and U16511 (N_16511,N_15941,N_15417);
nand U16512 (N_16512,N_15332,N_15699);
or U16513 (N_16513,N_15845,N_15791);
xnor U16514 (N_16514,N_15560,N_15594);
or U16515 (N_16515,N_15157,N_15478);
nor U16516 (N_16516,N_15787,N_15144);
or U16517 (N_16517,N_15346,N_15478);
nor U16518 (N_16518,N_15924,N_15014);
xnor U16519 (N_16519,N_15677,N_15096);
nor U16520 (N_16520,N_15095,N_15434);
or U16521 (N_16521,N_15536,N_15835);
nand U16522 (N_16522,N_15901,N_15985);
nor U16523 (N_16523,N_15865,N_15916);
nor U16524 (N_16524,N_15031,N_15217);
nand U16525 (N_16525,N_15878,N_15540);
and U16526 (N_16526,N_15864,N_15024);
nor U16527 (N_16527,N_15414,N_15160);
and U16528 (N_16528,N_15336,N_15868);
nor U16529 (N_16529,N_15518,N_15529);
nor U16530 (N_16530,N_15615,N_15986);
and U16531 (N_16531,N_15411,N_15746);
nor U16532 (N_16532,N_15650,N_15080);
nand U16533 (N_16533,N_15450,N_15221);
nand U16534 (N_16534,N_15053,N_15025);
nor U16535 (N_16535,N_15611,N_15652);
nand U16536 (N_16536,N_15909,N_15246);
nor U16537 (N_16537,N_15681,N_15746);
xor U16538 (N_16538,N_15963,N_15311);
and U16539 (N_16539,N_15981,N_15290);
or U16540 (N_16540,N_15510,N_15654);
nor U16541 (N_16541,N_15736,N_15876);
nor U16542 (N_16542,N_15378,N_15946);
nand U16543 (N_16543,N_15878,N_15663);
nand U16544 (N_16544,N_15965,N_15654);
nor U16545 (N_16545,N_15441,N_15722);
xor U16546 (N_16546,N_15316,N_15271);
nand U16547 (N_16547,N_15346,N_15871);
and U16548 (N_16548,N_15464,N_15350);
or U16549 (N_16549,N_15667,N_15893);
or U16550 (N_16550,N_15995,N_15197);
and U16551 (N_16551,N_15325,N_15722);
xor U16552 (N_16552,N_15437,N_15565);
nor U16553 (N_16553,N_15738,N_15913);
and U16554 (N_16554,N_15375,N_15590);
nand U16555 (N_16555,N_15289,N_15554);
xor U16556 (N_16556,N_15013,N_15914);
or U16557 (N_16557,N_15856,N_15041);
or U16558 (N_16558,N_15904,N_15352);
nor U16559 (N_16559,N_15235,N_15224);
nor U16560 (N_16560,N_15836,N_15711);
and U16561 (N_16561,N_15472,N_15984);
nand U16562 (N_16562,N_15386,N_15942);
nor U16563 (N_16563,N_15803,N_15189);
xnor U16564 (N_16564,N_15767,N_15277);
and U16565 (N_16565,N_15494,N_15359);
and U16566 (N_16566,N_15486,N_15048);
or U16567 (N_16567,N_15084,N_15234);
or U16568 (N_16568,N_15904,N_15975);
xnor U16569 (N_16569,N_15648,N_15519);
xnor U16570 (N_16570,N_15087,N_15521);
or U16571 (N_16571,N_15845,N_15125);
or U16572 (N_16572,N_15784,N_15568);
nor U16573 (N_16573,N_15601,N_15413);
nand U16574 (N_16574,N_15088,N_15762);
nand U16575 (N_16575,N_15132,N_15965);
and U16576 (N_16576,N_15509,N_15440);
nor U16577 (N_16577,N_15090,N_15367);
and U16578 (N_16578,N_15203,N_15870);
nand U16579 (N_16579,N_15257,N_15520);
xor U16580 (N_16580,N_15984,N_15245);
nor U16581 (N_16581,N_15191,N_15608);
and U16582 (N_16582,N_15739,N_15345);
xor U16583 (N_16583,N_15309,N_15414);
and U16584 (N_16584,N_15304,N_15143);
and U16585 (N_16585,N_15488,N_15434);
nor U16586 (N_16586,N_15530,N_15372);
nand U16587 (N_16587,N_15677,N_15267);
or U16588 (N_16588,N_15336,N_15295);
or U16589 (N_16589,N_15643,N_15229);
xor U16590 (N_16590,N_15905,N_15155);
or U16591 (N_16591,N_15815,N_15221);
nor U16592 (N_16592,N_15588,N_15571);
and U16593 (N_16593,N_15635,N_15675);
or U16594 (N_16594,N_15312,N_15510);
and U16595 (N_16595,N_15119,N_15361);
nor U16596 (N_16596,N_15116,N_15724);
nor U16597 (N_16597,N_15958,N_15816);
nand U16598 (N_16598,N_15391,N_15646);
nor U16599 (N_16599,N_15503,N_15657);
nand U16600 (N_16600,N_15271,N_15456);
nand U16601 (N_16601,N_15809,N_15413);
nor U16602 (N_16602,N_15186,N_15958);
and U16603 (N_16603,N_15298,N_15161);
nand U16604 (N_16604,N_15224,N_15048);
nor U16605 (N_16605,N_15195,N_15392);
xnor U16606 (N_16606,N_15568,N_15709);
or U16607 (N_16607,N_15173,N_15415);
xor U16608 (N_16608,N_15899,N_15457);
or U16609 (N_16609,N_15492,N_15306);
nand U16610 (N_16610,N_15381,N_15835);
or U16611 (N_16611,N_15273,N_15388);
nor U16612 (N_16612,N_15338,N_15757);
or U16613 (N_16613,N_15730,N_15478);
or U16614 (N_16614,N_15064,N_15449);
or U16615 (N_16615,N_15758,N_15303);
nand U16616 (N_16616,N_15340,N_15970);
or U16617 (N_16617,N_15612,N_15822);
nand U16618 (N_16618,N_15018,N_15334);
xor U16619 (N_16619,N_15562,N_15676);
xor U16620 (N_16620,N_15462,N_15751);
or U16621 (N_16621,N_15370,N_15952);
or U16622 (N_16622,N_15003,N_15491);
nor U16623 (N_16623,N_15418,N_15129);
and U16624 (N_16624,N_15985,N_15016);
and U16625 (N_16625,N_15727,N_15646);
and U16626 (N_16626,N_15681,N_15657);
nor U16627 (N_16627,N_15751,N_15431);
nor U16628 (N_16628,N_15613,N_15829);
and U16629 (N_16629,N_15095,N_15864);
xnor U16630 (N_16630,N_15753,N_15862);
or U16631 (N_16631,N_15022,N_15282);
nor U16632 (N_16632,N_15018,N_15365);
or U16633 (N_16633,N_15156,N_15889);
and U16634 (N_16634,N_15846,N_15040);
nor U16635 (N_16635,N_15898,N_15378);
nor U16636 (N_16636,N_15474,N_15972);
xor U16637 (N_16637,N_15361,N_15146);
nor U16638 (N_16638,N_15341,N_15670);
or U16639 (N_16639,N_15736,N_15618);
xnor U16640 (N_16640,N_15646,N_15017);
nor U16641 (N_16641,N_15094,N_15993);
and U16642 (N_16642,N_15971,N_15315);
and U16643 (N_16643,N_15218,N_15290);
and U16644 (N_16644,N_15741,N_15595);
or U16645 (N_16645,N_15060,N_15618);
or U16646 (N_16646,N_15432,N_15703);
and U16647 (N_16647,N_15162,N_15320);
and U16648 (N_16648,N_15649,N_15134);
xnor U16649 (N_16649,N_15947,N_15635);
and U16650 (N_16650,N_15278,N_15710);
and U16651 (N_16651,N_15571,N_15094);
or U16652 (N_16652,N_15717,N_15655);
nand U16653 (N_16653,N_15449,N_15075);
nor U16654 (N_16654,N_15440,N_15045);
nand U16655 (N_16655,N_15770,N_15276);
or U16656 (N_16656,N_15618,N_15262);
xor U16657 (N_16657,N_15486,N_15959);
or U16658 (N_16658,N_15824,N_15805);
or U16659 (N_16659,N_15097,N_15885);
or U16660 (N_16660,N_15531,N_15080);
nor U16661 (N_16661,N_15942,N_15865);
or U16662 (N_16662,N_15713,N_15583);
nand U16663 (N_16663,N_15551,N_15165);
xnor U16664 (N_16664,N_15591,N_15932);
nand U16665 (N_16665,N_15836,N_15487);
or U16666 (N_16666,N_15632,N_15217);
nor U16667 (N_16667,N_15007,N_15803);
nor U16668 (N_16668,N_15535,N_15001);
or U16669 (N_16669,N_15552,N_15056);
and U16670 (N_16670,N_15718,N_15505);
or U16671 (N_16671,N_15066,N_15757);
and U16672 (N_16672,N_15314,N_15238);
nor U16673 (N_16673,N_15926,N_15966);
xnor U16674 (N_16674,N_15370,N_15308);
nand U16675 (N_16675,N_15373,N_15468);
or U16676 (N_16676,N_15525,N_15888);
nor U16677 (N_16677,N_15626,N_15535);
xor U16678 (N_16678,N_15378,N_15371);
and U16679 (N_16679,N_15313,N_15512);
nand U16680 (N_16680,N_15187,N_15613);
nand U16681 (N_16681,N_15500,N_15795);
or U16682 (N_16682,N_15188,N_15635);
or U16683 (N_16683,N_15280,N_15686);
xor U16684 (N_16684,N_15949,N_15189);
nor U16685 (N_16685,N_15288,N_15514);
nand U16686 (N_16686,N_15659,N_15735);
xor U16687 (N_16687,N_15755,N_15692);
nor U16688 (N_16688,N_15311,N_15838);
nand U16689 (N_16689,N_15794,N_15897);
or U16690 (N_16690,N_15209,N_15635);
or U16691 (N_16691,N_15230,N_15595);
or U16692 (N_16692,N_15030,N_15708);
nor U16693 (N_16693,N_15241,N_15103);
xnor U16694 (N_16694,N_15732,N_15590);
and U16695 (N_16695,N_15434,N_15894);
nor U16696 (N_16696,N_15467,N_15465);
or U16697 (N_16697,N_15876,N_15322);
nand U16698 (N_16698,N_15604,N_15506);
nor U16699 (N_16699,N_15911,N_15240);
nor U16700 (N_16700,N_15877,N_15065);
or U16701 (N_16701,N_15548,N_15686);
or U16702 (N_16702,N_15645,N_15898);
nand U16703 (N_16703,N_15649,N_15459);
nor U16704 (N_16704,N_15447,N_15409);
or U16705 (N_16705,N_15388,N_15059);
xnor U16706 (N_16706,N_15901,N_15520);
and U16707 (N_16707,N_15290,N_15608);
nand U16708 (N_16708,N_15702,N_15657);
or U16709 (N_16709,N_15928,N_15053);
nor U16710 (N_16710,N_15189,N_15006);
nand U16711 (N_16711,N_15049,N_15142);
and U16712 (N_16712,N_15474,N_15354);
xor U16713 (N_16713,N_15157,N_15351);
or U16714 (N_16714,N_15007,N_15241);
nand U16715 (N_16715,N_15359,N_15455);
xor U16716 (N_16716,N_15724,N_15002);
nand U16717 (N_16717,N_15464,N_15189);
xor U16718 (N_16718,N_15586,N_15473);
xor U16719 (N_16719,N_15931,N_15223);
and U16720 (N_16720,N_15585,N_15540);
xor U16721 (N_16721,N_15325,N_15642);
and U16722 (N_16722,N_15412,N_15606);
nand U16723 (N_16723,N_15987,N_15849);
nand U16724 (N_16724,N_15065,N_15767);
xor U16725 (N_16725,N_15045,N_15681);
nand U16726 (N_16726,N_15217,N_15593);
nand U16727 (N_16727,N_15495,N_15999);
and U16728 (N_16728,N_15870,N_15616);
or U16729 (N_16729,N_15691,N_15675);
xor U16730 (N_16730,N_15476,N_15547);
nor U16731 (N_16731,N_15787,N_15649);
or U16732 (N_16732,N_15085,N_15856);
xor U16733 (N_16733,N_15358,N_15001);
and U16734 (N_16734,N_15734,N_15298);
nor U16735 (N_16735,N_15832,N_15133);
xnor U16736 (N_16736,N_15803,N_15302);
xor U16737 (N_16737,N_15013,N_15812);
nand U16738 (N_16738,N_15530,N_15731);
nand U16739 (N_16739,N_15234,N_15836);
xnor U16740 (N_16740,N_15001,N_15040);
nand U16741 (N_16741,N_15855,N_15092);
nand U16742 (N_16742,N_15118,N_15133);
nor U16743 (N_16743,N_15733,N_15197);
xnor U16744 (N_16744,N_15871,N_15314);
and U16745 (N_16745,N_15644,N_15667);
and U16746 (N_16746,N_15495,N_15391);
xnor U16747 (N_16747,N_15562,N_15205);
xnor U16748 (N_16748,N_15109,N_15451);
and U16749 (N_16749,N_15099,N_15698);
or U16750 (N_16750,N_15856,N_15975);
or U16751 (N_16751,N_15996,N_15257);
and U16752 (N_16752,N_15309,N_15343);
xor U16753 (N_16753,N_15750,N_15164);
nand U16754 (N_16754,N_15319,N_15998);
nand U16755 (N_16755,N_15339,N_15839);
and U16756 (N_16756,N_15310,N_15629);
and U16757 (N_16757,N_15935,N_15844);
nand U16758 (N_16758,N_15466,N_15367);
nand U16759 (N_16759,N_15741,N_15983);
or U16760 (N_16760,N_15058,N_15093);
and U16761 (N_16761,N_15820,N_15715);
and U16762 (N_16762,N_15582,N_15097);
nand U16763 (N_16763,N_15312,N_15756);
or U16764 (N_16764,N_15321,N_15738);
or U16765 (N_16765,N_15668,N_15413);
xor U16766 (N_16766,N_15056,N_15254);
or U16767 (N_16767,N_15675,N_15437);
xnor U16768 (N_16768,N_15916,N_15669);
and U16769 (N_16769,N_15710,N_15406);
xnor U16770 (N_16770,N_15783,N_15703);
xnor U16771 (N_16771,N_15268,N_15644);
or U16772 (N_16772,N_15274,N_15723);
nor U16773 (N_16773,N_15825,N_15002);
xor U16774 (N_16774,N_15495,N_15962);
nand U16775 (N_16775,N_15179,N_15860);
or U16776 (N_16776,N_15691,N_15758);
nand U16777 (N_16777,N_15142,N_15905);
nand U16778 (N_16778,N_15623,N_15076);
and U16779 (N_16779,N_15687,N_15479);
nand U16780 (N_16780,N_15652,N_15692);
nand U16781 (N_16781,N_15111,N_15521);
nand U16782 (N_16782,N_15526,N_15936);
or U16783 (N_16783,N_15405,N_15564);
xor U16784 (N_16784,N_15551,N_15627);
and U16785 (N_16785,N_15294,N_15635);
and U16786 (N_16786,N_15420,N_15799);
or U16787 (N_16787,N_15302,N_15162);
nand U16788 (N_16788,N_15865,N_15236);
nand U16789 (N_16789,N_15961,N_15015);
nand U16790 (N_16790,N_15667,N_15634);
or U16791 (N_16791,N_15752,N_15785);
nor U16792 (N_16792,N_15730,N_15271);
xor U16793 (N_16793,N_15782,N_15630);
or U16794 (N_16794,N_15698,N_15269);
nand U16795 (N_16795,N_15342,N_15561);
or U16796 (N_16796,N_15607,N_15093);
xor U16797 (N_16797,N_15217,N_15223);
nand U16798 (N_16798,N_15031,N_15804);
nor U16799 (N_16799,N_15175,N_15123);
nor U16800 (N_16800,N_15308,N_15670);
nand U16801 (N_16801,N_15259,N_15124);
xnor U16802 (N_16802,N_15087,N_15408);
xnor U16803 (N_16803,N_15004,N_15342);
nor U16804 (N_16804,N_15457,N_15152);
nand U16805 (N_16805,N_15613,N_15694);
nand U16806 (N_16806,N_15637,N_15011);
or U16807 (N_16807,N_15466,N_15301);
nor U16808 (N_16808,N_15260,N_15475);
and U16809 (N_16809,N_15128,N_15982);
and U16810 (N_16810,N_15034,N_15748);
nor U16811 (N_16811,N_15905,N_15112);
or U16812 (N_16812,N_15105,N_15484);
xnor U16813 (N_16813,N_15568,N_15159);
and U16814 (N_16814,N_15874,N_15365);
or U16815 (N_16815,N_15264,N_15710);
and U16816 (N_16816,N_15657,N_15393);
and U16817 (N_16817,N_15357,N_15535);
nor U16818 (N_16818,N_15408,N_15165);
or U16819 (N_16819,N_15419,N_15405);
xor U16820 (N_16820,N_15322,N_15696);
xnor U16821 (N_16821,N_15164,N_15539);
nand U16822 (N_16822,N_15265,N_15748);
or U16823 (N_16823,N_15106,N_15714);
xor U16824 (N_16824,N_15744,N_15835);
nand U16825 (N_16825,N_15175,N_15506);
xor U16826 (N_16826,N_15993,N_15544);
or U16827 (N_16827,N_15147,N_15860);
xor U16828 (N_16828,N_15289,N_15391);
nor U16829 (N_16829,N_15825,N_15259);
or U16830 (N_16830,N_15447,N_15771);
xor U16831 (N_16831,N_15151,N_15341);
nand U16832 (N_16832,N_15584,N_15522);
and U16833 (N_16833,N_15022,N_15123);
nand U16834 (N_16834,N_15976,N_15699);
nand U16835 (N_16835,N_15108,N_15258);
xnor U16836 (N_16836,N_15586,N_15545);
xnor U16837 (N_16837,N_15424,N_15213);
and U16838 (N_16838,N_15092,N_15645);
and U16839 (N_16839,N_15564,N_15910);
nand U16840 (N_16840,N_15211,N_15133);
nand U16841 (N_16841,N_15490,N_15098);
and U16842 (N_16842,N_15529,N_15722);
and U16843 (N_16843,N_15410,N_15080);
or U16844 (N_16844,N_15546,N_15392);
nand U16845 (N_16845,N_15423,N_15670);
nor U16846 (N_16846,N_15467,N_15395);
nand U16847 (N_16847,N_15142,N_15586);
xnor U16848 (N_16848,N_15575,N_15237);
nand U16849 (N_16849,N_15099,N_15244);
or U16850 (N_16850,N_15717,N_15402);
xor U16851 (N_16851,N_15470,N_15165);
nand U16852 (N_16852,N_15355,N_15081);
nor U16853 (N_16853,N_15758,N_15142);
or U16854 (N_16854,N_15685,N_15642);
or U16855 (N_16855,N_15311,N_15119);
nand U16856 (N_16856,N_15889,N_15676);
and U16857 (N_16857,N_15646,N_15597);
xnor U16858 (N_16858,N_15697,N_15751);
or U16859 (N_16859,N_15937,N_15228);
or U16860 (N_16860,N_15805,N_15435);
xnor U16861 (N_16861,N_15053,N_15908);
or U16862 (N_16862,N_15550,N_15456);
nor U16863 (N_16863,N_15888,N_15694);
nor U16864 (N_16864,N_15296,N_15863);
or U16865 (N_16865,N_15444,N_15619);
and U16866 (N_16866,N_15192,N_15284);
nand U16867 (N_16867,N_15769,N_15861);
nor U16868 (N_16868,N_15315,N_15942);
xnor U16869 (N_16869,N_15703,N_15618);
and U16870 (N_16870,N_15666,N_15516);
or U16871 (N_16871,N_15493,N_15809);
xnor U16872 (N_16872,N_15151,N_15208);
or U16873 (N_16873,N_15436,N_15272);
nor U16874 (N_16874,N_15895,N_15985);
xor U16875 (N_16875,N_15754,N_15634);
and U16876 (N_16876,N_15850,N_15471);
nand U16877 (N_16877,N_15584,N_15324);
nor U16878 (N_16878,N_15335,N_15911);
and U16879 (N_16879,N_15834,N_15703);
xnor U16880 (N_16880,N_15175,N_15683);
nor U16881 (N_16881,N_15472,N_15618);
xnor U16882 (N_16882,N_15299,N_15710);
xnor U16883 (N_16883,N_15698,N_15827);
and U16884 (N_16884,N_15147,N_15592);
xnor U16885 (N_16885,N_15059,N_15223);
nor U16886 (N_16886,N_15770,N_15605);
xnor U16887 (N_16887,N_15227,N_15515);
and U16888 (N_16888,N_15696,N_15984);
nor U16889 (N_16889,N_15856,N_15550);
nor U16890 (N_16890,N_15290,N_15802);
nand U16891 (N_16891,N_15268,N_15786);
or U16892 (N_16892,N_15235,N_15244);
or U16893 (N_16893,N_15384,N_15243);
or U16894 (N_16894,N_15954,N_15044);
and U16895 (N_16895,N_15239,N_15512);
nor U16896 (N_16896,N_15241,N_15569);
nand U16897 (N_16897,N_15479,N_15377);
xnor U16898 (N_16898,N_15251,N_15375);
nor U16899 (N_16899,N_15576,N_15648);
nor U16900 (N_16900,N_15290,N_15803);
nor U16901 (N_16901,N_15528,N_15651);
nor U16902 (N_16902,N_15599,N_15500);
and U16903 (N_16903,N_15506,N_15489);
and U16904 (N_16904,N_15484,N_15101);
and U16905 (N_16905,N_15857,N_15257);
xor U16906 (N_16906,N_15398,N_15402);
xor U16907 (N_16907,N_15332,N_15659);
nor U16908 (N_16908,N_15174,N_15029);
xor U16909 (N_16909,N_15242,N_15970);
nand U16910 (N_16910,N_15212,N_15224);
nor U16911 (N_16911,N_15694,N_15219);
nor U16912 (N_16912,N_15032,N_15920);
or U16913 (N_16913,N_15599,N_15404);
xnor U16914 (N_16914,N_15901,N_15362);
xor U16915 (N_16915,N_15927,N_15094);
or U16916 (N_16916,N_15823,N_15464);
and U16917 (N_16917,N_15452,N_15030);
nand U16918 (N_16918,N_15294,N_15274);
xnor U16919 (N_16919,N_15706,N_15354);
nand U16920 (N_16920,N_15770,N_15786);
and U16921 (N_16921,N_15017,N_15089);
and U16922 (N_16922,N_15822,N_15664);
nand U16923 (N_16923,N_15295,N_15689);
xor U16924 (N_16924,N_15946,N_15600);
xnor U16925 (N_16925,N_15007,N_15696);
and U16926 (N_16926,N_15028,N_15358);
and U16927 (N_16927,N_15201,N_15755);
nor U16928 (N_16928,N_15540,N_15754);
nor U16929 (N_16929,N_15452,N_15393);
xnor U16930 (N_16930,N_15954,N_15072);
nor U16931 (N_16931,N_15294,N_15577);
or U16932 (N_16932,N_15681,N_15579);
and U16933 (N_16933,N_15606,N_15965);
or U16934 (N_16934,N_15205,N_15329);
xnor U16935 (N_16935,N_15942,N_15449);
xnor U16936 (N_16936,N_15788,N_15198);
nor U16937 (N_16937,N_15745,N_15205);
or U16938 (N_16938,N_15185,N_15217);
nand U16939 (N_16939,N_15526,N_15177);
nor U16940 (N_16940,N_15368,N_15046);
xor U16941 (N_16941,N_15544,N_15668);
nand U16942 (N_16942,N_15464,N_15236);
nand U16943 (N_16943,N_15635,N_15610);
and U16944 (N_16944,N_15203,N_15786);
xor U16945 (N_16945,N_15536,N_15336);
nor U16946 (N_16946,N_15054,N_15792);
nand U16947 (N_16947,N_15650,N_15353);
nor U16948 (N_16948,N_15208,N_15683);
or U16949 (N_16949,N_15616,N_15517);
and U16950 (N_16950,N_15280,N_15951);
or U16951 (N_16951,N_15216,N_15526);
xnor U16952 (N_16952,N_15433,N_15726);
nand U16953 (N_16953,N_15289,N_15264);
or U16954 (N_16954,N_15919,N_15898);
or U16955 (N_16955,N_15691,N_15506);
or U16956 (N_16956,N_15716,N_15756);
nor U16957 (N_16957,N_15829,N_15060);
xnor U16958 (N_16958,N_15787,N_15953);
and U16959 (N_16959,N_15801,N_15318);
or U16960 (N_16960,N_15526,N_15004);
xor U16961 (N_16961,N_15060,N_15981);
xor U16962 (N_16962,N_15756,N_15742);
nand U16963 (N_16963,N_15461,N_15066);
and U16964 (N_16964,N_15154,N_15533);
nand U16965 (N_16965,N_15148,N_15771);
nor U16966 (N_16966,N_15480,N_15627);
and U16967 (N_16967,N_15603,N_15629);
and U16968 (N_16968,N_15939,N_15496);
or U16969 (N_16969,N_15472,N_15084);
nand U16970 (N_16970,N_15585,N_15300);
nor U16971 (N_16971,N_15877,N_15435);
xnor U16972 (N_16972,N_15881,N_15420);
nor U16973 (N_16973,N_15253,N_15163);
nand U16974 (N_16974,N_15790,N_15522);
and U16975 (N_16975,N_15366,N_15994);
xor U16976 (N_16976,N_15364,N_15450);
nand U16977 (N_16977,N_15671,N_15031);
xor U16978 (N_16978,N_15644,N_15221);
xor U16979 (N_16979,N_15219,N_15560);
and U16980 (N_16980,N_15021,N_15610);
nor U16981 (N_16981,N_15527,N_15866);
xor U16982 (N_16982,N_15626,N_15791);
xor U16983 (N_16983,N_15044,N_15602);
or U16984 (N_16984,N_15365,N_15788);
or U16985 (N_16985,N_15085,N_15940);
nand U16986 (N_16986,N_15853,N_15630);
nand U16987 (N_16987,N_15386,N_15953);
nand U16988 (N_16988,N_15257,N_15132);
nor U16989 (N_16989,N_15574,N_15998);
and U16990 (N_16990,N_15253,N_15077);
xnor U16991 (N_16991,N_15254,N_15765);
and U16992 (N_16992,N_15351,N_15890);
or U16993 (N_16993,N_15453,N_15034);
and U16994 (N_16994,N_15759,N_15454);
xnor U16995 (N_16995,N_15395,N_15824);
nor U16996 (N_16996,N_15596,N_15180);
or U16997 (N_16997,N_15443,N_15874);
or U16998 (N_16998,N_15825,N_15402);
nor U16999 (N_16999,N_15178,N_15464);
and U17000 (N_17000,N_16178,N_16062);
or U17001 (N_17001,N_16520,N_16260);
xor U17002 (N_17002,N_16265,N_16943);
or U17003 (N_17003,N_16866,N_16761);
xnor U17004 (N_17004,N_16810,N_16151);
and U17005 (N_17005,N_16752,N_16446);
nand U17006 (N_17006,N_16863,N_16014);
and U17007 (N_17007,N_16466,N_16921);
nor U17008 (N_17008,N_16830,N_16419);
xnor U17009 (N_17009,N_16267,N_16398);
or U17010 (N_17010,N_16378,N_16769);
and U17011 (N_17011,N_16462,N_16052);
or U17012 (N_17012,N_16624,N_16990);
or U17013 (N_17013,N_16524,N_16424);
nor U17014 (N_17014,N_16591,N_16428);
nor U17015 (N_17015,N_16147,N_16045);
or U17016 (N_17016,N_16031,N_16796);
or U17017 (N_17017,N_16289,N_16001);
nand U17018 (N_17018,N_16359,N_16538);
xor U17019 (N_17019,N_16926,N_16517);
xor U17020 (N_17020,N_16215,N_16636);
nor U17021 (N_17021,N_16756,N_16500);
and U17022 (N_17022,N_16741,N_16328);
nand U17023 (N_17023,N_16831,N_16518);
nor U17024 (N_17024,N_16808,N_16406);
and U17025 (N_17025,N_16806,N_16046);
nand U17026 (N_17026,N_16280,N_16374);
and U17027 (N_17027,N_16997,N_16129);
nand U17028 (N_17028,N_16706,N_16091);
and U17029 (N_17029,N_16043,N_16819);
xor U17030 (N_17030,N_16308,N_16656);
or U17031 (N_17031,N_16481,N_16627);
nand U17032 (N_17032,N_16931,N_16198);
xor U17033 (N_17033,N_16012,N_16329);
and U17034 (N_17034,N_16634,N_16357);
nand U17035 (N_17035,N_16017,N_16895);
nor U17036 (N_17036,N_16156,N_16413);
nor U17037 (N_17037,N_16107,N_16922);
or U17038 (N_17038,N_16429,N_16890);
or U17039 (N_17039,N_16897,N_16870);
xor U17040 (N_17040,N_16675,N_16586);
xnor U17041 (N_17041,N_16102,N_16485);
xor U17042 (N_17042,N_16900,N_16662);
xnor U17043 (N_17043,N_16940,N_16050);
nor U17044 (N_17044,N_16944,N_16281);
or U17045 (N_17045,N_16904,N_16303);
nand U17046 (N_17046,N_16099,N_16009);
nand U17047 (N_17047,N_16201,N_16425);
and U17048 (N_17048,N_16623,N_16019);
and U17049 (N_17049,N_16221,N_16165);
and U17050 (N_17050,N_16674,N_16189);
or U17051 (N_17051,N_16692,N_16381);
xnor U17052 (N_17052,N_16047,N_16440);
xor U17053 (N_17053,N_16456,N_16002);
and U17054 (N_17054,N_16746,N_16261);
and U17055 (N_17055,N_16074,N_16592);
nor U17056 (N_17056,N_16384,N_16392);
nor U17057 (N_17057,N_16506,N_16034);
nand U17058 (N_17058,N_16821,N_16210);
nor U17059 (N_17059,N_16803,N_16633);
and U17060 (N_17060,N_16909,N_16984);
nand U17061 (N_17061,N_16799,N_16710);
or U17062 (N_17062,N_16783,N_16118);
nor U17063 (N_17063,N_16457,N_16582);
or U17064 (N_17064,N_16812,N_16651);
or U17065 (N_17065,N_16575,N_16093);
or U17066 (N_17066,N_16365,N_16287);
nor U17067 (N_17067,N_16186,N_16266);
nor U17068 (N_17068,N_16055,N_16120);
nand U17069 (N_17069,N_16354,N_16076);
and U17070 (N_17070,N_16511,N_16671);
or U17071 (N_17071,N_16730,N_16916);
xnor U17072 (N_17072,N_16404,N_16113);
xor U17073 (N_17073,N_16753,N_16209);
nand U17074 (N_17074,N_16386,N_16548);
nand U17075 (N_17075,N_16484,N_16036);
nand U17076 (N_17076,N_16394,N_16935);
nand U17077 (N_17077,N_16859,N_16557);
xor U17078 (N_17078,N_16991,N_16884);
nor U17079 (N_17079,N_16180,N_16199);
and U17080 (N_17080,N_16134,N_16427);
or U17081 (N_17081,N_16324,N_16397);
nor U17082 (N_17082,N_16738,N_16925);
and U17083 (N_17083,N_16389,N_16809);
nand U17084 (N_17084,N_16259,N_16792);
nor U17085 (N_17085,N_16297,N_16025);
nor U17086 (N_17086,N_16436,N_16680);
nand U17087 (N_17087,N_16049,N_16593);
and U17088 (N_17088,N_16578,N_16679);
nor U17089 (N_17089,N_16691,N_16660);
or U17090 (N_17090,N_16021,N_16471);
nor U17091 (N_17091,N_16825,N_16777);
or U17092 (N_17092,N_16316,N_16455);
xnor U17093 (N_17093,N_16495,N_16733);
nor U17094 (N_17094,N_16066,N_16805);
and U17095 (N_17095,N_16232,N_16382);
nand U17096 (N_17096,N_16823,N_16696);
nand U17097 (N_17097,N_16993,N_16961);
or U17098 (N_17098,N_16764,N_16949);
nor U17099 (N_17099,N_16191,N_16228);
nor U17100 (N_17100,N_16835,N_16659);
or U17101 (N_17101,N_16095,N_16123);
xnor U17102 (N_17102,N_16273,N_16204);
nand U17103 (N_17103,N_16652,N_16958);
nor U17104 (N_17104,N_16370,N_16559);
and U17105 (N_17105,N_16326,N_16168);
or U17106 (N_17106,N_16644,N_16698);
nand U17107 (N_17107,N_16778,N_16040);
or U17108 (N_17108,N_16286,N_16820);
nor U17109 (N_17109,N_16807,N_16051);
nor U17110 (N_17110,N_16108,N_16097);
and U17111 (N_17111,N_16431,N_16241);
nor U17112 (N_17112,N_16525,N_16587);
and U17113 (N_17113,N_16405,N_16702);
xor U17114 (N_17114,N_16537,N_16829);
and U17115 (N_17115,N_16774,N_16448);
or U17116 (N_17116,N_16162,N_16463);
nor U17117 (N_17117,N_16639,N_16504);
xor U17118 (N_17118,N_16875,N_16514);
nand U17119 (N_17119,N_16606,N_16844);
and U17120 (N_17120,N_16860,N_16337);
nand U17121 (N_17121,N_16505,N_16409);
and U17122 (N_17122,N_16138,N_16729);
and U17123 (N_17123,N_16785,N_16945);
or U17124 (N_17124,N_16689,N_16125);
nand U17125 (N_17125,N_16197,N_16258);
xnor U17126 (N_17126,N_16565,N_16556);
and U17127 (N_17127,N_16747,N_16217);
or U17128 (N_17128,N_16270,N_16497);
xnor U17129 (N_17129,N_16772,N_16969);
xor U17130 (N_17130,N_16137,N_16968);
xnor U17131 (N_17131,N_16982,N_16194);
or U17132 (N_17132,N_16220,N_16699);
or U17133 (N_17133,N_16615,N_16004);
nand U17134 (N_17134,N_16603,N_16713);
nor U17135 (N_17135,N_16986,N_16219);
and U17136 (N_17136,N_16663,N_16084);
xor U17137 (N_17137,N_16832,N_16317);
xor U17138 (N_17138,N_16714,N_16187);
and U17139 (N_17139,N_16563,N_16192);
and U17140 (N_17140,N_16053,N_16254);
or U17141 (N_17141,N_16865,N_16590);
and U17142 (N_17142,N_16459,N_16833);
nor U17143 (N_17143,N_16535,N_16275);
and U17144 (N_17144,N_16750,N_16452);
xnor U17145 (N_17145,N_16722,N_16331);
or U17146 (N_17146,N_16848,N_16595);
and U17147 (N_17147,N_16348,N_16490);
nand U17148 (N_17148,N_16233,N_16414);
or U17149 (N_17149,N_16964,N_16762);
and U17150 (N_17150,N_16003,N_16748);
nand U17151 (N_17151,N_16188,N_16309);
and U17152 (N_17152,N_16248,N_16421);
xor U17153 (N_17153,N_16754,N_16979);
nor U17154 (N_17154,N_16387,N_16313);
nor U17155 (N_17155,N_16190,N_16090);
or U17156 (N_17156,N_16927,N_16127);
nand U17157 (N_17157,N_16901,N_16767);
nor U17158 (N_17158,N_16862,N_16549);
nand U17159 (N_17159,N_16024,N_16980);
xor U17160 (N_17160,N_16770,N_16006);
nor U17161 (N_17161,N_16998,N_16344);
or U17162 (N_17162,N_16728,N_16522);
xnor U17163 (N_17163,N_16030,N_16282);
nor U17164 (N_17164,N_16116,N_16298);
nand U17165 (N_17165,N_16887,N_16475);
and U17166 (N_17166,N_16487,N_16170);
xor U17167 (N_17167,N_16801,N_16655);
nand U17168 (N_17168,N_16195,N_16513);
or U17169 (N_17169,N_16584,N_16323);
nor U17170 (N_17170,N_16407,N_16938);
xnor U17171 (N_17171,N_16963,N_16044);
or U17172 (N_17172,N_16602,N_16932);
or U17173 (N_17173,N_16503,N_16380);
nor U17174 (N_17174,N_16683,N_16245);
xnor U17175 (N_17175,N_16027,N_16470);
nor U17176 (N_17176,N_16143,N_16760);
and U17177 (N_17177,N_16942,N_16898);
xor U17178 (N_17178,N_16972,N_16977);
xor U17179 (N_17179,N_16131,N_16061);
nand U17180 (N_17180,N_16521,N_16891);
or U17181 (N_17181,N_16672,N_16111);
or U17182 (N_17182,N_16849,N_16850);
nor U17183 (N_17183,N_16164,N_16202);
xnor U17184 (N_17184,N_16826,N_16564);
xnor U17185 (N_17185,N_16939,N_16872);
or U17186 (N_17186,N_16333,N_16492);
nor U17187 (N_17187,N_16928,N_16569);
nand U17188 (N_17188,N_16847,N_16836);
and U17189 (N_17189,N_16554,N_16447);
nand U17190 (N_17190,N_16902,N_16724);
xnor U17191 (N_17191,N_16815,N_16650);
nand U17192 (N_17192,N_16391,N_16717);
or U17193 (N_17193,N_16896,N_16811);
and U17194 (N_17194,N_16420,N_16923);
nand U17195 (N_17195,N_16816,N_16161);
nand U17196 (N_17196,N_16987,N_16976);
nand U17197 (N_17197,N_16960,N_16775);
nand U17198 (N_17198,N_16577,N_16876);
and U17199 (N_17199,N_16060,N_16899);
nand U17200 (N_17200,N_16782,N_16881);
nor U17201 (N_17201,N_16903,N_16566);
and U17202 (N_17202,N_16817,N_16828);
or U17203 (N_17203,N_16824,N_16172);
and U17204 (N_17204,N_16070,N_16843);
or U17205 (N_17205,N_16786,N_16618);
nor U17206 (N_17206,N_16892,N_16141);
nor U17207 (N_17207,N_16955,N_16794);
and U17208 (N_17208,N_16868,N_16718);
and U17209 (N_17209,N_16442,N_16948);
and U17210 (N_17210,N_16244,N_16920);
xnor U17211 (N_17211,N_16894,N_16771);
nand U17212 (N_17212,N_16768,N_16150);
and U17213 (N_17213,N_16763,N_16965);
nand U17214 (N_17214,N_16755,N_16112);
xnor U17215 (N_17215,N_16914,N_16562);
xor U17216 (N_17216,N_16915,N_16314);
and U17217 (N_17217,N_16104,N_16458);
and U17218 (N_17218,N_16700,N_16736);
nand U17219 (N_17219,N_16632,N_16597);
nor U17220 (N_17220,N_16364,N_16332);
and U17221 (N_17221,N_16598,N_16616);
xnor U17222 (N_17222,N_16918,N_16687);
nand U17223 (N_17223,N_16124,N_16276);
or U17224 (N_17224,N_16533,N_16797);
xnor U17225 (N_17225,N_16379,N_16092);
xnor U17226 (N_17226,N_16751,N_16115);
nand U17227 (N_17227,N_16100,N_16638);
and U17228 (N_17228,N_16039,N_16605);
nor U17229 (N_17229,N_16827,N_16515);
nor U17230 (N_17230,N_16128,N_16010);
nand U17231 (N_17231,N_16376,N_16437);
xnor U17232 (N_17232,N_16218,N_16295);
nand U17233 (N_17233,N_16681,N_16527);
nand U17234 (N_17234,N_16184,N_16101);
xnor U17235 (N_17235,N_16377,N_16403);
and U17236 (N_17236,N_16449,N_16739);
xor U17237 (N_17237,N_16529,N_16493);
and U17238 (N_17238,N_16056,N_16658);
xnor U17239 (N_17239,N_16476,N_16973);
and U17240 (N_17240,N_16396,N_16629);
or U17241 (N_17241,N_16791,N_16393);
or U17242 (N_17242,N_16838,N_16315);
or U17243 (N_17243,N_16139,N_16589);
nand U17244 (N_17244,N_16543,N_16934);
and U17245 (N_17245,N_16686,N_16028);
xor U17246 (N_17246,N_16356,N_16941);
nand U17247 (N_17247,N_16526,N_16426);
or U17248 (N_17248,N_16878,N_16226);
nand U17249 (N_17249,N_16306,N_16149);
or U17250 (N_17250,N_16212,N_16880);
nor U17251 (N_17251,N_16321,N_16041);
nand U17252 (N_17252,N_16999,N_16585);
or U17253 (N_17253,N_16647,N_16798);
xnor U17254 (N_17254,N_16694,N_16507);
and U17255 (N_17255,N_16469,N_16257);
nand U17256 (N_17256,N_16453,N_16290);
nor U17257 (N_17257,N_16974,N_16117);
or U17258 (N_17258,N_16087,N_16789);
nor U17259 (N_17259,N_16532,N_16110);
nor U17260 (N_17260,N_16292,N_16417);
or U17261 (N_17261,N_16441,N_16869);
or U17262 (N_17262,N_16358,N_16678);
and U17263 (N_17263,N_16708,N_16223);
xor U17264 (N_17264,N_16693,N_16677);
xor U17265 (N_17265,N_16203,N_16804);
and U17266 (N_17266,N_16947,N_16793);
nor U17267 (N_17267,N_16152,N_16278);
xor U17268 (N_17268,N_16343,N_16959);
and U17269 (N_17269,N_16547,N_16068);
xnor U17270 (N_17270,N_16300,N_16073);
nor U17271 (N_17271,N_16995,N_16008);
xnor U17272 (N_17272,N_16573,N_16766);
xnor U17273 (N_17273,N_16193,N_16788);
nand U17274 (N_17274,N_16596,N_16874);
or U17275 (N_17275,N_16307,N_16415);
nor U17276 (N_17276,N_16911,N_16322);
or U17277 (N_17277,N_16712,N_16933);
xor U17278 (N_17278,N_16016,N_16035);
nand U17279 (N_17279,N_16734,N_16122);
xnor U17280 (N_17280,N_16345,N_16879);
nand U17281 (N_17281,N_16304,N_16342);
and U17282 (N_17282,N_16867,N_16268);
nand U17283 (N_17283,N_16346,N_16886);
nor U17284 (N_17284,N_16749,N_16888);
and U17285 (N_17285,N_16893,N_16653);
nor U17286 (N_17286,N_16347,N_16235);
nand U17287 (N_17287,N_16086,N_16983);
nand U17288 (N_17288,N_16667,N_16758);
nand U17289 (N_17289,N_16351,N_16171);
or U17290 (N_17290,N_16038,N_16083);
xnor U17291 (N_17291,N_16214,N_16814);
xnor U17292 (N_17292,N_16568,N_16256);
xor U17293 (N_17293,N_16177,N_16970);
nor U17294 (N_17294,N_16697,N_16096);
and U17295 (N_17295,N_16445,N_16023);
nand U17296 (N_17296,N_16502,N_16133);
nor U17297 (N_17297,N_16341,N_16293);
nor U17298 (N_17298,N_16621,N_16580);
xnor U17299 (N_17299,N_16312,N_16858);
nor U17300 (N_17300,N_16033,N_16612);
xor U17301 (N_17301,N_16173,N_16013);
or U17302 (N_17302,N_16661,N_16334);
or U17303 (N_17303,N_16609,N_16930);
or U17304 (N_17304,N_16542,N_16103);
nor U17305 (N_17305,N_16200,N_16400);
nor U17306 (N_17306,N_16558,N_16081);
and U17307 (N_17307,N_16641,N_16026);
and U17308 (N_17308,N_16065,N_16205);
or U17309 (N_17309,N_16160,N_16480);
nand U17310 (N_17310,N_16642,N_16360);
nand U17311 (N_17311,N_16501,N_16119);
and U17312 (N_17312,N_16182,N_16673);
or U17313 (N_17313,N_16418,N_16350);
nand U17314 (N_17314,N_16423,N_16279);
xor U17315 (N_17315,N_16611,N_16508);
or U17316 (N_17316,N_16206,N_16401);
xnor U17317 (N_17317,N_16856,N_16723);
nand U17318 (N_17318,N_16438,N_16936);
and U17319 (N_17319,N_16688,N_16338);
nand U17320 (N_17320,N_16088,N_16029);
nand U17321 (N_17321,N_16631,N_16274);
xor U17322 (N_17322,N_16988,N_16684);
nor U17323 (N_17323,N_16759,N_16283);
nand U17324 (N_17324,N_16058,N_16069);
and U17325 (N_17325,N_16541,N_16250);
xnor U17326 (N_17326,N_16098,N_16208);
or U17327 (N_17327,N_16737,N_16264);
and U17328 (N_17328,N_16546,N_16225);
or U17329 (N_17329,N_16720,N_16601);
and U17330 (N_17330,N_16284,N_16311);
xor U17331 (N_17331,N_16227,N_16363);
nor U17332 (N_17332,N_16478,N_16594);
nand U17333 (N_17333,N_16159,N_16840);
xor U17334 (N_17334,N_16877,N_16599);
and U17335 (N_17335,N_16183,N_16757);
nand U17336 (N_17336,N_16037,N_16837);
nor U17337 (N_17337,N_16552,N_16465);
nor U17338 (N_17338,N_16294,N_16908);
nor U17339 (N_17339,N_16231,N_16079);
nor U17340 (N_17340,N_16721,N_16106);
or U17341 (N_17341,N_16255,N_16048);
xor U17342 (N_17342,N_16105,N_16919);
and U17343 (N_17343,N_16054,N_16145);
or U17344 (N_17344,N_16855,N_16251);
xnor U17345 (N_17345,N_16845,N_16534);
nor U17346 (N_17346,N_16649,N_16956);
xnor U17347 (N_17347,N_16906,N_16422);
or U17348 (N_17348,N_16579,N_16707);
nand U17349 (N_17349,N_16064,N_16645);
xnor U17350 (N_17350,N_16179,N_16953);
and U17351 (N_17351,N_16135,N_16648);
xor U17352 (N_17352,N_16510,N_16285);
or U17353 (N_17353,N_16800,N_16042);
or U17354 (N_17354,N_16236,N_16340);
nand U17355 (N_17355,N_16676,N_16207);
and U17356 (N_17356,N_16082,N_16369);
nor U17357 (N_17357,N_16690,N_16628);
xnor U17358 (N_17358,N_16864,N_16169);
nand U17359 (N_17359,N_16142,N_16301);
and U17360 (N_17360,N_16319,N_16174);
and U17361 (N_17361,N_16408,N_16715);
or U17362 (N_17362,N_16553,N_16157);
and U17363 (N_17363,N_16773,N_16581);
nor U17364 (N_17364,N_16243,N_16496);
or U17365 (N_17365,N_16985,N_16181);
or U17366 (N_17366,N_16460,N_16246);
nand U17367 (N_17367,N_16269,N_16834);
and U17368 (N_17368,N_16032,N_16727);
xor U17369 (N_17369,N_16851,N_16071);
or U17370 (N_17370,N_16946,N_16238);
xor U17371 (N_17371,N_16622,N_16555);
nand U17372 (N_17372,N_16719,N_16604);
nor U17373 (N_17373,N_16011,N_16957);
and U17374 (N_17374,N_16668,N_16528);
nor U17375 (N_17375,N_16637,N_16395);
xor U17376 (N_17376,N_16211,N_16560);
and U17377 (N_17377,N_16572,N_16551);
and U17378 (N_17378,N_16310,N_16952);
nor U17379 (N_17379,N_16372,N_16473);
nor U17380 (N_17380,N_16523,N_16852);
nand U17381 (N_17381,N_16185,N_16853);
nand U17382 (N_17382,N_16402,N_16912);
and U17383 (N_17383,N_16545,N_16873);
or U17384 (N_17384,N_16390,N_16277);
or U17385 (N_17385,N_16614,N_16339);
nand U17386 (N_17386,N_16239,N_16846);
nor U17387 (N_17387,N_16617,N_16608);
nor U17388 (N_17388,N_16917,N_16571);
nand U17389 (N_17389,N_16494,N_16263);
or U17390 (N_17390,N_16635,N_16516);
and U17391 (N_17391,N_16486,N_16388);
xor U17392 (N_17392,N_16253,N_16740);
or U17393 (N_17393,N_16444,N_16163);
nor U17394 (N_17394,N_16540,N_16630);
nand U17395 (N_17395,N_16962,N_16130);
or U17396 (N_17396,N_16654,N_16385);
nand U17397 (N_17397,N_16954,N_16155);
and U17398 (N_17398,N_16355,N_16467);
and U17399 (N_17399,N_16237,N_16726);
nand U17400 (N_17400,N_16709,N_16020);
and U17401 (N_17401,N_16743,N_16230);
nand U17402 (N_17402,N_16703,N_16981);
or U17403 (N_17403,N_16530,N_16583);
and U17404 (N_17404,N_16077,N_16489);
or U17405 (N_17405,N_16059,N_16861);
xnor U17406 (N_17406,N_16779,N_16937);
nor U17407 (N_17407,N_16144,N_16479);
and U17408 (N_17408,N_16154,N_16732);
nor U17409 (N_17409,N_16078,N_16781);
xor U17410 (N_17410,N_16765,N_16539);
nand U17411 (N_17411,N_16252,N_16576);
and U17412 (N_17412,N_16643,N_16291);
xor U17413 (N_17413,N_16913,N_16242);
xnor U17414 (N_17414,N_16005,N_16468);
or U17415 (N_17415,N_16439,N_16366);
or U17416 (N_17416,N_16416,N_16361);
nand U17417 (N_17417,N_16498,N_16491);
and U17418 (N_17418,N_16450,N_16625);
and U17419 (N_17419,N_16302,N_16536);
or U17420 (N_17420,N_16057,N_16213);
or U17421 (N_17421,N_16383,N_16109);
xnor U17422 (N_17422,N_16685,N_16978);
and U17423 (N_17423,N_16362,N_16335);
xnor U17424 (N_17424,N_16249,N_16842);
nor U17425 (N_17425,N_16950,N_16640);
nand U17426 (N_17426,N_16482,N_16018);
nor U17427 (N_17427,N_16132,N_16007);
nand U17428 (N_17428,N_16367,N_16588);
xnor U17429 (N_17429,N_16701,N_16499);
or U17430 (N_17430,N_16153,N_16889);
or U17431 (N_17431,N_16711,N_16085);
xor U17432 (N_17432,N_16435,N_16509);
nand U17433 (N_17433,N_16472,N_16240);
or U17434 (N_17434,N_16907,N_16063);
or U17435 (N_17435,N_16854,N_16776);
xnor U17436 (N_17436,N_16136,N_16464);
nand U17437 (N_17437,N_16550,N_16067);
or U17438 (N_17438,N_16705,N_16375);
nand U17439 (N_17439,N_16966,N_16780);
or U17440 (N_17440,N_16570,N_16607);
nor U17441 (N_17441,N_16318,N_16451);
xor U17442 (N_17442,N_16561,N_16657);
and U17443 (N_17443,N_16474,N_16905);
xnor U17444 (N_17444,N_16871,N_16325);
nand U17445 (N_17445,N_16461,N_16665);
nor U17446 (N_17446,N_16114,N_16790);
nand U17447 (N_17447,N_16196,N_16695);
or U17448 (N_17448,N_16994,N_16368);
or U17449 (N_17449,N_16094,N_16544);
xor U17450 (N_17450,N_16802,N_16735);
or U17451 (N_17451,N_16670,N_16666);
and U17452 (N_17452,N_16176,N_16742);
and U17453 (N_17453,N_16166,N_16704);
xnor U17454 (N_17454,N_16399,N_16813);
xor U17455 (N_17455,N_16600,N_16434);
xnor U17456 (N_17456,N_16975,N_16327);
and U17457 (N_17457,N_16075,N_16126);
or U17458 (N_17458,N_16626,N_16299);
nand U17459 (N_17459,N_16349,N_16610);
and U17460 (N_17460,N_16216,N_16352);
and U17461 (N_17461,N_16646,N_16234);
or U17462 (N_17462,N_16080,N_16613);
or U17463 (N_17463,N_16000,N_16430);
nor U17464 (N_17464,N_16787,N_16167);
or U17465 (N_17465,N_16519,N_16669);
xnor U17466 (N_17466,N_16619,N_16262);
xor U17467 (N_17467,N_16682,N_16229);
and U17468 (N_17468,N_16336,N_16784);
xor U17469 (N_17469,N_16433,N_16224);
nor U17470 (N_17470,N_16222,N_16443);
nor U17471 (N_17471,N_16140,N_16929);
or U17472 (N_17472,N_16924,N_16488);
xnor U17473 (N_17473,N_16967,N_16883);
xor U17474 (N_17474,N_16353,N_16882);
xnor U17475 (N_17475,N_16620,N_16158);
or U17476 (N_17476,N_16818,N_16664);
or U17477 (N_17477,N_16305,N_16483);
xor U17478 (N_17478,N_16731,N_16432);
xnor U17479 (N_17479,N_16795,N_16841);
and U17480 (N_17480,N_16996,N_16146);
nand U17481 (N_17481,N_16454,N_16885);
xor U17482 (N_17482,N_16330,N_16989);
xor U17483 (N_17483,N_16072,N_16531);
or U17484 (N_17484,N_16992,N_16022);
nand U17485 (N_17485,N_16247,N_16288);
and U17486 (N_17486,N_16015,N_16412);
xnor U17487 (N_17487,N_16320,N_16089);
xnor U17488 (N_17488,N_16822,N_16272);
or U17489 (N_17489,N_16951,N_16839);
nor U17490 (N_17490,N_16477,N_16574);
or U17491 (N_17491,N_16567,N_16857);
and U17492 (N_17492,N_16745,N_16716);
nor U17493 (N_17493,N_16910,N_16411);
nand U17494 (N_17494,N_16512,N_16744);
and U17495 (N_17495,N_16373,N_16410);
and U17496 (N_17496,N_16175,N_16148);
and U17497 (N_17497,N_16725,N_16271);
or U17498 (N_17498,N_16121,N_16296);
xor U17499 (N_17499,N_16971,N_16371);
or U17500 (N_17500,N_16565,N_16320);
xor U17501 (N_17501,N_16667,N_16915);
nand U17502 (N_17502,N_16300,N_16959);
xor U17503 (N_17503,N_16662,N_16174);
or U17504 (N_17504,N_16840,N_16334);
nor U17505 (N_17505,N_16816,N_16499);
nor U17506 (N_17506,N_16687,N_16630);
nand U17507 (N_17507,N_16878,N_16617);
or U17508 (N_17508,N_16693,N_16891);
xor U17509 (N_17509,N_16316,N_16105);
nand U17510 (N_17510,N_16493,N_16698);
xnor U17511 (N_17511,N_16740,N_16193);
or U17512 (N_17512,N_16772,N_16001);
nand U17513 (N_17513,N_16159,N_16936);
nand U17514 (N_17514,N_16127,N_16751);
and U17515 (N_17515,N_16148,N_16606);
and U17516 (N_17516,N_16593,N_16777);
or U17517 (N_17517,N_16953,N_16023);
nor U17518 (N_17518,N_16031,N_16295);
and U17519 (N_17519,N_16792,N_16568);
nor U17520 (N_17520,N_16632,N_16517);
nor U17521 (N_17521,N_16958,N_16035);
nor U17522 (N_17522,N_16875,N_16245);
nor U17523 (N_17523,N_16771,N_16074);
nor U17524 (N_17524,N_16144,N_16048);
xor U17525 (N_17525,N_16326,N_16190);
nor U17526 (N_17526,N_16961,N_16136);
or U17527 (N_17527,N_16227,N_16595);
xnor U17528 (N_17528,N_16464,N_16565);
nor U17529 (N_17529,N_16581,N_16490);
xnor U17530 (N_17530,N_16196,N_16435);
or U17531 (N_17531,N_16131,N_16779);
nor U17532 (N_17532,N_16527,N_16708);
or U17533 (N_17533,N_16407,N_16111);
nor U17534 (N_17534,N_16599,N_16402);
or U17535 (N_17535,N_16317,N_16452);
and U17536 (N_17536,N_16778,N_16532);
or U17537 (N_17537,N_16386,N_16206);
and U17538 (N_17538,N_16786,N_16975);
nor U17539 (N_17539,N_16913,N_16406);
nand U17540 (N_17540,N_16215,N_16930);
and U17541 (N_17541,N_16998,N_16841);
nor U17542 (N_17542,N_16573,N_16744);
or U17543 (N_17543,N_16835,N_16139);
or U17544 (N_17544,N_16644,N_16520);
xor U17545 (N_17545,N_16858,N_16395);
xor U17546 (N_17546,N_16012,N_16495);
nand U17547 (N_17547,N_16311,N_16392);
and U17548 (N_17548,N_16006,N_16654);
xor U17549 (N_17549,N_16169,N_16305);
nor U17550 (N_17550,N_16434,N_16048);
or U17551 (N_17551,N_16367,N_16974);
and U17552 (N_17552,N_16500,N_16496);
nand U17553 (N_17553,N_16411,N_16668);
xor U17554 (N_17554,N_16689,N_16716);
or U17555 (N_17555,N_16481,N_16829);
and U17556 (N_17556,N_16768,N_16039);
and U17557 (N_17557,N_16464,N_16708);
and U17558 (N_17558,N_16124,N_16193);
xor U17559 (N_17559,N_16563,N_16631);
nor U17560 (N_17560,N_16476,N_16018);
nor U17561 (N_17561,N_16731,N_16733);
and U17562 (N_17562,N_16289,N_16385);
and U17563 (N_17563,N_16079,N_16825);
or U17564 (N_17564,N_16846,N_16708);
nor U17565 (N_17565,N_16297,N_16249);
and U17566 (N_17566,N_16695,N_16546);
xnor U17567 (N_17567,N_16054,N_16786);
nor U17568 (N_17568,N_16706,N_16379);
nor U17569 (N_17569,N_16153,N_16569);
and U17570 (N_17570,N_16916,N_16442);
or U17571 (N_17571,N_16141,N_16124);
or U17572 (N_17572,N_16155,N_16969);
xnor U17573 (N_17573,N_16995,N_16880);
or U17574 (N_17574,N_16140,N_16902);
xnor U17575 (N_17575,N_16283,N_16030);
nand U17576 (N_17576,N_16324,N_16212);
or U17577 (N_17577,N_16540,N_16890);
or U17578 (N_17578,N_16349,N_16034);
xnor U17579 (N_17579,N_16166,N_16106);
nor U17580 (N_17580,N_16892,N_16165);
nand U17581 (N_17581,N_16416,N_16014);
nand U17582 (N_17582,N_16295,N_16183);
nor U17583 (N_17583,N_16317,N_16290);
or U17584 (N_17584,N_16420,N_16706);
or U17585 (N_17585,N_16196,N_16521);
xor U17586 (N_17586,N_16552,N_16596);
and U17587 (N_17587,N_16557,N_16941);
or U17588 (N_17588,N_16405,N_16455);
nand U17589 (N_17589,N_16476,N_16946);
and U17590 (N_17590,N_16427,N_16952);
nor U17591 (N_17591,N_16156,N_16742);
and U17592 (N_17592,N_16682,N_16771);
and U17593 (N_17593,N_16732,N_16052);
or U17594 (N_17594,N_16371,N_16413);
nor U17595 (N_17595,N_16376,N_16397);
or U17596 (N_17596,N_16767,N_16943);
xor U17597 (N_17597,N_16409,N_16236);
and U17598 (N_17598,N_16168,N_16918);
or U17599 (N_17599,N_16842,N_16711);
nor U17600 (N_17600,N_16291,N_16089);
nand U17601 (N_17601,N_16401,N_16993);
nor U17602 (N_17602,N_16926,N_16376);
nor U17603 (N_17603,N_16059,N_16021);
or U17604 (N_17604,N_16114,N_16058);
nand U17605 (N_17605,N_16102,N_16504);
or U17606 (N_17606,N_16067,N_16486);
xnor U17607 (N_17607,N_16581,N_16744);
nand U17608 (N_17608,N_16796,N_16301);
nor U17609 (N_17609,N_16234,N_16042);
or U17610 (N_17610,N_16158,N_16154);
nor U17611 (N_17611,N_16325,N_16313);
and U17612 (N_17612,N_16524,N_16041);
xor U17613 (N_17613,N_16069,N_16395);
xor U17614 (N_17614,N_16504,N_16489);
nand U17615 (N_17615,N_16189,N_16888);
nand U17616 (N_17616,N_16607,N_16748);
and U17617 (N_17617,N_16042,N_16045);
nand U17618 (N_17618,N_16234,N_16640);
or U17619 (N_17619,N_16861,N_16984);
nand U17620 (N_17620,N_16234,N_16418);
xnor U17621 (N_17621,N_16653,N_16470);
nand U17622 (N_17622,N_16884,N_16891);
or U17623 (N_17623,N_16958,N_16692);
and U17624 (N_17624,N_16753,N_16108);
and U17625 (N_17625,N_16987,N_16905);
nand U17626 (N_17626,N_16924,N_16032);
xor U17627 (N_17627,N_16207,N_16267);
nand U17628 (N_17628,N_16919,N_16088);
nor U17629 (N_17629,N_16573,N_16021);
xnor U17630 (N_17630,N_16377,N_16503);
xnor U17631 (N_17631,N_16343,N_16892);
or U17632 (N_17632,N_16357,N_16393);
nand U17633 (N_17633,N_16046,N_16758);
nand U17634 (N_17634,N_16836,N_16222);
nand U17635 (N_17635,N_16487,N_16896);
nand U17636 (N_17636,N_16021,N_16614);
and U17637 (N_17637,N_16495,N_16222);
or U17638 (N_17638,N_16132,N_16920);
nor U17639 (N_17639,N_16536,N_16197);
nand U17640 (N_17640,N_16887,N_16354);
xor U17641 (N_17641,N_16987,N_16488);
xor U17642 (N_17642,N_16324,N_16124);
or U17643 (N_17643,N_16064,N_16295);
xnor U17644 (N_17644,N_16402,N_16949);
nand U17645 (N_17645,N_16197,N_16675);
nand U17646 (N_17646,N_16287,N_16120);
nor U17647 (N_17647,N_16993,N_16642);
nand U17648 (N_17648,N_16799,N_16427);
nand U17649 (N_17649,N_16449,N_16586);
and U17650 (N_17650,N_16939,N_16350);
nand U17651 (N_17651,N_16014,N_16348);
xor U17652 (N_17652,N_16965,N_16216);
or U17653 (N_17653,N_16243,N_16619);
nand U17654 (N_17654,N_16223,N_16815);
or U17655 (N_17655,N_16665,N_16653);
and U17656 (N_17656,N_16072,N_16489);
or U17657 (N_17657,N_16199,N_16195);
and U17658 (N_17658,N_16911,N_16719);
nand U17659 (N_17659,N_16064,N_16788);
xnor U17660 (N_17660,N_16244,N_16227);
nand U17661 (N_17661,N_16307,N_16062);
and U17662 (N_17662,N_16970,N_16488);
or U17663 (N_17663,N_16764,N_16080);
nor U17664 (N_17664,N_16031,N_16496);
and U17665 (N_17665,N_16319,N_16536);
nor U17666 (N_17666,N_16196,N_16244);
xnor U17667 (N_17667,N_16270,N_16794);
or U17668 (N_17668,N_16084,N_16206);
nor U17669 (N_17669,N_16539,N_16500);
xnor U17670 (N_17670,N_16656,N_16848);
nand U17671 (N_17671,N_16856,N_16227);
and U17672 (N_17672,N_16643,N_16261);
nand U17673 (N_17673,N_16465,N_16198);
nor U17674 (N_17674,N_16698,N_16935);
or U17675 (N_17675,N_16871,N_16417);
nor U17676 (N_17676,N_16047,N_16783);
and U17677 (N_17677,N_16331,N_16979);
or U17678 (N_17678,N_16224,N_16758);
nand U17679 (N_17679,N_16974,N_16622);
xnor U17680 (N_17680,N_16198,N_16972);
nor U17681 (N_17681,N_16674,N_16593);
and U17682 (N_17682,N_16076,N_16237);
xnor U17683 (N_17683,N_16417,N_16300);
and U17684 (N_17684,N_16570,N_16714);
or U17685 (N_17685,N_16361,N_16478);
and U17686 (N_17686,N_16797,N_16669);
or U17687 (N_17687,N_16348,N_16604);
and U17688 (N_17688,N_16302,N_16067);
xnor U17689 (N_17689,N_16748,N_16402);
and U17690 (N_17690,N_16074,N_16082);
xnor U17691 (N_17691,N_16847,N_16679);
or U17692 (N_17692,N_16542,N_16411);
or U17693 (N_17693,N_16719,N_16695);
nor U17694 (N_17694,N_16603,N_16564);
or U17695 (N_17695,N_16316,N_16332);
xor U17696 (N_17696,N_16977,N_16791);
or U17697 (N_17697,N_16290,N_16643);
or U17698 (N_17698,N_16327,N_16349);
nor U17699 (N_17699,N_16985,N_16382);
xnor U17700 (N_17700,N_16911,N_16732);
nand U17701 (N_17701,N_16798,N_16535);
or U17702 (N_17702,N_16392,N_16877);
or U17703 (N_17703,N_16005,N_16080);
and U17704 (N_17704,N_16473,N_16111);
and U17705 (N_17705,N_16445,N_16661);
or U17706 (N_17706,N_16938,N_16266);
nand U17707 (N_17707,N_16150,N_16160);
and U17708 (N_17708,N_16300,N_16480);
nor U17709 (N_17709,N_16852,N_16917);
nand U17710 (N_17710,N_16996,N_16939);
nor U17711 (N_17711,N_16315,N_16904);
xnor U17712 (N_17712,N_16926,N_16626);
nor U17713 (N_17713,N_16455,N_16318);
or U17714 (N_17714,N_16381,N_16969);
nor U17715 (N_17715,N_16742,N_16907);
nand U17716 (N_17716,N_16557,N_16130);
nor U17717 (N_17717,N_16165,N_16548);
nor U17718 (N_17718,N_16822,N_16586);
xor U17719 (N_17719,N_16966,N_16898);
nand U17720 (N_17720,N_16285,N_16170);
xor U17721 (N_17721,N_16954,N_16305);
nand U17722 (N_17722,N_16020,N_16089);
nor U17723 (N_17723,N_16397,N_16014);
nand U17724 (N_17724,N_16607,N_16274);
or U17725 (N_17725,N_16643,N_16723);
xor U17726 (N_17726,N_16384,N_16506);
or U17727 (N_17727,N_16947,N_16511);
xnor U17728 (N_17728,N_16821,N_16379);
nor U17729 (N_17729,N_16832,N_16490);
xnor U17730 (N_17730,N_16723,N_16504);
nand U17731 (N_17731,N_16888,N_16327);
nand U17732 (N_17732,N_16428,N_16653);
nor U17733 (N_17733,N_16021,N_16134);
nor U17734 (N_17734,N_16606,N_16351);
nor U17735 (N_17735,N_16648,N_16814);
xor U17736 (N_17736,N_16020,N_16176);
nand U17737 (N_17737,N_16279,N_16202);
nor U17738 (N_17738,N_16889,N_16979);
xnor U17739 (N_17739,N_16972,N_16213);
xnor U17740 (N_17740,N_16759,N_16745);
nand U17741 (N_17741,N_16881,N_16773);
and U17742 (N_17742,N_16785,N_16615);
nor U17743 (N_17743,N_16141,N_16611);
nor U17744 (N_17744,N_16597,N_16668);
and U17745 (N_17745,N_16269,N_16996);
nand U17746 (N_17746,N_16607,N_16608);
nand U17747 (N_17747,N_16644,N_16534);
xor U17748 (N_17748,N_16035,N_16711);
and U17749 (N_17749,N_16319,N_16056);
xnor U17750 (N_17750,N_16362,N_16353);
nor U17751 (N_17751,N_16069,N_16316);
nand U17752 (N_17752,N_16750,N_16410);
nor U17753 (N_17753,N_16408,N_16225);
and U17754 (N_17754,N_16117,N_16450);
or U17755 (N_17755,N_16978,N_16476);
nor U17756 (N_17756,N_16414,N_16879);
and U17757 (N_17757,N_16129,N_16109);
nand U17758 (N_17758,N_16174,N_16262);
nor U17759 (N_17759,N_16608,N_16263);
nor U17760 (N_17760,N_16551,N_16444);
and U17761 (N_17761,N_16913,N_16453);
nand U17762 (N_17762,N_16275,N_16816);
or U17763 (N_17763,N_16170,N_16961);
xor U17764 (N_17764,N_16342,N_16415);
and U17765 (N_17765,N_16809,N_16572);
or U17766 (N_17766,N_16788,N_16458);
nand U17767 (N_17767,N_16287,N_16841);
nor U17768 (N_17768,N_16763,N_16786);
or U17769 (N_17769,N_16403,N_16780);
xnor U17770 (N_17770,N_16425,N_16557);
and U17771 (N_17771,N_16015,N_16558);
nor U17772 (N_17772,N_16683,N_16056);
xnor U17773 (N_17773,N_16113,N_16862);
nor U17774 (N_17774,N_16020,N_16521);
and U17775 (N_17775,N_16083,N_16366);
or U17776 (N_17776,N_16605,N_16493);
xor U17777 (N_17777,N_16260,N_16019);
nor U17778 (N_17778,N_16678,N_16808);
or U17779 (N_17779,N_16772,N_16620);
nor U17780 (N_17780,N_16444,N_16035);
xor U17781 (N_17781,N_16974,N_16535);
nand U17782 (N_17782,N_16632,N_16314);
nor U17783 (N_17783,N_16637,N_16082);
nand U17784 (N_17784,N_16360,N_16111);
nor U17785 (N_17785,N_16622,N_16985);
nor U17786 (N_17786,N_16535,N_16048);
or U17787 (N_17787,N_16148,N_16008);
xnor U17788 (N_17788,N_16214,N_16550);
or U17789 (N_17789,N_16189,N_16879);
xnor U17790 (N_17790,N_16410,N_16604);
or U17791 (N_17791,N_16447,N_16933);
and U17792 (N_17792,N_16157,N_16448);
nor U17793 (N_17793,N_16584,N_16824);
nor U17794 (N_17794,N_16874,N_16565);
or U17795 (N_17795,N_16261,N_16802);
and U17796 (N_17796,N_16694,N_16480);
and U17797 (N_17797,N_16849,N_16211);
nand U17798 (N_17798,N_16572,N_16273);
xor U17799 (N_17799,N_16665,N_16562);
or U17800 (N_17800,N_16015,N_16088);
nor U17801 (N_17801,N_16542,N_16102);
or U17802 (N_17802,N_16035,N_16327);
nor U17803 (N_17803,N_16128,N_16606);
xor U17804 (N_17804,N_16138,N_16869);
xnor U17805 (N_17805,N_16603,N_16050);
xor U17806 (N_17806,N_16127,N_16117);
or U17807 (N_17807,N_16992,N_16967);
and U17808 (N_17808,N_16185,N_16431);
and U17809 (N_17809,N_16180,N_16939);
nor U17810 (N_17810,N_16577,N_16497);
nand U17811 (N_17811,N_16074,N_16639);
and U17812 (N_17812,N_16405,N_16878);
and U17813 (N_17813,N_16823,N_16112);
nor U17814 (N_17814,N_16313,N_16586);
nand U17815 (N_17815,N_16791,N_16420);
or U17816 (N_17816,N_16037,N_16451);
and U17817 (N_17817,N_16481,N_16061);
nor U17818 (N_17818,N_16237,N_16319);
nor U17819 (N_17819,N_16828,N_16604);
or U17820 (N_17820,N_16055,N_16321);
nor U17821 (N_17821,N_16415,N_16000);
or U17822 (N_17822,N_16795,N_16279);
nor U17823 (N_17823,N_16549,N_16726);
nor U17824 (N_17824,N_16664,N_16355);
xor U17825 (N_17825,N_16368,N_16113);
xnor U17826 (N_17826,N_16356,N_16937);
nor U17827 (N_17827,N_16887,N_16014);
and U17828 (N_17828,N_16250,N_16006);
xor U17829 (N_17829,N_16737,N_16719);
and U17830 (N_17830,N_16712,N_16253);
or U17831 (N_17831,N_16462,N_16107);
nand U17832 (N_17832,N_16147,N_16656);
nand U17833 (N_17833,N_16165,N_16875);
and U17834 (N_17834,N_16167,N_16444);
xor U17835 (N_17835,N_16635,N_16725);
nor U17836 (N_17836,N_16098,N_16027);
nor U17837 (N_17837,N_16701,N_16421);
nor U17838 (N_17838,N_16895,N_16512);
nor U17839 (N_17839,N_16062,N_16416);
or U17840 (N_17840,N_16131,N_16185);
or U17841 (N_17841,N_16782,N_16272);
and U17842 (N_17842,N_16513,N_16830);
xor U17843 (N_17843,N_16605,N_16207);
or U17844 (N_17844,N_16615,N_16193);
nor U17845 (N_17845,N_16838,N_16313);
or U17846 (N_17846,N_16842,N_16950);
nand U17847 (N_17847,N_16537,N_16250);
nand U17848 (N_17848,N_16910,N_16874);
and U17849 (N_17849,N_16276,N_16545);
and U17850 (N_17850,N_16158,N_16716);
or U17851 (N_17851,N_16988,N_16923);
xor U17852 (N_17852,N_16627,N_16580);
nor U17853 (N_17853,N_16272,N_16132);
nand U17854 (N_17854,N_16342,N_16150);
nand U17855 (N_17855,N_16234,N_16160);
and U17856 (N_17856,N_16616,N_16102);
nand U17857 (N_17857,N_16976,N_16924);
and U17858 (N_17858,N_16752,N_16079);
and U17859 (N_17859,N_16053,N_16778);
nand U17860 (N_17860,N_16812,N_16495);
or U17861 (N_17861,N_16382,N_16977);
nand U17862 (N_17862,N_16061,N_16068);
nand U17863 (N_17863,N_16273,N_16276);
and U17864 (N_17864,N_16733,N_16310);
and U17865 (N_17865,N_16391,N_16083);
nor U17866 (N_17866,N_16301,N_16349);
xnor U17867 (N_17867,N_16014,N_16031);
nor U17868 (N_17868,N_16921,N_16641);
nand U17869 (N_17869,N_16437,N_16904);
nand U17870 (N_17870,N_16327,N_16108);
nor U17871 (N_17871,N_16875,N_16541);
xnor U17872 (N_17872,N_16257,N_16323);
or U17873 (N_17873,N_16624,N_16849);
and U17874 (N_17874,N_16010,N_16900);
nand U17875 (N_17875,N_16276,N_16077);
nor U17876 (N_17876,N_16836,N_16602);
nand U17877 (N_17877,N_16330,N_16885);
nand U17878 (N_17878,N_16898,N_16044);
nand U17879 (N_17879,N_16284,N_16716);
and U17880 (N_17880,N_16464,N_16660);
or U17881 (N_17881,N_16595,N_16999);
or U17882 (N_17882,N_16343,N_16108);
and U17883 (N_17883,N_16047,N_16172);
nor U17884 (N_17884,N_16088,N_16614);
or U17885 (N_17885,N_16632,N_16079);
xnor U17886 (N_17886,N_16599,N_16630);
nor U17887 (N_17887,N_16461,N_16649);
nand U17888 (N_17888,N_16065,N_16657);
nor U17889 (N_17889,N_16792,N_16701);
or U17890 (N_17890,N_16259,N_16926);
and U17891 (N_17891,N_16258,N_16874);
xor U17892 (N_17892,N_16646,N_16350);
nand U17893 (N_17893,N_16554,N_16980);
and U17894 (N_17894,N_16263,N_16229);
nand U17895 (N_17895,N_16178,N_16338);
nand U17896 (N_17896,N_16213,N_16403);
nand U17897 (N_17897,N_16499,N_16987);
or U17898 (N_17898,N_16387,N_16804);
xnor U17899 (N_17899,N_16089,N_16408);
or U17900 (N_17900,N_16974,N_16835);
xnor U17901 (N_17901,N_16636,N_16499);
nand U17902 (N_17902,N_16606,N_16459);
or U17903 (N_17903,N_16401,N_16869);
nor U17904 (N_17904,N_16207,N_16050);
nor U17905 (N_17905,N_16984,N_16980);
xnor U17906 (N_17906,N_16256,N_16569);
nor U17907 (N_17907,N_16851,N_16229);
nor U17908 (N_17908,N_16239,N_16683);
nor U17909 (N_17909,N_16570,N_16449);
nand U17910 (N_17910,N_16366,N_16894);
nor U17911 (N_17911,N_16591,N_16212);
nand U17912 (N_17912,N_16249,N_16679);
and U17913 (N_17913,N_16788,N_16129);
nand U17914 (N_17914,N_16764,N_16720);
xnor U17915 (N_17915,N_16603,N_16783);
nor U17916 (N_17916,N_16210,N_16823);
nand U17917 (N_17917,N_16196,N_16507);
and U17918 (N_17918,N_16400,N_16189);
nor U17919 (N_17919,N_16732,N_16245);
xor U17920 (N_17920,N_16000,N_16217);
xor U17921 (N_17921,N_16578,N_16481);
or U17922 (N_17922,N_16381,N_16960);
and U17923 (N_17923,N_16924,N_16391);
and U17924 (N_17924,N_16931,N_16137);
and U17925 (N_17925,N_16163,N_16226);
nor U17926 (N_17926,N_16137,N_16446);
and U17927 (N_17927,N_16909,N_16580);
nor U17928 (N_17928,N_16000,N_16581);
nor U17929 (N_17929,N_16834,N_16133);
and U17930 (N_17930,N_16171,N_16797);
nor U17931 (N_17931,N_16926,N_16035);
or U17932 (N_17932,N_16628,N_16296);
nand U17933 (N_17933,N_16911,N_16307);
or U17934 (N_17934,N_16704,N_16317);
and U17935 (N_17935,N_16704,N_16361);
and U17936 (N_17936,N_16578,N_16681);
and U17937 (N_17937,N_16278,N_16094);
nand U17938 (N_17938,N_16399,N_16403);
and U17939 (N_17939,N_16212,N_16946);
xor U17940 (N_17940,N_16445,N_16030);
or U17941 (N_17941,N_16911,N_16779);
xor U17942 (N_17942,N_16174,N_16800);
xor U17943 (N_17943,N_16442,N_16219);
nor U17944 (N_17944,N_16289,N_16973);
or U17945 (N_17945,N_16997,N_16720);
nand U17946 (N_17946,N_16564,N_16883);
or U17947 (N_17947,N_16742,N_16984);
nand U17948 (N_17948,N_16929,N_16004);
nand U17949 (N_17949,N_16138,N_16457);
nor U17950 (N_17950,N_16357,N_16882);
or U17951 (N_17951,N_16355,N_16964);
nor U17952 (N_17952,N_16190,N_16811);
or U17953 (N_17953,N_16086,N_16525);
nand U17954 (N_17954,N_16785,N_16123);
nand U17955 (N_17955,N_16883,N_16877);
nor U17956 (N_17956,N_16893,N_16630);
or U17957 (N_17957,N_16042,N_16547);
xnor U17958 (N_17958,N_16439,N_16382);
nand U17959 (N_17959,N_16189,N_16309);
or U17960 (N_17960,N_16516,N_16288);
nand U17961 (N_17961,N_16206,N_16495);
nor U17962 (N_17962,N_16531,N_16563);
and U17963 (N_17963,N_16904,N_16898);
nand U17964 (N_17964,N_16657,N_16722);
nand U17965 (N_17965,N_16119,N_16873);
and U17966 (N_17966,N_16923,N_16837);
nand U17967 (N_17967,N_16570,N_16527);
xor U17968 (N_17968,N_16576,N_16508);
xor U17969 (N_17969,N_16607,N_16800);
and U17970 (N_17970,N_16318,N_16489);
and U17971 (N_17971,N_16158,N_16204);
or U17972 (N_17972,N_16126,N_16494);
or U17973 (N_17973,N_16542,N_16858);
xnor U17974 (N_17974,N_16634,N_16338);
xor U17975 (N_17975,N_16273,N_16134);
nand U17976 (N_17976,N_16705,N_16385);
or U17977 (N_17977,N_16386,N_16687);
nand U17978 (N_17978,N_16905,N_16569);
nand U17979 (N_17979,N_16075,N_16722);
nand U17980 (N_17980,N_16977,N_16240);
nand U17981 (N_17981,N_16213,N_16552);
nand U17982 (N_17982,N_16890,N_16739);
xnor U17983 (N_17983,N_16335,N_16089);
xor U17984 (N_17984,N_16757,N_16727);
nor U17985 (N_17985,N_16182,N_16456);
and U17986 (N_17986,N_16157,N_16720);
and U17987 (N_17987,N_16859,N_16097);
nand U17988 (N_17988,N_16519,N_16366);
nand U17989 (N_17989,N_16760,N_16179);
nor U17990 (N_17990,N_16148,N_16291);
nand U17991 (N_17991,N_16976,N_16566);
or U17992 (N_17992,N_16035,N_16406);
nand U17993 (N_17993,N_16259,N_16301);
xor U17994 (N_17994,N_16796,N_16658);
xnor U17995 (N_17995,N_16550,N_16643);
and U17996 (N_17996,N_16209,N_16865);
nand U17997 (N_17997,N_16806,N_16922);
nand U17998 (N_17998,N_16308,N_16654);
nor U17999 (N_17999,N_16769,N_16358);
nand U18000 (N_18000,N_17400,N_17917);
nor U18001 (N_18001,N_17087,N_17742);
xor U18002 (N_18002,N_17422,N_17827);
xor U18003 (N_18003,N_17125,N_17820);
and U18004 (N_18004,N_17541,N_17090);
or U18005 (N_18005,N_17990,N_17774);
nand U18006 (N_18006,N_17977,N_17175);
xnor U18007 (N_18007,N_17950,N_17245);
nor U18008 (N_18008,N_17203,N_17532);
or U18009 (N_18009,N_17595,N_17849);
xor U18010 (N_18010,N_17451,N_17503);
xor U18011 (N_18011,N_17062,N_17094);
or U18012 (N_18012,N_17581,N_17225);
or U18013 (N_18013,N_17878,N_17993);
and U18014 (N_18014,N_17475,N_17297);
or U18015 (N_18015,N_17756,N_17624);
nor U18016 (N_18016,N_17221,N_17907);
and U18017 (N_18017,N_17835,N_17766);
and U18018 (N_18018,N_17998,N_17363);
xnor U18019 (N_18019,N_17416,N_17891);
or U18020 (N_18020,N_17874,N_17757);
xnor U18021 (N_18021,N_17957,N_17608);
xnor U18022 (N_18022,N_17722,N_17591);
nand U18023 (N_18023,N_17800,N_17684);
nor U18024 (N_18024,N_17191,N_17255);
and U18025 (N_18025,N_17882,N_17197);
and U18026 (N_18026,N_17702,N_17302);
and U18027 (N_18027,N_17754,N_17413);
nor U18028 (N_18028,N_17312,N_17710);
xnor U18029 (N_18029,N_17174,N_17831);
nor U18030 (N_18030,N_17238,N_17387);
and U18031 (N_18031,N_17158,N_17498);
xor U18032 (N_18032,N_17968,N_17740);
nor U18033 (N_18033,N_17785,N_17965);
xnor U18034 (N_18034,N_17036,N_17649);
nor U18035 (N_18035,N_17456,N_17585);
xor U18036 (N_18036,N_17060,N_17949);
nor U18037 (N_18037,N_17889,N_17574);
nand U18038 (N_18038,N_17868,N_17667);
and U18039 (N_18039,N_17788,N_17084);
nor U18040 (N_18040,N_17846,N_17228);
nor U18041 (N_18041,N_17226,N_17739);
nand U18042 (N_18042,N_17025,N_17274);
and U18043 (N_18043,N_17049,N_17142);
nand U18044 (N_18044,N_17336,N_17983);
and U18045 (N_18045,N_17510,N_17506);
and U18046 (N_18046,N_17706,N_17507);
nand U18047 (N_18047,N_17712,N_17470);
nand U18048 (N_18048,N_17743,N_17252);
or U18049 (N_18049,N_17737,N_17765);
or U18050 (N_18050,N_17641,N_17926);
xor U18051 (N_18051,N_17958,N_17732);
and U18052 (N_18052,N_17531,N_17139);
and U18053 (N_18053,N_17313,N_17651);
and U18054 (N_18054,N_17693,N_17857);
or U18055 (N_18055,N_17211,N_17935);
xnor U18056 (N_18056,N_17529,N_17279);
nand U18057 (N_18057,N_17376,N_17077);
and U18058 (N_18058,N_17303,N_17954);
and U18059 (N_18059,N_17332,N_17471);
nand U18060 (N_18060,N_17603,N_17898);
xor U18061 (N_18061,N_17844,N_17461);
and U18062 (N_18062,N_17130,N_17107);
and U18063 (N_18063,N_17559,N_17607);
nand U18064 (N_18064,N_17352,N_17789);
nor U18065 (N_18065,N_17096,N_17170);
and U18066 (N_18066,N_17964,N_17720);
or U18067 (N_18067,N_17782,N_17168);
nand U18068 (N_18068,N_17398,N_17896);
nand U18069 (N_18069,N_17551,N_17767);
nor U18070 (N_18070,N_17029,N_17584);
nor U18071 (N_18071,N_17658,N_17277);
or U18072 (N_18072,N_17802,N_17877);
nand U18073 (N_18073,N_17679,N_17455);
nand U18074 (N_18074,N_17910,N_17420);
and U18075 (N_18075,N_17458,N_17561);
xor U18076 (N_18076,N_17527,N_17848);
xnor U18077 (N_18077,N_17414,N_17148);
and U18078 (N_18078,N_17076,N_17617);
nor U18079 (N_18079,N_17521,N_17051);
nor U18080 (N_18080,N_17564,N_17755);
nand U18081 (N_18081,N_17150,N_17524);
nor U18082 (N_18082,N_17114,N_17216);
or U18083 (N_18083,N_17675,N_17281);
nand U18084 (N_18084,N_17932,N_17407);
xor U18085 (N_18085,N_17481,N_17262);
nand U18086 (N_18086,N_17640,N_17146);
or U18087 (N_18087,N_17880,N_17365);
or U18088 (N_18088,N_17929,N_17229);
or U18089 (N_18089,N_17061,N_17704);
xnor U18090 (N_18090,N_17236,N_17103);
nor U18091 (N_18091,N_17473,N_17560);
and U18092 (N_18092,N_17945,N_17396);
or U18093 (N_18093,N_17768,N_17557);
xnor U18094 (N_18094,N_17567,N_17695);
xor U18095 (N_18095,N_17786,N_17444);
xnor U18096 (N_18096,N_17052,N_17549);
nor U18097 (N_18097,N_17237,N_17545);
nor U18098 (N_18098,N_17323,N_17123);
nand U18099 (N_18099,N_17952,N_17673);
and U18100 (N_18100,N_17497,N_17402);
nand U18101 (N_18101,N_17777,N_17469);
xor U18102 (N_18102,N_17227,N_17292);
or U18103 (N_18103,N_17450,N_17568);
xnor U18104 (N_18104,N_17944,N_17657);
and U18105 (N_18105,N_17514,N_17477);
nand U18106 (N_18106,N_17465,N_17169);
nor U18107 (N_18107,N_17818,N_17707);
nor U18108 (N_18108,N_17258,N_17589);
and U18109 (N_18109,N_17593,N_17594);
nand U18110 (N_18110,N_17565,N_17794);
nor U18111 (N_18111,N_17875,N_17254);
xnor U18112 (N_18112,N_17747,N_17791);
and U18113 (N_18113,N_17689,N_17394);
xor U18114 (N_18114,N_17586,N_17535);
nand U18115 (N_18115,N_17733,N_17718);
and U18116 (N_18116,N_17962,N_17612);
and U18117 (N_18117,N_17727,N_17375);
and U18118 (N_18118,N_17263,N_17135);
or U18119 (N_18119,N_17068,N_17324);
and U18120 (N_18120,N_17256,N_17752);
nand U18121 (N_18121,N_17670,N_17663);
and U18122 (N_18122,N_17769,N_17172);
or U18123 (N_18123,N_17770,N_17329);
nand U18124 (N_18124,N_17643,N_17030);
and U18125 (N_18125,N_17692,N_17038);
xor U18126 (N_18126,N_17098,N_17655);
or U18127 (N_18127,N_17984,N_17486);
nor U18128 (N_18128,N_17569,N_17536);
xor U18129 (N_18129,N_17224,N_17017);
and U18130 (N_18130,N_17871,N_17086);
nand U18131 (N_18131,N_17071,N_17018);
xor U18132 (N_18132,N_17092,N_17424);
nor U18133 (N_18133,N_17326,N_17286);
or U18134 (N_18134,N_17632,N_17423);
xor U18135 (N_18135,N_17033,N_17709);
xor U18136 (N_18136,N_17816,N_17714);
or U18137 (N_18137,N_17374,N_17719);
nand U18138 (N_18138,N_17153,N_17276);
or U18139 (N_18139,N_17668,N_17886);
xor U18140 (N_18140,N_17070,N_17004);
xnor U18141 (N_18141,N_17577,N_17043);
or U18142 (N_18142,N_17867,N_17128);
nand U18143 (N_18143,N_17322,N_17911);
xor U18144 (N_18144,N_17852,N_17717);
or U18145 (N_18145,N_17853,N_17730);
nor U18146 (N_18146,N_17748,N_17308);
or U18147 (N_18147,N_17937,N_17337);
nand U18148 (N_18148,N_17399,N_17253);
nand U18149 (N_18149,N_17079,N_17404);
or U18150 (N_18150,N_17526,N_17434);
xor U18151 (N_18151,N_17384,N_17235);
nor U18152 (N_18152,N_17575,N_17966);
or U18153 (N_18153,N_17476,N_17055);
nand U18154 (N_18154,N_17464,N_17354);
nand U18155 (N_18155,N_17140,N_17341);
xnor U18156 (N_18156,N_17278,N_17190);
xnor U18157 (N_18157,N_17300,N_17188);
nor U18158 (N_18158,N_17397,N_17177);
nand U18159 (N_18159,N_17291,N_17466);
xnor U18160 (N_18160,N_17014,N_17922);
nand U18161 (N_18161,N_17345,N_17751);
nor U18162 (N_18162,N_17904,N_17259);
nand U18163 (N_18163,N_17677,N_17630);
or U18164 (N_18164,N_17895,N_17192);
nor U18165 (N_18165,N_17705,N_17888);
nor U18166 (N_18166,N_17750,N_17010);
or U18167 (N_18167,N_17468,N_17290);
or U18168 (N_18168,N_17563,N_17019);
nand U18169 (N_18169,N_17822,N_17296);
xor U18170 (N_18170,N_17588,N_17582);
nor U18171 (N_18171,N_17570,N_17264);
nor U18172 (N_18172,N_17951,N_17008);
nand U18173 (N_18173,N_17543,N_17115);
or U18174 (N_18174,N_17540,N_17537);
xor U18175 (N_18175,N_17523,N_17261);
xor U18176 (N_18176,N_17606,N_17916);
and U18177 (N_18177,N_17851,N_17515);
xor U18178 (N_18178,N_17894,N_17196);
or U18179 (N_18179,N_17257,N_17696);
or U18180 (N_18180,N_17002,N_17806);
or U18181 (N_18181,N_17362,N_17650);
nand U18182 (N_18182,N_17906,N_17771);
or U18183 (N_18183,N_17267,N_17132);
nor U18184 (N_18184,N_17187,N_17454);
nand U18185 (N_18185,N_17494,N_17654);
nor U18186 (N_18186,N_17311,N_17652);
xor U18187 (N_18187,N_17970,N_17202);
xnor U18188 (N_18188,N_17513,N_17035);
and U18189 (N_18189,N_17863,N_17293);
xnor U18190 (N_18190,N_17378,N_17905);
and U18191 (N_18191,N_17691,N_17830);
and U18192 (N_18192,N_17295,N_17900);
or U18193 (N_18193,N_17645,N_17854);
or U18194 (N_18194,N_17512,N_17441);
or U18195 (N_18195,N_17890,N_17386);
nor U18196 (N_18196,N_17307,N_17351);
nor U18197 (N_18197,N_17230,N_17596);
nand U18198 (N_18198,N_17088,N_17357);
nand U18199 (N_18199,N_17991,N_17484);
xnor U18200 (N_18200,N_17054,N_17104);
or U18201 (N_18201,N_17360,N_17266);
and U18202 (N_18202,N_17305,N_17304);
nor U18203 (N_18203,N_17181,N_17725);
or U18204 (N_18204,N_17735,N_17941);
xnor U18205 (N_18205,N_17686,N_17348);
and U18206 (N_18206,N_17698,N_17260);
nor U18207 (N_18207,N_17270,N_17919);
nand U18208 (N_18208,N_17199,N_17775);
xor U18209 (N_18209,N_17106,N_17249);
nand U18210 (N_18210,N_17412,N_17597);
and U18211 (N_18211,N_17636,N_17463);
nor U18212 (N_18212,N_17271,N_17493);
and U18213 (N_18213,N_17381,N_17328);
nor U18214 (N_18214,N_17823,N_17986);
xor U18215 (N_18215,N_17161,N_17611);
nand U18216 (N_18216,N_17152,N_17738);
xor U18217 (N_18217,N_17845,N_17085);
or U18218 (N_18218,N_17200,N_17600);
nand U18219 (N_18219,N_17244,N_17298);
xor U18220 (N_18220,N_17826,N_17997);
or U18221 (N_18221,N_17467,N_17836);
nor U18222 (N_18222,N_17946,N_17214);
xor U18223 (N_18223,N_17759,N_17343);
xnor U18224 (N_18224,N_17711,N_17566);
and U18225 (N_18225,N_17347,N_17495);
xor U18226 (N_18226,N_17832,N_17073);
nor U18227 (N_18227,N_17981,N_17438);
nand U18228 (N_18228,N_17969,N_17207);
or U18229 (N_18229,N_17417,N_17382);
nor U18230 (N_18230,N_17317,N_17440);
nor U18231 (N_18231,N_17330,N_17814);
or U18232 (N_18232,N_17961,N_17697);
or U18233 (N_18233,N_17869,N_17127);
or U18234 (N_18234,N_17599,N_17516);
or U18235 (N_18235,N_17173,N_17431);
xor U18236 (N_18236,N_17195,N_17027);
xor U18237 (N_18237,N_17368,N_17885);
nor U18238 (N_18238,N_17285,N_17314);
nand U18239 (N_18239,N_17519,N_17518);
and U18240 (N_18240,N_17231,N_17939);
xor U18241 (N_18241,N_17410,N_17306);
nand U18242 (N_18242,N_17508,N_17634);
and U18243 (N_18243,N_17186,N_17687);
nor U18244 (N_18244,N_17948,N_17690);
nand U18245 (N_18245,N_17275,N_17065);
and U18246 (N_18246,N_17700,N_17309);
and U18247 (N_18247,N_17862,N_17884);
nor U18248 (N_18248,N_17058,N_17547);
nor U18249 (N_18249,N_17373,N_17145);
and U18250 (N_18250,N_17979,N_17810);
nor U18251 (N_18251,N_17887,N_17223);
and U18252 (N_18252,N_17205,N_17320);
xnor U18253 (N_18253,N_17544,N_17415);
nor U18254 (N_18254,N_17380,N_17353);
or U18255 (N_18255,N_17683,N_17797);
xnor U18256 (N_18256,N_17390,N_17680);
nand U18257 (N_18257,N_17445,N_17623);
nand U18258 (N_18258,N_17517,N_17856);
or U18259 (N_18259,N_17621,N_17411);
and U18260 (N_18260,N_17914,N_17746);
nand U18261 (N_18261,N_17442,N_17425);
nand U18262 (N_18262,N_17108,N_17405);
xor U18263 (N_18263,N_17217,N_17095);
or U18264 (N_18264,N_17528,N_17478);
and U18265 (N_18265,N_17149,N_17918);
nand U18266 (N_18266,N_17960,N_17601);
nand U18267 (N_18267,N_17778,N_17699);
xor U18268 (N_18268,N_17385,N_17287);
or U18269 (N_18269,N_17427,N_17246);
nor U18270 (N_18270,N_17459,N_17934);
xnor U18271 (N_18271,N_17080,N_17164);
and U18272 (N_18272,N_17426,N_17821);
nand U18273 (N_18273,N_17028,N_17250);
nor U18274 (N_18274,N_17796,N_17901);
and U18275 (N_18275,N_17501,N_17803);
xor U18276 (N_18276,N_17485,N_17143);
xnor U18277 (N_18277,N_17182,N_17633);
nor U18278 (N_18278,N_17403,N_17248);
or U18279 (N_18279,N_17110,N_17940);
and U18280 (N_18280,N_17963,N_17653);
and U18281 (N_18281,N_17239,N_17022);
nand U18282 (N_18282,N_17676,N_17453);
and U18283 (N_18283,N_17121,N_17151);
or U18284 (N_18284,N_17784,N_17005);
nand U18285 (N_18285,N_17439,N_17915);
xor U18286 (N_18286,N_17003,N_17626);
xnor U18287 (N_18287,N_17590,N_17101);
nand U18288 (N_18288,N_17578,N_17489);
and U18289 (N_18289,N_17116,N_17674);
xnor U18290 (N_18290,N_17488,N_17480);
nand U18291 (N_18291,N_17602,N_17193);
and U18292 (N_18292,N_17576,N_17804);
nor U18293 (N_18293,N_17391,N_17452);
nor U18294 (N_18294,N_17120,N_17272);
or U18295 (N_18295,N_17971,N_17171);
and U18296 (N_18296,N_17069,N_17660);
and U18297 (N_18297,N_17001,N_17715);
or U18298 (N_18298,N_17758,N_17613);
or U18299 (N_18299,N_17629,N_17093);
xnor U18300 (N_18300,N_17105,N_17113);
or U18301 (N_18301,N_17909,N_17729);
xor U18302 (N_18302,N_17163,N_17533);
nand U18303 (N_18303,N_17841,N_17437);
nand U18304 (N_18304,N_17542,N_17638);
and U18305 (N_18305,N_17269,N_17622);
nor U18306 (N_18306,N_17923,N_17511);
and U18307 (N_18307,N_17956,N_17795);
xnor U18308 (N_18308,N_17864,N_17344);
nor U18309 (N_18309,N_17339,N_17047);
xor U18310 (N_18310,N_17793,N_17609);
nand U18311 (N_18311,N_17761,N_17358);
nand U18312 (N_18312,N_17598,N_17790);
xnor U18313 (N_18313,N_17472,N_17408);
nand U18314 (N_18314,N_17637,N_17075);
nor U18315 (N_18315,N_17037,N_17162);
nand U18316 (N_18316,N_17897,N_17999);
or U18317 (N_18317,N_17671,N_17974);
and U18318 (N_18318,N_17370,N_17813);
and U18319 (N_18319,N_17111,N_17615);
xnor U18320 (N_18320,N_17947,N_17372);
or U18321 (N_18321,N_17839,N_17801);
xnor U18322 (N_18322,N_17013,N_17708);
and U18323 (N_18323,N_17942,N_17741);
and U18324 (N_18324,N_17504,N_17166);
and U18325 (N_18325,N_17927,N_17861);
nand U18326 (N_18326,N_17490,N_17496);
and U18327 (N_18327,N_17315,N_17011);
nand U18328 (N_18328,N_17843,N_17024);
and U18329 (N_18329,N_17007,N_17350);
xnor U18330 (N_18330,N_17865,N_17432);
xnor U18331 (N_18331,N_17201,N_17222);
nand U18332 (N_18332,N_17118,N_17776);
and U18333 (N_18333,N_17760,N_17573);
xor U18334 (N_18334,N_17204,N_17953);
nor U18335 (N_18335,N_17701,N_17487);
nand U18336 (N_18336,N_17847,N_17097);
nand U18337 (N_18337,N_17367,N_17046);
nor U18338 (N_18338,N_17749,N_17234);
or U18339 (N_18339,N_17185,N_17383);
xor U18340 (N_18340,N_17931,N_17393);
or U18341 (N_18341,N_17479,N_17838);
nand U18342 (N_18342,N_17421,N_17763);
xnor U18343 (N_18343,N_17218,N_17783);
nand U18344 (N_18344,N_17798,N_17483);
and U18345 (N_18345,N_17012,N_17713);
and U18346 (N_18346,N_17183,N_17819);
or U18347 (N_18347,N_17000,N_17294);
and U18348 (N_18348,N_17474,N_17083);
xnor U18349 (N_18349,N_17457,N_17338);
nor U18350 (N_18350,N_17016,N_17842);
xnor U18351 (N_18351,N_17379,N_17091);
xor U18352 (N_18352,N_17418,N_17571);
xor U18353 (N_18353,N_17924,N_17505);
xor U18354 (N_18354,N_17833,N_17067);
nor U18355 (N_18355,N_17764,N_17872);
nand U18356 (N_18356,N_17122,N_17179);
nand U18357 (N_18357,N_17808,N_17447);
xnor U18358 (N_18358,N_17301,N_17936);
and U18359 (N_18359,N_17144,N_17592);
xnor U18360 (N_18360,N_17015,N_17388);
or U18361 (N_18361,N_17053,N_17781);
nand U18362 (N_18362,N_17074,N_17522);
or U18363 (N_18363,N_17265,N_17772);
xor U18364 (N_18364,N_17605,N_17136);
or U18365 (N_18365,N_17141,N_17546);
nor U18366 (N_18366,N_17042,N_17006);
nand U18367 (N_18367,N_17072,N_17066);
or U18368 (N_18368,N_17688,N_17359);
xnor U18369 (N_18369,N_17976,N_17892);
or U18370 (N_18370,N_17219,N_17395);
nor U18371 (N_18371,N_17552,N_17299);
xnor U18372 (N_18372,N_17627,N_17987);
and U18373 (N_18373,N_17041,N_17129);
and U18374 (N_18374,N_17647,N_17155);
nand U18375 (N_18375,N_17614,N_17639);
xor U18376 (N_18376,N_17938,N_17251);
nand U18377 (N_18377,N_17031,N_17855);
or U18378 (N_18378,N_17099,N_17428);
nand U18379 (N_18379,N_17021,N_17828);
or U18380 (N_18380,N_17619,N_17921);
xnor U18381 (N_18381,N_17534,N_17319);
nor U18382 (N_18382,N_17799,N_17694);
nand U18383 (N_18383,N_17762,N_17137);
nand U18384 (N_18384,N_17724,N_17980);
and U18385 (N_18385,N_17059,N_17930);
xor U18386 (N_18386,N_17661,N_17189);
nand U18387 (N_18387,N_17817,N_17208);
and U18388 (N_18388,N_17430,N_17809);
or U18389 (N_18389,N_17824,N_17134);
or U18390 (N_18390,N_17039,N_17126);
or U18391 (N_18391,N_17157,N_17050);
nor U18392 (N_18392,N_17736,N_17321);
nand U18393 (N_18393,N_17045,N_17023);
xor U18394 (N_18394,N_17180,N_17520);
xnor U18395 (N_18395,N_17879,N_17996);
and U18396 (N_18396,N_17233,N_17744);
or U18397 (N_18397,N_17184,N_17943);
nand U18398 (N_18398,N_17669,N_17635);
nand U18399 (N_18399,N_17063,N_17335);
xor U18400 (N_18400,N_17154,N_17903);
nand U18401 (N_18401,N_17355,N_17210);
nor U18402 (N_18402,N_17850,N_17401);
xnor U18403 (N_18403,N_17176,N_17716);
and U18404 (N_18404,N_17665,N_17100);
nand U18405 (N_18405,N_17333,N_17429);
nand U18406 (N_18406,N_17881,N_17815);
or U18407 (N_18407,N_17102,N_17048);
nor U18408 (N_18408,N_17811,N_17558);
xnor U18409 (N_18409,N_17131,N_17194);
xor U18410 (N_18410,N_17572,N_17975);
nand U18411 (N_18411,N_17978,N_17642);
and U18412 (N_18412,N_17579,N_17240);
xnor U18413 (N_18413,N_17371,N_17500);
and U18414 (N_18414,N_17325,N_17556);
or U18415 (N_18415,N_17369,N_17955);
and U18416 (N_18416,N_17913,N_17873);
and U18417 (N_18417,N_17446,N_17745);
and U18418 (N_18418,N_17082,N_17327);
and U18419 (N_18419,N_17726,N_17912);
xnor U18420 (N_18420,N_17268,N_17656);
nand U18421 (N_18421,N_17460,N_17112);
and U18422 (N_18422,N_17057,N_17628);
xor U18423 (N_18423,N_17883,N_17032);
xnor U18424 (N_18424,N_17550,N_17734);
or U18425 (N_18425,N_17812,N_17840);
nor U18426 (N_18426,N_17364,N_17644);
and U18427 (N_18427,N_17056,N_17138);
or U18428 (N_18428,N_17859,N_17773);
xor U18429 (N_18429,N_17982,N_17316);
nand U18430 (N_18430,N_17616,N_17356);
and U18431 (N_18431,N_17377,N_17805);
nand U18432 (N_18432,N_17555,N_17289);
nor U18433 (N_18433,N_17462,N_17449);
nand U18434 (N_18434,N_17985,N_17530);
and U18435 (N_18435,N_17212,N_17109);
and U18436 (N_18436,N_17925,N_17034);
or U18437 (N_18437,N_17241,N_17995);
nand U18438 (N_18438,N_17436,N_17198);
or U18439 (N_18439,N_17992,N_17731);
or U18440 (N_18440,N_17902,N_17928);
and U18441 (N_18441,N_17342,N_17435);
and U18442 (N_18442,N_17448,N_17988);
nor U18443 (N_18443,N_17443,N_17703);
and U18444 (N_18444,N_17213,N_17243);
and U18445 (N_18445,N_17721,N_17009);
xor U18446 (N_18446,N_17829,N_17664);
xnor U18447 (N_18447,N_17648,N_17866);
nand U18448 (N_18448,N_17499,N_17165);
nor U18449 (N_18449,N_17283,N_17780);
or U18450 (N_18450,N_17672,N_17119);
nor U18451 (N_18451,N_17419,N_17392);
nand U18452 (N_18452,N_17124,N_17610);
nand U18453 (N_18453,N_17220,N_17933);
nand U18454 (N_18454,N_17273,N_17681);
nor U18455 (N_18455,N_17792,N_17893);
nand U18456 (N_18456,N_17525,N_17078);
nor U18457 (N_18457,N_17482,N_17349);
nor U18458 (N_18458,N_17618,N_17834);
and U18459 (N_18459,N_17787,N_17020);
nor U18460 (N_18460,N_17334,N_17753);
and U18461 (N_18461,N_17666,N_17646);
and U18462 (N_18462,N_17860,N_17728);
xnor U18463 (N_18463,N_17625,N_17587);
xor U18464 (N_18464,N_17340,N_17361);
or U18465 (N_18465,N_17232,N_17807);
xor U18466 (N_18466,N_17026,N_17409);
or U18467 (N_18467,N_17662,N_17837);
nor U18468 (N_18468,N_17973,N_17994);
nand U18469 (N_18469,N_17583,N_17920);
and U18470 (N_18470,N_17509,N_17247);
and U18471 (N_18471,N_17659,N_17678);
nor U18472 (N_18472,N_17723,N_17282);
and U18473 (N_18473,N_17876,N_17160);
or U18474 (N_18474,N_17159,N_17089);
and U18475 (N_18475,N_17502,N_17331);
or U18476 (N_18476,N_17553,N_17366);
or U18477 (N_18477,N_17280,N_17117);
nand U18478 (N_18478,N_17554,N_17215);
or U18479 (N_18479,N_17081,N_17538);
or U18480 (N_18480,N_17631,N_17310);
and U18481 (N_18481,N_17989,N_17908);
or U18482 (N_18482,N_17147,N_17580);
nor U18483 (N_18483,N_17242,N_17548);
and U18484 (N_18484,N_17620,N_17682);
xnor U18485 (N_18485,N_17967,N_17156);
nand U18486 (N_18486,N_17539,N_17899);
or U18487 (N_18487,N_17491,N_17825);
nand U18488 (N_18488,N_17562,N_17959);
and U18489 (N_18489,N_17406,N_17133);
and U18490 (N_18490,N_17318,N_17433);
nand U18491 (N_18491,N_17064,N_17604);
or U18492 (N_18492,N_17288,N_17209);
xnor U18493 (N_18493,N_17779,N_17167);
or U18494 (N_18494,N_17389,N_17858);
nand U18495 (N_18495,N_17178,N_17206);
nor U18496 (N_18496,N_17972,N_17346);
nor U18497 (N_18497,N_17492,N_17685);
and U18498 (N_18498,N_17040,N_17284);
and U18499 (N_18499,N_17044,N_17870);
or U18500 (N_18500,N_17760,N_17412);
nand U18501 (N_18501,N_17247,N_17646);
xor U18502 (N_18502,N_17616,N_17731);
nor U18503 (N_18503,N_17866,N_17705);
nand U18504 (N_18504,N_17533,N_17460);
nand U18505 (N_18505,N_17633,N_17586);
or U18506 (N_18506,N_17405,N_17391);
nand U18507 (N_18507,N_17215,N_17699);
nor U18508 (N_18508,N_17721,N_17783);
and U18509 (N_18509,N_17006,N_17649);
or U18510 (N_18510,N_17472,N_17311);
nand U18511 (N_18511,N_17226,N_17036);
and U18512 (N_18512,N_17614,N_17917);
xnor U18513 (N_18513,N_17721,N_17218);
nand U18514 (N_18514,N_17331,N_17881);
xnor U18515 (N_18515,N_17268,N_17641);
or U18516 (N_18516,N_17887,N_17383);
xnor U18517 (N_18517,N_17583,N_17783);
or U18518 (N_18518,N_17603,N_17422);
nand U18519 (N_18519,N_17892,N_17875);
nor U18520 (N_18520,N_17806,N_17094);
and U18521 (N_18521,N_17697,N_17246);
nand U18522 (N_18522,N_17737,N_17833);
nor U18523 (N_18523,N_17365,N_17258);
or U18524 (N_18524,N_17551,N_17614);
and U18525 (N_18525,N_17430,N_17031);
or U18526 (N_18526,N_17326,N_17144);
nand U18527 (N_18527,N_17863,N_17990);
xor U18528 (N_18528,N_17303,N_17298);
or U18529 (N_18529,N_17023,N_17352);
and U18530 (N_18530,N_17824,N_17758);
and U18531 (N_18531,N_17340,N_17171);
nor U18532 (N_18532,N_17738,N_17296);
and U18533 (N_18533,N_17194,N_17403);
or U18534 (N_18534,N_17227,N_17912);
and U18535 (N_18535,N_17722,N_17590);
nand U18536 (N_18536,N_17241,N_17346);
nor U18537 (N_18537,N_17488,N_17355);
nor U18538 (N_18538,N_17514,N_17509);
nand U18539 (N_18539,N_17144,N_17866);
nand U18540 (N_18540,N_17372,N_17808);
xor U18541 (N_18541,N_17818,N_17158);
xor U18542 (N_18542,N_17926,N_17637);
nor U18543 (N_18543,N_17912,N_17607);
or U18544 (N_18544,N_17252,N_17861);
and U18545 (N_18545,N_17865,N_17278);
nor U18546 (N_18546,N_17431,N_17749);
and U18547 (N_18547,N_17354,N_17036);
nand U18548 (N_18548,N_17269,N_17185);
nor U18549 (N_18549,N_17609,N_17197);
and U18550 (N_18550,N_17097,N_17413);
and U18551 (N_18551,N_17948,N_17872);
nor U18552 (N_18552,N_17905,N_17170);
xnor U18553 (N_18553,N_17529,N_17420);
or U18554 (N_18554,N_17362,N_17059);
nor U18555 (N_18555,N_17764,N_17715);
nor U18556 (N_18556,N_17265,N_17481);
nor U18557 (N_18557,N_17040,N_17352);
or U18558 (N_18558,N_17839,N_17224);
or U18559 (N_18559,N_17649,N_17421);
xor U18560 (N_18560,N_17726,N_17555);
nand U18561 (N_18561,N_17191,N_17688);
xor U18562 (N_18562,N_17308,N_17840);
xor U18563 (N_18563,N_17518,N_17554);
and U18564 (N_18564,N_17760,N_17063);
and U18565 (N_18565,N_17620,N_17034);
nand U18566 (N_18566,N_17122,N_17106);
xor U18567 (N_18567,N_17973,N_17857);
xor U18568 (N_18568,N_17809,N_17788);
xnor U18569 (N_18569,N_17436,N_17509);
nor U18570 (N_18570,N_17050,N_17012);
or U18571 (N_18571,N_17763,N_17390);
nand U18572 (N_18572,N_17192,N_17873);
xnor U18573 (N_18573,N_17571,N_17406);
nor U18574 (N_18574,N_17742,N_17764);
and U18575 (N_18575,N_17318,N_17801);
xnor U18576 (N_18576,N_17303,N_17138);
nor U18577 (N_18577,N_17242,N_17796);
nor U18578 (N_18578,N_17246,N_17668);
nor U18579 (N_18579,N_17977,N_17882);
or U18580 (N_18580,N_17245,N_17495);
xor U18581 (N_18581,N_17458,N_17767);
nand U18582 (N_18582,N_17009,N_17478);
nor U18583 (N_18583,N_17522,N_17579);
nor U18584 (N_18584,N_17986,N_17185);
xor U18585 (N_18585,N_17532,N_17339);
and U18586 (N_18586,N_17814,N_17671);
and U18587 (N_18587,N_17411,N_17557);
and U18588 (N_18588,N_17088,N_17914);
nor U18589 (N_18589,N_17077,N_17947);
nor U18590 (N_18590,N_17294,N_17141);
nand U18591 (N_18591,N_17686,N_17023);
xor U18592 (N_18592,N_17802,N_17309);
nor U18593 (N_18593,N_17240,N_17891);
nor U18594 (N_18594,N_17498,N_17848);
and U18595 (N_18595,N_17530,N_17702);
or U18596 (N_18596,N_17627,N_17979);
and U18597 (N_18597,N_17167,N_17498);
nor U18598 (N_18598,N_17718,N_17765);
xor U18599 (N_18599,N_17003,N_17319);
xor U18600 (N_18600,N_17182,N_17809);
nand U18601 (N_18601,N_17696,N_17731);
xor U18602 (N_18602,N_17304,N_17756);
xor U18603 (N_18603,N_17300,N_17485);
nor U18604 (N_18604,N_17419,N_17426);
nor U18605 (N_18605,N_17771,N_17941);
or U18606 (N_18606,N_17413,N_17022);
or U18607 (N_18607,N_17955,N_17952);
and U18608 (N_18608,N_17417,N_17275);
or U18609 (N_18609,N_17313,N_17129);
nand U18610 (N_18610,N_17081,N_17643);
or U18611 (N_18611,N_17583,N_17548);
or U18612 (N_18612,N_17715,N_17849);
or U18613 (N_18613,N_17985,N_17804);
nor U18614 (N_18614,N_17244,N_17804);
nor U18615 (N_18615,N_17525,N_17820);
and U18616 (N_18616,N_17115,N_17564);
and U18617 (N_18617,N_17964,N_17656);
xor U18618 (N_18618,N_17080,N_17939);
nand U18619 (N_18619,N_17471,N_17960);
nand U18620 (N_18620,N_17672,N_17236);
xor U18621 (N_18621,N_17423,N_17441);
nand U18622 (N_18622,N_17600,N_17744);
and U18623 (N_18623,N_17316,N_17087);
xor U18624 (N_18624,N_17666,N_17357);
and U18625 (N_18625,N_17831,N_17630);
xnor U18626 (N_18626,N_17967,N_17281);
or U18627 (N_18627,N_17735,N_17358);
nand U18628 (N_18628,N_17220,N_17884);
nand U18629 (N_18629,N_17842,N_17892);
nand U18630 (N_18630,N_17288,N_17872);
or U18631 (N_18631,N_17338,N_17091);
nand U18632 (N_18632,N_17634,N_17176);
nor U18633 (N_18633,N_17045,N_17523);
nor U18634 (N_18634,N_17539,N_17671);
nor U18635 (N_18635,N_17386,N_17109);
nand U18636 (N_18636,N_17317,N_17512);
and U18637 (N_18637,N_17049,N_17648);
nor U18638 (N_18638,N_17280,N_17149);
and U18639 (N_18639,N_17883,N_17871);
or U18640 (N_18640,N_17375,N_17920);
nand U18641 (N_18641,N_17325,N_17901);
nor U18642 (N_18642,N_17578,N_17956);
or U18643 (N_18643,N_17762,N_17508);
nor U18644 (N_18644,N_17672,N_17460);
or U18645 (N_18645,N_17680,N_17135);
nor U18646 (N_18646,N_17911,N_17941);
and U18647 (N_18647,N_17370,N_17885);
nor U18648 (N_18648,N_17456,N_17974);
xnor U18649 (N_18649,N_17926,N_17103);
nand U18650 (N_18650,N_17241,N_17815);
or U18651 (N_18651,N_17445,N_17608);
nand U18652 (N_18652,N_17519,N_17465);
or U18653 (N_18653,N_17178,N_17278);
and U18654 (N_18654,N_17731,N_17276);
nand U18655 (N_18655,N_17061,N_17510);
or U18656 (N_18656,N_17770,N_17577);
nor U18657 (N_18657,N_17465,N_17742);
and U18658 (N_18658,N_17787,N_17941);
nand U18659 (N_18659,N_17638,N_17651);
or U18660 (N_18660,N_17818,N_17638);
nand U18661 (N_18661,N_17771,N_17579);
and U18662 (N_18662,N_17990,N_17223);
nand U18663 (N_18663,N_17844,N_17767);
nor U18664 (N_18664,N_17715,N_17526);
nand U18665 (N_18665,N_17577,N_17967);
nor U18666 (N_18666,N_17912,N_17123);
nor U18667 (N_18667,N_17362,N_17594);
nand U18668 (N_18668,N_17406,N_17248);
nor U18669 (N_18669,N_17886,N_17144);
and U18670 (N_18670,N_17593,N_17163);
nor U18671 (N_18671,N_17348,N_17028);
nand U18672 (N_18672,N_17421,N_17813);
and U18673 (N_18673,N_17973,N_17592);
and U18674 (N_18674,N_17265,N_17998);
or U18675 (N_18675,N_17594,N_17164);
or U18676 (N_18676,N_17184,N_17518);
nand U18677 (N_18677,N_17003,N_17431);
nand U18678 (N_18678,N_17285,N_17751);
nand U18679 (N_18679,N_17918,N_17126);
and U18680 (N_18680,N_17582,N_17433);
nand U18681 (N_18681,N_17172,N_17825);
nand U18682 (N_18682,N_17329,N_17622);
nor U18683 (N_18683,N_17077,N_17940);
xnor U18684 (N_18684,N_17462,N_17800);
or U18685 (N_18685,N_17118,N_17469);
and U18686 (N_18686,N_17080,N_17301);
nor U18687 (N_18687,N_17885,N_17324);
nand U18688 (N_18688,N_17576,N_17409);
and U18689 (N_18689,N_17943,N_17183);
nor U18690 (N_18690,N_17552,N_17000);
nand U18691 (N_18691,N_17255,N_17728);
or U18692 (N_18692,N_17339,N_17335);
or U18693 (N_18693,N_17225,N_17143);
nand U18694 (N_18694,N_17631,N_17373);
nor U18695 (N_18695,N_17237,N_17590);
or U18696 (N_18696,N_17785,N_17968);
or U18697 (N_18697,N_17089,N_17921);
and U18698 (N_18698,N_17081,N_17669);
and U18699 (N_18699,N_17380,N_17998);
nand U18700 (N_18700,N_17881,N_17731);
nor U18701 (N_18701,N_17715,N_17413);
and U18702 (N_18702,N_17150,N_17016);
nand U18703 (N_18703,N_17118,N_17659);
and U18704 (N_18704,N_17478,N_17755);
or U18705 (N_18705,N_17317,N_17498);
nand U18706 (N_18706,N_17472,N_17249);
or U18707 (N_18707,N_17890,N_17780);
nor U18708 (N_18708,N_17245,N_17389);
or U18709 (N_18709,N_17402,N_17078);
xor U18710 (N_18710,N_17337,N_17282);
xnor U18711 (N_18711,N_17200,N_17863);
and U18712 (N_18712,N_17691,N_17053);
nand U18713 (N_18713,N_17208,N_17527);
xnor U18714 (N_18714,N_17209,N_17159);
nand U18715 (N_18715,N_17904,N_17647);
or U18716 (N_18716,N_17147,N_17327);
nor U18717 (N_18717,N_17570,N_17397);
and U18718 (N_18718,N_17341,N_17785);
or U18719 (N_18719,N_17585,N_17232);
nor U18720 (N_18720,N_17860,N_17030);
nand U18721 (N_18721,N_17995,N_17730);
or U18722 (N_18722,N_17595,N_17776);
nor U18723 (N_18723,N_17996,N_17402);
nor U18724 (N_18724,N_17362,N_17091);
nand U18725 (N_18725,N_17800,N_17066);
xnor U18726 (N_18726,N_17060,N_17980);
nand U18727 (N_18727,N_17551,N_17031);
or U18728 (N_18728,N_17337,N_17969);
nand U18729 (N_18729,N_17678,N_17192);
or U18730 (N_18730,N_17529,N_17322);
nand U18731 (N_18731,N_17333,N_17848);
xor U18732 (N_18732,N_17821,N_17068);
or U18733 (N_18733,N_17324,N_17758);
xnor U18734 (N_18734,N_17864,N_17630);
or U18735 (N_18735,N_17978,N_17638);
xor U18736 (N_18736,N_17633,N_17038);
or U18737 (N_18737,N_17324,N_17476);
or U18738 (N_18738,N_17013,N_17639);
nor U18739 (N_18739,N_17902,N_17691);
nor U18740 (N_18740,N_17507,N_17808);
nand U18741 (N_18741,N_17607,N_17491);
or U18742 (N_18742,N_17493,N_17301);
nand U18743 (N_18743,N_17396,N_17961);
nand U18744 (N_18744,N_17701,N_17836);
or U18745 (N_18745,N_17654,N_17786);
xnor U18746 (N_18746,N_17988,N_17181);
xor U18747 (N_18747,N_17571,N_17438);
or U18748 (N_18748,N_17461,N_17059);
xnor U18749 (N_18749,N_17617,N_17867);
nor U18750 (N_18750,N_17234,N_17205);
xor U18751 (N_18751,N_17340,N_17191);
or U18752 (N_18752,N_17522,N_17104);
nor U18753 (N_18753,N_17505,N_17072);
xnor U18754 (N_18754,N_17030,N_17739);
xnor U18755 (N_18755,N_17112,N_17963);
nand U18756 (N_18756,N_17387,N_17027);
nor U18757 (N_18757,N_17925,N_17772);
nor U18758 (N_18758,N_17288,N_17007);
xor U18759 (N_18759,N_17905,N_17409);
nand U18760 (N_18760,N_17178,N_17325);
nor U18761 (N_18761,N_17333,N_17684);
and U18762 (N_18762,N_17227,N_17184);
and U18763 (N_18763,N_17725,N_17824);
and U18764 (N_18764,N_17950,N_17191);
and U18765 (N_18765,N_17146,N_17719);
and U18766 (N_18766,N_17648,N_17771);
nand U18767 (N_18767,N_17390,N_17828);
nand U18768 (N_18768,N_17930,N_17393);
and U18769 (N_18769,N_17077,N_17611);
xnor U18770 (N_18770,N_17175,N_17046);
or U18771 (N_18771,N_17019,N_17725);
xor U18772 (N_18772,N_17044,N_17257);
nand U18773 (N_18773,N_17029,N_17696);
and U18774 (N_18774,N_17198,N_17817);
xor U18775 (N_18775,N_17216,N_17947);
nand U18776 (N_18776,N_17266,N_17203);
xor U18777 (N_18777,N_17065,N_17145);
and U18778 (N_18778,N_17960,N_17554);
or U18779 (N_18779,N_17404,N_17179);
or U18780 (N_18780,N_17874,N_17586);
and U18781 (N_18781,N_17592,N_17523);
and U18782 (N_18782,N_17222,N_17988);
nand U18783 (N_18783,N_17772,N_17683);
and U18784 (N_18784,N_17502,N_17398);
or U18785 (N_18785,N_17446,N_17726);
or U18786 (N_18786,N_17260,N_17830);
nand U18787 (N_18787,N_17949,N_17946);
xor U18788 (N_18788,N_17961,N_17397);
or U18789 (N_18789,N_17584,N_17243);
or U18790 (N_18790,N_17803,N_17962);
xor U18791 (N_18791,N_17566,N_17635);
and U18792 (N_18792,N_17676,N_17473);
or U18793 (N_18793,N_17222,N_17555);
or U18794 (N_18794,N_17919,N_17910);
and U18795 (N_18795,N_17451,N_17577);
and U18796 (N_18796,N_17343,N_17626);
nand U18797 (N_18797,N_17193,N_17594);
and U18798 (N_18798,N_17980,N_17466);
and U18799 (N_18799,N_17711,N_17222);
and U18800 (N_18800,N_17572,N_17495);
or U18801 (N_18801,N_17009,N_17389);
and U18802 (N_18802,N_17502,N_17261);
or U18803 (N_18803,N_17629,N_17728);
xor U18804 (N_18804,N_17121,N_17270);
and U18805 (N_18805,N_17528,N_17204);
and U18806 (N_18806,N_17103,N_17344);
or U18807 (N_18807,N_17314,N_17556);
and U18808 (N_18808,N_17050,N_17972);
xnor U18809 (N_18809,N_17539,N_17118);
nor U18810 (N_18810,N_17059,N_17111);
and U18811 (N_18811,N_17248,N_17587);
nor U18812 (N_18812,N_17678,N_17720);
or U18813 (N_18813,N_17630,N_17215);
nand U18814 (N_18814,N_17716,N_17493);
nand U18815 (N_18815,N_17714,N_17406);
nand U18816 (N_18816,N_17019,N_17736);
nor U18817 (N_18817,N_17850,N_17119);
or U18818 (N_18818,N_17098,N_17011);
and U18819 (N_18819,N_17909,N_17321);
nand U18820 (N_18820,N_17655,N_17052);
nor U18821 (N_18821,N_17076,N_17474);
nand U18822 (N_18822,N_17506,N_17657);
and U18823 (N_18823,N_17588,N_17005);
nand U18824 (N_18824,N_17938,N_17701);
or U18825 (N_18825,N_17840,N_17347);
and U18826 (N_18826,N_17877,N_17694);
nand U18827 (N_18827,N_17437,N_17203);
xnor U18828 (N_18828,N_17201,N_17377);
nand U18829 (N_18829,N_17673,N_17693);
nand U18830 (N_18830,N_17530,N_17989);
nor U18831 (N_18831,N_17692,N_17172);
and U18832 (N_18832,N_17707,N_17120);
or U18833 (N_18833,N_17335,N_17205);
or U18834 (N_18834,N_17140,N_17296);
nand U18835 (N_18835,N_17943,N_17746);
nor U18836 (N_18836,N_17137,N_17934);
and U18837 (N_18837,N_17717,N_17981);
nor U18838 (N_18838,N_17515,N_17948);
nor U18839 (N_18839,N_17559,N_17184);
nand U18840 (N_18840,N_17418,N_17736);
nand U18841 (N_18841,N_17318,N_17490);
and U18842 (N_18842,N_17142,N_17538);
xnor U18843 (N_18843,N_17449,N_17150);
nor U18844 (N_18844,N_17391,N_17711);
xnor U18845 (N_18845,N_17567,N_17006);
nand U18846 (N_18846,N_17016,N_17732);
nand U18847 (N_18847,N_17105,N_17571);
nand U18848 (N_18848,N_17158,N_17143);
nor U18849 (N_18849,N_17385,N_17160);
nor U18850 (N_18850,N_17192,N_17117);
nand U18851 (N_18851,N_17956,N_17997);
nor U18852 (N_18852,N_17837,N_17329);
xor U18853 (N_18853,N_17337,N_17679);
and U18854 (N_18854,N_17339,N_17796);
nor U18855 (N_18855,N_17543,N_17989);
nor U18856 (N_18856,N_17201,N_17155);
nor U18857 (N_18857,N_17155,N_17944);
nor U18858 (N_18858,N_17001,N_17159);
nand U18859 (N_18859,N_17569,N_17483);
or U18860 (N_18860,N_17508,N_17837);
xor U18861 (N_18861,N_17460,N_17892);
nor U18862 (N_18862,N_17923,N_17565);
xor U18863 (N_18863,N_17698,N_17907);
or U18864 (N_18864,N_17411,N_17303);
and U18865 (N_18865,N_17416,N_17169);
xor U18866 (N_18866,N_17261,N_17170);
nor U18867 (N_18867,N_17471,N_17562);
nand U18868 (N_18868,N_17474,N_17904);
nor U18869 (N_18869,N_17897,N_17617);
nand U18870 (N_18870,N_17232,N_17330);
nor U18871 (N_18871,N_17002,N_17264);
nor U18872 (N_18872,N_17052,N_17205);
nor U18873 (N_18873,N_17148,N_17291);
or U18874 (N_18874,N_17920,N_17660);
xor U18875 (N_18875,N_17777,N_17659);
xnor U18876 (N_18876,N_17390,N_17949);
xnor U18877 (N_18877,N_17565,N_17786);
nor U18878 (N_18878,N_17398,N_17602);
or U18879 (N_18879,N_17304,N_17274);
or U18880 (N_18880,N_17630,N_17751);
nor U18881 (N_18881,N_17480,N_17278);
or U18882 (N_18882,N_17922,N_17490);
xor U18883 (N_18883,N_17999,N_17923);
nor U18884 (N_18884,N_17900,N_17682);
or U18885 (N_18885,N_17648,N_17610);
nand U18886 (N_18886,N_17539,N_17553);
and U18887 (N_18887,N_17167,N_17134);
and U18888 (N_18888,N_17667,N_17766);
nand U18889 (N_18889,N_17695,N_17911);
nand U18890 (N_18890,N_17493,N_17811);
xnor U18891 (N_18891,N_17824,N_17577);
nor U18892 (N_18892,N_17575,N_17571);
xnor U18893 (N_18893,N_17801,N_17804);
nand U18894 (N_18894,N_17607,N_17480);
and U18895 (N_18895,N_17552,N_17453);
nand U18896 (N_18896,N_17400,N_17587);
or U18897 (N_18897,N_17782,N_17965);
nand U18898 (N_18898,N_17463,N_17376);
nand U18899 (N_18899,N_17490,N_17435);
nand U18900 (N_18900,N_17727,N_17647);
and U18901 (N_18901,N_17457,N_17881);
xor U18902 (N_18902,N_17988,N_17952);
and U18903 (N_18903,N_17667,N_17422);
nand U18904 (N_18904,N_17700,N_17771);
nor U18905 (N_18905,N_17186,N_17340);
nand U18906 (N_18906,N_17085,N_17466);
and U18907 (N_18907,N_17559,N_17398);
or U18908 (N_18908,N_17617,N_17338);
nor U18909 (N_18909,N_17993,N_17593);
and U18910 (N_18910,N_17099,N_17310);
and U18911 (N_18911,N_17346,N_17489);
nor U18912 (N_18912,N_17780,N_17380);
nor U18913 (N_18913,N_17739,N_17221);
nor U18914 (N_18914,N_17914,N_17043);
and U18915 (N_18915,N_17902,N_17440);
or U18916 (N_18916,N_17242,N_17248);
nand U18917 (N_18917,N_17751,N_17842);
nor U18918 (N_18918,N_17978,N_17606);
and U18919 (N_18919,N_17806,N_17995);
or U18920 (N_18920,N_17609,N_17649);
and U18921 (N_18921,N_17845,N_17818);
or U18922 (N_18922,N_17086,N_17495);
and U18923 (N_18923,N_17693,N_17934);
nor U18924 (N_18924,N_17461,N_17267);
xnor U18925 (N_18925,N_17316,N_17095);
or U18926 (N_18926,N_17027,N_17619);
or U18927 (N_18927,N_17472,N_17621);
nor U18928 (N_18928,N_17974,N_17388);
xor U18929 (N_18929,N_17849,N_17685);
nand U18930 (N_18930,N_17044,N_17945);
and U18931 (N_18931,N_17920,N_17812);
and U18932 (N_18932,N_17950,N_17256);
and U18933 (N_18933,N_17795,N_17487);
nand U18934 (N_18934,N_17395,N_17390);
nor U18935 (N_18935,N_17952,N_17821);
xor U18936 (N_18936,N_17500,N_17035);
xnor U18937 (N_18937,N_17051,N_17878);
xor U18938 (N_18938,N_17995,N_17472);
and U18939 (N_18939,N_17774,N_17054);
nor U18940 (N_18940,N_17437,N_17696);
xnor U18941 (N_18941,N_17112,N_17726);
and U18942 (N_18942,N_17191,N_17447);
or U18943 (N_18943,N_17075,N_17442);
nor U18944 (N_18944,N_17628,N_17094);
or U18945 (N_18945,N_17187,N_17795);
nand U18946 (N_18946,N_17059,N_17719);
xor U18947 (N_18947,N_17512,N_17724);
or U18948 (N_18948,N_17460,N_17089);
xor U18949 (N_18949,N_17425,N_17780);
and U18950 (N_18950,N_17878,N_17620);
xor U18951 (N_18951,N_17928,N_17261);
nor U18952 (N_18952,N_17158,N_17444);
nor U18953 (N_18953,N_17387,N_17504);
xnor U18954 (N_18954,N_17093,N_17553);
or U18955 (N_18955,N_17590,N_17143);
nor U18956 (N_18956,N_17258,N_17502);
xor U18957 (N_18957,N_17154,N_17089);
xor U18958 (N_18958,N_17720,N_17654);
or U18959 (N_18959,N_17212,N_17257);
and U18960 (N_18960,N_17713,N_17039);
nand U18961 (N_18961,N_17716,N_17689);
and U18962 (N_18962,N_17785,N_17953);
nor U18963 (N_18963,N_17098,N_17418);
nor U18964 (N_18964,N_17970,N_17619);
nor U18965 (N_18965,N_17458,N_17681);
nand U18966 (N_18966,N_17392,N_17465);
and U18967 (N_18967,N_17071,N_17368);
or U18968 (N_18968,N_17545,N_17739);
or U18969 (N_18969,N_17996,N_17933);
xnor U18970 (N_18970,N_17424,N_17807);
nor U18971 (N_18971,N_17772,N_17289);
nor U18972 (N_18972,N_17373,N_17332);
or U18973 (N_18973,N_17041,N_17153);
xor U18974 (N_18974,N_17265,N_17241);
nor U18975 (N_18975,N_17323,N_17364);
xnor U18976 (N_18976,N_17259,N_17468);
and U18977 (N_18977,N_17052,N_17469);
and U18978 (N_18978,N_17333,N_17521);
nor U18979 (N_18979,N_17833,N_17561);
or U18980 (N_18980,N_17673,N_17130);
xnor U18981 (N_18981,N_17990,N_17989);
nand U18982 (N_18982,N_17842,N_17956);
nor U18983 (N_18983,N_17202,N_17751);
and U18984 (N_18984,N_17956,N_17275);
and U18985 (N_18985,N_17261,N_17423);
xnor U18986 (N_18986,N_17081,N_17310);
nor U18987 (N_18987,N_17083,N_17301);
or U18988 (N_18988,N_17619,N_17545);
or U18989 (N_18989,N_17642,N_17539);
xnor U18990 (N_18990,N_17173,N_17972);
nand U18991 (N_18991,N_17594,N_17809);
or U18992 (N_18992,N_17028,N_17365);
nor U18993 (N_18993,N_17678,N_17372);
nand U18994 (N_18994,N_17715,N_17889);
xor U18995 (N_18995,N_17077,N_17525);
or U18996 (N_18996,N_17869,N_17806);
nor U18997 (N_18997,N_17474,N_17998);
xnor U18998 (N_18998,N_17899,N_17710);
nor U18999 (N_18999,N_17434,N_17207);
and U19000 (N_19000,N_18087,N_18388);
nor U19001 (N_19001,N_18524,N_18231);
or U19002 (N_19002,N_18861,N_18465);
and U19003 (N_19003,N_18169,N_18393);
nand U19004 (N_19004,N_18698,N_18707);
xor U19005 (N_19005,N_18421,N_18064);
or U19006 (N_19006,N_18317,N_18450);
nand U19007 (N_19007,N_18301,N_18732);
nand U19008 (N_19008,N_18383,N_18044);
and U19009 (N_19009,N_18187,N_18831);
or U19010 (N_19010,N_18676,N_18077);
xnor U19011 (N_19011,N_18734,N_18254);
xnor U19012 (N_19012,N_18737,N_18931);
nor U19013 (N_19013,N_18036,N_18785);
nand U19014 (N_19014,N_18381,N_18017);
and U19015 (N_19015,N_18948,N_18360);
nand U19016 (N_19016,N_18350,N_18150);
or U19017 (N_19017,N_18043,N_18429);
xnor U19018 (N_19018,N_18533,N_18134);
nor U19019 (N_19019,N_18670,N_18438);
nand U19020 (N_19020,N_18509,N_18325);
nor U19021 (N_19021,N_18523,N_18274);
nor U19022 (N_19022,N_18113,N_18428);
xnor U19023 (N_19023,N_18129,N_18151);
or U19024 (N_19024,N_18655,N_18309);
xnor U19025 (N_19025,N_18105,N_18722);
nor U19026 (N_19026,N_18194,N_18690);
xnor U19027 (N_19027,N_18142,N_18654);
xnor U19028 (N_19028,N_18336,N_18426);
nor U19029 (N_19029,N_18100,N_18409);
nand U19030 (N_19030,N_18161,N_18266);
or U19031 (N_19031,N_18471,N_18294);
or U19032 (N_19032,N_18781,N_18770);
nor U19033 (N_19033,N_18673,N_18716);
nor U19034 (N_19034,N_18267,N_18636);
nor U19035 (N_19035,N_18516,N_18567);
and U19036 (N_19036,N_18678,N_18756);
and U19037 (N_19037,N_18282,N_18370);
xnor U19038 (N_19038,N_18920,N_18792);
or U19039 (N_19039,N_18957,N_18090);
nand U19040 (N_19040,N_18838,N_18034);
xnor U19041 (N_19041,N_18600,N_18379);
and U19042 (N_19042,N_18273,N_18102);
nand U19043 (N_19043,N_18940,N_18758);
nor U19044 (N_19044,N_18631,N_18369);
and U19045 (N_19045,N_18789,N_18629);
or U19046 (N_19046,N_18660,N_18641);
nor U19047 (N_19047,N_18444,N_18135);
nand U19048 (N_19048,N_18705,N_18612);
xor U19049 (N_19049,N_18445,N_18932);
and U19050 (N_19050,N_18053,N_18634);
and U19051 (N_19051,N_18299,N_18606);
xnor U19052 (N_19052,N_18796,N_18529);
nand U19053 (N_19053,N_18284,N_18063);
nor U19054 (N_19054,N_18961,N_18762);
nor U19055 (N_19055,N_18624,N_18632);
xor U19056 (N_19056,N_18000,N_18354);
and U19057 (N_19057,N_18846,N_18422);
nand U19058 (N_19058,N_18803,N_18452);
xor U19059 (N_19059,N_18318,N_18912);
nand U19060 (N_19060,N_18345,N_18688);
or U19061 (N_19061,N_18843,N_18917);
and U19062 (N_19062,N_18414,N_18699);
nand U19063 (N_19063,N_18595,N_18504);
nand U19064 (N_19064,N_18559,N_18853);
xnor U19065 (N_19065,N_18942,N_18158);
nor U19066 (N_19066,N_18442,N_18333);
nand U19067 (N_19067,N_18221,N_18390);
or U19068 (N_19068,N_18296,N_18331);
and U19069 (N_19069,N_18164,N_18435);
and U19070 (N_19070,N_18073,N_18585);
or U19071 (N_19071,N_18860,N_18922);
xnor U19072 (N_19072,N_18375,N_18479);
xnor U19073 (N_19073,N_18607,N_18462);
and U19074 (N_19074,N_18304,N_18014);
and U19075 (N_19075,N_18108,N_18786);
nand U19076 (N_19076,N_18481,N_18834);
nor U19077 (N_19077,N_18674,N_18235);
nand U19078 (N_19078,N_18996,N_18950);
nand U19079 (N_19079,N_18021,N_18328);
and U19080 (N_19080,N_18168,N_18742);
or U19081 (N_19081,N_18818,N_18569);
xnor U19082 (N_19082,N_18419,N_18866);
nand U19083 (N_19083,N_18425,N_18146);
xnor U19084 (N_19084,N_18128,N_18602);
or U19085 (N_19085,N_18233,N_18280);
xor U19086 (N_19086,N_18039,N_18209);
and U19087 (N_19087,N_18415,N_18764);
and U19088 (N_19088,N_18951,N_18248);
and U19089 (N_19089,N_18675,N_18116);
nor U19090 (N_19090,N_18778,N_18589);
or U19091 (N_19091,N_18788,N_18813);
and U19092 (N_19092,N_18122,N_18175);
and U19093 (N_19093,N_18069,N_18038);
xnor U19094 (N_19094,N_18171,N_18439);
nor U19095 (N_19095,N_18972,N_18577);
and U19096 (N_19096,N_18224,N_18976);
and U19097 (N_19097,N_18290,N_18198);
nand U19098 (N_19098,N_18059,N_18561);
or U19099 (N_19099,N_18658,N_18794);
xor U19100 (N_19100,N_18547,N_18828);
and U19101 (N_19101,N_18407,N_18287);
nor U19102 (N_19102,N_18588,N_18054);
nand U19103 (N_19103,N_18625,N_18747);
nor U19104 (N_19104,N_18736,N_18313);
or U19105 (N_19105,N_18526,N_18342);
and U19106 (N_19106,N_18033,N_18459);
and U19107 (N_19107,N_18195,N_18605);
nor U19108 (N_19108,N_18197,N_18847);
nor U19109 (N_19109,N_18238,N_18291);
or U19110 (N_19110,N_18941,N_18511);
and U19111 (N_19111,N_18928,N_18011);
or U19112 (N_19112,N_18619,N_18232);
nor U19113 (N_19113,N_18537,N_18825);
nor U19114 (N_19114,N_18946,N_18443);
and U19115 (N_19115,N_18045,N_18298);
and U19116 (N_19116,N_18423,N_18987);
nand U19117 (N_19117,N_18321,N_18215);
or U19118 (N_19118,N_18695,N_18293);
nor U19119 (N_19119,N_18540,N_18133);
xor U19120 (N_19120,N_18089,N_18637);
nand U19121 (N_19121,N_18316,N_18712);
xnor U19122 (N_19122,N_18289,N_18387);
or U19123 (N_19123,N_18130,N_18149);
nand U19124 (N_19124,N_18358,N_18052);
nor U19125 (N_19125,N_18012,N_18303);
xor U19126 (N_19126,N_18188,N_18018);
and U19127 (N_19127,N_18889,N_18178);
or U19128 (N_19128,N_18022,N_18103);
xnor U19129 (N_19129,N_18858,N_18728);
xor U19130 (N_19130,N_18009,N_18020);
xor U19131 (N_19131,N_18955,N_18708);
and U19132 (N_19132,N_18397,N_18802);
or U19133 (N_19133,N_18751,N_18019);
xnor U19134 (N_19134,N_18935,N_18867);
or U19135 (N_19135,N_18973,N_18251);
xor U19136 (N_19136,N_18353,N_18683);
nor U19137 (N_19137,N_18385,N_18242);
and U19138 (N_19138,N_18026,N_18687);
nor U19139 (N_19139,N_18906,N_18568);
or U19140 (N_19140,N_18630,N_18621);
and U19141 (N_19141,N_18677,N_18418);
and U19142 (N_19142,N_18189,N_18835);
nand U19143 (N_19143,N_18545,N_18686);
nor U19144 (N_19144,N_18320,N_18306);
nor U19145 (N_19145,N_18138,N_18801);
and U19146 (N_19146,N_18013,N_18220);
and U19147 (N_19147,N_18141,N_18148);
or U19148 (N_19148,N_18587,N_18964);
or U19149 (N_19149,N_18276,N_18469);
xor U19150 (N_19150,N_18863,N_18229);
xnor U19151 (N_19151,N_18015,N_18579);
xor U19152 (N_19152,N_18954,N_18112);
nand U19153 (N_19153,N_18900,N_18272);
xnor U19154 (N_19154,N_18528,N_18804);
xor U19155 (N_19155,N_18118,N_18978);
xnor U19156 (N_19156,N_18093,N_18190);
or U19157 (N_19157,N_18472,N_18985);
and U19158 (N_19158,N_18771,N_18633);
nor U19159 (N_19159,N_18639,N_18517);
xor U19160 (N_19160,N_18373,N_18115);
xnor U19161 (N_19161,N_18689,N_18875);
or U19162 (N_19162,N_18608,N_18650);
nor U19163 (N_19163,N_18894,N_18202);
or U19164 (N_19164,N_18721,N_18508);
and U19165 (N_19165,N_18498,N_18652);
and U19166 (N_19166,N_18056,N_18427);
xor U19167 (N_19167,N_18406,N_18389);
nand U19168 (N_19168,N_18004,N_18774);
or U19169 (N_19169,N_18307,N_18916);
nor U19170 (N_19170,N_18570,N_18919);
nor U19171 (N_19171,N_18692,N_18259);
or U19172 (N_19172,N_18213,N_18343);
and U19173 (N_19173,N_18147,N_18271);
nor U19174 (N_19174,N_18520,N_18177);
nor U19175 (N_19175,N_18971,N_18338);
xor U19176 (N_19176,N_18864,N_18827);
and U19177 (N_19177,N_18696,N_18656);
xnor U19178 (N_19178,N_18558,N_18880);
xnor U19179 (N_19179,N_18535,N_18902);
or U19180 (N_19180,N_18031,N_18024);
xnor U19181 (N_19181,N_18404,N_18706);
nand U19182 (N_19182,N_18349,N_18643);
or U19183 (N_19183,N_18352,N_18268);
xnor U19184 (N_19184,N_18058,N_18230);
or U19185 (N_19185,N_18448,N_18510);
and U19186 (N_19186,N_18876,N_18051);
nand U19187 (N_19187,N_18417,N_18709);
nor U19188 (N_19188,N_18960,N_18492);
and U19189 (N_19189,N_18275,N_18784);
nor U19190 (N_19190,N_18743,N_18735);
or U19191 (N_19191,N_18095,N_18560);
nor U19192 (N_19192,N_18974,N_18237);
xnor U19193 (N_19193,N_18967,N_18890);
nand U19194 (N_19194,N_18140,N_18200);
and U19195 (N_19195,N_18793,N_18490);
nand U19196 (N_19196,N_18206,N_18027);
and U19197 (N_19197,N_18779,N_18211);
nand U19198 (N_19198,N_18286,N_18071);
nand U19199 (N_19199,N_18653,N_18999);
or U19200 (N_19200,N_18505,N_18374);
nor U19201 (N_19201,N_18549,N_18981);
or U19202 (N_19202,N_18111,N_18433);
nor U19203 (N_19203,N_18424,N_18512);
nor U19204 (N_19204,N_18522,N_18649);
xor U19205 (N_19205,N_18196,N_18808);
xnor U19206 (N_19206,N_18185,N_18821);
and U19207 (N_19207,N_18944,N_18836);
nor U19208 (N_19208,N_18503,N_18700);
xor U19209 (N_19209,N_18346,N_18131);
or U19210 (N_19210,N_18088,N_18344);
or U19211 (N_19211,N_18485,N_18207);
or U19212 (N_19212,N_18183,N_18730);
and U19213 (N_19213,N_18302,N_18277);
nor U19214 (N_19214,N_18476,N_18155);
and U19215 (N_19215,N_18651,N_18401);
xnor U19216 (N_19216,N_18800,N_18092);
and U19217 (N_19217,N_18816,N_18319);
nor U19218 (N_19218,N_18873,N_18070);
and U19219 (N_19219,N_18893,N_18787);
and U19220 (N_19220,N_18556,N_18888);
xnor U19221 (N_19221,N_18430,N_18543);
nor U19222 (N_19222,N_18253,N_18123);
or U19223 (N_19223,N_18934,N_18578);
or U19224 (N_19224,N_18548,N_18852);
and U19225 (N_19225,N_18691,N_18635);
and U19226 (N_19226,N_18661,N_18480);
xnor U19227 (N_19227,N_18977,N_18250);
and U19228 (N_19228,N_18455,N_18312);
nand U19229 (N_19229,N_18574,N_18377);
xor U19230 (N_19230,N_18768,N_18008);
or U19231 (N_19231,N_18868,N_18798);
nand U19232 (N_19232,N_18005,N_18885);
or U19233 (N_19233,N_18182,N_18192);
and U19234 (N_19234,N_18519,N_18173);
nand U19235 (N_19235,N_18482,N_18534);
nor U19236 (N_19236,N_18084,N_18530);
and U19237 (N_19237,N_18101,N_18351);
xnor U19238 (N_19238,N_18822,N_18870);
xor U19239 (N_19239,N_18191,N_18878);
xor U19240 (N_19240,N_18361,N_18884);
nand U19241 (N_19241,N_18311,N_18127);
nand U19242 (N_19242,N_18887,N_18292);
nor U19243 (N_19243,N_18982,N_18616);
nand U19244 (N_19244,N_18174,N_18072);
or U19245 (N_19245,N_18094,N_18257);
nand U19246 (N_19246,N_18812,N_18667);
xor U19247 (N_19247,N_18693,N_18041);
nand U19248 (N_19248,N_18049,N_18965);
nor U19249 (N_19249,N_18850,N_18769);
and U19250 (N_19250,N_18162,N_18760);
and U19251 (N_19251,N_18791,N_18262);
or U19252 (N_19252,N_18217,N_18456);
nand U19253 (N_19253,N_18029,N_18557);
and U19254 (N_19254,N_18979,N_18753);
or U19255 (N_19255,N_18565,N_18943);
or U19256 (N_19256,N_18939,N_18288);
xnor U19257 (N_19257,N_18980,N_18823);
nor U19258 (N_19258,N_18413,N_18926);
nor U19259 (N_19259,N_18581,N_18380);
nand U19260 (N_19260,N_18119,N_18170);
or U19261 (N_19261,N_18341,N_18810);
nor U19262 (N_19262,N_18120,N_18348);
xor U19263 (N_19263,N_18305,N_18541);
and U19264 (N_19264,N_18368,N_18962);
nand U19265 (N_19265,N_18984,N_18615);
nand U19266 (N_19266,N_18367,N_18945);
nand U19267 (N_19267,N_18553,N_18820);
or U19268 (N_19268,N_18324,N_18933);
and U19269 (N_19269,N_18260,N_18359);
or U19270 (N_19270,N_18205,N_18256);
and U19271 (N_19271,N_18132,N_18061);
xnor U19272 (N_19272,N_18037,N_18062);
xor U19273 (N_19273,N_18703,N_18738);
and U19274 (N_19274,N_18269,N_18644);
and U19275 (N_19275,N_18405,N_18592);
xnor U19276 (N_19276,N_18486,N_18694);
or U19277 (N_19277,N_18844,N_18114);
nor U19278 (N_19278,N_18109,N_18335);
and U19279 (N_19279,N_18766,N_18872);
nand U19280 (N_19280,N_18614,N_18908);
xnor U19281 (N_19281,N_18672,N_18775);
nand U19282 (N_19282,N_18125,N_18881);
xnor U19283 (N_19283,N_18966,N_18782);
nor U19284 (N_19284,N_18222,N_18270);
nor U19285 (N_19285,N_18603,N_18204);
or U19286 (N_19286,N_18006,N_18468);
and U19287 (N_19287,N_18376,N_18583);
nor U19288 (N_19288,N_18921,N_18536);
nor U19289 (N_19289,N_18216,N_18153);
nor U19290 (N_19290,N_18117,N_18078);
and U19291 (N_19291,N_18842,N_18514);
xor U19292 (N_19292,N_18484,N_18487);
or U19293 (N_19293,N_18680,N_18930);
nor U19294 (N_19294,N_18573,N_18327);
or U19295 (N_19295,N_18493,N_18744);
xnor U19296 (N_19296,N_18532,N_18003);
xnor U19297 (N_19297,N_18483,N_18457);
xnor U19298 (N_19298,N_18797,N_18159);
nand U19299 (N_19299,N_18657,N_18028);
nand U19300 (N_19300,N_18461,N_18869);
nand U19301 (N_19301,N_18938,N_18586);
xnor U19302 (N_19302,N_18599,N_18555);
xnor U19303 (N_19303,N_18664,N_18710);
xor U19304 (N_19304,N_18829,N_18521);
and U19305 (N_19305,N_18400,N_18047);
or U19306 (N_19306,N_18899,N_18281);
nor U19307 (N_19307,N_18910,N_18773);
or U19308 (N_19308,N_18826,N_18862);
nand U19309 (N_19309,N_18470,N_18719);
nand U19310 (N_19310,N_18083,N_18139);
and U19311 (N_19311,N_18892,N_18136);
nand U19312 (N_19312,N_18824,N_18339);
and U19313 (N_19313,N_18640,N_18845);
or U19314 (N_19314,N_18068,N_18475);
nor U19315 (N_19315,N_18048,N_18865);
nor U19316 (N_19316,N_18886,N_18152);
nor U19317 (N_19317,N_18225,N_18332);
nor U19318 (N_19318,N_18154,N_18949);
or U19319 (N_19319,N_18563,N_18074);
xor U19320 (N_19320,N_18983,N_18371);
and U19321 (N_19321,N_18546,N_18975);
nand U19322 (N_19322,N_18219,N_18659);
nand U19323 (N_19323,N_18989,N_18193);
xor U19324 (N_19324,N_18249,N_18970);
nand U19325 (N_19325,N_18994,N_18176);
nand U19326 (N_19326,N_18107,N_18988);
xor U19327 (N_19327,N_18697,N_18110);
xnor U19328 (N_19328,N_18882,N_18626);
and U19329 (N_19329,N_18451,N_18628);
nand U19330 (N_19330,N_18066,N_18895);
xor U19331 (N_19331,N_18181,N_18076);
xnor U19332 (N_19332,N_18749,N_18763);
xnor U19333 (N_19333,N_18731,N_18571);
and U19334 (N_19334,N_18898,N_18620);
and U19335 (N_19335,N_18097,N_18780);
and U19336 (N_19336,N_18871,N_18507);
nor U19337 (N_19337,N_18167,N_18909);
and U19338 (N_19338,N_18584,N_18010);
xor U19339 (N_19339,N_18025,N_18372);
and U19340 (N_19340,N_18718,N_18564);
nor U19341 (N_19341,N_18576,N_18096);
nor U19342 (N_19342,N_18723,N_18366);
xnor U19343 (N_19343,N_18638,N_18308);
xor U19344 (N_19344,N_18160,N_18724);
and U19345 (N_19345,N_18488,N_18848);
and U19346 (N_19346,N_18007,N_18434);
xnor U19347 (N_19347,N_18704,N_18601);
and U19348 (N_19348,N_18214,N_18859);
nor U19349 (N_19349,N_18729,N_18610);
xnor U19350 (N_19350,N_18572,N_18740);
or U19351 (N_19351,N_18494,N_18879);
nor U19352 (N_19352,N_18145,N_18236);
xor U19353 (N_19353,N_18923,N_18799);
xnor U19354 (N_19354,N_18441,N_18609);
nor U19355 (N_19355,N_18086,N_18668);
nor U19356 (N_19356,N_18929,N_18958);
xor U19357 (N_19357,N_18410,N_18099);
nor U19358 (N_19358,N_18969,N_18226);
nand U19359 (N_19359,N_18463,N_18079);
and U19360 (N_19360,N_18364,N_18997);
or U19361 (N_19361,N_18499,N_18378);
nand U19362 (N_19362,N_18702,N_18685);
or U19363 (N_19363,N_18454,N_18314);
nand U19364 (N_19364,N_18464,N_18506);
nor U19365 (N_19365,N_18081,N_18727);
nand U19366 (N_19366,N_18566,N_18496);
xor U19367 (N_19367,N_18382,N_18937);
and U19368 (N_19368,N_18806,N_18648);
and U19369 (N_19369,N_18030,N_18542);
nor U19370 (N_19370,N_18085,N_18243);
nor U19371 (N_19371,N_18356,N_18877);
nand U19372 (N_19372,N_18953,N_18416);
nand U19373 (N_19373,N_18491,N_18412);
xnor U19374 (N_19374,N_18227,N_18765);
nor U19375 (N_19375,N_18777,N_18166);
and U19376 (N_19376,N_18671,N_18234);
nand U19377 (N_19377,N_18002,N_18622);
and U19378 (N_19378,N_18995,N_18437);
and U19379 (N_19379,N_18500,N_18901);
and U19380 (N_19380,N_18776,N_18395);
nor U19381 (N_19381,N_18746,N_18244);
nor U19382 (N_19382,N_18896,N_18340);
nand U19383 (N_19383,N_18184,N_18295);
or U19384 (N_19384,N_18913,N_18091);
or U19385 (N_19385,N_18538,N_18046);
xor U19386 (N_19386,N_18497,N_18098);
or U19387 (N_19387,N_18525,N_18172);
nor U19388 (N_19388,N_18050,N_18681);
nor U19389 (N_19389,N_18502,N_18790);
and U19390 (N_19390,N_18322,N_18905);
and U19391 (N_19391,N_18001,N_18082);
nand U19392 (N_19392,N_18725,N_18156);
and U19393 (N_19393,N_18252,N_18642);
or U19394 (N_19394,N_18391,N_18993);
nor U19395 (N_19395,N_18399,N_18246);
or U19396 (N_19396,N_18915,N_18726);
nor U19397 (N_19397,N_18241,N_18598);
or U19398 (N_19398,N_18927,N_18554);
and U19399 (N_19399,N_18701,N_18060);
or U19400 (N_19400,N_18513,N_18446);
and U19401 (N_19401,N_18596,N_18662);
nand U19402 (N_19402,N_18104,N_18362);
and U19403 (N_19403,N_18326,N_18208);
nor U19404 (N_19404,N_18990,N_18597);
xnor U19405 (N_19405,N_18992,N_18436);
nand U19406 (N_19406,N_18714,N_18180);
and U19407 (N_19407,N_18911,N_18411);
xnor U19408 (N_19408,N_18562,N_18330);
nor U19409 (N_19409,N_18466,N_18473);
or U19410 (N_19410,N_18203,N_18363);
nand U19411 (N_19411,N_18042,N_18402);
nand U19412 (N_19412,N_18265,N_18515);
nor U19413 (N_19413,N_18837,N_18539);
nor U19414 (N_19414,N_18285,N_18663);
or U19415 (N_19415,N_18240,N_18279);
or U19416 (N_19416,N_18550,N_18839);
and U19417 (N_19417,N_18495,N_18851);
nor U19418 (N_19418,N_18741,N_18715);
and U19419 (N_19419,N_18575,N_18647);
xnor U19420 (N_19420,N_18199,N_18936);
or U19421 (N_19421,N_18297,N_18925);
xor U19422 (N_19422,N_18106,N_18757);
or U19423 (N_19423,N_18431,N_18713);
nor U19424 (N_19424,N_18186,N_18665);
or U19425 (N_19425,N_18582,N_18748);
xnor U19426 (N_19426,N_18627,N_18239);
nand U19427 (N_19427,N_18717,N_18998);
or U19428 (N_19428,N_18223,N_18057);
nor U19429 (N_19429,N_18807,N_18126);
nor U19430 (N_19430,N_18856,N_18334);
and U19431 (N_19431,N_18329,N_18035);
and U19432 (N_19432,N_18258,N_18263);
nand U19433 (N_19433,N_18590,N_18604);
nor U19434 (N_19434,N_18323,N_18157);
nand U19435 (N_19435,N_18032,N_18067);
nand U19436 (N_19436,N_18874,N_18518);
xnor U19437 (N_19437,N_18392,N_18617);
xnor U19438 (N_19438,N_18750,N_18907);
nor U19439 (N_19439,N_18815,N_18477);
nor U19440 (N_19440,N_18347,N_18355);
nor U19441 (N_19441,N_18245,N_18959);
and U19442 (N_19442,N_18591,N_18761);
nand U19443 (N_19443,N_18300,N_18986);
and U19444 (N_19444,N_18179,N_18337);
and U19445 (N_19445,N_18201,N_18315);
xnor U19446 (N_19446,N_18733,N_18449);
nor U19447 (N_19447,N_18357,N_18551);
or U19448 (N_19448,N_18218,N_18819);
or U19449 (N_19449,N_18531,N_18720);
nor U19450 (N_19450,N_18833,N_18432);
and U19451 (N_19451,N_18857,N_18075);
nor U19452 (N_19452,N_18739,N_18283);
nor U19453 (N_19453,N_18403,N_18165);
nor U19454 (N_19454,N_18817,N_18552);
and U19455 (N_19455,N_18489,N_18121);
or U19456 (N_19456,N_18991,N_18593);
or U19457 (N_19457,N_18918,N_18623);
nor U19458 (N_19458,N_18830,N_18440);
and U19459 (N_19459,N_18016,N_18474);
xor U19460 (N_19460,N_18956,N_18924);
or U19461 (N_19461,N_18646,N_18767);
and U19462 (N_19462,N_18527,N_18023);
or U19463 (N_19463,N_18212,N_18228);
xor U19464 (N_19464,N_18682,N_18811);
nand U19465 (N_19465,N_18772,N_18754);
and U19466 (N_19466,N_18618,N_18752);
nand U19467 (N_19467,N_18613,N_18501);
or U19468 (N_19468,N_18947,N_18447);
xnor U19469 (N_19469,N_18143,N_18055);
or U19470 (N_19470,N_18903,N_18914);
or U19471 (N_19471,N_18645,N_18255);
and U19472 (N_19472,N_18261,N_18759);
nand U19473 (N_19473,N_18783,N_18124);
xor U19474 (N_19474,N_18755,N_18897);
or U19475 (N_19475,N_18420,N_18264);
or U19476 (N_19476,N_18210,N_18040);
xor U19477 (N_19477,N_18065,N_18883);
nor U19478 (N_19478,N_18580,N_18849);
xnor U19479 (N_19479,N_18904,N_18137);
xnor U19480 (N_19480,N_18669,N_18855);
nand U19481 (N_19481,N_18809,N_18666);
nand U19482 (N_19482,N_18795,N_18080);
nor U19483 (N_19483,N_18745,N_18386);
nand U19484 (N_19484,N_18394,N_18805);
and U19485 (N_19485,N_18891,N_18814);
or U19486 (N_19486,N_18453,N_18278);
nor U19487 (N_19487,N_18408,N_18163);
and U19488 (N_19488,N_18952,N_18832);
or U19489 (N_19489,N_18365,N_18478);
and U19490 (N_19490,N_18594,N_18458);
and U19491 (N_19491,N_18396,N_18611);
nand U19492 (N_19492,N_18854,N_18544);
nor U19493 (N_19493,N_18467,N_18684);
or U19494 (N_19494,N_18310,N_18460);
xnor U19495 (N_19495,N_18384,N_18398);
and U19496 (N_19496,N_18711,N_18963);
and U19497 (N_19497,N_18247,N_18841);
nor U19498 (N_19498,N_18679,N_18968);
nor U19499 (N_19499,N_18840,N_18144);
xnor U19500 (N_19500,N_18628,N_18081);
or U19501 (N_19501,N_18964,N_18644);
nor U19502 (N_19502,N_18224,N_18858);
or U19503 (N_19503,N_18584,N_18614);
or U19504 (N_19504,N_18388,N_18888);
nand U19505 (N_19505,N_18023,N_18004);
nand U19506 (N_19506,N_18152,N_18673);
xnor U19507 (N_19507,N_18615,N_18128);
nand U19508 (N_19508,N_18639,N_18760);
xor U19509 (N_19509,N_18847,N_18221);
or U19510 (N_19510,N_18535,N_18655);
nor U19511 (N_19511,N_18175,N_18809);
nor U19512 (N_19512,N_18168,N_18017);
and U19513 (N_19513,N_18822,N_18674);
xnor U19514 (N_19514,N_18672,N_18188);
nand U19515 (N_19515,N_18167,N_18466);
nand U19516 (N_19516,N_18917,N_18644);
and U19517 (N_19517,N_18991,N_18987);
or U19518 (N_19518,N_18335,N_18906);
or U19519 (N_19519,N_18052,N_18512);
nor U19520 (N_19520,N_18712,N_18165);
nor U19521 (N_19521,N_18218,N_18499);
xnor U19522 (N_19522,N_18946,N_18906);
nand U19523 (N_19523,N_18267,N_18067);
nand U19524 (N_19524,N_18362,N_18248);
nand U19525 (N_19525,N_18967,N_18453);
nor U19526 (N_19526,N_18321,N_18595);
and U19527 (N_19527,N_18950,N_18763);
nor U19528 (N_19528,N_18101,N_18345);
or U19529 (N_19529,N_18483,N_18717);
nand U19530 (N_19530,N_18689,N_18329);
xnor U19531 (N_19531,N_18897,N_18065);
nor U19532 (N_19532,N_18600,N_18423);
or U19533 (N_19533,N_18312,N_18712);
or U19534 (N_19534,N_18214,N_18359);
or U19535 (N_19535,N_18839,N_18306);
and U19536 (N_19536,N_18843,N_18840);
xnor U19537 (N_19537,N_18816,N_18886);
xor U19538 (N_19538,N_18465,N_18937);
nor U19539 (N_19539,N_18061,N_18328);
or U19540 (N_19540,N_18949,N_18132);
or U19541 (N_19541,N_18865,N_18446);
xor U19542 (N_19542,N_18131,N_18831);
and U19543 (N_19543,N_18558,N_18704);
and U19544 (N_19544,N_18192,N_18014);
and U19545 (N_19545,N_18043,N_18991);
xnor U19546 (N_19546,N_18850,N_18449);
xnor U19547 (N_19547,N_18781,N_18205);
nor U19548 (N_19548,N_18053,N_18093);
nand U19549 (N_19549,N_18504,N_18825);
xnor U19550 (N_19550,N_18422,N_18463);
nor U19551 (N_19551,N_18226,N_18995);
xor U19552 (N_19552,N_18873,N_18761);
and U19553 (N_19553,N_18866,N_18211);
nor U19554 (N_19554,N_18471,N_18161);
nor U19555 (N_19555,N_18113,N_18607);
and U19556 (N_19556,N_18512,N_18194);
nand U19557 (N_19557,N_18585,N_18390);
or U19558 (N_19558,N_18663,N_18276);
nand U19559 (N_19559,N_18617,N_18930);
nand U19560 (N_19560,N_18579,N_18924);
and U19561 (N_19561,N_18903,N_18681);
nand U19562 (N_19562,N_18796,N_18778);
xor U19563 (N_19563,N_18263,N_18757);
xor U19564 (N_19564,N_18683,N_18281);
or U19565 (N_19565,N_18347,N_18522);
or U19566 (N_19566,N_18330,N_18618);
nor U19567 (N_19567,N_18034,N_18589);
nor U19568 (N_19568,N_18481,N_18704);
or U19569 (N_19569,N_18203,N_18271);
nand U19570 (N_19570,N_18662,N_18384);
or U19571 (N_19571,N_18682,N_18730);
xnor U19572 (N_19572,N_18278,N_18903);
nand U19573 (N_19573,N_18473,N_18440);
nand U19574 (N_19574,N_18762,N_18530);
nor U19575 (N_19575,N_18595,N_18424);
nand U19576 (N_19576,N_18547,N_18851);
nor U19577 (N_19577,N_18838,N_18490);
nand U19578 (N_19578,N_18581,N_18742);
nor U19579 (N_19579,N_18976,N_18424);
nand U19580 (N_19580,N_18927,N_18440);
nand U19581 (N_19581,N_18189,N_18762);
nand U19582 (N_19582,N_18943,N_18924);
and U19583 (N_19583,N_18067,N_18136);
nand U19584 (N_19584,N_18929,N_18326);
nand U19585 (N_19585,N_18852,N_18702);
and U19586 (N_19586,N_18275,N_18232);
nand U19587 (N_19587,N_18469,N_18307);
and U19588 (N_19588,N_18116,N_18544);
xnor U19589 (N_19589,N_18918,N_18017);
and U19590 (N_19590,N_18442,N_18492);
or U19591 (N_19591,N_18601,N_18165);
nor U19592 (N_19592,N_18317,N_18075);
nor U19593 (N_19593,N_18824,N_18347);
or U19594 (N_19594,N_18911,N_18000);
nor U19595 (N_19595,N_18444,N_18579);
and U19596 (N_19596,N_18783,N_18958);
nand U19597 (N_19597,N_18251,N_18698);
nand U19598 (N_19598,N_18528,N_18809);
nand U19599 (N_19599,N_18164,N_18831);
and U19600 (N_19600,N_18008,N_18639);
nand U19601 (N_19601,N_18969,N_18132);
and U19602 (N_19602,N_18655,N_18205);
nand U19603 (N_19603,N_18102,N_18688);
nand U19604 (N_19604,N_18013,N_18887);
nor U19605 (N_19605,N_18337,N_18512);
xor U19606 (N_19606,N_18921,N_18666);
and U19607 (N_19607,N_18837,N_18486);
nor U19608 (N_19608,N_18275,N_18683);
nor U19609 (N_19609,N_18052,N_18213);
nor U19610 (N_19610,N_18341,N_18348);
xor U19611 (N_19611,N_18899,N_18077);
xor U19612 (N_19612,N_18129,N_18597);
nand U19613 (N_19613,N_18188,N_18627);
nor U19614 (N_19614,N_18911,N_18045);
or U19615 (N_19615,N_18822,N_18478);
nor U19616 (N_19616,N_18486,N_18421);
xnor U19617 (N_19617,N_18346,N_18264);
nand U19618 (N_19618,N_18593,N_18929);
or U19619 (N_19619,N_18113,N_18189);
nand U19620 (N_19620,N_18796,N_18668);
nand U19621 (N_19621,N_18925,N_18544);
or U19622 (N_19622,N_18143,N_18739);
nand U19623 (N_19623,N_18261,N_18644);
nor U19624 (N_19624,N_18392,N_18808);
nand U19625 (N_19625,N_18131,N_18214);
and U19626 (N_19626,N_18338,N_18315);
and U19627 (N_19627,N_18982,N_18307);
nand U19628 (N_19628,N_18430,N_18064);
nand U19629 (N_19629,N_18681,N_18649);
nor U19630 (N_19630,N_18300,N_18952);
or U19631 (N_19631,N_18102,N_18968);
and U19632 (N_19632,N_18567,N_18462);
xor U19633 (N_19633,N_18335,N_18924);
nor U19634 (N_19634,N_18333,N_18286);
xor U19635 (N_19635,N_18350,N_18637);
nand U19636 (N_19636,N_18240,N_18935);
and U19637 (N_19637,N_18860,N_18844);
and U19638 (N_19638,N_18001,N_18506);
or U19639 (N_19639,N_18874,N_18330);
or U19640 (N_19640,N_18070,N_18995);
xor U19641 (N_19641,N_18630,N_18059);
nor U19642 (N_19642,N_18186,N_18063);
or U19643 (N_19643,N_18561,N_18595);
xor U19644 (N_19644,N_18953,N_18509);
nand U19645 (N_19645,N_18296,N_18328);
or U19646 (N_19646,N_18442,N_18402);
xnor U19647 (N_19647,N_18108,N_18068);
xor U19648 (N_19648,N_18145,N_18619);
or U19649 (N_19649,N_18321,N_18988);
nor U19650 (N_19650,N_18305,N_18186);
xor U19651 (N_19651,N_18672,N_18147);
or U19652 (N_19652,N_18308,N_18289);
or U19653 (N_19653,N_18663,N_18414);
nor U19654 (N_19654,N_18893,N_18876);
xnor U19655 (N_19655,N_18477,N_18443);
nor U19656 (N_19656,N_18361,N_18651);
and U19657 (N_19657,N_18026,N_18815);
nand U19658 (N_19658,N_18314,N_18954);
xor U19659 (N_19659,N_18180,N_18051);
or U19660 (N_19660,N_18512,N_18422);
or U19661 (N_19661,N_18676,N_18642);
and U19662 (N_19662,N_18393,N_18840);
and U19663 (N_19663,N_18368,N_18780);
xor U19664 (N_19664,N_18665,N_18078);
or U19665 (N_19665,N_18376,N_18950);
nand U19666 (N_19666,N_18874,N_18479);
nand U19667 (N_19667,N_18971,N_18432);
nand U19668 (N_19668,N_18976,N_18672);
or U19669 (N_19669,N_18612,N_18139);
and U19670 (N_19670,N_18053,N_18602);
nor U19671 (N_19671,N_18085,N_18984);
and U19672 (N_19672,N_18540,N_18294);
nor U19673 (N_19673,N_18672,N_18522);
and U19674 (N_19674,N_18605,N_18079);
nand U19675 (N_19675,N_18663,N_18693);
nor U19676 (N_19676,N_18669,N_18283);
and U19677 (N_19677,N_18453,N_18029);
or U19678 (N_19678,N_18231,N_18730);
or U19679 (N_19679,N_18284,N_18865);
and U19680 (N_19680,N_18442,N_18166);
xor U19681 (N_19681,N_18550,N_18772);
xor U19682 (N_19682,N_18063,N_18743);
xnor U19683 (N_19683,N_18995,N_18728);
and U19684 (N_19684,N_18373,N_18619);
and U19685 (N_19685,N_18661,N_18419);
nor U19686 (N_19686,N_18462,N_18392);
and U19687 (N_19687,N_18843,N_18814);
nand U19688 (N_19688,N_18884,N_18266);
nor U19689 (N_19689,N_18069,N_18277);
or U19690 (N_19690,N_18478,N_18180);
nand U19691 (N_19691,N_18064,N_18393);
and U19692 (N_19692,N_18246,N_18780);
and U19693 (N_19693,N_18276,N_18656);
xor U19694 (N_19694,N_18278,N_18457);
nor U19695 (N_19695,N_18469,N_18039);
nor U19696 (N_19696,N_18778,N_18625);
nor U19697 (N_19697,N_18686,N_18258);
xor U19698 (N_19698,N_18176,N_18873);
or U19699 (N_19699,N_18486,N_18688);
nand U19700 (N_19700,N_18993,N_18220);
and U19701 (N_19701,N_18948,N_18282);
and U19702 (N_19702,N_18565,N_18444);
nand U19703 (N_19703,N_18644,N_18897);
nor U19704 (N_19704,N_18139,N_18185);
xnor U19705 (N_19705,N_18574,N_18431);
or U19706 (N_19706,N_18441,N_18169);
or U19707 (N_19707,N_18584,N_18535);
and U19708 (N_19708,N_18774,N_18416);
or U19709 (N_19709,N_18567,N_18928);
nor U19710 (N_19710,N_18003,N_18795);
and U19711 (N_19711,N_18080,N_18619);
and U19712 (N_19712,N_18786,N_18330);
and U19713 (N_19713,N_18649,N_18186);
and U19714 (N_19714,N_18474,N_18896);
and U19715 (N_19715,N_18029,N_18385);
xnor U19716 (N_19716,N_18735,N_18776);
nor U19717 (N_19717,N_18358,N_18258);
nand U19718 (N_19718,N_18531,N_18950);
xnor U19719 (N_19719,N_18742,N_18975);
nand U19720 (N_19720,N_18739,N_18723);
nand U19721 (N_19721,N_18337,N_18216);
nand U19722 (N_19722,N_18802,N_18222);
nor U19723 (N_19723,N_18433,N_18976);
xnor U19724 (N_19724,N_18066,N_18579);
and U19725 (N_19725,N_18224,N_18504);
nor U19726 (N_19726,N_18483,N_18270);
nand U19727 (N_19727,N_18360,N_18134);
and U19728 (N_19728,N_18168,N_18668);
xnor U19729 (N_19729,N_18933,N_18221);
xnor U19730 (N_19730,N_18639,N_18840);
and U19731 (N_19731,N_18609,N_18754);
nor U19732 (N_19732,N_18172,N_18885);
xnor U19733 (N_19733,N_18543,N_18712);
nor U19734 (N_19734,N_18042,N_18226);
nand U19735 (N_19735,N_18559,N_18715);
xor U19736 (N_19736,N_18506,N_18595);
or U19737 (N_19737,N_18153,N_18859);
nand U19738 (N_19738,N_18758,N_18425);
nor U19739 (N_19739,N_18624,N_18858);
or U19740 (N_19740,N_18896,N_18853);
nor U19741 (N_19741,N_18141,N_18216);
xor U19742 (N_19742,N_18580,N_18257);
nand U19743 (N_19743,N_18068,N_18927);
nand U19744 (N_19744,N_18350,N_18018);
nor U19745 (N_19745,N_18400,N_18901);
and U19746 (N_19746,N_18201,N_18657);
nor U19747 (N_19747,N_18189,N_18166);
and U19748 (N_19748,N_18805,N_18287);
nor U19749 (N_19749,N_18998,N_18843);
nand U19750 (N_19750,N_18717,N_18952);
nand U19751 (N_19751,N_18420,N_18438);
or U19752 (N_19752,N_18042,N_18583);
nor U19753 (N_19753,N_18584,N_18920);
and U19754 (N_19754,N_18981,N_18449);
or U19755 (N_19755,N_18381,N_18404);
nand U19756 (N_19756,N_18797,N_18078);
xnor U19757 (N_19757,N_18688,N_18572);
nor U19758 (N_19758,N_18392,N_18421);
nor U19759 (N_19759,N_18576,N_18552);
or U19760 (N_19760,N_18552,N_18177);
nand U19761 (N_19761,N_18121,N_18832);
nand U19762 (N_19762,N_18166,N_18462);
and U19763 (N_19763,N_18544,N_18370);
xor U19764 (N_19764,N_18539,N_18668);
and U19765 (N_19765,N_18270,N_18327);
xor U19766 (N_19766,N_18504,N_18188);
nor U19767 (N_19767,N_18193,N_18141);
nand U19768 (N_19768,N_18521,N_18680);
nand U19769 (N_19769,N_18915,N_18614);
nand U19770 (N_19770,N_18406,N_18533);
nand U19771 (N_19771,N_18124,N_18785);
and U19772 (N_19772,N_18920,N_18662);
and U19773 (N_19773,N_18732,N_18956);
or U19774 (N_19774,N_18836,N_18264);
xor U19775 (N_19775,N_18071,N_18859);
xnor U19776 (N_19776,N_18618,N_18371);
or U19777 (N_19777,N_18503,N_18064);
or U19778 (N_19778,N_18994,N_18267);
nor U19779 (N_19779,N_18027,N_18789);
nand U19780 (N_19780,N_18696,N_18063);
or U19781 (N_19781,N_18057,N_18893);
nand U19782 (N_19782,N_18438,N_18228);
or U19783 (N_19783,N_18353,N_18320);
nand U19784 (N_19784,N_18545,N_18886);
nand U19785 (N_19785,N_18574,N_18758);
nand U19786 (N_19786,N_18979,N_18831);
nand U19787 (N_19787,N_18627,N_18624);
or U19788 (N_19788,N_18657,N_18317);
or U19789 (N_19789,N_18242,N_18135);
xor U19790 (N_19790,N_18753,N_18920);
nor U19791 (N_19791,N_18565,N_18834);
or U19792 (N_19792,N_18434,N_18658);
xor U19793 (N_19793,N_18060,N_18159);
or U19794 (N_19794,N_18671,N_18749);
nand U19795 (N_19795,N_18752,N_18623);
nand U19796 (N_19796,N_18265,N_18529);
or U19797 (N_19797,N_18252,N_18311);
nor U19798 (N_19798,N_18077,N_18563);
or U19799 (N_19799,N_18399,N_18235);
or U19800 (N_19800,N_18255,N_18613);
nand U19801 (N_19801,N_18623,N_18848);
and U19802 (N_19802,N_18653,N_18599);
and U19803 (N_19803,N_18813,N_18773);
or U19804 (N_19804,N_18062,N_18966);
nand U19805 (N_19805,N_18464,N_18525);
nand U19806 (N_19806,N_18311,N_18805);
xnor U19807 (N_19807,N_18364,N_18543);
xnor U19808 (N_19808,N_18061,N_18519);
xor U19809 (N_19809,N_18095,N_18688);
and U19810 (N_19810,N_18396,N_18198);
and U19811 (N_19811,N_18062,N_18046);
or U19812 (N_19812,N_18372,N_18470);
nor U19813 (N_19813,N_18357,N_18219);
or U19814 (N_19814,N_18851,N_18361);
nor U19815 (N_19815,N_18689,N_18244);
nor U19816 (N_19816,N_18885,N_18677);
and U19817 (N_19817,N_18842,N_18178);
or U19818 (N_19818,N_18575,N_18915);
nand U19819 (N_19819,N_18085,N_18663);
and U19820 (N_19820,N_18066,N_18923);
xor U19821 (N_19821,N_18766,N_18393);
xnor U19822 (N_19822,N_18593,N_18845);
nand U19823 (N_19823,N_18864,N_18201);
and U19824 (N_19824,N_18492,N_18281);
or U19825 (N_19825,N_18151,N_18881);
nor U19826 (N_19826,N_18393,N_18912);
xnor U19827 (N_19827,N_18880,N_18571);
and U19828 (N_19828,N_18850,N_18147);
nand U19829 (N_19829,N_18187,N_18645);
or U19830 (N_19830,N_18505,N_18046);
nand U19831 (N_19831,N_18195,N_18247);
or U19832 (N_19832,N_18712,N_18282);
nor U19833 (N_19833,N_18183,N_18064);
nand U19834 (N_19834,N_18773,N_18635);
nor U19835 (N_19835,N_18395,N_18590);
nand U19836 (N_19836,N_18771,N_18183);
nand U19837 (N_19837,N_18542,N_18027);
or U19838 (N_19838,N_18098,N_18072);
or U19839 (N_19839,N_18196,N_18789);
xnor U19840 (N_19840,N_18613,N_18429);
nor U19841 (N_19841,N_18442,N_18620);
xor U19842 (N_19842,N_18668,N_18255);
nand U19843 (N_19843,N_18122,N_18023);
nor U19844 (N_19844,N_18725,N_18104);
nor U19845 (N_19845,N_18598,N_18156);
or U19846 (N_19846,N_18211,N_18280);
xnor U19847 (N_19847,N_18142,N_18517);
nor U19848 (N_19848,N_18211,N_18742);
xor U19849 (N_19849,N_18024,N_18631);
and U19850 (N_19850,N_18104,N_18176);
nand U19851 (N_19851,N_18607,N_18347);
and U19852 (N_19852,N_18311,N_18659);
nor U19853 (N_19853,N_18423,N_18966);
nand U19854 (N_19854,N_18709,N_18286);
nor U19855 (N_19855,N_18666,N_18820);
xor U19856 (N_19856,N_18131,N_18183);
or U19857 (N_19857,N_18470,N_18037);
nand U19858 (N_19858,N_18355,N_18586);
nor U19859 (N_19859,N_18550,N_18442);
and U19860 (N_19860,N_18955,N_18422);
or U19861 (N_19861,N_18461,N_18113);
xor U19862 (N_19862,N_18478,N_18576);
and U19863 (N_19863,N_18903,N_18937);
nor U19864 (N_19864,N_18442,N_18551);
and U19865 (N_19865,N_18212,N_18214);
nand U19866 (N_19866,N_18392,N_18929);
xnor U19867 (N_19867,N_18456,N_18286);
and U19868 (N_19868,N_18853,N_18089);
xor U19869 (N_19869,N_18334,N_18034);
or U19870 (N_19870,N_18687,N_18422);
xnor U19871 (N_19871,N_18409,N_18283);
and U19872 (N_19872,N_18334,N_18801);
nand U19873 (N_19873,N_18704,N_18399);
xor U19874 (N_19874,N_18979,N_18342);
nor U19875 (N_19875,N_18148,N_18479);
and U19876 (N_19876,N_18001,N_18527);
nor U19877 (N_19877,N_18177,N_18667);
xor U19878 (N_19878,N_18904,N_18876);
or U19879 (N_19879,N_18837,N_18034);
and U19880 (N_19880,N_18382,N_18797);
xnor U19881 (N_19881,N_18278,N_18272);
and U19882 (N_19882,N_18520,N_18243);
nor U19883 (N_19883,N_18882,N_18726);
and U19884 (N_19884,N_18789,N_18686);
nand U19885 (N_19885,N_18835,N_18435);
or U19886 (N_19886,N_18619,N_18315);
and U19887 (N_19887,N_18092,N_18343);
nor U19888 (N_19888,N_18657,N_18926);
nor U19889 (N_19889,N_18779,N_18427);
nand U19890 (N_19890,N_18401,N_18218);
or U19891 (N_19891,N_18027,N_18598);
or U19892 (N_19892,N_18831,N_18269);
and U19893 (N_19893,N_18320,N_18067);
nand U19894 (N_19894,N_18291,N_18024);
and U19895 (N_19895,N_18251,N_18156);
xor U19896 (N_19896,N_18737,N_18465);
nand U19897 (N_19897,N_18893,N_18353);
nor U19898 (N_19898,N_18328,N_18355);
nor U19899 (N_19899,N_18669,N_18738);
or U19900 (N_19900,N_18808,N_18164);
or U19901 (N_19901,N_18404,N_18891);
nor U19902 (N_19902,N_18618,N_18030);
nand U19903 (N_19903,N_18721,N_18023);
and U19904 (N_19904,N_18450,N_18303);
nand U19905 (N_19905,N_18917,N_18655);
and U19906 (N_19906,N_18954,N_18950);
nand U19907 (N_19907,N_18254,N_18976);
nor U19908 (N_19908,N_18439,N_18176);
or U19909 (N_19909,N_18723,N_18513);
or U19910 (N_19910,N_18708,N_18400);
or U19911 (N_19911,N_18149,N_18495);
and U19912 (N_19912,N_18023,N_18491);
xor U19913 (N_19913,N_18188,N_18186);
xor U19914 (N_19914,N_18602,N_18005);
nor U19915 (N_19915,N_18296,N_18503);
nand U19916 (N_19916,N_18795,N_18434);
xnor U19917 (N_19917,N_18556,N_18342);
nand U19918 (N_19918,N_18016,N_18991);
and U19919 (N_19919,N_18496,N_18593);
nor U19920 (N_19920,N_18414,N_18909);
nor U19921 (N_19921,N_18650,N_18817);
or U19922 (N_19922,N_18026,N_18611);
and U19923 (N_19923,N_18352,N_18118);
nor U19924 (N_19924,N_18697,N_18128);
and U19925 (N_19925,N_18492,N_18837);
nor U19926 (N_19926,N_18974,N_18163);
xor U19927 (N_19927,N_18865,N_18187);
and U19928 (N_19928,N_18170,N_18660);
or U19929 (N_19929,N_18242,N_18090);
and U19930 (N_19930,N_18675,N_18422);
nand U19931 (N_19931,N_18123,N_18561);
and U19932 (N_19932,N_18179,N_18777);
and U19933 (N_19933,N_18470,N_18108);
nor U19934 (N_19934,N_18238,N_18840);
nand U19935 (N_19935,N_18818,N_18505);
or U19936 (N_19936,N_18839,N_18814);
and U19937 (N_19937,N_18589,N_18544);
or U19938 (N_19938,N_18966,N_18079);
nand U19939 (N_19939,N_18606,N_18125);
or U19940 (N_19940,N_18548,N_18937);
xnor U19941 (N_19941,N_18303,N_18712);
xor U19942 (N_19942,N_18478,N_18854);
nor U19943 (N_19943,N_18801,N_18313);
xor U19944 (N_19944,N_18177,N_18897);
xnor U19945 (N_19945,N_18580,N_18673);
or U19946 (N_19946,N_18703,N_18635);
or U19947 (N_19947,N_18179,N_18849);
or U19948 (N_19948,N_18879,N_18157);
or U19949 (N_19949,N_18214,N_18690);
nand U19950 (N_19950,N_18476,N_18348);
xor U19951 (N_19951,N_18223,N_18747);
and U19952 (N_19952,N_18698,N_18036);
and U19953 (N_19953,N_18983,N_18334);
nand U19954 (N_19954,N_18136,N_18204);
xnor U19955 (N_19955,N_18759,N_18247);
xor U19956 (N_19956,N_18641,N_18537);
nand U19957 (N_19957,N_18548,N_18519);
nor U19958 (N_19958,N_18622,N_18613);
or U19959 (N_19959,N_18099,N_18239);
nand U19960 (N_19960,N_18098,N_18030);
nand U19961 (N_19961,N_18546,N_18303);
and U19962 (N_19962,N_18234,N_18323);
nor U19963 (N_19963,N_18732,N_18891);
nand U19964 (N_19964,N_18917,N_18170);
xnor U19965 (N_19965,N_18549,N_18093);
and U19966 (N_19966,N_18064,N_18040);
or U19967 (N_19967,N_18762,N_18234);
nor U19968 (N_19968,N_18746,N_18381);
nand U19969 (N_19969,N_18437,N_18149);
nand U19970 (N_19970,N_18499,N_18829);
nand U19971 (N_19971,N_18349,N_18625);
nor U19972 (N_19972,N_18656,N_18548);
nand U19973 (N_19973,N_18702,N_18742);
xnor U19974 (N_19974,N_18797,N_18824);
and U19975 (N_19975,N_18779,N_18503);
or U19976 (N_19976,N_18149,N_18612);
and U19977 (N_19977,N_18268,N_18876);
nand U19978 (N_19978,N_18806,N_18924);
nor U19979 (N_19979,N_18931,N_18248);
or U19980 (N_19980,N_18883,N_18576);
nand U19981 (N_19981,N_18167,N_18800);
nor U19982 (N_19982,N_18036,N_18506);
xor U19983 (N_19983,N_18522,N_18892);
or U19984 (N_19984,N_18176,N_18217);
or U19985 (N_19985,N_18892,N_18679);
nand U19986 (N_19986,N_18567,N_18210);
and U19987 (N_19987,N_18035,N_18769);
nor U19988 (N_19988,N_18923,N_18498);
and U19989 (N_19989,N_18700,N_18045);
xnor U19990 (N_19990,N_18894,N_18787);
xnor U19991 (N_19991,N_18209,N_18277);
nand U19992 (N_19992,N_18098,N_18961);
nor U19993 (N_19993,N_18144,N_18656);
xnor U19994 (N_19994,N_18813,N_18094);
xor U19995 (N_19995,N_18935,N_18457);
nand U19996 (N_19996,N_18945,N_18254);
or U19997 (N_19997,N_18860,N_18220);
or U19998 (N_19998,N_18537,N_18801);
xnor U19999 (N_19999,N_18293,N_18376);
or UO_0 (O_0,N_19023,N_19723);
and UO_1 (O_1,N_19059,N_19962);
nor UO_2 (O_2,N_19136,N_19538);
nor UO_3 (O_3,N_19809,N_19562);
nand UO_4 (O_4,N_19762,N_19260);
nand UO_5 (O_5,N_19544,N_19034);
nand UO_6 (O_6,N_19899,N_19098);
or UO_7 (O_7,N_19508,N_19579);
nor UO_8 (O_8,N_19408,N_19461);
or UO_9 (O_9,N_19469,N_19793);
nor UO_10 (O_10,N_19048,N_19534);
xnor UO_11 (O_11,N_19231,N_19772);
nor UO_12 (O_12,N_19557,N_19268);
nand UO_13 (O_13,N_19013,N_19889);
or UO_14 (O_14,N_19936,N_19853);
and UO_15 (O_15,N_19718,N_19797);
or UO_16 (O_16,N_19716,N_19810);
and UO_17 (O_17,N_19240,N_19632);
nor UO_18 (O_18,N_19886,N_19088);
nor UO_19 (O_19,N_19961,N_19942);
nand UO_20 (O_20,N_19804,N_19120);
xor UO_21 (O_21,N_19540,N_19873);
xnor UO_22 (O_22,N_19479,N_19841);
xor UO_23 (O_23,N_19280,N_19397);
and UO_24 (O_24,N_19801,N_19635);
nor UO_25 (O_25,N_19639,N_19426);
or UO_26 (O_26,N_19863,N_19791);
nand UO_27 (O_27,N_19262,N_19327);
xnor UO_28 (O_28,N_19456,N_19835);
or UO_29 (O_29,N_19702,N_19506);
nand UO_30 (O_30,N_19800,N_19432);
and UO_31 (O_31,N_19784,N_19173);
and UO_32 (O_32,N_19210,N_19149);
or UO_33 (O_33,N_19395,N_19293);
and UO_34 (O_34,N_19366,N_19451);
nand UO_35 (O_35,N_19085,N_19373);
xor UO_36 (O_36,N_19455,N_19228);
nor UO_37 (O_37,N_19255,N_19424);
and UO_38 (O_38,N_19980,N_19850);
nor UO_39 (O_39,N_19143,N_19565);
and UO_40 (O_40,N_19263,N_19539);
xor UO_41 (O_41,N_19106,N_19566);
xnor UO_42 (O_42,N_19200,N_19737);
or UO_43 (O_43,N_19514,N_19189);
nand UO_44 (O_44,N_19387,N_19249);
xor UO_45 (O_45,N_19065,N_19647);
xor UO_46 (O_46,N_19191,N_19711);
or UO_47 (O_47,N_19184,N_19125);
nand UO_48 (O_48,N_19206,N_19223);
or UO_49 (O_49,N_19049,N_19657);
or UO_50 (O_50,N_19473,N_19620);
and UO_51 (O_51,N_19522,N_19421);
nand UO_52 (O_52,N_19242,N_19156);
xor UO_53 (O_53,N_19821,N_19546);
xor UO_54 (O_54,N_19274,N_19478);
or UO_55 (O_55,N_19956,N_19217);
and UO_56 (O_56,N_19822,N_19337);
xor UO_57 (O_57,N_19795,N_19239);
or UO_58 (O_58,N_19827,N_19954);
nor UO_59 (O_59,N_19258,N_19484);
or UO_60 (O_60,N_19335,N_19693);
and UO_61 (O_61,N_19553,N_19887);
or UO_62 (O_62,N_19292,N_19178);
xor UO_63 (O_63,N_19837,N_19277);
xnor UO_64 (O_64,N_19081,N_19905);
or UO_65 (O_65,N_19398,N_19392);
xor UO_66 (O_66,N_19857,N_19053);
nor UO_67 (O_67,N_19133,N_19578);
xor UO_68 (O_68,N_19381,N_19113);
nor UO_69 (O_69,N_19589,N_19917);
nor UO_70 (O_70,N_19972,N_19749);
and UO_71 (O_71,N_19324,N_19529);
nand UO_72 (O_72,N_19952,N_19177);
xor UO_73 (O_73,N_19985,N_19115);
nor UO_74 (O_74,N_19743,N_19443);
xor UO_75 (O_75,N_19035,N_19636);
and UO_76 (O_76,N_19777,N_19535);
or UO_77 (O_77,N_19050,N_19384);
nand UO_78 (O_78,N_19330,N_19969);
xnor UO_79 (O_79,N_19163,N_19092);
nor UO_80 (O_80,N_19511,N_19660);
or UO_81 (O_81,N_19393,N_19353);
or UO_82 (O_82,N_19316,N_19041);
xor UO_83 (O_83,N_19714,N_19380);
nor UO_84 (O_84,N_19752,N_19666);
and UO_85 (O_85,N_19403,N_19089);
nor UO_86 (O_86,N_19364,N_19116);
nand UO_87 (O_87,N_19406,N_19493);
and UO_88 (O_88,N_19846,N_19076);
nor UO_89 (O_89,N_19569,N_19261);
or UO_90 (O_90,N_19164,N_19523);
xor UO_91 (O_91,N_19880,N_19336);
or UO_92 (O_92,N_19026,N_19998);
or UO_93 (O_93,N_19180,N_19778);
and UO_94 (O_94,N_19867,N_19269);
and UO_95 (O_95,N_19623,N_19814);
nand UO_96 (O_96,N_19874,N_19758);
nor UO_97 (O_97,N_19587,N_19742);
or UO_98 (O_98,N_19039,N_19012);
nand UO_99 (O_99,N_19607,N_19351);
and UO_100 (O_100,N_19297,N_19774);
or UO_101 (O_101,N_19645,N_19441);
or UO_102 (O_102,N_19400,N_19294);
xor UO_103 (O_103,N_19315,N_19314);
or UO_104 (O_104,N_19032,N_19947);
or UO_105 (O_105,N_19600,N_19829);
nand UO_106 (O_106,N_19188,N_19568);
or UO_107 (O_107,N_19573,N_19870);
or UO_108 (O_108,N_19134,N_19593);
and UO_109 (O_109,N_19219,N_19367);
or UO_110 (O_110,N_19649,N_19940);
and UO_111 (O_111,N_19344,N_19830);
nor UO_112 (O_112,N_19447,N_19572);
nor UO_113 (O_113,N_19900,N_19745);
xor UO_114 (O_114,N_19005,N_19927);
and UO_115 (O_115,N_19909,N_19014);
nand UO_116 (O_116,N_19211,N_19146);
and UO_117 (O_117,N_19064,N_19688);
and UO_118 (O_118,N_19295,N_19444);
or UO_119 (O_119,N_19348,N_19878);
nand UO_120 (O_120,N_19220,N_19779);
and UO_121 (O_121,N_19732,N_19665);
nand UO_122 (O_122,N_19983,N_19027);
or UO_123 (O_123,N_19320,N_19599);
and UO_124 (O_124,N_19279,N_19826);
xnor UO_125 (O_125,N_19613,N_19140);
nand UO_126 (O_126,N_19283,N_19057);
and UO_127 (O_127,N_19570,N_19077);
xnor UO_128 (O_128,N_19684,N_19914);
and UO_129 (O_129,N_19401,N_19243);
and UO_130 (O_130,N_19709,N_19806);
xnor UO_131 (O_131,N_19750,N_19273);
nor UO_132 (O_132,N_19360,N_19731);
and UO_133 (O_133,N_19706,N_19959);
nand UO_134 (O_134,N_19127,N_19250);
and UO_135 (O_135,N_19168,N_19021);
xor UO_136 (O_136,N_19734,N_19929);
and UO_137 (O_137,N_19984,N_19096);
xor UO_138 (O_138,N_19740,N_19641);
or UO_139 (O_139,N_19981,N_19072);
or UO_140 (O_140,N_19638,N_19298);
nor UO_141 (O_141,N_19198,N_19018);
nand UO_142 (O_142,N_19549,N_19042);
or UO_143 (O_143,N_19875,N_19640);
nand UO_144 (O_144,N_19241,N_19182);
nor UO_145 (O_145,N_19792,N_19884);
xor UO_146 (O_146,N_19307,N_19515);
and UO_147 (O_147,N_19513,N_19847);
nor UO_148 (O_148,N_19010,N_19996);
or UO_149 (O_149,N_19044,N_19661);
or UO_150 (O_150,N_19910,N_19414);
or UO_151 (O_151,N_19904,N_19434);
nor UO_152 (O_152,N_19347,N_19171);
nand UO_153 (O_153,N_19652,N_19111);
nand UO_154 (O_154,N_19449,N_19446);
nand UO_155 (O_155,N_19425,N_19525);
or UO_156 (O_156,N_19668,N_19248);
and UO_157 (O_157,N_19464,N_19063);
nand UO_158 (O_158,N_19375,N_19596);
nand UO_159 (O_159,N_19237,N_19119);
xor UO_160 (O_160,N_19533,N_19616);
nor UO_161 (O_161,N_19967,N_19585);
nand UO_162 (O_162,N_19350,N_19918);
nor UO_163 (O_163,N_19717,N_19396);
and UO_164 (O_164,N_19427,N_19062);
nor UO_165 (O_165,N_19973,N_19677);
xnor UO_166 (O_166,N_19445,N_19595);
xor UO_167 (O_167,N_19861,N_19453);
nor UO_168 (O_168,N_19654,N_19855);
xnor UO_169 (O_169,N_19704,N_19836);
nor UO_170 (O_170,N_19252,N_19517);
nor UO_171 (O_171,N_19915,N_19659);
nand UO_172 (O_172,N_19930,N_19378);
nor UO_173 (O_173,N_19524,N_19528);
and UO_174 (O_174,N_19169,N_19783);
xor UO_175 (O_175,N_19552,N_19377);
or UO_176 (O_176,N_19679,N_19877);
nand UO_177 (O_177,N_19839,N_19627);
or UO_178 (O_178,N_19142,N_19199);
or UO_179 (O_179,N_19055,N_19864);
or UO_180 (O_180,N_19158,N_19267);
and UO_181 (O_181,N_19520,N_19388);
or UO_182 (O_182,N_19457,N_19933);
and UO_183 (O_183,N_19003,N_19276);
and UO_184 (O_184,N_19270,N_19608);
and UO_185 (O_185,N_19022,N_19282);
and UO_186 (O_186,N_19467,N_19394);
xnor UO_187 (O_187,N_19082,N_19908);
nand UO_188 (O_188,N_19058,N_19201);
nand UO_189 (O_189,N_19968,N_19487);
nand UO_190 (O_190,N_19545,N_19083);
and UO_191 (O_191,N_19355,N_19037);
xor UO_192 (O_192,N_19687,N_19767);
nor UO_193 (O_193,N_19977,N_19409);
nor UO_194 (O_194,N_19953,N_19428);
nand UO_195 (O_195,N_19207,N_19695);
or UO_196 (O_196,N_19359,N_19819);
xnor UO_197 (O_197,N_19357,N_19193);
nor UO_198 (O_198,N_19713,N_19764);
xor UO_199 (O_199,N_19458,N_19747);
nor UO_200 (O_200,N_19680,N_19246);
or UO_201 (O_201,N_19681,N_19245);
and UO_202 (O_202,N_19785,N_19851);
nand UO_203 (O_203,N_19078,N_19112);
or UO_204 (O_204,N_19786,N_19871);
and UO_205 (O_205,N_19374,N_19489);
nor UO_206 (O_206,N_19233,N_19746);
nor UO_207 (O_207,N_19482,N_19937);
nor UO_208 (O_208,N_19526,N_19770);
and UO_209 (O_209,N_19564,N_19462);
nor UO_210 (O_210,N_19726,N_19454);
and UO_211 (O_211,N_19289,N_19868);
or UO_212 (O_212,N_19281,N_19581);
and UO_213 (O_213,N_19865,N_19622);
xor UO_214 (O_214,N_19707,N_19643);
and UO_215 (O_215,N_19235,N_19031);
and UO_216 (O_216,N_19893,N_19004);
and UO_217 (O_217,N_19744,N_19537);
xnor UO_218 (O_218,N_19015,N_19975);
nor UO_219 (O_219,N_19460,N_19730);
and UO_220 (O_220,N_19805,N_19033);
xor UO_221 (O_221,N_19610,N_19369);
nor UO_222 (O_222,N_19308,N_19556);
xor UO_223 (O_223,N_19071,N_19304);
xor UO_224 (O_224,N_19498,N_19637);
xor UO_225 (O_225,N_19187,N_19284);
and UO_226 (O_226,N_19019,N_19834);
and UO_227 (O_227,N_19820,N_19326);
and UO_228 (O_228,N_19329,N_19296);
xnor UO_229 (O_229,N_19046,N_19919);
xnor UO_230 (O_230,N_19601,N_19334);
nor UO_231 (O_231,N_19603,N_19025);
nand UO_232 (O_232,N_19621,N_19000);
xor UO_233 (O_233,N_19813,N_19222);
nand UO_234 (O_234,N_19594,N_19951);
xnor UO_235 (O_235,N_19766,N_19626);
nor UO_236 (O_236,N_19151,N_19694);
nor UO_237 (O_237,N_19002,N_19490);
nor UO_238 (O_238,N_19722,N_19205);
nor UO_239 (O_239,N_19856,N_19901);
nor UO_240 (O_240,N_19729,N_19322);
and UO_241 (O_241,N_19994,N_19036);
or UO_242 (O_242,N_19056,N_19885);
or UO_243 (O_243,N_19892,N_19943);
nand UO_244 (O_244,N_19488,N_19696);
xor UO_245 (O_245,N_19925,N_19509);
or UO_246 (O_246,N_19415,N_19780);
nand UO_247 (O_247,N_19903,N_19312);
nor UO_248 (O_248,N_19105,N_19087);
xor UO_249 (O_249,N_19093,N_19941);
nor UO_250 (O_250,N_19300,N_19618);
nor UO_251 (O_251,N_19674,N_19921);
nor UO_252 (O_252,N_19882,N_19765);
and UO_253 (O_253,N_19879,N_19038);
and UO_254 (O_254,N_19179,N_19160);
nand UO_255 (O_255,N_19876,N_19550);
nand UO_256 (O_256,N_19612,N_19831);
xor UO_257 (O_257,N_19362,N_19132);
xnor UO_258 (O_258,N_19130,N_19271);
nor UO_259 (O_259,N_19288,N_19107);
nor UO_260 (O_260,N_19802,N_19842);
xnor UO_261 (O_261,N_19964,N_19052);
nor UO_262 (O_262,N_19215,N_19794);
nor UO_263 (O_263,N_19928,N_19030);
nor UO_264 (O_264,N_19759,N_19577);
nand UO_265 (O_265,N_19960,N_19605);
and UO_266 (O_266,N_19790,N_19218);
and UO_267 (O_267,N_19185,N_19976);
or UO_268 (O_268,N_19463,N_19672);
xor UO_269 (O_269,N_19333,N_19939);
xor UO_270 (O_270,N_19376,N_19971);
or UO_271 (O_271,N_19580,N_19024);
xnor UO_272 (O_272,N_19824,N_19371);
nand UO_273 (O_273,N_19117,N_19989);
or UO_274 (O_274,N_19776,N_19771);
nand UO_275 (O_275,N_19020,N_19485);
or UO_276 (O_276,N_19705,N_19094);
nor UO_277 (O_277,N_19299,N_19633);
and UO_278 (O_278,N_19405,N_19150);
nand UO_279 (O_279,N_19195,N_19328);
or UO_280 (O_280,N_19208,N_19266);
xor UO_281 (O_281,N_19472,N_19650);
nor UO_282 (O_282,N_19194,N_19789);
and UO_283 (O_283,N_19285,N_19631);
or UO_284 (O_284,N_19979,N_19710);
and UO_285 (O_285,N_19763,N_19340);
nand UO_286 (O_286,N_19606,N_19306);
nand UO_287 (O_287,N_19817,N_19675);
nor UO_288 (O_288,N_19029,N_19074);
nand UO_289 (O_289,N_19435,N_19017);
xnor UO_290 (O_290,N_19574,N_19502);
and UO_291 (O_291,N_19591,N_19685);
nand UO_292 (O_292,N_19181,N_19399);
and UO_293 (O_293,N_19137,N_19229);
and UO_294 (O_294,N_19898,N_19363);
or UO_295 (O_295,N_19437,N_19097);
xnor UO_296 (O_296,N_19413,N_19175);
nor UO_297 (O_297,N_19828,N_19391);
and UO_298 (O_298,N_19440,N_19341);
or UO_299 (O_299,N_19738,N_19450);
and UO_300 (O_300,N_19844,N_19497);
or UO_301 (O_301,N_19833,N_19686);
nor UO_302 (O_302,N_19412,N_19128);
or UO_303 (O_303,N_19407,N_19518);
xor UO_304 (O_304,N_19495,N_19236);
nor UO_305 (O_305,N_19754,N_19547);
nor UO_306 (O_306,N_19852,N_19588);
xor UO_307 (O_307,N_19110,N_19895);
or UO_308 (O_308,N_19416,N_19070);
nor UO_309 (O_309,N_19075,N_19721);
nor UO_310 (O_310,N_19310,N_19386);
nor UO_311 (O_311,N_19530,N_19510);
nand UO_312 (O_312,N_19987,N_19658);
nor UO_313 (O_313,N_19719,N_19238);
nand UO_314 (O_314,N_19624,N_19992);
nor UO_315 (O_315,N_19512,N_19247);
xor UO_316 (O_316,N_19614,N_19272);
or UO_317 (O_317,N_19896,N_19483);
nor UO_318 (O_318,N_19803,N_19216);
nand UO_319 (O_319,N_19167,N_19257);
xnor UO_320 (O_320,N_19061,N_19339);
nand UO_321 (O_321,N_19318,N_19812);
nand UO_322 (O_322,N_19683,N_19760);
nand UO_323 (O_323,N_19183,N_19016);
nor UO_324 (O_324,N_19286,N_19091);
xnor UO_325 (O_325,N_19576,N_19028);
nand UO_326 (O_326,N_19197,N_19291);
nand UO_327 (O_327,N_19225,N_19007);
and UO_328 (O_328,N_19644,N_19551);
and UO_329 (O_329,N_19008,N_19648);
xor UO_330 (O_330,N_19869,N_19689);
nor UO_331 (O_331,N_19773,N_19741);
nand UO_332 (O_332,N_19265,N_19491);
nand UO_333 (O_333,N_19370,N_19358);
and UO_334 (O_334,N_19101,N_19838);
or UO_335 (O_335,N_19651,N_19698);
or UO_336 (O_336,N_19720,N_19253);
nor UO_337 (O_337,N_19438,N_19958);
or UO_338 (O_338,N_19906,N_19597);
and UO_339 (O_339,N_19911,N_19418);
or UO_340 (O_340,N_19410,N_19054);
or UO_341 (O_341,N_19978,N_19808);
nor UO_342 (O_342,N_19753,N_19963);
nand UO_343 (O_343,N_19990,N_19554);
or UO_344 (O_344,N_19368,N_19100);
nor UO_345 (O_345,N_19678,N_19944);
or UO_346 (O_346,N_19047,N_19126);
xnor UO_347 (O_347,N_19949,N_19474);
or UO_348 (O_348,N_19902,N_19172);
nand UO_349 (O_349,N_19932,N_19991);
nor UO_350 (O_350,N_19476,N_19433);
or UO_351 (O_351,N_19419,N_19924);
or UO_352 (O_352,N_19615,N_19848);
or UO_353 (O_353,N_19372,N_19586);
xnor UO_354 (O_354,N_19313,N_19145);
nand UO_355 (O_355,N_19221,N_19667);
nor UO_356 (O_356,N_19516,N_19118);
nor UO_357 (O_357,N_19768,N_19417);
nand UO_358 (O_358,N_19192,N_19646);
and UO_359 (O_359,N_19155,N_19148);
and UO_360 (O_360,N_19468,N_19302);
nand UO_361 (O_361,N_19931,N_19420);
or UO_362 (O_362,N_19798,N_19935);
nor UO_363 (O_363,N_19832,N_19402);
xnor UO_364 (O_364,N_19583,N_19602);
nand UO_365 (O_365,N_19494,N_19811);
or UO_366 (O_366,N_19575,N_19109);
and UO_367 (O_367,N_19673,N_19664);
and UO_368 (O_368,N_19244,N_19214);
xor UO_369 (O_369,N_19883,N_19733);
or UO_370 (O_370,N_19466,N_19825);
or UO_371 (O_371,N_19881,N_19114);
nand UO_372 (O_372,N_19701,N_19060);
nand UO_373 (O_373,N_19890,N_19095);
xor UO_374 (O_374,N_19170,N_19669);
nand UO_375 (O_375,N_19736,N_19655);
xnor UO_376 (O_376,N_19332,N_19986);
or UO_377 (O_377,N_19558,N_19066);
and UO_378 (O_378,N_19823,N_19213);
nor UO_379 (O_379,N_19354,N_19582);
or UO_380 (O_380,N_19727,N_19356);
nand UO_381 (O_381,N_19957,N_19390);
and UO_382 (O_382,N_19152,N_19411);
nor UO_383 (O_383,N_19922,N_19423);
and UO_384 (O_384,N_19287,N_19571);
or UO_385 (O_385,N_19712,N_19051);
nand UO_386 (O_386,N_19703,N_19159);
and UO_387 (O_387,N_19739,N_19227);
or UO_388 (O_388,N_19129,N_19611);
nor UO_389 (O_389,N_19692,N_19431);
or UO_390 (O_390,N_19212,N_19141);
nor UO_391 (O_391,N_19619,N_19226);
and UO_392 (O_392,N_19629,N_19452);
nand UO_393 (O_393,N_19290,N_19080);
or UO_394 (O_394,N_19548,N_19559);
nor UO_395 (O_395,N_19365,N_19135);
and UO_396 (O_396,N_19757,N_19592);
nand UO_397 (O_397,N_19671,N_19389);
or UO_398 (O_398,N_19543,N_19162);
and UO_399 (O_399,N_19124,N_19787);
and UO_400 (O_400,N_19174,N_19521);
or UO_401 (O_401,N_19816,N_19563);
xnor UO_402 (O_402,N_19974,N_19190);
nand UO_403 (O_403,N_19256,N_19946);
xor UO_404 (O_404,N_19011,N_19796);
nand UO_405 (O_405,N_19788,N_19642);
or UO_406 (O_406,N_19090,N_19323);
xor UO_407 (O_407,N_19486,N_19319);
nand UO_408 (O_408,N_19099,N_19699);
nor UO_409 (O_409,N_19436,N_19154);
nand UO_410 (O_410,N_19519,N_19379);
xnor UO_411 (O_411,N_19496,N_19532);
or UO_412 (O_412,N_19209,N_19492);
or UO_413 (O_413,N_19383,N_19912);
nor UO_414 (O_414,N_19001,N_19907);
xor UO_415 (O_415,N_19799,N_19843);
or UO_416 (O_416,N_19858,N_19309);
or UO_417 (O_417,N_19866,N_19480);
nand UO_418 (O_418,N_19009,N_19305);
xor UO_419 (O_419,N_19501,N_19232);
and UO_420 (O_420,N_19934,N_19735);
nor UO_421 (O_421,N_19815,N_19104);
or UO_422 (O_422,N_19555,N_19338);
xor UO_423 (O_423,N_19872,N_19429);
nand UO_424 (O_424,N_19470,N_19203);
or UO_425 (O_425,N_19728,N_19604);
and UO_426 (O_426,N_19849,N_19897);
xor UO_427 (O_427,N_19691,N_19948);
nor UO_428 (O_428,N_19542,N_19345);
nor UO_429 (O_429,N_19234,N_19067);
nor UO_430 (O_430,N_19663,N_19708);
or UO_431 (O_431,N_19700,N_19782);
xor UO_432 (O_432,N_19186,N_19751);
or UO_433 (O_433,N_19311,N_19769);
or UO_434 (O_434,N_19430,N_19131);
and UO_435 (O_435,N_19923,N_19157);
and UO_436 (O_436,N_19475,N_19818);
nor UO_437 (O_437,N_19916,N_19724);
or UO_438 (O_438,N_19196,N_19043);
nand UO_439 (O_439,N_19471,N_19690);
and UO_440 (O_440,N_19807,N_19697);
nand UO_441 (O_441,N_19560,N_19598);
nor UO_442 (O_442,N_19006,N_19982);
nand UO_443 (O_443,N_19301,N_19422);
and UO_444 (O_444,N_19781,N_19630);
and UO_445 (O_445,N_19259,N_19404);
xnor UO_446 (O_446,N_19503,N_19541);
nand UO_447 (O_447,N_19343,N_19166);
and UO_448 (O_448,N_19346,N_19845);
nor UO_449 (O_449,N_19955,N_19670);
or UO_450 (O_450,N_19913,N_19352);
xor UO_451 (O_451,N_19993,N_19504);
and UO_452 (O_452,N_19349,N_19122);
and UO_453 (O_453,N_19465,N_19755);
or UO_454 (O_454,N_19995,N_19086);
and UO_455 (O_455,N_19303,N_19628);
nand UO_456 (O_456,N_19123,N_19481);
xnor UO_457 (O_457,N_19859,N_19945);
and UO_458 (O_458,N_19331,N_19361);
and UO_459 (O_459,N_19342,N_19584);
nand UO_460 (O_460,N_19715,N_19448);
nand UO_461 (O_461,N_19138,N_19775);
nor UO_462 (O_462,N_19988,N_19121);
xnor UO_463 (O_463,N_19108,N_19144);
or UO_464 (O_464,N_19997,N_19891);
nand UO_465 (O_465,N_19966,N_19153);
and UO_466 (O_466,N_19068,N_19860);
xor UO_467 (O_467,N_19325,N_19165);
and UO_468 (O_468,N_19748,N_19970);
nand UO_469 (O_469,N_19254,N_19317);
xnor UO_470 (O_470,N_19999,N_19888);
nor UO_471 (O_471,N_19204,N_19477);
nand UO_472 (O_472,N_19567,N_19536);
xnor UO_473 (O_473,N_19862,N_19499);
xnor UO_474 (O_474,N_19069,N_19590);
xor UO_475 (O_475,N_19459,N_19264);
nand UO_476 (O_476,N_19625,N_19894);
or UO_477 (O_477,N_19531,N_19617);
nand UO_478 (O_478,N_19382,N_19176);
or UO_479 (O_479,N_19224,N_19926);
and UO_480 (O_480,N_19965,N_19500);
nand UO_481 (O_481,N_19102,N_19938);
nor UO_482 (O_482,N_19161,N_19725);
xor UO_483 (O_483,N_19662,N_19442);
or UO_484 (O_484,N_19653,N_19854);
and UO_485 (O_485,N_19656,N_19079);
and UO_486 (O_486,N_19439,N_19147);
nand UO_487 (O_487,N_19634,N_19676);
and UO_488 (O_488,N_19385,N_19321);
or UO_489 (O_489,N_19609,N_19761);
nor UO_490 (O_490,N_19251,N_19505);
xor UO_491 (O_491,N_19202,N_19920);
nor UO_492 (O_492,N_19073,N_19756);
nand UO_493 (O_493,N_19040,N_19275);
xor UO_494 (O_494,N_19084,N_19045);
or UO_495 (O_495,N_19950,N_19139);
xor UO_496 (O_496,N_19507,N_19230);
nor UO_497 (O_497,N_19561,N_19278);
or UO_498 (O_498,N_19840,N_19682);
nor UO_499 (O_499,N_19103,N_19527);
nor UO_500 (O_500,N_19225,N_19932);
and UO_501 (O_501,N_19629,N_19841);
nand UO_502 (O_502,N_19484,N_19502);
nor UO_503 (O_503,N_19461,N_19044);
nand UO_504 (O_504,N_19850,N_19394);
and UO_505 (O_505,N_19569,N_19373);
nor UO_506 (O_506,N_19296,N_19607);
and UO_507 (O_507,N_19414,N_19280);
and UO_508 (O_508,N_19040,N_19644);
xor UO_509 (O_509,N_19083,N_19322);
and UO_510 (O_510,N_19930,N_19366);
nor UO_511 (O_511,N_19703,N_19016);
and UO_512 (O_512,N_19290,N_19407);
nand UO_513 (O_513,N_19025,N_19680);
or UO_514 (O_514,N_19532,N_19801);
nand UO_515 (O_515,N_19288,N_19577);
and UO_516 (O_516,N_19320,N_19143);
nor UO_517 (O_517,N_19753,N_19778);
nor UO_518 (O_518,N_19906,N_19393);
xor UO_519 (O_519,N_19903,N_19688);
xnor UO_520 (O_520,N_19019,N_19633);
or UO_521 (O_521,N_19625,N_19764);
and UO_522 (O_522,N_19425,N_19715);
nor UO_523 (O_523,N_19240,N_19401);
nor UO_524 (O_524,N_19509,N_19620);
and UO_525 (O_525,N_19541,N_19646);
and UO_526 (O_526,N_19606,N_19339);
and UO_527 (O_527,N_19450,N_19778);
xnor UO_528 (O_528,N_19612,N_19053);
nor UO_529 (O_529,N_19058,N_19944);
and UO_530 (O_530,N_19276,N_19102);
nor UO_531 (O_531,N_19035,N_19657);
or UO_532 (O_532,N_19870,N_19198);
nand UO_533 (O_533,N_19843,N_19023);
xor UO_534 (O_534,N_19195,N_19019);
nand UO_535 (O_535,N_19623,N_19688);
and UO_536 (O_536,N_19762,N_19030);
or UO_537 (O_537,N_19387,N_19748);
xnor UO_538 (O_538,N_19575,N_19053);
nand UO_539 (O_539,N_19534,N_19320);
nand UO_540 (O_540,N_19303,N_19495);
nor UO_541 (O_541,N_19602,N_19063);
nand UO_542 (O_542,N_19908,N_19431);
nand UO_543 (O_543,N_19299,N_19859);
nor UO_544 (O_544,N_19702,N_19541);
and UO_545 (O_545,N_19363,N_19000);
nor UO_546 (O_546,N_19519,N_19783);
and UO_547 (O_547,N_19821,N_19848);
or UO_548 (O_548,N_19826,N_19801);
and UO_549 (O_549,N_19439,N_19565);
or UO_550 (O_550,N_19328,N_19253);
and UO_551 (O_551,N_19701,N_19486);
or UO_552 (O_552,N_19609,N_19285);
nor UO_553 (O_553,N_19688,N_19102);
nand UO_554 (O_554,N_19178,N_19884);
nor UO_555 (O_555,N_19700,N_19482);
nor UO_556 (O_556,N_19908,N_19129);
nor UO_557 (O_557,N_19894,N_19731);
nor UO_558 (O_558,N_19350,N_19959);
or UO_559 (O_559,N_19945,N_19896);
and UO_560 (O_560,N_19960,N_19673);
or UO_561 (O_561,N_19491,N_19653);
nor UO_562 (O_562,N_19689,N_19498);
and UO_563 (O_563,N_19068,N_19273);
nand UO_564 (O_564,N_19832,N_19594);
xor UO_565 (O_565,N_19382,N_19342);
xnor UO_566 (O_566,N_19156,N_19438);
xor UO_567 (O_567,N_19987,N_19553);
nand UO_568 (O_568,N_19280,N_19141);
nand UO_569 (O_569,N_19485,N_19627);
nand UO_570 (O_570,N_19918,N_19131);
nand UO_571 (O_571,N_19160,N_19682);
and UO_572 (O_572,N_19760,N_19955);
nand UO_573 (O_573,N_19149,N_19970);
and UO_574 (O_574,N_19275,N_19313);
nor UO_575 (O_575,N_19640,N_19769);
or UO_576 (O_576,N_19133,N_19587);
nor UO_577 (O_577,N_19100,N_19439);
nand UO_578 (O_578,N_19733,N_19020);
nand UO_579 (O_579,N_19661,N_19524);
nand UO_580 (O_580,N_19692,N_19358);
and UO_581 (O_581,N_19805,N_19089);
nand UO_582 (O_582,N_19333,N_19961);
xnor UO_583 (O_583,N_19791,N_19387);
or UO_584 (O_584,N_19173,N_19171);
nor UO_585 (O_585,N_19239,N_19326);
and UO_586 (O_586,N_19076,N_19789);
or UO_587 (O_587,N_19221,N_19760);
nand UO_588 (O_588,N_19637,N_19393);
and UO_589 (O_589,N_19605,N_19096);
nor UO_590 (O_590,N_19412,N_19798);
nor UO_591 (O_591,N_19714,N_19327);
nor UO_592 (O_592,N_19494,N_19576);
and UO_593 (O_593,N_19036,N_19061);
and UO_594 (O_594,N_19124,N_19683);
and UO_595 (O_595,N_19207,N_19527);
nand UO_596 (O_596,N_19936,N_19569);
xnor UO_597 (O_597,N_19484,N_19494);
and UO_598 (O_598,N_19253,N_19186);
or UO_599 (O_599,N_19526,N_19352);
nand UO_600 (O_600,N_19499,N_19917);
nand UO_601 (O_601,N_19245,N_19019);
nor UO_602 (O_602,N_19132,N_19514);
nand UO_603 (O_603,N_19108,N_19486);
nor UO_604 (O_604,N_19447,N_19642);
or UO_605 (O_605,N_19976,N_19262);
or UO_606 (O_606,N_19991,N_19305);
nor UO_607 (O_607,N_19379,N_19357);
nor UO_608 (O_608,N_19976,N_19975);
nor UO_609 (O_609,N_19016,N_19518);
and UO_610 (O_610,N_19308,N_19092);
xnor UO_611 (O_611,N_19012,N_19865);
xnor UO_612 (O_612,N_19629,N_19648);
nor UO_613 (O_613,N_19867,N_19653);
nand UO_614 (O_614,N_19840,N_19400);
and UO_615 (O_615,N_19676,N_19349);
nand UO_616 (O_616,N_19652,N_19964);
or UO_617 (O_617,N_19687,N_19676);
nand UO_618 (O_618,N_19424,N_19019);
or UO_619 (O_619,N_19842,N_19297);
nand UO_620 (O_620,N_19236,N_19209);
xor UO_621 (O_621,N_19409,N_19050);
nor UO_622 (O_622,N_19097,N_19757);
xnor UO_623 (O_623,N_19089,N_19572);
nor UO_624 (O_624,N_19912,N_19601);
and UO_625 (O_625,N_19939,N_19549);
and UO_626 (O_626,N_19838,N_19481);
and UO_627 (O_627,N_19017,N_19784);
and UO_628 (O_628,N_19775,N_19906);
xor UO_629 (O_629,N_19011,N_19914);
or UO_630 (O_630,N_19767,N_19707);
nand UO_631 (O_631,N_19753,N_19459);
xnor UO_632 (O_632,N_19832,N_19250);
and UO_633 (O_633,N_19634,N_19503);
nand UO_634 (O_634,N_19568,N_19499);
or UO_635 (O_635,N_19457,N_19017);
nor UO_636 (O_636,N_19559,N_19188);
nand UO_637 (O_637,N_19458,N_19822);
nor UO_638 (O_638,N_19944,N_19689);
nor UO_639 (O_639,N_19082,N_19952);
xnor UO_640 (O_640,N_19596,N_19240);
or UO_641 (O_641,N_19302,N_19989);
nand UO_642 (O_642,N_19229,N_19472);
xor UO_643 (O_643,N_19518,N_19373);
or UO_644 (O_644,N_19394,N_19137);
and UO_645 (O_645,N_19690,N_19803);
nand UO_646 (O_646,N_19161,N_19364);
nand UO_647 (O_647,N_19248,N_19030);
xnor UO_648 (O_648,N_19994,N_19069);
and UO_649 (O_649,N_19942,N_19432);
xor UO_650 (O_650,N_19379,N_19925);
nor UO_651 (O_651,N_19424,N_19794);
and UO_652 (O_652,N_19680,N_19931);
and UO_653 (O_653,N_19151,N_19224);
xor UO_654 (O_654,N_19049,N_19549);
nor UO_655 (O_655,N_19699,N_19994);
or UO_656 (O_656,N_19905,N_19764);
and UO_657 (O_657,N_19310,N_19922);
and UO_658 (O_658,N_19897,N_19816);
or UO_659 (O_659,N_19458,N_19487);
and UO_660 (O_660,N_19859,N_19501);
nor UO_661 (O_661,N_19875,N_19334);
nor UO_662 (O_662,N_19415,N_19524);
xor UO_663 (O_663,N_19887,N_19042);
or UO_664 (O_664,N_19775,N_19763);
or UO_665 (O_665,N_19436,N_19711);
and UO_666 (O_666,N_19872,N_19861);
and UO_667 (O_667,N_19292,N_19216);
nor UO_668 (O_668,N_19928,N_19104);
nor UO_669 (O_669,N_19143,N_19025);
or UO_670 (O_670,N_19492,N_19440);
or UO_671 (O_671,N_19520,N_19157);
nand UO_672 (O_672,N_19231,N_19140);
or UO_673 (O_673,N_19871,N_19104);
and UO_674 (O_674,N_19380,N_19152);
or UO_675 (O_675,N_19192,N_19027);
nor UO_676 (O_676,N_19265,N_19413);
nand UO_677 (O_677,N_19390,N_19447);
nand UO_678 (O_678,N_19338,N_19992);
or UO_679 (O_679,N_19557,N_19244);
or UO_680 (O_680,N_19813,N_19511);
nor UO_681 (O_681,N_19835,N_19863);
and UO_682 (O_682,N_19523,N_19034);
and UO_683 (O_683,N_19313,N_19069);
nor UO_684 (O_684,N_19393,N_19686);
nand UO_685 (O_685,N_19470,N_19337);
nand UO_686 (O_686,N_19368,N_19130);
xor UO_687 (O_687,N_19209,N_19980);
nand UO_688 (O_688,N_19119,N_19123);
nor UO_689 (O_689,N_19455,N_19919);
or UO_690 (O_690,N_19022,N_19444);
or UO_691 (O_691,N_19925,N_19762);
nor UO_692 (O_692,N_19721,N_19437);
xor UO_693 (O_693,N_19143,N_19698);
nor UO_694 (O_694,N_19635,N_19088);
xor UO_695 (O_695,N_19512,N_19744);
nand UO_696 (O_696,N_19531,N_19935);
xnor UO_697 (O_697,N_19828,N_19423);
nand UO_698 (O_698,N_19818,N_19078);
nor UO_699 (O_699,N_19584,N_19158);
nor UO_700 (O_700,N_19831,N_19489);
xor UO_701 (O_701,N_19057,N_19105);
xnor UO_702 (O_702,N_19011,N_19674);
nor UO_703 (O_703,N_19092,N_19150);
and UO_704 (O_704,N_19128,N_19029);
nor UO_705 (O_705,N_19020,N_19711);
nand UO_706 (O_706,N_19409,N_19119);
and UO_707 (O_707,N_19906,N_19412);
and UO_708 (O_708,N_19076,N_19324);
and UO_709 (O_709,N_19565,N_19616);
xnor UO_710 (O_710,N_19107,N_19095);
and UO_711 (O_711,N_19968,N_19129);
nand UO_712 (O_712,N_19431,N_19521);
or UO_713 (O_713,N_19512,N_19403);
and UO_714 (O_714,N_19868,N_19695);
nand UO_715 (O_715,N_19434,N_19014);
nor UO_716 (O_716,N_19180,N_19418);
nor UO_717 (O_717,N_19351,N_19591);
nor UO_718 (O_718,N_19706,N_19526);
xor UO_719 (O_719,N_19762,N_19891);
xnor UO_720 (O_720,N_19261,N_19881);
nor UO_721 (O_721,N_19301,N_19839);
nand UO_722 (O_722,N_19089,N_19188);
and UO_723 (O_723,N_19545,N_19219);
or UO_724 (O_724,N_19159,N_19670);
nand UO_725 (O_725,N_19221,N_19240);
nand UO_726 (O_726,N_19377,N_19948);
and UO_727 (O_727,N_19906,N_19466);
nand UO_728 (O_728,N_19978,N_19488);
nor UO_729 (O_729,N_19042,N_19102);
nor UO_730 (O_730,N_19320,N_19008);
nor UO_731 (O_731,N_19451,N_19420);
and UO_732 (O_732,N_19884,N_19819);
xnor UO_733 (O_733,N_19260,N_19854);
nor UO_734 (O_734,N_19300,N_19301);
or UO_735 (O_735,N_19355,N_19767);
nor UO_736 (O_736,N_19444,N_19973);
or UO_737 (O_737,N_19523,N_19230);
nand UO_738 (O_738,N_19094,N_19100);
or UO_739 (O_739,N_19161,N_19994);
xor UO_740 (O_740,N_19714,N_19468);
or UO_741 (O_741,N_19789,N_19445);
xor UO_742 (O_742,N_19990,N_19159);
or UO_743 (O_743,N_19802,N_19265);
nand UO_744 (O_744,N_19148,N_19590);
xnor UO_745 (O_745,N_19679,N_19124);
xor UO_746 (O_746,N_19442,N_19834);
nand UO_747 (O_747,N_19381,N_19755);
nand UO_748 (O_748,N_19286,N_19567);
xor UO_749 (O_749,N_19461,N_19956);
nand UO_750 (O_750,N_19666,N_19866);
and UO_751 (O_751,N_19238,N_19099);
xnor UO_752 (O_752,N_19963,N_19413);
nand UO_753 (O_753,N_19249,N_19833);
nand UO_754 (O_754,N_19088,N_19247);
and UO_755 (O_755,N_19318,N_19006);
or UO_756 (O_756,N_19026,N_19834);
nand UO_757 (O_757,N_19892,N_19241);
or UO_758 (O_758,N_19794,N_19327);
xnor UO_759 (O_759,N_19412,N_19604);
or UO_760 (O_760,N_19374,N_19473);
nor UO_761 (O_761,N_19274,N_19869);
or UO_762 (O_762,N_19215,N_19424);
xor UO_763 (O_763,N_19071,N_19022);
or UO_764 (O_764,N_19505,N_19824);
xor UO_765 (O_765,N_19789,N_19803);
or UO_766 (O_766,N_19883,N_19933);
xor UO_767 (O_767,N_19188,N_19283);
and UO_768 (O_768,N_19651,N_19058);
or UO_769 (O_769,N_19412,N_19706);
or UO_770 (O_770,N_19883,N_19034);
nand UO_771 (O_771,N_19939,N_19235);
nand UO_772 (O_772,N_19203,N_19448);
and UO_773 (O_773,N_19682,N_19301);
nand UO_774 (O_774,N_19631,N_19932);
xor UO_775 (O_775,N_19964,N_19612);
nand UO_776 (O_776,N_19981,N_19717);
nor UO_777 (O_777,N_19254,N_19120);
nand UO_778 (O_778,N_19827,N_19431);
nor UO_779 (O_779,N_19707,N_19741);
or UO_780 (O_780,N_19957,N_19659);
xnor UO_781 (O_781,N_19556,N_19390);
xor UO_782 (O_782,N_19897,N_19109);
or UO_783 (O_783,N_19182,N_19210);
and UO_784 (O_784,N_19692,N_19618);
xor UO_785 (O_785,N_19369,N_19750);
nor UO_786 (O_786,N_19429,N_19220);
or UO_787 (O_787,N_19972,N_19727);
xnor UO_788 (O_788,N_19586,N_19885);
xor UO_789 (O_789,N_19975,N_19559);
xnor UO_790 (O_790,N_19120,N_19072);
xnor UO_791 (O_791,N_19597,N_19568);
xor UO_792 (O_792,N_19393,N_19379);
and UO_793 (O_793,N_19383,N_19036);
or UO_794 (O_794,N_19174,N_19526);
or UO_795 (O_795,N_19846,N_19823);
and UO_796 (O_796,N_19609,N_19834);
and UO_797 (O_797,N_19545,N_19890);
xor UO_798 (O_798,N_19188,N_19354);
and UO_799 (O_799,N_19209,N_19315);
or UO_800 (O_800,N_19188,N_19183);
and UO_801 (O_801,N_19998,N_19390);
nand UO_802 (O_802,N_19369,N_19000);
nand UO_803 (O_803,N_19324,N_19668);
nand UO_804 (O_804,N_19486,N_19995);
or UO_805 (O_805,N_19096,N_19272);
and UO_806 (O_806,N_19033,N_19947);
xnor UO_807 (O_807,N_19673,N_19696);
xor UO_808 (O_808,N_19439,N_19715);
nand UO_809 (O_809,N_19891,N_19741);
xnor UO_810 (O_810,N_19622,N_19889);
or UO_811 (O_811,N_19596,N_19842);
xor UO_812 (O_812,N_19322,N_19721);
xnor UO_813 (O_813,N_19876,N_19152);
xnor UO_814 (O_814,N_19369,N_19777);
and UO_815 (O_815,N_19998,N_19286);
nor UO_816 (O_816,N_19584,N_19894);
nand UO_817 (O_817,N_19663,N_19255);
nor UO_818 (O_818,N_19578,N_19901);
or UO_819 (O_819,N_19504,N_19195);
nand UO_820 (O_820,N_19370,N_19555);
xor UO_821 (O_821,N_19112,N_19075);
and UO_822 (O_822,N_19433,N_19377);
or UO_823 (O_823,N_19798,N_19253);
xnor UO_824 (O_824,N_19612,N_19401);
xnor UO_825 (O_825,N_19766,N_19038);
and UO_826 (O_826,N_19399,N_19972);
nor UO_827 (O_827,N_19089,N_19960);
xnor UO_828 (O_828,N_19315,N_19217);
and UO_829 (O_829,N_19389,N_19962);
nor UO_830 (O_830,N_19243,N_19589);
xor UO_831 (O_831,N_19049,N_19516);
and UO_832 (O_832,N_19698,N_19968);
or UO_833 (O_833,N_19908,N_19269);
or UO_834 (O_834,N_19695,N_19398);
nor UO_835 (O_835,N_19428,N_19559);
or UO_836 (O_836,N_19202,N_19052);
xnor UO_837 (O_837,N_19450,N_19795);
xor UO_838 (O_838,N_19213,N_19469);
xor UO_839 (O_839,N_19085,N_19750);
xor UO_840 (O_840,N_19130,N_19789);
or UO_841 (O_841,N_19743,N_19406);
and UO_842 (O_842,N_19475,N_19743);
or UO_843 (O_843,N_19929,N_19702);
nand UO_844 (O_844,N_19245,N_19350);
or UO_845 (O_845,N_19609,N_19832);
nor UO_846 (O_846,N_19646,N_19585);
xor UO_847 (O_847,N_19237,N_19220);
xor UO_848 (O_848,N_19584,N_19544);
nor UO_849 (O_849,N_19006,N_19507);
xor UO_850 (O_850,N_19438,N_19787);
nor UO_851 (O_851,N_19783,N_19288);
nand UO_852 (O_852,N_19963,N_19285);
or UO_853 (O_853,N_19711,N_19586);
nor UO_854 (O_854,N_19641,N_19119);
xnor UO_855 (O_855,N_19948,N_19680);
xor UO_856 (O_856,N_19906,N_19237);
or UO_857 (O_857,N_19027,N_19222);
or UO_858 (O_858,N_19092,N_19107);
nand UO_859 (O_859,N_19490,N_19634);
nor UO_860 (O_860,N_19808,N_19190);
and UO_861 (O_861,N_19064,N_19352);
xor UO_862 (O_862,N_19566,N_19358);
and UO_863 (O_863,N_19438,N_19120);
nor UO_864 (O_864,N_19849,N_19367);
nor UO_865 (O_865,N_19154,N_19329);
or UO_866 (O_866,N_19774,N_19650);
nor UO_867 (O_867,N_19215,N_19691);
nor UO_868 (O_868,N_19603,N_19276);
or UO_869 (O_869,N_19590,N_19825);
nand UO_870 (O_870,N_19436,N_19560);
or UO_871 (O_871,N_19690,N_19900);
xnor UO_872 (O_872,N_19030,N_19894);
and UO_873 (O_873,N_19138,N_19607);
nor UO_874 (O_874,N_19940,N_19389);
nand UO_875 (O_875,N_19101,N_19356);
and UO_876 (O_876,N_19694,N_19290);
nor UO_877 (O_877,N_19382,N_19495);
xnor UO_878 (O_878,N_19773,N_19985);
and UO_879 (O_879,N_19602,N_19256);
xnor UO_880 (O_880,N_19495,N_19951);
and UO_881 (O_881,N_19565,N_19614);
or UO_882 (O_882,N_19491,N_19012);
nand UO_883 (O_883,N_19340,N_19769);
xnor UO_884 (O_884,N_19659,N_19159);
or UO_885 (O_885,N_19035,N_19876);
nor UO_886 (O_886,N_19667,N_19808);
xnor UO_887 (O_887,N_19855,N_19540);
or UO_888 (O_888,N_19039,N_19454);
nor UO_889 (O_889,N_19507,N_19968);
and UO_890 (O_890,N_19096,N_19337);
nand UO_891 (O_891,N_19437,N_19239);
nor UO_892 (O_892,N_19688,N_19139);
and UO_893 (O_893,N_19020,N_19264);
nand UO_894 (O_894,N_19615,N_19910);
nor UO_895 (O_895,N_19050,N_19666);
xnor UO_896 (O_896,N_19099,N_19083);
nor UO_897 (O_897,N_19839,N_19577);
nand UO_898 (O_898,N_19122,N_19543);
xnor UO_899 (O_899,N_19320,N_19102);
nor UO_900 (O_900,N_19899,N_19532);
or UO_901 (O_901,N_19168,N_19733);
and UO_902 (O_902,N_19843,N_19826);
or UO_903 (O_903,N_19299,N_19596);
xor UO_904 (O_904,N_19062,N_19747);
nand UO_905 (O_905,N_19392,N_19619);
nand UO_906 (O_906,N_19701,N_19580);
or UO_907 (O_907,N_19164,N_19558);
xnor UO_908 (O_908,N_19998,N_19107);
nor UO_909 (O_909,N_19095,N_19795);
and UO_910 (O_910,N_19834,N_19001);
xor UO_911 (O_911,N_19574,N_19816);
and UO_912 (O_912,N_19896,N_19116);
and UO_913 (O_913,N_19403,N_19870);
nand UO_914 (O_914,N_19360,N_19596);
nand UO_915 (O_915,N_19276,N_19420);
nand UO_916 (O_916,N_19743,N_19971);
and UO_917 (O_917,N_19271,N_19320);
or UO_918 (O_918,N_19248,N_19762);
nand UO_919 (O_919,N_19001,N_19630);
nor UO_920 (O_920,N_19592,N_19242);
or UO_921 (O_921,N_19272,N_19645);
or UO_922 (O_922,N_19362,N_19149);
nand UO_923 (O_923,N_19606,N_19298);
and UO_924 (O_924,N_19153,N_19049);
nor UO_925 (O_925,N_19012,N_19613);
nor UO_926 (O_926,N_19818,N_19721);
or UO_927 (O_927,N_19642,N_19653);
nor UO_928 (O_928,N_19022,N_19666);
xnor UO_929 (O_929,N_19777,N_19663);
or UO_930 (O_930,N_19756,N_19398);
and UO_931 (O_931,N_19656,N_19928);
and UO_932 (O_932,N_19971,N_19753);
and UO_933 (O_933,N_19618,N_19534);
and UO_934 (O_934,N_19664,N_19864);
nand UO_935 (O_935,N_19742,N_19376);
nand UO_936 (O_936,N_19297,N_19379);
or UO_937 (O_937,N_19989,N_19428);
nor UO_938 (O_938,N_19079,N_19350);
and UO_939 (O_939,N_19858,N_19011);
nand UO_940 (O_940,N_19871,N_19469);
nor UO_941 (O_941,N_19677,N_19239);
xnor UO_942 (O_942,N_19045,N_19724);
xnor UO_943 (O_943,N_19845,N_19624);
and UO_944 (O_944,N_19655,N_19615);
xor UO_945 (O_945,N_19277,N_19251);
nand UO_946 (O_946,N_19006,N_19589);
and UO_947 (O_947,N_19517,N_19989);
xnor UO_948 (O_948,N_19150,N_19984);
nand UO_949 (O_949,N_19907,N_19582);
or UO_950 (O_950,N_19834,N_19067);
or UO_951 (O_951,N_19408,N_19175);
nor UO_952 (O_952,N_19661,N_19225);
nand UO_953 (O_953,N_19447,N_19972);
nor UO_954 (O_954,N_19492,N_19651);
and UO_955 (O_955,N_19463,N_19996);
nand UO_956 (O_956,N_19777,N_19928);
nor UO_957 (O_957,N_19240,N_19912);
or UO_958 (O_958,N_19922,N_19847);
nand UO_959 (O_959,N_19063,N_19696);
xor UO_960 (O_960,N_19459,N_19187);
nor UO_961 (O_961,N_19193,N_19239);
xnor UO_962 (O_962,N_19407,N_19499);
nor UO_963 (O_963,N_19500,N_19936);
xor UO_964 (O_964,N_19505,N_19551);
nand UO_965 (O_965,N_19647,N_19795);
and UO_966 (O_966,N_19322,N_19554);
and UO_967 (O_967,N_19101,N_19430);
and UO_968 (O_968,N_19820,N_19877);
xor UO_969 (O_969,N_19124,N_19974);
and UO_970 (O_970,N_19824,N_19329);
or UO_971 (O_971,N_19360,N_19876);
or UO_972 (O_972,N_19692,N_19323);
nand UO_973 (O_973,N_19649,N_19066);
nand UO_974 (O_974,N_19423,N_19386);
xor UO_975 (O_975,N_19060,N_19552);
and UO_976 (O_976,N_19629,N_19347);
nand UO_977 (O_977,N_19019,N_19998);
nor UO_978 (O_978,N_19803,N_19292);
xor UO_979 (O_979,N_19146,N_19956);
and UO_980 (O_980,N_19356,N_19654);
xnor UO_981 (O_981,N_19460,N_19546);
nor UO_982 (O_982,N_19187,N_19028);
nand UO_983 (O_983,N_19255,N_19123);
nor UO_984 (O_984,N_19444,N_19680);
nor UO_985 (O_985,N_19904,N_19793);
nor UO_986 (O_986,N_19825,N_19546);
nand UO_987 (O_987,N_19975,N_19749);
and UO_988 (O_988,N_19054,N_19768);
or UO_989 (O_989,N_19009,N_19337);
and UO_990 (O_990,N_19913,N_19119);
and UO_991 (O_991,N_19258,N_19186);
nand UO_992 (O_992,N_19498,N_19291);
nand UO_993 (O_993,N_19268,N_19427);
and UO_994 (O_994,N_19764,N_19951);
and UO_995 (O_995,N_19645,N_19400);
nand UO_996 (O_996,N_19283,N_19579);
and UO_997 (O_997,N_19738,N_19001);
nand UO_998 (O_998,N_19047,N_19706);
xnor UO_999 (O_999,N_19781,N_19703);
xor UO_1000 (O_1000,N_19064,N_19119);
nor UO_1001 (O_1001,N_19935,N_19092);
nor UO_1002 (O_1002,N_19072,N_19269);
xor UO_1003 (O_1003,N_19348,N_19224);
or UO_1004 (O_1004,N_19708,N_19392);
xnor UO_1005 (O_1005,N_19033,N_19811);
xnor UO_1006 (O_1006,N_19153,N_19037);
and UO_1007 (O_1007,N_19016,N_19326);
xor UO_1008 (O_1008,N_19360,N_19619);
or UO_1009 (O_1009,N_19514,N_19055);
or UO_1010 (O_1010,N_19271,N_19038);
and UO_1011 (O_1011,N_19486,N_19530);
nor UO_1012 (O_1012,N_19457,N_19692);
nand UO_1013 (O_1013,N_19409,N_19438);
and UO_1014 (O_1014,N_19746,N_19061);
or UO_1015 (O_1015,N_19780,N_19146);
nand UO_1016 (O_1016,N_19955,N_19211);
or UO_1017 (O_1017,N_19120,N_19919);
nor UO_1018 (O_1018,N_19021,N_19663);
or UO_1019 (O_1019,N_19402,N_19129);
and UO_1020 (O_1020,N_19884,N_19465);
and UO_1021 (O_1021,N_19710,N_19921);
nand UO_1022 (O_1022,N_19358,N_19590);
and UO_1023 (O_1023,N_19192,N_19554);
nand UO_1024 (O_1024,N_19927,N_19685);
and UO_1025 (O_1025,N_19547,N_19088);
xnor UO_1026 (O_1026,N_19344,N_19847);
and UO_1027 (O_1027,N_19420,N_19467);
nand UO_1028 (O_1028,N_19572,N_19183);
or UO_1029 (O_1029,N_19600,N_19157);
nor UO_1030 (O_1030,N_19553,N_19050);
nor UO_1031 (O_1031,N_19225,N_19192);
and UO_1032 (O_1032,N_19505,N_19982);
nor UO_1033 (O_1033,N_19883,N_19908);
nand UO_1034 (O_1034,N_19137,N_19438);
nor UO_1035 (O_1035,N_19507,N_19379);
nand UO_1036 (O_1036,N_19696,N_19315);
nor UO_1037 (O_1037,N_19412,N_19664);
xnor UO_1038 (O_1038,N_19415,N_19352);
and UO_1039 (O_1039,N_19320,N_19754);
nand UO_1040 (O_1040,N_19265,N_19730);
and UO_1041 (O_1041,N_19625,N_19390);
and UO_1042 (O_1042,N_19003,N_19682);
nor UO_1043 (O_1043,N_19118,N_19426);
nor UO_1044 (O_1044,N_19209,N_19707);
nand UO_1045 (O_1045,N_19793,N_19262);
nand UO_1046 (O_1046,N_19206,N_19582);
or UO_1047 (O_1047,N_19265,N_19941);
and UO_1048 (O_1048,N_19346,N_19801);
nor UO_1049 (O_1049,N_19238,N_19373);
or UO_1050 (O_1050,N_19158,N_19048);
nand UO_1051 (O_1051,N_19048,N_19876);
and UO_1052 (O_1052,N_19656,N_19410);
nor UO_1053 (O_1053,N_19070,N_19715);
nor UO_1054 (O_1054,N_19788,N_19345);
nor UO_1055 (O_1055,N_19647,N_19270);
and UO_1056 (O_1056,N_19712,N_19726);
or UO_1057 (O_1057,N_19647,N_19452);
nand UO_1058 (O_1058,N_19558,N_19754);
and UO_1059 (O_1059,N_19736,N_19321);
and UO_1060 (O_1060,N_19854,N_19440);
and UO_1061 (O_1061,N_19537,N_19791);
xnor UO_1062 (O_1062,N_19791,N_19219);
xor UO_1063 (O_1063,N_19283,N_19808);
and UO_1064 (O_1064,N_19186,N_19350);
nand UO_1065 (O_1065,N_19580,N_19546);
and UO_1066 (O_1066,N_19152,N_19197);
or UO_1067 (O_1067,N_19568,N_19506);
and UO_1068 (O_1068,N_19723,N_19059);
xnor UO_1069 (O_1069,N_19259,N_19724);
nand UO_1070 (O_1070,N_19825,N_19929);
nor UO_1071 (O_1071,N_19467,N_19339);
nand UO_1072 (O_1072,N_19798,N_19942);
nand UO_1073 (O_1073,N_19017,N_19781);
and UO_1074 (O_1074,N_19156,N_19044);
xor UO_1075 (O_1075,N_19784,N_19362);
nor UO_1076 (O_1076,N_19733,N_19299);
nand UO_1077 (O_1077,N_19041,N_19949);
and UO_1078 (O_1078,N_19226,N_19184);
nor UO_1079 (O_1079,N_19164,N_19329);
nor UO_1080 (O_1080,N_19512,N_19486);
or UO_1081 (O_1081,N_19884,N_19694);
or UO_1082 (O_1082,N_19935,N_19683);
nand UO_1083 (O_1083,N_19529,N_19071);
nor UO_1084 (O_1084,N_19750,N_19541);
and UO_1085 (O_1085,N_19910,N_19285);
nor UO_1086 (O_1086,N_19113,N_19138);
nor UO_1087 (O_1087,N_19312,N_19022);
and UO_1088 (O_1088,N_19523,N_19394);
nor UO_1089 (O_1089,N_19418,N_19469);
and UO_1090 (O_1090,N_19133,N_19385);
or UO_1091 (O_1091,N_19468,N_19970);
xnor UO_1092 (O_1092,N_19302,N_19120);
and UO_1093 (O_1093,N_19747,N_19602);
and UO_1094 (O_1094,N_19311,N_19778);
nor UO_1095 (O_1095,N_19962,N_19517);
and UO_1096 (O_1096,N_19724,N_19177);
xnor UO_1097 (O_1097,N_19691,N_19098);
nor UO_1098 (O_1098,N_19423,N_19715);
nor UO_1099 (O_1099,N_19497,N_19639);
xnor UO_1100 (O_1100,N_19148,N_19143);
and UO_1101 (O_1101,N_19634,N_19550);
nor UO_1102 (O_1102,N_19521,N_19802);
xnor UO_1103 (O_1103,N_19704,N_19327);
and UO_1104 (O_1104,N_19276,N_19351);
xnor UO_1105 (O_1105,N_19954,N_19285);
nand UO_1106 (O_1106,N_19072,N_19844);
nor UO_1107 (O_1107,N_19926,N_19640);
and UO_1108 (O_1108,N_19828,N_19780);
nor UO_1109 (O_1109,N_19221,N_19401);
xor UO_1110 (O_1110,N_19638,N_19356);
nor UO_1111 (O_1111,N_19826,N_19479);
and UO_1112 (O_1112,N_19667,N_19204);
nor UO_1113 (O_1113,N_19878,N_19975);
and UO_1114 (O_1114,N_19938,N_19578);
nor UO_1115 (O_1115,N_19053,N_19978);
xnor UO_1116 (O_1116,N_19608,N_19884);
or UO_1117 (O_1117,N_19118,N_19555);
or UO_1118 (O_1118,N_19584,N_19715);
nand UO_1119 (O_1119,N_19488,N_19841);
nand UO_1120 (O_1120,N_19278,N_19316);
or UO_1121 (O_1121,N_19567,N_19115);
nand UO_1122 (O_1122,N_19778,N_19714);
or UO_1123 (O_1123,N_19541,N_19061);
nor UO_1124 (O_1124,N_19259,N_19231);
or UO_1125 (O_1125,N_19391,N_19741);
and UO_1126 (O_1126,N_19381,N_19416);
nand UO_1127 (O_1127,N_19068,N_19459);
nand UO_1128 (O_1128,N_19863,N_19473);
nand UO_1129 (O_1129,N_19492,N_19281);
xnor UO_1130 (O_1130,N_19259,N_19954);
nor UO_1131 (O_1131,N_19807,N_19248);
or UO_1132 (O_1132,N_19849,N_19611);
or UO_1133 (O_1133,N_19824,N_19459);
nand UO_1134 (O_1134,N_19016,N_19319);
or UO_1135 (O_1135,N_19664,N_19584);
nand UO_1136 (O_1136,N_19327,N_19776);
or UO_1137 (O_1137,N_19781,N_19100);
or UO_1138 (O_1138,N_19177,N_19020);
and UO_1139 (O_1139,N_19359,N_19303);
nand UO_1140 (O_1140,N_19018,N_19187);
or UO_1141 (O_1141,N_19506,N_19491);
nor UO_1142 (O_1142,N_19540,N_19486);
xnor UO_1143 (O_1143,N_19790,N_19516);
or UO_1144 (O_1144,N_19147,N_19405);
nand UO_1145 (O_1145,N_19970,N_19929);
and UO_1146 (O_1146,N_19861,N_19716);
nor UO_1147 (O_1147,N_19229,N_19982);
nand UO_1148 (O_1148,N_19088,N_19180);
nand UO_1149 (O_1149,N_19002,N_19559);
and UO_1150 (O_1150,N_19819,N_19521);
nand UO_1151 (O_1151,N_19971,N_19290);
nand UO_1152 (O_1152,N_19109,N_19881);
xor UO_1153 (O_1153,N_19382,N_19726);
and UO_1154 (O_1154,N_19042,N_19883);
nand UO_1155 (O_1155,N_19687,N_19754);
and UO_1156 (O_1156,N_19812,N_19246);
nor UO_1157 (O_1157,N_19249,N_19282);
or UO_1158 (O_1158,N_19333,N_19297);
and UO_1159 (O_1159,N_19502,N_19893);
or UO_1160 (O_1160,N_19360,N_19385);
nor UO_1161 (O_1161,N_19201,N_19295);
xor UO_1162 (O_1162,N_19230,N_19447);
nor UO_1163 (O_1163,N_19882,N_19080);
xor UO_1164 (O_1164,N_19836,N_19567);
nand UO_1165 (O_1165,N_19656,N_19245);
nor UO_1166 (O_1166,N_19967,N_19076);
or UO_1167 (O_1167,N_19919,N_19110);
or UO_1168 (O_1168,N_19913,N_19110);
nand UO_1169 (O_1169,N_19992,N_19846);
nand UO_1170 (O_1170,N_19838,N_19158);
xor UO_1171 (O_1171,N_19721,N_19941);
and UO_1172 (O_1172,N_19363,N_19657);
nor UO_1173 (O_1173,N_19525,N_19980);
or UO_1174 (O_1174,N_19828,N_19829);
xnor UO_1175 (O_1175,N_19721,N_19517);
xor UO_1176 (O_1176,N_19731,N_19405);
or UO_1177 (O_1177,N_19864,N_19847);
nand UO_1178 (O_1178,N_19714,N_19538);
nor UO_1179 (O_1179,N_19714,N_19165);
nand UO_1180 (O_1180,N_19894,N_19127);
or UO_1181 (O_1181,N_19825,N_19857);
and UO_1182 (O_1182,N_19151,N_19143);
xnor UO_1183 (O_1183,N_19714,N_19073);
xor UO_1184 (O_1184,N_19205,N_19582);
xnor UO_1185 (O_1185,N_19694,N_19396);
and UO_1186 (O_1186,N_19318,N_19200);
nor UO_1187 (O_1187,N_19259,N_19618);
and UO_1188 (O_1188,N_19284,N_19126);
xnor UO_1189 (O_1189,N_19442,N_19757);
nor UO_1190 (O_1190,N_19501,N_19235);
xor UO_1191 (O_1191,N_19503,N_19065);
xnor UO_1192 (O_1192,N_19099,N_19887);
nor UO_1193 (O_1193,N_19147,N_19800);
or UO_1194 (O_1194,N_19799,N_19086);
and UO_1195 (O_1195,N_19786,N_19904);
xnor UO_1196 (O_1196,N_19260,N_19123);
and UO_1197 (O_1197,N_19556,N_19140);
or UO_1198 (O_1198,N_19751,N_19531);
xor UO_1199 (O_1199,N_19441,N_19205);
xor UO_1200 (O_1200,N_19570,N_19503);
nand UO_1201 (O_1201,N_19247,N_19019);
nand UO_1202 (O_1202,N_19285,N_19982);
nand UO_1203 (O_1203,N_19569,N_19424);
nand UO_1204 (O_1204,N_19708,N_19885);
and UO_1205 (O_1205,N_19728,N_19036);
nand UO_1206 (O_1206,N_19703,N_19561);
nor UO_1207 (O_1207,N_19662,N_19776);
or UO_1208 (O_1208,N_19333,N_19184);
nor UO_1209 (O_1209,N_19084,N_19898);
and UO_1210 (O_1210,N_19238,N_19513);
nor UO_1211 (O_1211,N_19906,N_19204);
xor UO_1212 (O_1212,N_19629,N_19977);
nor UO_1213 (O_1213,N_19013,N_19637);
or UO_1214 (O_1214,N_19026,N_19762);
and UO_1215 (O_1215,N_19887,N_19272);
or UO_1216 (O_1216,N_19360,N_19981);
xor UO_1217 (O_1217,N_19966,N_19148);
nor UO_1218 (O_1218,N_19813,N_19344);
or UO_1219 (O_1219,N_19090,N_19452);
nand UO_1220 (O_1220,N_19229,N_19233);
and UO_1221 (O_1221,N_19451,N_19244);
nand UO_1222 (O_1222,N_19782,N_19836);
and UO_1223 (O_1223,N_19600,N_19437);
nand UO_1224 (O_1224,N_19674,N_19266);
xnor UO_1225 (O_1225,N_19013,N_19039);
nand UO_1226 (O_1226,N_19963,N_19209);
and UO_1227 (O_1227,N_19875,N_19624);
nor UO_1228 (O_1228,N_19581,N_19900);
or UO_1229 (O_1229,N_19701,N_19951);
xnor UO_1230 (O_1230,N_19772,N_19943);
nor UO_1231 (O_1231,N_19462,N_19248);
xor UO_1232 (O_1232,N_19294,N_19050);
nor UO_1233 (O_1233,N_19178,N_19785);
nor UO_1234 (O_1234,N_19776,N_19230);
nor UO_1235 (O_1235,N_19072,N_19265);
nand UO_1236 (O_1236,N_19419,N_19333);
xor UO_1237 (O_1237,N_19874,N_19985);
xor UO_1238 (O_1238,N_19374,N_19387);
nand UO_1239 (O_1239,N_19361,N_19073);
nor UO_1240 (O_1240,N_19622,N_19037);
xnor UO_1241 (O_1241,N_19339,N_19978);
xnor UO_1242 (O_1242,N_19838,N_19999);
xor UO_1243 (O_1243,N_19000,N_19231);
nor UO_1244 (O_1244,N_19213,N_19061);
and UO_1245 (O_1245,N_19147,N_19046);
nand UO_1246 (O_1246,N_19636,N_19509);
xnor UO_1247 (O_1247,N_19587,N_19031);
nor UO_1248 (O_1248,N_19446,N_19974);
or UO_1249 (O_1249,N_19606,N_19194);
or UO_1250 (O_1250,N_19094,N_19408);
nor UO_1251 (O_1251,N_19130,N_19125);
and UO_1252 (O_1252,N_19275,N_19813);
and UO_1253 (O_1253,N_19048,N_19783);
or UO_1254 (O_1254,N_19603,N_19330);
and UO_1255 (O_1255,N_19307,N_19398);
xnor UO_1256 (O_1256,N_19478,N_19861);
nand UO_1257 (O_1257,N_19832,N_19128);
nor UO_1258 (O_1258,N_19183,N_19074);
and UO_1259 (O_1259,N_19246,N_19872);
nor UO_1260 (O_1260,N_19375,N_19311);
nand UO_1261 (O_1261,N_19194,N_19528);
nor UO_1262 (O_1262,N_19489,N_19928);
xnor UO_1263 (O_1263,N_19720,N_19579);
nand UO_1264 (O_1264,N_19816,N_19860);
nand UO_1265 (O_1265,N_19918,N_19276);
and UO_1266 (O_1266,N_19291,N_19413);
xnor UO_1267 (O_1267,N_19815,N_19313);
or UO_1268 (O_1268,N_19970,N_19853);
nor UO_1269 (O_1269,N_19266,N_19668);
xor UO_1270 (O_1270,N_19132,N_19946);
nor UO_1271 (O_1271,N_19518,N_19000);
xnor UO_1272 (O_1272,N_19994,N_19341);
nand UO_1273 (O_1273,N_19657,N_19295);
xnor UO_1274 (O_1274,N_19127,N_19096);
xor UO_1275 (O_1275,N_19323,N_19836);
or UO_1276 (O_1276,N_19178,N_19522);
or UO_1277 (O_1277,N_19552,N_19097);
or UO_1278 (O_1278,N_19181,N_19426);
nor UO_1279 (O_1279,N_19469,N_19318);
nor UO_1280 (O_1280,N_19179,N_19718);
nor UO_1281 (O_1281,N_19462,N_19512);
xnor UO_1282 (O_1282,N_19767,N_19799);
nand UO_1283 (O_1283,N_19755,N_19271);
or UO_1284 (O_1284,N_19133,N_19559);
nand UO_1285 (O_1285,N_19743,N_19499);
and UO_1286 (O_1286,N_19322,N_19158);
nor UO_1287 (O_1287,N_19681,N_19968);
xnor UO_1288 (O_1288,N_19857,N_19787);
and UO_1289 (O_1289,N_19279,N_19889);
and UO_1290 (O_1290,N_19242,N_19998);
or UO_1291 (O_1291,N_19131,N_19042);
nand UO_1292 (O_1292,N_19437,N_19874);
xor UO_1293 (O_1293,N_19499,N_19044);
nand UO_1294 (O_1294,N_19898,N_19995);
nand UO_1295 (O_1295,N_19426,N_19513);
xnor UO_1296 (O_1296,N_19613,N_19338);
xor UO_1297 (O_1297,N_19560,N_19246);
nor UO_1298 (O_1298,N_19918,N_19578);
nand UO_1299 (O_1299,N_19869,N_19402);
or UO_1300 (O_1300,N_19118,N_19976);
and UO_1301 (O_1301,N_19993,N_19359);
xor UO_1302 (O_1302,N_19369,N_19088);
nand UO_1303 (O_1303,N_19790,N_19490);
xor UO_1304 (O_1304,N_19413,N_19690);
or UO_1305 (O_1305,N_19970,N_19992);
nand UO_1306 (O_1306,N_19042,N_19267);
nor UO_1307 (O_1307,N_19712,N_19985);
xor UO_1308 (O_1308,N_19936,N_19741);
or UO_1309 (O_1309,N_19219,N_19520);
and UO_1310 (O_1310,N_19101,N_19591);
xor UO_1311 (O_1311,N_19233,N_19935);
nand UO_1312 (O_1312,N_19388,N_19110);
nor UO_1313 (O_1313,N_19243,N_19453);
xnor UO_1314 (O_1314,N_19461,N_19347);
nor UO_1315 (O_1315,N_19559,N_19278);
nand UO_1316 (O_1316,N_19033,N_19698);
xnor UO_1317 (O_1317,N_19258,N_19009);
nor UO_1318 (O_1318,N_19192,N_19937);
nor UO_1319 (O_1319,N_19723,N_19586);
nor UO_1320 (O_1320,N_19895,N_19781);
or UO_1321 (O_1321,N_19025,N_19560);
or UO_1322 (O_1322,N_19332,N_19118);
xnor UO_1323 (O_1323,N_19047,N_19365);
xor UO_1324 (O_1324,N_19881,N_19399);
or UO_1325 (O_1325,N_19999,N_19073);
nor UO_1326 (O_1326,N_19345,N_19611);
nand UO_1327 (O_1327,N_19195,N_19205);
and UO_1328 (O_1328,N_19384,N_19490);
and UO_1329 (O_1329,N_19216,N_19550);
or UO_1330 (O_1330,N_19379,N_19285);
and UO_1331 (O_1331,N_19805,N_19993);
xor UO_1332 (O_1332,N_19609,N_19995);
or UO_1333 (O_1333,N_19434,N_19343);
xor UO_1334 (O_1334,N_19637,N_19191);
nand UO_1335 (O_1335,N_19663,N_19985);
xor UO_1336 (O_1336,N_19271,N_19567);
and UO_1337 (O_1337,N_19101,N_19044);
xor UO_1338 (O_1338,N_19945,N_19986);
nor UO_1339 (O_1339,N_19469,N_19292);
nor UO_1340 (O_1340,N_19205,N_19890);
xor UO_1341 (O_1341,N_19093,N_19705);
nand UO_1342 (O_1342,N_19587,N_19401);
nand UO_1343 (O_1343,N_19926,N_19869);
nand UO_1344 (O_1344,N_19583,N_19063);
nor UO_1345 (O_1345,N_19931,N_19287);
and UO_1346 (O_1346,N_19026,N_19216);
nand UO_1347 (O_1347,N_19866,N_19749);
xor UO_1348 (O_1348,N_19930,N_19490);
xor UO_1349 (O_1349,N_19105,N_19832);
or UO_1350 (O_1350,N_19001,N_19303);
nor UO_1351 (O_1351,N_19163,N_19004);
xnor UO_1352 (O_1352,N_19798,N_19618);
xnor UO_1353 (O_1353,N_19764,N_19552);
nand UO_1354 (O_1354,N_19234,N_19748);
nand UO_1355 (O_1355,N_19276,N_19583);
nor UO_1356 (O_1356,N_19144,N_19347);
and UO_1357 (O_1357,N_19577,N_19291);
or UO_1358 (O_1358,N_19908,N_19827);
nor UO_1359 (O_1359,N_19834,N_19304);
or UO_1360 (O_1360,N_19317,N_19872);
nand UO_1361 (O_1361,N_19708,N_19037);
and UO_1362 (O_1362,N_19912,N_19372);
and UO_1363 (O_1363,N_19316,N_19391);
and UO_1364 (O_1364,N_19395,N_19926);
or UO_1365 (O_1365,N_19660,N_19273);
nand UO_1366 (O_1366,N_19879,N_19778);
or UO_1367 (O_1367,N_19005,N_19330);
xor UO_1368 (O_1368,N_19009,N_19808);
nand UO_1369 (O_1369,N_19447,N_19438);
nor UO_1370 (O_1370,N_19002,N_19192);
nor UO_1371 (O_1371,N_19482,N_19097);
and UO_1372 (O_1372,N_19922,N_19073);
or UO_1373 (O_1373,N_19501,N_19361);
xnor UO_1374 (O_1374,N_19898,N_19353);
xnor UO_1375 (O_1375,N_19144,N_19871);
or UO_1376 (O_1376,N_19861,N_19510);
or UO_1377 (O_1377,N_19845,N_19515);
nor UO_1378 (O_1378,N_19491,N_19101);
nand UO_1379 (O_1379,N_19220,N_19703);
nor UO_1380 (O_1380,N_19649,N_19600);
and UO_1381 (O_1381,N_19089,N_19492);
nand UO_1382 (O_1382,N_19284,N_19015);
xor UO_1383 (O_1383,N_19402,N_19000);
xnor UO_1384 (O_1384,N_19813,N_19459);
or UO_1385 (O_1385,N_19371,N_19692);
nand UO_1386 (O_1386,N_19046,N_19280);
and UO_1387 (O_1387,N_19727,N_19656);
nand UO_1388 (O_1388,N_19128,N_19346);
xnor UO_1389 (O_1389,N_19886,N_19691);
nand UO_1390 (O_1390,N_19328,N_19820);
nor UO_1391 (O_1391,N_19848,N_19634);
nor UO_1392 (O_1392,N_19959,N_19984);
nor UO_1393 (O_1393,N_19770,N_19773);
nand UO_1394 (O_1394,N_19488,N_19659);
xnor UO_1395 (O_1395,N_19957,N_19088);
or UO_1396 (O_1396,N_19560,N_19955);
nor UO_1397 (O_1397,N_19120,N_19106);
and UO_1398 (O_1398,N_19473,N_19928);
or UO_1399 (O_1399,N_19541,N_19314);
or UO_1400 (O_1400,N_19000,N_19245);
xnor UO_1401 (O_1401,N_19786,N_19475);
or UO_1402 (O_1402,N_19195,N_19210);
xnor UO_1403 (O_1403,N_19898,N_19674);
nand UO_1404 (O_1404,N_19791,N_19365);
and UO_1405 (O_1405,N_19973,N_19101);
or UO_1406 (O_1406,N_19696,N_19664);
nor UO_1407 (O_1407,N_19225,N_19550);
or UO_1408 (O_1408,N_19124,N_19887);
or UO_1409 (O_1409,N_19695,N_19571);
nor UO_1410 (O_1410,N_19773,N_19082);
and UO_1411 (O_1411,N_19054,N_19100);
and UO_1412 (O_1412,N_19824,N_19062);
xnor UO_1413 (O_1413,N_19409,N_19454);
nor UO_1414 (O_1414,N_19328,N_19568);
and UO_1415 (O_1415,N_19723,N_19493);
xnor UO_1416 (O_1416,N_19734,N_19117);
and UO_1417 (O_1417,N_19093,N_19184);
nand UO_1418 (O_1418,N_19300,N_19318);
xnor UO_1419 (O_1419,N_19277,N_19616);
xor UO_1420 (O_1420,N_19047,N_19096);
nand UO_1421 (O_1421,N_19257,N_19319);
or UO_1422 (O_1422,N_19756,N_19271);
nor UO_1423 (O_1423,N_19805,N_19067);
xor UO_1424 (O_1424,N_19748,N_19576);
xor UO_1425 (O_1425,N_19297,N_19895);
nand UO_1426 (O_1426,N_19638,N_19770);
or UO_1427 (O_1427,N_19825,N_19021);
and UO_1428 (O_1428,N_19648,N_19413);
or UO_1429 (O_1429,N_19230,N_19550);
nand UO_1430 (O_1430,N_19013,N_19832);
nand UO_1431 (O_1431,N_19279,N_19206);
xor UO_1432 (O_1432,N_19877,N_19850);
or UO_1433 (O_1433,N_19906,N_19215);
nand UO_1434 (O_1434,N_19120,N_19457);
and UO_1435 (O_1435,N_19540,N_19902);
nand UO_1436 (O_1436,N_19159,N_19933);
xor UO_1437 (O_1437,N_19819,N_19479);
and UO_1438 (O_1438,N_19217,N_19174);
nor UO_1439 (O_1439,N_19847,N_19706);
or UO_1440 (O_1440,N_19748,N_19163);
xor UO_1441 (O_1441,N_19394,N_19259);
nand UO_1442 (O_1442,N_19440,N_19808);
nand UO_1443 (O_1443,N_19580,N_19696);
and UO_1444 (O_1444,N_19191,N_19945);
xor UO_1445 (O_1445,N_19739,N_19757);
nor UO_1446 (O_1446,N_19835,N_19057);
nor UO_1447 (O_1447,N_19846,N_19607);
and UO_1448 (O_1448,N_19463,N_19673);
or UO_1449 (O_1449,N_19778,N_19256);
nand UO_1450 (O_1450,N_19113,N_19930);
or UO_1451 (O_1451,N_19491,N_19936);
nand UO_1452 (O_1452,N_19101,N_19859);
or UO_1453 (O_1453,N_19636,N_19671);
nor UO_1454 (O_1454,N_19526,N_19923);
or UO_1455 (O_1455,N_19230,N_19115);
xnor UO_1456 (O_1456,N_19360,N_19208);
xor UO_1457 (O_1457,N_19277,N_19318);
and UO_1458 (O_1458,N_19257,N_19610);
nor UO_1459 (O_1459,N_19848,N_19998);
nor UO_1460 (O_1460,N_19154,N_19100);
and UO_1461 (O_1461,N_19377,N_19778);
or UO_1462 (O_1462,N_19010,N_19444);
or UO_1463 (O_1463,N_19125,N_19829);
or UO_1464 (O_1464,N_19938,N_19438);
nor UO_1465 (O_1465,N_19507,N_19648);
nor UO_1466 (O_1466,N_19135,N_19251);
nor UO_1467 (O_1467,N_19970,N_19653);
or UO_1468 (O_1468,N_19624,N_19893);
or UO_1469 (O_1469,N_19751,N_19687);
and UO_1470 (O_1470,N_19104,N_19891);
nor UO_1471 (O_1471,N_19525,N_19274);
nand UO_1472 (O_1472,N_19590,N_19592);
nor UO_1473 (O_1473,N_19608,N_19750);
nand UO_1474 (O_1474,N_19816,N_19177);
and UO_1475 (O_1475,N_19936,N_19567);
xnor UO_1476 (O_1476,N_19865,N_19222);
and UO_1477 (O_1477,N_19173,N_19557);
and UO_1478 (O_1478,N_19916,N_19094);
and UO_1479 (O_1479,N_19630,N_19654);
or UO_1480 (O_1480,N_19685,N_19517);
nand UO_1481 (O_1481,N_19114,N_19248);
xor UO_1482 (O_1482,N_19518,N_19862);
nand UO_1483 (O_1483,N_19454,N_19430);
or UO_1484 (O_1484,N_19694,N_19232);
and UO_1485 (O_1485,N_19004,N_19837);
or UO_1486 (O_1486,N_19427,N_19258);
xor UO_1487 (O_1487,N_19149,N_19161);
or UO_1488 (O_1488,N_19514,N_19929);
and UO_1489 (O_1489,N_19832,N_19708);
nand UO_1490 (O_1490,N_19950,N_19897);
xor UO_1491 (O_1491,N_19339,N_19808);
nand UO_1492 (O_1492,N_19495,N_19094);
nor UO_1493 (O_1493,N_19958,N_19190);
nor UO_1494 (O_1494,N_19514,N_19826);
nand UO_1495 (O_1495,N_19279,N_19449);
nand UO_1496 (O_1496,N_19507,N_19917);
xor UO_1497 (O_1497,N_19112,N_19643);
and UO_1498 (O_1498,N_19790,N_19992);
nand UO_1499 (O_1499,N_19680,N_19684);
nor UO_1500 (O_1500,N_19140,N_19830);
nand UO_1501 (O_1501,N_19480,N_19828);
xnor UO_1502 (O_1502,N_19176,N_19185);
and UO_1503 (O_1503,N_19468,N_19321);
nand UO_1504 (O_1504,N_19135,N_19200);
nand UO_1505 (O_1505,N_19177,N_19865);
xnor UO_1506 (O_1506,N_19028,N_19810);
nand UO_1507 (O_1507,N_19984,N_19949);
and UO_1508 (O_1508,N_19679,N_19215);
and UO_1509 (O_1509,N_19348,N_19486);
nor UO_1510 (O_1510,N_19345,N_19958);
nor UO_1511 (O_1511,N_19458,N_19975);
nand UO_1512 (O_1512,N_19891,N_19896);
nand UO_1513 (O_1513,N_19658,N_19615);
xor UO_1514 (O_1514,N_19884,N_19123);
nor UO_1515 (O_1515,N_19314,N_19578);
nor UO_1516 (O_1516,N_19776,N_19272);
nor UO_1517 (O_1517,N_19772,N_19408);
nor UO_1518 (O_1518,N_19732,N_19307);
and UO_1519 (O_1519,N_19205,N_19887);
nand UO_1520 (O_1520,N_19240,N_19884);
and UO_1521 (O_1521,N_19274,N_19675);
nor UO_1522 (O_1522,N_19365,N_19230);
nor UO_1523 (O_1523,N_19110,N_19152);
nand UO_1524 (O_1524,N_19558,N_19899);
nand UO_1525 (O_1525,N_19360,N_19990);
nand UO_1526 (O_1526,N_19484,N_19524);
and UO_1527 (O_1527,N_19524,N_19500);
or UO_1528 (O_1528,N_19830,N_19714);
xor UO_1529 (O_1529,N_19555,N_19898);
or UO_1530 (O_1530,N_19217,N_19696);
and UO_1531 (O_1531,N_19616,N_19353);
or UO_1532 (O_1532,N_19108,N_19870);
nor UO_1533 (O_1533,N_19218,N_19748);
and UO_1534 (O_1534,N_19267,N_19025);
nor UO_1535 (O_1535,N_19132,N_19418);
nand UO_1536 (O_1536,N_19951,N_19230);
or UO_1537 (O_1537,N_19391,N_19025);
nor UO_1538 (O_1538,N_19501,N_19564);
and UO_1539 (O_1539,N_19945,N_19688);
nor UO_1540 (O_1540,N_19993,N_19125);
and UO_1541 (O_1541,N_19102,N_19963);
or UO_1542 (O_1542,N_19584,N_19640);
or UO_1543 (O_1543,N_19549,N_19266);
nor UO_1544 (O_1544,N_19409,N_19400);
nand UO_1545 (O_1545,N_19999,N_19127);
nor UO_1546 (O_1546,N_19818,N_19098);
and UO_1547 (O_1547,N_19645,N_19816);
xnor UO_1548 (O_1548,N_19932,N_19619);
and UO_1549 (O_1549,N_19592,N_19402);
nand UO_1550 (O_1550,N_19923,N_19502);
xor UO_1551 (O_1551,N_19329,N_19136);
xnor UO_1552 (O_1552,N_19623,N_19969);
nor UO_1553 (O_1553,N_19104,N_19343);
nor UO_1554 (O_1554,N_19107,N_19280);
and UO_1555 (O_1555,N_19985,N_19717);
or UO_1556 (O_1556,N_19143,N_19539);
nor UO_1557 (O_1557,N_19233,N_19683);
or UO_1558 (O_1558,N_19692,N_19813);
and UO_1559 (O_1559,N_19133,N_19851);
and UO_1560 (O_1560,N_19828,N_19132);
xor UO_1561 (O_1561,N_19077,N_19121);
xor UO_1562 (O_1562,N_19319,N_19869);
and UO_1563 (O_1563,N_19287,N_19541);
and UO_1564 (O_1564,N_19443,N_19349);
xnor UO_1565 (O_1565,N_19560,N_19201);
or UO_1566 (O_1566,N_19846,N_19789);
nand UO_1567 (O_1567,N_19837,N_19563);
and UO_1568 (O_1568,N_19807,N_19754);
and UO_1569 (O_1569,N_19555,N_19145);
nor UO_1570 (O_1570,N_19839,N_19935);
or UO_1571 (O_1571,N_19739,N_19643);
and UO_1572 (O_1572,N_19029,N_19547);
xor UO_1573 (O_1573,N_19414,N_19855);
nand UO_1574 (O_1574,N_19432,N_19475);
and UO_1575 (O_1575,N_19179,N_19175);
xnor UO_1576 (O_1576,N_19266,N_19811);
nor UO_1577 (O_1577,N_19964,N_19443);
nor UO_1578 (O_1578,N_19037,N_19859);
xnor UO_1579 (O_1579,N_19768,N_19686);
xor UO_1580 (O_1580,N_19805,N_19030);
nor UO_1581 (O_1581,N_19751,N_19456);
xor UO_1582 (O_1582,N_19476,N_19443);
and UO_1583 (O_1583,N_19710,N_19676);
and UO_1584 (O_1584,N_19383,N_19037);
xor UO_1585 (O_1585,N_19721,N_19379);
xor UO_1586 (O_1586,N_19897,N_19213);
xor UO_1587 (O_1587,N_19089,N_19446);
and UO_1588 (O_1588,N_19194,N_19370);
or UO_1589 (O_1589,N_19226,N_19264);
nor UO_1590 (O_1590,N_19642,N_19397);
nor UO_1591 (O_1591,N_19418,N_19086);
or UO_1592 (O_1592,N_19292,N_19200);
nand UO_1593 (O_1593,N_19786,N_19850);
or UO_1594 (O_1594,N_19632,N_19690);
xnor UO_1595 (O_1595,N_19895,N_19820);
or UO_1596 (O_1596,N_19699,N_19173);
nand UO_1597 (O_1597,N_19555,N_19756);
xor UO_1598 (O_1598,N_19475,N_19993);
or UO_1599 (O_1599,N_19290,N_19074);
and UO_1600 (O_1600,N_19572,N_19793);
or UO_1601 (O_1601,N_19910,N_19679);
nand UO_1602 (O_1602,N_19735,N_19409);
xor UO_1603 (O_1603,N_19125,N_19948);
nand UO_1604 (O_1604,N_19997,N_19394);
nor UO_1605 (O_1605,N_19664,N_19076);
nor UO_1606 (O_1606,N_19117,N_19905);
xor UO_1607 (O_1607,N_19855,N_19084);
nor UO_1608 (O_1608,N_19350,N_19596);
nand UO_1609 (O_1609,N_19679,N_19960);
nor UO_1610 (O_1610,N_19332,N_19868);
nor UO_1611 (O_1611,N_19746,N_19735);
xnor UO_1612 (O_1612,N_19644,N_19166);
nand UO_1613 (O_1613,N_19938,N_19366);
xnor UO_1614 (O_1614,N_19724,N_19941);
or UO_1615 (O_1615,N_19600,N_19127);
and UO_1616 (O_1616,N_19853,N_19371);
nor UO_1617 (O_1617,N_19395,N_19879);
nand UO_1618 (O_1618,N_19899,N_19876);
nor UO_1619 (O_1619,N_19873,N_19579);
or UO_1620 (O_1620,N_19957,N_19080);
nor UO_1621 (O_1621,N_19204,N_19189);
or UO_1622 (O_1622,N_19380,N_19871);
nand UO_1623 (O_1623,N_19444,N_19793);
or UO_1624 (O_1624,N_19947,N_19847);
and UO_1625 (O_1625,N_19019,N_19988);
nand UO_1626 (O_1626,N_19894,N_19562);
nor UO_1627 (O_1627,N_19203,N_19812);
nor UO_1628 (O_1628,N_19767,N_19908);
nor UO_1629 (O_1629,N_19314,N_19750);
and UO_1630 (O_1630,N_19148,N_19851);
and UO_1631 (O_1631,N_19956,N_19429);
nor UO_1632 (O_1632,N_19500,N_19038);
nor UO_1633 (O_1633,N_19674,N_19322);
nor UO_1634 (O_1634,N_19395,N_19636);
nor UO_1635 (O_1635,N_19358,N_19850);
nand UO_1636 (O_1636,N_19241,N_19733);
and UO_1637 (O_1637,N_19658,N_19181);
nor UO_1638 (O_1638,N_19275,N_19061);
xnor UO_1639 (O_1639,N_19894,N_19129);
nor UO_1640 (O_1640,N_19799,N_19511);
or UO_1641 (O_1641,N_19961,N_19927);
xor UO_1642 (O_1642,N_19926,N_19955);
and UO_1643 (O_1643,N_19216,N_19049);
and UO_1644 (O_1644,N_19670,N_19315);
or UO_1645 (O_1645,N_19992,N_19384);
nor UO_1646 (O_1646,N_19490,N_19267);
and UO_1647 (O_1647,N_19746,N_19994);
and UO_1648 (O_1648,N_19299,N_19150);
and UO_1649 (O_1649,N_19953,N_19594);
and UO_1650 (O_1650,N_19063,N_19145);
or UO_1651 (O_1651,N_19483,N_19885);
xnor UO_1652 (O_1652,N_19929,N_19526);
nor UO_1653 (O_1653,N_19206,N_19431);
nand UO_1654 (O_1654,N_19649,N_19729);
and UO_1655 (O_1655,N_19708,N_19087);
xor UO_1656 (O_1656,N_19551,N_19864);
nand UO_1657 (O_1657,N_19509,N_19643);
nand UO_1658 (O_1658,N_19283,N_19857);
and UO_1659 (O_1659,N_19981,N_19416);
nor UO_1660 (O_1660,N_19986,N_19264);
or UO_1661 (O_1661,N_19621,N_19473);
and UO_1662 (O_1662,N_19740,N_19695);
and UO_1663 (O_1663,N_19143,N_19077);
or UO_1664 (O_1664,N_19156,N_19835);
nand UO_1665 (O_1665,N_19184,N_19978);
or UO_1666 (O_1666,N_19111,N_19222);
and UO_1667 (O_1667,N_19791,N_19751);
and UO_1668 (O_1668,N_19444,N_19070);
nor UO_1669 (O_1669,N_19729,N_19555);
and UO_1670 (O_1670,N_19575,N_19659);
or UO_1671 (O_1671,N_19492,N_19824);
xor UO_1672 (O_1672,N_19801,N_19644);
nor UO_1673 (O_1673,N_19854,N_19640);
nor UO_1674 (O_1674,N_19311,N_19770);
or UO_1675 (O_1675,N_19408,N_19040);
or UO_1676 (O_1676,N_19294,N_19964);
nor UO_1677 (O_1677,N_19682,N_19422);
nor UO_1678 (O_1678,N_19855,N_19232);
nand UO_1679 (O_1679,N_19983,N_19719);
nor UO_1680 (O_1680,N_19916,N_19880);
xnor UO_1681 (O_1681,N_19778,N_19922);
nand UO_1682 (O_1682,N_19328,N_19142);
nor UO_1683 (O_1683,N_19077,N_19111);
nand UO_1684 (O_1684,N_19816,N_19825);
nand UO_1685 (O_1685,N_19004,N_19682);
xnor UO_1686 (O_1686,N_19397,N_19974);
nor UO_1687 (O_1687,N_19502,N_19365);
xor UO_1688 (O_1688,N_19375,N_19956);
xnor UO_1689 (O_1689,N_19570,N_19444);
and UO_1690 (O_1690,N_19161,N_19586);
xnor UO_1691 (O_1691,N_19237,N_19500);
nand UO_1692 (O_1692,N_19252,N_19552);
xnor UO_1693 (O_1693,N_19075,N_19989);
and UO_1694 (O_1694,N_19286,N_19082);
and UO_1695 (O_1695,N_19891,N_19329);
xor UO_1696 (O_1696,N_19092,N_19943);
nand UO_1697 (O_1697,N_19157,N_19512);
nor UO_1698 (O_1698,N_19306,N_19156);
and UO_1699 (O_1699,N_19995,N_19792);
nand UO_1700 (O_1700,N_19715,N_19401);
nand UO_1701 (O_1701,N_19247,N_19249);
xnor UO_1702 (O_1702,N_19328,N_19606);
or UO_1703 (O_1703,N_19348,N_19853);
nand UO_1704 (O_1704,N_19912,N_19856);
and UO_1705 (O_1705,N_19791,N_19963);
or UO_1706 (O_1706,N_19198,N_19354);
nor UO_1707 (O_1707,N_19713,N_19585);
or UO_1708 (O_1708,N_19585,N_19275);
nand UO_1709 (O_1709,N_19863,N_19891);
nor UO_1710 (O_1710,N_19063,N_19367);
xnor UO_1711 (O_1711,N_19204,N_19434);
nor UO_1712 (O_1712,N_19147,N_19137);
and UO_1713 (O_1713,N_19104,N_19365);
and UO_1714 (O_1714,N_19327,N_19227);
and UO_1715 (O_1715,N_19896,N_19985);
nand UO_1716 (O_1716,N_19792,N_19121);
and UO_1717 (O_1717,N_19020,N_19333);
nand UO_1718 (O_1718,N_19523,N_19031);
nor UO_1719 (O_1719,N_19192,N_19791);
or UO_1720 (O_1720,N_19319,N_19328);
nor UO_1721 (O_1721,N_19668,N_19563);
and UO_1722 (O_1722,N_19952,N_19660);
nor UO_1723 (O_1723,N_19081,N_19079);
nor UO_1724 (O_1724,N_19201,N_19456);
or UO_1725 (O_1725,N_19900,N_19739);
xor UO_1726 (O_1726,N_19169,N_19243);
nor UO_1727 (O_1727,N_19330,N_19248);
nor UO_1728 (O_1728,N_19102,N_19004);
or UO_1729 (O_1729,N_19622,N_19233);
nor UO_1730 (O_1730,N_19533,N_19716);
xor UO_1731 (O_1731,N_19522,N_19828);
xor UO_1732 (O_1732,N_19889,N_19220);
or UO_1733 (O_1733,N_19206,N_19289);
or UO_1734 (O_1734,N_19708,N_19101);
nor UO_1735 (O_1735,N_19132,N_19749);
nand UO_1736 (O_1736,N_19993,N_19529);
or UO_1737 (O_1737,N_19626,N_19325);
nor UO_1738 (O_1738,N_19608,N_19480);
and UO_1739 (O_1739,N_19445,N_19249);
nand UO_1740 (O_1740,N_19292,N_19853);
nand UO_1741 (O_1741,N_19285,N_19389);
and UO_1742 (O_1742,N_19377,N_19595);
nor UO_1743 (O_1743,N_19122,N_19403);
nand UO_1744 (O_1744,N_19239,N_19225);
or UO_1745 (O_1745,N_19207,N_19219);
nor UO_1746 (O_1746,N_19624,N_19081);
or UO_1747 (O_1747,N_19185,N_19838);
and UO_1748 (O_1748,N_19266,N_19881);
nor UO_1749 (O_1749,N_19267,N_19013);
and UO_1750 (O_1750,N_19253,N_19102);
nand UO_1751 (O_1751,N_19328,N_19676);
or UO_1752 (O_1752,N_19087,N_19185);
nor UO_1753 (O_1753,N_19789,N_19055);
nand UO_1754 (O_1754,N_19032,N_19072);
or UO_1755 (O_1755,N_19867,N_19499);
xnor UO_1756 (O_1756,N_19971,N_19995);
nor UO_1757 (O_1757,N_19039,N_19544);
nand UO_1758 (O_1758,N_19202,N_19594);
nor UO_1759 (O_1759,N_19004,N_19382);
nand UO_1760 (O_1760,N_19994,N_19392);
nor UO_1761 (O_1761,N_19764,N_19429);
nand UO_1762 (O_1762,N_19706,N_19774);
nor UO_1763 (O_1763,N_19888,N_19301);
xnor UO_1764 (O_1764,N_19641,N_19118);
nand UO_1765 (O_1765,N_19345,N_19769);
nand UO_1766 (O_1766,N_19333,N_19530);
nand UO_1767 (O_1767,N_19781,N_19112);
and UO_1768 (O_1768,N_19095,N_19621);
and UO_1769 (O_1769,N_19813,N_19254);
nor UO_1770 (O_1770,N_19636,N_19869);
nor UO_1771 (O_1771,N_19134,N_19893);
nand UO_1772 (O_1772,N_19008,N_19193);
xor UO_1773 (O_1773,N_19706,N_19681);
or UO_1774 (O_1774,N_19130,N_19772);
or UO_1775 (O_1775,N_19878,N_19048);
nand UO_1776 (O_1776,N_19967,N_19326);
and UO_1777 (O_1777,N_19372,N_19306);
nor UO_1778 (O_1778,N_19253,N_19980);
nor UO_1779 (O_1779,N_19777,N_19166);
nand UO_1780 (O_1780,N_19041,N_19011);
nor UO_1781 (O_1781,N_19785,N_19799);
nand UO_1782 (O_1782,N_19638,N_19666);
nand UO_1783 (O_1783,N_19469,N_19993);
nor UO_1784 (O_1784,N_19822,N_19075);
nor UO_1785 (O_1785,N_19433,N_19284);
nor UO_1786 (O_1786,N_19149,N_19049);
xor UO_1787 (O_1787,N_19764,N_19916);
and UO_1788 (O_1788,N_19240,N_19670);
and UO_1789 (O_1789,N_19046,N_19260);
nor UO_1790 (O_1790,N_19803,N_19440);
and UO_1791 (O_1791,N_19519,N_19906);
nor UO_1792 (O_1792,N_19553,N_19906);
nand UO_1793 (O_1793,N_19743,N_19084);
or UO_1794 (O_1794,N_19446,N_19230);
or UO_1795 (O_1795,N_19376,N_19773);
xnor UO_1796 (O_1796,N_19246,N_19664);
nor UO_1797 (O_1797,N_19716,N_19275);
nand UO_1798 (O_1798,N_19263,N_19184);
nor UO_1799 (O_1799,N_19771,N_19523);
nand UO_1800 (O_1800,N_19155,N_19472);
or UO_1801 (O_1801,N_19167,N_19147);
or UO_1802 (O_1802,N_19418,N_19612);
or UO_1803 (O_1803,N_19860,N_19763);
nand UO_1804 (O_1804,N_19805,N_19755);
nand UO_1805 (O_1805,N_19472,N_19697);
nor UO_1806 (O_1806,N_19205,N_19177);
and UO_1807 (O_1807,N_19025,N_19613);
nand UO_1808 (O_1808,N_19578,N_19167);
nor UO_1809 (O_1809,N_19885,N_19931);
and UO_1810 (O_1810,N_19230,N_19056);
nor UO_1811 (O_1811,N_19432,N_19304);
nor UO_1812 (O_1812,N_19534,N_19183);
nand UO_1813 (O_1813,N_19426,N_19792);
and UO_1814 (O_1814,N_19750,N_19293);
nor UO_1815 (O_1815,N_19072,N_19566);
and UO_1816 (O_1816,N_19478,N_19061);
and UO_1817 (O_1817,N_19326,N_19976);
and UO_1818 (O_1818,N_19173,N_19291);
or UO_1819 (O_1819,N_19529,N_19549);
and UO_1820 (O_1820,N_19178,N_19193);
nor UO_1821 (O_1821,N_19741,N_19585);
nand UO_1822 (O_1822,N_19401,N_19779);
and UO_1823 (O_1823,N_19266,N_19801);
nor UO_1824 (O_1824,N_19694,N_19581);
xor UO_1825 (O_1825,N_19277,N_19795);
or UO_1826 (O_1826,N_19781,N_19541);
nand UO_1827 (O_1827,N_19806,N_19202);
nand UO_1828 (O_1828,N_19091,N_19403);
or UO_1829 (O_1829,N_19760,N_19993);
and UO_1830 (O_1830,N_19084,N_19103);
or UO_1831 (O_1831,N_19644,N_19516);
or UO_1832 (O_1832,N_19763,N_19743);
xnor UO_1833 (O_1833,N_19103,N_19003);
or UO_1834 (O_1834,N_19202,N_19246);
nor UO_1835 (O_1835,N_19466,N_19732);
nand UO_1836 (O_1836,N_19389,N_19415);
xnor UO_1837 (O_1837,N_19218,N_19622);
nand UO_1838 (O_1838,N_19298,N_19814);
nor UO_1839 (O_1839,N_19241,N_19414);
nand UO_1840 (O_1840,N_19354,N_19500);
nand UO_1841 (O_1841,N_19313,N_19110);
nand UO_1842 (O_1842,N_19357,N_19342);
nand UO_1843 (O_1843,N_19149,N_19329);
and UO_1844 (O_1844,N_19808,N_19920);
xor UO_1845 (O_1845,N_19574,N_19192);
nand UO_1846 (O_1846,N_19110,N_19743);
xnor UO_1847 (O_1847,N_19613,N_19100);
nor UO_1848 (O_1848,N_19766,N_19046);
xor UO_1849 (O_1849,N_19490,N_19294);
nand UO_1850 (O_1850,N_19276,N_19225);
nand UO_1851 (O_1851,N_19586,N_19640);
nand UO_1852 (O_1852,N_19433,N_19259);
xnor UO_1853 (O_1853,N_19024,N_19213);
or UO_1854 (O_1854,N_19469,N_19137);
or UO_1855 (O_1855,N_19732,N_19429);
xnor UO_1856 (O_1856,N_19829,N_19106);
or UO_1857 (O_1857,N_19746,N_19297);
and UO_1858 (O_1858,N_19133,N_19718);
nand UO_1859 (O_1859,N_19616,N_19946);
xor UO_1860 (O_1860,N_19861,N_19760);
xnor UO_1861 (O_1861,N_19181,N_19092);
xor UO_1862 (O_1862,N_19999,N_19375);
xnor UO_1863 (O_1863,N_19896,N_19051);
or UO_1864 (O_1864,N_19562,N_19968);
or UO_1865 (O_1865,N_19129,N_19883);
or UO_1866 (O_1866,N_19783,N_19879);
xnor UO_1867 (O_1867,N_19178,N_19880);
nor UO_1868 (O_1868,N_19532,N_19716);
xor UO_1869 (O_1869,N_19950,N_19303);
nor UO_1870 (O_1870,N_19056,N_19674);
or UO_1871 (O_1871,N_19732,N_19035);
nand UO_1872 (O_1872,N_19015,N_19188);
and UO_1873 (O_1873,N_19118,N_19699);
or UO_1874 (O_1874,N_19790,N_19430);
or UO_1875 (O_1875,N_19254,N_19275);
xor UO_1876 (O_1876,N_19809,N_19244);
and UO_1877 (O_1877,N_19826,N_19199);
or UO_1878 (O_1878,N_19450,N_19624);
nand UO_1879 (O_1879,N_19831,N_19055);
and UO_1880 (O_1880,N_19915,N_19348);
or UO_1881 (O_1881,N_19536,N_19470);
xor UO_1882 (O_1882,N_19526,N_19358);
or UO_1883 (O_1883,N_19868,N_19723);
xor UO_1884 (O_1884,N_19079,N_19903);
nor UO_1885 (O_1885,N_19303,N_19639);
and UO_1886 (O_1886,N_19299,N_19110);
nor UO_1887 (O_1887,N_19509,N_19505);
xor UO_1888 (O_1888,N_19692,N_19969);
nand UO_1889 (O_1889,N_19281,N_19038);
nand UO_1890 (O_1890,N_19942,N_19471);
nand UO_1891 (O_1891,N_19723,N_19166);
and UO_1892 (O_1892,N_19105,N_19656);
and UO_1893 (O_1893,N_19618,N_19269);
xor UO_1894 (O_1894,N_19650,N_19515);
and UO_1895 (O_1895,N_19845,N_19206);
nand UO_1896 (O_1896,N_19721,N_19726);
or UO_1897 (O_1897,N_19740,N_19413);
or UO_1898 (O_1898,N_19929,N_19633);
nand UO_1899 (O_1899,N_19878,N_19588);
xor UO_1900 (O_1900,N_19381,N_19011);
xor UO_1901 (O_1901,N_19246,N_19959);
and UO_1902 (O_1902,N_19478,N_19163);
nand UO_1903 (O_1903,N_19159,N_19878);
or UO_1904 (O_1904,N_19685,N_19816);
and UO_1905 (O_1905,N_19377,N_19965);
xnor UO_1906 (O_1906,N_19034,N_19037);
and UO_1907 (O_1907,N_19258,N_19896);
nand UO_1908 (O_1908,N_19189,N_19736);
xor UO_1909 (O_1909,N_19390,N_19651);
nor UO_1910 (O_1910,N_19145,N_19711);
nand UO_1911 (O_1911,N_19606,N_19388);
or UO_1912 (O_1912,N_19936,N_19509);
or UO_1913 (O_1913,N_19763,N_19883);
nand UO_1914 (O_1914,N_19166,N_19967);
or UO_1915 (O_1915,N_19381,N_19906);
and UO_1916 (O_1916,N_19719,N_19274);
nor UO_1917 (O_1917,N_19278,N_19634);
and UO_1918 (O_1918,N_19913,N_19046);
and UO_1919 (O_1919,N_19811,N_19305);
and UO_1920 (O_1920,N_19797,N_19509);
nor UO_1921 (O_1921,N_19603,N_19385);
nor UO_1922 (O_1922,N_19353,N_19646);
or UO_1923 (O_1923,N_19085,N_19616);
and UO_1924 (O_1924,N_19568,N_19454);
nand UO_1925 (O_1925,N_19842,N_19664);
or UO_1926 (O_1926,N_19351,N_19116);
nor UO_1927 (O_1927,N_19026,N_19659);
or UO_1928 (O_1928,N_19349,N_19350);
nand UO_1929 (O_1929,N_19973,N_19859);
and UO_1930 (O_1930,N_19562,N_19093);
nand UO_1931 (O_1931,N_19926,N_19799);
and UO_1932 (O_1932,N_19478,N_19912);
nand UO_1933 (O_1933,N_19112,N_19976);
nor UO_1934 (O_1934,N_19856,N_19114);
nor UO_1935 (O_1935,N_19968,N_19854);
nand UO_1936 (O_1936,N_19993,N_19297);
xor UO_1937 (O_1937,N_19651,N_19636);
or UO_1938 (O_1938,N_19738,N_19093);
and UO_1939 (O_1939,N_19536,N_19532);
and UO_1940 (O_1940,N_19523,N_19990);
or UO_1941 (O_1941,N_19796,N_19662);
nor UO_1942 (O_1942,N_19121,N_19179);
and UO_1943 (O_1943,N_19075,N_19515);
and UO_1944 (O_1944,N_19871,N_19154);
nand UO_1945 (O_1945,N_19307,N_19304);
nand UO_1946 (O_1946,N_19308,N_19811);
xnor UO_1947 (O_1947,N_19388,N_19047);
and UO_1948 (O_1948,N_19245,N_19983);
nand UO_1949 (O_1949,N_19947,N_19929);
xor UO_1950 (O_1950,N_19997,N_19190);
nand UO_1951 (O_1951,N_19755,N_19424);
xnor UO_1952 (O_1952,N_19633,N_19151);
xor UO_1953 (O_1953,N_19528,N_19467);
xnor UO_1954 (O_1954,N_19259,N_19526);
and UO_1955 (O_1955,N_19897,N_19769);
xor UO_1956 (O_1956,N_19705,N_19175);
xor UO_1957 (O_1957,N_19892,N_19691);
or UO_1958 (O_1958,N_19491,N_19144);
or UO_1959 (O_1959,N_19529,N_19025);
xnor UO_1960 (O_1960,N_19704,N_19799);
xor UO_1961 (O_1961,N_19581,N_19416);
xnor UO_1962 (O_1962,N_19522,N_19532);
nand UO_1963 (O_1963,N_19059,N_19337);
nand UO_1964 (O_1964,N_19775,N_19077);
nand UO_1965 (O_1965,N_19564,N_19949);
xnor UO_1966 (O_1966,N_19400,N_19719);
nor UO_1967 (O_1967,N_19570,N_19919);
xor UO_1968 (O_1968,N_19431,N_19058);
or UO_1969 (O_1969,N_19162,N_19319);
or UO_1970 (O_1970,N_19731,N_19984);
and UO_1971 (O_1971,N_19328,N_19954);
or UO_1972 (O_1972,N_19960,N_19163);
xnor UO_1973 (O_1973,N_19538,N_19832);
nand UO_1974 (O_1974,N_19588,N_19895);
and UO_1975 (O_1975,N_19993,N_19746);
nand UO_1976 (O_1976,N_19879,N_19698);
nor UO_1977 (O_1977,N_19863,N_19429);
or UO_1978 (O_1978,N_19188,N_19505);
or UO_1979 (O_1979,N_19759,N_19773);
or UO_1980 (O_1980,N_19647,N_19507);
nand UO_1981 (O_1981,N_19219,N_19292);
or UO_1982 (O_1982,N_19526,N_19254);
nand UO_1983 (O_1983,N_19683,N_19332);
and UO_1984 (O_1984,N_19965,N_19735);
nor UO_1985 (O_1985,N_19437,N_19113);
nand UO_1986 (O_1986,N_19200,N_19778);
nor UO_1987 (O_1987,N_19545,N_19743);
or UO_1988 (O_1988,N_19473,N_19996);
nor UO_1989 (O_1989,N_19637,N_19607);
nand UO_1990 (O_1990,N_19413,N_19435);
nor UO_1991 (O_1991,N_19552,N_19240);
and UO_1992 (O_1992,N_19342,N_19616);
xor UO_1993 (O_1993,N_19092,N_19649);
nor UO_1994 (O_1994,N_19216,N_19101);
xor UO_1995 (O_1995,N_19385,N_19574);
nand UO_1996 (O_1996,N_19224,N_19322);
nor UO_1997 (O_1997,N_19138,N_19335);
and UO_1998 (O_1998,N_19382,N_19975);
nor UO_1999 (O_1999,N_19119,N_19020);
xnor UO_2000 (O_2000,N_19567,N_19602);
and UO_2001 (O_2001,N_19523,N_19272);
xnor UO_2002 (O_2002,N_19066,N_19640);
nor UO_2003 (O_2003,N_19300,N_19496);
xnor UO_2004 (O_2004,N_19049,N_19873);
xnor UO_2005 (O_2005,N_19706,N_19055);
and UO_2006 (O_2006,N_19558,N_19543);
xnor UO_2007 (O_2007,N_19659,N_19457);
nor UO_2008 (O_2008,N_19255,N_19279);
xnor UO_2009 (O_2009,N_19866,N_19393);
xnor UO_2010 (O_2010,N_19816,N_19952);
xnor UO_2011 (O_2011,N_19054,N_19281);
and UO_2012 (O_2012,N_19084,N_19775);
nor UO_2013 (O_2013,N_19269,N_19250);
xnor UO_2014 (O_2014,N_19427,N_19585);
nor UO_2015 (O_2015,N_19816,N_19391);
nor UO_2016 (O_2016,N_19533,N_19520);
nand UO_2017 (O_2017,N_19066,N_19035);
xnor UO_2018 (O_2018,N_19927,N_19615);
or UO_2019 (O_2019,N_19557,N_19639);
nor UO_2020 (O_2020,N_19316,N_19500);
nor UO_2021 (O_2021,N_19174,N_19224);
and UO_2022 (O_2022,N_19603,N_19221);
and UO_2023 (O_2023,N_19002,N_19929);
and UO_2024 (O_2024,N_19315,N_19665);
nand UO_2025 (O_2025,N_19310,N_19563);
and UO_2026 (O_2026,N_19670,N_19197);
xnor UO_2027 (O_2027,N_19797,N_19822);
xnor UO_2028 (O_2028,N_19160,N_19192);
and UO_2029 (O_2029,N_19148,N_19968);
and UO_2030 (O_2030,N_19113,N_19358);
and UO_2031 (O_2031,N_19603,N_19601);
or UO_2032 (O_2032,N_19504,N_19832);
xnor UO_2033 (O_2033,N_19943,N_19019);
and UO_2034 (O_2034,N_19568,N_19880);
xor UO_2035 (O_2035,N_19573,N_19707);
or UO_2036 (O_2036,N_19420,N_19215);
xor UO_2037 (O_2037,N_19859,N_19337);
and UO_2038 (O_2038,N_19906,N_19335);
or UO_2039 (O_2039,N_19047,N_19581);
and UO_2040 (O_2040,N_19424,N_19348);
and UO_2041 (O_2041,N_19888,N_19033);
nand UO_2042 (O_2042,N_19898,N_19067);
and UO_2043 (O_2043,N_19986,N_19779);
nor UO_2044 (O_2044,N_19820,N_19572);
xor UO_2045 (O_2045,N_19629,N_19210);
and UO_2046 (O_2046,N_19063,N_19099);
and UO_2047 (O_2047,N_19470,N_19181);
or UO_2048 (O_2048,N_19286,N_19582);
or UO_2049 (O_2049,N_19213,N_19646);
xnor UO_2050 (O_2050,N_19456,N_19188);
nor UO_2051 (O_2051,N_19311,N_19526);
and UO_2052 (O_2052,N_19975,N_19922);
xor UO_2053 (O_2053,N_19191,N_19030);
or UO_2054 (O_2054,N_19023,N_19018);
nor UO_2055 (O_2055,N_19730,N_19487);
and UO_2056 (O_2056,N_19318,N_19791);
and UO_2057 (O_2057,N_19010,N_19525);
xor UO_2058 (O_2058,N_19815,N_19128);
nand UO_2059 (O_2059,N_19625,N_19007);
and UO_2060 (O_2060,N_19776,N_19749);
xnor UO_2061 (O_2061,N_19228,N_19431);
or UO_2062 (O_2062,N_19027,N_19644);
and UO_2063 (O_2063,N_19424,N_19688);
and UO_2064 (O_2064,N_19176,N_19250);
or UO_2065 (O_2065,N_19371,N_19584);
nand UO_2066 (O_2066,N_19257,N_19743);
and UO_2067 (O_2067,N_19076,N_19352);
and UO_2068 (O_2068,N_19076,N_19269);
nand UO_2069 (O_2069,N_19160,N_19612);
nor UO_2070 (O_2070,N_19791,N_19358);
or UO_2071 (O_2071,N_19607,N_19566);
xor UO_2072 (O_2072,N_19558,N_19668);
nand UO_2073 (O_2073,N_19312,N_19062);
nand UO_2074 (O_2074,N_19857,N_19557);
or UO_2075 (O_2075,N_19068,N_19783);
nor UO_2076 (O_2076,N_19404,N_19329);
and UO_2077 (O_2077,N_19205,N_19567);
and UO_2078 (O_2078,N_19042,N_19897);
or UO_2079 (O_2079,N_19544,N_19540);
or UO_2080 (O_2080,N_19623,N_19175);
and UO_2081 (O_2081,N_19035,N_19202);
nor UO_2082 (O_2082,N_19760,N_19697);
nand UO_2083 (O_2083,N_19317,N_19783);
xnor UO_2084 (O_2084,N_19392,N_19501);
nor UO_2085 (O_2085,N_19598,N_19446);
nor UO_2086 (O_2086,N_19980,N_19989);
and UO_2087 (O_2087,N_19277,N_19159);
or UO_2088 (O_2088,N_19107,N_19963);
nand UO_2089 (O_2089,N_19868,N_19537);
xor UO_2090 (O_2090,N_19205,N_19512);
and UO_2091 (O_2091,N_19680,N_19113);
nand UO_2092 (O_2092,N_19297,N_19132);
xor UO_2093 (O_2093,N_19654,N_19549);
xnor UO_2094 (O_2094,N_19621,N_19044);
nor UO_2095 (O_2095,N_19004,N_19416);
nand UO_2096 (O_2096,N_19757,N_19177);
and UO_2097 (O_2097,N_19393,N_19050);
nor UO_2098 (O_2098,N_19447,N_19549);
nor UO_2099 (O_2099,N_19452,N_19691);
nand UO_2100 (O_2100,N_19076,N_19743);
nor UO_2101 (O_2101,N_19884,N_19313);
and UO_2102 (O_2102,N_19518,N_19541);
or UO_2103 (O_2103,N_19305,N_19742);
and UO_2104 (O_2104,N_19696,N_19749);
nand UO_2105 (O_2105,N_19521,N_19641);
nor UO_2106 (O_2106,N_19215,N_19179);
and UO_2107 (O_2107,N_19424,N_19269);
nor UO_2108 (O_2108,N_19486,N_19157);
nor UO_2109 (O_2109,N_19789,N_19851);
nand UO_2110 (O_2110,N_19230,N_19588);
or UO_2111 (O_2111,N_19508,N_19528);
xor UO_2112 (O_2112,N_19370,N_19353);
or UO_2113 (O_2113,N_19655,N_19268);
nor UO_2114 (O_2114,N_19137,N_19963);
xor UO_2115 (O_2115,N_19337,N_19750);
nand UO_2116 (O_2116,N_19305,N_19488);
nor UO_2117 (O_2117,N_19554,N_19845);
nand UO_2118 (O_2118,N_19565,N_19746);
xor UO_2119 (O_2119,N_19364,N_19641);
or UO_2120 (O_2120,N_19783,N_19937);
nor UO_2121 (O_2121,N_19052,N_19298);
nand UO_2122 (O_2122,N_19573,N_19896);
nand UO_2123 (O_2123,N_19040,N_19718);
or UO_2124 (O_2124,N_19331,N_19146);
or UO_2125 (O_2125,N_19099,N_19017);
and UO_2126 (O_2126,N_19027,N_19508);
xnor UO_2127 (O_2127,N_19110,N_19577);
nor UO_2128 (O_2128,N_19254,N_19552);
or UO_2129 (O_2129,N_19294,N_19183);
nor UO_2130 (O_2130,N_19567,N_19647);
nand UO_2131 (O_2131,N_19323,N_19501);
or UO_2132 (O_2132,N_19375,N_19720);
or UO_2133 (O_2133,N_19473,N_19798);
nor UO_2134 (O_2134,N_19031,N_19654);
and UO_2135 (O_2135,N_19816,N_19294);
nand UO_2136 (O_2136,N_19223,N_19836);
and UO_2137 (O_2137,N_19107,N_19169);
or UO_2138 (O_2138,N_19145,N_19342);
or UO_2139 (O_2139,N_19211,N_19900);
and UO_2140 (O_2140,N_19105,N_19804);
or UO_2141 (O_2141,N_19926,N_19925);
and UO_2142 (O_2142,N_19234,N_19682);
and UO_2143 (O_2143,N_19252,N_19059);
and UO_2144 (O_2144,N_19744,N_19908);
nand UO_2145 (O_2145,N_19840,N_19045);
or UO_2146 (O_2146,N_19441,N_19535);
nor UO_2147 (O_2147,N_19828,N_19243);
or UO_2148 (O_2148,N_19445,N_19590);
and UO_2149 (O_2149,N_19405,N_19657);
or UO_2150 (O_2150,N_19364,N_19949);
and UO_2151 (O_2151,N_19300,N_19889);
and UO_2152 (O_2152,N_19937,N_19006);
and UO_2153 (O_2153,N_19074,N_19241);
nor UO_2154 (O_2154,N_19411,N_19451);
and UO_2155 (O_2155,N_19107,N_19152);
or UO_2156 (O_2156,N_19973,N_19778);
and UO_2157 (O_2157,N_19310,N_19044);
nand UO_2158 (O_2158,N_19386,N_19444);
and UO_2159 (O_2159,N_19210,N_19880);
xnor UO_2160 (O_2160,N_19199,N_19338);
nand UO_2161 (O_2161,N_19878,N_19845);
nand UO_2162 (O_2162,N_19486,N_19232);
xor UO_2163 (O_2163,N_19663,N_19739);
nor UO_2164 (O_2164,N_19071,N_19687);
xor UO_2165 (O_2165,N_19378,N_19744);
nand UO_2166 (O_2166,N_19232,N_19255);
or UO_2167 (O_2167,N_19298,N_19797);
nand UO_2168 (O_2168,N_19733,N_19149);
nor UO_2169 (O_2169,N_19558,N_19783);
or UO_2170 (O_2170,N_19840,N_19203);
xor UO_2171 (O_2171,N_19348,N_19846);
or UO_2172 (O_2172,N_19697,N_19938);
and UO_2173 (O_2173,N_19834,N_19074);
xnor UO_2174 (O_2174,N_19538,N_19689);
xnor UO_2175 (O_2175,N_19402,N_19756);
or UO_2176 (O_2176,N_19825,N_19319);
xnor UO_2177 (O_2177,N_19664,N_19532);
nand UO_2178 (O_2178,N_19237,N_19995);
nor UO_2179 (O_2179,N_19785,N_19224);
and UO_2180 (O_2180,N_19793,N_19337);
or UO_2181 (O_2181,N_19649,N_19907);
nor UO_2182 (O_2182,N_19266,N_19309);
or UO_2183 (O_2183,N_19964,N_19140);
or UO_2184 (O_2184,N_19688,N_19813);
nand UO_2185 (O_2185,N_19749,N_19709);
and UO_2186 (O_2186,N_19125,N_19127);
nor UO_2187 (O_2187,N_19471,N_19752);
nand UO_2188 (O_2188,N_19075,N_19485);
or UO_2189 (O_2189,N_19573,N_19680);
nor UO_2190 (O_2190,N_19658,N_19895);
xor UO_2191 (O_2191,N_19466,N_19225);
nor UO_2192 (O_2192,N_19937,N_19988);
or UO_2193 (O_2193,N_19220,N_19271);
xnor UO_2194 (O_2194,N_19964,N_19379);
and UO_2195 (O_2195,N_19245,N_19548);
nand UO_2196 (O_2196,N_19561,N_19489);
nand UO_2197 (O_2197,N_19188,N_19961);
or UO_2198 (O_2198,N_19206,N_19651);
nor UO_2199 (O_2199,N_19479,N_19213);
and UO_2200 (O_2200,N_19147,N_19145);
and UO_2201 (O_2201,N_19760,N_19016);
xnor UO_2202 (O_2202,N_19835,N_19999);
and UO_2203 (O_2203,N_19123,N_19037);
nand UO_2204 (O_2204,N_19282,N_19739);
nor UO_2205 (O_2205,N_19115,N_19904);
nand UO_2206 (O_2206,N_19871,N_19382);
xor UO_2207 (O_2207,N_19041,N_19934);
and UO_2208 (O_2208,N_19612,N_19721);
and UO_2209 (O_2209,N_19219,N_19389);
and UO_2210 (O_2210,N_19705,N_19339);
and UO_2211 (O_2211,N_19890,N_19359);
xor UO_2212 (O_2212,N_19927,N_19163);
and UO_2213 (O_2213,N_19467,N_19089);
and UO_2214 (O_2214,N_19758,N_19857);
and UO_2215 (O_2215,N_19929,N_19808);
xnor UO_2216 (O_2216,N_19083,N_19220);
xnor UO_2217 (O_2217,N_19508,N_19753);
xor UO_2218 (O_2218,N_19079,N_19571);
nand UO_2219 (O_2219,N_19469,N_19555);
nand UO_2220 (O_2220,N_19644,N_19077);
nand UO_2221 (O_2221,N_19097,N_19630);
xnor UO_2222 (O_2222,N_19483,N_19200);
xor UO_2223 (O_2223,N_19291,N_19916);
nand UO_2224 (O_2224,N_19108,N_19034);
or UO_2225 (O_2225,N_19842,N_19773);
nor UO_2226 (O_2226,N_19942,N_19224);
or UO_2227 (O_2227,N_19232,N_19897);
nand UO_2228 (O_2228,N_19055,N_19839);
or UO_2229 (O_2229,N_19799,N_19585);
or UO_2230 (O_2230,N_19646,N_19682);
xnor UO_2231 (O_2231,N_19834,N_19211);
xnor UO_2232 (O_2232,N_19981,N_19039);
and UO_2233 (O_2233,N_19487,N_19267);
nor UO_2234 (O_2234,N_19622,N_19604);
or UO_2235 (O_2235,N_19539,N_19677);
xnor UO_2236 (O_2236,N_19683,N_19789);
and UO_2237 (O_2237,N_19080,N_19015);
nor UO_2238 (O_2238,N_19099,N_19535);
nor UO_2239 (O_2239,N_19408,N_19058);
or UO_2240 (O_2240,N_19024,N_19332);
nor UO_2241 (O_2241,N_19852,N_19034);
xnor UO_2242 (O_2242,N_19656,N_19641);
and UO_2243 (O_2243,N_19405,N_19134);
xor UO_2244 (O_2244,N_19031,N_19205);
nand UO_2245 (O_2245,N_19909,N_19227);
or UO_2246 (O_2246,N_19727,N_19550);
xnor UO_2247 (O_2247,N_19136,N_19378);
or UO_2248 (O_2248,N_19499,N_19757);
nand UO_2249 (O_2249,N_19714,N_19993);
nand UO_2250 (O_2250,N_19687,N_19156);
and UO_2251 (O_2251,N_19931,N_19073);
nor UO_2252 (O_2252,N_19336,N_19535);
or UO_2253 (O_2253,N_19923,N_19481);
nor UO_2254 (O_2254,N_19892,N_19070);
nand UO_2255 (O_2255,N_19804,N_19731);
nor UO_2256 (O_2256,N_19732,N_19632);
and UO_2257 (O_2257,N_19502,N_19126);
nand UO_2258 (O_2258,N_19969,N_19546);
xor UO_2259 (O_2259,N_19415,N_19728);
xnor UO_2260 (O_2260,N_19519,N_19654);
nor UO_2261 (O_2261,N_19754,N_19469);
or UO_2262 (O_2262,N_19455,N_19532);
and UO_2263 (O_2263,N_19400,N_19080);
and UO_2264 (O_2264,N_19753,N_19619);
xnor UO_2265 (O_2265,N_19658,N_19527);
nor UO_2266 (O_2266,N_19255,N_19713);
nand UO_2267 (O_2267,N_19860,N_19020);
xnor UO_2268 (O_2268,N_19743,N_19150);
and UO_2269 (O_2269,N_19875,N_19479);
and UO_2270 (O_2270,N_19582,N_19592);
and UO_2271 (O_2271,N_19527,N_19624);
or UO_2272 (O_2272,N_19761,N_19057);
and UO_2273 (O_2273,N_19653,N_19749);
nand UO_2274 (O_2274,N_19777,N_19056);
nor UO_2275 (O_2275,N_19029,N_19641);
and UO_2276 (O_2276,N_19917,N_19320);
or UO_2277 (O_2277,N_19830,N_19491);
or UO_2278 (O_2278,N_19688,N_19290);
xnor UO_2279 (O_2279,N_19904,N_19694);
xnor UO_2280 (O_2280,N_19565,N_19121);
nor UO_2281 (O_2281,N_19255,N_19484);
or UO_2282 (O_2282,N_19412,N_19693);
and UO_2283 (O_2283,N_19901,N_19955);
or UO_2284 (O_2284,N_19053,N_19388);
and UO_2285 (O_2285,N_19494,N_19487);
nor UO_2286 (O_2286,N_19767,N_19237);
nand UO_2287 (O_2287,N_19787,N_19231);
nor UO_2288 (O_2288,N_19953,N_19820);
xnor UO_2289 (O_2289,N_19308,N_19550);
or UO_2290 (O_2290,N_19961,N_19166);
and UO_2291 (O_2291,N_19976,N_19491);
nor UO_2292 (O_2292,N_19228,N_19668);
xnor UO_2293 (O_2293,N_19870,N_19373);
nand UO_2294 (O_2294,N_19788,N_19760);
nor UO_2295 (O_2295,N_19844,N_19267);
xnor UO_2296 (O_2296,N_19544,N_19351);
or UO_2297 (O_2297,N_19414,N_19429);
nand UO_2298 (O_2298,N_19159,N_19488);
nand UO_2299 (O_2299,N_19251,N_19764);
and UO_2300 (O_2300,N_19012,N_19266);
nand UO_2301 (O_2301,N_19136,N_19982);
nand UO_2302 (O_2302,N_19158,N_19877);
nor UO_2303 (O_2303,N_19137,N_19433);
or UO_2304 (O_2304,N_19381,N_19102);
or UO_2305 (O_2305,N_19581,N_19547);
nor UO_2306 (O_2306,N_19389,N_19466);
xor UO_2307 (O_2307,N_19974,N_19796);
or UO_2308 (O_2308,N_19213,N_19648);
nor UO_2309 (O_2309,N_19647,N_19202);
nand UO_2310 (O_2310,N_19089,N_19204);
and UO_2311 (O_2311,N_19056,N_19424);
nand UO_2312 (O_2312,N_19696,N_19117);
and UO_2313 (O_2313,N_19308,N_19219);
xor UO_2314 (O_2314,N_19390,N_19344);
xor UO_2315 (O_2315,N_19167,N_19699);
nor UO_2316 (O_2316,N_19886,N_19907);
xor UO_2317 (O_2317,N_19591,N_19108);
or UO_2318 (O_2318,N_19128,N_19150);
and UO_2319 (O_2319,N_19190,N_19373);
nand UO_2320 (O_2320,N_19560,N_19520);
or UO_2321 (O_2321,N_19562,N_19853);
xor UO_2322 (O_2322,N_19098,N_19905);
and UO_2323 (O_2323,N_19256,N_19939);
nand UO_2324 (O_2324,N_19457,N_19736);
or UO_2325 (O_2325,N_19129,N_19802);
xor UO_2326 (O_2326,N_19560,N_19105);
nor UO_2327 (O_2327,N_19495,N_19121);
and UO_2328 (O_2328,N_19831,N_19359);
and UO_2329 (O_2329,N_19766,N_19703);
xor UO_2330 (O_2330,N_19839,N_19220);
nor UO_2331 (O_2331,N_19648,N_19176);
and UO_2332 (O_2332,N_19275,N_19947);
nand UO_2333 (O_2333,N_19559,N_19201);
and UO_2334 (O_2334,N_19886,N_19044);
nand UO_2335 (O_2335,N_19255,N_19975);
nand UO_2336 (O_2336,N_19750,N_19307);
xnor UO_2337 (O_2337,N_19395,N_19729);
xor UO_2338 (O_2338,N_19466,N_19625);
nor UO_2339 (O_2339,N_19715,N_19900);
or UO_2340 (O_2340,N_19232,N_19099);
xnor UO_2341 (O_2341,N_19221,N_19467);
nor UO_2342 (O_2342,N_19624,N_19239);
nor UO_2343 (O_2343,N_19139,N_19753);
nor UO_2344 (O_2344,N_19891,N_19776);
xor UO_2345 (O_2345,N_19867,N_19835);
and UO_2346 (O_2346,N_19588,N_19143);
nand UO_2347 (O_2347,N_19264,N_19147);
nor UO_2348 (O_2348,N_19522,N_19839);
or UO_2349 (O_2349,N_19743,N_19405);
xor UO_2350 (O_2350,N_19472,N_19000);
nor UO_2351 (O_2351,N_19190,N_19793);
xor UO_2352 (O_2352,N_19044,N_19781);
nand UO_2353 (O_2353,N_19722,N_19449);
xnor UO_2354 (O_2354,N_19963,N_19147);
and UO_2355 (O_2355,N_19687,N_19083);
xor UO_2356 (O_2356,N_19647,N_19181);
nand UO_2357 (O_2357,N_19606,N_19890);
and UO_2358 (O_2358,N_19541,N_19656);
or UO_2359 (O_2359,N_19211,N_19341);
and UO_2360 (O_2360,N_19567,N_19729);
nand UO_2361 (O_2361,N_19384,N_19623);
or UO_2362 (O_2362,N_19200,N_19283);
nand UO_2363 (O_2363,N_19961,N_19874);
xor UO_2364 (O_2364,N_19070,N_19115);
or UO_2365 (O_2365,N_19597,N_19270);
or UO_2366 (O_2366,N_19693,N_19649);
or UO_2367 (O_2367,N_19257,N_19600);
and UO_2368 (O_2368,N_19854,N_19975);
xor UO_2369 (O_2369,N_19101,N_19380);
nand UO_2370 (O_2370,N_19567,N_19783);
nand UO_2371 (O_2371,N_19044,N_19980);
and UO_2372 (O_2372,N_19634,N_19066);
and UO_2373 (O_2373,N_19773,N_19839);
and UO_2374 (O_2374,N_19078,N_19365);
or UO_2375 (O_2375,N_19188,N_19706);
nor UO_2376 (O_2376,N_19274,N_19004);
xnor UO_2377 (O_2377,N_19827,N_19516);
nand UO_2378 (O_2378,N_19568,N_19730);
and UO_2379 (O_2379,N_19099,N_19312);
or UO_2380 (O_2380,N_19608,N_19727);
or UO_2381 (O_2381,N_19366,N_19995);
nor UO_2382 (O_2382,N_19916,N_19333);
nand UO_2383 (O_2383,N_19494,N_19263);
or UO_2384 (O_2384,N_19676,N_19321);
nand UO_2385 (O_2385,N_19033,N_19183);
nand UO_2386 (O_2386,N_19973,N_19538);
and UO_2387 (O_2387,N_19981,N_19891);
nand UO_2388 (O_2388,N_19066,N_19172);
xor UO_2389 (O_2389,N_19675,N_19594);
nand UO_2390 (O_2390,N_19168,N_19225);
nor UO_2391 (O_2391,N_19006,N_19445);
nor UO_2392 (O_2392,N_19096,N_19812);
nor UO_2393 (O_2393,N_19652,N_19890);
nor UO_2394 (O_2394,N_19955,N_19704);
xor UO_2395 (O_2395,N_19717,N_19820);
nand UO_2396 (O_2396,N_19141,N_19288);
nand UO_2397 (O_2397,N_19673,N_19862);
or UO_2398 (O_2398,N_19787,N_19430);
and UO_2399 (O_2399,N_19442,N_19150);
nand UO_2400 (O_2400,N_19812,N_19844);
and UO_2401 (O_2401,N_19497,N_19045);
xnor UO_2402 (O_2402,N_19530,N_19930);
nor UO_2403 (O_2403,N_19650,N_19135);
or UO_2404 (O_2404,N_19996,N_19313);
xor UO_2405 (O_2405,N_19900,N_19076);
nand UO_2406 (O_2406,N_19384,N_19767);
xnor UO_2407 (O_2407,N_19964,N_19541);
nor UO_2408 (O_2408,N_19312,N_19910);
and UO_2409 (O_2409,N_19307,N_19491);
or UO_2410 (O_2410,N_19879,N_19009);
nor UO_2411 (O_2411,N_19117,N_19721);
nor UO_2412 (O_2412,N_19864,N_19382);
and UO_2413 (O_2413,N_19469,N_19812);
nand UO_2414 (O_2414,N_19279,N_19426);
nor UO_2415 (O_2415,N_19916,N_19536);
nor UO_2416 (O_2416,N_19959,N_19490);
or UO_2417 (O_2417,N_19673,N_19336);
or UO_2418 (O_2418,N_19599,N_19249);
xnor UO_2419 (O_2419,N_19895,N_19235);
or UO_2420 (O_2420,N_19975,N_19034);
or UO_2421 (O_2421,N_19268,N_19185);
or UO_2422 (O_2422,N_19568,N_19613);
or UO_2423 (O_2423,N_19152,N_19350);
nand UO_2424 (O_2424,N_19053,N_19243);
or UO_2425 (O_2425,N_19174,N_19413);
xnor UO_2426 (O_2426,N_19303,N_19712);
nand UO_2427 (O_2427,N_19670,N_19222);
nand UO_2428 (O_2428,N_19679,N_19357);
and UO_2429 (O_2429,N_19997,N_19149);
xor UO_2430 (O_2430,N_19991,N_19006);
xnor UO_2431 (O_2431,N_19365,N_19410);
nand UO_2432 (O_2432,N_19809,N_19063);
nand UO_2433 (O_2433,N_19587,N_19484);
or UO_2434 (O_2434,N_19369,N_19374);
nand UO_2435 (O_2435,N_19909,N_19489);
and UO_2436 (O_2436,N_19979,N_19971);
xor UO_2437 (O_2437,N_19971,N_19362);
nand UO_2438 (O_2438,N_19698,N_19733);
xor UO_2439 (O_2439,N_19298,N_19951);
and UO_2440 (O_2440,N_19077,N_19346);
xnor UO_2441 (O_2441,N_19545,N_19233);
and UO_2442 (O_2442,N_19715,N_19242);
xor UO_2443 (O_2443,N_19529,N_19948);
and UO_2444 (O_2444,N_19116,N_19843);
nor UO_2445 (O_2445,N_19365,N_19543);
nand UO_2446 (O_2446,N_19678,N_19212);
nand UO_2447 (O_2447,N_19515,N_19336);
nor UO_2448 (O_2448,N_19987,N_19210);
and UO_2449 (O_2449,N_19567,N_19424);
nand UO_2450 (O_2450,N_19614,N_19476);
xor UO_2451 (O_2451,N_19414,N_19283);
or UO_2452 (O_2452,N_19750,N_19014);
or UO_2453 (O_2453,N_19449,N_19702);
nor UO_2454 (O_2454,N_19235,N_19693);
nor UO_2455 (O_2455,N_19199,N_19258);
nand UO_2456 (O_2456,N_19000,N_19030);
nand UO_2457 (O_2457,N_19886,N_19442);
or UO_2458 (O_2458,N_19699,N_19387);
and UO_2459 (O_2459,N_19087,N_19387);
nor UO_2460 (O_2460,N_19941,N_19993);
nor UO_2461 (O_2461,N_19311,N_19355);
and UO_2462 (O_2462,N_19225,N_19817);
and UO_2463 (O_2463,N_19943,N_19891);
nand UO_2464 (O_2464,N_19613,N_19081);
or UO_2465 (O_2465,N_19213,N_19813);
nand UO_2466 (O_2466,N_19485,N_19575);
xor UO_2467 (O_2467,N_19346,N_19764);
or UO_2468 (O_2468,N_19777,N_19927);
and UO_2469 (O_2469,N_19534,N_19529);
nor UO_2470 (O_2470,N_19120,N_19935);
or UO_2471 (O_2471,N_19580,N_19073);
xnor UO_2472 (O_2472,N_19838,N_19436);
xnor UO_2473 (O_2473,N_19813,N_19391);
nor UO_2474 (O_2474,N_19356,N_19938);
nor UO_2475 (O_2475,N_19100,N_19156);
and UO_2476 (O_2476,N_19740,N_19847);
or UO_2477 (O_2477,N_19893,N_19384);
nor UO_2478 (O_2478,N_19382,N_19919);
nor UO_2479 (O_2479,N_19731,N_19892);
xnor UO_2480 (O_2480,N_19128,N_19175);
nand UO_2481 (O_2481,N_19786,N_19795);
xor UO_2482 (O_2482,N_19816,N_19408);
nand UO_2483 (O_2483,N_19514,N_19819);
xor UO_2484 (O_2484,N_19976,N_19636);
nand UO_2485 (O_2485,N_19614,N_19475);
xor UO_2486 (O_2486,N_19170,N_19466);
nand UO_2487 (O_2487,N_19727,N_19823);
nand UO_2488 (O_2488,N_19770,N_19449);
or UO_2489 (O_2489,N_19462,N_19828);
or UO_2490 (O_2490,N_19292,N_19286);
and UO_2491 (O_2491,N_19976,N_19540);
nor UO_2492 (O_2492,N_19127,N_19750);
nor UO_2493 (O_2493,N_19155,N_19956);
xor UO_2494 (O_2494,N_19098,N_19896);
nor UO_2495 (O_2495,N_19318,N_19364);
xor UO_2496 (O_2496,N_19113,N_19691);
xor UO_2497 (O_2497,N_19849,N_19105);
xor UO_2498 (O_2498,N_19896,N_19872);
xnor UO_2499 (O_2499,N_19737,N_19584);
endmodule