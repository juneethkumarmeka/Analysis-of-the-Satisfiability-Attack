module basic_2500_25000_3000_8_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
xor U0 (N_0,In_2005,In_1646);
nor U1 (N_1,In_1345,In_860);
xor U2 (N_2,In_1248,In_2245);
xnor U3 (N_3,In_1264,In_2289);
nand U4 (N_4,In_1288,In_971);
and U5 (N_5,In_2096,In_1903);
nor U6 (N_6,In_1647,In_870);
or U7 (N_7,In_684,In_1204);
nand U8 (N_8,In_425,In_1403);
and U9 (N_9,In_752,In_168);
nor U10 (N_10,In_667,In_743);
or U11 (N_11,In_1486,In_337);
nand U12 (N_12,In_138,In_145);
or U13 (N_13,In_915,In_2380);
xnor U14 (N_14,In_2423,In_243);
or U15 (N_15,In_569,In_783);
and U16 (N_16,In_2435,In_744);
xnor U17 (N_17,In_836,In_1103);
and U18 (N_18,In_1769,In_1088);
nand U19 (N_19,In_375,In_2480);
and U20 (N_20,In_906,In_115);
xnor U21 (N_21,In_1621,In_1377);
and U22 (N_22,In_705,In_938);
or U23 (N_23,In_1851,In_1032);
xor U24 (N_24,In_1447,In_703);
xnor U25 (N_25,In_2071,In_1161);
and U26 (N_26,In_294,In_1073);
nand U27 (N_27,In_355,In_1152);
or U28 (N_28,In_1594,In_1808);
nor U29 (N_29,In_1240,In_1316);
and U30 (N_30,In_1538,In_348);
and U31 (N_31,In_873,In_704);
nor U32 (N_32,In_1816,In_741);
xnor U33 (N_33,In_1572,In_2156);
xnor U34 (N_34,In_2193,In_366);
xnor U35 (N_35,In_600,In_2291);
or U36 (N_36,In_1492,In_940);
and U37 (N_37,In_1253,In_680);
nor U38 (N_38,In_1059,In_1221);
or U39 (N_39,In_791,In_211);
or U40 (N_40,In_1443,In_2276);
or U41 (N_41,In_968,In_245);
nor U42 (N_42,In_1626,In_112);
and U43 (N_43,In_1305,In_2161);
and U44 (N_44,In_2269,In_1975);
nand U45 (N_45,In_2310,In_332);
nand U46 (N_46,In_2229,In_2349);
nand U47 (N_47,In_2141,In_1746);
nor U48 (N_48,In_1219,In_660);
xor U49 (N_49,In_86,In_444);
nor U50 (N_50,In_160,In_1148);
xnor U51 (N_51,In_577,In_333);
nand U52 (N_52,In_161,In_402);
or U53 (N_53,In_963,In_874);
nor U54 (N_54,In_338,In_946);
or U55 (N_55,In_1418,In_351);
and U56 (N_56,In_1990,In_2);
nor U57 (N_57,In_1434,In_1295);
xor U58 (N_58,In_169,In_2208);
and U59 (N_59,In_345,In_1153);
nor U60 (N_60,In_1213,In_1757);
nor U61 (N_61,In_397,In_1733);
and U62 (N_62,In_1593,In_1158);
nor U63 (N_63,In_923,In_682);
xor U64 (N_64,In_730,In_507);
and U65 (N_65,In_1765,In_1795);
nor U66 (N_66,In_1421,In_1337);
nand U67 (N_67,In_1832,In_1179);
xor U68 (N_68,In_742,In_2397);
and U69 (N_69,In_1883,In_1466);
or U70 (N_70,In_64,In_2183);
nand U71 (N_71,In_573,In_1802);
and U72 (N_72,In_532,In_1748);
or U73 (N_73,In_1869,In_1672);
and U74 (N_74,In_2084,In_1237);
and U75 (N_75,In_1653,In_1732);
and U76 (N_76,In_1373,In_1215);
nand U77 (N_77,In_369,In_1102);
nor U78 (N_78,In_2032,In_2317);
nand U79 (N_79,In_346,In_620);
nor U80 (N_80,In_1125,In_1112);
and U81 (N_81,In_2260,In_256);
and U82 (N_82,In_1984,In_2469);
nor U83 (N_83,In_1871,In_624);
nand U84 (N_84,In_719,In_1028);
or U85 (N_85,In_598,In_1035);
xor U86 (N_86,In_1521,In_962);
nand U87 (N_87,In_371,In_1674);
and U88 (N_88,In_238,In_1796);
nand U89 (N_89,In_150,In_2266);
nand U90 (N_90,In_1624,In_1906);
and U91 (N_91,In_526,In_392);
or U92 (N_92,In_651,In_1986);
nand U93 (N_93,In_608,In_480);
nor U94 (N_94,In_972,In_307);
and U95 (N_95,In_1806,In_258);
xnor U96 (N_96,In_1685,In_988);
and U97 (N_97,In_1114,In_1864);
or U98 (N_98,In_415,In_90);
and U99 (N_99,In_534,In_39);
or U100 (N_100,In_776,In_30);
xnor U101 (N_101,In_1529,In_996);
xnor U102 (N_102,In_2297,In_517);
nand U103 (N_103,In_1056,In_1319);
nand U104 (N_104,In_678,In_1657);
and U105 (N_105,In_2192,In_2267);
or U106 (N_106,In_1634,In_297);
nand U107 (N_107,In_565,In_62);
and U108 (N_108,In_913,In_622);
nor U109 (N_109,In_875,In_77);
or U110 (N_110,In_716,In_1972);
and U111 (N_111,In_840,In_1294);
nor U112 (N_112,In_1923,In_357);
or U113 (N_113,In_1696,In_1049);
nor U114 (N_114,In_897,In_1242);
xor U115 (N_115,In_2130,In_553);
nor U116 (N_116,In_1914,In_949);
and U117 (N_117,In_2366,In_945);
nand U118 (N_118,In_961,In_1278);
nand U119 (N_119,In_1321,In_2172);
or U120 (N_120,In_1489,In_1054);
and U121 (N_121,In_1362,In_2114);
nand U122 (N_122,In_1884,In_1484);
or U123 (N_123,In_203,In_1519);
and U124 (N_124,In_769,In_74);
nor U125 (N_125,In_125,In_1145);
or U126 (N_126,In_1544,In_457);
and U127 (N_127,In_1605,In_802);
nor U128 (N_128,In_1235,In_2036);
nand U129 (N_129,In_723,In_2018);
nand U130 (N_130,In_95,In_1710);
or U131 (N_131,In_1252,In_1222);
xnor U132 (N_132,In_1353,In_811);
xor U133 (N_133,In_1055,In_126);
and U134 (N_134,In_685,In_2122);
xnor U135 (N_135,In_1239,In_134);
nor U136 (N_136,In_489,In_1488);
nor U137 (N_137,In_1867,In_388);
or U138 (N_138,In_2424,In_2217);
or U139 (N_139,In_1142,In_649);
xnor U140 (N_140,In_433,In_2418);
xor U141 (N_141,In_1351,In_310);
and U142 (N_142,In_1042,In_1683);
xor U143 (N_143,In_1854,In_37);
and U144 (N_144,In_772,In_1981);
xnor U145 (N_145,In_1899,In_1428);
xor U146 (N_146,In_1960,In_855);
and U147 (N_147,In_2097,In_352);
xnor U148 (N_148,In_326,In_1737);
nor U149 (N_149,In_379,In_473);
nor U150 (N_150,In_1614,In_656);
or U151 (N_151,In_1013,In_2497);
and U152 (N_152,In_560,In_2187);
nor U153 (N_153,In_623,In_225);
xor U154 (N_154,In_1458,In_826);
nand U155 (N_155,In_885,In_314);
xor U156 (N_156,In_2033,In_277);
nand U157 (N_157,In_2194,In_676);
and U158 (N_158,In_627,In_136);
nor U159 (N_159,In_2292,In_1812);
and U160 (N_160,In_1731,In_468);
nand U161 (N_161,In_2109,In_774);
nor U162 (N_162,In_985,In_1713);
nand U163 (N_163,In_2155,In_2102);
and U164 (N_164,In_775,In_2198);
nor U165 (N_165,In_1437,In_2024);
or U166 (N_166,In_1568,In_202);
or U167 (N_167,In_2386,In_148);
nor U168 (N_168,In_761,In_1740);
nor U169 (N_169,In_2359,In_2333);
or U170 (N_170,In_2439,In_1781);
xnor U171 (N_171,In_852,In_1875);
and U172 (N_172,In_91,In_2414);
nand U173 (N_173,In_699,In_274);
or U174 (N_174,In_2206,In_1452);
nor U175 (N_175,In_1279,In_308);
xnor U176 (N_176,In_1936,In_470);
nor U177 (N_177,In_872,In_683);
or U178 (N_178,In_1645,In_1904);
and U179 (N_179,In_1131,In_982);
xnor U180 (N_180,In_531,In_2280);
xnor U181 (N_181,In_2026,In_59);
nand U182 (N_182,In_2288,In_1225);
nand U183 (N_183,In_666,In_34);
xor U184 (N_184,In_1128,In_1394);
and U185 (N_185,In_1885,In_389);
nor U186 (N_186,In_2093,In_149);
nor U187 (N_187,In_1172,In_2107);
or U188 (N_188,In_1790,In_1756);
or U189 (N_189,In_548,In_19);
nand U190 (N_190,In_459,In_1971);
and U191 (N_191,In_1217,In_2105);
xor U192 (N_192,In_530,In_1108);
nor U193 (N_193,In_2283,In_2474);
xnor U194 (N_194,In_2328,In_143);
nor U195 (N_195,In_1119,In_32);
nor U196 (N_196,In_993,In_861);
nor U197 (N_197,In_1251,In_135);
xnor U198 (N_198,In_1214,In_2143);
or U199 (N_199,In_1075,In_48);
xor U200 (N_200,In_173,In_1202);
nand U201 (N_201,In_1203,In_1993);
and U202 (N_202,In_1697,In_267);
nand U203 (N_203,In_2368,In_1775);
nand U204 (N_204,In_2204,In_1389);
xnor U205 (N_205,In_1630,In_1040);
nand U206 (N_206,In_1270,In_157);
nand U207 (N_207,In_639,In_215);
nand U208 (N_208,In_2309,In_606);
nand U209 (N_209,In_2028,In_268);
xor U210 (N_210,In_2274,In_970);
or U211 (N_211,In_1123,In_2210);
or U212 (N_212,In_2466,In_1773);
and U213 (N_213,In_2235,In_163);
or U214 (N_214,In_1510,In_2484);
xnor U215 (N_215,In_103,In_2056);
or U216 (N_216,In_427,In_794);
nand U217 (N_217,In_1706,In_190);
xnor U218 (N_218,In_728,In_1965);
nor U219 (N_219,In_401,In_732);
and U220 (N_220,In_1818,In_2050);
xnor U221 (N_221,In_374,In_1335);
nor U222 (N_222,In_919,In_1589);
or U223 (N_223,In_1845,In_284);
or U224 (N_224,In_1648,In_1004);
nor U225 (N_225,In_2383,In_1226);
nand U226 (N_226,In_543,In_814);
xor U227 (N_227,In_803,In_1949);
and U228 (N_228,In_564,In_165);
xnor U229 (N_229,In_386,In_650);
or U230 (N_230,In_2181,In_1760);
or U231 (N_231,In_572,In_692);
or U232 (N_232,In_1552,In_408);
and U233 (N_233,In_2408,In_898);
or U234 (N_234,In_780,In_1664);
nor U235 (N_235,In_833,In_1220);
or U236 (N_236,In_1528,In_1018);
and U237 (N_237,In_674,In_1243);
or U238 (N_238,In_856,In_465);
or U239 (N_239,In_1411,In_1537);
or U240 (N_240,In_986,In_1363);
nand U241 (N_241,In_1536,In_954);
and U242 (N_242,In_2174,In_479);
and U243 (N_243,In_1559,In_264);
nor U244 (N_244,In_2259,In_2016);
or U245 (N_245,In_197,In_756);
nor U246 (N_246,In_1768,In_1491);
xor U247 (N_247,In_464,In_2158);
xor U248 (N_248,In_2085,In_1482);
nand U249 (N_249,In_1878,In_2293);
xor U250 (N_250,In_935,In_147);
xnor U251 (N_251,In_1038,In_1586);
xor U252 (N_252,In_411,In_2008);
and U253 (N_253,In_2341,In_1450);
and U254 (N_254,In_1750,In_1763);
nand U255 (N_255,In_1066,In_194);
nor U256 (N_256,In_1419,In_1563);
nand U257 (N_257,In_475,In_1144);
xor U258 (N_258,In_488,In_2263);
nand U259 (N_259,In_2479,In_551);
xor U260 (N_260,In_1606,In_1620);
and U261 (N_261,In_1957,In_429);
nor U262 (N_262,In_1725,In_1406);
nand U263 (N_263,In_2092,In_1346);
nand U264 (N_264,In_1498,In_10);
xor U265 (N_265,In_1177,In_370);
and U266 (N_266,In_2055,In_1192);
xnor U267 (N_267,In_1456,In_1550);
nand U268 (N_268,In_485,In_504);
nor U269 (N_269,In_1314,In_2299);
or U270 (N_270,In_1897,In_2154);
nand U271 (N_271,In_178,In_325);
or U272 (N_272,In_1942,In_1716);
nor U273 (N_273,In_1116,In_1472);
and U274 (N_274,In_2118,In_80);
xnor U275 (N_275,In_1539,In_1205);
xor U276 (N_276,In_2081,In_1069);
or U277 (N_277,In_854,In_1663);
and U278 (N_278,In_377,In_2087);
or U279 (N_279,In_2251,In_463);
nand U280 (N_280,In_2099,In_394);
nand U281 (N_281,In_361,In_96);
and U282 (N_282,In_1186,In_1931);
xnor U283 (N_283,In_2040,In_722);
nand U284 (N_284,In_2072,In_1771);
nand U285 (N_285,In_2275,In_1627);
nand U286 (N_286,In_1497,In_2391);
xor U287 (N_287,In_1755,In_2031);
xor U288 (N_288,In_35,In_1613);
xnor U289 (N_289,In_269,In_196);
nor U290 (N_290,In_304,In_1920);
nor U291 (N_291,In_79,In_98);
nand U292 (N_292,In_525,In_94);
xor U293 (N_293,In_120,In_983);
nor U294 (N_294,In_55,In_24);
or U295 (N_295,In_367,In_1064);
and U296 (N_296,In_438,In_3);
and U297 (N_297,In_2231,In_285);
or U298 (N_298,In_1892,In_1228);
xor U299 (N_299,In_1231,In_220);
or U300 (N_300,In_12,In_1405);
or U301 (N_301,In_1670,In_1457);
nor U302 (N_302,In_2381,In_2074);
nand U303 (N_303,In_2134,In_1797);
and U304 (N_304,In_275,In_450);
xnor U305 (N_305,In_1284,In_2488);
nor U306 (N_306,In_812,In_449);
or U307 (N_307,In_2436,In_767);
nor U308 (N_308,In_601,In_492);
xor U309 (N_309,In_1978,In_440);
xnor U310 (N_310,In_1465,In_907);
xnor U311 (N_311,In_1198,In_1595);
or U312 (N_312,In_579,In_4);
or U313 (N_313,In_439,In_1535);
xnor U314 (N_314,In_296,In_1842);
nor U315 (N_315,In_133,In_1794);
nor U316 (N_316,In_1005,In_524);
or U317 (N_317,In_186,In_1616);
or U318 (N_318,In_2468,In_1381);
nor U319 (N_319,In_528,In_430);
nand U320 (N_320,In_1293,In_2253);
or U321 (N_321,In_409,In_2401);
or U322 (N_322,In_960,In_629);
or U323 (N_323,In_259,In_626);
nor U324 (N_324,In_300,In_555);
or U325 (N_325,In_2052,In_1147);
and U326 (N_326,In_1666,In_97);
or U327 (N_327,In_476,In_632);
nor U328 (N_328,In_1318,In_1436);
xor U329 (N_329,In_2047,In_1197);
nor U330 (N_330,In_2116,In_2077);
or U331 (N_331,In_11,In_1622);
and U332 (N_332,In_2153,In_384);
or U333 (N_333,In_2473,In_410);
and U334 (N_334,In_21,In_1998);
and U335 (N_335,In_491,In_1749);
and U336 (N_336,In_1809,In_1302);
nand U337 (N_337,In_1860,In_1100);
nand U338 (N_338,In_2111,In_1992);
nand U339 (N_339,In_57,In_1598);
xnor U340 (N_340,In_942,In_434);
and U341 (N_341,In_1558,In_981);
nand U342 (N_342,In_1573,In_69);
nor U343 (N_343,In_956,In_2377);
xor U344 (N_344,In_2419,In_76);
xor U345 (N_345,In_1250,In_1890);
nor U346 (N_346,In_2409,In_2278);
or U347 (N_347,In_1615,In_844);
or U348 (N_348,In_1409,In_1009);
nor U349 (N_349,In_175,In_2321);
and U350 (N_350,In_1565,In_234);
and U351 (N_351,In_1888,In_85);
nand U352 (N_352,In_1227,In_317);
nand U353 (N_353,In_2449,In_92);
nor U354 (N_354,In_1777,In_1951);
nor U355 (N_355,In_7,In_1120);
xnor U356 (N_356,In_1868,In_928);
xnor U357 (N_357,In_25,In_1303);
and U358 (N_358,In_107,In_407);
or U359 (N_359,In_1926,In_733);
nand U360 (N_360,In_1174,In_1139);
and U361 (N_361,In_664,In_1045);
or U362 (N_362,In_1224,In_336);
xor U363 (N_363,In_1037,In_65);
xor U364 (N_364,In_246,In_2110);
xor U365 (N_365,In_460,In_817);
nor U366 (N_366,In_927,In_224);
or U367 (N_367,In_349,In_690);
xor U368 (N_368,In_1676,In_1358);
and U369 (N_369,In_1584,In_110);
or U370 (N_370,In_545,In_2443);
and U371 (N_371,In_414,In_1126);
xnor U372 (N_372,In_1862,In_1300);
and U373 (N_373,In_1404,In_1506);
nand U374 (N_374,In_869,In_1171);
or U375 (N_375,In_2205,In_2037);
or U376 (N_376,In_1199,In_1911);
or U377 (N_377,In_1829,In_689);
nand U378 (N_378,In_1308,In_1642);
nand U379 (N_379,In_240,In_1633);
xnor U380 (N_380,In_558,In_2164);
nor U381 (N_381,In_2338,In_201);
or U382 (N_382,In_755,In_2490);
and U383 (N_383,In_484,In_2442);
nand U384 (N_384,In_1822,In_795);
or U385 (N_385,In_1791,In_2195);
nand U386 (N_386,In_1933,In_1720);
xnor U387 (N_387,In_1977,In_1234);
or U388 (N_388,In_2002,In_2127);
or U389 (N_389,In_237,In_291);
and U390 (N_390,In_420,In_2207);
or U391 (N_391,In_2203,In_1785);
or U392 (N_392,In_2222,In_1130);
xnor U393 (N_393,In_2322,In_1701);
xnor U394 (N_394,In_342,In_1063);
or U395 (N_395,In_2133,In_887);
and U396 (N_396,In_2169,In_750);
and U397 (N_397,In_373,In_1833);
nor U398 (N_398,In_14,In_2382);
nand U399 (N_399,In_1813,In_2370);
and U400 (N_400,In_1591,In_700);
nand U401 (N_401,In_1574,In_857);
or U402 (N_402,In_890,In_2124);
nor U403 (N_403,In_2434,In_659);
and U404 (N_404,In_736,In_663);
nand U405 (N_405,In_806,In_2290);
or U406 (N_406,In_720,In_1527);
xor U407 (N_407,In_88,In_482);
nor U408 (N_408,In_951,In_105);
and U409 (N_409,In_1872,In_754);
nor U410 (N_410,In_1792,In_1208);
nor U411 (N_411,In_1087,In_762);
nand U412 (N_412,In_426,In_1093);
nand U413 (N_413,In_2398,In_2330);
and U414 (N_414,In_747,In_739);
and U415 (N_415,In_1863,In_1410);
nor U416 (N_416,In_209,In_254);
nand U417 (N_417,In_2249,In_1582);
xor U418 (N_418,In_1569,In_2219);
and U419 (N_419,In_1651,In_896);
or U420 (N_420,In_1764,In_1695);
and U421 (N_421,In_1612,In_1985);
nor U422 (N_422,In_2481,In_839);
nor U423 (N_423,In_512,In_2065);
nand U424 (N_424,In_1641,In_1398);
or U425 (N_425,In_1420,In_980);
nor U426 (N_426,In_937,In_1072);
or U427 (N_427,In_1354,In_1661);
nor U428 (N_428,In_15,In_1030);
and U429 (N_429,In_933,In_2117);
nor U430 (N_430,In_2277,In_2371);
xnor U431 (N_431,In_1415,In_745);
xnor U432 (N_432,In_1499,In_977);
nor U433 (N_433,In_538,In_283);
nand U434 (N_434,In_2350,In_1585);
xnor U435 (N_435,In_523,In_2302);
nor U436 (N_436,In_2363,In_2129);
or U437 (N_437,In_1638,In_1530);
nand U438 (N_438,In_289,In_1979);
or U439 (N_439,In_354,In_1124);
or U440 (N_440,In_1655,In_654);
nor U441 (N_441,In_1273,In_1392);
and U442 (N_442,In_2066,In_18);
xor U443 (N_443,In_1324,In_1579);
or U444 (N_444,In_195,In_1907);
xor U445 (N_445,In_1441,In_1372);
xor U446 (N_446,In_171,In_1094);
or U447 (N_447,In_1334,In_185);
nor U448 (N_448,In_1857,In_1068);
or U449 (N_449,In_1266,In_151);
and U450 (N_450,In_726,In_816);
nand U451 (N_451,In_2182,In_1508);
nand U452 (N_452,In_1079,In_156);
or U453 (N_453,In_453,In_158);
xor U454 (N_454,In_1083,In_1898);
and U455 (N_455,In_500,In_1438);
xnor U456 (N_456,In_541,In_1385);
nand U457 (N_457,In_1210,In_778);
and U458 (N_458,In_2175,In_2369);
or U459 (N_459,In_405,In_423);
and U460 (N_460,In_216,In_604);
or U461 (N_461,In_1060,In_693);
and U462 (N_462,In_454,In_1677);
or U463 (N_463,In_1592,In_1515);
nand U464 (N_464,In_1678,In_686);
and U465 (N_465,In_2335,In_1935);
xnor U466 (N_466,In_1330,In_2360);
nor U467 (N_467,In_698,In_1798);
nand U468 (N_468,In_1597,In_805);
nor U469 (N_469,In_422,In_2270);
and U470 (N_470,In_2459,In_1181);
nor U471 (N_471,In_2011,In_1136);
and U472 (N_472,In_1659,In_2021);
or U473 (N_473,In_497,In_1767);
or U474 (N_474,In_1257,In_1782);
xnor U475 (N_475,In_2426,In_2345);
nand U476 (N_476,In_1846,In_1039);
xor U477 (N_477,In_2445,In_226);
and U478 (N_478,In_2044,In_413);
nor U479 (N_479,In_2160,In_213);
or U480 (N_480,In_1386,In_1850);
xnor U481 (N_481,In_2104,In_735);
xor U482 (N_482,In_1912,In_1928);
nor U483 (N_483,In_1831,In_1290);
nor U484 (N_484,In_562,In_2342);
nor U485 (N_485,In_461,In_2347);
and U486 (N_486,In_669,In_1555);
and U487 (N_487,In_1910,In_2493);
nand U488 (N_488,In_1369,In_1950);
nand U489 (N_489,In_114,In_841);
or U490 (N_490,In_609,In_1588);
nand U491 (N_491,In_1,In_637);
xor U492 (N_492,In_2273,In_2250);
nand U493 (N_493,In_2010,In_1859);
xnor U494 (N_494,In_1715,In_1887);
nor U495 (N_495,In_1067,In_2168);
and U496 (N_496,In_571,In_1129);
xnor U497 (N_497,In_272,In_518);
and U498 (N_498,In_1717,In_2144);
nand U499 (N_499,In_1435,In_1604);
nor U500 (N_500,In_318,In_1400);
and U501 (N_501,In_1336,In_328);
nand U502 (N_502,In_1402,In_939);
and U503 (N_503,In_1417,In_758);
nand U504 (N_504,In_2471,In_1272);
nor U505 (N_505,In_1668,In_42);
xor U506 (N_506,In_0,In_286);
nand U507 (N_507,In_172,In_1522);
nand U508 (N_508,In_323,In_44);
nor U509 (N_509,In_1722,In_2049);
nor U510 (N_510,In_832,In_1448);
or U511 (N_511,In_2252,In_1397);
nand U512 (N_512,In_1459,In_1034);
nor U513 (N_513,In_2150,In_496);
or U514 (N_514,In_979,In_1804);
nand U515 (N_515,In_1766,In_1881);
nand U516 (N_516,In_672,In_2396);
xnor U517 (N_517,In_2390,In_1727);
nor U518 (N_518,In_2486,In_1339);
nor U519 (N_519,In_1311,In_1095);
and U520 (N_520,In_200,In_2025);
and U521 (N_521,In_987,In_2197);
and U522 (N_522,In_1444,In_909);
xor U523 (N_523,In_123,In_2112);
nor U524 (N_524,In_2413,In_712);
nor U525 (N_525,In_1044,In_1667);
nor U526 (N_526,In_152,In_1835);
or U527 (N_527,In_1033,In_1378);
nand U528 (N_528,In_1523,In_1654);
nand U529 (N_529,In_2073,In_729);
nand U530 (N_530,In_1602,In_603);
xnor U531 (N_531,In_1927,In_2325);
and U532 (N_532,In_2046,In_590);
nor U533 (N_533,In_1980,In_2220);
xnor U534 (N_534,In_1107,In_1274);
or U535 (N_535,In_1939,In_1724);
nand U536 (N_536,In_591,In_1455);
or U537 (N_537,In_1943,In_2315);
and U538 (N_538,In_1940,In_2076);
or U539 (N_539,In_20,In_193);
nand U540 (N_540,In_859,In_1163);
and U541 (N_541,In_490,In_49);
nor U542 (N_542,In_846,In_1006);
or U543 (N_543,In_1649,In_320);
and U544 (N_544,In_941,In_575);
nor U545 (N_545,In_1921,In_2137);
nand U546 (N_546,In_164,In_1296);
nand U547 (N_547,In_1090,In_1635);
nand U548 (N_548,In_1577,In_867);
nor U549 (N_549,In_1560,In_2454);
nand U550 (N_550,In_1629,In_2147);
xnor U551 (N_551,In_1905,In_1480);
nor U552 (N_552,In_451,In_381);
nand U553 (N_553,In_2063,In_1317);
xor U554 (N_554,In_1375,In_2331);
nand U555 (N_555,In_250,In_1729);
or U556 (N_556,In_830,In_483);
nor U557 (N_557,In_2152,In_1247);
nand U558 (N_558,In_1800,In_1241);
xnor U559 (N_559,In_631,In_702);
nor U560 (N_560,In_1430,In_102);
xor U561 (N_561,In_47,In_821);
and U562 (N_562,In_2470,In_153);
nand U563 (N_563,In_137,In_31);
nor U564 (N_564,In_997,In_1132);
nand U565 (N_565,In_673,In_1901);
and U566 (N_566,In_499,In_52);
nand U567 (N_567,In_1470,In_1700);
nor U568 (N_568,In_1557,In_1786);
nand U569 (N_569,In_1886,In_1451);
or U570 (N_570,In_119,In_1384);
or U571 (N_571,In_262,In_2232);
nor U572 (N_572,In_912,In_2254);
nor U573 (N_573,In_315,In_1277);
xor U574 (N_574,In_749,In_1759);
or U575 (N_575,In_638,In_2432);
nand U576 (N_576,In_807,In_452);
xnor U577 (N_577,In_810,In_455);
or U578 (N_578,In_2421,In_260);
xnor U579 (N_579,In_1896,In_694);
or U580 (N_580,In_1462,In_944);
nor U581 (N_581,In_883,In_967);
nand U582 (N_582,In_501,In_952);
or U583 (N_583,In_2326,In_593);
and U584 (N_584,In_1464,In_244);
nand U585 (N_585,In_1807,In_2392);
and U586 (N_586,In_509,In_2246);
xnor U587 (N_587,In_2394,In_170);
or U588 (N_588,In_2248,In_1164);
nand U589 (N_589,In_2307,In_969);
and U590 (N_590,In_222,In_2091);
nand U591 (N_591,In_45,In_1946);
xnor U592 (N_592,In_975,In_777);
nand U593 (N_593,In_1051,In_1513);
or U594 (N_594,In_613,In_1996);
xnor U595 (N_595,In_1439,In_1256);
or U596 (N_596,In_2221,In_901);
nor U597 (N_597,In_1160,In_882);
nor U598 (N_598,In_442,In_356);
and U599 (N_599,In_934,In_124);
or U600 (N_600,In_1709,In_1267);
and U601 (N_601,In_1446,In_281);
nand U602 (N_602,In_820,In_327);
nor U603 (N_603,In_1954,In_261);
xnor U604 (N_604,In_557,In_331);
and U605 (N_605,In_2188,In_446);
nand U606 (N_606,In_677,In_615);
xor U607 (N_607,In_22,In_1216);
nand U608 (N_608,In_441,In_910);
nor U609 (N_609,In_1422,In_1471);
or U610 (N_610,In_1870,In_255);
xnor U611 (N_611,In_2279,In_2101);
or U612 (N_612,In_378,In_2375);
xor U613 (N_613,In_176,In_1526);
or U614 (N_614,In_834,In_2012);
nand U615 (N_615,In_311,In_991);
nand U616 (N_616,In_1825,In_2355);
nand U617 (N_617,In_1865,In_2201);
nor U618 (N_618,In_2405,In_585);
nand U619 (N_619,In_1982,In_848);
and U620 (N_620,In_2190,In_582);
nand U621 (N_621,In_1542,In_687);
nor U622 (N_622,In_782,In_1680);
or U623 (N_623,In_198,In_2014);
and U624 (N_624,In_2265,In_2399);
or U625 (N_625,In_2344,In_1997);
or U626 (N_626,In_83,In_516);
nor U627 (N_627,In_587,In_2444);
nand U628 (N_628,In_2115,In_104);
xor U629 (N_629,In_1427,In_2300);
nand U630 (N_630,In_113,In_1233);
xor U631 (N_631,In_2281,In_646);
or U632 (N_632,In_948,In_1826);
nor U633 (N_633,In_1485,In_1947);
nor U634 (N_634,In_205,In_1024);
xnor U635 (N_635,In_1632,In_574);
xor U636 (N_636,In_652,In_1600);
xor U637 (N_637,In_1137,In_1304);
xnor U638 (N_638,In_2180,In_1313);
or U639 (N_639,In_1698,In_1754);
and U640 (N_640,In_709,In_1691);
nand U641 (N_641,In_1570,In_1991);
and U642 (N_642,In_2485,In_1858);
nand U643 (N_643,In_594,In_99);
and U644 (N_644,In_556,In_28);
and U645 (N_645,In_614,In_447);
or U646 (N_646,In_230,In_1077);
nand U647 (N_647,In_445,In_1207);
nor U648 (N_648,In_1070,In_628);
nor U649 (N_649,In_1020,In_1511);
and U650 (N_650,In_1873,In_2216);
xor U651 (N_651,In_2057,In_228);
nand U652 (N_652,In_1938,In_520);
nand U653 (N_653,In_1046,In_1603);
nor U654 (N_654,In_1953,In_1643);
or U655 (N_655,In_1236,In_845);
and U656 (N_656,In_1431,In_128);
or U657 (N_657,In_2038,In_2162);
xnor U658 (N_658,In_1084,In_2015);
nor U659 (N_659,In_372,In_456);
or U660 (N_660,In_2173,In_303);
and U661 (N_661,In_1966,In_2119);
xor U662 (N_662,In_2385,In_1291);
and U663 (N_663,In_458,In_1637);
nor U664 (N_664,In_181,In_1900);
or U665 (N_665,In_362,In_865);
nor U666 (N_666,In_1162,In_2125);
xor U667 (N_667,In_1200,In_1682);
and U668 (N_668,In_365,In_1503);
xor U669 (N_669,In_1824,In_2319);
xor U670 (N_670,In_2428,In_1355);
xnor U671 (N_671,In_1509,In_2492);
or U672 (N_672,In_1671,In_957);
nor U673 (N_673,In_1611,In_618);
nor U674 (N_674,In_319,In_1549);
nand U675 (N_675,In_502,In_2411);
nand U676 (N_676,In_835,In_132);
xnor U677 (N_677,In_708,In_404);
or U678 (N_678,In_584,In_218);
nor U679 (N_679,In_1348,In_592);
nand U680 (N_680,In_1803,In_1115);
nand U681 (N_681,In_1176,In_1855);
nand U682 (N_682,In_1686,In_248);
xnor U683 (N_683,In_1309,In_825);
nor U684 (N_684,In_305,In_263);
and U685 (N_685,In_1817,In_2058);
xnor U686 (N_686,In_353,In_1787);
xnor U687 (N_687,In_1891,In_2166);
nand U688 (N_688,In_731,In_1955);
and U689 (N_689,In_2261,In_2061);
xor U690 (N_690,In_1918,In_1952);
and U691 (N_691,In_68,In_630);
nor U692 (N_692,In_206,In_129);
and U693 (N_693,In_419,In_1932);
and U694 (N_694,In_1361,In_1778);
or U695 (N_695,In_1350,In_1423);
or U696 (N_696,In_1016,In_359);
nor U697 (N_697,In_1490,In_1925);
nand U698 (N_698,In_2415,In_2343);
nor U699 (N_699,In_838,In_2465);
xnor U700 (N_700,In_1945,In_1323);
xor U701 (N_701,In_78,In_610);
or U702 (N_702,In_568,In_1151);
nor U703 (N_703,In_1742,In_1244);
and U704 (N_704,In_931,In_1880);
nor U705 (N_705,In_223,In_2007);
nor U706 (N_706,In_2362,In_140);
nand U707 (N_707,In_2496,In_436);
xor U708 (N_708,In_2009,In_1333);
or U709 (N_709,In_1481,In_2446);
nand U710 (N_710,In_1735,In_581);
nand U711 (N_711,In_2327,In_2447);
or U712 (N_712,In_1571,In_508);
and U713 (N_713,In_1930,In_2233);
and U714 (N_714,In_1331,In_1547);
nand U715 (N_715,In_605,In_2030);
nor U716 (N_716,In_71,In_1968);
xnor U717 (N_717,In_994,In_1367);
or U718 (N_718,In_1827,In_67);
and U719 (N_719,In_2431,In_1956);
nand U720 (N_720,In_1098,In_586);
or U721 (N_721,In_282,In_462);
or U722 (N_722,In_1245,In_786);
nand U723 (N_723,In_2346,In_894);
or U724 (N_724,In_1660,In_1679);
xor U725 (N_725,In_1944,In_721);
and U726 (N_726,In_1665,In_1282);
or U727 (N_727,In_1368,In_214);
nand U728 (N_728,In_809,In_2365);
nand U729 (N_729,In_1728,In_2123);
nor U730 (N_730,In_1623,In_1662);
and U731 (N_731,In_1382,In_768);
xor U732 (N_732,In_1607,In_1533);
or U733 (N_733,In_1356,In_253);
nor U734 (N_734,In_1141,In_1387);
xnor U735 (N_735,In_671,In_533);
xor U736 (N_736,In_2475,In_1478);
and U737 (N_737,In_486,In_118);
or U738 (N_738,In_1327,In_668);
or U739 (N_739,In_1140,In_1601);
nand U740 (N_740,In_760,In_2053);
nand U741 (N_741,In_495,In_2467);
or U742 (N_742,In_1479,In_1919);
nand U743 (N_743,In_661,In_418);
and U744 (N_744,In_2196,In_1587);
xor U745 (N_745,In_1111,In_29);
nand U746 (N_746,In_863,In_616);
or U747 (N_747,In_1146,In_1567);
nand U748 (N_748,In_1843,In_400);
xnor U749 (N_749,In_1118,In_868);
nor U750 (N_750,In_1487,In_1500);
or U751 (N_751,In_2089,In_494);
nand U752 (N_752,In_2146,In_1189);
or U753 (N_753,In_753,In_210);
or U754 (N_754,In_1454,In_580);
xor U755 (N_755,In_1719,In_929);
nand U756 (N_756,In_1328,In_2272);
or U757 (N_757,In_1058,In_2287);
and U758 (N_758,In_1483,In_1134);
or U759 (N_759,In_313,In_990);
and U760 (N_760,In_1967,In_765);
and U761 (N_761,In_1149,In_1206);
and U762 (N_762,In_2149,In_566);
xor U763 (N_763,In_943,In_1262);
nor U764 (N_764,In_1379,In_958);
xnor U765 (N_765,In_1201,In_1774);
nor U766 (N_766,In_322,In_1596);
nor U767 (N_767,In_1089,In_2211);
xnor U768 (N_768,In_893,In_2083);
or U769 (N_769,In_2303,In_1714);
nand U770 (N_770,In_1959,In_781);
xor U771 (N_771,In_184,In_187);
or U772 (N_772,In_911,In_563);
nor U773 (N_773,In_1783,In_1275);
or U774 (N_774,In_1449,In_1618);
nand U775 (N_775,In_448,In_180);
and U776 (N_776,In_1758,In_2136);
nor U777 (N_777,In_1036,In_514);
and U778 (N_778,In_416,In_395);
and U779 (N_779,In_1578,In_368);
and U780 (N_780,In_2264,In_212);
and U781 (N_781,In_2336,In_101);
xor U782 (N_782,In_1652,In_1699);
and U783 (N_783,In_1534,In_2427);
or U784 (N_784,In_2139,In_725);
and U785 (N_785,In_544,In_1516);
nand U786 (N_786,In_1017,In_554);
nand U787 (N_787,In_36,In_583);
nor U788 (N_788,In_61,In_1086);
nand U789 (N_789,In_27,In_2440);
nor U790 (N_790,In_635,In_1265);
and U791 (N_791,In_1010,In_1453);
or U792 (N_792,In_204,In_1071);
nor U793 (N_793,In_13,In_1929);
nand U794 (N_794,In_1789,In_219);
xnor U795 (N_795,In_89,In_2086);
and U796 (N_796,In_247,In_2131);
and U797 (N_797,In_1514,In_1788);
nand U798 (N_798,In_1026,In_644);
and U799 (N_799,In_472,In_142);
and U800 (N_800,In_822,In_493);
nor U801 (N_801,In_2499,In_1543);
nand U802 (N_802,In_1043,In_1052);
nand U803 (N_803,In_889,In_1364);
and U804 (N_804,In_324,In_344);
nand U805 (N_805,In_808,In_1298);
nor U806 (N_806,In_1011,In_2388);
nor U807 (N_807,In_1703,In_2163);
nor U808 (N_808,In_1280,In_1540);
and U809 (N_809,In_239,In_1532);
nor U810 (N_810,In_515,In_321);
nand U811 (N_811,In_796,In_1751);
nand U812 (N_812,In_691,In_1002);
xnor U813 (N_813,In_642,In_2489);
xor U814 (N_814,In_658,In_2237);
and U815 (N_815,In_1390,In_2354);
xnor U816 (N_816,In_2039,In_785);
xor U817 (N_817,In_1076,In_1167);
xor U818 (N_818,In_973,In_797);
nand U819 (N_819,In_2013,In_208);
nor U820 (N_820,In_1922,In_2478);
nor U821 (N_821,In_273,In_2157);
xor U822 (N_822,In_799,In_976);
and U823 (N_823,In_570,In_1964);
xor U824 (N_824,In_1836,In_340);
xor U825 (N_825,In_1619,In_2226);
or U826 (N_826,In_876,In_1909);
nand U827 (N_827,In_2441,In_2456);
or U828 (N_828,In_607,In_2364);
and U829 (N_829,In_521,In_1467);
xor U830 (N_830,In_1793,In_2498);
nor U831 (N_831,In_895,In_309);
or U832 (N_832,In_793,In_1583);
nand U833 (N_833,In_2145,In_2348);
xor U834 (N_834,In_1061,In_299);
nand U835 (N_835,In_1640,In_858);
nand U836 (N_836,In_2311,In_657);
nand U837 (N_837,In_1109,In_1187);
xor U838 (N_838,In_1844,In_2268);
or U839 (N_839,In_383,In_276);
and U840 (N_840,In_899,In_1000);
or U841 (N_841,In_1477,In_189);
nand U842 (N_842,In_2202,In_2017);
nor U843 (N_843,In_306,In_697);
or U844 (N_844,In_695,In_1576);
nand U845 (N_845,In_1315,In_1562);
nand U846 (N_846,In_1625,In_2294);
nand U847 (N_847,In_636,In_17);
and U848 (N_848,In_2179,In_2410);
xnor U849 (N_849,In_376,In_2138);
or U850 (N_850,In_1580,In_167);
nor U851 (N_851,In_1376,In_1631);
xor U852 (N_852,In_2329,In_2034);
nand U853 (N_853,In_2060,In_862);
xor U854 (N_854,In_1517,In_1135);
nand U855 (N_855,In_2059,In_1399);
nor U856 (N_856,In_1876,In_51);
nand U857 (N_857,In_595,In_1723);
nand U858 (N_858,In_995,In_288);
and U859 (N_859,In_1504,In_681);
nor U860 (N_860,In_249,In_1110);
nor U861 (N_861,In_2296,In_301);
nor U862 (N_862,In_46,In_1025);
nand U863 (N_863,In_1080,In_1776);
xor U864 (N_864,In_2135,In_2448);
nor U865 (N_865,In_539,In_1432);
and U866 (N_866,In_707,In_1117);
nand U867 (N_867,In_1012,In_412);
nor U868 (N_868,In_763,In_188);
nand U869 (N_869,In_2258,In_347);
or U870 (N_870,In_1310,In_878);
xnor U871 (N_871,In_2384,In_1424);
and U872 (N_872,In_1143,In_1524);
and U873 (N_873,In_828,In_891);
xor U874 (N_874,In_527,In_1254);
xnor U875 (N_875,In_437,In_207);
or U876 (N_876,In_879,In_1178);
nor U877 (N_877,In_903,In_2243);
nor U878 (N_878,In_106,In_2400);
xor U879 (N_879,In_819,In_421);
or U880 (N_880,In_1639,In_2228);
xnor U881 (N_881,In_908,In_1496);
xor U882 (N_882,In_1994,In_655);
nor U883 (N_883,In_252,In_382);
or U884 (N_884,In_2452,In_922);
nand U885 (N_885,In_1092,In_278);
xor U886 (N_886,In_1113,In_435);
and U887 (N_887,In_1312,In_1268);
and U888 (N_888,In_1799,In_93);
or U889 (N_889,In_2334,In_2165);
or U890 (N_890,In_1681,In_2438);
or U891 (N_891,In_621,In_1306);
or U892 (N_892,In_602,In_1983);
xnor U893 (N_893,In_662,In_1352);
nand U894 (N_894,In_837,In_1366);
and U895 (N_895,In_880,In_1770);
nand U896 (N_896,In_1209,In_1097);
or U897 (N_897,In_813,In_1617);
and U898 (N_898,In_329,In_1525);
nand U899 (N_899,In_271,In_1704);
nand U900 (N_900,In_2041,In_715);
or U901 (N_901,In_1819,In_2494);
or U902 (N_902,In_930,In_2437);
and U903 (N_903,In_2301,In_2477);
xnor U904 (N_904,In_1561,In_2352);
and U905 (N_905,In_1823,In_1246);
xor U906 (N_906,In_2357,In_688);
nand U907 (N_907,In_1190,In_1779);
nor U908 (N_908,In_2054,In_1810);
and U909 (N_909,In_1255,In_902);
nand U910 (N_910,In_888,In_1031);
nor U911 (N_911,In_1269,In_884);
or U912 (N_912,In_2458,In_2372);
nor U913 (N_913,In_955,In_63);
nand U914 (N_914,In_2214,In_2191);
xor U915 (N_915,In_316,In_696);
nand U916 (N_916,In_1848,In_800);
xnor U917 (N_917,In_1461,In_964);
and U918 (N_918,In_1180,In_2463);
and U919 (N_919,In_850,In_2286);
xnor U920 (N_920,In_1772,In_1184);
nand U921 (N_921,In_1154,In_474);
or U922 (N_922,In_2420,In_1692);
nor U923 (N_923,In_1307,In_597);
and U924 (N_924,In_1271,In_2070);
nand U925 (N_925,In_1170,In_478);
nor U926 (N_926,In_487,In_1047);
xor U927 (N_927,In_2412,In_2103);
and U928 (N_928,In_1195,In_2404);
or U929 (N_929,In_1074,In_2004);
or U930 (N_930,In_2043,In_1837);
nand U931 (N_931,In_2213,In_1739);
or U932 (N_932,In_1738,In_1821);
nand U933 (N_933,In_33,In_2062);
and U934 (N_934,In_1734,In_1707);
nor U935 (N_935,In_1958,In_2142);
nand U936 (N_936,In_23,In_1463);
xnor U937 (N_937,In_2068,In_1122);
or U938 (N_938,In_1941,In_1469);
xnor U939 (N_939,In_280,In_302);
xnor U940 (N_940,In_864,In_1599);
and U941 (N_941,In_233,In_1258);
or U942 (N_942,In_298,In_1105);
nand U943 (N_943,In_100,In_926);
xor U944 (N_944,In_917,In_1566);
and U945 (N_945,In_2128,In_1001);
xnor U946 (N_946,In_1260,In_235);
nand U947 (N_947,In_2209,In_2491);
and U948 (N_948,In_1507,In_1948);
or U949 (N_949,In_2022,In_2460);
xor U950 (N_950,In_1974,In_757);
or U951 (N_951,In_2257,In_2495);
or U952 (N_952,In_2113,In_53);
or U953 (N_953,In_1344,In_1752);
xor U954 (N_954,In_1062,In_547);
and U955 (N_955,In_1708,In_936);
nand U956 (N_956,In_737,In_2003);
or U957 (N_957,In_2020,In_2298);
xor U958 (N_958,In_2215,In_1127);
and U959 (N_959,In_1021,In_1877);
or U960 (N_960,In_387,In_892);
xnor U961 (N_961,In_1475,In_510);
nand U962 (N_962,In_350,In_2379);
or U963 (N_963,In_70,In_82);
xnor U964 (N_964,In_1325,In_611);
xor U965 (N_965,In_466,In_2374);
xnor U966 (N_966,In_827,In_1893);
and U967 (N_967,In_900,In_2430);
nand U968 (N_968,In_916,In_1828);
nand U969 (N_969,In_1169,In_1360);
or U970 (N_970,In_1834,In_748);
and U971 (N_971,In_588,In_334);
xnor U972 (N_972,In_241,In_229);
or U973 (N_973,In_1520,In_2200);
xor U974 (N_974,In_242,In_1546);
nor U975 (N_975,In_1065,In_2029);
xor U976 (N_976,In_469,In_701);
and U977 (N_977,In_1349,In_2453);
nor U978 (N_978,In_779,In_1853);
nor U979 (N_979,In_818,In_116);
and U980 (N_980,In_1761,In_2340);
or U981 (N_981,In_2224,In_824);
nor U982 (N_982,In_567,In_424);
nor U983 (N_983,In_706,In_2241);
nor U984 (N_984,In_1297,In_1425);
or U985 (N_985,In_2389,In_1104);
or U986 (N_986,In_312,In_2006);
or U987 (N_987,In_2027,In_121);
nor U988 (N_988,In_2472,In_1610);
and U989 (N_989,In_471,In_1445);
and U990 (N_990,In_1223,In_1495);
nand U991 (N_991,In_1041,In_2476);
nand U992 (N_992,In_1022,In_1924);
or U993 (N_993,In_2308,In_155);
xor U994 (N_994,In_746,In_665);
nand U995 (N_995,In_1917,In_1292);
and U996 (N_996,In_921,In_1784);
and U997 (N_997,In_2271,In_2403);
and U998 (N_998,In_1380,In_2393);
nor U999 (N_999,In_784,In_974);
nand U1000 (N_1000,In_1096,In_790);
or U1001 (N_1001,In_2483,In_2457);
and U1002 (N_1002,In_2212,In_117);
or U1003 (N_1003,In_1564,In_1391);
nor U1004 (N_1004,In_2042,In_38);
or U1005 (N_1005,In_257,In_2387);
xnor U1006 (N_1006,In_853,In_1408);
nor U1007 (N_1007,In_50,In_1628);
nor U1008 (N_1008,In_1357,In_648);
xnor U1009 (N_1009,In_503,In_1014);
and U1010 (N_1010,In_1078,In_1099);
or U1011 (N_1011,In_2218,In_1155);
nand U1012 (N_1012,In_1007,In_1332);
and U1013 (N_1013,In_2230,In_162);
nand U1014 (N_1014,In_1693,In_2075);
and U1015 (N_1015,In_2225,In_1359);
and U1016 (N_1016,In_1556,In_360);
xor U1017 (N_1017,In_1838,In_1961);
and U1018 (N_1018,In_959,In_932);
nor U1019 (N_1019,In_2373,In_139);
xnor U1020 (N_1020,In_251,In_1553);
and U1021 (N_1021,In_403,In_41);
and U1022 (N_1022,In_396,In_1401);
nand U1023 (N_1023,In_2186,In_2048);
nor U1024 (N_1024,In_2455,In_26);
nor U1025 (N_1025,In_1085,In_589);
nor U1026 (N_1026,In_1830,In_1913);
or U1027 (N_1027,In_1027,In_2240);
xnor U1028 (N_1028,In_1744,In_431);
and U1029 (N_1029,In_341,In_1702);
or U1030 (N_1030,In_1320,In_2001);
xor U1031 (N_1031,In_519,In_2244);
and U1032 (N_1032,In_1518,In_1175);
xnor U1033 (N_1033,In_1133,In_815);
and U1034 (N_1034,In_1493,In_54);
nor U1035 (N_1035,In_1745,In_1501);
or U1036 (N_1036,In_2482,In_1287);
or U1037 (N_1037,In_2023,In_2247);
or U1038 (N_1038,In_1973,In_1541);
xnor U1039 (N_1039,In_2306,In_619);
xnor U1040 (N_1040,In_1370,In_2314);
or U1041 (N_1041,In_1711,In_1894);
and U1042 (N_1042,In_2285,In_724);
nand U1043 (N_1043,In_481,In_2051);
and U1044 (N_1044,In_2189,In_1590);
or U1045 (N_1045,In_1839,In_1191);
xnor U1046 (N_1046,In_1468,In_953);
or U1047 (N_1047,In_905,In_1395);
and U1048 (N_1048,In_6,In_174);
xor U1049 (N_1049,In_1341,In_1747);
nor U1050 (N_1050,In_2378,In_734);
nor U1051 (N_1051,In_111,In_385);
nor U1052 (N_1052,In_1393,In_2199);
or U1053 (N_1053,In_1008,In_1416);
and U1054 (N_1054,In_2367,In_290);
nand U1055 (N_1055,In_713,In_2064);
xnor U1056 (N_1056,In_1050,In_1365);
and U1057 (N_1057,In_60,In_1505);
and U1058 (N_1058,In_1029,In_1969);
xnor U1059 (N_1059,In_393,In_182);
nand U1060 (N_1060,In_335,In_84);
nor U1061 (N_1061,In_1138,In_443);
nor U1062 (N_1062,In_1229,In_2256);
xnor U1063 (N_1063,In_1963,In_2433);
nand U1064 (N_1064,In_498,In_1841);
xor U1065 (N_1065,In_2069,In_851);
and U1066 (N_1066,In_191,In_914);
nand U1067 (N_1067,In_1879,In_2416);
or U1068 (N_1068,In_1283,In_535);
nand U1069 (N_1069,In_1343,In_1805);
and U1070 (N_1070,In_2227,In_1753);
or U1071 (N_1071,In_1193,In_643);
and U1072 (N_1072,In_1347,In_2332);
nor U1073 (N_1073,In_829,In_641);
nand U1074 (N_1074,In_904,In_1502);
xnor U1075 (N_1075,In_2312,In_1286);
nor U1076 (N_1076,In_1548,In_550);
nor U1077 (N_1077,In_1383,In_1721);
and U1078 (N_1078,In_2148,In_1166);
or U1079 (N_1079,In_505,In_1165);
nor U1080 (N_1080,In_1433,In_2098);
and U1081 (N_1081,In_1970,In_2035);
xor U1082 (N_1082,In_823,In_1440);
or U1083 (N_1083,In_2079,In_1053);
nand U1084 (N_1084,In_740,In_1730);
nor U1085 (N_1085,In_842,In_1329);
or U1086 (N_1086,In_2337,In_56);
nor U1087 (N_1087,In_843,In_1426);
nand U1088 (N_1088,In_2316,In_1815);
and U1089 (N_1089,In_2167,In_1081);
xor U1090 (N_1090,In_886,In_1413);
nor U1091 (N_1091,In_87,In_599);
and U1092 (N_1092,In_1852,In_166);
nand U1093 (N_1093,In_788,In_766);
nor U1094 (N_1094,In_711,In_984);
nor U1095 (N_1095,In_131,In_270);
nor U1096 (N_1096,In_390,In_710);
xnor U1097 (N_1097,In_634,In_1259);
nand U1098 (N_1098,In_266,In_2313);
xnor U1099 (N_1099,In_1575,In_199);
nand U1100 (N_1100,In_1196,In_1388);
xnor U1101 (N_1101,In_1608,In_66);
nor U1102 (N_1102,In_477,In_804);
and U1103 (N_1103,In_1895,In_2177);
and U1104 (N_1104,In_2242,In_1889);
xnor U1105 (N_1105,In_2170,In_2082);
nor U1106 (N_1106,In_992,In_773);
xor U1107 (N_1107,In_2238,In_232);
or U1108 (N_1108,In_2100,In_647);
or U1109 (N_1109,In_792,In_2407);
and U1110 (N_1110,In_633,In_675);
or U1111 (N_1111,In_1412,In_265);
nand U1112 (N_1112,In_1687,In_540);
nand U1113 (N_1113,In_1473,In_1856);
nand U1114 (N_1114,In_2402,In_108);
nand U1115 (N_1115,In_1281,In_2067);
or U1116 (N_1116,In_1820,In_144);
or U1117 (N_1117,In_2121,In_292);
or U1118 (N_1118,In_1342,In_625);
or U1119 (N_1119,In_576,In_2429);
xnor U1120 (N_1120,In_343,In_989);
or U1121 (N_1121,In_522,In_2178);
and U1122 (N_1122,In_428,In_330);
nor U1123 (N_1123,In_2184,In_1015);
nand U1124 (N_1124,In_1581,In_217);
nand U1125 (N_1125,In_2090,In_787);
or U1126 (N_1126,In_2106,In_231);
xnor U1127 (N_1127,In_670,In_1545);
xnor U1128 (N_1128,In_1238,In_529);
nand U1129 (N_1129,In_1551,In_2464);
and U1130 (N_1130,In_1690,In_1211);
or U1131 (N_1131,In_1374,In_2159);
and U1132 (N_1132,In_506,In_81);
nor U1133 (N_1133,In_141,In_1650);
and U1134 (N_1134,In_1494,In_1999);
nor U1135 (N_1135,In_1442,In_1159);
xor U1136 (N_1136,In_578,In_640);
and U1137 (N_1137,In_679,In_1554);
xnor U1138 (N_1138,In_717,In_2234);
or U1139 (N_1139,In_1937,In_8);
xnor U1140 (N_1140,In_920,In_177);
or U1141 (N_1141,In_2078,In_1414);
and U1142 (N_1142,In_866,In_764);
xnor U1143 (N_1143,In_770,In_653);
or U1144 (N_1144,In_1989,In_1811);
nand U1145 (N_1145,In_2185,In_552);
nand U1146 (N_1146,In_2462,In_2295);
nor U1147 (N_1147,In_1669,In_279);
xor U1148 (N_1148,In_751,In_881);
xnor U1149 (N_1149,In_1474,In_596);
nor U1150 (N_1150,In_1902,In_2323);
nor U1151 (N_1151,In_542,In_1866);
or U1152 (N_1152,In_1276,In_2236);
and U1153 (N_1153,In_1644,In_1840);
and U1154 (N_1154,In_1658,In_1743);
nor U1155 (N_1155,In_1849,In_1407);
nand U1156 (N_1156,In_2361,In_1157);
nand U1157 (N_1157,In_1091,In_1915);
or U1158 (N_1158,In_1182,In_1874);
or U1159 (N_1159,In_1741,In_432);
nor U1160 (N_1160,In_831,In_1694);
nand U1161 (N_1161,In_1656,In_1285);
or U1162 (N_1162,In_549,In_1976);
nor U1163 (N_1163,In_467,In_2120);
nor U1164 (N_1164,In_2318,In_513);
and U1165 (N_1165,In_965,In_847);
nor U1166 (N_1166,In_1249,In_925);
nor U1167 (N_1167,In_2088,In_1301);
and U1168 (N_1168,In_1987,In_406);
nand U1169 (N_1169,In_2353,In_339);
nand U1170 (N_1170,In_536,In_417);
and U1171 (N_1171,In_2417,In_2395);
or U1172 (N_1172,In_849,In_2176);
or U1173 (N_1173,In_2356,In_1326);
nor U1174 (N_1174,In_2282,In_399);
or U1175 (N_1175,In_364,In_2223);
nand U1176 (N_1176,In_2339,In_2095);
nand U1177 (N_1177,In_1289,In_1995);
nor U1178 (N_1178,In_1962,In_1726);
xor U1179 (N_1179,In_43,In_398);
xnor U1180 (N_1180,In_1218,In_40);
and U1181 (N_1181,In_1689,In_154);
or U1182 (N_1182,In_877,In_2451);
nand U1183 (N_1183,In_130,In_1736);
nand U1184 (N_1184,In_1688,In_1636);
nand U1185 (N_1185,In_771,In_363);
and U1186 (N_1186,In_2324,In_1101);
nor U1187 (N_1187,In_2000,In_789);
and U1188 (N_1188,In_1121,In_1396);
nand U1189 (N_1189,In_73,In_1512);
xor U1190 (N_1190,In_1150,In_1261);
nor U1191 (N_1191,In_179,In_2151);
nand U1192 (N_1192,In_1762,In_2304);
or U1193 (N_1193,In_1673,In_295);
nor U1194 (N_1194,In_714,In_72);
nand U1195 (N_1195,In_918,In_1263);
or U1196 (N_1196,In_236,In_2305);
nor U1197 (N_1197,In_1882,In_16);
xor U1198 (N_1198,In_1684,In_999);
and U1199 (N_1199,In_561,In_2320);
or U1200 (N_1200,In_1173,In_537);
nor U1201 (N_1201,In_645,In_2450);
nand U1202 (N_1202,In_947,In_2108);
and U1203 (N_1203,In_2094,In_1048);
and U1204 (N_1204,In_801,In_1338);
xor U1205 (N_1205,In_1156,In_1232);
nand U1206 (N_1206,In_380,In_612);
nand U1207 (N_1207,In_5,In_2132);
xnor U1208 (N_1208,In_1712,In_2376);
xor U1209 (N_1209,In_287,In_759);
or U1210 (N_1210,In_2422,In_1212);
nand U1211 (N_1211,In_2461,In_978);
or U1212 (N_1212,In_109,In_511);
xor U1213 (N_1213,In_966,In_1185);
and U1214 (N_1214,In_227,In_1847);
nor U1215 (N_1215,In_718,In_1429);
nor U1216 (N_1216,In_2045,In_221);
and U1217 (N_1217,In_1814,In_1019);
and U1218 (N_1218,In_1460,In_192);
nor U1219 (N_1219,In_2140,In_1988);
nor U1220 (N_1220,In_1908,In_2425);
nand U1221 (N_1221,In_2262,In_1340);
xnor U1222 (N_1222,In_1183,In_146);
nand U1223 (N_1223,In_1168,In_950);
nand U1224 (N_1224,In_2171,In_1230);
xor U1225 (N_1225,In_1934,In_2351);
nor U1226 (N_1226,In_1609,In_293);
xnor U1227 (N_1227,In_1082,In_122);
nand U1228 (N_1228,In_798,In_1371);
or U1229 (N_1229,In_127,In_9);
nand U1230 (N_1230,In_727,In_1106);
or U1231 (N_1231,In_2406,In_871);
xor U1232 (N_1232,In_738,In_546);
xnor U1233 (N_1233,In_2487,In_1531);
and U1234 (N_1234,In_58,In_998);
nor U1235 (N_1235,In_2019,In_559);
nand U1236 (N_1236,In_75,In_2239);
nor U1237 (N_1237,In_159,In_1194);
or U1238 (N_1238,In_2126,In_1322);
xor U1239 (N_1239,In_1705,In_1675);
and U1240 (N_1240,In_391,In_1023);
or U1241 (N_1241,In_2284,In_358);
xor U1242 (N_1242,In_924,In_2358);
nand U1243 (N_1243,In_1476,In_1861);
xnor U1244 (N_1244,In_1801,In_1916);
nand U1245 (N_1245,In_1718,In_617);
xor U1246 (N_1246,In_2080,In_1057);
xnor U1247 (N_1247,In_1780,In_1003);
nor U1248 (N_1248,In_2255,In_1188);
and U1249 (N_1249,In_1299,In_183);
nor U1250 (N_1250,In_349,In_1130);
nand U1251 (N_1251,In_644,In_805);
xnor U1252 (N_1252,In_1895,In_1119);
nor U1253 (N_1253,In_1165,In_1964);
nor U1254 (N_1254,In_1649,In_66);
nor U1255 (N_1255,In_515,In_1104);
or U1256 (N_1256,In_1848,In_114);
xor U1257 (N_1257,In_1217,In_309);
nand U1258 (N_1258,In_2089,In_1241);
xnor U1259 (N_1259,In_681,In_379);
or U1260 (N_1260,In_1043,In_233);
nand U1261 (N_1261,In_2212,In_2403);
nand U1262 (N_1262,In_2047,In_1933);
nor U1263 (N_1263,In_1709,In_1376);
nor U1264 (N_1264,In_595,In_2418);
nor U1265 (N_1265,In_2476,In_589);
or U1266 (N_1266,In_1098,In_123);
nor U1267 (N_1267,In_587,In_1835);
xnor U1268 (N_1268,In_1063,In_1751);
nor U1269 (N_1269,In_185,In_1654);
nand U1270 (N_1270,In_1961,In_2392);
nor U1271 (N_1271,In_2310,In_164);
xnor U1272 (N_1272,In_637,In_1440);
nor U1273 (N_1273,In_1190,In_380);
xor U1274 (N_1274,In_32,In_1609);
nor U1275 (N_1275,In_1571,In_1130);
or U1276 (N_1276,In_1272,In_2351);
xor U1277 (N_1277,In_1546,In_2358);
nand U1278 (N_1278,In_2494,In_2063);
xnor U1279 (N_1279,In_1613,In_518);
nor U1280 (N_1280,In_2179,In_110);
nor U1281 (N_1281,In_473,In_630);
or U1282 (N_1282,In_862,In_747);
nor U1283 (N_1283,In_887,In_241);
nor U1284 (N_1284,In_1025,In_486);
nor U1285 (N_1285,In_2418,In_899);
and U1286 (N_1286,In_791,In_1040);
nor U1287 (N_1287,In_1636,In_1917);
nand U1288 (N_1288,In_1037,In_164);
nor U1289 (N_1289,In_537,In_2388);
or U1290 (N_1290,In_2015,In_96);
nand U1291 (N_1291,In_36,In_1500);
nor U1292 (N_1292,In_1780,In_1509);
nor U1293 (N_1293,In_1396,In_113);
and U1294 (N_1294,In_1288,In_1578);
nand U1295 (N_1295,In_1619,In_1785);
and U1296 (N_1296,In_1483,In_2494);
and U1297 (N_1297,In_1103,In_207);
nand U1298 (N_1298,In_133,In_1452);
and U1299 (N_1299,In_1300,In_1026);
nand U1300 (N_1300,In_354,In_1853);
and U1301 (N_1301,In_1541,In_8);
xnor U1302 (N_1302,In_2111,In_1608);
nand U1303 (N_1303,In_1500,In_1916);
nand U1304 (N_1304,In_1116,In_2497);
nand U1305 (N_1305,In_781,In_420);
xor U1306 (N_1306,In_620,In_1113);
xor U1307 (N_1307,In_767,In_675);
or U1308 (N_1308,In_944,In_595);
xnor U1309 (N_1309,In_1117,In_867);
xnor U1310 (N_1310,In_1012,In_1299);
nand U1311 (N_1311,In_1335,In_88);
and U1312 (N_1312,In_253,In_1006);
xor U1313 (N_1313,In_247,In_1105);
xor U1314 (N_1314,In_1144,In_836);
xnor U1315 (N_1315,In_964,In_337);
or U1316 (N_1316,In_100,In_2399);
nand U1317 (N_1317,In_786,In_523);
nor U1318 (N_1318,In_289,In_1484);
nand U1319 (N_1319,In_1463,In_2085);
nand U1320 (N_1320,In_2147,In_1460);
nor U1321 (N_1321,In_1149,In_1154);
and U1322 (N_1322,In_1657,In_1920);
nand U1323 (N_1323,In_1772,In_2377);
nand U1324 (N_1324,In_790,In_810);
or U1325 (N_1325,In_965,In_1771);
or U1326 (N_1326,In_2128,In_2146);
and U1327 (N_1327,In_332,In_1060);
or U1328 (N_1328,In_16,In_1668);
xor U1329 (N_1329,In_252,In_1292);
nand U1330 (N_1330,In_2497,In_1575);
nand U1331 (N_1331,In_2057,In_267);
xor U1332 (N_1332,In_2159,In_1205);
or U1333 (N_1333,In_1865,In_739);
nand U1334 (N_1334,In_465,In_975);
and U1335 (N_1335,In_1471,In_1358);
nand U1336 (N_1336,In_689,In_725);
nor U1337 (N_1337,In_1791,In_242);
nor U1338 (N_1338,In_1676,In_1830);
and U1339 (N_1339,In_492,In_1361);
nand U1340 (N_1340,In_2122,In_1385);
or U1341 (N_1341,In_888,In_1104);
xor U1342 (N_1342,In_700,In_933);
nand U1343 (N_1343,In_2459,In_1830);
and U1344 (N_1344,In_15,In_2138);
and U1345 (N_1345,In_2254,In_888);
or U1346 (N_1346,In_1920,In_2298);
nand U1347 (N_1347,In_1861,In_2419);
nor U1348 (N_1348,In_1725,In_189);
nor U1349 (N_1349,In_548,In_1372);
xnor U1350 (N_1350,In_1923,In_872);
and U1351 (N_1351,In_440,In_345);
xor U1352 (N_1352,In_1596,In_607);
or U1353 (N_1353,In_1314,In_1082);
and U1354 (N_1354,In_1889,In_1909);
nand U1355 (N_1355,In_1578,In_1446);
xnor U1356 (N_1356,In_906,In_526);
xnor U1357 (N_1357,In_2357,In_2301);
and U1358 (N_1358,In_173,In_1173);
nor U1359 (N_1359,In_536,In_2302);
and U1360 (N_1360,In_1,In_991);
xnor U1361 (N_1361,In_1939,In_1716);
or U1362 (N_1362,In_2491,In_1180);
nand U1363 (N_1363,In_220,In_1679);
nand U1364 (N_1364,In_2299,In_516);
and U1365 (N_1365,In_247,In_717);
nand U1366 (N_1366,In_1130,In_1517);
and U1367 (N_1367,In_1759,In_1334);
nand U1368 (N_1368,In_1351,In_660);
and U1369 (N_1369,In_784,In_962);
nor U1370 (N_1370,In_766,In_1386);
nor U1371 (N_1371,In_2209,In_373);
nand U1372 (N_1372,In_1086,In_150);
nand U1373 (N_1373,In_567,In_1545);
and U1374 (N_1374,In_1401,In_2062);
and U1375 (N_1375,In_882,In_359);
nor U1376 (N_1376,In_1,In_311);
and U1377 (N_1377,In_713,In_164);
or U1378 (N_1378,In_1102,In_1516);
xnor U1379 (N_1379,In_779,In_760);
or U1380 (N_1380,In_1268,In_882);
nor U1381 (N_1381,In_432,In_873);
nand U1382 (N_1382,In_2121,In_365);
nand U1383 (N_1383,In_1886,In_260);
and U1384 (N_1384,In_2399,In_388);
nand U1385 (N_1385,In_843,In_389);
or U1386 (N_1386,In_550,In_1167);
xor U1387 (N_1387,In_2277,In_1224);
or U1388 (N_1388,In_28,In_1485);
nand U1389 (N_1389,In_2339,In_2220);
xor U1390 (N_1390,In_109,In_1014);
nand U1391 (N_1391,In_2047,In_945);
and U1392 (N_1392,In_703,In_1135);
xnor U1393 (N_1393,In_2489,In_1284);
xor U1394 (N_1394,In_1976,In_1220);
and U1395 (N_1395,In_2337,In_1625);
nand U1396 (N_1396,In_2084,In_1181);
nand U1397 (N_1397,In_1531,In_1296);
and U1398 (N_1398,In_2045,In_2002);
nand U1399 (N_1399,In_494,In_2456);
nand U1400 (N_1400,In_1252,In_613);
nand U1401 (N_1401,In_1961,In_227);
nand U1402 (N_1402,In_2421,In_962);
nand U1403 (N_1403,In_823,In_1937);
and U1404 (N_1404,In_582,In_257);
and U1405 (N_1405,In_908,In_921);
nor U1406 (N_1406,In_1667,In_1349);
xor U1407 (N_1407,In_2493,In_391);
xnor U1408 (N_1408,In_1343,In_1671);
nand U1409 (N_1409,In_1679,In_2224);
xor U1410 (N_1410,In_1976,In_1572);
nand U1411 (N_1411,In_2201,In_668);
and U1412 (N_1412,In_2319,In_818);
xor U1413 (N_1413,In_1355,In_1450);
nand U1414 (N_1414,In_505,In_2160);
nand U1415 (N_1415,In_1231,In_1585);
or U1416 (N_1416,In_1887,In_630);
and U1417 (N_1417,In_549,In_1498);
xor U1418 (N_1418,In_1082,In_2044);
nor U1419 (N_1419,In_1806,In_690);
and U1420 (N_1420,In_1575,In_683);
nor U1421 (N_1421,In_339,In_97);
or U1422 (N_1422,In_1183,In_809);
xnor U1423 (N_1423,In_340,In_1226);
nor U1424 (N_1424,In_2244,In_1010);
xor U1425 (N_1425,In_1797,In_397);
and U1426 (N_1426,In_98,In_223);
nor U1427 (N_1427,In_1903,In_741);
xor U1428 (N_1428,In_510,In_27);
nand U1429 (N_1429,In_1271,In_1922);
or U1430 (N_1430,In_1874,In_1431);
or U1431 (N_1431,In_2198,In_2156);
nor U1432 (N_1432,In_2295,In_333);
or U1433 (N_1433,In_1404,In_1728);
or U1434 (N_1434,In_93,In_2485);
nor U1435 (N_1435,In_2394,In_1894);
and U1436 (N_1436,In_1631,In_2465);
xnor U1437 (N_1437,In_1905,In_1257);
nor U1438 (N_1438,In_2114,In_127);
and U1439 (N_1439,In_2282,In_1964);
xnor U1440 (N_1440,In_54,In_1461);
nand U1441 (N_1441,In_2459,In_794);
nor U1442 (N_1442,In_1335,In_957);
xnor U1443 (N_1443,In_2266,In_2376);
nor U1444 (N_1444,In_893,In_2441);
or U1445 (N_1445,In_5,In_2135);
and U1446 (N_1446,In_327,In_938);
nand U1447 (N_1447,In_1103,In_1713);
xor U1448 (N_1448,In_2463,In_27);
nand U1449 (N_1449,In_1246,In_1325);
and U1450 (N_1450,In_1643,In_1842);
nand U1451 (N_1451,In_921,In_1308);
or U1452 (N_1452,In_2208,In_255);
or U1453 (N_1453,In_2302,In_598);
nand U1454 (N_1454,In_2490,In_1828);
nor U1455 (N_1455,In_159,In_1524);
or U1456 (N_1456,In_1411,In_1244);
nor U1457 (N_1457,In_850,In_1452);
and U1458 (N_1458,In_2247,In_915);
xnor U1459 (N_1459,In_1804,In_0);
nand U1460 (N_1460,In_95,In_2416);
or U1461 (N_1461,In_1635,In_1573);
or U1462 (N_1462,In_1568,In_168);
nand U1463 (N_1463,In_929,In_1981);
nor U1464 (N_1464,In_190,In_906);
nor U1465 (N_1465,In_1720,In_1250);
or U1466 (N_1466,In_890,In_1951);
nor U1467 (N_1467,In_2016,In_775);
nor U1468 (N_1468,In_1292,In_507);
or U1469 (N_1469,In_1729,In_2443);
nor U1470 (N_1470,In_2163,In_1179);
xor U1471 (N_1471,In_1795,In_2411);
nand U1472 (N_1472,In_2211,In_431);
nand U1473 (N_1473,In_916,In_1551);
and U1474 (N_1474,In_63,In_1424);
or U1475 (N_1475,In_2258,In_1763);
xnor U1476 (N_1476,In_682,In_530);
or U1477 (N_1477,In_1654,In_1856);
or U1478 (N_1478,In_2456,In_2219);
nor U1479 (N_1479,In_67,In_1276);
and U1480 (N_1480,In_496,In_1971);
nand U1481 (N_1481,In_2156,In_2440);
xnor U1482 (N_1482,In_660,In_1033);
or U1483 (N_1483,In_1182,In_700);
nand U1484 (N_1484,In_858,In_1711);
or U1485 (N_1485,In_1652,In_364);
nand U1486 (N_1486,In_715,In_371);
or U1487 (N_1487,In_1744,In_2080);
or U1488 (N_1488,In_1536,In_1492);
nand U1489 (N_1489,In_1346,In_2211);
nor U1490 (N_1490,In_1821,In_1207);
or U1491 (N_1491,In_673,In_1814);
nand U1492 (N_1492,In_2105,In_1288);
and U1493 (N_1493,In_1580,In_1705);
or U1494 (N_1494,In_2326,In_937);
nor U1495 (N_1495,In_466,In_176);
xor U1496 (N_1496,In_1682,In_2117);
and U1497 (N_1497,In_187,In_1820);
and U1498 (N_1498,In_2084,In_1767);
and U1499 (N_1499,In_1896,In_2398);
xor U1500 (N_1500,In_1648,In_1963);
and U1501 (N_1501,In_562,In_2468);
nand U1502 (N_1502,In_1266,In_1332);
nand U1503 (N_1503,In_2435,In_886);
and U1504 (N_1504,In_1409,In_1149);
nand U1505 (N_1505,In_57,In_1628);
or U1506 (N_1506,In_705,In_960);
nor U1507 (N_1507,In_785,In_2123);
nor U1508 (N_1508,In_2332,In_2084);
or U1509 (N_1509,In_2220,In_2068);
nand U1510 (N_1510,In_286,In_2191);
or U1511 (N_1511,In_2233,In_1261);
xor U1512 (N_1512,In_774,In_410);
nand U1513 (N_1513,In_1481,In_1910);
nor U1514 (N_1514,In_1802,In_21);
nor U1515 (N_1515,In_123,In_1781);
xor U1516 (N_1516,In_1031,In_1927);
nor U1517 (N_1517,In_2434,In_213);
nor U1518 (N_1518,In_1123,In_78);
xnor U1519 (N_1519,In_1051,In_2487);
or U1520 (N_1520,In_243,In_1969);
nand U1521 (N_1521,In_401,In_869);
and U1522 (N_1522,In_905,In_2412);
xnor U1523 (N_1523,In_1866,In_550);
xor U1524 (N_1524,In_1748,In_1507);
nand U1525 (N_1525,In_528,In_2041);
and U1526 (N_1526,In_2094,In_572);
and U1527 (N_1527,In_1017,In_1577);
nand U1528 (N_1528,In_1949,In_2195);
or U1529 (N_1529,In_1765,In_45);
xor U1530 (N_1530,In_820,In_81);
or U1531 (N_1531,In_319,In_1314);
and U1532 (N_1532,In_270,In_1694);
nand U1533 (N_1533,In_2361,In_2277);
nor U1534 (N_1534,In_719,In_1789);
and U1535 (N_1535,In_965,In_1221);
nand U1536 (N_1536,In_770,In_513);
xnor U1537 (N_1537,In_589,In_1315);
or U1538 (N_1538,In_1777,In_215);
nand U1539 (N_1539,In_2010,In_738);
nand U1540 (N_1540,In_2194,In_1859);
nor U1541 (N_1541,In_2027,In_1894);
xnor U1542 (N_1542,In_1343,In_1595);
and U1543 (N_1543,In_424,In_2113);
and U1544 (N_1544,In_1770,In_253);
nand U1545 (N_1545,In_1551,In_2202);
xor U1546 (N_1546,In_565,In_889);
nand U1547 (N_1547,In_1857,In_1262);
nand U1548 (N_1548,In_774,In_209);
nand U1549 (N_1549,In_2227,In_1061);
nor U1550 (N_1550,In_1663,In_1079);
or U1551 (N_1551,In_642,In_1295);
and U1552 (N_1552,In_2487,In_462);
nand U1553 (N_1553,In_994,In_1837);
or U1554 (N_1554,In_1674,In_160);
or U1555 (N_1555,In_1567,In_1516);
and U1556 (N_1556,In_2392,In_2081);
xor U1557 (N_1557,In_1142,In_1522);
or U1558 (N_1558,In_1691,In_1260);
xor U1559 (N_1559,In_2288,In_1862);
nor U1560 (N_1560,In_481,In_482);
nor U1561 (N_1561,In_1251,In_2036);
nor U1562 (N_1562,In_2272,In_726);
xor U1563 (N_1563,In_1545,In_347);
nor U1564 (N_1564,In_1186,In_1387);
xnor U1565 (N_1565,In_1772,In_1247);
or U1566 (N_1566,In_695,In_1055);
nor U1567 (N_1567,In_2221,In_1841);
nor U1568 (N_1568,In_1853,In_1352);
nand U1569 (N_1569,In_1216,In_1391);
nor U1570 (N_1570,In_2140,In_2047);
or U1571 (N_1571,In_438,In_2429);
xor U1572 (N_1572,In_1355,In_525);
nor U1573 (N_1573,In_1125,In_318);
nor U1574 (N_1574,In_770,In_72);
and U1575 (N_1575,In_2132,In_790);
xnor U1576 (N_1576,In_1755,In_1854);
and U1577 (N_1577,In_1872,In_1983);
nand U1578 (N_1578,In_2469,In_1816);
nor U1579 (N_1579,In_1195,In_1313);
xnor U1580 (N_1580,In_1030,In_581);
nor U1581 (N_1581,In_1447,In_1412);
nand U1582 (N_1582,In_1077,In_1581);
or U1583 (N_1583,In_2060,In_1106);
nor U1584 (N_1584,In_478,In_1504);
nand U1585 (N_1585,In_332,In_459);
nand U1586 (N_1586,In_615,In_699);
and U1587 (N_1587,In_1379,In_1463);
and U1588 (N_1588,In_347,In_1128);
nor U1589 (N_1589,In_1506,In_1992);
or U1590 (N_1590,In_707,In_698);
nand U1591 (N_1591,In_108,In_16);
and U1592 (N_1592,In_2157,In_383);
and U1593 (N_1593,In_1437,In_947);
nand U1594 (N_1594,In_2384,In_2368);
and U1595 (N_1595,In_1105,In_1209);
nor U1596 (N_1596,In_1774,In_2252);
nor U1597 (N_1597,In_571,In_2102);
and U1598 (N_1598,In_1145,In_1994);
and U1599 (N_1599,In_1825,In_2347);
xnor U1600 (N_1600,In_49,In_108);
nand U1601 (N_1601,In_1142,In_2282);
nand U1602 (N_1602,In_198,In_1047);
xor U1603 (N_1603,In_1052,In_391);
and U1604 (N_1604,In_309,In_1509);
and U1605 (N_1605,In_1222,In_2280);
xor U1606 (N_1606,In_1353,In_2293);
and U1607 (N_1607,In_235,In_2405);
xor U1608 (N_1608,In_1420,In_1576);
and U1609 (N_1609,In_905,In_950);
and U1610 (N_1610,In_2349,In_641);
and U1611 (N_1611,In_1771,In_477);
nand U1612 (N_1612,In_1068,In_1981);
xor U1613 (N_1613,In_1749,In_1148);
nor U1614 (N_1614,In_648,In_254);
nand U1615 (N_1615,In_835,In_1675);
xor U1616 (N_1616,In_2360,In_2140);
or U1617 (N_1617,In_1743,In_2238);
nand U1618 (N_1618,In_1516,In_208);
or U1619 (N_1619,In_524,In_2449);
nor U1620 (N_1620,In_1540,In_585);
and U1621 (N_1621,In_774,In_2378);
nand U1622 (N_1622,In_1709,In_1518);
or U1623 (N_1623,In_2340,In_849);
or U1624 (N_1624,In_1150,In_492);
nor U1625 (N_1625,In_1419,In_1809);
nand U1626 (N_1626,In_1292,In_2065);
nor U1627 (N_1627,In_626,In_708);
nor U1628 (N_1628,In_2378,In_1551);
and U1629 (N_1629,In_431,In_1343);
xor U1630 (N_1630,In_771,In_1050);
or U1631 (N_1631,In_2100,In_2398);
nand U1632 (N_1632,In_374,In_2226);
and U1633 (N_1633,In_240,In_965);
nor U1634 (N_1634,In_508,In_250);
nor U1635 (N_1635,In_1955,In_822);
nand U1636 (N_1636,In_1566,In_937);
xor U1637 (N_1637,In_57,In_1504);
and U1638 (N_1638,In_105,In_2151);
nor U1639 (N_1639,In_657,In_2171);
and U1640 (N_1640,In_2366,In_2447);
nor U1641 (N_1641,In_707,In_12);
nand U1642 (N_1642,In_1538,In_2201);
and U1643 (N_1643,In_2474,In_2366);
or U1644 (N_1644,In_1228,In_2381);
xnor U1645 (N_1645,In_496,In_1321);
and U1646 (N_1646,In_1593,In_1138);
and U1647 (N_1647,In_244,In_1825);
or U1648 (N_1648,In_2452,In_1560);
and U1649 (N_1649,In_102,In_1036);
and U1650 (N_1650,In_2210,In_676);
or U1651 (N_1651,In_365,In_1577);
xor U1652 (N_1652,In_222,In_1751);
and U1653 (N_1653,In_1922,In_667);
nand U1654 (N_1654,In_1796,In_182);
nor U1655 (N_1655,In_1135,In_2031);
nand U1656 (N_1656,In_802,In_1871);
nand U1657 (N_1657,In_712,In_1092);
xor U1658 (N_1658,In_1021,In_1529);
and U1659 (N_1659,In_1793,In_1926);
nand U1660 (N_1660,In_1088,In_2467);
nand U1661 (N_1661,In_1187,In_1526);
nor U1662 (N_1662,In_2198,In_1445);
nand U1663 (N_1663,In_155,In_1867);
nand U1664 (N_1664,In_1071,In_511);
nor U1665 (N_1665,In_837,In_729);
and U1666 (N_1666,In_30,In_1533);
and U1667 (N_1667,In_1024,In_1468);
nor U1668 (N_1668,In_1427,In_1714);
xor U1669 (N_1669,In_406,In_722);
nand U1670 (N_1670,In_1461,In_1191);
nor U1671 (N_1671,In_171,In_48);
nand U1672 (N_1672,In_1273,In_1272);
xor U1673 (N_1673,In_125,In_1215);
and U1674 (N_1674,In_1603,In_168);
or U1675 (N_1675,In_843,In_937);
xnor U1676 (N_1676,In_1431,In_2254);
nand U1677 (N_1677,In_1214,In_199);
or U1678 (N_1678,In_546,In_1728);
or U1679 (N_1679,In_1654,In_2000);
or U1680 (N_1680,In_2265,In_62);
or U1681 (N_1681,In_1050,In_41);
and U1682 (N_1682,In_1231,In_1004);
or U1683 (N_1683,In_819,In_766);
or U1684 (N_1684,In_397,In_1259);
xnor U1685 (N_1685,In_2358,In_240);
xor U1686 (N_1686,In_941,In_1155);
nand U1687 (N_1687,In_2061,In_425);
xnor U1688 (N_1688,In_1924,In_1465);
nor U1689 (N_1689,In_635,In_1199);
nand U1690 (N_1690,In_1941,In_818);
nor U1691 (N_1691,In_1863,In_417);
or U1692 (N_1692,In_666,In_2412);
xnor U1693 (N_1693,In_881,In_410);
or U1694 (N_1694,In_1869,In_2359);
xnor U1695 (N_1695,In_2367,In_978);
and U1696 (N_1696,In_277,In_273);
or U1697 (N_1697,In_704,In_538);
nand U1698 (N_1698,In_2183,In_1502);
xnor U1699 (N_1699,In_1770,In_2098);
nand U1700 (N_1700,In_493,In_381);
nor U1701 (N_1701,In_1849,In_693);
or U1702 (N_1702,In_1606,In_21);
nand U1703 (N_1703,In_283,In_639);
or U1704 (N_1704,In_1650,In_34);
and U1705 (N_1705,In_1848,In_1434);
or U1706 (N_1706,In_1695,In_1279);
nand U1707 (N_1707,In_518,In_568);
nand U1708 (N_1708,In_174,In_2427);
or U1709 (N_1709,In_1992,In_298);
nand U1710 (N_1710,In_668,In_1833);
nor U1711 (N_1711,In_2105,In_1146);
xnor U1712 (N_1712,In_1181,In_1295);
and U1713 (N_1713,In_1378,In_32);
nor U1714 (N_1714,In_347,In_1085);
xor U1715 (N_1715,In_1549,In_252);
or U1716 (N_1716,In_1539,In_1250);
or U1717 (N_1717,In_2332,In_279);
or U1718 (N_1718,In_759,In_268);
xnor U1719 (N_1719,In_282,In_1865);
nand U1720 (N_1720,In_1189,In_390);
xor U1721 (N_1721,In_1591,In_2277);
xnor U1722 (N_1722,In_732,In_1278);
nand U1723 (N_1723,In_1517,In_2119);
or U1724 (N_1724,In_941,In_2115);
or U1725 (N_1725,In_1424,In_479);
nand U1726 (N_1726,In_1063,In_1207);
nor U1727 (N_1727,In_727,In_509);
or U1728 (N_1728,In_661,In_282);
nor U1729 (N_1729,In_170,In_2414);
nand U1730 (N_1730,In_1990,In_1261);
nor U1731 (N_1731,In_2217,In_533);
xor U1732 (N_1732,In_25,In_2219);
nand U1733 (N_1733,In_1476,In_537);
nand U1734 (N_1734,In_118,In_2101);
nand U1735 (N_1735,In_496,In_834);
or U1736 (N_1736,In_578,In_516);
or U1737 (N_1737,In_582,In_2151);
xor U1738 (N_1738,In_108,In_854);
or U1739 (N_1739,In_657,In_1019);
and U1740 (N_1740,In_2187,In_1382);
and U1741 (N_1741,In_94,In_866);
and U1742 (N_1742,In_2344,In_388);
nand U1743 (N_1743,In_2400,In_396);
nand U1744 (N_1744,In_114,In_2381);
nor U1745 (N_1745,In_2084,In_120);
and U1746 (N_1746,In_1233,In_1729);
nor U1747 (N_1747,In_895,In_1131);
nor U1748 (N_1748,In_1033,In_760);
nor U1749 (N_1749,In_1565,In_2304);
nor U1750 (N_1750,In_1309,In_514);
and U1751 (N_1751,In_1177,In_1629);
xnor U1752 (N_1752,In_88,In_1352);
xnor U1753 (N_1753,In_546,In_1929);
nand U1754 (N_1754,In_1218,In_874);
and U1755 (N_1755,In_2446,In_182);
nor U1756 (N_1756,In_947,In_1321);
xor U1757 (N_1757,In_2355,In_2235);
xor U1758 (N_1758,In_1046,In_438);
or U1759 (N_1759,In_1338,In_1569);
and U1760 (N_1760,In_2358,In_2176);
and U1761 (N_1761,In_824,In_1898);
xor U1762 (N_1762,In_398,In_1213);
nor U1763 (N_1763,In_2323,In_1733);
nor U1764 (N_1764,In_180,In_89);
or U1765 (N_1765,In_1270,In_1121);
or U1766 (N_1766,In_2303,In_2366);
and U1767 (N_1767,In_2226,In_1327);
nor U1768 (N_1768,In_259,In_704);
xnor U1769 (N_1769,In_1804,In_1777);
and U1770 (N_1770,In_2181,In_1492);
nand U1771 (N_1771,In_270,In_826);
nand U1772 (N_1772,In_1105,In_2231);
xor U1773 (N_1773,In_940,In_1216);
nor U1774 (N_1774,In_1267,In_13);
xor U1775 (N_1775,In_92,In_17);
xnor U1776 (N_1776,In_2334,In_1577);
and U1777 (N_1777,In_1168,In_1239);
nor U1778 (N_1778,In_349,In_730);
nand U1779 (N_1779,In_1431,In_1241);
nor U1780 (N_1780,In_439,In_1214);
xnor U1781 (N_1781,In_1113,In_1061);
nor U1782 (N_1782,In_2387,In_1682);
nand U1783 (N_1783,In_755,In_2394);
nand U1784 (N_1784,In_22,In_2213);
nand U1785 (N_1785,In_1515,In_755);
nand U1786 (N_1786,In_684,In_3);
nand U1787 (N_1787,In_2123,In_1295);
xnor U1788 (N_1788,In_1543,In_1584);
and U1789 (N_1789,In_2406,In_1611);
nor U1790 (N_1790,In_664,In_192);
or U1791 (N_1791,In_1399,In_2104);
xor U1792 (N_1792,In_2253,In_1922);
or U1793 (N_1793,In_1118,In_2453);
xor U1794 (N_1794,In_1863,In_2133);
nand U1795 (N_1795,In_848,In_576);
nor U1796 (N_1796,In_933,In_226);
nor U1797 (N_1797,In_109,In_375);
or U1798 (N_1798,In_1961,In_1744);
or U1799 (N_1799,In_1602,In_656);
nor U1800 (N_1800,In_1831,In_2223);
nor U1801 (N_1801,In_319,In_793);
nor U1802 (N_1802,In_2118,In_1841);
nor U1803 (N_1803,In_119,In_1468);
nor U1804 (N_1804,In_1216,In_2217);
nand U1805 (N_1805,In_2415,In_318);
and U1806 (N_1806,In_973,In_86);
and U1807 (N_1807,In_1339,In_893);
xnor U1808 (N_1808,In_2384,In_1374);
nor U1809 (N_1809,In_2121,In_38);
or U1810 (N_1810,In_1311,In_474);
and U1811 (N_1811,In_676,In_687);
xnor U1812 (N_1812,In_1630,In_1062);
nor U1813 (N_1813,In_2004,In_791);
nor U1814 (N_1814,In_152,In_2184);
xnor U1815 (N_1815,In_572,In_1273);
and U1816 (N_1816,In_1649,In_1782);
xor U1817 (N_1817,In_1375,In_907);
xor U1818 (N_1818,In_1456,In_1158);
and U1819 (N_1819,In_363,In_193);
xor U1820 (N_1820,In_242,In_1499);
nor U1821 (N_1821,In_593,In_19);
and U1822 (N_1822,In_1377,In_1085);
xnor U1823 (N_1823,In_1785,In_1399);
xnor U1824 (N_1824,In_2119,In_2230);
and U1825 (N_1825,In_2312,In_141);
or U1826 (N_1826,In_2439,In_785);
nor U1827 (N_1827,In_760,In_1068);
nand U1828 (N_1828,In_2144,In_457);
nand U1829 (N_1829,In_682,In_1652);
and U1830 (N_1830,In_400,In_1667);
nand U1831 (N_1831,In_1289,In_1725);
xor U1832 (N_1832,In_1699,In_392);
xor U1833 (N_1833,In_1274,In_2344);
xnor U1834 (N_1834,In_1044,In_1751);
xnor U1835 (N_1835,In_1750,In_2162);
nand U1836 (N_1836,In_1300,In_2041);
and U1837 (N_1837,In_2488,In_882);
or U1838 (N_1838,In_1468,In_1077);
and U1839 (N_1839,In_1808,In_2125);
nand U1840 (N_1840,In_1872,In_174);
xor U1841 (N_1841,In_2273,In_2104);
nand U1842 (N_1842,In_2140,In_2242);
xor U1843 (N_1843,In_1403,In_526);
xor U1844 (N_1844,In_1867,In_949);
nand U1845 (N_1845,In_1388,In_1566);
and U1846 (N_1846,In_2268,In_2466);
nand U1847 (N_1847,In_630,In_1635);
nand U1848 (N_1848,In_1427,In_1811);
or U1849 (N_1849,In_214,In_1597);
or U1850 (N_1850,In_867,In_2239);
or U1851 (N_1851,In_114,In_1969);
xor U1852 (N_1852,In_148,In_2169);
and U1853 (N_1853,In_4,In_2054);
nand U1854 (N_1854,In_1509,In_530);
and U1855 (N_1855,In_395,In_1995);
and U1856 (N_1856,In_708,In_355);
and U1857 (N_1857,In_1441,In_517);
nor U1858 (N_1858,In_233,In_1332);
nor U1859 (N_1859,In_1138,In_1655);
xnor U1860 (N_1860,In_1606,In_1433);
or U1861 (N_1861,In_1685,In_428);
nor U1862 (N_1862,In_365,In_640);
nor U1863 (N_1863,In_1642,In_2021);
nor U1864 (N_1864,In_509,In_1468);
nor U1865 (N_1865,In_1278,In_147);
nor U1866 (N_1866,In_1043,In_210);
nand U1867 (N_1867,In_2243,In_607);
nor U1868 (N_1868,In_1382,In_434);
and U1869 (N_1869,In_840,In_156);
or U1870 (N_1870,In_1516,In_1845);
nand U1871 (N_1871,In_1274,In_1702);
xor U1872 (N_1872,In_474,In_2264);
nor U1873 (N_1873,In_1113,In_1634);
xnor U1874 (N_1874,In_1505,In_73);
nand U1875 (N_1875,In_302,In_909);
nand U1876 (N_1876,In_2016,In_573);
and U1877 (N_1877,In_1332,In_1649);
xnor U1878 (N_1878,In_876,In_1738);
nand U1879 (N_1879,In_905,In_2259);
nand U1880 (N_1880,In_399,In_904);
nor U1881 (N_1881,In_1346,In_1812);
xnor U1882 (N_1882,In_1692,In_679);
nand U1883 (N_1883,In_1757,In_1557);
xnor U1884 (N_1884,In_2171,In_1025);
and U1885 (N_1885,In_1312,In_2143);
or U1886 (N_1886,In_518,In_596);
or U1887 (N_1887,In_1740,In_1415);
or U1888 (N_1888,In_1103,In_463);
or U1889 (N_1889,In_1815,In_1927);
nand U1890 (N_1890,In_11,In_1122);
or U1891 (N_1891,In_2196,In_2250);
or U1892 (N_1892,In_1043,In_1337);
and U1893 (N_1893,In_69,In_807);
or U1894 (N_1894,In_2008,In_1882);
xnor U1895 (N_1895,In_1233,In_1016);
nor U1896 (N_1896,In_787,In_1349);
nand U1897 (N_1897,In_302,In_382);
nand U1898 (N_1898,In_1192,In_1856);
nand U1899 (N_1899,In_351,In_1732);
xor U1900 (N_1900,In_1987,In_1495);
xnor U1901 (N_1901,In_2036,In_2425);
and U1902 (N_1902,In_1461,In_1304);
and U1903 (N_1903,In_1169,In_1853);
xor U1904 (N_1904,In_1326,In_944);
nor U1905 (N_1905,In_2259,In_1972);
nor U1906 (N_1906,In_1772,In_1630);
and U1907 (N_1907,In_1138,In_1820);
or U1908 (N_1908,In_234,In_2001);
and U1909 (N_1909,In_1141,In_2443);
xnor U1910 (N_1910,In_2208,In_179);
nand U1911 (N_1911,In_292,In_2130);
or U1912 (N_1912,In_553,In_35);
xnor U1913 (N_1913,In_2336,In_1373);
nor U1914 (N_1914,In_2425,In_1900);
nand U1915 (N_1915,In_2101,In_1106);
xor U1916 (N_1916,In_2343,In_1792);
nor U1917 (N_1917,In_2033,In_746);
nor U1918 (N_1918,In_2321,In_1071);
or U1919 (N_1919,In_708,In_1273);
and U1920 (N_1920,In_1437,In_1430);
xor U1921 (N_1921,In_2486,In_2461);
nand U1922 (N_1922,In_868,In_1853);
or U1923 (N_1923,In_1058,In_407);
xor U1924 (N_1924,In_492,In_789);
and U1925 (N_1925,In_2040,In_2071);
nand U1926 (N_1926,In_2165,In_375);
and U1927 (N_1927,In_1291,In_259);
or U1928 (N_1928,In_2313,In_1758);
or U1929 (N_1929,In_440,In_1484);
nor U1930 (N_1930,In_2411,In_507);
nor U1931 (N_1931,In_1515,In_1431);
and U1932 (N_1932,In_1193,In_2377);
nand U1933 (N_1933,In_1828,In_1420);
or U1934 (N_1934,In_562,In_846);
nand U1935 (N_1935,In_580,In_1947);
nand U1936 (N_1936,In_2041,In_2008);
nor U1937 (N_1937,In_1423,In_1946);
or U1938 (N_1938,In_2128,In_1435);
or U1939 (N_1939,In_1208,In_1986);
and U1940 (N_1940,In_671,In_1521);
and U1941 (N_1941,In_877,In_982);
nor U1942 (N_1942,In_232,In_320);
and U1943 (N_1943,In_33,In_2286);
xnor U1944 (N_1944,In_1438,In_497);
or U1945 (N_1945,In_613,In_1730);
and U1946 (N_1946,In_1294,In_1744);
nand U1947 (N_1947,In_1839,In_2160);
or U1948 (N_1948,In_684,In_1642);
or U1949 (N_1949,In_2313,In_515);
nand U1950 (N_1950,In_2346,In_509);
nor U1951 (N_1951,In_199,In_53);
and U1952 (N_1952,In_2276,In_974);
xor U1953 (N_1953,In_1746,In_361);
nor U1954 (N_1954,In_53,In_2214);
and U1955 (N_1955,In_342,In_833);
nor U1956 (N_1956,In_796,In_823);
and U1957 (N_1957,In_2065,In_109);
xor U1958 (N_1958,In_1538,In_2233);
and U1959 (N_1959,In_2391,In_2264);
nand U1960 (N_1960,In_934,In_225);
nor U1961 (N_1961,In_2436,In_405);
and U1962 (N_1962,In_1822,In_1299);
xnor U1963 (N_1963,In_1596,In_484);
nor U1964 (N_1964,In_946,In_2231);
and U1965 (N_1965,In_2181,In_31);
nand U1966 (N_1966,In_534,In_1821);
nand U1967 (N_1967,In_37,In_1077);
nor U1968 (N_1968,In_1537,In_1687);
xnor U1969 (N_1969,In_374,In_1488);
and U1970 (N_1970,In_2029,In_1432);
or U1971 (N_1971,In_1106,In_87);
xnor U1972 (N_1972,In_1778,In_2431);
nor U1973 (N_1973,In_96,In_1834);
or U1974 (N_1974,In_1711,In_2081);
nand U1975 (N_1975,In_1813,In_323);
or U1976 (N_1976,In_990,In_1211);
xnor U1977 (N_1977,In_681,In_630);
xor U1978 (N_1978,In_1112,In_1649);
nand U1979 (N_1979,In_313,In_691);
xor U1980 (N_1980,In_983,In_493);
or U1981 (N_1981,In_1078,In_1378);
nor U1982 (N_1982,In_775,In_1104);
and U1983 (N_1983,In_683,In_1990);
or U1984 (N_1984,In_370,In_419);
and U1985 (N_1985,In_2223,In_947);
or U1986 (N_1986,In_216,In_159);
and U1987 (N_1987,In_1864,In_123);
xnor U1988 (N_1988,In_1100,In_598);
nor U1989 (N_1989,In_1768,In_2392);
nor U1990 (N_1990,In_317,In_1336);
xnor U1991 (N_1991,In_1697,In_2187);
xnor U1992 (N_1992,In_1987,In_2397);
and U1993 (N_1993,In_354,In_1071);
or U1994 (N_1994,In_350,In_903);
nor U1995 (N_1995,In_97,In_1268);
or U1996 (N_1996,In_1159,In_245);
or U1997 (N_1997,In_1312,In_1239);
nand U1998 (N_1998,In_2279,In_658);
nor U1999 (N_1999,In_795,In_1093);
xor U2000 (N_2000,In_829,In_1900);
nor U2001 (N_2001,In_121,In_1033);
and U2002 (N_2002,In_1299,In_2351);
xnor U2003 (N_2003,In_33,In_2321);
nand U2004 (N_2004,In_2024,In_589);
or U2005 (N_2005,In_194,In_2325);
nor U2006 (N_2006,In_2253,In_1678);
or U2007 (N_2007,In_2068,In_930);
nor U2008 (N_2008,In_2071,In_1196);
xor U2009 (N_2009,In_2454,In_1649);
nor U2010 (N_2010,In_1413,In_1039);
nor U2011 (N_2011,In_217,In_477);
nand U2012 (N_2012,In_1265,In_400);
nand U2013 (N_2013,In_814,In_544);
nand U2014 (N_2014,In_90,In_1057);
xnor U2015 (N_2015,In_701,In_202);
nand U2016 (N_2016,In_1206,In_1383);
and U2017 (N_2017,In_1601,In_926);
xnor U2018 (N_2018,In_2084,In_2036);
xor U2019 (N_2019,In_1580,In_101);
xnor U2020 (N_2020,In_1191,In_1904);
and U2021 (N_2021,In_1023,In_1412);
and U2022 (N_2022,In_1276,In_1378);
and U2023 (N_2023,In_965,In_2203);
and U2024 (N_2024,In_674,In_1897);
or U2025 (N_2025,In_1917,In_1637);
or U2026 (N_2026,In_1427,In_609);
nand U2027 (N_2027,In_709,In_210);
and U2028 (N_2028,In_557,In_2113);
or U2029 (N_2029,In_41,In_453);
nor U2030 (N_2030,In_561,In_2343);
nor U2031 (N_2031,In_540,In_1774);
or U2032 (N_2032,In_2321,In_956);
nor U2033 (N_2033,In_579,In_146);
or U2034 (N_2034,In_426,In_493);
or U2035 (N_2035,In_158,In_2212);
xor U2036 (N_2036,In_1757,In_1907);
xor U2037 (N_2037,In_1906,In_970);
xnor U2038 (N_2038,In_2424,In_2150);
and U2039 (N_2039,In_1229,In_717);
or U2040 (N_2040,In_1085,In_1699);
nand U2041 (N_2041,In_730,In_352);
xor U2042 (N_2042,In_568,In_2271);
and U2043 (N_2043,In_355,In_2246);
xnor U2044 (N_2044,In_1504,In_2013);
or U2045 (N_2045,In_1952,In_1630);
nor U2046 (N_2046,In_326,In_1663);
nand U2047 (N_2047,In_2292,In_502);
nand U2048 (N_2048,In_1446,In_2410);
nand U2049 (N_2049,In_1447,In_2030);
nor U2050 (N_2050,In_380,In_1897);
xnor U2051 (N_2051,In_967,In_1105);
or U2052 (N_2052,In_2357,In_92);
nor U2053 (N_2053,In_1215,In_1427);
nand U2054 (N_2054,In_1561,In_495);
nor U2055 (N_2055,In_1982,In_2052);
or U2056 (N_2056,In_1357,In_1407);
nand U2057 (N_2057,In_564,In_195);
nand U2058 (N_2058,In_1638,In_502);
nand U2059 (N_2059,In_2325,In_733);
nor U2060 (N_2060,In_1231,In_264);
and U2061 (N_2061,In_1987,In_1763);
or U2062 (N_2062,In_1765,In_561);
and U2063 (N_2063,In_662,In_1617);
nor U2064 (N_2064,In_1797,In_194);
nand U2065 (N_2065,In_1910,In_390);
nor U2066 (N_2066,In_2160,In_1243);
nand U2067 (N_2067,In_1798,In_2305);
nor U2068 (N_2068,In_273,In_2132);
or U2069 (N_2069,In_1997,In_313);
nand U2070 (N_2070,In_1814,In_1065);
xor U2071 (N_2071,In_1384,In_1080);
or U2072 (N_2072,In_1023,In_2226);
and U2073 (N_2073,In_836,In_534);
xor U2074 (N_2074,In_17,In_1289);
and U2075 (N_2075,In_308,In_164);
or U2076 (N_2076,In_1424,In_1580);
nand U2077 (N_2077,In_358,In_155);
nand U2078 (N_2078,In_102,In_2295);
xnor U2079 (N_2079,In_819,In_2325);
nor U2080 (N_2080,In_2210,In_657);
or U2081 (N_2081,In_1187,In_277);
xor U2082 (N_2082,In_662,In_1481);
nand U2083 (N_2083,In_922,In_1464);
or U2084 (N_2084,In_2439,In_1674);
or U2085 (N_2085,In_1189,In_1493);
or U2086 (N_2086,In_112,In_2318);
or U2087 (N_2087,In_914,In_1504);
and U2088 (N_2088,In_1117,In_1625);
nor U2089 (N_2089,In_2115,In_1004);
xor U2090 (N_2090,In_1368,In_545);
nand U2091 (N_2091,In_1772,In_971);
xnor U2092 (N_2092,In_1347,In_1137);
or U2093 (N_2093,In_884,In_536);
nor U2094 (N_2094,In_1787,In_1027);
and U2095 (N_2095,In_1277,In_2057);
nor U2096 (N_2096,In_783,In_1244);
and U2097 (N_2097,In_1874,In_750);
and U2098 (N_2098,In_1000,In_1797);
or U2099 (N_2099,In_174,In_1209);
and U2100 (N_2100,In_2384,In_1842);
or U2101 (N_2101,In_1906,In_242);
or U2102 (N_2102,In_899,In_1807);
nand U2103 (N_2103,In_701,In_1083);
nor U2104 (N_2104,In_1112,In_415);
and U2105 (N_2105,In_1161,In_1699);
nor U2106 (N_2106,In_891,In_475);
nand U2107 (N_2107,In_1586,In_1519);
xor U2108 (N_2108,In_749,In_445);
and U2109 (N_2109,In_7,In_710);
nand U2110 (N_2110,In_960,In_672);
or U2111 (N_2111,In_411,In_2005);
and U2112 (N_2112,In_2442,In_586);
and U2113 (N_2113,In_2245,In_1534);
nor U2114 (N_2114,In_1269,In_67);
nor U2115 (N_2115,In_339,In_2274);
nand U2116 (N_2116,In_637,In_652);
nand U2117 (N_2117,In_1596,In_432);
and U2118 (N_2118,In_1196,In_1438);
nor U2119 (N_2119,In_1114,In_1072);
nand U2120 (N_2120,In_1238,In_921);
nor U2121 (N_2121,In_1768,In_366);
nand U2122 (N_2122,In_1119,In_687);
xor U2123 (N_2123,In_1126,In_458);
and U2124 (N_2124,In_166,In_53);
or U2125 (N_2125,In_2155,In_1649);
nor U2126 (N_2126,In_1517,In_1803);
xor U2127 (N_2127,In_2111,In_1561);
and U2128 (N_2128,In_173,In_1136);
and U2129 (N_2129,In_1715,In_2428);
xor U2130 (N_2130,In_818,In_1296);
and U2131 (N_2131,In_945,In_817);
or U2132 (N_2132,In_1363,In_2316);
xor U2133 (N_2133,In_1732,In_758);
or U2134 (N_2134,In_1993,In_485);
nor U2135 (N_2135,In_477,In_1517);
nand U2136 (N_2136,In_2316,In_1020);
nor U2137 (N_2137,In_1220,In_2337);
xnor U2138 (N_2138,In_758,In_1571);
nand U2139 (N_2139,In_631,In_1797);
nor U2140 (N_2140,In_1657,In_1705);
xor U2141 (N_2141,In_1185,In_1193);
nand U2142 (N_2142,In_2310,In_1795);
and U2143 (N_2143,In_40,In_1844);
xnor U2144 (N_2144,In_297,In_682);
xor U2145 (N_2145,In_887,In_2094);
xor U2146 (N_2146,In_274,In_1931);
and U2147 (N_2147,In_1048,In_14);
or U2148 (N_2148,In_337,In_1604);
nand U2149 (N_2149,In_191,In_1619);
xnor U2150 (N_2150,In_633,In_2168);
xnor U2151 (N_2151,In_2070,In_2356);
nor U2152 (N_2152,In_51,In_1932);
and U2153 (N_2153,In_427,In_1091);
or U2154 (N_2154,In_1204,In_1368);
or U2155 (N_2155,In_2058,In_2130);
nor U2156 (N_2156,In_1277,In_768);
xnor U2157 (N_2157,In_912,In_638);
nor U2158 (N_2158,In_1378,In_364);
and U2159 (N_2159,In_560,In_2468);
and U2160 (N_2160,In_1693,In_78);
nor U2161 (N_2161,In_2483,In_2019);
nor U2162 (N_2162,In_779,In_2073);
and U2163 (N_2163,In_2056,In_1879);
xor U2164 (N_2164,In_463,In_402);
nand U2165 (N_2165,In_928,In_1786);
or U2166 (N_2166,In_1545,In_916);
or U2167 (N_2167,In_948,In_1801);
and U2168 (N_2168,In_777,In_1239);
xor U2169 (N_2169,In_1297,In_812);
xor U2170 (N_2170,In_2153,In_2426);
nor U2171 (N_2171,In_1341,In_1027);
nand U2172 (N_2172,In_278,In_2031);
and U2173 (N_2173,In_55,In_1849);
xnor U2174 (N_2174,In_1221,In_2468);
nand U2175 (N_2175,In_1552,In_517);
nand U2176 (N_2176,In_2021,In_1138);
nor U2177 (N_2177,In_454,In_2008);
or U2178 (N_2178,In_133,In_309);
and U2179 (N_2179,In_1795,In_307);
or U2180 (N_2180,In_753,In_2454);
and U2181 (N_2181,In_2035,In_2290);
nor U2182 (N_2182,In_59,In_58);
and U2183 (N_2183,In_1995,In_1655);
or U2184 (N_2184,In_825,In_530);
and U2185 (N_2185,In_35,In_701);
and U2186 (N_2186,In_455,In_1173);
xnor U2187 (N_2187,In_1327,In_1304);
nand U2188 (N_2188,In_850,In_2207);
nand U2189 (N_2189,In_504,In_2407);
nand U2190 (N_2190,In_954,In_124);
nand U2191 (N_2191,In_1024,In_478);
xor U2192 (N_2192,In_339,In_2108);
and U2193 (N_2193,In_1209,In_1815);
nand U2194 (N_2194,In_1441,In_333);
nand U2195 (N_2195,In_2460,In_582);
or U2196 (N_2196,In_610,In_41);
xnor U2197 (N_2197,In_1902,In_2022);
nor U2198 (N_2198,In_2286,In_1060);
xor U2199 (N_2199,In_369,In_1005);
nand U2200 (N_2200,In_2403,In_2167);
xor U2201 (N_2201,In_1667,In_2243);
nor U2202 (N_2202,In_2247,In_2321);
xnor U2203 (N_2203,In_421,In_1401);
xnor U2204 (N_2204,In_2438,In_1858);
xor U2205 (N_2205,In_967,In_1706);
and U2206 (N_2206,In_1573,In_147);
nand U2207 (N_2207,In_101,In_364);
or U2208 (N_2208,In_367,In_627);
xor U2209 (N_2209,In_251,In_1345);
and U2210 (N_2210,In_1090,In_1103);
nand U2211 (N_2211,In_1259,In_1239);
and U2212 (N_2212,In_1338,In_1161);
or U2213 (N_2213,In_2010,In_2001);
xnor U2214 (N_2214,In_1421,In_126);
xnor U2215 (N_2215,In_15,In_2437);
and U2216 (N_2216,In_208,In_482);
xnor U2217 (N_2217,In_532,In_1856);
nor U2218 (N_2218,In_344,In_1956);
nor U2219 (N_2219,In_1338,In_1260);
xnor U2220 (N_2220,In_677,In_701);
and U2221 (N_2221,In_1646,In_1596);
xnor U2222 (N_2222,In_2268,In_1146);
and U2223 (N_2223,In_249,In_1543);
or U2224 (N_2224,In_2121,In_842);
or U2225 (N_2225,In_2062,In_1682);
xor U2226 (N_2226,In_1056,In_1445);
and U2227 (N_2227,In_1389,In_1705);
nand U2228 (N_2228,In_409,In_69);
or U2229 (N_2229,In_335,In_1105);
nor U2230 (N_2230,In_382,In_2237);
xor U2231 (N_2231,In_347,In_2);
xor U2232 (N_2232,In_652,In_1988);
xnor U2233 (N_2233,In_510,In_2296);
nor U2234 (N_2234,In_2220,In_1550);
or U2235 (N_2235,In_885,In_893);
nand U2236 (N_2236,In_1824,In_1007);
or U2237 (N_2237,In_1137,In_1696);
xnor U2238 (N_2238,In_2044,In_1023);
nand U2239 (N_2239,In_680,In_430);
nor U2240 (N_2240,In_646,In_644);
nand U2241 (N_2241,In_878,In_2250);
or U2242 (N_2242,In_1729,In_1812);
nor U2243 (N_2243,In_1413,In_1983);
xnor U2244 (N_2244,In_1829,In_1111);
or U2245 (N_2245,In_1770,In_505);
or U2246 (N_2246,In_1365,In_909);
nor U2247 (N_2247,In_664,In_1623);
nor U2248 (N_2248,In_1811,In_41);
nor U2249 (N_2249,In_1947,In_2380);
xnor U2250 (N_2250,In_763,In_93);
xor U2251 (N_2251,In_941,In_539);
xor U2252 (N_2252,In_539,In_992);
xnor U2253 (N_2253,In_556,In_2063);
nand U2254 (N_2254,In_1444,In_1533);
xnor U2255 (N_2255,In_1089,In_662);
xor U2256 (N_2256,In_126,In_306);
or U2257 (N_2257,In_2397,In_1830);
nor U2258 (N_2258,In_1363,In_1063);
nor U2259 (N_2259,In_660,In_2428);
or U2260 (N_2260,In_1015,In_1176);
or U2261 (N_2261,In_1586,In_2294);
and U2262 (N_2262,In_1179,In_15);
xnor U2263 (N_2263,In_1219,In_1501);
nor U2264 (N_2264,In_2216,In_2339);
or U2265 (N_2265,In_1206,In_1288);
nand U2266 (N_2266,In_1401,In_1623);
xor U2267 (N_2267,In_1388,In_1631);
or U2268 (N_2268,In_370,In_1377);
nor U2269 (N_2269,In_2420,In_956);
xor U2270 (N_2270,In_53,In_556);
nand U2271 (N_2271,In_1790,In_1967);
and U2272 (N_2272,In_222,In_789);
or U2273 (N_2273,In_1077,In_2200);
nor U2274 (N_2274,In_1723,In_471);
nor U2275 (N_2275,In_1888,In_1447);
xor U2276 (N_2276,In_1364,In_2346);
nor U2277 (N_2277,In_628,In_1768);
or U2278 (N_2278,In_49,In_1799);
and U2279 (N_2279,In_2466,In_1001);
xnor U2280 (N_2280,In_1529,In_1015);
nor U2281 (N_2281,In_81,In_1379);
or U2282 (N_2282,In_750,In_2496);
nand U2283 (N_2283,In_662,In_705);
xor U2284 (N_2284,In_1213,In_294);
nor U2285 (N_2285,In_2411,In_265);
and U2286 (N_2286,In_481,In_1559);
nor U2287 (N_2287,In_585,In_1275);
nor U2288 (N_2288,In_1344,In_1930);
xnor U2289 (N_2289,In_2226,In_1951);
nand U2290 (N_2290,In_1318,In_399);
nor U2291 (N_2291,In_130,In_68);
nor U2292 (N_2292,In_1266,In_1785);
nor U2293 (N_2293,In_866,In_560);
and U2294 (N_2294,In_201,In_2477);
or U2295 (N_2295,In_1000,In_2215);
nor U2296 (N_2296,In_1229,In_1106);
nor U2297 (N_2297,In_2245,In_815);
nor U2298 (N_2298,In_587,In_522);
or U2299 (N_2299,In_806,In_915);
or U2300 (N_2300,In_865,In_1122);
and U2301 (N_2301,In_1084,In_626);
and U2302 (N_2302,In_1491,In_1569);
and U2303 (N_2303,In_2290,In_116);
xor U2304 (N_2304,In_678,In_1860);
xnor U2305 (N_2305,In_1679,In_614);
nand U2306 (N_2306,In_345,In_754);
and U2307 (N_2307,In_722,In_1044);
nand U2308 (N_2308,In_1499,In_714);
nor U2309 (N_2309,In_400,In_1726);
or U2310 (N_2310,In_1351,In_1428);
nor U2311 (N_2311,In_2162,In_1150);
or U2312 (N_2312,In_2303,In_2383);
nor U2313 (N_2313,In_296,In_538);
xor U2314 (N_2314,In_774,In_2183);
xor U2315 (N_2315,In_170,In_788);
xnor U2316 (N_2316,In_1185,In_2223);
and U2317 (N_2317,In_546,In_121);
and U2318 (N_2318,In_2173,In_337);
nor U2319 (N_2319,In_602,In_931);
xor U2320 (N_2320,In_2365,In_2095);
nand U2321 (N_2321,In_264,In_1699);
nand U2322 (N_2322,In_1746,In_671);
or U2323 (N_2323,In_1363,In_698);
and U2324 (N_2324,In_1650,In_2009);
nor U2325 (N_2325,In_2223,In_386);
and U2326 (N_2326,In_611,In_884);
nor U2327 (N_2327,In_712,In_1325);
xor U2328 (N_2328,In_1343,In_2402);
or U2329 (N_2329,In_877,In_1991);
nand U2330 (N_2330,In_765,In_1832);
or U2331 (N_2331,In_2275,In_790);
nand U2332 (N_2332,In_1988,In_2369);
nand U2333 (N_2333,In_1004,In_2095);
nor U2334 (N_2334,In_415,In_700);
xnor U2335 (N_2335,In_263,In_2370);
and U2336 (N_2336,In_1861,In_1508);
and U2337 (N_2337,In_1729,In_1036);
and U2338 (N_2338,In_1431,In_1051);
and U2339 (N_2339,In_1536,In_1419);
xnor U2340 (N_2340,In_389,In_464);
or U2341 (N_2341,In_927,In_1782);
nand U2342 (N_2342,In_2369,In_2290);
and U2343 (N_2343,In_793,In_1634);
or U2344 (N_2344,In_1363,In_775);
nand U2345 (N_2345,In_537,In_272);
or U2346 (N_2346,In_1603,In_1149);
or U2347 (N_2347,In_211,In_1695);
xor U2348 (N_2348,In_1808,In_1957);
nor U2349 (N_2349,In_1851,In_1383);
nand U2350 (N_2350,In_621,In_265);
and U2351 (N_2351,In_218,In_1323);
or U2352 (N_2352,In_249,In_1293);
or U2353 (N_2353,In_1203,In_1386);
nor U2354 (N_2354,In_1740,In_2335);
nand U2355 (N_2355,In_1285,In_1288);
or U2356 (N_2356,In_2451,In_2061);
and U2357 (N_2357,In_633,In_2089);
and U2358 (N_2358,In_1166,In_1113);
xor U2359 (N_2359,In_1296,In_970);
nor U2360 (N_2360,In_307,In_1206);
nor U2361 (N_2361,In_1393,In_266);
and U2362 (N_2362,In_2373,In_1428);
nor U2363 (N_2363,In_1388,In_1462);
xnor U2364 (N_2364,In_190,In_409);
and U2365 (N_2365,In_209,In_1336);
or U2366 (N_2366,In_626,In_1965);
nor U2367 (N_2367,In_2465,In_1225);
and U2368 (N_2368,In_168,In_2175);
nand U2369 (N_2369,In_2036,In_274);
xor U2370 (N_2370,In_1040,In_2026);
nand U2371 (N_2371,In_180,In_1961);
xnor U2372 (N_2372,In_409,In_765);
and U2373 (N_2373,In_632,In_2132);
or U2374 (N_2374,In_278,In_72);
nand U2375 (N_2375,In_867,In_1879);
nor U2376 (N_2376,In_2431,In_939);
and U2377 (N_2377,In_387,In_949);
xnor U2378 (N_2378,In_1374,In_68);
nand U2379 (N_2379,In_1817,In_1281);
nand U2380 (N_2380,In_220,In_535);
nand U2381 (N_2381,In_1950,In_2458);
and U2382 (N_2382,In_1599,In_198);
or U2383 (N_2383,In_2158,In_1342);
and U2384 (N_2384,In_189,In_55);
nand U2385 (N_2385,In_1697,In_2269);
nor U2386 (N_2386,In_298,In_1686);
nor U2387 (N_2387,In_304,In_676);
or U2388 (N_2388,In_572,In_1983);
nand U2389 (N_2389,In_1536,In_2196);
or U2390 (N_2390,In_2398,In_88);
xor U2391 (N_2391,In_578,In_240);
and U2392 (N_2392,In_219,In_983);
nor U2393 (N_2393,In_547,In_2265);
nor U2394 (N_2394,In_1516,In_1827);
nor U2395 (N_2395,In_1422,In_1595);
or U2396 (N_2396,In_419,In_1578);
or U2397 (N_2397,In_1791,In_404);
or U2398 (N_2398,In_1288,In_1609);
and U2399 (N_2399,In_25,In_239);
or U2400 (N_2400,In_1062,In_914);
xor U2401 (N_2401,In_1365,In_1220);
xnor U2402 (N_2402,In_646,In_2394);
or U2403 (N_2403,In_1597,In_349);
xnor U2404 (N_2404,In_1513,In_1735);
xnor U2405 (N_2405,In_2369,In_446);
and U2406 (N_2406,In_298,In_542);
xnor U2407 (N_2407,In_1081,In_1705);
nand U2408 (N_2408,In_1192,In_455);
xnor U2409 (N_2409,In_784,In_263);
xor U2410 (N_2410,In_625,In_1790);
or U2411 (N_2411,In_1134,In_2107);
xor U2412 (N_2412,In_2196,In_1815);
nor U2413 (N_2413,In_2148,In_452);
nor U2414 (N_2414,In_1917,In_1504);
nand U2415 (N_2415,In_932,In_1133);
and U2416 (N_2416,In_1524,In_87);
and U2417 (N_2417,In_375,In_2346);
xor U2418 (N_2418,In_178,In_1542);
xnor U2419 (N_2419,In_356,In_2348);
and U2420 (N_2420,In_1573,In_1026);
or U2421 (N_2421,In_1040,In_1358);
xnor U2422 (N_2422,In_2216,In_839);
or U2423 (N_2423,In_91,In_1427);
nand U2424 (N_2424,In_1388,In_2497);
nand U2425 (N_2425,In_805,In_1833);
or U2426 (N_2426,In_437,In_694);
nor U2427 (N_2427,In_1871,In_489);
xnor U2428 (N_2428,In_2322,In_383);
xnor U2429 (N_2429,In_1831,In_957);
xnor U2430 (N_2430,In_576,In_1494);
xor U2431 (N_2431,In_110,In_516);
nor U2432 (N_2432,In_1039,In_770);
nor U2433 (N_2433,In_2298,In_109);
xnor U2434 (N_2434,In_567,In_752);
xor U2435 (N_2435,In_625,In_586);
nor U2436 (N_2436,In_1562,In_1593);
or U2437 (N_2437,In_1656,In_1943);
and U2438 (N_2438,In_441,In_1835);
nor U2439 (N_2439,In_1384,In_10);
nor U2440 (N_2440,In_1236,In_849);
or U2441 (N_2441,In_2302,In_2458);
nor U2442 (N_2442,In_2022,In_1119);
xnor U2443 (N_2443,In_732,In_1244);
and U2444 (N_2444,In_1327,In_456);
nor U2445 (N_2445,In_621,In_1514);
and U2446 (N_2446,In_880,In_1617);
and U2447 (N_2447,In_952,In_1417);
nand U2448 (N_2448,In_1833,In_880);
nor U2449 (N_2449,In_713,In_1652);
nand U2450 (N_2450,In_20,In_244);
nor U2451 (N_2451,In_1967,In_1301);
xnor U2452 (N_2452,In_532,In_2181);
xnor U2453 (N_2453,In_1448,In_1080);
or U2454 (N_2454,In_1256,In_555);
or U2455 (N_2455,In_69,In_379);
or U2456 (N_2456,In_1924,In_1282);
and U2457 (N_2457,In_229,In_64);
xnor U2458 (N_2458,In_2264,In_863);
nor U2459 (N_2459,In_1511,In_1101);
xor U2460 (N_2460,In_1647,In_2128);
and U2461 (N_2461,In_718,In_887);
nor U2462 (N_2462,In_2222,In_882);
nand U2463 (N_2463,In_555,In_1505);
xor U2464 (N_2464,In_2466,In_1279);
nand U2465 (N_2465,In_1937,In_439);
nor U2466 (N_2466,In_2036,In_2);
nand U2467 (N_2467,In_1676,In_150);
nand U2468 (N_2468,In_97,In_387);
nor U2469 (N_2469,In_2117,In_1838);
xnor U2470 (N_2470,In_1807,In_448);
and U2471 (N_2471,In_1964,In_2242);
nor U2472 (N_2472,In_339,In_1880);
and U2473 (N_2473,In_1807,In_1126);
nand U2474 (N_2474,In_1588,In_1130);
nor U2475 (N_2475,In_1069,In_781);
and U2476 (N_2476,In_2446,In_914);
xnor U2477 (N_2477,In_2018,In_888);
or U2478 (N_2478,In_685,In_715);
nand U2479 (N_2479,In_801,In_2211);
nor U2480 (N_2480,In_1153,In_288);
nor U2481 (N_2481,In_447,In_1406);
nand U2482 (N_2482,In_498,In_1727);
or U2483 (N_2483,In_272,In_892);
nand U2484 (N_2484,In_1648,In_1285);
xor U2485 (N_2485,In_137,In_2176);
nand U2486 (N_2486,In_1749,In_89);
nand U2487 (N_2487,In_2160,In_72);
or U2488 (N_2488,In_990,In_1322);
nor U2489 (N_2489,In_1220,In_665);
or U2490 (N_2490,In_796,In_1573);
and U2491 (N_2491,In_1754,In_188);
or U2492 (N_2492,In_2039,In_2048);
nor U2493 (N_2493,In_1654,In_2346);
and U2494 (N_2494,In_1683,In_2047);
xnor U2495 (N_2495,In_2400,In_1814);
nand U2496 (N_2496,In_1196,In_287);
nor U2497 (N_2497,In_597,In_1723);
nand U2498 (N_2498,In_143,In_124);
nor U2499 (N_2499,In_1226,In_630);
and U2500 (N_2500,In_604,In_1070);
xnor U2501 (N_2501,In_110,In_534);
nand U2502 (N_2502,In_124,In_2250);
or U2503 (N_2503,In_1365,In_1448);
xnor U2504 (N_2504,In_939,In_2201);
or U2505 (N_2505,In_276,In_49);
nand U2506 (N_2506,In_1710,In_1867);
and U2507 (N_2507,In_733,In_2217);
xnor U2508 (N_2508,In_2390,In_1988);
or U2509 (N_2509,In_1635,In_2323);
nand U2510 (N_2510,In_679,In_1259);
nand U2511 (N_2511,In_209,In_1920);
xor U2512 (N_2512,In_2135,In_2395);
and U2513 (N_2513,In_2246,In_2157);
or U2514 (N_2514,In_54,In_2189);
or U2515 (N_2515,In_650,In_584);
xor U2516 (N_2516,In_2492,In_755);
xor U2517 (N_2517,In_275,In_816);
or U2518 (N_2518,In_1229,In_1774);
nor U2519 (N_2519,In_934,In_1061);
and U2520 (N_2520,In_62,In_120);
or U2521 (N_2521,In_1589,In_1437);
or U2522 (N_2522,In_2009,In_251);
nand U2523 (N_2523,In_266,In_2176);
and U2524 (N_2524,In_1185,In_1153);
nand U2525 (N_2525,In_661,In_315);
or U2526 (N_2526,In_635,In_2173);
xnor U2527 (N_2527,In_1980,In_1081);
nor U2528 (N_2528,In_2288,In_1904);
or U2529 (N_2529,In_842,In_1209);
and U2530 (N_2530,In_539,In_178);
nor U2531 (N_2531,In_1551,In_2499);
xor U2532 (N_2532,In_156,In_395);
nand U2533 (N_2533,In_282,In_477);
or U2534 (N_2534,In_610,In_370);
xor U2535 (N_2535,In_1632,In_1637);
nor U2536 (N_2536,In_1552,In_1352);
or U2537 (N_2537,In_1366,In_1358);
and U2538 (N_2538,In_1664,In_982);
nand U2539 (N_2539,In_2350,In_1925);
xor U2540 (N_2540,In_417,In_312);
nor U2541 (N_2541,In_2017,In_2491);
or U2542 (N_2542,In_2152,In_33);
xor U2543 (N_2543,In_273,In_1417);
or U2544 (N_2544,In_350,In_2112);
and U2545 (N_2545,In_1185,In_68);
or U2546 (N_2546,In_18,In_710);
nor U2547 (N_2547,In_831,In_2234);
nor U2548 (N_2548,In_2285,In_358);
nor U2549 (N_2549,In_1566,In_1258);
or U2550 (N_2550,In_1075,In_2022);
xor U2551 (N_2551,In_1559,In_1691);
nor U2552 (N_2552,In_1254,In_920);
or U2553 (N_2553,In_1679,In_1413);
xor U2554 (N_2554,In_452,In_319);
nor U2555 (N_2555,In_1993,In_1933);
xnor U2556 (N_2556,In_1322,In_1250);
xor U2557 (N_2557,In_1390,In_543);
and U2558 (N_2558,In_1779,In_1557);
nor U2559 (N_2559,In_159,In_1925);
xnor U2560 (N_2560,In_322,In_1227);
or U2561 (N_2561,In_1315,In_1608);
nor U2562 (N_2562,In_2073,In_747);
xnor U2563 (N_2563,In_1518,In_48);
xor U2564 (N_2564,In_1644,In_282);
xor U2565 (N_2565,In_1526,In_2401);
nor U2566 (N_2566,In_113,In_1908);
or U2567 (N_2567,In_92,In_269);
or U2568 (N_2568,In_2198,In_713);
nor U2569 (N_2569,In_1654,In_551);
nand U2570 (N_2570,In_574,In_1660);
or U2571 (N_2571,In_1266,In_454);
xnor U2572 (N_2572,In_341,In_37);
nand U2573 (N_2573,In_266,In_431);
or U2574 (N_2574,In_1521,In_1467);
and U2575 (N_2575,In_1165,In_1059);
or U2576 (N_2576,In_2108,In_321);
or U2577 (N_2577,In_1699,In_1654);
nand U2578 (N_2578,In_1500,In_358);
and U2579 (N_2579,In_336,In_282);
or U2580 (N_2580,In_1139,In_128);
xor U2581 (N_2581,In_523,In_2160);
nor U2582 (N_2582,In_1744,In_1674);
and U2583 (N_2583,In_1093,In_2224);
nor U2584 (N_2584,In_1187,In_953);
xnor U2585 (N_2585,In_1319,In_612);
xor U2586 (N_2586,In_828,In_846);
nand U2587 (N_2587,In_2095,In_1921);
nand U2588 (N_2588,In_1148,In_2082);
nor U2589 (N_2589,In_1078,In_1723);
or U2590 (N_2590,In_219,In_111);
or U2591 (N_2591,In_1910,In_2301);
and U2592 (N_2592,In_2207,In_429);
and U2593 (N_2593,In_1494,In_165);
nor U2594 (N_2594,In_1453,In_1858);
xor U2595 (N_2595,In_725,In_1703);
xnor U2596 (N_2596,In_1522,In_2106);
xor U2597 (N_2597,In_302,In_1530);
nand U2598 (N_2598,In_1206,In_1121);
nor U2599 (N_2599,In_934,In_2455);
nor U2600 (N_2600,In_282,In_2081);
nand U2601 (N_2601,In_1288,In_1432);
and U2602 (N_2602,In_2143,In_257);
nand U2603 (N_2603,In_320,In_1979);
nand U2604 (N_2604,In_5,In_1415);
and U2605 (N_2605,In_371,In_1437);
xnor U2606 (N_2606,In_2379,In_1981);
and U2607 (N_2607,In_2183,In_697);
xor U2608 (N_2608,In_1427,In_737);
or U2609 (N_2609,In_1573,In_782);
or U2610 (N_2610,In_1118,In_1069);
nand U2611 (N_2611,In_1450,In_760);
nor U2612 (N_2612,In_1021,In_1373);
nand U2613 (N_2613,In_1409,In_534);
nand U2614 (N_2614,In_387,In_324);
xor U2615 (N_2615,In_459,In_2204);
nand U2616 (N_2616,In_815,In_692);
nand U2617 (N_2617,In_1661,In_1407);
nand U2618 (N_2618,In_1791,In_1540);
nor U2619 (N_2619,In_1199,In_390);
or U2620 (N_2620,In_5,In_39);
and U2621 (N_2621,In_1688,In_132);
or U2622 (N_2622,In_835,In_726);
nor U2623 (N_2623,In_1434,In_525);
xnor U2624 (N_2624,In_468,In_932);
or U2625 (N_2625,In_1098,In_1409);
xnor U2626 (N_2626,In_907,In_1299);
xor U2627 (N_2627,In_1083,In_1440);
and U2628 (N_2628,In_511,In_1603);
or U2629 (N_2629,In_1245,In_6);
nand U2630 (N_2630,In_2119,In_1449);
and U2631 (N_2631,In_161,In_520);
or U2632 (N_2632,In_2284,In_2427);
and U2633 (N_2633,In_1042,In_1171);
nor U2634 (N_2634,In_1603,In_531);
xnor U2635 (N_2635,In_1098,In_823);
and U2636 (N_2636,In_366,In_809);
or U2637 (N_2637,In_1765,In_697);
and U2638 (N_2638,In_788,In_518);
and U2639 (N_2639,In_2354,In_1130);
and U2640 (N_2640,In_1109,In_2256);
or U2641 (N_2641,In_944,In_678);
nand U2642 (N_2642,In_74,In_2423);
and U2643 (N_2643,In_1463,In_1284);
or U2644 (N_2644,In_830,In_578);
nor U2645 (N_2645,In_2059,In_1587);
xnor U2646 (N_2646,In_2449,In_1690);
nor U2647 (N_2647,In_746,In_332);
xnor U2648 (N_2648,In_651,In_126);
or U2649 (N_2649,In_1982,In_14);
or U2650 (N_2650,In_339,In_771);
nor U2651 (N_2651,In_2287,In_945);
and U2652 (N_2652,In_1762,In_1225);
or U2653 (N_2653,In_46,In_762);
nand U2654 (N_2654,In_184,In_1237);
and U2655 (N_2655,In_600,In_350);
nand U2656 (N_2656,In_716,In_587);
or U2657 (N_2657,In_904,In_1590);
nand U2658 (N_2658,In_823,In_261);
xnor U2659 (N_2659,In_102,In_1566);
or U2660 (N_2660,In_73,In_2254);
and U2661 (N_2661,In_1492,In_1452);
nand U2662 (N_2662,In_1101,In_2003);
nand U2663 (N_2663,In_1046,In_2095);
or U2664 (N_2664,In_20,In_861);
xor U2665 (N_2665,In_1927,In_2273);
nor U2666 (N_2666,In_578,In_2032);
or U2667 (N_2667,In_1114,In_2030);
or U2668 (N_2668,In_1714,In_1636);
xor U2669 (N_2669,In_1217,In_1490);
nor U2670 (N_2670,In_1759,In_374);
nor U2671 (N_2671,In_396,In_1361);
and U2672 (N_2672,In_1026,In_859);
nand U2673 (N_2673,In_527,In_2045);
nand U2674 (N_2674,In_1577,In_1788);
and U2675 (N_2675,In_1489,In_401);
and U2676 (N_2676,In_2009,In_198);
and U2677 (N_2677,In_1259,In_2447);
nand U2678 (N_2678,In_75,In_2466);
and U2679 (N_2679,In_2031,In_2483);
and U2680 (N_2680,In_1127,In_801);
and U2681 (N_2681,In_349,In_1883);
and U2682 (N_2682,In_584,In_1347);
and U2683 (N_2683,In_581,In_2027);
or U2684 (N_2684,In_844,In_147);
xnor U2685 (N_2685,In_1770,In_1086);
and U2686 (N_2686,In_1953,In_2339);
and U2687 (N_2687,In_2234,In_1568);
xor U2688 (N_2688,In_1892,In_2095);
or U2689 (N_2689,In_1121,In_1405);
nor U2690 (N_2690,In_1218,In_2217);
nor U2691 (N_2691,In_192,In_267);
nand U2692 (N_2692,In_1276,In_586);
nand U2693 (N_2693,In_619,In_1102);
or U2694 (N_2694,In_2424,In_1105);
and U2695 (N_2695,In_654,In_1852);
nor U2696 (N_2696,In_2247,In_516);
nand U2697 (N_2697,In_707,In_278);
or U2698 (N_2698,In_262,In_1124);
and U2699 (N_2699,In_1756,In_1763);
nor U2700 (N_2700,In_1116,In_1685);
nor U2701 (N_2701,In_2032,In_571);
and U2702 (N_2702,In_2078,In_2344);
nand U2703 (N_2703,In_1665,In_1217);
xnor U2704 (N_2704,In_1439,In_235);
xor U2705 (N_2705,In_586,In_662);
nand U2706 (N_2706,In_1036,In_843);
xnor U2707 (N_2707,In_2078,In_1808);
xnor U2708 (N_2708,In_2391,In_2090);
or U2709 (N_2709,In_44,In_1164);
nor U2710 (N_2710,In_2229,In_2427);
or U2711 (N_2711,In_2401,In_509);
xnor U2712 (N_2712,In_645,In_2067);
nor U2713 (N_2713,In_1199,In_939);
nand U2714 (N_2714,In_2141,In_1257);
nor U2715 (N_2715,In_491,In_1239);
and U2716 (N_2716,In_326,In_2);
nand U2717 (N_2717,In_2238,In_813);
nand U2718 (N_2718,In_1729,In_2195);
nor U2719 (N_2719,In_1242,In_2458);
nand U2720 (N_2720,In_1849,In_1348);
nand U2721 (N_2721,In_2477,In_2498);
nor U2722 (N_2722,In_646,In_711);
xor U2723 (N_2723,In_1688,In_1539);
or U2724 (N_2724,In_2432,In_975);
nand U2725 (N_2725,In_877,In_2162);
xnor U2726 (N_2726,In_843,In_53);
and U2727 (N_2727,In_590,In_1351);
and U2728 (N_2728,In_897,In_1633);
xnor U2729 (N_2729,In_1505,In_580);
nor U2730 (N_2730,In_1033,In_1369);
nand U2731 (N_2731,In_568,In_1565);
xnor U2732 (N_2732,In_1773,In_851);
nor U2733 (N_2733,In_1229,In_550);
nand U2734 (N_2734,In_534,In_12);
and U2735 (N_2735,In_741,In_911);
nor U2736 (N_2736,In_886,In_180);
nor U2737 (N_2737,In_2268,In_891);
nor U2738 (N_2738,In_169,In_739);
nor U2739 (N_2739,In_94,In_2290);
or U2740 (N_2740,In_1606,In_339);
xnor U2741 (N_2741,In_907,In_2344);
or U2742 (N_2742,In_579,In_743);
and U2743 (N_2743,In_955,In_2168);
nor U2744 (N_2744,In_2116,In_488);
and U2745 (N_2745,In_33,In_1891);
nand U2746 (N_2746,In_503,In_820);
xnor U2747 (N_2747,In_2117,In_250);
and U2748 (N_2748,In_790,In_765);
nor U2749 (N_2749,In_68,In_1580);
xnor U2750 (N_2750,In_665,In_197);
xor U2751 (N_2751,In_455,In_2012);
or U2752 (N_2752,In_1396,In_690);
or U2753 (N_2753,In_2455,In_2470);
or U2754 (N_2754,In_1834,In_1851);
nor U2755 (N_2755,In_2484,In_627);
nor U2756 (N_2756,In_1723,In_311);
and U2757 (N_2757,In_2437,In_1264);
nor U2758 (N_2758,In_2270,In_2032);
nand U2759 (N_2759,In_934,In_1771);
nor U2760 (N_2760,In_2048,In_2163);
and U2761 (N_2761,In_1701,In_970);
xor U2762 (N_2762,In_394,In_2126);
and U2763 (N_2763,In_2477,In_2111);
nand U2764 (N_2764,In_1166,In_1811);
and U2765 (N_2765,In_1860,In_1833);
xnor U2766 (N_2766,In_253,In_1702);
xor U2767 (N_2767,In_1883,In_327);
or U2768 (N_2768,In_678,In_964);
xnor U2769 (N_2769,In_1624,In_1160);
nor U2770 (N_2770,In_1904,In_121);
nor U2771 (N_2771,In_2356,In_996);
nand U2772 (N_2772,In_113,In_1087);
nand U2773 (N_2773,In_18,In_430);
xnor U2774 (N_2774,In_2227,In_1913);
nor U2775 (N_2775,In_239,In_2336);
nor U2776 (N_2776,In_581,In_1028);
nor U2777 (N_2777,In_209,In_1313);
nand U2778 (N_2778,In_508,In_1260);
xnor U2779 (N_2779,In_369,In_2451);
or U2780 (N_2780,In_2090,In_324);
nand U2781 (N_2781,In_2455,In_964);
and U2782 (N_2782,In_1622,In_264);
nor U2783 (N_2783,In_2007,In_2104);
and U2784 (N_2784,In_1877,In_1106);
nand U2785 (N_2785,In_964,In_59);
or U2786 (N_2786,In_751,In_1204);
nand U2787 (N_2787,In_1946,In_143);
nand U2788 (N_2788,In_881,In_807);
and U2789 (N_2789,In_1122,In_2009);
xor U2790 (N_2790,In_319,In_739);
and U2791 (N_2791,In_849,In_1979);
or U2792 (N_2792,In_2344,In_1024);
xnor U2793 (N_2793,In_13,In_2465);
nand U2794 (N_2794,In_1865,In_2451);
xor U2795 (N_2795,In_1818,In_147);
and U2796 (N_2796,In_1792,In_83);
nand U2797 (N_2797,In_2233,In_1663);
or U2798 (N_2798,In_1850,In_990);
and U2799 (N_2799,In_581,In_1074);
and U2800 (N_2800,In_2006,In_22);
nor U2801 (N_2801,In_409,In_399);
nor U2802 (N_2802,In_801,In_642);
nand U2803 (N_2803,In_2224,In_318);
nand U2804 (N_2804,In_1231,In_1326);
nand U2805 (N_2805,In_935,In_217);
nor U2806 (N_2806,In_575,In_2033);
or U2807 (N_2807,In_2051,In_566);
nand U2808 (N_2808,In_1312,In_2352);
or U2809 (N_2809,In_1497,In_943);
nand U2810 (N_2810,In_1693,In_1723);
nand U2811 (N_2811,In_2039,In_1778);
or U2812 (N_2812,In_99,In_1564);
nand U2813 (N_2813,In_360,In_629);
and U2814 (N_2814,In_294,In_945);
xor U2815 (N_2815,In_1494,In_1337);
and U2816 (N_2816,In_1258,In_1921);
or U2817 (N_2817,In_399,In_1413);
and U2818 (N_2818,In_462,In_1022);
and U2819 (N_2819,In_2176,In_1926);
nor U2820 (N_2820,In_1375,In_211);
nand U2821 (N_2821,In_2239,In_414);
nand U2822 (N_2822,In_1608,In_2103);
and U2823 (N_2823,In_318,In_910);
nor U2824 (N_2824,In_1634,In_743);
nand U2825 (N_2825,In_98,In_3);
nor U2826 (N_2826,In_847,In_598);
nor U2827 (N_2827,In_1005,In_1908);
nor U2828 (N_2828,In_1193,In_854);
nor U2829 (N_2829,In_1910,In_291);
or U2830 (N_2830,In_1768,In_295);
xnor U2831 (N_2831,In_702,In_575);
xnor U2832 (N_2832,In_1663,In_2426);
nor U2833 (N_2833,In_133,In_72);
xnor U2834 (N_2834,In_784,In_902);
xnor U2835 (N_2835,In_1282,In_1478);
xor U2836 (N_2836,In_509,In_2055);
xnor U2837 (N_2837,In_425,In_303);
or U2838 (N_2838,In_286,In_2457);
xor U2839 (N_2839,In_1483,In_2440);
or U2840 (N_2840,In_188,In_576);
nand U2841 (N_2841,In_1174,In_1436);
nand U2842 (N_2842,In_2091,In_2190);
nor U2843 (N_2843,In_69,In_1189);
or U2844 (N_2844,In_1549,In_1985);
xor U2845 (N_2845,In_2479,In_2139);
or U2846 (N_2846,In_1760,In_191);
nor U2847 (N_2847,In_132,In_2495);
nor U2848 (N_2848,In_2255,In_2499);
nor U2849 (N_2849,In_1537,In_2066);
xnor U2850 (N_2850,In_712,In_42);
and U2851 (N_2851,In_714,In_190);
or U2852 (N_2852,In_665,In_2257);
nand U2853 (N_2853,In_548,In_1087);
nor U2854 (N_2854,In_1904,In_439);
nor U2855 (N_2855,In_1555,In_761);
or U2856 (N_2856,In_2111,In_1210);
and U2857 (N_2857,In_1717,In_641);
xor U2858 (N_2858,In_1406,In_1904);
xnor U2859 (N_2859,In_2428,In_422);
and U2860 (N_2860,In_228,In_1962);
and U2861 (N_2861,In_1514,In_1390);
nand U2862 (N_2862,In_117,In_620);
nor U2863 (N_2863,In_441,In_1421);
xnor U2864 (N_2864,In_1299,In_1197);
xor U2865 (N_2865,In_1688,In_1283);
and U2866 (N_2866,In_669,In_51);
or U2867 (N_2867,In_992,In_2064);
nor U2868 (N_2868,In_1174,In_580);
nand U2869 (N_2869,In_283,In_1359);
or U2870 (N_2870,In_1287,In_2414);
nand U2871 (N_2871,In_1908,In_1802);
nor U2872 (N_2872,In_719,In_2164);
or U2873 (N_2873,In_1177,In_2300);
nor U2874 (N_2874,In_1159,In_1179);
or U2875 (N_2875,In_2155,In_449);
nand U2876 (N_2876,In_781,In_409);
or U2877 (N_2877,In_1914,In_965);
nor U2878 (N_2878,In_1374,In_1903);
nand U2879 (N_2879,In_1726,In_2409);
nor U2880 (N_2880,In_2380,In_1207);
nor U2881 (N_2881,In_1583,In_1215);
nor U2882 (N_2882,In_905,In_2367);
nand U2883 (N_2883,In_1791,In_1684);
xnor U2884 (N_2884,In_1528,In_1726);
or U2885 (N_2885,In_1271,In_1211);
nand U2886 (N_2886,In_1846,In_163);
nand U2887 (N_2887,In_1188,In_2421);
and U2888 (N_2888,In_347,In_2483);
nor U2889 (N_2889,In_53,In_299);
or U2890 (N_2890,In_1606,In_1334);
nor U2891 (N_2891,In_2101,In_2179);
and U2892 (N_2892,In_480,In_2330);
nand U2893 (N_2893,In_979,In_2278);
and U2894 (N_2894,In_343,In_679);
or U2895 (N_2895,In_2395,In_1994);
xnor U2896 (N_2896,In_210,In_1978);
and U2897 (N_2897,In_1272,In_1415);
or U2898 (N_2898,In_724,In_900);
xor U2899 (N_2899,In_999,In_1967);
and U2900 (N_2900,In_2090,In_2007);
or U2901 (N_2901,In_812,In_1656);
nand U2902 (N_2902,In_2279,In_1680);
or U2903 (N_2903,In_1384,In_839);
and U2904 (N_2904,In_2306,In_2231);
or U2905 (N_2905,In_273,In_677);
nand U2906 (N_2906,In_1605,In_2343);
nor U2907 (N_2907,In_996,In_969);
nor U2908 (N_2908,In_337,In_2057);
or U2909 (N_2909,In_694,In_2297);
xnor U2910 (N_2910,In_1640,In_224);
nor U2911 (N_2911,In_539,In_1298);
or U2912 (N_2912,In_167,In_580);
nor U2913 (N_2913,In_662,In_319);
and U2914 (N_2914,In_2443,In_2273);
or U2915 (N_2915,In_775,In_1552);
nand U2916 (N_2916,In_556,In_88);
or U2917 (N_2917,In_2069,In_379);
nor U2918 (N_2918,In_1714,In_9);
or U2919 (N_2919,In_2490,In_1511);
nand U2920 (N_2920,In_1175,In_294);
nand U2921 (N_2921,In_972,In_1177);
xor U2922 (N_2922,In_1346,In_273);
or U2923 (N_2923,In_283,In_1562);
nor U2924 (N_2924,In_1102,In_548);
nor U2925 (N_2925,In_1237,In_2098);
nor U2926 (N_2926,In_646,In_1652);
nand U2927 (N_2927,In_2275,In_921);
xor U2928 (N_2928,In_1367,In_346);
nand U2929 (N_2929,In_430,In_2155);
or U2930 (N_2930,In_2211,In_1040);
xnor U2931 (N_2931,In_1301,In_1604);
xor U2932 (N_2932,In_1189,In_2029);
xor U2933 (N_2933,In_846,In_272);
or U2934 (N_2934,In_1879,In_583);
nand U2935 (N_2935,In_1733,In_1314);
nand U2936 (N_2936,In_797,In_1906);
and U2937 (N_2937,In_1724,In_88);
xor U2938 (N_2938,In_832,In_176);
and U2939 (N_2939,In_2342,In_186);
or U2940 (N_2940,In_1014,In_283);
nand U2941 (N_2941,In_1679,In_573);
nor U2942 (N_2942,In_2069,In_2208);
nor U2943 (N_2943,In_937,In_1054);
and U2944 (N_2944,In_2450,In_370);
or U2945 (N_2945,In_226,In_1117);
nor U2946 (N_2946,In_2342,In_763);
nor U2947 (N_2947,In_80,In_1147);
xnor U2948 (N_2948,In_2018,In_1992);
xor U2949 (N_2949,In_1533,In_2050);
and U2950 (N_2950,In_1595,In_2137);
nand U2951 (N_2951,In_130,In_1310);
xor U2952 (N_2952,In_405,In_1689);
xor U2953 (N_2953,In_838,In_851);
nand U2954 (N_2954,In_272,In_1320);
nand U2955 (N_2955,In_1194,In_1387);
nor U2956 (N_2956,In_560,In_16);
nor U2957 (N_2957,In_2036,In_810);
xor U2958 (N_2958,In_84,In_136);
and U2959 (N_2959,In_370,In_1216);
nor U2960 (N_2960,In_2157,In_593);
or U2961 (N_2961,In_1383,In_861);
nor U2962 (N_2962,In_1105,In_2229);
nor U2963 (N_2963,In_890,In_1511);
or U2964 (N_2964,In_2115,In_1416);
nor U2965 (N_2965,In_197,In_1340);
or U2966 (N_2966,In_600,In_90);
nand U2967 (N_2967,In_1403,In_1150);
xor U2968 (N_2968,In_1923,In_2495);
nor U2969 (N_2969,In_806,In_1826);
nor U2970 (N_2970,In_458,In_1843);
and U2971 (N_2971,In_2144,In_2404);
or U2972 (N_2972,In_1614,In_650);
xor U2973 (N_2973,In_1285,In_1130);
xnor U2974 (N_2974,In_409,In_1436);
and U2975 (N_2975,In_705,In_2122);
nor U2976 (N_2976,In_111,In_1182);
nand U2977 (N_2977,In_1683,In_1122);
nor U2978 (N_2978,In_1131,In_1782);
xnor U2979 (N_2979,In_1727,In_1009);
nand U2980 (N_2980,In_586,In_2029);
nor U2981 (N_2981,In_72,In_1181);
nor U2982 (N_2982,In_1460,In_2397);
xor U2983 (N_2983,In_1832,In_202);
nand U2984 (N_2984,In_400,In_1432);
nor U2985 (N_2985,In_910,In_2290);
xor U2986 (N_2986,In_89,In_1546);
nand U2987 (N_2987,In_1581,In_808);
xor U2988 (N_2988,In_1929,In_1007);
nand U2989 (N_2989,In_12,In_430);
nor U2990 (N_2990,In_416,In_1172);
xor U2991 (N_2991,In_1800,In_1136);
and U2992 (N_2992,In_356,In_2026);
xor U2993 (N_2993,In_850,In_102);
nand U2994 (N_2994,In_1686,In_2268);
or U2995 (N_2995,In_2106,In_362);
nor U2996 (N_2996,In_1250,In_986);
xor U2997 (N_2997,In_134,In_2456);
nor U2998 (N_2998,In_2247,In_120);
nor U2999 (N_2999,In_119,In_921);
nand U3000 (N_3000,In_278,In_1677);
and U3001 (N_3001,In_683,In_2076);
nor U3002 (N_3002,In_2008,In_174);
and U3003 (N_3003,In_1237,In_576);
nor U3004 (N_3004,In_2106,In_186);
or U3005 (N_3005,In_881,In_525);
nand U3006 (N_3006,In_1361,In_893);
nor U3007 (N_3007,In_2301,In_1626);
nor U3008 (N_3008,In_2405,In_731);
xor U3009 (N_3009,In_17,In_1776);
nand U3010 (N_3010,In_2049,In_1407);
nand U3011 (N_3011,In_1203,In_1613);
and U3012 (N_3012,In_1809,In_40);
nor U3013 (N_3013,In_1174,In_537);
or U3014 (N_3014,In_910,In_537);
xnor U3015 (N_3015,In_733,In_382);
and U3016 (N_3016,In_628,In_1889);
xnor U3017 (N_3017,In_876,In_61);
nor U3018 (N_3018,In_1421,In_1808);
xnor U3019 (N_3019,In_1411,In_692);
nand U3020 (N_3020,In_236,In_846);
and U3021 (N_3021,In_1697,In_1733);
and U3022 (N_3022,In_2289,In_617);
nand U3023 (N_3023,In_1409,In_454);
nor U3024 (N_3024,In_2341,In_2470);
nand U3025 (N_3025,In_2025,In_521);
nor U3026 (N_3026,In_80,In_351);
nand U3027 (N_3027,In_1408,In_530);
xor U3028 (N_3028,In_1415,In_211);
nor U3029 (N_3029,In_1062,In_1245);
or U3030 (N_3030,In_2081,In_2077);
nand U3031 (N_3031,In_253,In_231);
or U3032 (N_3032,In_2437,In_779);
xnor U3033 (N_3033,In_1946,In_1192);
nand U3034 (N_3034,In_529,In_962);
xnor U3035 (N_3035,In_2135,In_1765);
nor U3036 (N_3036,In_2050,In_1060);
nor U3037 (N_3037,In_27,In_163);
nor U3038 (N_3038,In_126,In_1383);
or U3039 (N_3039,In_835,In_468);
nand U3040 (N_3040,In_155,In_696);
nor U3041 (N_3041,In_2162,In_905);
nor U3042 (N_3042,In_720,In_914);
xor U3043 (N_3043,In_627,In_1915);
or U3044 (N_3044,In_1791,In_1278);
xor U3045 (N_3045,In_269,In_1717);
nand U3046 (N_3046,In_2027,In_1206);
xnor U3047 (N_3047,In_1230,In_1133);
xor U3048 (N_3048,In_491,In_1646);
nand U3049 (N_3049,In_272,In_691);
or U3050 (N_3050,In_965,In_817);
or U3051 (N_3051,In_1126,In_2062);
or U3052 (N_3052,In_1406,In_1932);
xor U3053 (N_3053,In_564,In_1473);
and U3054 (N_3054,In_1796,In_1862);
and U3055 (N_3055,In_2071,In_1715);
or U3056 (N_3056,In_2421,In_1078);
xnor U3057 (N_3057,In_1509,In_1544);
nor U3058 (N_3058,In_2267,In_1690);
xnor U3059 (N_3059,In_2439,In_190);
nor U3060 (N_3060,In_532,In_284);
and U3061 (N_3061,In_1780,In_680);
xor U3062 (N_3062,In_1439,In_1688);
xnor U3063 (N_3063,In_1495,In_551);
or U3064 (N_3064,In_186,In_2085);
xnor U3065 (N_3065,In_727,In_1810);
nand U3066 (N_3066,In_2352,In_841);
xnor U3067 (N_3067,In_1770,In_2258);
and U3068 (N_3068,In_1172,In_455);
or U3069 (N_3069,In_1638,In_1810);
nor U3070 (N_3070,In_1428,In_1128);
xor U3071 (N_3071,In_1100,In_377);
or U3072 (N_3072,In_2148,In_1584);
nor U3073 (N_3073,In_1658,In_1605);
nor U3074 (N_3074,In_570,In_904);
xor U3075 (N_3075,In_2356,In_1217);
nor U3076 (N_3076,In_2398,In_1233);
or U3077 (N_3077,In_1054,In_1468);
or U3078 (N_3078,In_110,In_2316);
or U3079 (N_3079,In_1085,In_1011);
and U3080 (N_3080,In_701,In_1809);
and U3081 (N_3081,In_1121,In_1356);
or U3082 (N_3082,In_544,In_568);
nand U3083 (N_3083,In_657,In_488);
and U3084 (N_3084,In_2376,In_2093);
nand U3085 (N_3085,In_821,In_376);
and U3086 (N_3086,In_2315,In_1984);
nor U3087 (N_3087,In_2472,In_1402);
or U3088 (N_3088,In_2059,In_1631);
and U3089 (N_3089,In_2427,In_281);
xor U3090 (N_3090,In_2466,In_1600);
xor U3091 (N_3091,In_881,In_2486);
and U3092 (N_3092,In_577,In_477);
xnor U3093 (N_3093,In_184,In_2488);
nand U3094 (N_3094,In_2416,In_1963);
nand U3095 (N_3095,In_2031,In_1023);
nor U3096 (N_3096,In_198,In_2222);
or U3097 (N_3097,In_1371,In_250);
and U3098 (N_3098,In_1015,In_1789);
or U3099 (N_3099,In_1558,In_579);
nand U3100 (N_3100,In_728,In_541);
xnor U3101 (N_3101,In_2358,In_1570);
and U3102 (N_3102,In_561,In_1390);
or U3103 (N_3103,In_1016,In_1188);
or U3104 (N_3104,In_1991,In_1383);
or U3105 (N_3105,In_225,In_1391);
or U3106 (N_3106,In_1557,In_1694);
nand U3107 (N_3107,In_172,In_170);
nand U3108 (N_3108,In_501,In_1322);
nor U3109 (N_3109,In_921,In_2350);
or U3110 (N_3110,In_852,In_1347);
nand U3111 (N_3111,In_1976,In_2480);
xor U3112 (N_3112,In_1193,In_366);
nand U3113 (N_3113,In_2167,In_1063);
nor U3114 (N_3114,In_2029,In_1628);
and U3115 (N_3115,In_1369,In_2196);
nor U3116 (N_3116,In_2414,In_1891);
or U3117 (N_3117,In_213,In_880);
nor U3118 (N_3118,In_886,In_2493);
xor U3119 (N_3119,In_766,In_2438);
xnor U3120 (N_3120,In_696,In_740);
and U3121 (N_3121,In_430,In_932);
xnor U3122 (N_3122,In_1965,In_2392);
xor U3123 (N_3123,In_1198,In_211);
nand U3124 (N_3124,In_1784,In_1412);
nor U3125 (N_3125,N_1834,N_310);
or U3126 (N_3126,N_423,N_2647);
nor U3127 (N_3127,N_1076,N_1072);
xnor U3128 (N_3128,N_2192,N_2215);
or U3129 (N_3129,N_2404,N_2528);
nand U3130 (N_3130,N_945,N_1039);
or U3131 (N_3131,N_348,N_234);
or U3132 (N_3132,N_1276,N_3093);
and U3133 (N_3133,N_2257,N_1503);
or U3134 (N_3134,N_827,N_1677);
nand U3135 (N_3135,N_1051,N_1931);
and U3136 (N_3136,N_216,N_2115);
xnor U3137 (N_3137,N_1242,N_867);
or U3138 (N_3138,N_2961,N_2889);
nor U3139 (N_3139,N_1544,N_1794);
nand U3140 (N_3140,N_1690,N_2207);
or U3141 (N_3141,N_3066,N_1380);
or U3142 (N_3142,N_682,N_2332);
and U3143 (N_3143,N_1762,N_1118);
nor U3144 (N_3144,N_613,N_703);
and U3145 (N_3145,N_2414,N_695);
or U3146 (N_3146,N_1841,N_670);
nand U3147 (N_3147,N_2034,N_1129);
xnor U3148 (N_3148,N_453,N_2331);
nor U3149 (N_3149,N_1732,N_2452);
xor U3150 (N_3150,N_1650,N_2521);
nor U3151 (N_3151,N_2083,N_3046);
nor U3152 (N_3152,N_865,N_1100);
nor U3153 (N_3153,N_2727,N_1054);
or U3154 (N_3154,N_757,N_1745);
xor U3155 (N_3155,N_491,N_1562);
nand U3156 (N_3156,N_2847,N_17);
nand U3157 (N_3157,N_1969,N_1226);
or U3158 (N_3158,N_2478,N_2537);
or U3159 (N_3159,N_2976,N_2305);
xnor U3160 (N_3160,N_1678,N_1481);
nor U3161 (N_3161,N_242,N_1000);
xor U3162 (N_3162,N_967,N_1556);
or U3163 (N_3163,N_2206,N_2068);
nor U3164 (N_3164,N_1087,N_1924);
xor U3165 (N_3165,N_1530,N_718);
and U3166 (N_3166,N_590,N_1236);
nand U3167 (N_3167,N_2916,N_2669);
nand U3168 (N_3168,N_2686,N_306);
nand U3169 (N_3169,N_3035,N_1784);
or U3170 (N_3170,N_155,N_1894);
and U3171 (N_3171,N_959,N_2822);
xnor U3172 (N_3172,N_10,N_2360);
and U3173 (N_3173,N_2955,N_136);
or U3174 (N_3174,N_298,N_2952);
nor U3175 (N_3175,N_2935,N_2598);
xnor U3176 (N_3176,N_968,N_1662);
nand U3177 (N_3177,N_924,N_2557);
or U3178 (N_3178,N_475,N_557);
nand U3179 (N_3179,N_2433,N_773);
xnor U3180 (N_3180,N_1336,N_1608);
nand U3181 (N_3181,N_50,N_1280);
nor U3182 (N_3182,N_2474,N_1714);
and U3183 (N_3183,N_434,N_1907);
or U3184 (N_3184,N_2428,N_3028);
nor U3185 (N_3185,N_2698,N_1793);
nor U3186 (N_3186,N_2202,N_544);
or U3187 (N_3187,N_189,N_1009);
or U3188 (N_3188,N_3088,N_2562);
nor U3189 (N_3189,N_1861,N_327);
or U3190 (N_3190,N_2405,N_828);
and U3191 (N_3191,N_1422,N_1399);
and U3192 (N_3192,N_2185,N_1539);
nor U3193 (N_3193,N_848,N_2074);
nor U3194 (N_3194,N_631,N_2133);
and U3195 (N_3195,N_1059,N_2431);
nand U3196 (N_3196,N_1810,N_283);
nor U3197 (N_3197,N_368,N_846);
nand U3198 (N_3198,N_1642,N_2888);
and U3199 (N_3199,N_742,N_1141);
nor U3200 (N_3200,N_320,N_2760);
nor U3201 (N_3201,N_2950,N_122);
and U3202 (N_3202,N_82,N_1869);
nor U3203 (N_3203,N_984,N_2212);
xor U3204 (N_3204,N_2210,N_179);
and U3205 (N_3205,N_1484,N_204);
nand U3206 (N_3206,N_2560,N_173);
xnor U3207 (N_3207,N_1990,N_1575);
xor U3208 (N_3208,N_2366,N_861);
or U3209 (N_3209,N_2132,N_450);
and U3210 (N_3210,N_1876,N_2681);
nor U3211 (N_3211,N_1055,N_1030);
nor U3212 (N_3212,N_352,N_547);
nor U3213 (N_3213,N_3026,N_2939);
nor U3214 (N_3214,N_151,N_738);
nor U3215 (N_3215,N_1047,N_2788);
nand U3216 (N_3216,N_958,N_812);
and U3217 (N_3217,N_2350,N_796);
or U3218 (N_3218,N_2846,N_1266);
and U3219 (N_3219,N_1023,N_885);
or U3220 (N_3220,N_2737,N_2188);
and U3221 (N_3221,N_3075,N_2695);
or U3222 (N_3222,N_2195,N_676);
or U3223 (N_3223,N_85,N_272);
and U3224 (N_3224,N_1623,N_1614);
nand U3225 (N_3225,N_2714,N_2593);
nor U3226 (N_3226,N_473,N_42);
or U3227 (N_3227,N_728,N_2403);
xor U3228 (N_3228,N_1361,N_3098);
nand U3229 (N_3229,N_1154,N_2694);
nand U3230 (N_3230,N_2777,N_2325);
nor U3231 (N_3231,N_1597,N_1081);
xnor U3232 (N_3232,N_2757,N_2592);
nand U3233 (N_3233,N_2584,N_585);
or U3234 (N_3234,N_1582,N_1884);
nor U3235 (N_3235,N_2928,N_2143);
and U3236 (N_3236,N_1769,N_1619);
and U3237 (N_3237,N_747,N_1148);
and U3238 (N_3238,N_312,N_2527);
xnor U3239 (N_3239,N_1557,N_2774);
nand U3240 (N_3240,N_2545,N_1203);
or U3241 (N_3241,N_595,N_2796);
nand U3242 (N_3242,N_2627,N_1167);
nor U3243 (N_3243,N_2067,N_1808);
or U3244 (N_3244,N_79,N_2178);
nand U3245 (N_3245,N_2785,N_3071);
xor U3246 (N_3246,N_1815,N_607);
nand U3247 (N_3247,N_369,N_1947);
nor U3248 (N_3248,N_1408,N_1574);
xor U3249 (N_3249,N_2026,N_142);
or U3250 (N_3250,N_1913,N_1656);
xor U3251 (N_3251,N_560,N_3103);
nor U3252 (N_3252,N_1162,N_981);
and U3253 (N_3253,N_2589,N_2709);
or U3254 (N_3254,N_183,N_1938);
xor U3255 (N_3255,N_1112,N_1842);
nor U3256 (N_3256,N_233,N_1144);
nand U3257 (N_3257,N_1653,N_1818);
nand U3258 (N_3258,N_2493,N_2089);
nand U3259 (N_3259,N_2055,N_1865);
nand U3260 (N_3260,N_2073,N_2851);
xor U3261 (N_3261,N_2021,N_2652);
nand U3262 (N_3262,N_530,N_292);
or U3263 (N_3263,N_688,N_3116);
nor U3264 (N_3264,N_144,N_2665);
and U3265 (N_3265,N_2276,N_1224);
xor U3266 (N_3266,N_1331,N_208);
or U3267 (N_3267,N_1168,N_668);
xor U3268 (N_3268,N_1528,N_328);
or U3269 (N_3269,N_1795,N_2158);
nand U3270 (N_3270,N_1026,N_806);
and U3271 (N_3271,N_2632,N_1968);
and U3272 (N_3272,N_1560,N_1073);
xor U3273 (N_3273,N_1207,N_2876);
xnor U3274 (N_3274,N_2603,N_2313);
xor U3275 (N_3275,N_2731,N_1731);
xor U3276 (N_3276,N_58,N_2138);
xnor U3277 (N_3277,N_3003,N_1123);
nor U3278 (N_3278,N_1074,N_158);
or U3279 (N_3279,N_3091,N_3045);
or U3280 (N_3280,N_2969,N_2062);
nor U3281 (N_3281,N_1812,N_2582);
and U3282 (N_3282,N_3086,N_790);
and U3283 (N_3283,N_2800,N_2135);
xor U3284 (N_3284,N_337,N_1259);
nor U3285 (N_3285,N_197,N_1857);
xnor U3286 (N_3286,N_1316,N_513);
and U3287 (N_3287,N_1724,N_2358);
or U3288 (N_3288,N_316,N_2623);
or U3289 (N_3289,N_1668,N_1327);
or U3290 (N_3290,N_3019,N_2836);
or U3291 (N_3291,N_830,N_553);
xnor U3292 (N_3292,N_1751,N_1358);
and U3293 (N_3293,N_1944,N_933);
nor U3294 (N_3294,N_148,N_2444);
and U3295 (N_3295,N_236,N_2136);
xnor U3296 (N_3296,N_115,N_159);
xnor U3297 (N_3297,N_3070,N_2465);
nor U3298 (N_3298,N_1634,N_874);
nand U3299 (N_3299,N_594,N_97);
nor U3300 (N_3300,N_1282,N_521);
nor U3301 (N_3301,N_3033,N_1015);
and U3302 (N_3302,N_2372,N_1521);
xor U3303 (N_3303,N_531,N_1204);
nor U3304 (N_3304,N_2570,N_1791);
nor U3305 (N_3305,N_2490,N_2124);
xor U3306 (N_3306,N_3117,N_819);
nor U3307 (N_3307,N_1273,N_200);
nor U3308 (N_3308,N_2738,N_1723);
and U3309 (N_3309,N_226,N_2112);
and U3310 (N_3310,N_2586,N_2713);
nand U3311 (N_3311,N_1355,N_1993);
xor U3312 (N_3312,N_1719,N_105);
xor U3313 (N_3313,N_1255,N_1488);
or U3314 (N_3314,N_3011,N_350);
nor U3315 (N_3315,N_1237,N_411);
nor U3316 (N_3316,N_1752,N_2007);
and U3317 (N_3317,N_811,N_1500);
and U3318 (N_3318,N_2919,N_510);
nor U3319 (N_3319,N_534,N_894);
or U3320 (N_3320,N_1285,N_660);
or U3321 (N_3321,N_744,N_3085);
nor U3322 (N_3322,N_537,N_2349);
or U3323 (N_3323,N_2640,N_232);
xor U3324 (N_3324,N_1421,N_1542);
or U3325 (N_3325,N_1624,N_1104);
and U3326 (N_3326,N_2411,N_2913);
nand U3327 (N_3327,N_2538,N_3015);
or U3328 (N_3328,N_1502,N_2971);
or U3329 (N_3329,N_1048,N_2753);
and U3330 (N_3330,N_1707,N_460);
nor U3331 (N_3331,N_2575,N_418);
and U3332 (N_3332,N_931,N_302);
nor U3333 (N_3333,N_2381,N_2259);
nor U3334 (N_3334,N_223,N_224);
xor U3335 (N_3335,N_1197,N_3067);
and U3336 (N_3336,N_2687,N_1753);
nand U3337 (N_3337,N_414,N_363);
nand U3338 (N_3338,N_624,N_509);
xnor U3339 (N_3339,N_2447,N_1790);
xor U3340 (N_3340,N_2953,N_3054);
nor U3341 (N_3341,N_57,N_1314);
and U3342 (N_3342,N_2535,N_2364);
nor U3343 (N_3343,N_2013,N_2689);
nor U3344 (N_3344,N_55,N_2701);
or U3345 (N_3345,N_1457,N_504);
xnor U3346 (N_3346,N_1786,N_113);
nor U3347 (N_3347,N_943,N_1549);
and U3348 (N_3348,N_2253,N_2371);
and U3349 (N_3349,N_2036,N_30);
nor U3350 (N_3350,N_1291,N_2790);
and U3351 (N_3351,N_2131,N_1710);
xnor U3352 (N_3352,N_722,N_3021);
xnor U3353 (N_3353,N_215,N_2100);
xnor U3354 (N_3354,N_3030,N_2455);
or U3355 (N_3355,N_1417,N_1238);
nor U3356 (N_3356,N_2732,N_1366);
and U3357 (N_3357,N_1407,N_2972);
nand U3358 (N_3358,N_571,N_1078);
nor U3359 (N_3359,N_1892,N_1700);
nand U3360 (N_3360,N_2284,N_1085);
nor U3361 (N_3361,N_1288,N_195);
or U3362 (N_3362,N_1778,N_2436);
nor U3363 (N_3363,N_2715,N_1367);
xor U3364 (N_3364,N_1587,N_2962);
nor U3365 (N_3365,N_2235,N_1183);
and U3366 (N_3366,N_3059,N_2311);
nor U3367 (N_3367,N_381,N_1836);
nor U3368 (N_3368,N_2032,N_290);
or U3369 (N_3369,N_225,N_2384);
xor U3370 (N_3370,N_2984,N_2921);
nand U3371 (N_3371,N_1979,N_3051);
or U3372 (N_3372,N_1303,N_1832);
xnor U3373 (N_3373,N_2064,N_1186);
xor U3374 (N_3374,N_1974,N_1086);
or U3375 (N_3375,N_634,N_1362);
xor U3376 (N_3376,N_2113,N_1837);
or U3377 (N_3377,N_1669,N_386);
or U3378 (N_3378,N_743,N_1915);
nor U3379 (N_3379,N_2053,N_291);
nand U3380 (N_3380,N_1657,N_755);
nand U3381 (N_3381,N_2617,N_3002);
nand U3382 (N_3382,N_2407,N_2469);
xnor U3383 (N_3383,N_459,N_2883);
xor U3384 (N_3384,N_2168,N_12);
nand U3385 (N_3385,N_338,N_2383);
or U3386 (N_3386,N_2502,N_1935);
xnor U3387 (N_3387,N_1701,N_1694);
and U3388 (N_3388,N_2967,N_2045);
or U3389 (N_3389,N_2837,N_2227);
xnor U3390 (N_3390,N_487,N_3050);
and U3391 (N_3391,N_1191,N_1532);
xnor U3392 (N_3392,N_2905,N_1982);
xnor U3393 (N_3393,N_2515,N_34);
or U3394 (N_3394,N_2468,N_2056);
xnor U3395 (N_3395,N_2862,N_376);
nand U3396 (N_3396,N_648,N_205);
nor U3397 (N_3397,N_2223,N_1340);
and U3398 (N_3398,N_2000,N_2659);
nor U3399 (N_3399,N_1391,N_870);
and U3400 (N_3400,N_2925,N_1430);
nand U3401 (N_3401,N_2075,N_1729);
nor U3402 (N_3402,N_2492,N_45);
nor U3403 (N_3403,N_2773,N_2899);
xor U3404 (N_3404,N_1205,N_987);
and U3405 (N_3405,N_791,N_1056);
and U3406 (N_3406,N_3121,N_1216);
nor U3407 (N_3407,N_3065,N_1089);
xnor U3408 (N_3408,N_1372,N_1595);
or U3409 (N_3409,N_145,N_13);
xor U3410 (N_3410,N_564,N_1965);
nand U3411 (N_3411,N_2475,N_2375);
nand U3412 (N_3412,N_2299,N_1010);
and U3413 (N_3413,N_813,N_2173);
xnor U3414 (N_3414,N_3100,N_3009);
nor U3415 (N_3415,N_156,N_2496);
nand U3416 (N_3416,N_734,N_2674);
xnor U3417 (N_3417,N_11,N_431);
xor U3418 (N_3418,N_857,N_1149);
xnor U3419 (N_3419,N_2139,N_446);
nor U3420 (N_3420,N_696,N_253);
nand U3421 (N_3421,N_1275,N_1737);
or U3422 (N_3422,N_1838,N_977);
and U3423 (N_3423,N_2618,N_18);
nor U3424 (N_3424,N_2278,N_96);
nand U3425 (N_3425,N_3052,N_889);
xor U3426 (N_3426,N_1647,N_355);
or U3427 (N_3427,N_1501,N_1166);
nand U3428 (N_3428,N_726,N_2038);
xor U3429 (N_3429,N_1526,N_1802);
nand U3430 (N_3430,N_367,N_2301);
nand U3431 (N_3431,N_1598,N_2164);
nand U3432 (N_3432,N_1559,N_763);
xnor U3433 (N_3433,N_212,N_90);
or U3434 (N_3434,N_3076,N_2480);
xor U3435 (N_3435,N_2323,N_1651);
and U3436 (N_3436,N_1515,N_1290);
and U3437 (N_3437,N_2711,N_230);
xnor U3438 (N_3438,N_2230,N_1635);
or U3439 (N_3439,N_927,N_323);
and U3440 (N_3440,N_821,N_2606);
or U3441 (N_3441,N_3041,N_1696);
xor U3442 (N_3442,N_1001,N_714);
nor U3443 (N_3443,N_1214,N_2427);
nand U3444 (N_3444,N_3037,N_2547);
nand U3445 (N_3445,N_497,N_1561);
xnor U3446 (N_3446,N_2690,N_1767);
nor U3447 (N_3447,N_1992,N_1171);
or U3448 (N_3448,N_63,N_1264);
and U3449 (N_3449,N_1016,N_991);
xnor U3450 (N_3450,N_2426,N_2927);
xnor U3451 (N_3451,N_2109,N_3027);
nor U3452 (N_3452,N_206,N_2569);
or U3453 (N_3453,N_725,N_1995);
nand U3454 (N_3454,N_997,N_3007);
nand U3455 (N_3455,N_797,N_972);
or U3456 (N_3456,N_1411,N_702);
and U3457 (N_3457,N_3048,N_2146);
nor U3458 (N_3458,N_617,N_1017);
and U3459 (N_3459,N_1375,N_31);
nor U3460 (N_3460,N_1736,N_3064);
nor U3461 (N_3461,N_853,N_1024);
xnor U3462 (N_3462,N_2848,N_1486);
xnor U3463 (N_3463,N_2079,N_149);
or U3464 (N_3464,N_3084,N_238);
xnor U3465 (N_3465,N_1493,N_2450);
and U3466 (N_3466,N_1828,N_2126);
nand U3467 (N_3467,N_2845,N_2033);
or U3468 (N_3468,N_745,N_787);
nor U3469 (N_3469,N_3113,N_103);
xnor U3470 (N_3470,N_915,N_2550);
and U3471 (N_3471,N_400,N_831);
or U3472 (N_3472,N_217,N_1343);
xor U3473 (N_3473,N_1579,N_3031);
nand U3474 (N_3474,N_2890,N_604);
nand U3475 (N_3475,N_2050,N_2499);
and U3476 (N_3476,N_667,N_1035);
or U3477 (N_3477,N_2887,N_1543);
nand U3478 (N_3478,N_2319,N_265);
xnor U3479 (N_3479,N_1441,N_603);
xnor U3480 (N_3480,N_1936,N_1458);
nor U3481 (N_3481,N_2746,N_1202);
xor U3482 (N_3482,N_425,N_1322);
nor U3483 (N_3483,N_1052,N_772);
or U3484 (N_3484,N_2051,N_1269);
or U3485 (N_3485,N_599,N_1178);
or U3486 (N_3486,N_2810,N_199);
or U3487 (N_3487,N_731,N_1512);
and U3488 (N_3488,N_656,N_1354);
nand U3489 (N_3489,N_1094,N_371);
nand U3490 (N_3490,N_1856,N_2965);
or U3491 (N_3491,N_2802,N_2438);
or U3492 (N_3492,N_1325,N_1095);
or U3493 (N_3493,N_168,N_228);
nor U3494 (N_3494,N_2183,N_880);
or U3495 (N_3495,N_1849,N_2997);
xnor U3496 (N_3496,N_1041,N_626);
xor U3497 (N_3497,N_3080,N_2662);
or U3498 (N_3498,N_454,N_289);
nand U3499 (N_3499,N_2645,N_2816);
xor U3500 (N_3500,N_808,N_2565);
nor U3501 (N_3501,N_691,N_1402);
and U3502 (N_3502,N_519,N_1212);
nor U3503 (N_3503,N_1703,N_2811);
nor U3504 (N_3504,N_250,N_508);
and U3505 (N_3505,N_588,N_740);
and U3506 (N_3506,N_2260,N_2915);
xnor U3507 (N_3507,N_960,N_1064);
xnor U3508 (N_3508,N_1092,N_466);
xor U3509 (N_3509,N_2957,N_1955);
or U3510 (N_3510,N_1676,N_782);
nor U3511 (N_3511,N_789,N_1644);
nand U3512 (N_3512,N_2680,N_137);
or U3513 (N_3513,N_2642,N_429);
and U3514 (N_3514,N_1169,N_2162);
nand U3515 (N_3515,N_1612,N_1939);
xnor U3516 (N_3516,N_2147,N_334);
nand U3517 (N_3517,N_3092,N_51);
and U3518 (N_3518,N_946,N_1855);
nor U3519 (N_3519,N_1188,N_2236);
and U3520 (N_3520,N_1444,N_107);
or U3521 (N_3521,N_1760,N_1545);
xnor U3522 (N_3522,N_2893,N_264);
nor U3523 (N_3523,N_1378,N_858);
and U3524 (N_3524,N_1179,N_1899);
or U3525 (N_3525,N_175,N_2076);
and U3526 (N_3526,N_1195,N_1840);
nand U3527 (N_3527,N_1406,N_1240);
nand U3528 (N_3528,N_1413,N_207);
nor U3529 (N_3529,N_1241,N_124);
xnor U3530 (N_3530,N_563,N_441);
or U3531 (N_3531,N_1514,N_655);
nand U3532 (N_3532,N_2599,N_980);
or U3533 (N_3533,N_1210,N_820);
xor U3534 (N_3534,N_930,N_176);
xnor U3535 (N_3535,N_1415,N_2548);
nor U3536 (N_3536,N_1431,N_282);
xor U3537 (N_3537,N_1022,N_2318);
nand U3538 (N_3538,N_1117,N_1629);
and U3539 (N_3539,N_1034,N_1495);
xor U3540 (N_3540,N_93,N_2445);
nand U3541 (N_3541,N_2166,N_1593);
and U3542 (N_3542,N_1172,N_1305);
xor U3543 (N_3543,N_2370,N_1872);
or U3544 (N_3544,N_374,N_2664);
or U3545 (N_3545,N_1230,N_3104);
and U3546 (N_3546,N_2010,N_1005);
and U3547 (N_3547,N_1972,N_1875);
or U3548 (N_3548,N_2351,N_221);
nand U3549 (N_3549,N_92,N_707);
and U3550 (N_3550,N_2317,N_1775);
nor U3551 (N_3551,N_1967,N_2382);
and U3552 (N_3552,N_2879,N_2839);
nor U3553 (N_3553,N_2795,N_1800);
nor U3554 (N_3554,N_2233,N_2125);
xor U3555 (N_3555,N_6,N_2242);
and U3556 (N_3556,N_1780,N_976);
and U3557 (N_3557,N_140,N_1228);
nor U3558 (N_3558,N_1783,N_2703);
nand U3559 (N_3559,N_1213,N_2844);
nand U3560 (N_3560,N_1712,N_698);
nand U3561 (N_3561,N_412,N_1976);
nor U3562 (N_3562,N_2441,N_186);
nand U3563 (N_3563,N_300,N_1941);
or U3564 (N_3564,N_1374,N_464);
and U3565 (N_3565,N_2184,N_854);
nand U3566 (N_3566,N_301,N_2170);
nor U3567 (N_3567,N_3112,N_1263);
or U3568 (N_3568,N_583,N_3036);
and U3569 (N_3569,N_280,N_1182);
or U3570 (N_3570,N_1817,N_1874);
xor U3571 (N_3571,N_1645,N_2285);
or U3572 (N_3572,N_1173,N_2340);
xnor U3573 (N_3573,N_793,N_1341);
and U3574 (N_3574,N_342,N_1125);
nand U3575 (N_3575,N_100,N_2926);
xor U3576 (N_3576,N_3082,N_2339);
and U3577 (N_3577,N_1401,N_1814);
nor U3578 (N_3578,N_2274,N_315);
and U3579 (N_3579,N_56,N_488);
xnor U3580 (N_3580,N_860,N_2872);
or U3581 (N_3581,N_1844,N_1720);
nor U3582 (N_3582,N_776,N_689);
and U3583 (N_3583,N_729,N_161);
and U3584 (N_3584,N_3023,N_2204);
and U3585 (N_3585,N_2047,N_1519);
xor U3586 (N_3586,N_2220,N_2216);
and U3587 (N_3587,N_2602,N_2673);
nor U3588 (N_3588,N_2858,N_849);
and U3589 (N_3589,N_1439,N_2095);
and U3590 (N_3590,N_506,N_1352);
and U3591 (N_3591,N_2761,N_1697);
or U3592 (N_3592,N_1334,N_1473);
nor U3593 (N_3593,N_1098,N_3083);
and U3594 (N_3594,N_2546,N_2282);
and U3595 (N_3595,N_1061,N_2798);
xnor U3596 (N_3596,N_1893,N_979);
nor U3597 (N_3597,N_426,N_2416);
and U3598 (N_3598,N_2574,N_2415);
nor U3599 (N_3599,N_886,N_2422);
xnor U3600 (N_3600,N_1069,N_493);
or U3601 (N_3601,N_7,N_2308);
nor U3602 (N_3602,N_611,N_2729);
nor U3603 (N_3603,N_1547,N_146);
nor U3604 (N_3604,N_2255,N_3020);
and U3605 (N_3605,N_1588,N_2941);
nor U3606 (N_3606,N_2161,N_3072);
and U3607 (N_3607,N_1467,N_1294);
xor U3608 (N_3608,N_920,N_294);
nor U3609 (N_3609,N_1895,N_2990);
or U3610 (N_3610,N_3069,N_106);
and U3611 (N_3611,N_2857,N_884);
xnor U3612 (N_3612,N_1492,N_2832);
and U3613 (N_3613,N_2254,N_299);
nand U3614 (N_3614,N_913,N_349);
nor U3615 (N_3615,N_47,N_2217);
or U3616 (N_3616,N_2150,N_2486);
xnor U3617 (N_3617,N_1445,N_678);
or U3618 (N_3618,N_1432,N_1020);
nand U3619 (N_3619,N_2945,N_2566);
nand U3620 (N_3620,N_2190,N_2591);
nand U3621 (N_3621,N_612,N_2262);
nand U3622 (N_3622,N_1854,N_2094);
and U3623 (N_3623,N_1106,N_247);
and U3624 (N_3624,N_2718,N_2630);
nand U3625 (N_3625,N_2651,N_1320);
xnor U3626 (N_3626,N_482,N_2688);
or U3627 (N_3627,N_2504,N_545);
nand U3628 (N_3628,N_1446,N_1797);
nand U3629 (N_3629,N_2831,N_2172);
nor U3630 (N_3630,N_2408,N_2970);
and U3631 (N_3631,N_774,N_3094);
or U3632 (N_3632,N_872,N_2544);
or U3633 (N_3633,N_484,N_2749);
and U3634 (N_3634,N_1119,N_518);
and U3635 (N_3635,N_2221,N_1958);
nor U3636 (N_3636,N_1338,N_1693);
xnor U3637 (N_3637,N_2559,N_2612);
xor U3638 (N_3638,N_1755,N_2175);
or U3639 (N_3639,N_1239,N_2556);
and U3640 (N_3640,N_1096,N_608);
nor U3641 (N_3641,N_2022,N_472);
or U3642 (N_3642,N_2144,N_1727);
and U3643 (N_3643,N_1006,N_2692);
nand U3644 (N_3644,N_1037,N_2768);
nand U3645 (N_3645,N_1134,N_2341);
or U3646 (N_3646,N_753,N_675);
xnor U3647 (N_3647,N_2122,N_399);
or U3648 (N_3648,N_3106,N_850);
xor U3649 (N_3649,N_940,N_1128);
xor U3650 (N_3650,N_941,N_844);
nor U3651 (N_3651,N_2097,N_2487);
or U3652 (N_3652,N_2611,N_971);
xnor U3653 (N_3653,N_1909,N_1927);
nand U3654 (N_3654,N_2828,N_1008);
and U3655 (N_3655,N_416,N_527);
nand U3656 (N_3656,N_2609,N_1573);
xnor U3657 (N_3657,N_1548,N_2634);
and U3658 (N_3658,N_3043,N_1116);
and U3659 (N_3659,N_520,N_2506);
and U3660 (N_3660,N_1920,N_67);
nor U3661 (N_3661,N_1741,N_962);
and U3662 (N_3662,N_1991,N_129);
nand U3663 (N_3663,N_1747,N_1507);
nand U3664 (N_3664,N_331,N_2245);
or U3665 (N_3665,N_2838,N_786);
nand U3666 (N_3666,N_1739,N_2733);
xnor U3667 (N_3667,N_2155,N_2361);
nor U3668 (N_3668,N_2648,N_2093);
xnor U3669 (N_3669,N_1371,N_1578);
and U3670 (N_3670,N_1258,N_1520);
and U3671 (N_3671,N_1138,N_2672);
nor U3672 (N_3672,N_576,N_784);
or U3673 (N_3673,N_119,N_2386);
and U3674 (N_3674,N_694,N_2080);
nor U3675 (N_3675,N_2649,N_109);
nand U3676 (N_3676,N_1975,N_1978);
or U3677 (N_3677,N_1209,N_584);
xor U3678 (N_3678,N_288,N_1296);
nand U3679 (N_3679,N_1725,N_2211);
xor U3680 (N_3680,N_2644,N_3055);
nor U3681 (N_3681,N_2482,N_2336);
and U3682 (N_3682,N_2882,N_53);
nor U3683 (N_3683,N_1429,N_49);
xnor U3684 (N_3684,N_2141,N_1585);
or U3685 (N_3685,N_2993,N_2290);
or U3686 (N_3686,N_154,N_2104);
nor U3687 (N_3687,N_2082,N_1813);
nor U3688 (N_3688,N_2542,N_1261);
or U3689 (N_3689,N_2054,N_528);
nor U3690 (N_3690,N_2697,N_2866);
xnor U3691 (N_3691,N_512,N_2049);
xnor U3692 (N_3692,N_2121,N_14);
xnor U3693 (N_3693,N_98,N_816);
and U3694 (N_3694,N_71,N_2410);
nand U3695 (N_3695,N_804,N_891);
xnor U3696 (N_3696,N_1454,N_641);
or U3697 (N_3697,N_3124,N_606);
or U3698 (N_3698,N_1898,N_573);
nor U3699 (N_3699,N_2006,N_2996);
xor U3700 (N_3700,N_815,N_975);
xnor U3701 (N_3701,N_1803,N_2440);
and U3702 (N_3702,N_2661,N_1373);
or U3703 (N_3703,N_543,N_359);
or U3704 (N_3704,N_756,N_1572);
xor U3705 (N_3705,N_3081,N_2902);
nor U3706 (N_3706,N_1133,N_485);
and U3707 (N_3707,N_2061,N_2028);
and U3708 (N_3708,N_476,N_26);
or U3709 (N_3709,N_2875,N_1554);
nand U3710 (N_3710,N_1664,N_1475);
nor U3711 (N_3711,N_2189,N_22);
and U3712 (N_3712,N_2771,N_952);
xnor U3713 (N_3713,N_2011,N_2199);
nand U3714 (N_3714,N_1531,N_800);
nand U3715 (N_3715,N_2776,N_1953);
nand U3716 (N_3716,N_799,N_1393);
xor U3717 (N_3717,N_2417,N_1254);
nand U3718 (N_3718,N_2507,N_2069);
xnor U3719 (N_3719,N_2903,N_2933);
nand U3720 (N_3720,N_1866,N_802);
and U3721 (N_3721,N_633,N_3013);
nor U3722 (N_3722,N_1771,N_141);
nand U3723 (N_3723,N_680,N_2914);
or U3724 (N_3724,N_2809,N_192);
nand U3725 (N_3725,N_798,N_254);
nor U3726 (N_3726,N_957,N_3097);
nand U3727 (N_3727,N_2526,N_1835);
and U3728 (N_3728,N_447,N_502);
nand U3729 (N_3729,N_3123,N_1306);
or U3730 (N_3730,N_2145,N_70);
and U3731 (N_3731,N_669,N_343);
nand U3732 (N_3732,N_1313,N_3017);
xor U3733 (N_3733,N_1200,N_1185);
nand U3734 (N_3734,N_2854,N_1396);
nand U3735 (N_3735,N_2085,N_2442);
nand U3736 (N_3736,N_1638,N_2454);
nand U3737 (N_3737,N_2014,N_1925);
or U3738 (N_3738,N_1427,N_1699);
xor U3739 (N_3739,N_2898,N_978);
xor U3740 (N_3740,N_706,N_1346);
nand U3741 (N_3741,N_2676,N_2432);
and U3742 (N_3742,N_318,N_2395);
nor U3743 (N_3743,N_2306,N_1137);
nor U3744 (N_3744,N_2081,N_1220);
or U3745 (N_3745,N_181,N_1449);
nand U3746 (N_3746,N_522,N_2418);
nor U3747 (N_3747,N_1270,N_2389);
nor U3748 (N_3748,N_764,N_618);
xor U3749 (N_3749,N_1451,N_1196);
nor U3750 (N_3750,N_1663,N_896);
nand U3751 (N_3751,N_1773,N_1097);
xnor U3752 (N_3752,N_2043,N_1702);
or U3753 (N_3753,N_1067,N_1342);
nor U3754 (N_3754,N_202,N_94);
nand U3755 (N_3755,N_988,N_1926);
or U3756 (N_3756,N_869,N_2741);
nand U3757 (N_3757,N_1627,N_1659);
nand U3758 (N_3758,N_2191,N_898);
nor U3759 (N_3759,N_2458,N_640);
nor U3760 (N_3760,N_1307,N_1324);
nor U3761 (N_3761,N_1807,N_2353);
and U3762 (N_3762,N_2813,N_572);
nand U3763 (N_3763,N_1190,N_1630);
or U3764 (N_3764,N_1628,N_2600);
or U3765 (N_3765,N_313,N_2088);
or U3766 (N_3766,N_2338,N_888);
xor U3767 (N_3767,N_2020,N_851);
and U3768 (N_3768,N_356,N_2376);
nand U3769 (N_3769,N_1253,N_2671);
xnor U3770 (N_3770,N_1244,N_1416);
xor U3771 (N_3771,N_2637,N_1606);
nor U3772 (N_3772,N_748,N_1465);
xnor U3773 (N_3773,N_1879,N_1621);
nor U3774 (N_3774,N_2987,N_2932);
nand U3775 (N_3775,N_1330,N_1274);
and U3776 (N_3776,N_1136,N_1508);
nor U3777 (N_3777,N_3056,N_2485);
nor U3778 (N_3778,N_2725,N_1045);
nor U3779 (N_3779,N_629,N_1509);
and U3780 (N_3780,N_500,N_2120);
nand U3781 (N_3781,N_171,N_2759);
or U3782 (N_3782,N_916,N_2307);
xor U3783 (N_3783,N_162,N_3024);
nand U3784 (N_3784,N_2237,N_2208);
xnor U3785 (N_3785,N_1897,N_131);
xor U3786 (N_3786,N_2739,N_1683);
and U3787 (N_3787,N_569,N_1985);
nor U3788 (N_3788,N_1877,N_1912);
nor U3789 (N_3789,N_1538,N_1735);
nand U3790 (N_3790,N_2078,N_759);
xor U3791 (N_3791,N_492,N_1505);
or U3792 (N_3792,N_285,N_1156);
nor U3793 (N_3793,N_710,N_2533);
and U3794 (N_3794,N_855,N_2657);
nor U3795 (N_3795,N_468,N_392);
nand U3796 (N_3796,N_366,N_214);
nand U3797 (N_3797,N_1632,N_907);
nand U3798 (N_3798,N_2201,N_1293);
xnor U3799 (N_3799,N_1929,N_2829);
and U3800 (N_3800,N_1121,N_2116);
or U3801 (N_3801,N_965,N_1262);
and U3802 (N_3802,N_2954,N_147);
nor U3803 (N_3803,N_1038,N_2629);
or U3804 (N_3804,N_248,N_541);
and U3805 (N_3805,N_213,N_1234);
xnor U3806 (N_3806,N_2250,N_2387);
nand U3807 (N_3807,N_2959,N_1381);
or U3808 (N_3808,N_390,N_2460);
xor U3809 (N_3809,N_715,N_746);
or U3810 (N_3810,N_3040,N_2706);
and U3811 (N_3811,N_1551,N_2541);
xnor U3812 (N_3812,N_2198,N_868);
and U3813 (N_3813,N_227,N_2754);
and U3814 (N_3814,N_2024,N_1333);
and U3815 (N_3815,N_2986,N_657);
or U3816 (N_3816,N_542,N_566);
or U3817 (N_3817,N_1999,N_1260);
nand U3818 (N_3818,N_2782,N_436);
xnor U3819 (N_3819,N_835,N_1728);
or U3820 (N_3820,N_1319,N_2048);
xor U3821 (N_3821,N_391,N_2246);
or U3822 (N_3822,N_1027,N_733);
xor U3823 (N_3823,N_1850,N_1948);
and U3824 (N_3824,N_2620,N_911);
and U3825 (N_3825,N_955,N_1610);
xnor U3826 (N_3826,N_1695,N_2596);
xor U3827 (N_3827,N_483,N_2484);
and U3828 (N_3828,N_2103,N_1717);
or U3829 (N_3829,N_1705,N_2196);
xnor U3830 (N_3830,N_3062,N_1708);
or U3831 (N_3831,N_567,N_2616);
xnor U3832 (N_3832,N_3110,N_3005);
or U3833 (N_3833,N_1523,N_2187);
nor U3834 (N_3834,N_2169,N_2786);
or U3835 (N_3835,N_378,N_2098);
nand U3836 (N_3836,N_2820,N_439);
and U3837 (N_3837,N_1471,N_2086);
nand U3838 (N_3838,N_2163,N_2529);
xor U3839 (N_3839,N_2641,N_708);
nand U3840 (N_3840,N_127,N_203);
nand U3841 (N_3841,N_1271,N_2142);
or U3842 (N_3842,N_1923,N_2391);
xnor U3843 (N_3843,N_1298,N_2716);
xnor U3844 (N_3844,N_2397,N_2071);
nand U3845 (N_3845,N_15,N_2429);
or U3846 (N_3846,N_2769,N_1896);
nor U3847 (N_3847,N_1880,N_2859);
or U3848 (N_3848,N_1256,N_2239);
or U3849 (N_3849,N_2156,N_2378);
nand U3850 (N_3850,N_1646,N_2751);
xor U3851 (N_3851,N_2747,N_132);
nand U3852 (N_3852,N_396,N_319);
xor U3853 (N_3853,N_1726,N_1649);
xnor U3854 (N_3854,N_2390,N_1660);
xnor U3855 (N_3855,N_658,N_2722);
nor U3856 (N_3856,N_1181,N_1636);
xor U3857 (N_3857,N_1933,N_1386);
and U3858 (N_3858,N_1460,N_2500);
xor U3859 (N_3859,N_2251,N_2865);
nor U3860 (N_3860,N_2218,N_275);
nand U3861 (N_3861,N_32,N_1083);
xnor U3862 (N_3862,N_2252,N_2398);
nand U3863 (N_3863,N_1364,N_692);
nor U3864 (N_3864,N_2877,N_1553);
xor U3865 (N_3865,N_758,N_1321);
nor U3866 (N_3866,N_2453,N_421);
xor U3867 (N_3867,N_1227,N_2522);
nor U3868 (N_3868,N_1286,N_5);
or U3869 (N_3869,N_2880,N_3058);
or U3870 (N_3870,N_550,N_474);
and U3871 (N_3871,N_128,N_1640);
nand U3872 (N_3872,N_2462,N_2801);
nor U3873 (N_3873,N_1641,N_1480);
xor U3874 (N_3874,N_1289,N_1217);
xor U3875 (N_3875,N_2852,N_3068);
and U3876 (N_3876,N_1973,N_160);
or U3877 (N_3877,N_783,N_2797);
and U3878 (N_3878,N_1349,N_1616);
and U3879 (N_3879,N_1107,N_2193);
nor U3880 (N_3880,N_516,N_1157);
nand U3881 (N_3881,N_2322,N_2087);
nand U3882 (N_3882,N_1146,N_24);
nor U3883 (N_3883,N_3114,N_284);
xor U3884 (N_3884,N_2646,N_912);
nor U3885 (N_3885,N_1801,N_825);
and U3886 (N_3886,N_1090,N_1193);
or U3887 (N_3887,N_2756,N_330);
or U3888 (N_3888,N_2543,N_654);
nand U3889 (N_3889,N_2868,N_1989);
and U3890 (N_3890,N_407,N_856);
or U3891 (N_3891,N_2778,N_1718);
nand U3892 (N_3892,N_2149,N_1670);
or U3893 (N_3893,N_1820,N_2437);
nand U3894 (N_3894,N_2784,N_3115);
nand U3895 (N_3895,N_2633,N_2978);
and U3896 (N_3896,N_1474,N_2148);
and U3897 (N_3897,N_2588,N_2911);
nand U3898 (N_3898,N_810,N_901);
nor U3899 (N_3899,N_762,N_3047);
nand U3900 (N_3900,N_372,N_1626);
nand U3901 (N_3901,N_1785,N_1594);
nand U3902 (N_3902,N_614,N_2752);
nor U3903 (N_3903,N_1919,N_2579);
nand U3904 (N_3904,N_273,N_134);
xnor U3905 (N_3905,N_2958,N_627);
xor U3906 (N_3906,N_351,N_2909);
nor U3907 (N_3907,N_1101,N_339);
or U3908 (N_3908,N_1435,N_268);
or U3909 (N_3909,N_260,N_517);
nor U3910 (N_3910,N_2878,N_1028);
xor U3911 (N_3911,N_3042,N_2842);
and U3912 (N_3912,N_2232,N_841);
nand U3913 (N_3913,N_2793,N_2907);
xor U3914 (N_3914,N_1040,N_2923);
nor U3915 (N_3915,N_2908,N_3016);
xnor U3916 (N_3916,N_2489,N_501);
nand U3917 (N_3917,N_43,N_1715);
xor U3918 (N_3918,N_2734,N_28);
and U3919 (N_3919,N_736,N_647);
and U3920 (N_3920,N_1198,N_1764);
and U3921 (N_3921,N_2153,N_478);
or U3922 (N_3922,N_685,N_266);
nand U3923 (N_3923,N_2684,N_1438);
xor U3924 (N_3924,N_833,N_2658);
nor U3925 (N_3925,N_469,N_2041);
or U3926 (N_3926,N_2058,N_2553);
nand U3927 (N_3927,N_437,N_1963);
or U3928 (N_3928,N_2421,N_910);
or U3929 (N_3929,N_1332,N_1344);
xnor U3930 (N_3930,N_2302,N_878);
xor U3931 (N_3931,N_2874,N_1208);
xor U3932 (N_3932,N_2508,N_852);
xor U3933 (N_3933,N_1603,N_1382);
xor U3934 (N_3934,N_2892,N_3095);
nand U3935 (N_3935,N_1788,N_1410);
and U3936 (N_3936,N_1385,N_683);
nand U3937 (N_3937,N_2779,N_95);
and U3938 (N_3938,N_108,N_1019);
and U3939 (N_3939,N_2619,N_1108);
nand U3940 (N_3940,N_674,N_311);
xnor U3941 (N_3941,N_3053,N_845);
or U3942 (N_3942,N_2726,N_847);
nor U3943 (N_3943,N_2512,N_2918);
and U3944 (N_3944,N_903,N_2457);
nor U3945 (N_3945,N_1472,N_781);
or U3946 (N_3946,N_982,N_2275);
or U3947 (N_3947,N_1297,N_166);
and U3948 (N_3948,N_408,N_2117);
or U3949 (N_3949,N_123,N_1535);
nor U3950 (N_3950,N_1232,N_536);
or U3951 (N_3951,N_3105,N_2850);
or U3952 (N_3952,N_1738,N_2736);
xnor U3953 (N_3953,N_2412,N_2663);
nand U3954 (N_3954,N_2763,N_1317);
nor U3955 (N_3955,N_1637,N_663);
xor U3956 (N_3956,N_3107,N_1225);
nand U3957 (N_3957,N_1462,N_2585);
xor U3958 (N_3958,N_295,N_2912);
nand U3959 (N_3959,N_2682,N_1223);
xor U3960 (N_3960,N_1611,N_2379);
nand U3961 (N_3961,N_393,N_1951);
nor U3962 (N_3962,N_2964,N_2608);
nand U3963 (N_3963,N_918,N_1682);
nand U3964 (N_3964,N_2922,N_625);
nand U3965 (N_3965,N_596,N_1025);
xor U3966 (N_3966,N_2975,N_2551);
or U3967 (N_3967,N_1949,N_430);
nand U3968 (N_3968,N_823,N_1299);
nor U3969 (N_3969,N_795,N_2704);
and U3970 (N_3970,N_2856,N_362);
nand U3971 (N_3971,N_2540,N_1353);
or U3972 (N_3972,N_1765,N_2705);
and U3973 (N_3973,N_2345,N_2781);
or U3974 (N_3974,N_388,N_2084);
or U3975 (N_3975,N_837,N_3000);
nand U3976 (N_3976,N_737,N_1405);
and U3977 (N_3977,N_1122,N_1115);
nor U3978 (N_3978,N_54,N_1243);
xnor U3979 (N_3979,N_1590,N_2219);
xnor U3980 (N_3980,N_2561,N_2573);
and U3981 (N_3981,N_174,N_1631);
or U3982 (N_3982,N_2293,N_1890);
or U3983 (N_3983,N_1577,N_1452);
and U3984 (N_3984,N_1679,N_48);
nor U3985 (N_3985,N_2430,N_2762);
xor U3986 (N_3986,N_2514,N_1153);
and U3987 (N_3987,N_237,N_322);
or U3988 (N_3988,N_494,N_2770);
nor U3989 (N_3989,N_471,N_1618);
and U3990 (N_3990,N_2717,N_2425);
nand U3991 (N_3991,N_1589,N_2281);
or U3992 (N_3992,N_1395,N_686);
and U3993 (N_3993,N_693,N_499);
nor U3994 (N_3994,N_2904,N_2288);
xor U3995 (N_3995,N_1398,N_548);
or U3996 (N_3996,N_1811,N_1124);
xor U3997 (N_3997,N_68,N_440);
nor U3998 (N_3998,N_785,N_1552);
nand U3999 (N_3999,N_1394,N_2435);
xnor U4000 (N_4000,N_1885,N_1206);
nand U4001 (N_4001,N_438,N_2294);
nand U4002 (N_4002,N_2948,N_2326);
nor U4003 (N_4003,N_754,N_1930);
nand U4004 (N_4004,N_3057,N_2300);
nor U4005 (N_4005,N_2167,N_1165);
and U4006 (N_4006,N_2668,N_2310);
nand U4007 (N_4007,N_919,N_1326);
nand U4008 (N_4008,N_210,N_586);
xor U4009 (N_4009,N_3038,N_2271);
or U4010 (N_4010,N_2571,N_354);
nand U4011 (N_4011,N_1805,N_1249);
xnor U4012 (N_4012,N_555,N_2333);
and U4013 (N_4013,N_836,N_2814);
and U4014 (N_4014,N_1758,N_769);
nand U4015 (N_4015,N_251,N_2985);
and U4016 (N_4016,N_2509,N_523);
and U4017 (N_4017,N_60,N_2091);
and U4018 (N_4018,N_1248,N_1591);
and U4019 (N_4019,N_914,N_2601);
nand U4020 (N_4020,N_3096,N_1971);
or U4021 (N_4021,N_344,N_1900);
and U4022 (N_4022,N_1478,N_180);
or U4023 (N_4023,N_1824,N_1688);
or U4024 (N_4024,N_2685,N_1954);
or U4025 (N_4025,N_1846,N_2849);
xor U4026 (N_4026,N_921,N_2650);
or U4027 (N_4027,N_1743,N_20);
nand U4028 (N_4028,N_2511,N_373);
xnor U4029 (N_4029,N_1776,N_651);
xor U4030 (N_4030,N_2973,N_1105);
xnor U4031 (N_4031,N_1940,N_1960);
or U4032 (N_4032,N_2448,N_456);
nand U4033 (N_4033,N_602,N_635);
nand U4034 (N_4034,N_1311,N_642);
nor U4035 (N_4035,N_1359,N_1233);
nand U4036 (N_4036,N_2775,N_859);
nor U4037 (N_4037,N_2352,N_814);
nor U4038 (N_4038,N_2016,N_2209);
xnor U4039 (N_4039,N_2044,N_1080);
or U4040 (N_4040,N_385,N_2894);
nand U4041 (N_4041,N_2249,N_1887);
xnor U4042 (N_4042,N_2334,N_383);
nor U4043 (N_4043,N_765,N_2399);
nand U4044 (N_4044,N_110,N_2977);
and U4045 (N_4045,N_37,N_1109);
nor U4046 (N_4046,N_2004,N_909);
xor U4047 (N_4047,N_3032,N_1964);
nor U4048 (N_4048,N_2027,N_681);
xnor U4049 (N_4049,N_1369,N_1215);
nor U4050 (N_4050,N_1370,N_2256);
xnor U4051 (N_4051,N_2549,N_1348);
nand U4052 (N_4052,N_2934,N_2742);
nand U4053 (N_4053,N_877,N_2228);
nand U4054 (N_4054,N_405,N_2244);
and U4055 (N_4055,N_3022,N_574);
xnor U4056 (N_4056,N_2983,N_1763);
and U4057 (N_4057,N_2881,N_935);
or U4058 (N_4058,N_2400,N_2743);
xor U4059 (N_4059,N_2108,N_1250);
xor U4060 (N_4060,N_1499,N_1746);
nand U4061 (N_4061,N_117,N_244);
xnor U4062 (N_4062,N_2342,N_458);
or U4063 (N_4063,N_370,N_598);
nand U4064 (N_4064,N_2530,N_568);
nor U4065 (N_4065,N_1093,N_1267);
xor U4066 (N_4066,N_906,N_1527);
nand U4067 (N_4067,N_1068,N_1826);
xnor U4068 (N_4068,N_2517,N_1639);
xor U4069 (N_4069,N_2002,N_2765);
and U4070 (N_4070,N_269,N_1529);
nor U4071 (N_4071,N_1777,N_2134);
and U4072 (N_4072,N_1425,N_554);
or U4073 (N_4073,N_990,N_256);
nand U4074 (N_4074,N_2607,N_231);
nand U4075 (N_4075,N_2581,N_2401);
xor U4076 (N_4076,N_730,N_1113);
nor U4077 (N_4077,N_2459,N_1111);
nand U4078 (N_4078,N_2873,N_882);
nand U4079 (N_4079,N_552,N_579);
nand U4080 (N_4080,N_2179,N_267);
nor U4081 (N_4081,N_3077,N_1862);
nor U4082 (N_4082,N_2577,N_1189);
xor U4083 (N_4083,N_2367,N_2750);
or U4084 (N_4084,N_2023,N_1091);
xor U4085 (N_4085,N_2966,N_324);
and U4086 (N_4086,N_1605,N_2597);
xor U4087 (N_4087,N_2516,N_2241);
xnor U4088 (N_4088,N_1424,N_1716);
nand U4089 (N_4089,N_1540,N_2266);
xor U4090 (N_4090,N_3004,N_126);
or U4091 (N_4091,N_2292,N_274);
xor U4092 (N_4092,N_2471,N_2072);
or U4093 (N_4093,N_133,N_863);
nor U4094 (N_4094,N_135,N_286);
xor U4095 (N_4095,N_503,N_1691);
nor U4096 (N_4096,N_1470,N_1863);
nor U4097 (N_4097,N_1565,N_546);
xor U4098 (N_4098,N_387,N_3061);
xor U4099 (N_4099,N_89,N_84);
xnor U4100 (N_4100,N_2864,N_1744);
or U4101 (N_4101,N_1304,N_2643);
nand U4102 (N_4102,N_2029,N_2654);
nand U4103 (N_4103,N_246,N_69);
nand U4104 (N_4104,N_61,N_3001);
nor U4105 (N_4105,N_1592,N_1295);
nor U4106 (N_4106,N_1833,N_1789);
nand U4107 (N_4107,N_525,N_2886);
nand U4108 (N_4108,N_610,N_1761);
nor U4109 (N_4109,N_2248,N_198);
or U4110 (N_4110,N_1674,N_788);
nand U4111 (N_4111,N_2015,N_1517);
nor U4112 (N_4112,N_623,N_1852);
xor U4113 (N_4113,N_2683,N_2901);
nor U4114 (N_4114,N_3120,N_2497);
or U4115 (N_4115,N_1680,N_498);
nor U4116 (N_4116,N_632,N_448);
or U4117 (N_4117,N_2930,N_2123);
nand U4118 (N_4118,N_2693,N_1706);
and U4119 (N_4119,N_2466,N_271);
nor U4120 (N_4120,N_2678,N_1567);
and U4121 (N_4121,N_2291,N_1323);
or U4122 (N_4122,N_2702,N_1079);
and U4123 (N_4123,N_1569,N_751);
or U4124 (N_4124,N_761,N_413);
xor U4125 (N_4125,N_2467,N_461);
or U4126 (N_4126,N_1222,N_2994);
nand U4127 (N_4127,N_191,N_2481);
xor U4128 (N_4128,N_196,N_644);
xnor U4129 (N_4129,N_2835,N_1966);
or U4130 (N_4130,N_996,N_2615);
nand U4131 (N_4131,N_2413,N_1671);
xor U4132 (N_4132,N_983,N_1155);
nand U4133 (N_4133,N_1806,N_1158);
nor U4134 (N_4134,N_143,N_1345);
nand U4135 (N_4135,N_182,N_2005);
xor U4136 (N_4136,N_2677,N_2025);
nor U4137 (N_4137,N_2989,N_2177);
nor U4138 (N_4138,N_395,N_2446);
nand U4139 (N_4139,N_1404,N_241);
nand U4140 (N_4140,N_336,N_701);
nor U4141 (N_4141,N_2181,N_2264);
and U4142 (N_4142,N_1360,N_2119);
and U4143 (N_4143,N_2396,N_636);
xor U4144 (N_4144,N_3118,N_993);
or U4145 (N_4145,N_2443,N_1997);
or U4146 (N_4146,N_1821,N_1252);
xor U4147 (N_4147,N_1312,N_989);
nand U4148 (N_4148,N_462,N_380);
nand U4149 (N_4149,N_74,N_1021);
nand U4150 (N_4150,N_653,N_477);
and U4151 (N_4151,N_2315,N_2343);
nor U4152 (N_4152,N_361,N_2287);
xor U4153 (N_4153,N_511,N_2280);
nor U4154 (N_4154,N_1392,N_1147);
xnor U4155 (N_4155,N_445,N_3122);
or U4156 (N_4156,N_77,N_2712);
nand U4157 (N_4157,N_2707,N_2197);
and U4158 (N_4158,N_646,N_2194);
nor U4159 (N_4159,N_1132,N_2789);
or U4160 (N_4160,N_2943,N_75);
nor U4161 (N_4161,N_2439,N_360);
or U4162 (N_4162,N_1871,N_580);
or U4163 (N_4163,N_1221,N_52);
nand U4164 (N_4164,N_1889,N_1770);
xor U4165 (N_4165,N_1103,N_2982);
and U4166 (N_4166,N_1604,N_2491);
nand U4167 (N_4167,N_1003,N_593);
xnor U4168 (N_4168,N_2159,N_839);
or U4169 (N_4169,N_257,N_535);
and U4170 (N_4170,N_1910,N_433);
xor U4171 (N_4171,N_194,N_1563);
nand U4172 (N_4172,N_887,N_1959);
nand U4173 (N_4173,N_900,N_1942);
nor U4174 (N_4174,N_1600,N_964);
xnor U4175 (N_4175,N_2708,N_88);
or U4176 (N_4176,N_2346,N_2152);
or U4177 (N_4177,N_1661,N_1917);
nor U4178 (N_4178,N_1063,N_1187);
xnor U4179 (N_4179,N_671,N_1219);
nor U4180 (N_4180,N_1060,N_1943);
xor U4181 (N_4181,N_2748,N_276);
and U4182 (N_4182,N_1337,N_259);
xor U4183 (N_4183,N_1908,N_1994);
and U4184 (N_4184,N_1878,N_3102);
xor U4185 (N_4185,N_78,N_1388);
nand U4186 (N_4186,N_717,N_1011);
nand U4187 (N_4187,N_538,N_1798);
nor U4188 (N_4188,N_2402,N_2621);
and U4189 (N_4189,N_1464,N_561);
nor U4190 (N_4190,N_2578,N_193);
or U4191 (N_4191,N_1996,N_1453);
xnor U4192 (N_4192,N_3079,N_2320);
and U4193 (N_4193,N_81,N_893);
and U4194 (N_4194,N_25,N_1174);
nand U4195 (N_4195,N_1292,N_419);
or U4196 (N_4196,N_2273,N_995);
and U4197 (N_4197,N_29,N_1140);
or U4198 (N_4198,N_2656,N_2885);
and U4199 (N_4199,N_444,N_1873);
nor U4200 (N_4200,N_643,N_73);
xor U4201 (N_4201,N_1175,N_2001);
xnor U4202 (N_4202,N_766,N_287);
nor U4203 (N_4203,N_2812,N_2171);
or U4204 (N_4204,N_2423,N_777);
and U4205 (N_4205,N_1904,N_2286);
nor U4206 (N_4206,N_121,N_102);
and U4207 (N_4207,N_951,N_184);
xnor U4208 (N_4208,N_665,N_1170);
and U4209 (N_4209,N_2476,N_2344);
nand U4210 (N_4210,N_2337,N_389);
nand U4211 (N_4211,N_577,N_2362);
xnor U4212 (N_4212,N_2622,N_2017);
nand U4213 (N_4213,N_1376,N_401);
or U4214 (N_4214,N_705,N_1987);
xor U4215 (N_4215,N_1126,N_1469);
nor U4216 (N_4216,N_1309,N_922);
nand U4217 (N_4217,N_2213,N_1300);
and U4218 (N_4218,N_185,N_169);
and U4219 (N_4219,N_2243,N_116);
or U4220 (N_4220,N_1365,N_222);
or U4221 (N_4221,N_1804,N_2174);
and U4222 (N_4222,N_897,N_2377);
or U4223 (N_4223,N_2420,N_1356);
or U4224 (N_4224,N_44,N_2363);
nand U4225 (N_4225,N_1318,N_526);
nand U4226 (N_4226,N_936,N_1409);
or U4227 (N_4227,N_1403,N_353);
or U4228 (N_4228,N_2815,N_1459);
nor U4229 (N_4229,N_1504,N_954);
nor U4230 (N_4230,N_923,N_1071);
nand U4231 (N_4231,N_2238,N_1272);
or U4232 (N_4232,N_3063,N_1139);
nand U4233 (N_4233,N_245,N_1442);
nand U4234 (N_4234,N_589,N_803);
nand U4235 (N_4235,N_3087,N_966);
xor U4236 (N_4236,N_1420,N_279);
nor U4237 (N_4237,N_1922,N_1434);
nor U4238 (N_4238,N_1891,N_505);
and U4239 (N_4239,N_2691,N_427);
nand U4240 (N_4240,N_1033,N_309);
or U4241 (N_4241,N_719,N_1468);
nor U4242 (N_4242,N_875,N_2479);
nor U4243 (N_4243,N_3078,N_76);
xor U4244 (N_4244,N_2335,N_3119);
xnor U4245 (N_4245,N_1902,N_2639);
nand U4246 (N_4246,N_3012,N_1482);
nand U4247 (N_4247,N_308,N_402);
nand U4248 (N_4248,N_377,N_2834);
or U4249 (N_4249,N_2105,N_1436);
nor U4250 (N_4250,N_262,N_1400);
nand U4251 (N_4251,N_659,N_985);
nor U4252 (N_4252,N_873,N_2374);
nand U4253 (N_4253,N_1819,N_834);
nand U4254 (N_4254,N_335,N_2804);
or U4255 (N_4255,N_1620,N_630);
xor U4256 (N_4256,N_1988,N_794);
and U4257 (N_4257,N_822,N_1130);
or U4258 (N_4258,N_1882,N_925);
nand U4259 (N_4259,N_3060,N_432);
nor U4260 (N_4260,N_2827,N_620);
nand U4261 (N_4261,N_2980,N_357);
xor U4262 (N_4262,N_1102,N_1654);
xnor U4263 (N_4263,N_235,N_1281);
or U4264 (N_4264,N_1257,N_278);
nand U4265 (N_4265,N_1479,N_1937);
xnor U4266 (N_4266,N_480,N_219);
or U4267 (N_4267,N_2942,N_881);
and U4268 (N_4268,N_1301,N_1932);
and U4269 (N_4269,N_403,N_792);
and U4270 (N_4270,N_1084,N_829);
nand U4271 (N_4271,N_457,N_1730);
nand U4272 (N_4272,N_486,N_778);
nor U4273 (N_4273,N_1643,N_2505);
nor U4274 (N_4274,N_2099,N_2567);
xnor U4275 (N_4275,N_1487,N_240);
xor U4276 (N_4276,N_2638,N_917);
xnor U4277 (N_4277,N_2518,N_329);
xor U4278 (N_4278,N_2940,N_2700);
or U4279 (N_4279,N_2464,N_664);
nand U4280 (N_4280,N_973,N_1192);
nand U4281 (N_4281,N_2424,N_296);
or U4282 (N_4282,N_112,N_59);
or U4283 (N_4283,N_16,N_1287);
xor U4284 (N_4284,N_382,N_375);
nand U4285 (N_4285,N_3049,N_732);
nor U4286 (N_4286,N_1018,N_1986);
nand U4287 (N_4287,N_1970,N_1859);
and U4288 (N_4288,N_1308,N_1983);
or U4289 (N_4289,N_556,N_1957);
nand U4290 (N_4290,N_2297,N_672);
and U4291 (N_4291,N_2008,N_2513);
nor U4292 (N_4292,N_2359,N_2956);
xor U4293 (N_4293,N_890,N_398);
nor U4294 (N_4294,N_1576,N_3090);
xnor U4295 (N_4295,N_2614,N_739);
xnor U4296 (N_4296,N_2721,N_1673);
xnor U4297 (N_4297,N_2520,N_1284);
and U4298 (N_4298,N_2394,N_1581);
and U4299 (N_4299,N_101,N_2594);
nand U4300 (N_4300,N_229,N_2917);
nand U4301 (N_4301,N_2670,N_3099);
nand U4302 (N_4302,N_1277,N_2205);
nand U4303 (N_4303,N_470,N_2066);
nand U4304 (N_4304,N_1906,N_2824);
nor U4305 (N_4305,N_1476,N_2477);
and U4306 (N_4306,N_2304,N_1916);
nand U4307 (N_4307,N_801,N_950);
xor U4308 (N_4308,N_3034,N_325);
or U4309 (N_4309,N_1058,N_2610);
nor U4310 (N_4310,N_948,N_2498);
or U4311 (N_4311,N_2463,N_934);
nand U4312 (N_4312,N_258,N_347);
or U4313 (N_4313,N_1733,N_963);
or U4314 (N_4314,N_1881,N_1754);
and U4315 (N_4315,N_2277,N_297);
nor U4316 (N_4316,N_1412,N_2380);
xor U4317 (N_4317,N_1245,N_1);
xnor U4318 (N_4318,N_2805,N_892);
nand U4319 (N_4319,N_2519,N_2931);
or U4320 (N_4320,N_609,N_704);
xor U4321 (N_4321,N_2060,N_2059);
xnor U4322 (N_4322,N_2624,N_1315);
and U4323 (N_4323,N_2628,N_1830);
xnor U4324 (N_4324,N_2483,N_2102);
xnor U4325 (N_4325,N_83,N_243);
and U4326 (N_4326,N_2449,N_969);
and U4327 (N_4327,N_1161,N_1698);
nor U4328 (N_4328,N_507,N_1748);
and U4329 (N_4329,N_591,N_768);
and U4330 (N_4330,N_1456,N_157);
nand U4331 (N_4331,N_397,N_2679);
xor U4332 (N_4332,N_2316,N_455);
or U4333 (N_4333,N_2817,N_1829);
xor U4334 (N_4334,N_2936,N_2910);
or U4335 (N_4335,N_270,N_1711);
xnor U4336 (N_4336,N_1749,N_2803);
or U4337 (N_4337,N_2140,N_1722);
or U4338 (N_4338,N_2488,N_2735);
xor U4339 (N_4339,N_712,N_1049);
nand U4340 (N_4340,N_2960,N_1858);
nand U4341 (N_4341,N_1448,N_2298);
xor U4342 (N_4342,N_2906,N_1050);
or U4343 (N_4343,N_33,N_1586);
nand U4344 (N_4344,N_592,N_1546);
nor U4345 (N_4345,N_1099,N_1466);
and U4346 (N_4346,N_2855,N_1601);
xor U4347 (N_4347,N_304,N_3010);
or U4348 (N_4348,N_2327,N_415);
and U4349 (N_4349,N_9,N_1127);
xnor U4350 (N_4350,N_2451,N_587);
nor U4351 (N_4351,N_443,N_650);
and U4352 (N_4352,N_883,N_2314);
nand U4353 (N_4353,N_2328,N_1463);
nor U4354 (N_4354,N_2576,N_64);
or U4355 (N_4355,N_2265,N_2070);
nand U4356 (N_4356,N_2699,N_1870);
nor U4357 (N_4357,N_1247,N_1570);
nand U4358 (N_4358,N_211,N_1613);
or U4359 (N_4359,N_2580,N_2461);
and U4360 (N_4360,N_1847,N_38);
xor U4361 (N_4361,N_2840,N_1843);
nand U4362 (N_4362,N_1159,N_1684);
or U4363 (N_4363,N_2564,N_2758);
or U4364 (N_4364,N_305,N_178);
and U4365 (N_4365,N_1046,N_3006);
or U4366 (N_4366,N_406,N_1672);
or U4367 (N_4367,N_1599,N_779);
or U4368 (N_4368,N_700,N_2039);
and U4369 (N_4369,N_575,N_1822);
nor U4370 (N_4370,N_2728,N_23);
nor U4371 (N_4371,N_2,N_1418);
and U4372 (N_4372,N_2929,N_1516);
and U4373 (N_4373,N_2092,N_3074);
xor U4374 (N_4374,N_2283,N_2495);
and U4375 (N_4375,N_562,N_2745);
and U4376 (N_4376,N_2063,N_239);
or U4377 (N_4377,N_1692,N_321);
nand U4378 (N_4378,N_994,N_1792);
xnor U4379 (N_4379,N_605,N_2860);
nor U4380 (N_4380,N_3014,N_2587);
nor U4381 (N_4381,N_1533,N_2295);
xnor U4382 (N_4382,N_615,N_2613);
nor U4383 (N_4383,N_2794,N_760);
and U4384 (N_4384,N_2999,N_807);
and U4385 (N_4385,N_1888,N_1689);
nand U4386 (N_4386,N_87,N_1756);
and U4387 (N_4387,N_420,N_1602);
nand U4388 (N_4388,N_1658,N_1853);
xnor U4389 (N_4389,N_949,N_720);
xnor U4390 (N_4390,N_2992,N_928);
and U4391 (N_4391,N_1013,N_939);
nor U4392 (N_4392,N_2653,N_1278);
or U4393 (N_4393,N_2869,N_1796);
nor U4394 (N_4394,N_961,N_998);
xnor U4395 (N_4395,N_422,N_2373);
nand U4396 (N_4396,N_8,N_165);
and U4397 (N_4397,N_2826,N_2118);
or U4398 (N_4398,N_1568,N_559);
xor U4399 (N_4399,N_4,N_2870);
nor U4400 (N_4400,N_490,N_452);
xor U4401 (N_4401,N_1310,N_2012);
and U4402 (N_4402,N_1142,N_167);
nor U4403 (N_4403,N_1721,N_2604);
xor U4404 (N_4404,N_2065,N_1053);
or U4405 (N_4405,N_1177,N_723);
xor U4406 (N_4406,N_2532,N_2186);
or U4407 (N_4407,N_1580,N_2224);
or U4408 (N_4408,N_2365,N_394);
xnor U4409 (N_4409,N_1934,N_1114);
xnor U4410 (N_4410,N_358,N_2963);
nor U4411 (N_4411,N_2035,N_2470);
nor U4412 (N_4412,N_2037,N_1851);
and U4413 (N_4413,N_770,N_1766);
or U4414 (N_4414,N_2539,N_1075);
nand U4415 (N_4415,N_41,N_1827);
xor U4416 (N_4416,N_1687,N_986);
and U4417 (N_4417,N_999,N_1740);
nor U4418 (N_4418,N_2101,N_1625);
nand U4419 (N_4419,N_1918,N_130);
nand U4420 (N_4420,N_2536,N_2057);
nor U4421 (N_4421,N_2261,N_2494);
or U4422 (N_4422,N_332,N_177);
xnor U4423 (N_4423,N_2200,N_1461);
nor U4424 (N_4424,N_673,N_690);
nor U4425 (N_4425,N_2819,N_1511);
xor U4426 (N_4426,N_824,N_201);
and U4427 (N_4427,N_1368,N_775);
xor U4428 (N_4428,N_65,N_449);
and U4429 (N_4429,N_697,N_1652);
nand U4430 (N_4430,N_970,N_929);
xnor U4431 (N_4431,N_1781,N_2388);
nand U4432 (N_4432,N_1541,N_1283);
and U4433 (N_4433,N_947,N_805);
nor U4434 (N_4434,N_1809,N_2129);
nor U4435 (N_4435,N_1759,N_2821);
xnor U4436 (N_4436,N_1363,N_944);
nor U4437 (N_4437,N_435,N_597);
nor U4438 (N_4438,N_1901,N_684);
xor U4439 (N_4439,N_379,N_1506);
nor U4440 (N_4440,N_2818,N_1044);
nor U4441 (N_4441,N_2472,N_1675);
and U4442 (N_4442,N_1831,N_2938);
nor U4443 (N_4443,N_2720,N_1012);
nor U4444 (N_4444,N_1945,N_163);
and U4445 (N_4445,N_314,N_2312);
or U4446 (N_4446,N_2531,N_2807);
or U4447 (N_4447,N_2296,N_2631);
xor U4448 (N_4448,N_699,N_190);
xor U4449 (N_4449,N_1437,N_1143);
nand U4450 (N_4450,N_1757,N_549);
xnor U4451 (N_4451,N_1328,N_1489);
nand U4452 (N_4452,N_1685,N_1246);
or U4453 (N_4453,N_2787,N_1160);
nand U4454 (N_4454,N_2766,N_2524);
nand U4455 (N_4455,N_1648,N_780);
nor U4456 (N_4456,N_876,N_1235);
or U4457 (N_4457,N_2154,N_871);
and U4458 (N_4458,N_638,N_1980);
xor U4459 (N_4459,N_410,N_622);
nand U4460 (N_4460,N_1681,N_1447);
xnor U4461 (N_4461,N_2525,N_2666);
xor U4462 (N_4462,N_255,N_2937);
and U4463 (N_4463,N_2861,N_2583);
and U4464 (N_4464,N_1201,N_540);
or U4465 (N_4465,N_2843,N_0);
xnor U4466 (N_4466,N_2605,N_409);
and U4467 (N_4467,N_2625,N_2409);
xor U4468 (N_4468,N_2040,N_1704);
xor U4469 (N_4469,N_600,N_1558);
nor U4470 (N_4470,N_104,N_649);
xnor U4471 (N_4471,N_1510,N_2077);
nand U4472 (N_4472,N_153,N_902);
nand U4473 (N_4473,N_578,N_1779);
and U4474 (N_4474,N_1070,N_2501);
nand U4475 (N_4475,N_404,N_2419);
nand U4476 (N_4476,N_1525,N_1860);
xor U4477 (N_4477,N_570,N_1839);
nor U4478 (N_4478,N_1946,N_1609);
nand U4479 (N_4479,N_721,N_172);
nand U4480 (N_4480,N_1709,N_62);
and U4481 (N_4481,N_1110,N_1555);
nand U4482 (N_4482,N_2019,N_35);
or U4483 (N_4483,N_539,N_1787);
xor U4484 (N_4484,N_1497,N_817);
or U4485 (N_4485,N_2944,N_2554);
or U4486 (N_4486,N_489,N_1524);
nand U4487 (N_4487,N_138,N_346);
or U4488 (N_4488,N_467,N_1782);
or U4489 (N_4489,N_2799,N_341);
or U4490 (N_4490,N_2289,N_942);
xnor U4491 (N_4491,N_2552,N_2806);
or U4492 (N_4492,N_1799,N_1135);
or U4493 (N_4493,N_711,N_1163);
and U4494 (N_4494,N_465,N_3);
or U4495 (N_4495,N_1419,N_218);
or U4496 (N_4496,N_2127,N_1440);
or U4497 (N_4497,N_1816,N_442);
nor U4498 (N_4498,N_1131,N_838);
nand U4499 (N_4499,N_261,N_1522);
and U4500 (N_4500,N_735,N_1428);
or U4501 (N_4501,N_1950,N_2823);
or U4502 (N_4502,N_2744,N_3109);
nand U4503 (N_4503,N_2231,N_2369);
nand U4504 (N_4504,N_2568,N_1302);
xor U4505 (N_4505,N_1268,N_220);
and U4506 (N_4506,N_2755,N_2740);
or U4507 (N_4507,N_1617,N_514);
xor U4508 (N_4508,N_1379,N_1211);
and U4509 (N_4509,N_1229,N_1383);
nor U4510 (N_4510,N_662,N_3018);
or U4511 (N_4511,N_3101,N_3029);
or U4512 (N_4512,N_39,N_2106);
nor U4513 (N_4513,N_1450,N_826);
nand U4514 (N_4514,N_1534,N_1184);
xnor U4515 (N_4515,N_2157,N_2924);
nor U4516 (N_4516,N_2981,N_1883);
nor U4517 (N_4517,N_1455,N_637);
or U4518 (N_4518,N_1377,N_2229);
or U4519 (N_4519,N_1007,N_1339);
or U4520 (N_4520,N_1329,N_2730);
and U4521 (N_4521,N_2107,N_1977);
or U4522 (N_4522,N_188,N_1571);
or U4523 (N_4523,N_2660,N_1667);
nand U4524 (N_4524,N_2180,N_1911);
nand U4525 (N_4525,N_1956,N_2090);
nor U4526 (N_4526,N_2355,N_2635);
or U4527 (N_4527,N_2321,N_1596);
xnor U4528 (N_4528,N_621,N_263);
and U4529 (N_4529,N_1550,N_424);
and U4530 (N_4530,N_2949,N_2636);
nor U4531 (N_4531,N_2456,N_2867);
nor U4532 (N_4532,N_2247,N_479);
xnor U4533 (N_4533,N_1384,N_1768);
xor U4534 (N_4534,N_992,N_840);
and U4535 (N_4535,N_1498,N_2176);
or U4536 (N_4536,N_1145,N_899);
nand U4537 (N_4537,N_2767,N_767);
and U4538 (N_4538,N_2130,N_741);
xnor U4539 (N_4539,N_2947,N_2696);
or U4540 (N_4540,N_2808,N_80);
xor U4541 (N_4541,N_417,N_1057);
xnor U4542 (N_4542,N_2825,N_2052);
xor U4543 (N_4543,N_2534,N_1357);
nor U4544 (N_4544,N_601,N_2268);
nand U4545 (N_4545,N_551,N_307);
and U4546 (N_4546,N_565,N_2128);
nand U4547 (N_4547,N_2368,N_1032);
xnor U4548 (N_4548,N_3089,N_713);
nor U4549 (N_4549,N_1390,N_2626);
xnor U4550 (N_4550,N_1774,N_340);
nor U4551 (N_4551,N_533,N_1998);
nor U4552 (N_4552,N_1564,N_628);
or U4553 (N_4553,N_2841,N_2234);
xor U4554 (N_4554,N_2723,N_2309);
and U4555 (N_4555,N_2780,N_384);
or U4556 (N_4556,N_3039,N_2354);
nor U4557 (N_4557,N_581,N_1062);
and U4558 (N_4558,N_1265,N_1615);
and U4559 (N_4559,N_2523,N_1864);
nand U4560 (N_4560,N_365,N_2988);
xnor U4561 (N_4561,N_1607,N_463);
nor U4562 (N_4562,N_908,N_2269);
nand U4563 (N_4563,N_1496,N_66);
and U4564 (N_4564,N_1042,N_2792);
xnor U4565 (N_4565,N_2030,N_1513);
or U4566 (N_4566,N_2900,N_1622);
nor U4567 (N_4567,N_2871,N_2783);
nand U4568 (N_4568,N_953,N_293);
xor U4569 (N_4569,N_170,N_2991);
nor U4570 (N_4570,N_2946,N_974);
xor U4571 (N_4571,N_677,N_842);
nand U4572 (N_4572,N_364,N_86);
xor U4573 (N_4573,N_40,N_1477);
nand U4574 (N_4574,N_1029,N_1082);
nand U4575 (N_4575,N_428,N_1218);
and U4576 (N_4576,N_582,N_1961);
and U4577 (N_4577,N_2710,N_1742);
and U4578 (N_4578,N_2979,N_2675);
and U4579 (N_4579,N_2240,N_727);
and U4580 (N_4580,N_303,N_515);
nor U4581 (N_4581,N_111,N_666);
nand U4582 (N_4582,N_2226,N_2724);
nor U4583 (N_4583,N_1914,N_2590);
and U4584 (N_4584,N_120,N_2096);
xnor U4585 (N_4585,N_709,N_2203);
xor U4586 (N_4586,N_2137,N_2995);
or U4587 (N_4587,N_866,N_1077);
or U4588 (N_4588,N_2347,N_326);
or U4589 (N_4589,N_2393,N_750);
and U4590 (N_4590,N_1335,N_99);
nand U4591 (N_4591,N_645,N_524);
nor U4592 (N_4592,N_3108,N_2968);
nor U4593 (N_4593,N_716,N_1423);
nor U4594 (N_4594,N_2356,N_2258);
and U4595 (N_4595,N_496,N_2863);
and U4596 (N_4596,N_2920,N_2263);
nor U4597 (N_4597,N_1397,N_2110);
or U4598 (N_4598,N_209,N_1962);
nor U4599 (N_4599,N_2031,N_1347);
xnor U4600 (N_4600,N_1984,N_2272);
nor U4601 (N_4601,N_1387,N_1867);
and U4602 (N_4602,N_2719,N_317);
nor U4603 (N_4603,N_2473,N_749);
nor U4604 (N_4604,N_2270,N_36);
nand U4605 (N_4605,N_2830,N_1176);
nor U4606 (N_4606,N_2225,N_2357);
and U4607 (N_4607,N_3025,N_1491);
nor U4608 (N_4608,N_2348,N_843);
nand U4609 (N_4609,N_3044,N_1031);
or U4610 (N_4610,N_2998,N_1665);
xor U4611 (N_4611,N_926,N_956);
nor U4612 (N_4612,N_532,N_345);
and U4613 (N_4613,N_1414,N_2895);
and U4614 (N_4614,N_1088,N_932);
xor U4615 (N_4615,N_2267,N_1014);
or U4616 (N_4616,N_1350,N_1151);
nand U4617 (N_4617,N_2558,N_895);
xor U4618 (N_4618,N_2974,N_864);
nand U4619 (N_4619,N_1120,N_679);
nor U4620 (N_4620,N_1518,N_1536);
nor U4621 (N_4621,N_1483,N_249);
nand U4622 (N_4622,N_187,N_832);
nand U4623 (N_4623,N_2406,N_639);
nand U4624 (N_4624,N_2279,N_114);
or U4625 (N_4625,N_1886,N_2385);
xor U4626 (N_4626,N_1065,N_1194);
xor U4627 (N_4627,N_2833,N_125);
nand U4628 (N_4628,N_2884,N_2303);
xor U4629 (N_4629,N_1905,N_1584);
xnor U4630 (N_4630,N_2764,N_1231);
nand U4631 (N_4631,N_2655,N_1494);
xor U4632 (N_4632,N_1666,N_2434);
nand U4633 (N_4633,N_1981,N_3111);
xor U4634 (N_4634,N_2772,N_91);
or U4635 (N_4635,N_46,N_150);
xor U4636 (N_4636,N_1036,N_752);
or U4637 (N_4637,N_72,N_1686);
nand U4638 (N_4638,N_2009,N_2510);
nand U4639 (N_4639,N_652,N_1868);
xnor U4640 (N_4640,N_2003,N_2555);
xor U4641 (N_4641,N_1150,N_724);
xor U4642 (N_4642,N_879,N_2896);
xor U4643 (N_4643,N_27,N_1433);
nand U4644 (N_4644,N_1633,N_2572);
and U4645 (N_4645,N_164,N_2182);
nand U4646 (N_4646,N_1199,N_2165);
nand U4647 (N_4647,N_1443,N_2324);
and U4648 (N_4648,N_558,N_1251);
and U4649 (N_4649,N_2330,N_118);
and U4650 (N_4650,N_1845,N_1180);
nor U4651 (N_4651,N_661,N_1485);
xnor U4652 (N_4652,N_2042,N_1772);
xor U4653 (N_4653,N_2392,N_1825);
nor U4654 (N_4654,N_1655,N_2503);
and U4655 (N_4655,N_1066,N_3008);
nor U4656 (N_4656,N_495,N_2160);
nor U4657 (N_4657,N_2853,N_862);
nor U4658 (N_4658,N_252,N_938);
nor U4659 (N_4659,N_1043,N_1152);
and U4660 (N_4660,N_19,N_1583);
nand U4661 (N_4661,N_1389,N_1713);
xnor U4662 (N_4662,N_2111,N_2891);
xnor U4663 (N_4663,N_2595,N_2791);
xnor U4664 (N_4664,N_818,N_2897);
nand U4665 (N_4665,N_2151,N_905);
nand U4666 (N_4666,N_2046,N_1164);
and U4667 (N_4667,N_771,N_1903);
or U4668 (N_4668,N_277,N_21);
or U4669 (N_4669,N_1426,N_1823);
xor U4670 (N_4670,N_2214,N_3073);
or U4671 (N_4671,N_529,N_1734);
and U4672 (N_4672,N_2114,N_904);
nor U4673 (N_4673,N_2951,N_1921);
nor U4674 (N_4674,N_333,N_1952);
and U4675 (N_4675,N_1750,N_451);
nand U4676 (N_4676,N_1566,N_619);
and U4677 (N_4677,N_481,N_1004);
and U4678 (N_4678,N_1537,N_616);
xnor U4679 (N_4679,N_2222,N_687);
nor U4680 (N_4680,N_1490,N_1279);
and U4681 (N_4681,N_2018,N_281);
nor U4682 (N_4682,N_1351,N_1848);
nand U4683 (N_4683,N_1928,N_2329);
xnor U4684 (N_4684,N_809,N_139);
xnor U4685 (N_4685,N_2667,N_937);
xnor U4686 (N_4686,N_2563,N_152);
xnor U4687 (N_4687,N_1002,N_1722);
nand U4688 (N_4688,N_2226,N_102);
nand U4689 (N_4689,N_2621,N_1294);
xor U4690 (N_4690,N_92,N_1381);
nand U4691 (N_4691,N_687,N_2050);
xnor U4692 (N_4692,N_1479,N_2627);
nand U4693 (N_4693,N_2353,N_1348);
nand U4694 (N_4694,N_743,N_1807);
xor U4695 (N_4695,N_2561,N_404);
xor U4696 (N_4696,N_378,N_3049);
or U4697 (N_4697,N_2736,N_1776);
nand U4698 (N_4698,N_981,N_938);
nand U4699 (N_4699,N_1342,N_1121);
or U4700 (N_4700,N_798,N_861);
xnor U4701 (N_4701,N_2050,N_875);
xor U4702 (N_4702,N_2719,N_635);
and U4703 (N_4703,N_911,N_762);
or U4704 (N_4704,N_1174,N_143);
xnor U4705 (N_4705,N_2472,N_2702);
xnor U4706 (N_4706,N_82,N_243);
nand U4707 (N_4707,N_2614,N_1010);
and U4708 (N_4708,N_605,N_725);
nor U4709 (N_4709,N_2526,N_2492);
and U4710 (N_4710,N_172,N_2073);
and U4711 (N_4711,N_2128,N_1418);
xor U4712 (N_4712,N_2778,N_466);
and U4713 (N_4713,N_1386,N_1367);
nand U4714 (N_4714,N_755,N_1812);
nand U4715 (N_4715,N_1754,N_560);
xor U4716 (N_4716,N_797,N_524);
or U4717 (N_4717,N_2958,N_1711);
nand U4718 (N_4718,N_1257,N_164);
xor U4719 (N_4719,N_2051,N_57);
nand U4720 (N_4720,N_1150,N_1076);
and U4721 (N_4721,N_170,N_190);
nor U4722 (N_4722,N_1077,N_466);
nand U4723 (N_4723,N_1107,N_1945);
nor U4724 (N_4724,N_486,N_967);
nand U4725 (N_4725,N_4,N_257);
xor U4726 (N_4726,N_2267,N_1003);
or U4727 (N_4727,N_2354,N_2518);
nand U4728 (N_4728,N_2547,N_200);
and U4729 (N_4729,N_336,N_2111);
and U4730 (N_4730,N_2353,N_2746);
nand U4731 (N_4731,N_791,N_1808);
or U4732 (N_4732,N_1606,N_2930);
nor U4733 (N_4733,N_85,N_338);
xnor U4734 (N_4734,N_632,N_3112);
nor U4735 (N_4735,N_1236,N_1735);
and U4736 (N_4736,N_496,N_2316);
nand U4737 (N_4737,N_2137,N_1939);
xor U4738 (N_4738,N_2592,N_126);
xor U4739 (N_4739,N_668,N_1298);
nor U4740 (N_4740,N_2408,N_2877);
or U4741 (N_4741,N_2291,N_849);
xnor U4742 (N_4742,N_224,N_3021);
xor U4743 (N_4743,N_397,N_1374);
and U4744 (N_4744,N_2784,N_181);
or U4745 (N_4745,N_2482,N_324);
and U4746 (N_4746,N_1822,N_1083);
or U4747 (N_4747,N_1850,N_1292);
nand U4748 (N_4748,N_1076,N_683);
nor U4749 (N_4749,N_650,N_91);
nand U4750 (N_4750,N_2039,N_198);
xor U4751 (N_4751,N_3097,N_2119);
nor U4752 (N_4752,N_663,N_3044);
nand U4753 (N_4753,N_643,N_2868);
xor U4754 (N_4754,N_2377,N_601);
nand U4755 (N_4755,N_2025,N_1249);
nand U4756 (N_4756,N_234,N_1959);
nor U4757 (N_4757,N_2378,N_123);
xor U4758 (N_4758,N_162,N_1275);
or U4759 (N_4759,N_102,N_443);
or U4760 (N_4760,N_2060,N_374);
or U4761 (N_4761,N_431,N_2675);
xnor U4762 (N_4762,N_2562,N_1644);
xnor U4763 (N_4763,N_2264,N_1670);
nand U4764 (N_4764,N_2692,N_890);
or U4765 (N_4765,N_2628,N_1457);
nor U4766 (N_4766,N_216,N_2819);
or U4767 (N_4767,N_980,N_1700);
or U4768 (N_4768,N_1120,N_143);
and U4769 (N_4769,N_1418,N_2513);
or U4770 (N_4770,N_758,N_1497);
nand U4771 (N_4771,N_2124,N_2004);
or U4772 (N_4772,N_2118,N_2238);
or U4773 (N_4773,N_1130,N_1720);
xor U4774 (N_4774,N_2233,N_1393);
nor U4775 (N_4775,N_750,N_1954);
nand U4776 (N_4776,N_1435,N_1273);
nand U4777 (N_4777,N_1787,N_916);
xor U4778 (N_4778,N_177,N_2274);
xor U4779 (N_4779,N_775,N_3108);
or U4780 (N_4780,N_921,N_2712);
nor U4781 (N_4781,N_1998,N_1222);
nand U4782 (N_4782,N_2033,N_2233);
nor U4783 (N_4783,N_46,N_2451);
or U4784 (N_4784,N_2751,N_3122);
xnor U4785 (N_4785,N_1147,N_2157);
nand U4786 (N_4786,N_2984,N_1762);
xor U4787 (N_4787,N_2230,N_1416);
or U4788 (N_4788,N_1837,N_2562);
xnor U4789 (N_4789,N_2327,N_1262);
or U4790 (N_4790,N_2249,N_2999);
or U4791 (N_4791,N_2501,N_3000);
xor U4792 (N_4792,N_1052,N_12);
nand U4793 (N_4793,N_1803,N_2898);
nor U4794 (N_4794,N_924,N_869);
nor U4795 (N_4795,N_3081,N_1764);
or U4796 (N_4796,N_1229,N_1526);
or U4797 (N_4797,N_2523,N_2950);
or U4798 (N_4798,N_1447,N_1020);
nor U4799 (N_4799,N_271,N_3077);
xnor U4800 (N_4800,N_501,N_2197);
nand U4801 (N_4801,N_2857,N_2004);
and U4802 (N_4802,N_1997,N_386);
xor U4803 (N_4803,N_2035,N_2097);
nand U4804 (N_4804,N_431,N_1135);
nor U4805 (N_4805,N_2282,N_2334);
nor U4806 (N_4806,N_1433,N_1788);
nand U4807 (N_4807,N_461,N_1548);
nor U4808 (N_4808,N_332,N_579);
nor U4809 (N_4809,N_2186,N_1392);
nand U4810 (N_4810,N_275,N_2501);
nand U4811 (N_4811,N_2609,N_2500);
or U4812 (N_4812,N_1979,N_2131);
and U4813 (N_4813,N_265,N_2035);
nor U4814 (N_4814,N_1874,N_2827);
nor U4815 (N_4815,N_1407,N_995);
nor U4816 (N_4816,N_906,N_1136);
xor U4817 (N_4817,N_2833,N_351);
and U4818 (N_4818,N_1161,N_490);
or U4819 (N_4819,N_1114,N_1695);
or U4820 (N_4820,N_1586,N_577);
nor U4821 (N_4821,N_65,N_1343);
or U4822 (N_4822,N_54,N_2969);
or U4823 (N_4823,N_1123,N_1874);
xor U4824 (N_4824,N_2910,N_2316);
xnor U4825 (N_4825,N_2307,N_2468);
nand U4826 (N_4826,N_1824,N_149);
nor U4827 (N_4827,N_373,N_1546);
nor U4828 (N_4828,N_301,N_750);
or U4829 (N_4829,N_254,N_1291);
and U4830 (N_4830,N_510,N_363);
nor U4831 (N_4831,N_1101,N_970);
nand U4832 (N_4832,N_74,N_1573);
nand U4833 (N_4833,N_2925,N_1613);
xor U4834 (N_4834,N_915,N_826);
nand U4835 (N_4835,N_634,N_2306);
xnor U4836 (N_4836,N_2552,N_2597);
or U4837 (N_4837,N_134,N_104);
nand U4838 (N_4838,N_1127,N_1144);
nand U4839 (N_4839,N_72,N_457);
and U4840 (N_4840,N_2493,N_1750);
nor U4841 (N_4841,N_114,N_926);
nor U4842 (N_4842,N_1902,N_2413);
nand U4843 (N_4843,N_2077,N_2838);
nor U4844 (N_4844,N_377,N_2419);
nand U4845 (N_4845,N_302,N_2510);
nand U4846 (N_4846,N_529,N_3064);
or U4847 (N_4847,N_2392,N_636);
nor U4848 (N_4848,N_1817,N_2201);
nand U4849 (N_4849,N_2736,N_1780);
xnor U4850 (N_4850,N_2794,N_2574);
xnor U4851 (N_4851,N_1445,N_1217);
nor U4852 (N_4852,N_723,N_801);
and U4853 (N_4853,N_1548,N_940);
nand U4854 (N_4854,N_1468,N_3071);
nand U4855 (N_4855,N_1164,N_1510);
nand U4856 (N_4856,N_599,N_2723);
nand U4857 (N_4857,N_1194,N_2423);
or U4858 (N_4858,N_2084,N_2904);
xnor U4859 (N_4859,N_493,N_1908);
or U4860 (N_4860,N_1855,N_2014);
nand U4861 (N_4861,N_2175,N_214);
xor U4862 (N_4862,N_1284,N_413);
nor U4863 (N_4863,N_2095,N_2467);
nand U4864 (N_4864,N_1297,N_40);
nand U4865 (N_4865,N_1887,N_181);
xnor U4866 (N_4866,N_1264,N_2833);
nor U4867 (N_4867,N_1888,N_181);
xor U4868 (N_4868,N_1962,N_2933);
or U4869 (N_4869,N_755,N_1924);
nand U4870 (N_4870,N_196,N_2674);
xor U4871 (N_4871,N_1052,N_1070);
nor U4872 (N_4872,N_557,N_2906);
or U4873 (N_4873,N_1811,N_714);
nand U4874 (N_4874,N_2080,N_158);
or U4875 (N_4875,N_2943,N_832);
nand U4876 (N_4876,N_687,N_1734);
or U4877 (N_4877,N_390,N_2890);
nand U4878 (N_4878,N_2843,N_2686);
xor U4879 (N_4879,N_1726,N_2234);
nor U4880 (N_4880,N_2824,N_1312);
and U4881 (N_4881,N_2007,N_2250);
nand U4882 (N_4882,N_209,N_508);
nand U4883 (N_4883,N_1651,N_1582);
nand U4884 (N_4884,N_1335,N_2370);
nand U4885 (N_4885,N_336,N_1858);
nand U4886 (N_4886,N_731,N_2711);
xnor U4887 (N_4887,N_2646,N_1902);
nor U4888 (N_4888,N_1588,N_1710);
or U4889 (N_4889,N_2397,N_933);
nor U4890 (N_4890,N_1664,N_1360);
nor U4891 (N_4891,N_1803,N_2926);
nand U4892 (N_4892,N_2416,N_1675);
nor U4893 (N_4893,N_2218,N_1976);
nor U4894 (N_4894,N_2167,N_303);
nor U4895 (N_4895,N_1373,N_2473);
nor U4896 (N_4896,N_1298,N_207);
or U4897 (N_4897,N_1610,N_2720);
or U4898 (N_4898,N_1004,N_333);
xor U4899 (N_4899,N_854,N_1216);
and U4900 (N_4900,N_361,N_3085);
and U4901 (N_4901,N_818,N_1607);
and U4902 (N_4902,N_1582,N_458);
xor U4903 (N_4903,N_1485,N_2939);
xnor U4904 (N_4904,N_2355,N_2653);
xor U4905 (N_4905,N_1195,N_1908);
nand U4906 (N_4906,N_596,N_2791);
and U4907 (N_4907,N_1336,N_1896);
or U4908 (N_4908,N_827,N_3107);
xor U4909 (N_4909,N_1610,N_1428);
or U4910 (N_4910,N_501,N_2460);
and U4911 (N_4911,N_2708,N_412);
xor U4912 (N_4912,N_2954,N_2187);
and U4913 (N_4913,N_372,N_67);
nand U4914 (N_4914,N_3114,N_1776);
or U4915 (N_4915,N_1700,N_1072);
and U4916 (N_4916,N_2128,N_1040);
or U4917 (N_4917,N_1335,N_1739);
nor U4918 (N_4918,N_701,N_2591);
and U4919 (N_4919,N_240,N_2150);
or U4920 (N_4920,N_2938,N_1029);
nand U4921 (N_4921,N_2571,N_875);
xor U4922 (N_4922,N_350,N_2535);
xor U4923 (N_4923,N_1179,N_1948);
or U4924 (N_4924,N_260,N_104);
and U4925 (N_4925,N_121,N_2241);
nor U4926 (N_4926,N_2887,N_2643);
nor U4927 (N_4927,N_936,N_2011);
nand U4928 (N_4928,N_1640,N_2629);
and U4929 (N_4929,N_1845,N_1374);
and U4930 (N_4930,N_29,N_731);
or U4931 (N_4931,N_403,N_2780);
nor U4932 (N_4932,N_1121,N_2987);
or U4933 (N_4933,N_712,N_2686);
or U4934 (N_4934,N_1794,N_2290);
xor U4935 (N_4935,N_3098,N_581);
nand U4936 (N_4936,N_1878,N_1061);
and U4937 (N_4937,N_1235,N_1874);
xnor U4938 (N_4938,N_1327,N_1573);
xor U4939 (N_4939,N_1281,N_2314);
nor U4940 (N_4940,N_401,N_1546);
nor U4941 (N_4941,N_2643,N_1632);
nand U4942 (N_4942,N_2803,N_2332);
and U4943 (N_4943,N_2871,N_282);
xor U4944 (N_4944,N_2968,N_2874);
nand U4945 (N_4945,N_2041,N_100);
xor U4946 (N_4946,N_2922,N_1223);
nor U4947 (N_4947,N_2591,N_2718);
nand U4948 (N_4948,N_3028,N_756);
nor U4949 (N_4949,N_2850,N_105);
or U4950 (N_4950,N_1057,N_1178);
and U4951 (N_4951,N_1499,N_346);
and U4952 (N_4952,N_2026,N_629);
or U4953 (N_4953,N_313,N_2508);
xnor U4954 (N_4954,N_2148,N_554);
xnor U4955 (N_4955,N_1489,N_1143);
xor U4956 (N_4956,N_26,N_831);
nand U4957 (N_4957,N_1327,N_1932);
nand U4958 (N_4958,N_1552,N_1911);
nor U4959 (N_4959,N_2712,N_2308);
or U4960 (N_4960,N_2034,N_2004);
or U4961 (N_4961,N_487,N_689);
and U4962 (N_4962,N_1108,N_543);
or U4963 (N_4963,N_2843,N_658);
xnor U4964 (N_4964,N_914,N_1523);
or U4965 (N_4965,N_1791,N_1945);
and U4966 (N_4966,N_1822,N_1433);
and U4967 (N_4967,N_2426,N_258);
nand U4968 (N_4968,N_1457,N_703);
and U4969 (N_4969,N_1876,N_472);
nand U4970 (N_4970,N_2299,N_410);
or U4971 (N_4971,N_1541,N_1258);
xor U4972 (N_4972,N_1075,N_413);
and U4973 (N_4973,N_2984,N_2596);
nand U4974 (N_4974,N_224,N_1458);
xor U4975 (N_4975,N_2095,N_2129);
nand U4976 (N_4976,N_1132,N_1356);
and U4977 (N_4977,N_716,N_1167);
and U4978 (N_4978,N_391,N_1414);
and U4979 (N_4979,N_2113,N_1882);
nand U4980 (N_4980,N_2175,N_2796);
nor U4981 (N_4981,N_895,N_372);
and U4982 (N_4982,N_2935,N_1184);
or U4983 (N_4983,N_2622,N_1997);
nor U4984 (N_4984,N_1807,N_1296);
nand U4985 (N_4985,N_369,N_1808);
or U4986 (N_4986,N_2465,N_900);
nor U4987 (N_4987,N_1664,N_2331);
nand U4988 (N_4988,N_2154,N_2836);
and U4989 (N_4989,N_129,N_1691);
or U4990 (N_4990,N_1237,N_315);
and U4991 (N_4991,N_772,N_1582);
and U4992 (N_4992,N_2203,N_25);
and U4993 (N_4993,N_2072,N_554);
xnor U4994 (N_4994,N_868,N_1931);
nand U4995 (N_4995,N_2578,N_119);
or U4996 (N_4996,N_1119,N_1342);
nor U4997 (N_4997,N_213,N_1053);
nor U4998 (N_4998,N_45,N_1649);
nor U4999 (N_4999,N_2831,N_1945);
or U5000 (N_5000,N_1311,N_3);
nand U5001 (N_5001,N_183,N_1539);
and U5002 (N_5002,N_211,N_1340);
and U5003 (N_5003,N_429,N_107);
xor U5004 (N_5004,N_589,N_1119);
and U5005 (N_5005,N_1868,N_3087);
or U5006 (N_5006,N_191,N_1738);
and U5007 (N_5007,N_1240,N_2032);
and U5008 (N_5008,N_346,N_944);
xor U5009 (N_5009,N_360,N_2257);
xor U5010 (N_5010,N_3076,N_2350);
nand U5011 (N_5011,N_380,N_1229);
or U5012 (N_5012,N_329,N_2723);
xor U5013 (N_5013,N_417,N_2658);
nor U5014 (N_5014,N_1362,N_925);
or U5015 (N_5015,N_2397,N_1553);
and U5016 (N_5016,N_61,N_1786);
or U5017 (N_5017,N_751,N_2638);
or U5018 (N_5018,N_2532,N_1052);
nor U5019 (N_5019,N_2929,N_1541);
nor U5020 (N_5020,N_2076,N_595);
xnor U5021 (N_5021,N_229,N_735);
xnor U5022 (N_5022,N_875,N_365);
or U5023 (N_5023,N_129,N_2249);
xnor U5024 (N_5024,N_2017,N_3069);
nand U5025 (N_5025,N_382,N_1289);
nand U5026 (N_5026,N_1261,N_619);
xor U5027 (N_5027,N_258,N_834);
nand U5028 (N_5028,N_2702,N_3070);
nor U5029 (N_5029,N_2067,N_279);
or U5030 (N_5030,N_772,N_2738);
nor U5031 (N_5031,N_2585,N_149);
nor U5032 (N_5032,N_706,N_2797);
or U5033 (N_5033,N_2356,N_151);
nand U5034 (N_5034,N_2783,N_1987);
xnor U5035 (N_5035,N_1583,N_1191);
and U5036 (N_5036,N_2021,N_3049);
nor U5037 (N_5037,N_2365,N_1236);
and U5038 (N_5038,N_936,N_2140);
nand U5039 (N_5039,N_1272,N_228);
nand U5040 (N_5040,N_1676,N_2249);
and U5041 (N_5041,N_953,N_2386);
or U5042 (N_5042,N_2513,N_1378);
xnor U5043 (N_5043,N_148,N_1704);
nand U5044 (N_5044,N_2809,N_43);
nor U5045 (N_5045,N_2326,N_1747);
nor U5046 (N_5046,N_1366,N_681);
or U5047 (N_5047,N_3,N_364);
xnor U5048 (N_5048,N_2972,N_1253);
and U5049 (N_5049,N_1751,N_2012);
nand U5050 (N_5050,N_2837,N_1003);
or U5051 (N_5051,N_1463,N_2415);
nor U5052 (N_5052,N_2400,N_911);
and U5053 (N_5053,N_179,N_434);
or U5054 (N_5054,N_2670,N_2083);
xor U5055 (N_5055,N_1955,N_1095);
nor U5056 (N_5056,N_1555,N_1554);
xor U5057 (N_5057,N_1070,N_2619);
nor U5058 (N_5058,N_601,N_867);
nor U5059 (N_5059,N_2288,N_814);
and U5060 (N_5060,N_50,N_753);
xor U5061 (N_5061,N_2224,N_2553);
nor U5062 (N_5062,N_662,N_1856);
xnor U5063 (N_5063,N_2555,N_2078);
xor U5064 (N_5064,N_510,N_1406);
or U5065 (N_5065,N_1213,N_2949);
or U5066 (N_5066,N_2857,N_1437);
nor U5067 (N_5067,N_1856,N_1131);
or U5068 (N_5068,N_2486,N_840);
xor U5069 (N_5069,N_664,N_2751);
nand U5070 (N_5070,N_2633,N_1296);
or U5071 (N_5071,N_1799,N_466);
nand U5072 (N_5072,N_1893,N_1415);
or U5073 (N_5073,N_2949,N_1395);
and U5074 (N_5074,N_815,N_1642);
xnor U5075 (N_5075,N_1008,N_204);
nand U5076 (N_5076,N_437,N_1603);
and U5077 (N_5077,N_2402,N_2811);
nor U5078 (N_5078,N_1205,N_1070);
nand U5079 (N_5079,N_647,N_2413);
or U5080 (N_5080,N_1928,N_3029);
nand U5081 (N_5081,N_671,N_1771);
or U5082 (N_5082,N_3086,N_2695);
and U5083 (N_5083,N_2723,N_325);
and U5084 (N_5084,N_331,N_587);
nand U5085 (N_5085,N_732,N_2641);
or U5086 (N_5086,N_341,N_1169);
and U5087 (N_5087,N_1204,N_3102);
xor U5088 (N_5088,N_20,N_1853);
or U5089 (N_5089,N_2724,N_1690);
nand U5090 (N_5090,N_982,N_2321);
or U5091 (N_5091,N_641,N_1660);
or U5092 (N_5092,N_169,N_155);
and U5093 (N_5093,N_3029,N_1022);
and U5094 (N_5094,N_1475,N_385);
xor U5095 (N_5095,N_1385,N_94);
xnor U5096 (N_5096,N_110,N_3087);
nor U5097 (N_5097,N_2531,N_371);
nor U5098 (N_5098,N_1648,N_709);
or U5099 (N_5099,N_1476,N_659);
nand U5100 (N_5100,N_1878,N_2188);
or U5101 (N_5101,N_2914,N_2539);
nor U5102 (N_5102,N_3041,N_157);
nand U5103 (N_5103,N_795,N_3087);
nand U5104 (N_5104,N_2343,N_1556);
and U5105 (N_5105,N_1592,N_1449);
nor U5106 (N_5106,N_1450,N_2400);
nor U5107 (N_5107,N_1232,N_657);
or U5108 (N_5108,N_1182,N_41);
nor U5109 (N_5109,N_904,N_284);
nor U5110 (N_5110,N_536,N_362);
or U5111 (N_5111,N_1111,N_2767);
nor U5112 (N_5112,N_116,N_2981);
nand U5113 (N_5113,N_1723,N_506);
and U5114 (N_5114,N_845,N_217);
and U5115 (N_5115,N_1652,N_35);
or U5116 (N_5116,N_2192,N_123);
nor U5117 (N_5117,N_1141,N_2988);
nor U5118 (N_5118,N_1254,N_1395);
xor U5119 (N_5119,N_1163,N_2736);
xnor U5120 (N_5120,N_1122,N_997);
nor U5121 (N_5121,N_1776,N_1044);
nand U5122 (N_5122,N_1672,N_1187);
and U5123 (N_5123,N_537,N_463);
or U5124 (N_5124,N_1236,N_130);
nand U5125 (N_5125,N_1962,N_1567);
or U5126 (N_5126,N_2054,N_2246);
or U5127 (N_5127,N_2372,N_2729);
xnor U5128 (N_5128,N_2151,N_2110);
and U5129 (N_5129,N_2687,N_2919);
or U5130 (N_5130,N_3111,N_28);
or U5131 (N_5131,N_99,N_2813);
xor U5132 (N_5132,N_1557,N_777);
and U5133 (N_5133,N_121,N_221);
xor U5134 (N_5134,N_3025,N_302);
and U5135 (N_5135,N_641,N_1658);
or U5136 (N_5136,N_1302,N_2060);
nand U5137 (N_5137,N_832,N_1954);
and U5138 (N_5138,N_1711,N_561);
or U5139 (N_5139,N_2198,N_919);
or U5140 (N_5140,N_1609,N_1771);
nor U5141 (N_5141,N_2851,N_2105);
or U5142 (N_5142,N_2955,N_2357);
nand U5143 (N_5143,N_949,N_697);
xnor U5144 (N_5144,N_613,N_1623);
and U5145 (N_5145,N_1470,N_2935);
and U5146 (N_5146,N_2844,N_1143);
nor U5147 (N_5147,N_2435,N_1911);
and U5148 (N_5148,N_1720,N_1589);
nand U5149 (N_5149,N_2541,N_1517);
or U5150 (N_5150,N_250,N_1721);
xor U5151 (N_5151,N_1161,N_1499);
and U5152 (N_5152,N_182,N_1745);
and U5153 (N_5153,N_1491,N_897);
or U5154 (N_5154,N_1617,N_688);
or U5155 (N_5155,N_1331,N_1418);
nor U5156 (N_5156,N_1228,N_1731);
nand U5157 (N_5157,N_1896,N_160);
xnor U5158 (N_5158,N_1301,N_1428);
xnor U5159 (N_5159,N_1559,N_2390);
and U5160 (N_5160,N_2796,N_2981);
nor U5161 (N_5161,N_807,N_2194);
nor U5162 (N_5162,N_1580,N_1631);
xor U5163 (N_5163,N_2623,N_2119);
xor U5164 (N_5164,N_1596,N_2284);
or U5165 (N_5165,N_1210,N_1379);
nor U5166 (N_5166,N_3031,N_1047);
nand U5167 (N_5167,N_1875,N_1965);
or U5168 (N_5168,N_2034,N_1820);
xor U5169 (N_5169,N_2964,N_2368);
and U5170 (N_5170,N_1527,N_608);
and U5171 (N_5171,N_1036,N_78);
nor U5172 (N_5172,N_2705,N_1414);
and U5173 (N_5173,N_3123,N_1871);
or U5174 (N_5174,N_1806,N_510);
nand U5175 (N_5175,N_383,N_1935);
or U5176 (N_5176,N_489,N_2129);
xor U5177 (N_5177,N_1948,N_2959);
nor U5178 (N_5178,N_877,N_1312);
or U5179 (N_5179,N_1058,N_2434);
and U5180 (N_5180,N_698,N_2481);
or U5181 (N_5181,N_1837,N_381);
xor U5182 (N_5182,N_482,N_626);
and U5183 (N_5183,N_598,N_3088);
or U5184 (N_5184,N_1078,N_1951);
or U5185 (N_5185,N_2703,N_2544);
xor U5186 (N_5186,N_1864,N_82);
xnor U5187 (N_5187,N_2685,N_1721);
nor U5188 (N_5188,N_3077,N_1078);
nand U5189 (N_5189,N_1627,N_41);
xor U5190 (N_5190,N_1760,N_2625);
nor U5191 (N_5191,N_511,N_143);
nand U5192 (N_5192,N_1494,N_429);
nand U5193 (N_5193,N_2397,N_932);
nor U5194 (N_5194,N_2109,N_2611);
and U5195 (N_5195,N_2424,N_455);
xor U5196 (N_5196,N_1348,N_2930);
xnor U5197 (N_5197,N_2258,N_1727);
nor U5198 (N_5198,N_2034,N_2157);
nor U5199 (N_5199,N_2919,N_1853);
or U5200 (N_5200,N_3095,N_2071);
nand U5201 (N_5201,N_3076,N_2056);
or U5202 (N_5202,N_841,N_2006);
nor U5203 (N_5203,N_1555,N_1391);
nand U5204 (N_5204,N_1072,N_1933);
and U5205 (N_5205,N_373,N_1810);
or U5206 (N_5206,N_1021,N_72);
and U5207 (N_5207,N_1613,N_169);
nand U5208 (N_5208,N_2563,N_1309);
or U5209 (N_5209,N_1034,N_1277);
nor U5210 (N_5210,N_882,N_2563);
or U5211 (N_5211,N_2518,N_1162);
xor U5212 (N_5212,N_172,N_2899);
or U5213 (N_5213,N_752,N_1995);
nor U5214 (N_5214,N_2010,N_2812);
or U5215 (N_5215,N_1345,N_2648);
xor U5216 (N_5216,N_2086,N_2749);
and U5217 (N_5217,N_1254,N_3084);
xnor U5218 (N_5218,N_479,N_2241);
xor U5219 (N_5219,N_729,N_2378);
or U5220 (N_5220,N_2136,N_1297);
nor U5221 (N_5221,N_1510,N_2772);
nor U5222 (N_5222,N_554,N_939);
nor U5223 (N_5223,N_1603,N_57);
nor U5224 (N_5224,N_421,N_3094);
or U5225 (N_5225,N_638,N_2649);
xor U5226 (N_5226,N_1233,N_384);
nor U5227 (N_5227,N_1399,N_1811);
nor U5228 (N_5228,N_2202,N_1208);
and U5229 (N_5229,N_1127,N_1225);
xor U5230 (N_5230,N_1817,N_817);
xor U5231 (N_5231,N_2532,N_2743);
xnor U5232 (N_5232,N_1595,N_2125);
and U5233 (N_5233,N_1003,N_615);
nor U5234 (N_5234,N_2240,N_2700);
xor U5235 (N_5235,N_1933,N_2117);
xnor U5236 (N_5236,N_499,N_1241);
xor U5237 (N_5237,N_2528,N_2792);
or U5238 (N_5238,N_99,N_924);
and U5239 (N_5239,N_1090,N_2304);
or U5240 (N_5240,N_2513,N_2113);
nor U5241 (N_5241,N_1294,N_180);
nor U5242 (N_5242,N_3074,N_1983);
or U5243 (N_5243,N_1218,N_2633);
and U5244 (N_5244,N_1175,N_1488);
xor U5245 (N_5245,N_1408,N_777);
nand U5246 (N_5246,N_308,N_206);
nor U5247 (N_5247,N_1177,N_1128);
xor U5248 (N_5248,N_667,N_2778);
nor U5249 (N_5249,N_618,N_3087);
xor U5250 (N_5250,N_2847,N_2689);
nor U5251 (N_5251,N_1145,N_1101);
nand U5252 (N_5252,N_2450,N_2996);
nand U5253 (N_5253,N_1,N_1361);
nor U5254 (N_5254,N_32,N_1535);
or U5255 (N_5255,N_815,N_1128);
nor U5256 (N_5256,N_1901,N_1751);
nor U5257 (N_5257,N_2298,N_2230);
xor U5258 (N_5258,N_832,N_1497);
nand U5259 (N_5259,N_1329,N_1182);
nand U5260 (N_5260,N_1284,N_829);
nand U5261 (N_5261,N_2167,N_1222);
and U5262 (N_5262,N_1618,N_2223);
nand U5263 (N_5263,N_1121,N_307);
xnor U5264 (N_5264,N_440,N_2368);
or U5265 (N_5265,N_40,N_738);
nand U5266 (N_5266,N_2537,N_3046);
and U5267 (N_5267,N_2625,N_2569);
or U5268 (N_5268,N_1407,N_943);
nand U5269 (N_5269,N_2917,N_2309);
nor U5270 (N_5270,N_1720,N_2486);
xor U5271 (N_5271,N_1605,N_118);
xnor U5272 (N_5272,N_1180,N_647);
xor U5273 (N_5273,N_1507,N_968);
nand U5274 (N_5274,N_1862,N_1069);
or U5275 (N_5275,N_2996,N_449);
nand U5276 (N_5276,N_2169,N_181);
and U5277 (N_5277,N_2612,N_934);
nor U5278 (N_5278,N_55,N_111);
or U5279 (N_5279,N_968,N_1083);
xnor U5280 (N_5280,N_152,N_2947);
and U5281 (N_5281,N_775,N_2690);
or U5282 (N_5282,N_3124,N_2595);
or U5283 (N_5283,N_1223,N_1000);
or U5284 (N_5284,N_2776,N_1707);
or U5285 (N_5285,N_10,N_2732);
nand U5286 (N_5286,N_3121,N_2645);
nand U5287 (N_5287,N_1848,N_286);
nor U5288 (N_5288,N_1650,N_623);
or U5289 (N_5289,N_1777,N_2145);
or U5290 (N_5290,N_3089,N_960);
xnor U5291 (N_5291,N_122,N_1685);
nand U5292 (N_5292,N_1163,N_1997);
nand U5293 (N_5293,N_1398,N_1887);
or U5294 (N_5294,N_1241,N_1275);
nand U5295 (N_5295,N_1771,N_2637);
nor U5296 (N_5296,N_2554,N_1258);
xnor U5297 (N_5297,N_1611,N_2318);
or U5298 (N_5298,N_391,N_39);
xnor U5299 (N_5299,N_1822,N_1663);
nand U5300 (N_5300,N_389,N_936);
xnor U5301 (N_5301,N_2475,N_3073);
or U5302 (N_5302,N_2215,N_1367);
and U5303 (N_5303,N_2289,N_1292);
nand U5304 (N_5304,N_790,N_2044);
and U5305 (N_5305,N_2913,N_2704);
nor U5306 (N_5306,N_1832,N_155);
xnor U5307 (N_5307,N_1086,N_1248);
nor U5308 (N_5308,N_246,N_2964);
nor U5309 (N_5309,N_2515,N_918);
xnor U5310 (N_5310,N_1450,N_2869);
xnor U5311 (N_5311,N_1762,N_194);
nor U5312 (N_5312,N_838,N_1017);
nand U5313 (N_5313,N_1851,N_2607);
xnor U5314 (N_5314,N_2107,N_1193);
nand U5315 (N_5315,N_1202,N_1952);
nand U5316 (N_5316,N_288,N_3091);
nor U5317 (N_5317,N_1648,N_915);
nand U5318 (N_5318,N_1311,N_543);
nand U5319 (N_5319,N_9,N_1209);
xor U5320 (N_5320,N_1675,N_1878);
and U5321 (N_5321,N_1676,N_308);
or U5322 (N_5322,N_1747,N_2051);
xor U5323 (N_5323,N_1033,N_766);
nor U5324 (N_5324,N_1647,N_588);
and U5325 (N_5325,N_2571,N_2248);
nor U5326 (N_5326,N_2904,N_2807);
and U5327 (N_5327,N_2461,N_2638);
xnor U5328 (N_5328,N_1871,N_775);
and U5329 (N_5329,N_1986,N_1023);
xor U5330 (N_5330,N_568,N_1056);
xor U5331 (N_5331,N_1113,N_1111);
or U5332 (N_5332,N_1663,N_2843);
nor U5333 (N_5333,N_1140,N_2452);
and U5334 (N_5334,N_79,N_986);
nand U5335 (N_5335,N_1504,N_565);
xor U5336 (N_5336,N_2776,N_2152);
nand U5337 (N_5337,N_2123,N_1722);
nor U5338 (N_5338,N_1919,N_2927);
and U5339 (N_5339,N_615,N_213);
nor U5340 (N_5340,N_245,N_287);
nand U5341 (N_5341,N_1583,N_2808);
nor U5342 (N_5342,N_907,N_1273);
nor U5343 (N_5343,N_2279,N_4);
xor U5344 (N_5344,N_2939,N_912);
and U5345 (N_5345,N_777,N_1160);
nand U5346 (N_5346,N_2226,N_402);
xnor U5347 (N_5347,N_577,N_1870);
xnor U5348 (N_5348,N_1829,N_522);
and U5349 (N_5349,N_570,N_2912);
or U5350 (N_5350,N_61,N_2577);
xnor U5351 (N_5351,N_2200,N_1755);
nand U5352 (N_5352,N_457,N_846);
or U5353 (N_5353,N_2084,N_1416);
xor U5354 (N_5354,N_666,N_804);
and U5355 (N_5355,N_489,N_237);
xor U5356 (N_5356,N_2960,N_1708);
nand U5357 (N_5357,N_2702,N_659);
nand U5358 (N_5358,N_1700,N_1967);
and U5359 (N_5359,N_1045,N_2966);
and U5360 (N_5360,N_424,N_185);
and U5361 (N_5361,N_2462,N_1715);
and U5362 (N_5362,N_185,N_1083);
nor U5363 (N_5363,N_2009,N_2871);
nand U5364 (N_5364,N_846,N_504);
xor U5365 (N_5365,N_1175,N_308);
xnor U5366 (N_5366,N_1795,N_1036);
nand U5367 (N_5367,N_119,N_792);
and U5368 (N_5368,N_633,N_750);
and U5369 (N_5369,N_1825,N_2956);
or U5370 (N_5370,N_2942,N_1587);
nor U5371 (N_5371,N_2504,N_2022);
and U5372 (N_5372,N_842,N_1083);
nand U5373 (N_5373,N_2810,N_658);
or U5374 (N_5374,N_2555,N_1564);
nand U5375 (N_5375,N_1146,N_788);
xnor U5376 (N_5376,N_1877,N_2036);
and U5377 (N_5377,N_1799,N_1721);
nand U5378 (N_5378,N_130,N_2300);
xnor U5379 (N_5379,N_1010,N_744);
nand U5380 (N_5380,N_406,N_1825);
or U5381 (N_5381,N_2094,N_941);
nand U5382 (N_5382,N_606,N_2411);
nand U5383 (N_5383,N_1406,N_2907);
xor U5384 (N_5384,N_1032,N_2612);
xor U5385 (N_5385,N_3045,N_1631);
nor U5386 (N_5386,N_2079,N_1817);
nor U5387 (N_5387,N_1903,N_1782);
and U5388 (N_5388,N_2808,N_2624);
nand U5389 (N_5389,N_1266,N_2678);
nor U5390 (N_5390,N_2532,N_3119);
nor U5391 (N_5391,N_718,N_539);
xor U5392 (N_5392,N_2999,N_2898);
nor U5393 (N_5393,N_1450,N_1966);
and U5394 (N_5394,N_582,N_1647);
or U5395 (N_5395,N_2072,N_711);
or U5396 (N_5396,N_2121,N_424);
xnor U5397 (N_5397,N_1497,N_1090);
or U5398 (N_5398,N_55,N_1286);
nand U5399 (N_5399,N_1692,N_550);
or U5400 (N_5400,N_2639,N_701);
xor U5401 (N_5401,N_2507,N_342);
nor U5402 (N_5402,N_1726,N_380);
and U5403 (N_5403,N_1487,N_1483);
or U5404 (N_5404,N_587,N_2838);
or U5405 (N_5405,N_1389,N_1733);
or U5406 (N_5406,N_635,N_231);
xor U5407 (N_5407,N_2858,N_2277);
nor U5408 (N_5408,N_456,N_1837);
or U5409 (N_5409,N_2502,N_1824);
nand U5410 (N_5410,N_1118,N_1175);
nor U5411 (N_5411,N_1650,N_2046);
xor U5412 (N_5412,N_2688,N_89);
xor U5413 (N_5413,N_524,N_1484);
nand U5414 (N_5414,N_1024,N_3106);
nor U5415 (N_5415,N_1601,N_1516);
nor U5416 (N_5416,N_1362,N_58);
nor U5417 (N_5417,N_1999,N_2185);
and U5418 (N_5418,N_2691,N_1505);
nand U5419 (N_5419,N_249,N_216);
xor U5420 (N_5420,N_1908,N_1809);
nor U5421 (N_5421,N_1891,N_1869);
or U5422 (N_5422,N_94,N_1516);
or U5423 (N_5423,N_3049,N_868);
or U5424 (N_5424,N_1334,N_2176);
and U5425 (N_5425,N_431,N_2272);
xnor U5426 (N_5426,N_764,N_3018);
nor U5427 (N_5427,N_2209,N_991);
nand U5428 (N_5428,N_2888,N_913);
nand U5429 (N_5429,N_367,N_561);
or U5430 (N_5430,N_2223,N_1640);
nand U5431 (N_5431,N_2313,N_2728);
nor U5432 (N_5432,N_3059,N_2147);
and U5433 (N_5433,N_2014,N_2512);
or U5434 (N_5434,N_2543,N_2755);
and U5435 (N_5435,N_2257,N_3049);
nor U5436 (N_5436,N_2095,N_1173);
and U5437 (N_5437,N_967,N_15);
and U5438 (N_5438,N_1848,N_1395);
and U5439 (N_5439,N_1983,N_1179);
nor U5440 (N_5440,N_2578,N_2414);
and U5441 (N_5441,N_2952,N_1935);
xnor U5442 (N_5442,N_2606,N_1650);
or U5443 (N_5443,N_673,N_1027);
nor U5444 (N_5444,N_1546,N_1242);
and U5445 (N_5445,N_742,N_1888);
and U5446 (N_5446,N_1477,N_1865);
nand U5447 (N_5447,N_1194,N_1216);
or U5448 (N_5448,N_28,N_1604);
nand U5449 (N_5449,N_2321,N_2180);
and U5450 (N_5450,N_1478,N_1349);
or U5451 (N_5451,N_1777,N_830);
and U5452 (N_5452,N_775,N_903);
nand U5453 (N_5453,N_2387,N_1616);
nor U5454 (N_5454,N_314,N_1244);
or U5455 (N_5455,N_2988,N_1696);
xor U5456 (N_5456,N_1840,N_2541);
xor U5457 (N_5457,N_1808,N_172);
or U5458 (N_5458,N_658,N_1810);
nor U5459 (N_5459,N_2188,N_2395);
nand U5460 (N_5460,N_799,N_481);
or U5461 (N_5461,N_677,N_2485);
and U5462 (N_5462,N_2082,N_1623);
xnor U5463 (N_5463,N_36,N_770);
xnor U5464 (N_5464,N_1443,N_870);
or U5465 (N_5465,N_3077,N_1636);
nor U5466 (N_5466,N_901,N_6);
nor U5467 (N_5467,N_501,N_1132);
nand U5468 (N_5468,N_1635,N_1959);
nand U5469 (N_5469,N_2142,N_11);
nor U5470 (N_5470,N_2809,N_2255);
nor U5471 (N_5471,N_1049,N_1026);
and U5472 (N_5472,N_373,N_330);
nor U5473 (N_5473,N_1378,N_1379);
and U5474 (N_5474,N_3048,N_2471);
xnor U5475 (N_5475,N_2718,N_262);
and U5476 (N_5476,N_46,N_855);
and U5477 (N_5477,N_1481,N_2196);
or U5478 (N_5478,N_1496,N_2334);
and U5479 (N_5479,N_1226,N_1909);
xor U5480 (N_5480,N_955,N_238);
xor U5481 (N_5481,N_517,N_254);
xor U5482 (N_5482,N_1964,N_120);
nor U5483 (N_5483,N_2786,N_1384);
xor U5484 (N_5484,N_694,N_2874);
and U5485 (N_5485,N_629,N_258);
nand U5486 (N_5486,N_2398,N_848);
xnor U5487 (N_5487,N_2080,N_1532);
nor U5488 (N_5488,N_2896,N_1786);
nand U5489 (N_5489,N_1139,N_1861);
or U5490 (N_5490,N_1705,N_1406);
and U5491 (N_5491,N_1110,N_474);
nand U5492 (N_5492,N_458,N_2324);
nor U5493 (N_5493,N_1595,N_904);
and U5494 (N_5494,N_2304,N_2244);
or U5495 (N_5495,N_1951,N_2285);
nand U5496 (N_5496,N_915,N_2649);
and U5497 (N_5497,N_1482,N_2092);
or U5498 (N_5498,N_1241,N_1557);
or U5499 (N_5499,N_1695,N_1359);
nor U5500 (N_5500,N_1930,N_68);
xor U5501 (N_5501,N_1,N_2549);
and U5502 (N_5502,N_36,N_696);
nand U5503 (N_5503,N_2262,N_2916);
and U5504 (N_5504,N_576,N_1555);
and U5505 (N_5505,N_890,N_1555);
and U5506 (N_5506,N_2093,N_1721);
or U5507 (N_5507,N_953,N_1435);
nand U5508 (N_5508,N_1571,N_1700);
and U5509 (N_5509,N_69,N_712);
xnor U5510 (N_5510,N_2528,N_3047);
and U5511 (N_5511,N_1524,N_737);
xor U5512 (N_5512,N_974,N_2515);
or U5513 (N_5513,N_523,N_1758);
or U5514 (N_5514,N_2469,N_358);
nand U5515 (N_5515,N_238,N_2943);
nor U5516 (N_5516,N_2642,N_368);
or U5517 (N_5517,N_2694,N_94);
or U5518 (N_5518,N_2677,N_48);
or U5519 (N_5519,N_2437,N_2591);
nand U5520 (N_5520,N_2324,N_2671);
and U5521 (N_5521,N_1414,N_1614);
nor U5522 (N_5522,N_1862,N_1743);
xor U5523 (N_5523,N_2028,N_667);
nand U5524 (N_5524,N_1357,N_640);
and U5525 (N_5525,N_2572,N_2603);
and U5526 (N_5526,N_1588,N_580);
nor U5527 (N_5527,N_1619,N_1766);
nand U5528 (N_5528,N_1437,N_2866);
and U5529 (N_5529,N_501,N_158);
xnor U5530 (N_5530,N_1234,N_654);
xor U5531 (N_5531,N_1912,N_1327);
xnor U5532 (N_5532,N_1517,N_639);
nand U5533 (N_5533,N_675,N_2553);
nand U5534 (N_5534,N_3043,N_1367);
and U5535 (N_5535,N_2227,N_845);
and U5536 (N_5536,N_1088,N_140);
and U5537 (N_5537,N_1722,N_801);
nor U5538 (N_5538,N_1474,N_1987);
nand U5539 (N_5539,N_1099,N_326);
xor U5540 (N_5540,N_885,N_1670);
and U5541 (N_5541,N_2269,N_1703);
and U5542 (N_5542,N_2162,N_2793);
xor U5543 (N_5543,N_1780,N_2267);
nor U5544 (N_5544,N_2965,N_1859);
xnor U5545 (N_5545,N_491,N_1619);
nand U5546 (N_5546,N_115,N_2648);
or U5547 (N_5547,N_938,N_851);
and U5548 (N_5548,N_884,N_1738);
and U5549 (N_5549,N_2829,N_707);
nor U5550 (N_5550,N_401,N_2231);
nand U5551 (N_5551,N_529,N_884);
or U5552 (N_5552,N_2576,N_2604);
or U5553 (N_5553,N_3083,N_1643);
and U5554 (N_5554,N_1189,N_2600);
nand U5555 (N_5555,N_3067,N_2488);
and U5556 (N_5556,N_1817,N_587);
and U5557 (N_5557,N_2833,N_2796);
and U5558 (N_5558,N_2620,N_1237);
xnor U5559 (N_5559,N_2403,N_64);
and U5560 (N_5560,N_2220,N_274);
and U5561 (N_5561,N_835,N_795);
xor U5562 (N_5562,N_2019,N_1135);
or U5563 (N_5563,N_1789,N_1927);
and U5564 (N_5564,N_2100,N_159);
or U5565 (N_5565,N_2705,N_429);
nor U5566 (N_5566,N_564,N_1249);
or U5567 (N_5567,N_1574,N_573);
xor U5568 (N_5568,N_2542,N_3069);
and U5569 (N_5569,N_1035,N_241);
xor U5570 (N_5570,N_1735,N_2905);
and U5571 (N_5571,N_303,N_2985);
or U5572 (N_5572,N_1991,N_271);
and U5573 (N_5573,N_469,N_2625);
xnor U5574 (N_5574,N_106,N_955);
xnor U5575 (N_5575,N_1869,N_204);
and U5576 (N_5576,N_344,N_451);
and U5577 (N_5577,N_2839,N_12);
xor U5578 (N_5578,N_2906,N_1186);
nor U5579 (N_5579,N_1314,N_2149);
and U5580 (N_5580,N_1602,N_355);
xor U5581 (N_5581,N_2244,N_1209);
nor U5582 (N_5582,N_2869,N_900);
and U5583 (N_5583,N_34,N_2276);
nand U5584 (N_5584,N_1817,N_41);
and U5585 (N_5585,N_328,N_453);
nor U5586 (N_5586,N_12,N_2588);
and U5587 (N_5587,N_938,N_175);
and U5588 (N_5588,N_2385,N_3124);
xor U5589 (N_5589,N_2554,N_849);
nand U5590 (N_5590,N_3006,N_2612);
xor U5591 (N_5591,N_232,N_1657);
xnor U5592 (N_5592,N_1887,N_2894);
or U5593 (N_5593,N_1725,N_873);
nor U5594 (N_5594,N_2045,N_461);
nor U5595 (N_5595,N_2028,N_1078);
and U5596 (N_5596,N_1514,N_581);
and U5597 (N_5597,N_999,N_2914);
or U5598 (N_5598,N_1868,N_1177);
and U5599 (N_5599,N_2418,N_691);
xnor U5600 (N_5600,N_1749,N_41);
xor U5601 (N_5601,N_15,N_601);
xnor U5602 (N_5602,N_2861,N_2005);
or U5603 (N_5603,N_1517,N_773);
and U5604 (N_5604,N_2027,N_155);
nand U5605 (N_5605,N_505,N_2089);
nand U5606 (N_5606,N_2219,N_984);
or U5607 (N_5607,N_911,N_2855);
nor U5608 (N_5608,N_376,N_901);
or U5609 (N_5609,N_906,N_322);
nand U5610 (N_5610,N_172,N_280);
nor U5611 (N_5611,N_605,N_1651);
nand U5612 (N_5612,N_1310,N_1250);
xnor U5613 (N_5613,N_365,N_527);
or U5614 (N_5614,N_931,N_1263);
and U5615 (N_5615,N_1967,N_377);
or U5616 (N_5616,N_1675,N_1653);
or U5617 (N_5617,N_2702,N_2365);
and U5618 (N_5618,N_418,N_309);
xnor U5619 (N_5619,N_658,N_1935);
or U5620 (N_5620,N_2211,N_1580);
nor U5621 (N_5621,N_2563,N_2861);
nor U5622 (N_5622,N_2043,N_511);
and U5623 (N_5623,N_369,N_1732);
nand U5624 (N_5624,N_375,N_2856);
nand U5625 (N_5625,N_1266,N_86);
nor U5626 (N_5626,N_2748,N_1304);
nor U5627 (N_5627,N_125,N_1092);
nand U5628 (N_5628,N_2395,N_2055);
and U5629 (N_5629,N_2177,N_1995);
nand U5630 (N_5630,N_1260,N_116);
and U5631 (N_5631,N_227,N_1455);
xor U5632 (N_5632,N_2131,N_2568);
and U5633 (N_5633,N_2795,N_2050);
or U5634 (N_5634,N_371,N_2325);
or U5635 (N_5635,N_1062,N_715);
nor U5636 (N_5636,N_1124,N_1620);
nand U5637 (N_5637,N_1806,N_2409);
xnor U5638 (N_5638,N_2063,N_2804);
and U5639 (N_5639,N_61,N_90);
nand U5640 (N_5640,N_1198,N_92);
nor U5641 (N_5641,N_351,N_1127);
and U5642 (N_5642,N_2432,N_2573);
or U5643 (N_5643,N_1404,N_1435);
or U5644 (N_5644,N_1278,N_605);
nor U5645 (N_5645,N_1007,N_1275);
nor U5646 (N_5646,N_1716,N_442);
and U5647 (N_5647,N_548,N_1515);
nand U5648 (N_5648,N_228,N_1478);
xor U5649 (N_5649,N_1352,N_2401);
xor U5650 (N_5650,N_1700,N_798);
or U5651 (N_5651,N_1746,N_415);
or U5652 (N_5652,N_1422,N_533);
and U5653 (N_5653,N_488,N_2678);
nor U5654 (N_5654,N_277,N_2966);
nand U5655 (N_5655,N_201,N_1122);
xnor U5656 (N_5656,N_703,N_2252);
nor U5657 (N_5657,N_184,N_3036);
or U5658 (N_5658,N_2435,N_1845);
or U5659 (N_5659,N_849,N_1044);
xor U5660 (N_5660,N_1118,N_741);
nor U5661 (N_5661,N_1855,N_1387);
or U5662 (N_5662,N_116,N_3006);
and U5663 (N_5663,N_2869,N_950);
or U5664 (N_5664,N_2512,N_1711);
nand U5665 (N_5665,N_1158,N_2774);
or U5666 (N_5666,N_1660,N_2311);
xnor U5667 (N_5667,N_356,N_1044);
and U5668 (N_5668,N_27,N_1303);
nand U5669 (N_5669,N_1294,N_1631);
xnor U5670 (N_5670,N_2705,N_2728);
or U5671 (N_5671,N_1844,N_1964);
xor U5672 (N_5672,N_2287,N_2119);
nand U5673 (N_5673,N_2663,N_2049);
nor U5674 (N_5674,N_1151,N_1782);
or U5675 (N_5675,N_2505,N_2695);
xor U5676 (N_5676,N_1631,N_642);
nand U5677 (N_5677,N_1469,N_1390);
nor U5678 (N_5678,N_1084,N_2801);
nor U5679 (N_5679,N_2610,N_2595);
xnor U5680 (N_5680,N_1997,N_417);
nand U5681 (N_5681,N_444,N_2735);
xnor U5682 (N_5682,N_1998,N_2404);
or U5683 (N_5683,N_2344,N_169);
xor U5684 (N_5684,N_1880,N_3055);
xnor U5685 (N_5685,N_2789,N_812);
nor U5686 (N_5686,N_210,N_422);
and U5687 (N_5687,N_958,N_370);
and U5688 (N_5688,N_1456,N_1073);
or U5689 (N_5689,N_243,N_1967);
nor U5690 (N_5690,N_902,N_1444);
xnor U5691 (N_5691,N_1526,N_1628);
or U5692 (N_5692,N_2522,N_1576);
or U5693 (N_5693,N_2048,N_3097);
xor U5694 (N_5694,N_2018,N_1508);
or U5695 (N_5695,N_473,N_1838);
or U5696 (N_5696,N_2422,N_1186);
xor U5697 (N_5697,N_1713,N_2637);
nor U5698 (N_5698,N_441,N_359);
and U5699 (N_5699,N_553,N_2584);
and U5700 (N_5700,N_1608,N_2512);
and U5701 (N_5701,N_2308,N_2843);
and U5702 (N_5702,N_1232,N_2667);
nor U5703 (N_5703,N_2014,N_123);
nand U5704 (N_5704,N_2816,N_1548);
nand U5705 (N_5705,N_2892,N_1155);
nor U5706 (N_5706,N_418,N_2543);
nor U5707 (N_5707,N_1494,N_2472);
nand U5708 (N_5708,N_1501,N_1404);
xnor U5709 (N_5709,N_2499,N_3122);
nand U5710 (N_5710,N_1999,N_462);
nor U5711 (N_5711,N_600,N_207);
nand U5712 (N_5712,N_1226,N_1373);
and U5713 (N_5713,N_2802,N_1786);
xor U5714 (N_5714,N_1831,N_1990);
xor U5715 (N_5715,N_740,N_1797);
or U5716 (N_5716,N_955,N_2231);
nand U5717 (N_5717,N_2659,N_1879);
or U5718 (N_5718,N_1891,N_182);
xnor U5719 (N_5719,N_808,N_2864);
and U5720 (N_5720,N_101,N_1335);
xnor U5721 (N_5721,N_2477,N_656);
xor U5722 (N_5722,N_2711,N_1141);
or U5723 (N_5723,N_2075,N_135);
nor U5724 (N_5724,N_1821,N_813);
nor U5725 (N_5725,N_442,N_2407);
and U5726 (N_5726,N_993,N_1706);
or U5727 (N_5727,N_2375,N_241);
xnor U5728 (N_5728,N_744,N_829);
xor U5729 (N_5729,N_2400,N_760);
nor U5730 (N_5730,N_346,N_405);
or U5731 (N_5731,N_1534,N_3080);
xor U5732 (N_5732,N_1153,N_805);
nand U5733 (N_5733,N_1679,N_2262);
nand U5734 (N_5734,N_3017,N_1412);
xnor U5735 (N_5735,N_1849,N_1977);
xor U5736 (N_5736,N_1645,N_2982);
or U5737 (N_5737,N_2764,N_1957);
nor U5738 (N_5738,N_215,N_2557);
nand U5739 (N_5739,N_1410,N_2978);
nand U5740 (N_5740,N_2158,N_1024);
and U5741 (N_5741,N_1195,N_1508);
and U5742 (N_5742,N_1578,N_1796);
nand U5743 (N_5743,N_1558,N_957);
or U5744 (N_5744,N_3036,N_2540);
nor U5745 (N_5745,N_757,N_1352);
and U5746 (N_5746,N_327,N_1603);
and U5747 (N_5747,N_2721,N_349);
or U5748 (N_5748,N_253,N_2228);
xor U5749 (N_5749,N_1980,N_34);
or U5750 (N_5750,N_1833,N_2796);
nand U5751 (N_5751,N_663,N_2095);
nand U5752 (N_5752,N_2858,N_512);
and U5753 (N_5753,N_1990,N_1075);
xor U5754 (N_5754,N_265,N_1172);
nor U5755 (N_5755,N_923,N_2961);
or U5756 (N_5756,N_838,N_542);
nor U5757 (N_5757,N_251,N_911);
nor U5758 (N_5758,N_525,N_1363);
nand U5759 (N_5759,N_1127,N_2806);
and U5760 (N_5760,N_1006,N_2636);
nand U5761 (N_5761,N_2722,N_1343);
nand U5762 (N_5762,N_3064,N_3060);
nand U5763 (N_5763,N_2370,N_1948);
nand U5764 (N_5764,N_382,N_981);
nand U5765 (N_5765,N_2918,N_3103);
nor U5766 (N_5766,N_427,N_806);
xnor U5767 (N_5767,N_1060,N_1338);
xor U5768 (N_5768,N_2415,N_2492);
and U5769 (N_5769,N_1469,N_1814);
nor U5770 (N_5770,N_2559,N_2452);
xor U5771 (N_5771,N_101,N_983);
and U5772 (N_5772,N_2382,N_1502);
nor U5773 (N_5773,N_2211,N_498);
or U5774 (N_5774,N_881,N_1561);
nand U5775 (N_5775,N_448,N_1012);
xor U5776 (N_5776,N_574,N_86);
xnor U5777 (N_5777,N_1970,N_2443);
nor U5778 (N_5778,N_2179,N_2628);
nand U5779 (N_5779,N_2824,N_1160);
nor U5780 (N_5780,N_3005,N_2487);
xor U5781 (N_5781,N_2560,N_2107);
and U5782 (N_5782,N_1087,N_1058);
and U5783 (N_5783,N_1448,N_426);
or U5784 (N_5784,N_746,N_117);
nor U5785 (N_5785,N_884,N_1183);
or U5786 (N_5786,N_2091,N_1270);
xor U5787 (N_5787,N_98,N_1943);
xor U5788 (N_5788,N_1230,N_2163);
xnor U5789 (N_5789,N_2648,N_2022);
nand U5790 (N_5790,N_1730,N_706);
xnor U5791 (N_5791,N_1770,N_1357);
nand U5792 (N_5792,N_2878,N_1527);
nor U5793 (N_5793,N_3000,N_1201);
xnor U5794 (N_5794,N_2809,N_2682);
nor U5795 (N_5795,N_1466,N_623);
and U5796 (N_5796,N_1778,N_1045);
xor U5797 (N_5797,N_2694,N_1203);
or U5798 (N_5798,N_1040,N_2319);
xor U5799 (N_5799,N_736,N_792);
nand U5800 (N_5800,N_1465,N_2408);
and U5801 (N_5801,N_1551,N_2683);
nor U5802 (N_5802,N_2762,N_2538);
or U5803 (N_5803,N_614,N_2710);
nor U5804 (N_5804,N_2622,N_1674);
and U5805 (N_5805,N_1084,N_1472);
nand U5806 (N_5806,N_1958,N_2030);
or U5807 (N_5807,N_538,N_2484);
nand U5808 (N_5808,N_2688,N_2150);
nand U5809 (N_5809,N_2669,N_1935);
nand U5810 (N_5810,N_782,N_2403);
and U5811 (N_5811,N_1088,N_1376);
nand U5812 (N_5812,N_1495,N_394);
or U5813 (N_5813,N_75,N_252);
and U5814 (N_5814,N_1272,N_331);
nand U5815 (N_5815,N_2527,N_307);
xnor U5816 (N_5816,N_2798,N_2378);
and U5817 (N_5817,N_166,N_1559);
or U5818 (N_5818,N_1486,N_2048);
xnor U5819 (N_5819,N_150,N_1338);
and U5820 (N_5820,N_2134,N_1808);
nand U5821 (N_5821,N_404,N_2666);
nand U5822 (N_5822,N_1295,N_2402);
xnor U5823 (N_5823,N_2246,N_1846);
xor U5824 (N_5824,N_771,N_114);
and U5825 (N_5825,N_2854,N_1253);
or U5826 (N_5826,N_187,N_540);
nand U5827 (N_5827,N_277,N_2567);
or U5828 (N_5828,N_1302,N_1977);
or U5829 (N_5829,N_2267,N_466);
xor U5830 (N_5830,N_2666,N_573);
nor U5831 (N_5831,N_1351,N_2852);
nor U5832 (N_5832,N_895,N_1465);
or U5833 (N_5833,N_527,N_1004);
nand U5834 (N_5834,N_1164,N_376);
nand U5835 (N_5835,N_1472,N_344);
and U5836 (N_5836,N_2459,N_3099);
and U5837 (N_5837,N_1227,N_2553);
xnor U5838 (N_5838,N_1391,N_1899);
nor U5839 (N_5839,N_2597,N_2372);
and U5840 (N_5840,N_783,N_406);
or U5841 (N_5841,N_882,N_2994);
nand U5842 (N_5842,N_2903,N_2537);
or U5843 (N_5843,N_2596,N_2024);
xor U5844 (N_5844,N_681,N_551);
nand U5845 (N_5845,N_1684,N_2136);
nor U5846 (N_5846,N_1178,N_578);
xor U5847 (N_5847,N_1131,N_264);
and U5848 (N_5848,N_3088,N_1957);
nor U5849 (N_5849,N_2552,N_810);
or U5850 (N_5850,N_1790,N_2989);
xor U5851 (N_5851,N_486,N_2601);
nor U5852 (N_5852,N_2156,N_3112);
or U5853 (N_5853,N_1390,N_1195);
nor U5854 (N_5854,N_2193,N_1852);
and U5855 (N_5855,N_2576,N_3052);
and U5856 (N_5856,N_1007,N_3051);
nor U5857 (N_5857,N_2552,N_2679);
xnor U5858 (N_5858,N_830,N_2369);
nand U5859 (N_5859,N_646,N_1238);
xor U5860 (N_5860,N_755,N_2615);
and U5861 (N_5861,N_2680,N_3045);
xor U5862 (N_5862,N_2690,N_1649);
xor U5863 (N_5863,N_948,N_1591);
or U5864 (N_5864,N_1836,N_810);
nor U5865 (N_5865,N_1311,N_2034);
or U5866 (N_5866,N_2715,N_3022);
nand U5867 (N_5867,N_1167,N_2960);
nand U5868 (N_5868,N_1285,N_1995);
nor U5869 (N_5869,N_1670,N_1817);
nor U5870 (N_5870,N_668,N_2464);
and U5871 (N_5871,N_2114,N_1744);
xnor U5872 (N_5872,N_1145,N_2777);
nor U5873 (N_5873,N_1763,N_3084);
xor U5874 (N_5874,N_1403,N_1813);
nand U5875 (N_5875,N_2216,N_1534);
and U5876 (N_5876,N_698,N_1332);
xor U5877 (N_5877,N_1445,N_2206);
nor U5878 (N_5878,N_2923,N_1047);
nor U5879 (N_5879,N_2019,N_2058);
nor U5880 (N_5880,N_343,N_2169);
and U5881 (N_5881,N_1198,N_1768);
nor U5882 (N_5882,N_108,N_1793);
xnor U5883 (N_5883,N_1384,N_1414);
or U5884 (N_5884,N_2358,N_485);
and U5885 (N_5885,N_508,N_1285);
or U5886 (N_5886,N_1343,N_1505);
nand U5887 (N_5887,N_1684,N_2740);
nand U5888 (N_5888,N_2751,N_2951);
and U5889 (N_5889,N_2850,N_817);
nand U5890 (N_5890,N_2871,N_474);
nand U5891 (N_5891,N_2748,N_2987);
nand U5892 (N_5892,N_1228,N_625);
or U5893 (N_5893,N_1296,N_2058);
or U5894 (N_5894,N_3010,N_2920);
xor U5895 (N_5895,N_2427,N_362);
and U5896 (N_5896,N_2225,N_407);
and U5897 (N_5897,N_1095,N_7);
or U5898 (N_5898,N_965,N_1944);
nand U5899 (N_5899,N_3019,N_704);
xnor U5900 (N_5900,N_450,N_957);
nand U5901 (N_5901,N_1133,N_1659);
or U5902 (N_5902,N_2978,N_2811);
and U5903 (N_5903,N_2770,N_1161);
nor U5904 (N_5904,N_711,N_2827);
and U5905 (N_5905,N_149,N_1033);
nor U5906 (N_5906,N_510,N_55);
or U5907 (N_5907,N_95,N_2854);
nor U5908 (N_5908,N_1013,N_1130);
xnor U5909 (N_5909,N_1049,N_2936);
nand U5910 (N_5910,N_192,N_1659);
nand U5911 (N_5911,N_2244,N_177);
or U5912 (N_5912,N_2292,N_2772);
nor U5913 (N_5913,N_1229,N_1054);
xnor U5914 (N_5914,N_856,N_2182);
or U5915 (N_5915,N_619,N_2476);
nor U5916 (N_5916,N_2277,N_1393);
or U5917 (N_5917,N_1803,N_2004);
or U5918 (N_5918,N_2505,N_1246);
or U5919 (N_5919,N_677,N_3102);
or U5920 (N_5920,N_1989,N_1102);
and U5921 (N_5921,N_607,N_148);
and U5922 (N_5922,N_325,N_1446);
nand U5923 (N_5923,N_184,N_1290);
nor U5924 (N_5924,N_51,N_2206);
and U5925 (N_5925,N_2954,N_1402);
nor U5926 (N_5926,N_608,N_1119);
xnor U5927 (N_5927,N_324,N_2281);
and U5928 (N_5928,N_2953,N_1068);
nor U5929 (N_5929,N_2426,N_2322);
xor U5930 (N_5930,N_623,N_1561);
nor U5931 (N_5931,N_1784,N_1945);
nor U5932 (N_5932,N_2015,N_786);
nand U5933 (N_5933,N_2933,N_2591);
xnor U5934 (N_5934,N_920,N_1598);
or U5935 (N_5935,N_1787,N_2745);
or U5936 (N_5936,N_453,N_1090);
or U5937 (N_5937,N_1547,N_165);
nor U5938 (N_5938,N_1089,N_768);
nor U5939 (N_5939,N_2020,N_3016);
and U5940 (N_5940,N_1223,N_351);
xnor U5941 (N_5941,N_162,N_2757);
nor U5942 (N_5942,N_862,N_1422);
and U5943 (N_5943,N_607,N_1061);
or U5944 (N_5944,N_2153,N_1947);
or U5945 (N_5945,N_199,N_1187);
and U5946 (N_5946,N_174,N_2519);
or U5947 (N_5947,N_1583,N_26);
nand U5948 (N_5948,N_396,N_1229);
nand U5949 (N_5949,N_2600,N_206);
nand U5950 (N_5950,N_3101,N_1400);
xnor U5951 (N_5951,N_2244,N_1667);
xor U5952 (N_5952,N_3022,N_1573);
nor U5953 (N_5953,N_2701,N_404);
and U5954 (N_5954,N_292,N_1389);
or U5955 (N_5955,N_230,N_1643);
nand U5956 (N_5956,N_639,N_3011);
and U5957 (N_5957,N_987,N_2179);
nor U5958 (N_5958,N_2955,N_1983);
xor U5959 (N_5959,N_407,N_1784);
or U5960 (N_5960,N_76,N_103);
or U5961 (N_5961,N_285,N_365);
nor U5962 (N_5962,N_2705,N_1426);
nor U5963 (N_5963,N_2891,N_3084);
or U5964 (N_5964,N_1146,N_2153);
nand U5965 (N_5965,N_63,N_924);
nor U5966 (N_5966,N_2475,N_2940);
xnor U5967 (N_5967,N_2202,N_650);
and U5968 (N_5968,N_1745,N_1972);
nand U5969 (N_5969,N_1040,N_1935);
nor U5970 (N_5970,N_3048,N_1845);
xnor U5971 (N_5971,N_1501,N_2676);
or U5972 (N_5972,N_1270,N_2181);
or U5973 (N_5973,N_2756,N_619);
and U5974 (N_5974,N_482,N_762);
nor U5975 (N_5975,N_1115,N_1847);
and U5976 (N_5976,N_935,N_2160);
nand U5977 (N_5977,N_96,N_2533);
nor U5978 (N_5978,N_2820,N_175);
or U5979 (N_5979,N_2530,N_593);
nor U5980 (N_5980,N_342,N_596);
nor U5981 (N_5981,N_1784,N_1404);
nand U5982 (N_5982,N_2007,N_460);
nor U5983 (N_5983,N_1225,N_77);
nand U5984 (N_5984,N_2830,N_1688);
nor U5985 (N_5985,N_416,N_1016);
nand U5986 (N_5986,N_718,N_983);
nand U5987 (N_5987,N_2531,N_1139);
nand U5988 (N_5988,N_1972,N_2850);
or U5989 (N_5989,N_2760,N_976);
xnor U5990 (N_5990,N_1499,N_885);
or U5991 (N_5991,N_671,N_1619);
nor U5992 (N_5992,N_922,N_2164);
or U5993 (N_5993,N_626,N_2079);
xor U5994 (N_5994,N_1989,N_461);
nand U5995 (N_5995,N_2003,N_2983);
nand U5996 (N_5996,N_2102,N_1344);
nor U5997 (N_5997,N_408,N_806);
nor U5998 (N_5998,N_2265,N_2834);
nor U5999 (N_5999,N_475,N_1265);
or U6000 (N_6000,N_87,N_1322);
and U6001 (N_6001,N_1734,N_1542);
and U6002 (N_6002,N_186,N_452);
nand U6003 (N_6003,N_372,N_412);
or U6004 (N_6004,N_2566,N_1851);
or U6005 (N_6005,N_2613,N_1324);
nand U6006 (N_6006,N_20,N_354);
or U6007 (N_6007,N_741,N_2349);
nor U6008 (N_6008,N_934,N_1487);
nand U6009 (N_6009,N_3111,N_2954);
nand U6010 (N_6010,N_2396,N_1475);
xnor U6011 (N_6011,N_2624,N_1903);
nor U6012 (N_6012,N_1846,N_2165);
and U6013 (N_6013,N_481,N_2481);
or U6014 (N_6014,N_1757,N_694);
or U6015 (N_6015,N_1155,N_1984);
nor U6016 (N_6016,N_681,N_525);
xor U6017 (N_6017,N_1371,N_1722);
nor U6018 (N_6018,N_1076,N_3112);
nand U6019 (N_6019,N_1457,N_2420);
or U6020 (N_6020,N_2384,N_1718);
xor U6021 (N_6021,N_2544,N_404);
nand U6022 (N_6022,N_1438,N_2090);
or U6023 (N_6023,N_1643,N_1650);
nor U6024 (N_6024,N_2574,N_389);
xnor U6025 (N_6025,N_2193,N_220);
and U6026 (N_6026,N_1099,N_2327);
xor U6027 (N_6027,N_2384,N_2233);
or U6028 (N_6028,N_1899,N_574);
nor U6029 (N_6029,N_1179,N_2363);
nor U6030 (N_6030,N_695,N_1100);
or U6031 (N_6031,N_333,N_3005);
nand U6032 (N_6032,N_2897,N_550);
xor U6033 (N_6033,N_2526,N_2849);
xor U6034 (N_6034,N_301,N_1381);
nand U6035 (N_6035,N_1981,N_2865);
and U6036 (N_6036,N_3059,N_2816);
nand U6037 (N_6037,N_771,N_3117);
or U6038 (N_6038,N_2243,N_2272);
or U6039 (N_6039,N_999,N_1024);
nand U6040 (N_6040,N_1367,N_1661);
or U6041 (N_6041,N_327,N_2248);
nor U6042 (N_6042,N_1599,N_2030);
and U6043 (N_6043,N_3002,N_1128);
nand U6044 (N_6044,N_2581,N_159);
nand U6045 (N_6045,N_2377,N_1688);
or U6046 (N_6046,N_1885,N_578);
nand U6047 (N_6047,N_2026,N_814);
nand U6048 (N_6048,N_360,N_2379);
nor U6049 (N_6049,N_1932,N_533);
or U6050 (N_6050,N_862,N_2496);
xnor U6051 (N_6051,N_2336,N_688);
xor U6052 (N_6052,N_1702,N_18);
nand U6053 (N_6053,N_2260,N_2032);
nor U6054 (N_6054,N_1660,N_8);
nor U6055 (N_6055,N_483,N_3012);
and U6056 (N_6056,N_684,N_555);
nor U6057 (N_6057,N_1445,N_2456);
and U6058 (N_6058,N_2392,N_1405);
and U6059 (N_6059,N_2144,N_2630);
nand U6060 (N_6060,N_707,N_2400);
or U6061 (N_6061,N_608,N_2859);
nand U6062 (N_6062,N_2326,N_1909);
nand U6063 (N_6063,N_2602,N_1142);
xor U6064 (N_6064,N_964,N_2833);
xor U6065 (N_6065,N_2222,N_1042);
or U6066 (N_6066,N_2464,N_1835);
xnor U6067 (N_6067,N_299,N_1293);
and U6068 (N_6068,N_28,N_32);
and U6069 (N_6069,N_3123,N_718);
or U6070 (N_6070,N_150,N_1694);
nand U6071 (N_6071,N_1194,N_1108);
and U6072 (N_6072,N_1944,N_2623);
or U6073 (N_6073,N_1617,N_143);
nand U6074 (N_6074,N_2131,N_382);
nand U6075 (N_6075,N_517,N_2284);
xnor U6076 (N_6076,N_1890,N_2869);
xnor U6077 (N_6077,N_1848,N_1034);
nand U6078 (N_6078,N_1625,N_1461);
or U6079 (N_6079,N_205,N_2357);
nand U6080 (N_6080,N_2073,N_2953);
nand U6081 (N_6081,N_1676,N_12);
or U6082 (N_6082,N_1752,N_1903);
xor U6083 (N_6083,N_2623,N_439);
or U6084 (N_6084,N_2838,N_1383);
or U6085 (N_6085,N_1548,N_1097);
or U6086 (N_6086,N_2494,N_1624);
nand U6087 (N_6087,N_2679,N_1651);
and U6088 (N_6088,N_2118,N_2494);
nand U6089 (N_6089,N_2122,N_179);
or U6090 (N_6090,N_563,N_1128);
or U6091 (N_6091,N_1633,N_2990);
and U6092 (N_6092,N_982,N_164);
nand U6093 (N_6093,N_2250,N_1649);
or U6094 (N_6094,N_2806,N_1009);
or U6095 (N_6095,N_2676,N_2520);
or U6096 (N_6096,N_257,N_481);
nor U6097 (N_6097,N_1760,N_905);
xnor U6098 (N_6098,N_486,N_2498);
nor U6099 (N_6099,N_1040,N_2177);
xor U6100 (N_6100,N_1018,N_1869);
nand U6101 (N_6101,N_2586,N_1481);
nand U6102 (N_6102,N_417,N_1147);
or U6103 (N_6103,N_2662,N_347);
nor U6104 (N_6104,N_812,N_3016);
nand U6105 (N_6105,N_1995,N_2071);
nor U6106 (N_6106,N_1014,N_121);
nor U6107 (N_6107,N_18,N_1359);
nor U6108 (N_6108,N_1753,N_1460);
xor U6109 (N_6109,N_2049,N_206);
nand U6110 (N_6110,N_3124,N_932);
and U6111 (N_6111,N_2699,N_1535);
or U6112 (N_6112,N_1629,N_2345);
xor U6113 (N_6113,N_2571,N_334);
nor U6114 (N_6114,N_200,N_3001);
and U6115 (N_6115,N_403,N_2033);
nor U6116 (N_6116,N_1218,N_1863);
xor U6117 (N_6117,N_2443,N_1284);
xnor U6118 (N_6118,N_359,N_853);
nand U6119 (N_6119,N_2569,N_1835);
and U6120 (N_6120,N_2157,N_1440);
nand U6121 (N_6121,N_2326,N_590);
xnor U6122 (N_6122,N_1682,N_1128);
nand U6123 (N_6123,N_661,N_1581);
and U6124 (N_6124,N_1702,N_1202);
xnor U6125 (N_6125,N_1076,N_510);
and U6126 (N_6126,N_1756,N_269);
nor U6127 (N_6127,N_2182,N_500);
xor U6128 (N_6128,N_997,N_1270);
nor U6129 (N_6129,N_2909,N_987);
nand U6130 (N_6130,N_1605,N_2436);
nand U6131 (N_6131,N_2151,N_1739);
or U6132 (N_6132,N_233,N_2733);
nor U6133 (N_6133,N_3016,N_2605);
xnor U6134 (N_6134,N_1105,N_2768);
nand U6135 (N_6135,N_736,N_39);
nand U6136 (N_6136,N_686,N_2702);
nand U6137 (N_6137,N_3090,N_2358);
or U6138 (N_6138,N_55,N_952);
and U6139 (N_6139,N_1501,N_200);
and U6140 (N_6140,N_1212,N_2401);
xnor U6141 (N_6141,N_660,N_2218);
nand U6142 (N_6142,N_1873,N_553);
nand U6143 (N_6143,N_627,N_24);
xor U6144 (N_6144,N_1765,N_2979);
or U6145 (N_6145,N_2704,N_2064);
nor U6146 (N_6146,N_987,N_2846);
nor U6147 (N_6147,N_2863,N_455);
or U6148 (N_6148,N_1751,N_2132);
xnor U6149 (N_6149,N_1453,N_2831);
xnor U6150 (N_6150,N_2544,N_1417);
nand U6151 (N_6151,N_2582,N_2585);
nor U6152 (N_6152,N_343,N_356);
nor U6153 (N_6153,N_2113,N_251);
nand U6154 (N_6154,N_2577,N_1576);
or U6155 (N_6155,N_675,N_360);
and U6156 (N_6156,N_922,N_1829);
nand U6157 (N_6157,N_1078,N_2684);
nand U6158 (N_6158,N_2413,N_3085);
or U6159 (N_6159,N_425,N_1447);
or U6160 (N_6160,N_778,N_3050);
and U6161 (N_6161,N_2889,N_946);
xnor U6162 (N_6162,N_939,N_420);
and U6163 (N_6163,N_59,N_1585);
xor U6164 (N_6164,N_2203,N_3107);
or U6165 (N_6165,N_2873,N_7);
xnor U6166 (N_6166,N_1046,N_2042);
and U6167 (N_6167,N_1349,N_2540);
xnor U6168 (N_6168,N_2232,N_105);
or U6169 (N_6169,N_2833,N_2565);
nand U6170 (N_6170,N_877,N_328);
nand U6171 (N_6171,N_2389,N_1001);
nand U6172 (N_6172,N_996,N_987);
nor U6173 (N_6173,N_1223,N_1807);
and U6174 (N_6174,N_1922,N_1464);
or U6175 (N_6175,N_2348,N_845);
nand U6176 (N_6176,N_1461,N_1898);
nand U6177 (N_6177,N_2783,N_1158);
or U6178 (N_6178,N_1663,N_453);
nand U6179 (N_6179,N_1455,N_2921);
nor U6180 (N_6180,N_3003,N_1491);
xnor U6181 (N_6181,N_630,N_2078);
nand U6182 (N_6182,N_1227,N_1670);
and U6183 (N_6183,N_279,N_1381);
xnor U6184 (N_6184,N_2427,N_2068);
xnor U6185 (N_6185,N_2487,N_2091);
nor U6186 (N_6186,N_129,N_9);
and U6187 (N_6187,N_2923,N_3043);
xor U6188 (N_6188,N_2711,N_1359);
xnor U6189 (N_6189,N_976,N_2970);
or U6190 (N_6190,N_1005,N_808);
xnor U6191 (N_6191,N_1612,N_236);
xor U6192 (N_6192,N_2203,N_216);
nand U6193 (N_6193,N_1144,N_914);
or U6194 (N_6194,N_741,N_1158);
and U6195 (N_6195,N_3022,N_2452);
and U6196 (N_6196,N_1915,N_2142);
nand U6197 (N_6197,N_28,N_1066);
nor U6198 (N_6198,N_2639,N_1927);
or U6199 (N_6199,N_1512,N_1464);
or U6200 (N_6200,N_2030,N_2588);
and U6201 (N_6201,N_2252,N_913);
or U6202 (N_6202,N_2757,N_565);
or U6203 (N_6203,N_2675,N_1519);
and U6204 (N_6204,N_1867,N_1139);
nor U6205 (N_6205,N_2657,N_2900);
or U6206 (N_6206,N_2533,N_2121);
and U6207 (N_6207,N_2726,N_2566);
and U6208 (N_6208,N_820,N_1708);
or U6209 (N_6209,N_2486,N_70);
or U6210 (N_6210,N_1935,N_1140);
or U6211 (N_6211,N_2936,N_1206);
xor U6212 (N_6212,N_2284,N_3036);
xnor U6213 (N_6213,N_687,N_3017);
and U6214 (N_6214,N_1487,N_1372);
xnor U6215 (N_6215,N_1032,N_289);
or U6216 (N_6216,N_1411,N_2891);
nor U6217 (N_6217,N_2118,N_2128);
nor U6218 (N_6218,N_2069,N_717);
and U6219 (N_6219,N_1710,N_406);
nand U6220 (N_6220,N_586,N_1243);
or U6221 (N_6221,N_2138,N_2582);
and U6222 (N_6222,N_1360,N_2180);
nor U6223 (N_6223,N_2257,N_1761);
or U6224 (N_6224,N_1646,N_48);
nand U6225 (N_6225,N_3092,N_63);
nor U6226 (N_6226,N_94,N_1224);
nor U6227 (N_6227,N_580,N_561);
nand U6228 (N_6228,N_452,N_1336);
or U6229 (N_6229,N_2023,N_264);
and U6230 (N_6230,N_36,N_1789);
xnor U6231 (N_6231,N_1208,N_259);
and U6232 (N_6232,N_690,N_2343);
and U6233 (N_6233,N_2689,N_482);
and U6234 (N_6234,N_7,N_31);
xnor U6235 (N_6235,N_458,N_612);
and U6236 (N_6236,N_1849,N_224);
or U6237 (N_6237,N_2166,N_33);
xnor U6238 (N_6238,N_556,N_284);
nor U6239 (N_6239,N_649,N_2161);
xor U6240 (N_6240,N_86,N_679);
or U6241 (N_6241,N_2464,N_2068);
nand U6242 (N_6242,N_1567,N_2672);
xor U6243 (N_6243,N_1362,N_1052);
nor U6244 (N_6244,N_775,N_1062);
xnor U6245 (N_6245,N_317,N_2232);
nor U6246 (N_6246,N_2004,N_824);
nor U6247 (N_6247,N_1787,N_1536);
nand U6248 (N_6248,N_32,N_2093);
nand U6249 (N_6249,N_1345,N_209);
nor U6250 (N_6250,N_3962,N_3955);
nor U6251 (N_6251,N_4669,N_5499);
nor U6252 (N_6252,N_5650,N_5856);
or U6253 (N_6253,N_5232,N_3267);
nor U6254 (N_6254,N_4282,N_3211);
xnor U6255 (N_6255,N_5323,N_4143);
or U6256 (N_6256,N_5713,N_3829);
nand U6257 (N_6257,N_3863,N_4808);
or U6258 (N_6258,N_4363,N_5906);
or U6259 (N_6259,N_3397,N_3920);
nand U6260 (N_6260,N_4259,N_4526);
and U6261 (N_6261,N_3581,N_3885);
and U6262 (N_6262,N_4329,N_4599);
nor U6263 (N_6263,N_3242,N_5596);
xor U6264 (N_6264,N_3391,N_4077);
and U6265 (N_6265,N_4045,N_3159);
or U6266 (N_6266,N_6036,N_3860);
or U6267 (N_6267,N_3518,N_3934);
nor U6268 (N_6268,N_6192,N_4798);
nor U6269 (N_6269,N_5791,N_5172);
nor U6270 (N_6270,N_3879,N_4192);
or U6271 (N_6271,N_3866,N_4863);
nand U6272 (N_6272,N_4425,N_5070);
nor U6273 (N_6273,N_4279,N_4032);
nor U6274 (N_6274,N_5851,N_4223);
nor U6275 (N_6275,N_5628,N_4439);
and U6276 (N_6276,N_3439,N_5029);
nor U6277 (N_6277,N_5349,N_5413);
xnor U6278 (N_6278,N_5289,N_3737);
nor U6279 (N_6279,N_3653,N_5089);
xor U6280 (N_6280,N_3595,N_5110);
and U6281 (N_6281,N_6007,N_3608);
nand U6282 (N_6282,N_5076,N_3620);
nor U6283 (N_6283,N_6043,N_4637);
nor U6284 (N_6284,N_5062,N_3407);
nor U6285 (N_6285,N_4294,N_4281);
nand U6286 (N_6286,N_3871,N_5137);
and U6287 (N_6287,N_5724,N_3149);
and U6288 (N_6288,N_3983,N_5935);
xor U6289 (N_6289,N_6085,N_5972);
or U6290 (N_6290,N_5468,N_4759);
or U6291 (N_6291,N_5126,N_4544);
or U6292 (N_6292,N_3827,N_6119);
or U6293 (N_6293,N_6012,N_3346);
xnor U6294 (N_6294,N_3836,N_5819);
nand U6295 (N_6295,N_4309,N_3999);
nor U6296 (N_6296,N_6199,N_5486);
or U6297 (N_6297,N_3698,N_3393);
and U6298 (N_6298,N_4980,N_4597);
and U6299 (N_6299,N_4606,N_3560);
xnor U6300 (N_6300,N_4810,N_3190);
or U6301 (N_6301,N_5773,N_3508);
nor U6302 (N_6302,N_5585,N_5097);
and U6303 (N_6303,N_5244,N_6161);
and U6304 (N_6304,N_4763,N_5708);
nand U6305 (N_6305,N_4495,N_3376);
and U6306 (N_6306,N_5634,N_4400);
and U6307 (N_6307,N_5396,N_3457);
xor U6308 (N_6308,N_4401,N_3201);
and U6309 (N_6309,N_5037,N_3740);
and U6310 (N_6310,N_5430,N_4058);
xor U6311 (N_6311,N_5604,N_4125);
or U6312 (N_6312,N_4678,N_6134);
and U6313 (N_6313,N_6246,N_3640);
nand U6314 (N_6314,N_3754,N_3292);
and U6315 (N_6315,N_4043,N_4289);
nor U6316 (N_6316,N_4629,N_5250);
and U6317 (N_6317,N_5259,N_3806);
xor U6318 (N_6318,N_3990,N_5941);
or U6319 (N_6319,N_5868,N_4604);
xor U6320 (N_6320,N_4452,N_5831);
and U6321 (N_6321,N_4454,N_4009);
xnor U6322 (N_6322,N_4037,N_3938);
nor U6323 (N_6323,N_4002,N_5385);
nand U6324 (N_6324,N_4104,N_3730);
nand U6325 (N_6325,N_3630,N_4179);
nor U6326 (N_6326,N_5912,N_3358);
and U6327 (N_6327,N_4121,N_4940);
nand U6328 (N_6328,N_5140,N_3789);
and U6329 (N_6329,N_4438,N_5878);
and U6330 (N_6330,N_4951,N_6080);
or U6331 (N_6331,N_4031,N_5154);
nand U6332 (N_6332,N_6178,N_3576);
nor U6333 (N_6333,N_4713,N_4506);
and U6334 (N_6334,N_6213,N_5788);
nand U6335 (N_6335,N_3338,N_6060);
xor U6336 (N_6336,N_6099,N_5228);
xor U6337 (N_6337,N_3341,N_6028);
and U6338 (N_6338,N_4487,N_3588);
or U6339 (N_6339,N_5745,N_5810);
nand U6340 (N_6340,N_3734,N_6015);
and U6341 (N_6341,N_4057,N_5237);
xnor U6342 (N_6342,N_4614,N_3366);
nor U6343 (N_6343,N_6106,N_4735);
or U6344 (N_6344,N_4985,N_3335);
xnor U6345 (N_6345,N_4543,N_3417);
nor U6346 (N_6346,N_4233,N_5759);
nand U6347 (N_6347,N_4308,N_3131);
nand U6348 (N_6348,N_4446,N_4736);
or U6349 (N_6349,N_5007,N_5488);
or U6350 (N_6350,N_3982,N_3347);
and U6351 (N_6351,N_5644,N_4268);
xor U6352 (N_6352,N_5740,N_5956);
nand U6353 (N_6353,N_5083,N_5229);
nor U6354 (N_6354,N_3174,N_4467);
or U6355 (N_6355,N_5735,N_5808);
nand U6356 (N_6356,N_5290,N_3995);
or U6357 (N_6357,N_4062,N_4296);
nor U6358 (N_6358,N_3258,N_3558);
xnor U6359 (N_6359,N_3125,N_5513);
nor U6360 (N_6360,N_4670,N_4335);
nand U6361 (N_6361,N_4626,N_4571);
or U6362 (N_6362,N_4768,N_4398);
xnor U6363 (N_6363,N_3644,N_4803);
nand U6364 (N_6364,N_5509,N_3849);
nor U6365 (N_6365,N_3651,N_3128);
and U6366 (N_6366,N_4159,N_5254);
or U6367 (N_6367,N_3168,N_4065);
xor U6368 (N_6368,N_4396,N_3799);
nand U6369 (N_6369,N_5103,N_5325);
xor U6370 (N_6370,N_6035,N_3780);
nor U6371 (N_6371,N_3485,N_5755);
or U6372 (N_6372,N_4402,N_3848);
nor U6373 (N_6373,N_3276,N_5838);
and U6374 (N_6374,N_4357,N_5960);
xnor U6375 (N_6375,N_6139,N_3898);
or U6376 (N_6376,N_5741,N_3781);
xnor U6377 (N_6377,N_3513,N_4496);
nand U6378 (N_6378,N_5682,N_3418);
or U6379 (N_6379,N_5982,N_5291);
nor U6380 (N_6380,N_3900,N_5054);
or U6381 (N_6381,N_5109,N_4246);
xor U6382 (N_6382,N_6046,N_4051);
xnor U6383 (N_6383,N_4237,N_4576);
xor U6384 (N_6384,N_4177,N_4094);
or U6385 (N_6385,N_3176,N_5382);
xnor U6386 (N_6386,N_5936,N_4587);
nand U6387 (N_6387,N_4146,N_5583);
or U6388 (N_6388,N_3833,N_4845);
nand U6389 (N_6389,N_4039,N_6075);
or U6390 (N_6390,N_6077,N_3818);
nand U6391 (N_6391,N_4727,N_3476);
xnor U6392 (N_6392,N_6102,N_5777);
xnor U6393 (N_6393,N_3456,N_5948);
nand U6394 (N_6394,N_5093,N_3923);
and U6395 (N_6395,N_6222,N_6150);
and U6396 (N_6396,N_5836,N_4564);
xor U6397 (N_6397,N_3590,N_5113);
xor U6398 (N_6398,N_4144,N_5647);
nand U6399 (N_6399,N_5309,N_5204);
or U6400 (N_6400,N_3205,N_3804);
and U6401 (N_6401,N_4119,N_5171);
xor U6402 (N_6402,N_5961,N_3636);
nor U6403 (N_6403,N_3895,N_3615);
nand U6404 (N_6404,N_4910,N_5099);
nor U6405 (N_6405,N_4026,N_3197);
or U6406 (N_6406,N_4310,N_5580);
and U6407 (N_6407,N_5293,N_3728);
or U6408 (N_6408,N_4962,N_3770);
nand U6409 (N_6409,N_4064,N_6048);
nor U6410 (N_6410,N_3252,N_3707);
nor U6411 (N_6411,N_3474,N_3275);
xor U6412 (N_6412,N_5623,N_4858);
and U6413 (N_6413,N_5132,N_3237);
nand U6414 (N_6414,N_5920,N_4277);
nand U6415 (N_6415,N_5267,N_4802);
nand U6416 (N_6416,N_4372,N_4134);
nand U6417 (N_6417,N_5142,N_5192);
nor U6418 (N_6418,N_4163,N_4287);
nand U6419 (N_6419,N_4076,N_5698);
nand U6420 (N_6420,N_5241,N_6142);
and U6421 (N_6421,N_4381,N_4020);
xor U6422 (N_6422,N_4038,N_3148);
xor U6423 (N_6423,N_5279,N_5532);
xor U6424 (N_6424,N_3514,N_4515);
nand U6425 (N_6425,N_5129,N_5928);
xor U6426 (N_6426,N_5220,N_5921);
nor U6427 (N_6427,N_3160,N_4346);
nor U6428 (N_6428,N_3984,N_4389);
xor U6429 (N_6429,N_5150,N_3154);
or U6430 (N_6430,N_3910,N_4965);
nor U6431 (N_6431,N_4998,N_5749);
nor U6432 (N_6432,N_4750,N_3175);
nor U6433 (N_6433,N_4646,N_4572);
nor U6434 (N_6434,N_3771,N_4238);
nor U6435 (N_6435,N_3844,N_4241);
and U6436 (N_6436,N_4405,N_4332);
nand U6437 (N_6437,N_5876,N_5200);
xnor U6438 (N_6438,N_4416,N_3941);
nor U6439 (N_6439,N_3388,N_3579);
nand U6440 (N_6440,N_3214,N_5832);
and U6441 (N_6441,N_5642,N_4099);
nand U6442 (N_6442,N_4753,N_3629);
nand U6443 (N_6443,N_5009,N_4014);
and U6444 (N_6444,N_5575,N_4874);
xor U6445 (N_6445,N_3127,N_4362);
nor U6446 (N_6446,N_5752,N_4929);
or U6447 (N_6447,N_3892,N_5760);
xnor U6448 (N_6448,N_5169,N_3759);
xnor U6449 (N_6449,N_5315,N_5611);
nor U6450 (N_6450,N_4554,N_4538);
and U6451 (N_6451,N_3178,N_3989);
nor U6452 (N_6452,N_3956,N_5010);
or U6453 (N_6453,N_3297,N_5023);
nor U6454 (N_6454,N_3419,N_5577);
nand U6455 (N_6455,N_4377,N_3310);
or U6456 (N_6456,N_4541,N_4741);
nor U6457 (N_6457,N_4240,N_3427);
xor U6458 (N_6458,N_5034,N_4973);
xor U6459 (N_6459,N_6066,N_6182);
and U6460 (N_6460,N_3230,N_4876);
or U6461 (N_6461,N_5535,N_5873);
xor U6462 (N_6462,N_4843,N_5633);
or U6463 (N_6463,N_5081,N_4726);
or U6464 (N_6464,N_3313,N_6074);
or U6465 (N_6465,N_6189,N_4537);
or U6466 (N_6466,N_4354,N_4872);
xnor U6467 (N_6467,N_5612,N_4050);
xor U6468 (N_6468,N_4434,N_3426);
or U6469 (N_6469,N_5043,N_4024);
nor U6470 (N_6470,N_4790,N_4138);
and U6471 (N_6471,N_5201,N_5122);
nor U6472 (N_6472,N_5545,N_4431);
nand U6473 (N_6473,N_4285,N_3890);
xor U6474 (N_6474,N_4658,N_3279);
and U6475 (N_6475,N_5608,N_5701);
nand U6476 (N_6476,N_5304,N_4857);
nand U6477 (N_6477,N_5094,N_5319);
xnor U6478 (N_6478,N_3626,N_4818);
nor U6479 (N_6479,N_3855,N_5227);
xnor U6480 (N_6480,N_4918,N_4437);
nand U6481 (N_6481,N_5959,N_5915);
xnor U6482 (N_6482,N_3975,N_3501);
nor U6483 (N_6483,N_5216,N_3834);
xor U6484 (N_6484,N_5834,N_6073);
xor U6485 (N_6485,N_5340,N_5953);
nor U6486 (N_6486,N_4114,N_3339);
nand U6487 (N_6487,N_4673,N_3839);
nand U6488 (N_6488,N_3449,N_3538);
or U6489 (N_6489,N_4888,N_3673);
or U6490 (N_6490,N_4687,N_6173);
xnor U6491 (N_6491,N_5531,N_4414);
nand U6492 (N_6492,N_3304,N_4262);
xnor U6493 (N_6493,N_4008,N_5722);
nand U6494 (N_6494,N_3546,N_3343);
and U6495 (N_6495,N_4822,N_3927);
nand U6496 (N_6496,N_3696,N_5406);
or U6497 (N_6497,N_5747,N_5782);
or U6498 (N_6498,N_4005,N_3389);
nor U6499 (N_6499,N_3210,N_3869);
nand U6500 (N_6500,N_5733,N_4707);
nand U6501 (N_6501,N_4620,N_4862);
nand U6502 (N_6502,N_3566,N_4089);
and U6503 (N_6503,N_4110,N_3464);
xor U6504 (N_6504,N_5994,N_3878);
or U6505 (N_6505,N_5742,N_4084);
nand U6506 (N_6506,N_5166,N_5729);
nor U6507 (N_6507,N_5886,N_3370);
or U6508 (N_6508,N_5805,N_5648);
or U6509 (N_6509,N_6013,N_3202);
and U6510 (N_6510,N_3675,N_5449);
xnor U6511 (N_6511,N_4088,N_4482);
and U6512 (N_6512,N_4216,N_3659);
or U6513 (N_6513,N_5840,N_6176);
or U6514 (N_6514,N_3598,N_4767);
and U6515 (N_6515,N_4636,N_5073);
or U6516 (N_6516,N_3606,N_4981);
xnor U6517 (N_6517,N_3460,N_3811);
nor U6518 (N_6518,N_3935,N_4519);
or U6519 (N_6519,N_5591,N_5434);
nand U6520 (N_6520,N_3667,N_3716);
or U6521 (N_6521,N_3355,N_5390);
and U6522 (N_6522,N_3243,N_4536);
or U6523 (N_6523,N_4080,N_5374);
nand U6524 (N_6524,N_5802,N_5860);
or U6525 (N_6525,N_5669,N_5700);
or U6526 (N_6526,N_4469,N_3932);
xor U6527 (N_6527,N_3200,N_4601);
and U6528 (N_6528,N_3583,N_4214);
nand U6529 (N_6529,N_5523,N_5990);
and U6530 (N_6530,N_4397,N_3263);
and U6531 (N_6531,N_6041,N_4807);
nor U6532 (N_6532,N_3585,N_5639);
nor U6533 (N_6533,N_4926,N_4001);
and U6534 (N_6534,N_4718,N_5621);
nor U6535 (N_6535,N_3374,N_5662);
xnor U6536 (N_6536,N_5947,N_5756);
nor U6537 (N_6537,N_6061,N_3877);
xor U6538 (N_6538,N_3520,N_5436);
and U6539 (N_6539,N_6067,N_5493);
xnor U6540 (N_6540,N_3163,N_3798);
and U6541 (N_6541,N_5170,N_4117);
and U6542 (N_6542,N_5426,N_4324);
nand U6543 (N_6543,N_4896,N_3628);
or U6544 (N_6544,N_5550,N_3563);
nand U6545 (N_6545,N_3847,N_5746);
nand U6546 (N_6546,N_5461,N_4004);
nor U6547 (N_6547,N_3461,N_3968);
nand U6548 (N_6548,N_5125,N_5260);
nor U6549 (N_6549,N_4960,N_4817);
and U6550 (N_6550,N_4685,N_5275);
nand U6551 (N_6551,N_5173,N_4352);
nand U6552 (N_6552,N_4333,N_5276);
nand U6553 (N_6553,N_4663,N_3348);
or U6554 (N_6554,N_5992,N_5217);
xnor U6555 (N_6555,N_5401,N_3532);
xnor U6556 (N_6556,N_5653,N_4447);
xnor U6557 (N_6557,N_3515,N_3140);
and U6558 (N_6558,N_5078,N_6023);
xnor U6559 (N_6559,N_3238,N_4343);
nor U6560 (N_6560,N_5570,N_4725);
or U6561 (N_6561,N_3592,N_4945);
xnor U6562 (N_6562,N_6056,N_5632);
nor U6563 (N_6563,N_6183,N_3749);
or U6564 (N_6564,N_5999,N_5578);
and U6565 (N_6565,N_5177,N_3580);
nor U6566 (N_6566,N_5636,N_5333);
nor U6567 (N_6567,N_5167,N_3674);
or U6568 (N_6568,N_5444,N_5312);
xor U6569 (N_6569,N_5183,N_5019);
and U6570 (N_6570,N_5557,N_3250);
nor U6571 (N_6571,N_3881,N_5600);
nor U6572 (N_6572,N_4589,N_4605);
or U6573 (N_6573,N_4877,N_4665);
nor U6574 (N_6574,N_5822,N_4625);
nor U6575 (N_6575,N_5984,N_6138);
and U6576 (N_6576,N_5651,N_4194);
nor U6577 (N_6577,N_5770,N_5280);
nand U6578 (N_6578,N_6201,N_4970);
or U6579 (N_6579,N_3828,N_3790);
xor U6580 (N_6580,N_3188,N_4303);
or U6581 (N_6581,N_4832,N_5904);
nor U6582 (N_6582,N_3795,N_4697);
nand U6583 (N_6583,N_3684,N_5067);
nand U6584 (N_6584,N_5442,N_6208);
nand U6585 (N_6585,N_5606,N_5041);
and U6586 (N_6586,N_4201,N_3782);
or U6587 (N_6587,N_4695,N_5929);
nor U6588 (N_6588,N_6093,N_3721);
or U6589 (N_6589,N_3484,N_3356);
nor U6590 (N_6590,N_6127,N_4488);
xor U6591 (N_6591,N_3886,N_4860);
xnor U6592 (N_6592,N_4299,N_5336);
nor U6593 (N_6593,N_5869,N_4947);
nor U6594 (N_6594,N_5652,N_3976);
and U6595 (N_6595,N_3255,N_3785);
nand U6596 (N_6596,N_6242,N_4327);
and U6597 (N_6597,N_5341,N_5607);
nand U6598 (N_6598,N_3948,N_4445);
or U6599 (N_6599,N_4886,N_4473);
nor U6600 (N_6600,N_4920,N_5123);
or U6601 (N_6601,N_4996,N_4430);
nor U6602 (N_6602,N_4100,N_4046);
and U6603 (N_6603,N_4856,N_5222);
or U6604 (N_6604,N_3981,N_6070);
nor U6605 (N_6605,N_3413,N_5505);
and U6606 (N_6606,N_5190,N_5894);
or U6607 (N_6607,N_3224,N_5605);
and U6608 (N_6608,N_4567,N_5437);
or U6609 (N_6609,N_3711,N_4603);
xnor U6610 (N_6610,N_3565,N_4272);
xnor U6611 (N_6611,N_3195,N_3246);
nand U6612 (N_6612,N_4632,N_5405);
and U6613 (N_6613,N_3233,N_4200);
nand U6614 (N_6614,N_4645,N_6137);
nor U6615 (N_6615,N_4251,N_4513);
and U6616 (N_6616,N_3564,N_3405);
or U6617 (N_6617,N_6230,N_3908);
or U6618 (N_6618,N_3854,N_5983);
xnor U6619 (N_6619,N_3499,N_6057);
and U6620 (N_6620,N_3302,N_5556);
xnor U6621 (N_6621,N_5875,N_3952);
or U6622 (N_6622,N_6218,N_5448);
and U6623 (N_6623,N_5817,N_3777);
and U6624 (N_6624,N_5900,N_3153);
xnor U6625 (N_6625,N_5416,N_4212);
nor U6626 (N_6626,N_4471,N_4185);
nor U6627 (N_6627,N_4992,N_4879);
or U6628 (N_6628,N_4484,N_6006);
nand U6629 (N_6629,N_5358,N_3745);
nor U6630 (N_6630,N_4356,N_5625);
nand U6631 (N_6631,N_5627,N_4859);
nor U6632 (N_6632,N_4149,N_5506);
nand U6633 (N_6633,N_3800,N_5485);
and U6634 (N_6634,N_3151,N_5616);
nand U6635 (N_6635,N_6110,N_5039);
and U6636 (N_6636,N_4854,N_5744);
nor U6637 (N_6637,N_3286,N_4635);
nor U6638 (N_6638,N_5823,N_3398);
xnor U6639 (N_6639,N_5579,N_4115);
nand U6640 (N_6640,N_5008,N_6122);
nor U6641 (N_6641,N_5922,N_4894);
and U6642 (N_6642,N_3979,N_3375);
or U6643 (N_6643,N_4267,N_4561);
nand U6644 (N_6644,N_5618,N_5438);
and U6645 (N_6645,N_3282,N_5695);
xor U6646 (N_6646,N_4740,N_6063);
and U6647 (N_6647,N_3248,N_5049);
xnor U6648 (N_6648,N_5656,N_6162);
xor U6649 (N_6649,N_3787,N_4930);
and U6650 (N_6650,N_5364,N_4805);
xor U6651 (N_6651,N_4771,N_3961);
xor U6652 (N_6652,N_5320,N_3571);
and U6653 (N_6653,N_4855,N_4497);
or U6654 (N_6654,N_5757,N_5558);
and U6655 (N_6655,N_4738,N_5298);
or U6656 (N_6656,N_6129,N_4704);
and U6657 (N_6657,N_5957,N_6207);
or U6658 (N_6658,N_5775,N_3473);
or U6659 (N_6659,N_5356,N_4948);
nor U6660 (N_6660,N_3519,N_5723);
and U6661 (N_6661,N_4588,N_5974);
xnor U6662 (N_6662,N_3488,N_6221);
nor U6663 (N_6663,N_5696,N_4562);
or U6664 (N_6664,N_5910,N_3949);
nor U6665 (N_6665,N_4153,N_6053);
or U6666 (N_6666,N_3340,N_4033);
nor U6667 (N_6667,N_5517,N_4780);
nor U6668 (N_6668,N_5459,N_3319);
or U6669 (N_6669,N_3940,N_5288);
nor U6670 (N_6670,N_5421,N_5111);
nor U6671 (N_6671,N_4978,N_6232);
xor U6672 (N_6672,N_6026,N_4501);
nand U6673 (N_6673,N_4385,N_4834);
and U6674 (N_6674,N_4528,N_6160);
and U6675 (N_6675,N_5381,N_6032);
nand U6676 (N_6676,N_5403,N_5731);
xor U6677 (N_6677,N_3601,N_5326);
or U6678 (N_6678,N_3656,N_3289);
xnor U6679 (N_6679,N_4577,N_6079);
and U6680 (N_6680,N_5680,N_4412);
nand U6681 (N_6681,N_3695,N_4969);
or U6682 (N_6682,N_3776,N_3171);
or U6683 (N_6683,N_4443,N_4475);
nand U6684 (N_6684,N_4905,N_5883);
and U6685 (N_6685,N_4989,N_4022);
or U6686 (N_6686,N_4871,N_3821);
or U6687 (N_6687,N_5131,N_5763);
nor U6688 (N_6688,N_4764,N_4762);
xor U6689 (N_6689,N_6090,N_3451);
nor U6690 (N_6690,N_5311,N_6168);
xor U6691 (N_6691,N_3820,N_3685);
and U6692 (N_6692,N_5563,N_3308);
or U6693 (N_6693,N_3801,N_5626);
nor U6694 (N_6694,N_5958,N_5539);
xnor U6695 (N_6695,N_5512,N_5386);
xnor U6696 (N_6696,N_5828,N_6198);
or U6697 (N_6697,N_3166,N_4092);
nor U6698 (N_6698,N_4427,N_5511);
nor U6699 (N_6699,N_4461,N_4451);
or U6700 (N_6700,N_4770,N_3572);
and U6701 (N_6701,N_5807,N_3550);
or U6702 (N_6702,N_6130,N_3998);
and U6703 (N_6703,N_3368,N_4647);
nor U6704 (N_6704,N_5524,N_4984);
nand U6705 (N_6705,N_3323,N_4339);
or U6706 (N_6706,N_5792,N_4173);
or U6707 (N_6707,N_3991,N_4158);
nand U6708 (N_6708,N_4429,N_3503);
nand U6709 (N_6709,N_5473,N_5354);
and U6710 (N_6710,N_4786,N_4508);
xor U6711 (N_6711,N_5677,N_3494);
and U6712 (N_6712,N_3504,N_6153);
and U6713 (N_6713,N_3281,N_4476);
or U6714 (N_6714,N_4690,N_5453);
xnor U6715 (N_6715,N_5933,N_3134);
xnor U6716 (N_6716,N_4180,N_6054);
xnor U6717 (N_6717,N_4922,N_3602);
xnor U6718 (N_6718,N_3316,N_5898);
nor U6719 (N_6719,N_3783,N_5339);
and U6720 (N_6720,N_4566,N_3322);
or U6721 (N_6721,N_5977,N_3187);
nor U6722 (N_6722,N_4677,N_3317);
and U6723 (N_6723,N_4480,N_4183);
and U6724 (N_6724,N_4379,N_4003);
or U6725 (N_6725,N_4231,N_3650);
nor U6726 (N_6726,N_4680,N_5527);
nor U6727 (N_6727,N_4982,N_4974);
xor U6728 (N_6728,N_4191,N_5771);
nand U6729 (N_6729,N_3573,N_3215);
xnor U6730 (N_6730,N_4866,N_5263);
xnor U6731 (N_6731,N_3345,N_5568);
nand U6732 (N_6732,N_3902,N_3996);
nand U6733 (N_6733,N_4893,N_5294);
nand U6734 (N_6734,N_5681,N_4952);
nand U6735 (N_6735,N_5397,N_4732);
and U6736 (N_6736,N_5937,N_4055);
nand U6737 (N_6737,N_3665,N_5712);
nand U6738 (N_6738,N_6109,N_6017);
nor U6739 (N_6739,N_6155,N_5016);
xor U6740 (N_6740,N_5938,N_5353);
nor U6741 (N_6741,N_4581,N_3823);
and U6742 (N_6742,N_4028,N_5661);
nor U6743 (N_6743,N_3192,N_3360);
or U6744 (N_6744,N_4007,N_3733);
xor U6745 (N_6745,N_5955,N_3880);
and U6746 (N_6746,N_6247,N_4844);
or U6747 (N_6747,N_3138,N_4242);
nand U6748 (N_6748,N_3137,N_4784);
or U6749 (N_6749,N_4986,N_5998);
nand U6750 (N_6750,N_3765,N_4491);
and U6751 (N_6751,N_3325,N_5199);
xnor U6752 (N_6752,N_3332,N_4934);
nor U6753 (N_6753,N_5240,N_5417);
xor U6754 (N_6754,N_5544,N_4164);
nor U6755 (N_6755,N_5063,N_6163);
nor U6756 (N_6756,N_4916,N_3865);
and U6757 (N_6757,N_4322,N_5065);
nor U6758 (N_6758,N_6194,N_4371);
or U6759 (N_6759,N_5826,N_5362);
nand U6760 (N_6760,N_3150,N_5683);
xor U6761 (N_6761,N_6167,N_4331);
and U6762 (N_6762,N_5145,N_5458);
and U6763 (N_6763,N_5986,N_3570);
nor U6764 (N_6764,N_4071,N_5197);
nand U6765 (N_6765,N_4304,N_3220);
and U6766 (N_6766,N_3856,N_4837);
or U6767 (N_6767,N_5985,N_4107);
and U6768 (N_6768,N_4326,N_5945);
nor U6769 (N_6769,N_4901,N_3784);
xor U6770 (N_6770,N_3305,N_4456);
xor U6771 (N_6771,N_3509,N_4895);
and U6772 (N_6772,N_3157,N_5026);
xnor U6773 (N_6773,N_4345,N_4234);
nand U6774 (N_6774,N_3363,N_5489);
or U6775 (N_6775,N_6159,N_3529);
nand U6776 (N_6776,N_3859,N_5514);
or U6777 (N_6777,N_4615,N_3162);
nor U6778 (N_6778,N_5660,N_5973);
xnor U6779 (N_6779,N_4025,N_4155);
or U6780 (N_6780,N_4956,N_4529);
nor U6781 (N_6781,N_5051,N_4885);
nand U6782 (N_6782,N_4909,N_4552);
or U6783 (N_6783,N_4426,N_5032);
nand U6784 (N_6784,N_5482,N_3467);
nor U6785 (N_6785,N_4527,N_6095);
nand U6786 (N_6786,N_3625,N_5268);
nor U6787 (N_6787,N_3324,N_3372);
nand U6788 (N_6788,N_4642,N_3307);
nor U6789 (N_6789,N_5889,N_4098);
nor U6790 (N_6790,N_5435,N_3290);
or U6791 (N_6791,N_6111,N_3198);
and U6792 (N_6792,N_3390,N_3496);
nor U6793 (N_6793,N_6236,N_3184);
nor U6794 (N_6794,N_5377,N_5491);
or U6795 (N_6795,N_6022,N_3219);
nand U6796 (N_6796,N_4878,N_5631);
and U6797 (N_6797,N_3971,N_3964);
nand U6798 (N_6798,N_4399,N_5164);
and U6799 (N_6799,N_3654,N_5736);
or U6800 (N_6800,N_5300,N_3870);
or U6801 (N_6801,N_5939,N_5270);
or U6802 (N_6802,N_5086,N_3403);
or U6803 (N_6803,N_3627,N_4424);
nor U6804 (N_6804,N_5143,N_5913);
nor U6805 (N_6805,N_4809,N_4551);
or U6806 (N_6806,N_3973,N_5693);
nand U6807 (N_6807,N_4307,N_4067);
and U6808 (N_6808,N_4518,N_5286);
nor U6809 (N_6809,N_3158,N_3686);
nand U6810 (N_6810,N_3235,N_5987);
and U6811 (N_6811,N_3130,N_4631);
and U6812 (N_6812,N_4435,N_4162);
and U6813 (N_6813,N_5467,N_6125);
and U6814 (N_6814,N_4696,N_5483);
and U6815 (N_6815,N_4791,N_4840);
and U6816 (N_6816,N_4311,N_5710);
nand U6817 (N_6817,N_6187,N_4550);
nor U6818 (N_6818,N_3760,N_6158);
or U6819 (N_6819,N_5720,N_5209);
nor U6820 (N_6820,N_3652,N_6169);
or U6821 (N_6821,N_4648,N_4364);
nor U6822 (N_6822,N_4321,N_3472);
and U6823 (N_6823,N_3542,N_4157);
and U6824 (N_6824,N_3425,N_4968);
nand U6825 (N_6825,N_4788,N_5451);
and U6826 (N_6826,N_4082,N_3622);
nor U6827 (N_6827,N_3462,N_6200);
or U6828 (N_6828,N_5715,N_6069);
and U6829 (N_6829,N_3295,N_4101);
nor U6830 (N_6830,N_5717,N_5899);
nor U6831 (N_6831,N_4072,N_5951);
nand U6832 (N_6832,N_5471,N_4344);
or U6833 (N_6833,N_4761,N_5050);
and U6834 (N_6834,N_4717,N_4702);
nand U6835 (N_6835,N_3265,N_3778);
xor U6836 (N_6836,N_4111,N_3891);
and U6837 (N_6837,N_3873,N_5589);
xnor U6838 (N_6838,N_3517,N_4902);
xor U6839 (N_6839,N_6094,N_4999);
xnor U6840 (N_6840,N_3875,N_3502);
xor U6841 (N_6841,N_3199,N_5727);
nand U6842 (N_6842,N_5441,N_3455);
or U6843 (N_6843,N_5033,N_5017);
or U6844 (N_6844,N_3574,N_5096);
nor U6845 (N_6845,N_4386,N_4560);
and U6846 (N_6846,N_3788,N_5447);
and U6847 (N_6847,N_4066,N_6091);
nor U6848 (N_6848,N_3767,N_4199);
nand U6849 (N_6849,N_5691,N_5888);
xor U6850 (N_6850,N_3300,N_4779);
nor U6851 (N_6851,N_5186,N_5013);
or U6852 (N_6852,N_5574,N_4244);
nand U6853 (N_6853,N_3612,N_5533);
nand U6854 (N_6854,N_5813,N_3541);
or U6855 (N_6855,N_5787,N_5649);
nand U6856 (N_6856,N_4250,N_5077);
xnor U6857 (N_6857,N_4286,N_3277);
nand U6858 (N_6858,N_5163,N_3831);
or U6859 (N_6859,N_4457,N_4306);
or U6860 (N_6860,N_6175,N_4503);
nand U6861 (N_6861,N_5969,N_5785);
nand U6862 (N_6862,N_5784,N_3763);
or U6863 (N_6863,N_5100,N_3642);
nor U6864 (N_6864,N_6118,N_3161);
nor U6865 (N_6865,N_5178,N_3344);
nor U6866 (N_6866,N_5345,N_5484);
xor U6867 (N_6867,N_4773,N_5141);
or U6868 (N_6868,N_4291,N_4351);
xnor U6869 (N_6869,N_5538,N_4574);
nand U6870 (N_6870,N_3846,N_5849);
nor U6871 (N_6871,N_6133,N_5988);
xor U6872 (N_6872,N_5399,N_3619);
nand U6873 (N_6873,N_4085,N_5927);
and U6874 (N_6874,N_3683,N_4093);
xnor U6875 (N_6875,N_3400,N_4584);
or U6876 (N_6876,N_3732,N_4875);
nand U6877 (N_6877,N_3896,N_6003);
and U6878 (N_6878,N_4068,N_5864);
xnor U6879 (N_6879,N_4490,N_4824);
nor U6880 (N_6880,N_5566,N_5375);
nor U6881 (N_6881,N_5146,N_4463);
nor U6882 (N_6882,N_4181,N_4142);
and U6883 (N_6883,N_4300,N_6039);
nand U6884 (N_6884,N_4374,N_4721);
xor U6885 (N_6885,N_3206,N_4706);
xor U6886 (N_6886,N_3662,N_5112);
xor U6887 (N_6887,N_4936,N_5954);
xnor U6888 (N_6888,N_5498,N_3512);
nand U6889 (N_6889,N_6027,N_5398);
nor U6890 (N_6890,N_5641,N_3369);
or U6891 (N_6891,N_4522,N_3303);
or U6892 (N_6892,N_4821,N_5714);
nand U6893 (N_6893,N_6040,N_5857);
xor U6894 (N_6894,N_4147,N_5748);
nand U6895 (N_6895,N_5175,N_5546);
xor U6896 (N_6896,N_5387,N_4075);
or U6897 (N_6897,N_4757,N_4778);
xnor U6898 (N_6898,N_4792,N_4123);
nand U6899 (N_6899,N_5283,N_5404);
or U6900 (N_6900,N_3445,N_3803);
or U6901 (N_6901,N_5835,N_6243);
and U6902 (N_6902,N_4959,N_4851);
and U6903 (N_6903,N_3769,N_5902);
xor U6904 (N_6904,N_6157,N_6064);
nor U6905 (N_6905,N_4220,N_5092);
nand U6906 (N_6906,N_4983,N_5181);
or U6907 (N_6907,N_5562,N_3697);
nand U6908 (N_6908,N_4229,N_5803);
or U6909 (N_6909,N_3431,N_5573);
and U6910 (N_6910,N_4747,N_3977);
nand U6911 (N_6911,N_4018,N_4955);
xor U6912 (N_6912,N_5269,N_4760);
xnor U6913 (N_6913,N_5622,N_4853);
and U6914 (N_6914,N_3555,N_6231);
xor U6915 (N_6915,N_5331,N_3471);
and U6916 (N_6916,N_3852,N_5466);
or U6917 (N_6917,N_3539,N_5025);
nor U6918 (N_6918,N_5045,N_3647);
xnor U6919 (N_6919,N_3208,N_4565);
or U6920 (N_6920,N_4297,N_6037);
nand U6921 (N_6921,N_6084,N_5271);
nor U6922 (N_6922,N_3218,N_4613);
and U6923 (N_6923,N_5496,N_5522);
nand U6924 (N_6924,N_3634,N_3589);
and U6925 (N_6925,N_6191,N_4472);
or U6926 (N_6926,N_5207,N_5128);
xor U6927 (N_6927,N_4384,N_5343);
and U6928 (N_6928,N_4338,N_6216);
and U6929 (N_6929,N_4172,N_6058);
xor U6930 (N_6930,N_6100,N_5159);
nor U6931 (N_6931,N_5247,N_3942);
and U6932 (N_6932,N_3386,N_5106);
and U6933 (N_6933,N_3719,N_5182);
xnor U6934 (N_6934,N_4466,N_4382);
nand U6935 (N_6935,N_5335,N_5411);
nand U6936 (N_6936,N_6217,N_4919);
xor U6937 (N_6937,N_5079,N_5786);
or U6938 (N_6938,N_5135,N_5460);
and U6939 (N_6939,N_5006,N_5764);
nand U6940 (N_6940,N_5425,N_3470);
and U6941 (N_6941,N_6154,N_5882);
or U6942 (N_6942,N_4932,N_3373);
and U6943 (N_6943,N_4585,N_5452);
xnor U6944 (N_6944,N_4942,N_3648);
nor U6945 (N_6945,N_4765,N_5423);
nor U6946 (N_6946,N_6087,N_4972);
nor U6947 (N_6947,N_5214,N_4668);
and U6948 (N_6948,N_4073,N_5351);
or U6949 (N_6949,N_5964,N_4021);
xnor U6950 (N_6950,N_5303,N_4317);
and U6951 (N_6951,N_5863,N_3434);
xnor U6952 (N_6952,N_6146,N_5160);
or U6953 (N_6953,N_3194,N_3835);
or U6954 (N_6954,N_4534,N_3251);
nor U6955 (N_6955,N_4198,N_3280);
or U6956 (N_6956,N_3943,N_4165);
nor U6957 (N_6957,N_3480,N_3946);
and U6958 (N_6958,N_3681,N_4976);
nor U6959 (N_6959,N_5962,N_6092);
and U6960 (N_6960,N_3758,N_4376);
or U6961 (N_6961,N_4776,N_5314);
nand U6962 (N_6962,N_5584,N_3523);
or U6963 (N_6963,N_4411,N_4868);
or U6964 (N_6964,N_5040,N_4660);
nor U6965 (N_6965,N_5750,N_3411);
and U6966 (N_6966,N_4204,N_5620);
and U6967 (N_6967,N_3262,N_5495);
xnor U6968 (N_6968,N_4782,N_4823);
xor U6969 (N_6969,N_4393,N_6011);
xnor U6970 (N_6970,N_6042,N_4775);
nand U6971 (N_6971,N_5324,N_5261);
or U6972 (N_6972,N_4124,N_4010);
or U6973 (N_6973,N_3524,N_5870);
and U6974 (N_6974,N_3337,N_4671);
or U6975 (N_6975,N_4048,N_3186);
or U6976 (N_6976,N_4530,N_5976);
nand U6977 (N_6977,N_4320,N_5370);
or U6978 (N_6978,N_6029,N_5243);
xor U6979 (N_6979,N_5853,N_5038);
nand U6980 (N_6980,N_3475,N_5887);
xnor U6981 (N_6981,N_3193,N_3676);
nand U6982 (N_6982,N_4305,N_3172);
xor U6983 (N_6983,N_3320,N_4319);
or U6984 (N_6984,N_5187,N_5091);
nand U6985 (N_6985,N_4794,N_3378);
and U6986 (N_6986,N_5881,N_4641);
xnor U6987 (N_6987,N_3757,N_4975);
or U6988 (N_6988,N_4899,N_5609);
and U6989 (N_6989,N_3333,N_4908);
and U6990 (N_6990,N_5248,N_3294);
xor U6991 (N_6991,N_5518,N_4301);
and U6992 (N_6992,N_3216,N_5185);
nand U6993 (N_6993,N_3936,N_4095);
nor U6994 (N_6994,N_4913,N_5690);
nand U6995 (N_6995,N_3953,N_4781);
xor U6996 (N_6996,N_4361,N_3424);
xnor U6997 (N_6997,N_6193,N_3381);
or U6998 (N_6998,N_3259,N_3918);
nand U6999 (N_6999,N_4656,N_3567);
and U7000 (N_7000,N_3819,N_4979);
or U7001 (N_7001,N_5932,N_5149);
nor U7002 (N_7002,N_5281,N_3465);
or U7003 (N_7003,N_5360,N_5355);
nor U7004 (N_7004,N_6086,N_3670);
nor U7005 (N_7005,N_3753,N_4903);
and U7006 (N_7006,N_4015,N_5087);
nor U7007 (N_7007,N_5795,N_4370);
nor U7008 (N_7008,N_3505,N_4602);
and U7009 (N_7009,N_4442,N_4053);
and U7010 (N_7010,N_3522,N_5012);
nor U7011 (N_7011,N_5844,N_4505);
or U7012 (N_7012,N_3139,N_3189);
nor U7013 (N_7013,N_3669,N_6083);
nand U7014 (N_7014,N_6072,N_4944);
nor U7015 (N_7015,N_3997,N_3762);
nor U7016 (N_7016,N_5000,N_5981);
nor U7017 (N_7017,N_5024,N_5107);
or U7018 (N_7018,N_6031,N_5213);
and U7019 (N_7019,N_4106,N_5191);
xor U7020 (N_7020,N_5980,N_5119);
nand U7021 (N_7021,N_5376,N_4674);
nor U7022 (N_7022,N_5284,N_5211);
nand U7023 (N_7023,N_5072,N_3796);
or U7024 (N_7024,N_3718,N_5098);
and U7025 (N_7025,N_6195,N_5510);
and U7026 (N_7026,N_3987,N_3483);
xnor U7027 (N_7027,N_3637,N_4532);
or U7028 (N_7028,N_5060,N_6249);
nand U7029 (N_7029,N_3450,N_5069);
and U7030 (N_7030,N_5551,N_3658);
xnor U7031 (N_7031,N_3704,N_5258);
and U7032 (N_7032,N_5116,N_4481);
nand U7033 (N_7033,N_5058,N_5667);
nand U7034 (N_7034,N_4880,N_5157);
and U7035 (N_7035,N_3362,N_5890);
nand U7036 (N_7036,N_5725,N_4553);
xor U7037 (N_7037,N_3768,N_6186);
and U7038 (N_7038,N_4812,N_3293);
or U7039 (N_7039,N_5848,N_5837);
nand U7040 (N_7040,N_5603,N_3921);
nand U7041 (N_7041,N_4190,N_3887);
and U7042 (N_7042,N_4662,N_3677);
nand U7043 (N_7043,N_3575,N_5908);
nand U7044 (N_7044,N_4616,N_4731);
nor U7045 (N_7045,N_3387,N_3406);
nand U7046 (N_7046,N_4793,N_4949);
or U7047 (N_7047,N_4407,N_3631);
xor U7048 (N_7048,N_6215,N_3709);
xor U7049 (N_7049,N_6136,N_3287);
nor U7050 (N_7050,N_3618,N_4766);
and U7051 (N_7051,N_4140,N_3569);
or U7052 (N_7052,N_5738,N_4360);
and U7053 (N_7053,N_5588,N_4128);
or U7054 (N_7054,N_3750,N_3679);
nor U7055 (N_7055,N_4507,N_3551);
and U7056 (N_7056,N_5408,N_4621);
nand U7057 (N_7057,N_4019,N_4276);
nand U7058 (N_7058,N_5654,N_3692);
nand U7059 (N_7059,N_5610,N_5858);
nand U7060 (N_7060,N_4699,N_5602);
or U7061 (N_7061,N_3314,N_5372);
and U7062 (N_7062,N_4630,N_3399);
and U7063 (N_7063,N_5850,N_5867);
nor U7064 (N_7064,N_5365,N_5685);
or U7065 (N_7065,N_3632,N_3705);
or U7066 (N_7066,N_5646,N_4257);
and U7067 (N_7067,N_4689,N_5501);
or U7068 (N_7068,N_6010,N_3965);
nor U7069 (N_7069,N_5637,N_4109);
nor U7070 (N_7070,N_4865,N_5395);
nor U7071 (N_7071,N_5357,N_4924);
nand U7072 (N_7072,N_5011,N_5780);
nor U7073 (N_7073,N_5599,N_4723);
nand U7074 (N_7074,N_3511,N_5402);
nand U7075 (N_7075,N_4742,N_3797);
or U7076 (N_7076,N_5564,N_3738);
or U7077 (N_7077,N_3245,N_5554);
nand U7078 (N_7078,N_3296,N_3239);
or U7079 (N_7079,N_3516,N_3554);
nand U7080 (N_7080,N_3331,N_3623);
xor U7081 (N_7081,N_4745,N_5706);
or U7082 (N_7082,N_5842,N_3227);
xnor U7083 (N_7083,N_5478,N_6209);
nor U7084 (N_7084,N_4349,N_3906);
nor U7085 (N_7085,N_4280,N_4450);
xnor U7086 (N_7086,N_6233,N_4820);
nand U7087 (N_7087,N_4545,N_5565);
and U7088 (N_7088,N_5302,N_3395);
nor U7089 (N_7089,N_5919,N_4210);
or U7090 (N_7090,N_4743,N_5678);
nand U7091 (N_7091,N_5151,N_4698);
nand U7092 (N_7092,N_4988,N_5342);
nand U7093 (N_7093,N_4789,N_5165);
xor U7094 (N_7094,N_6135,N_4269);
nor U7095 (N_7095,N_5018,N_6052);
and U7096 (N_7096,N_3350,N_3329);
nor U7097 (N_7097,N_3851,N_3917);
xor U7098 (N_7098,N_5379,N_4870);
nor U7099 (N_7099,N_6002,N_5475);
or U7100 (N_7100,N_4811,N_5670);
nor U7101 (N_7101,N_3703,N_3525);
xnor U7102 (N_7102,N_4254,N_6103);
xor U7103 (N_7103,N_4593,N_3463);
xnor U7104 (N_7104,N_4408,N_5368);
or U7105 (N_7105,N_6059,N_5970);
or U7106 (N_7106,N_5085,N_4248);
nand U7107 (N_7107,N_4224,N_5824);
or U7108 (N_7108,N_3951,N_6196);
nand U7109 (N_7109,N_4404,N_5893);
xnor U7110 (N_7110,N_5236,N_3888);
and U7111 (N_7111,N_6181,N_4365);
or U7112 (N_7112,N_5202,N_4935);
and U7113 (N_7113,N_5909,N_5056);
xnor U7114 (N_7114,N_6024,N_6088);
or U7115 (N_7115,N_6004,N_4966);
and U7116 (N_7116,N_5115,N_4263);
xnor U7117 (N_7117,N_5176,N_5002);
nand U7118 (N_7118,N_4422,N_4869);
nand U7119 (N_7119,N_3947,N_3993);
and U7120 (N_7120,N_5940,N_5758);
and U7121 (N_7121,N_6234,N_6225);
and U7122 (N_7122,N_3169,N_5774);
xor U7123 (N_7123,N_5555,N_4047);
and U7124 (N_7124,N_3437,N_5586);
or U7125 (N_7125,N_3334,N_5071);
nand U7126 (N_7126,N_3147,N_5761);
nor U7127 (N_7127,N_5776,N_4828);
and U7128 (N_7128,N_5549,N_3191);
or U7129 (N_7129,N_5102,N_4737);
or U7130 (N_7130,N_5233,N_5424);
nor U7131 (N_7131,N_4441,N_6185);
or U7132 (N_7132,N_4059,N_3557);
or U7133 (N_7133,N_5839,N_4156);
nor U7134 (N_7134,N_3495,N_5443);
nand U7135 (N_7135,N_3700,N_4547);
nand U7136 (N_7136,N_5440,N_4226);
nand U7137 (N_7137,N_3969,N_4245);
xor U7138 (N_7138,N_4915,N_4215);
and U7139 (N_7139,N_5543,N_3714);
nor U7140 (N_7140,N_4341,N_5234);
and U7141 (N_7141,N_3850,N_3578);
xnor U7142 (N_7142,N_5224,N_5525);
nand U7143 (N_7143,N_3257,N_3444);
nand U7144 (N_7144,N_5212,N_5391);
and U7145 (N_7145,N_4611,N_3416);
nor U7146 (N_7146,N_5481,N_3822);
nand U7147 (N_7147,N_5316,N_3741);
nor U7148 (N_7148,N_3664,N_4034);
nor U7149 (N_7149,N_3394,N_5843);
nor U7150 (N_7150,N_4617,N_3751);
nor U7151 (N_7151,N_3766,N_3786);
nor U7152 (N_7152,N_3678,N_4849);
or U7153 (N_7153,N_4806,N_3807);
nor U7154 (N_7154,N_4122,N_4644);
or U7155 (N_7155,N_4131,N_4705);
nor U7156 (N_7156,N_3458,N_5995);
xnor U7157 (N_7157,N_4734,N_5322);
or U7158 (N_7158,N_5455,N_4219);
nand U7159 (N_7159,N_5930,N_4937);
xnor U7160 (N_7160,N_4000,N_3641);
and U7161 (N_7161,N_3933,N_6033);
xnor U7162 (N_7162,N_4197,N_3830);
xnor U7163 (N_7163,N_4313,N_5952);
or U7164 (N_7164,N_5594,N_3155);
xnor U7165 (N_7165,N_5694,N_3306);
nor U7166 (N_7166,N_5412,N_5257);
nor U7167 (N_7167,N_3438,N_5422);
nand U7168 (N_7168,N_5221,N_4440);
or U7169 (N_7169,N_5118,N_3809);
nor U7170 (N_7170,N_4933,N_4049);
and U7171 (N_7171,N_4754,N_5179);
nor U7172 (N_7172,N_5668,N_5854);
xnor U7173 (N_7173,N_4042,N_4369);
or U7174 (N_7174,N_4898,N_3409);
xnor U7175 (N_7175,N_4549,N_5035);
nor U7176 (N_7176,N_4086,N_4108);
nor U7177 (N_7177,N_5158,N_4887);
and U7178 (N_7178,N_5389,N_5433);
nand U7179 (N_7179,N_3919,N_4749);
and U7180 (N_7180,N_4733,N_4882);
nand U7181 (N_7181,N_5934,N_4799);
xnor U7182 (N_7182,N_3481,N_5673);
nor U7183 (N_7183,N_5245,N_4275);
and U7184 (N_7184,N_5847,N_5997);
and U7185 (N_7185,N_4683,N_5918);
or U7186 (N_7186,N_5230,N_3298);
and U7187 (N_7187,N_5463,N_3950);
or U7188 (N_7188,N_4006,N_4995);
and U7189 (N_7189,N_5477,N_5560);
nand U7190 (N_7190,N_4628,N_3915);
and U7191 (N_7191,N_4746,N_4692);
or U7192 (N_7192,N_5540,N_4116);
and U7193 (N_7193,N_4176,N_3288);
and U7194 (N_7194,N_4274,N_4419);
or U7195 (N_7195,N_3144,N_6030);
or U7196 (N_7196,N_6068,N_4769);
or U7197 (N_7197,N_5783,N_3351);
or U7198 (N_7198,N_4716,N_3858);
nand U7199 (N_7199,N_4358,N_3720);
nor U7200 (N_7200,N_3816,N_4516);
or U7201 (N_7201,N_4795,N_3440);
or U7202 (N_7202,N_3774,N_4711);
or U7203 (N_7203,N_3129,N_5830);
nor U7204 (N_7204,N_6241,N_3992);
nand U7205 (N_7205,N_3553,N_4373);
xnor U7206 (N_7206,N_4864,N_5779);
nor U7207 (N_7207,N_4112,N_3929);
nor U7208 (N_7208,N_3808,N_4105);
nor U7209 (N_7209,N_6115,N_3826);
and U7210 (N_7210,N_5841,N_3274);
nor U7211 (N_7211,N_5895,N_4273);
or U7212 (N_7212,N_4539,N_5529);
or U7213 (N_7213,N_4607,N_3825);
and U7214 (N_7214,N_4213,N_3722);
xor U7215 (N_7215,N_5253,N_4170);
or U7216 (N_7216,N_5246,N_3556);
xnor U7217 (N_7217,N_4221,N_3225);
and U7218 (N_7218,N_4334,N_4533);
and U7219 (N_7219,N_4954,N_4052);
and U7220 (N_7220,N_4881,N_5420);
nor U7221 (N_7221,N_5476,N_4521);
and U7222 (N_7222,N_5659,N_4380);
nand U7223 (N_7223,N_5911,N_3978);
xnor U7224 (N_7224,N_4751,N_5439);
and U7225 (N_7225,N_3180,N_5716);
nor U7226 (N_7226,N_4624,N_5262);
and U7227 (N_7227,N_5635,N_6239);
xnor U7228 (N_7228,N_4582,N_3884);
or U7229 (N_7229,N_4391,N_4342);
xor U7230 (N_7230,N_4030,N_3327);
nand U7231 (N_7231,N_4270,N_4298);
xnor U7232 (N_7232,N_5282,N_3903);
xor U7233 (N_7233,N_4829,N_6228);
and U7234 (N_7234,N_4659,N_3315);
and U7235 (N_7235,N_3181,N_5046);
and U7236 (N_7236,N_4136,N_6020);
nor U7237 (N_7237,N_5821,N_5516);
and U7238 (N_7238,N_5697,N_3268);
and U7239 (N_7239,N_4479,N_3510);
or U7240 (N_7240,N_4417,N_4785);
nor U7241 (N_7241,N_4148,N_4113);
xnor U7242 (N_7242,N_3645,N_3974);
or U7243 (N_7243,N_5903,N_4596);
nand U7244 (N_7244,N_3385,N_5055);
or U7245 (N_7245,N_5833,N_4255);
xnor U7246 (N_7246,N_4253,N_6096);
nand U7247 (N_7247,N_4492,N_6045);
or U7248 (N_7248,N_5614,N_5427);
nor U7249 (N_7249,N_5801,N_4654);
nand U7250 (N_7250,N_5162,N_3666);
nor U7251 (N_7251,N_4694,N_4827);
xor U7252 (N_7252,N_3493,N_4892);
nor U7253 (N_7253,N_3599,N_6021);
nand U7254 (N_7254,N_3284,N_5719);
xnor U7255 (N_7255,N_4686,N_5743);
nand U7256 (N_7256,N_3928,N_4186);
nand U7257 (N_7257,N_5814,N_5778);
nand U7258 (N_7258,N_3559,N_3164);
xor U7259 (N_7259,N_4284,N_4772);
or U7260 (N_7260,N_4188,N_4264);
or U7261 (N_7261,N_5597,N_6117);
nand U7262 (N_7262,N_4608,N_4135);
nor U7263 (N_7263,N_5180,N_4184);
nand U7264 (N_7264,N_4957,N_4102);
nand U7265 (N_7265,N_4835,N_4283);
nand U7266 (N_7266,N_5492,N_3253);
xnor U7267 (N_7267,N_5901,N_3610);
nor U7268 (N_7268,N_5593,N_4618);
nand U7269 (N_7269,N_4436,N_4266);
or U7270 (N_7270,N_3729,N_5963);
nor U7271 (N_7271,N_3183,N_5075);
or U7272 (N_7272,N_4977,N_3549);
nand U7273 (N_7273,N_3260,N_3552);
and U7274 (N_7274,N_6179,N_5829);
nor U7275 (N_7275,N_5914,N_3365);
nand U7276 (N_7276,N_5765,N_5699);
nor U7277 (N_7277,N_5196,N_3146);
nor U7278 (N_7278,N_6205,N_3607);
nand U7279 (N_7279,N_3775,N_4189);
and U7280 (N_7280,N_4347,N_5772);
or U7281 (N_7281,N_6104,N_5615);
nor U7282 (N_7282,N_4044,N_4787);
or U7283 (N_7283,N_6108,N_5344);
or U7284 (N_7284,N_5534,N_4394);
or U7285 (N_7285,N_4485,N_3872);
nor U7286 (N_7286,N_5692,N_6171);
xor U7287 (N_7287,N_5136,N_3907);
nor U7288 (N_7288,N_3382,N_3448);
and U7289 (N_7289,N_4838,N_5630);
xnor U7290 (N_7290,N_3545,N_3459);
nand U7291 (N_7291,N_5663,N_4535);
xor U7292 (N_7292,N_5028,N_5194);
and U7293 (N_7293,N_3840,N_5595);
nor U7294 (N_7294,N_5528,N_5308);
and U7295 (N_7295,N_4651,N_3479);
or U7296 (N_7296,N_3421,N_3468);
xor U7297 (N_7297,N_5203,N_5541);
and U7298 (N_7298,N_5338,N_5968);
nor U7299 (N_7299,N_4418,N_4744);
nand U7300 (N_7300,N_4016,N_5474);
or U7301 (N_7301,N_3264,N_3661);
nor U7302 (N_7302,N_4971,N_3617);
xnor U7303 (N_7303,N_6203,N_5494);
and U7304 (N_7304,N_3486,N_4464);
and U7305 (N_7305,N_5057,N_5059);
xnor U7306 (N_7306,N_3894,N_3269);
xor U7307 (N_7307,N_4243,N_4682);
xor U7308 (N_7308,N_3755,N_5332);
nor U7309 (N_7309,N_5737,N_4943);
and U7310 (N_7310,N_4205,N_5272);
and U7311 (N_7311,N_4709,N_5871);
xor U7312 (N_7312,N_5703,N_6126);
nor U7313 (N_7313,N_4710,N_4167);
nand U7314 (N_7314,N_5905,N_4236);
and U7315 (N_7315,N_5235,N_3142);
nand U7316 (N_7316,N_6001,N_4013);
xor U7317 (N_7317,N_3845,N_3540);
xor U7318 (N_7318,N_5287,N_5277);
nor U7319 (N_7319,N_5108,N_3680);
nor U7320 (N_7320,N_3708,N_3883);
and U7321 (N_7321,N_4207,N_5226);
and U7322 (N_7322,N_4355,N_5462);
nor U7323 (N_7323,N_5769,N_4852);
xnor U7324 (N_7324,N_5156,N_5352);
and U7325 (N_7325,N_5521,N_5369);
nand U7326 (N_7326,N_4315,N_3301);
nand U7327 (N_7327,N_5350,N_4575);
nand U7328 (N_7328,N_5897,N_5456);
nand U7329 (N_7329,N_3185,N_5020);
nand U7330 (N_7330,N_3613,N_5409);
nor U7331 (N_7331,N_3752,N_5686);
and U7332 (N_7332,N_4295,N_5121);
xor U7333 (N_7333,N_4774,N_6202);
nor U7334 (N_7334,N_3217,N_3412);
nand U7335 (N_7335,N_4160,N_5383);
xnor U7336 (N_7336,N_5292,N_3668);
nand U7337 (N_7337,N_6025,N_5084);
nor U7338 (N_7338,N_5732,N_5195);
xor U7339 (N_7339,N_4748,N_6219);
and U7340 (N_7340,N_3988,N_6081);
and U7341 (N_7341,N_5497,N_5503);
nor U7342 (N_7342,N_3466,N_4150);
and U7343 (N_7343,N_5684,N_4993);
or U7344 (N_7344,N_5215,N_3384);
xnor U7345 (N_7345,N_3963,N_5762);
nand U7346 (N_7346,N_4083,N_4990);
and U7347 (N_7347,N_4831,N_3954);
xnor U7348 (N_7348,N_4525,N_4531);
xor U7349 (N_7349,N_5966,N_4350);
xor U7350 (N_7350,N_4502,N_4494);
xor U7351 (N_7351,N_3793,N_5553);
nor U7352 (N_7352,N_6248,N_4600);
or U7353 (N_7353,N_3931,N_4939);
or U7354 (N_7354,N_4061,N_5310);
nor U7355 (N_7355,N_4175,N_4166);
nor U7356 (N_7356,N_5674,N_5931);
or U7357 (N_7357,N_5431,N_5027);
nor U7358 (N_7358,N_6120,N_3367);
or U7359 (N_7359,N_4861,N_6105);
nor U7360 (N_7360,N_4261,N_4847);
or U7361 (N_7361,N_4228,N_4209);
xor U7362 (N_7362,N_4169,N_6190);
and U7363 (N_7363,N_5330,N_3497);
nor U7364 (N_7364,N_4610,N_4178);
or U7365 (N_7365,N_5450,N_3743);
xor U7366 (N_7366,N_3727,N_3428);
and U7367 (N_7367,N_5297,N_5155);
xor U7368 (N_7368,N_5022,N_4739);
nand U7369 (N_7369,N_3321,N_3299);
xor U7370 (N_7370,N_3136,N_5334);
xnor U7371 (N_7371,N_5465,N_3152);
and U7372 (N_7372,N_5993,N_5689);
and U7373 (N_7373,N_5865,N_4474);
or U7374 (N_7374,N_3478,N_6212);
nand U7375 (N_7375,N_3173,N_3747);
xnor U7376 (N_7376,N_4612,N_5048);
nor U7377 (N_7377,N_4927,N_3687);
xor U7378 (N_7378,N_4950,N_4359);
or U7379 (N_7379,N_3671,N_5705);
nor U7380 (N_7380,N_3939,N_4378);
and U7381 (N_7381,N_3371,N_5133);
or U7382 (N_7382,N_5846,N_3841);
xor U7383 (N_7383,N_5138,N_3420);
xor U7384 (N_7384,N_4830,N_6223);
nand U7385 (N_7385,N_4819,N_5464);
xnor U7386 (N_7386,N_4137,N_3498);
nor U7387 (N_7387,N_3408,N_6101);
xnor U7388 (N_7388,N_3349,N_3838);
and U7389 (N_7389,N_4797,N_5242);
nand U7390 (N_7390,N_4517,N_5946);
nor U7391 (N_7391,N_3813,N_5337);
or U7392 (N_7392,N_3547,N_5739);
nand U7393 (N_7393,N_4925,N_6145);
nand U7394 (N_7394,N_3311,N_5429);
and U7395 (N_7395,N_4558,N_4997);
and U7396 (N_7396,N_4730,N_4029);
nand U7397 (N_7397,N_3655,N_4720);
nor U7398 (N_7398,N_4078,N_3609);
nand U7399 (N_7399,N_4230,N_4667);
xnor U7400 (N_7400,N_5052,N_6112);
nor U7401 (N_7401,N_6227,N_4675);
nand U7402 (N_7402,N_5880,N_5613);
nand U7403 (N_7403,N_3802,N_5907);
nor U7404 (N_7404,N_3593,N_5571);
nor U7405 (N_7405,N_4688,N_3435);
nand U7406 (N_7406,N_5530,N_6076);
and U7407 (N_7407,N_6124,N_3490);
or U7408 (N_7408,N_5329,N_5515);
or U7409 (N_7409,N_5380,N_3867);
nor U7410 (N_7410,N_4889,N_5127);
or U7411 (N_7411,N_4462,N_5790);
and U7412 (N_7412,N_3967,N_4410);
xor U7413 (N_7413,N_4679,N_4841);
and U7414 (N_7414,N_3591,N_5885);
nor U7415 (N_7415,N_6082,N_4290);
or U7416 (N_7416,N_4070,N_5753);
and U7417 (N_7417,N_5174,N_3244);
and U7418 (N_7418,N_4923,N_3487);
xnor U7419 (N_7419,N_5666,N_5153);
and U7420 (N_7420,N_4661,N_4483);
nand U7421 (N_7421,N_4154,N_5082);
nor U7422 (N_7422,N_5001,N_4722);
nand U7423 (N_7423,N_3586,N_3725);
nor U7424 (N_7424,N_5884,N_3326);
and U7425 (N_7425,N_5658,N_4921);
and U7426 (N_7426,N_4825,N_5074);
or U7427 (N_7427,N_4252,N_3209);
nor U7428 (N_7428,N_6113,N_3283);
xnor U7429 (N_7429,N_3660,N_5707);
nor U7430 (N_7430,N_6000,N_5266);
and U7431 (N_7431,N_6210,N_4728);
nor U7432 (N_7432,N_5704,N_3336);
nor U7433 (N_7433,N_4655,N_3611);
xor U7434 (N_7434,N_4758,N_6078);
xnor U7435 (N_7435,N_5624,N_3761);
nor U7436 (N_7436,N_3278,N_5363);
nand U7437 (N_7437,N_3814,N_4465);
xor U7438 (N_7438,N_4815,N_3196);
nand U7439 (N_7439,N_5665,N_6014);
nand U7440 (N_7440,N_4638,N_3489);
nand U7441 (N_7441,N_5572,N_6114);
and U7442 (N_7442,N_5480,N_3824);
xor U7443 (N_7443,N_4514,N_3794);
xor U7444 (N_7444,N_4592,N_3177);
and U7445 (N_7445,N_4348,N_3561);
or U7446 (N_7446,N_5675,N_4366);
and U7447 (N_7447,N_5239,N_4813);
nand U7448 (N_7448,N_4247,N_5671);
nor U7449 (N_7449,N_3904,N_5859);
or U7450 (N_7450,N_3986,N_4470);
and U7451 (N_7451,N_5114,N_5042);
or U7452 (N_7452,N_3231,N_3635);
nor U7453 (N_7453,N_4666,N_3584);
xnor U7454 (N_7454,N_3713,N_6197);
or U7455 (N_7455,N_5088,N_5218);
and U7456 (N_7456,N_5547,N_6049);
and U7457 (N_7457,N_3568,N_5730);
nor U7458 (N_7458,N_5971,N_3600);
and U7459 (N_7459,N_4755,N_4500);
nor U7460 (N_7460,N_4187,N_5949);
nor U7461 (N_7461,N_4195,N_3477);
nand U7462 (N_7462,N_3604,N_4196);
nor U7463 (N_7463,N_3577,N_4557);
nand U7464 (N_7464,N_5617,N_5005);
and U7465 (N_7465,N_4783,N_4293);
and U7466 (N_7466,N_3141,N_6098);
or U7467 (N_7467,N_5809,N_3972);
nand U7468 (N_7468,N_6166,N_4801);
nor U7469 (N_7469,N_6141,N_3710);
xor U7470 (N_7470,N_4292,N_3271);
and U7471 (N_7471,N_3868,N_4579);
or U7472 (N_7472,N_5942,N_5044);
or U7473 (N_7473,N_5989,N_4130);
or U7474 (N_7474,N_4278,N_5872);
nand U7475 (N_7475,N_6019,N_3832);
xnor U7476 (N_7476,N_3415,N_4145);
and U7477 (N_7477,N_5457,N_4510);
xor U7478 (N_7478,N_5470,N_3735);
or U7479 (N_7479,N_3534,N_5866);
nand U7480 (N_7480,N_5219,N_4816);
xnor U7481 (N_7481,N_3506,N_4318);
nor U7482 (N_7482,N_4103,N_3926);
or U7483 (N_7483,N_5861,N_5168);
and U7484 (N_7484,N_5124,N_5520);
xor U7485 (N_7485,N_4423,N_4961);
nor U7486 (N_7486,N_3853,N_5101);
and U7487 (N_7487,N_3352,N_3446);
nand U7488 (N_7488,N_4218,N_4151);
nand U7489 (N_7489,N_4578,N_3889);
and U7490 (N_7490,N_4777,N_5734);
and U7491 (N_7491,N_4035,N_5251);
xnor U7492 (N_7492,N_3922,N_4486);
or U7493 (N_7493,N_4963,N_3605);
nor U7494 (N_7494,N_5502,N_5711);
nor U7495 (N_7495,N_4609,N_5147);
xnor U7496 (N_7496,N_5567,N_3764);
or U7497 (N_7497,N_6224,N_4523);
and U7498 (N_7498,N_4724,N_5812);
and U7499 (N_7499,N_3254,N_3223);
xor U7500 (N_7500,N_4556,N_3402);
and U7501 (N_7501,N_6211,N_3266);
nor U7502 (N_7502,N_4912,N_4193);
nand U7503 (N_7503,N_3817,N_6170);
and U7504 (N_7504,N_4012,N_4540);
and U7505 (N_7505,N_5924,N_4256);
and U7506 (N_7506,N_4120,N_6132);
nand U7507 (N_7507,N_4842,N_4217);
nand U7508 (N_7508,N_6038,N_4511);
or U7509 (N_7509,N_5799,N_5134);
or U7510 (N_7510,N_3447,N_3717);
nor U7511 (N_7511,N_4595,N_5507);
nand U7512 (N_7512,N_3882,N_4884);
xnor U7513 (N_7513,N_4368,N_4498);
xnor U7514 (N_7514,N_3772,N_4627);
or U7515 (N_7515,N_4141,N_3649);
nand U7516 (N_7516,N_5414,N_5148);
nand U7517 (N_7517,N_4403,N_3874);
or U7518 (N_7518,N_4524,N_4848);
xor U7519 (N_7519,N_5638,N_6018);
nor U7520 (N_7520,N_5152,N_3985);
or U7521 (N_7521,N_4455,N_5252);
or U7522 (N_7522,N_5548,N_5979);
xnor U7523 (N_7523,N_5446,N_3548);
xnor U7524 (N_7524,N_3646,N_4850);
and U7525 (N_7525,N_4684,N_5015);
and U7526 (N_7526,N_5295,N_5321);
nor U7527 (N_7527,N_5407,N_3430);
and U7528 (N_7528,N_6220,N_3994);
nor U7529 (N_7529,N_5392,N_3843);
nand U7530 (N_7530,N_4056,N_6206);
xnor U7531 (N_7531,N_6147,N_4563);
and U7532 (N_7532,N_6172,N_5274);
or U7533 (N_7533,N_5359,N_3911);
nand U7534 (N_7534,N_4994,N_4239);
xnor U7535 (N_7535,N_4127,N_4559);
xnor U7536 (N_7536,N_4703,N_5587);
or U7537 (N_7537,N_6148,N_6229);
or U7538 (N_7538,N_3410,N_3226);
and U7539 (N_7539,N_5306,N_4458);
nand U7540 (N_7540,N_3582,N_3536);
nand U7541 (N_7541,N_5798,N_3712);
and U7542 (N_7542,N_5536,N_5278);
nor U7543 (N_7543,N_5225,N_3454);
xnor U7544 (N_7544,N_4330,N_5879);
nor U7545 (N_7545,N_4650,N_5265);
nor U7546 (N_7546,N_6065,N_5569);
or U7547 (N_7547,N_3453,N_3857);
and U7548 (N_7548,N_4420,N_4701);
or U7549 (N_7549,N_4074,N_6121);
xnor U7550 (N_7550,N_3862,N_4161);
and U7551 (N_7551,N_3724,N_3285);
nand U7552 (N_7552,N_5797,N_5815);
nand U7553 (N_7553,N_5896,N_5542);
or U7554 (N_7554,N_3945,N_4208);
xnor U7555 (N_7555,N_3756,N_4392);
nand U7556 (N_7556,N_5526,N_3897);
nand U7557 (N_7557,N_6051,N_5104);
nand U7558 (N_7558,N_5031,N_5068);
nand U7559 (N_7559,N_3597,N_3133);
nand U7560 (N_7560,N_4542,N_3232);
and U7561 (N_7561,N_4390,N_3357);
and U7562 (N_7562,N_5751,N_5709);
or U7563 (N_7563,N_4873,N_4041);
or U7564 (N_7564,N_3207,N_3702);
xnor U7565 (N_7565,N_5393,N_4337);
xor U7566 (N_7566,N_5264,N_3731);
nand U7567 (N_7567,N_3126,N_6047);
and U7568 (N_7568,N_4712,N_3723);
or U7569 (N_7569,N_4081,N_3328);
or U7570 (N_7570,N_4152,N_3143);
or U7571 (N_7571,N_4904,N_3179);
or U7572 (N_7572,N_4555,N_3535);
or U7573 (N_7573,N_5943,N_4091);
and U7574 (N_7574,N_5996,N_3234);
and U7575 (N_7575,N_3810,N_3500);
or U7576 (N_7576,N_6044,N_4657);
and U7577 (N_7577,N_3912,N_3452);
xor U7578 (N_7578,N_4225,N_6009);
or U7579 (N_7579,N_3937,N_3531);
nand U7580 (N_7580,N_3742,N_3396);
or U7581 (N_7581,N_5891,N_4097);
nand U7582 (N_7582,N_4800,N_3544);
xnor U7583 (N_7583,N_5592,N_5793);
or U7584 (N_7584,N_3442,N_5794);
nor U7585 (N_7585,N_5454,N_4958);
xnor U7586 (N_7586,N_5367,N_5804);
or U7587 (N_7587,N_6156,N_3507);
nor U7588 (N_7588,N_3958,N_5299);
nand U7589 (N_7589,N_5796,N_4917);
xor U7590 (N_7590,N_3528,N_4652);
and U7591 (N_7591,N_4568,N_4911);
or U7592 (N_7592,N_5061,N_3663);
nor U7593 (N_7593,N_6097,N_5347);
nand U7594 (N_7594,N_3204,N_3247);
or U7595 (N_7595,N_5766,N_3693);
and U7596 (N_7596,N_4087,N_6177);
or U7597 (N_7597,N_4249,N_3688);
nand U7598 (N_7598,N_4693,N_6235);
xor U7599 (N_7599,N_5806,N_5394);
xnor U7600 (N_7600,N_5679,N_5978);
or U7601 (N_7601,N_6244,N_6116);
or U7602 (N_7602,N_4691,N_5317);
xor U7603 (N_7603,N_5965,N_5348);
nor U7604 (N_7604,N_3901,N_5080);
nand U7605 (N_7605,N_5874,N_4938);
or U7606 (N_7606,N_4839,N_3526);
or U7607 (N_7607,N_4643,N_5967);
nor U7608 (N_7608,N_5328,N_4700);
xor U7609 (N_7609,N_3624,N_4325);
and U7610 (N_7610,N_5561,N_4672);
and U7611 (N_7611,N_4489,N_4591);
nand U7612 (N_7612,N_3657,N_5418);
nor U7613 (N_7613,N_3639,N_3562);
xnor U7614 (N_7614,N_3229,N_3353);
or U7615 (N_7615,N_3864,N_3222);
nand U7616 (N_7616,N_5030,N_3861);
xnor U7617 (N_7617,N_5818,N_5223);
nor U7618 (N_7618,N_5917,N_3423);
nor U7619 (N_7619,N_3361,N_3521);
nor U7620 (N_7620,N_3165,N_3441);
xor U7621 (N_7621,N_3914,N_6184);
nor U7622 (N_7622,N_5206,N_6188);
and U7623 (N_7623,N_4681,N_6062);
nand U7624 (N_7624,N_3256,N_6240);
nor U7625 (N_7625,N_6245,N_5205);
or U7626 (N_7626,N_4312,N_6050);
and U7627 (N_7627,N_4118,N_4265);
nor U7628 (N_7628,N_3706,N_4409);
xor U7629 (N_7629,N_6149,N_5926);
nand U7630 (N_7630,N_4756,N_4367);
nor U7631 (N_7631,N_3812,N_5361);
nand U7632 (N_7632,N_5537,N_5296);
nand U7633 (N_7633,N_4570,N_5629);
nor U7634 (N_7634,N_4928,N_4653);
nand U7635 (N_7635,N_3491,N_3132);
nand U7636 (N_7636,N_5432,N_4096);
nor U7637 (N_7637,N_3815,N_4235);
xor U7638 (N_7638,N_3638,N_5004);
xor U7639 (N_7639,N_4340,N_5384);
nor U7640 (N_7640,N_3443,N_5184);
and U7641 (N_7641,N_5827,N_3739);
and U7642 (N_7642,N_5053,N_3876);
nand U7643 (N_7643,N_3272,N_3135);
nand U7644 (N_7644,N_4395,N_6143);
nand U7645 (N_7645,N_4336,N_4079);
nand U7646 (N_7646,N_3241,N_4548);
or U7647 (N_7647,N_5419,N_4583);
nand U7648 (N_7648,N_3899,N_5189);
and U7649 (N_7649,N_6174,N_5256);
xnor U7650 (N_7650,N_5117,N_5469);
or U7651 (N_7651,N_4664,N_5021);
xor U7652 (N_7652,N_5500,N_3924);
nand U7653 (N_7653,N_4090,N_4222);
and U7654 (N_7654,N_5855,N_5479);
and U7655 (N_7655,N_4891,N_4168);
nand U7656 (N_7656,N_5672,N_3145);
nand U7657 (N_7657,N_5047,N_4897);
and U7658 (N_7658,N_6164,N_5781);
nor U7659 (N_7659,N_4715,N_5327);
nor U7660 (N_7660,N_4987,N_4953);
and U7661 (N_7661,N_3249,N_5095);
nand U7662 (N_7662,N_3240,N_4906);
and U7663 (N_7663,N_5991,N_4499);
nor U7664 (N_7664,N_3359,N_5307);
nor U7665 (N_7665,N_5664,N_4433);
nand U7666 (N_7666,N_3156,N_3909);
and U7667 (N_7667,N_4060,N_3925);
nand U7668 (N_7668,N_5066,N_5130);
and U7669 (N_7669,N_3603,N_5301);
and U7670 (N_7670,N_3691,N_3643);
and U7671 (N_7671,N_4967,N_3791);
or U7672 (N_7672,N_4314,N_6128);
nor U7673 (N_7673,N_5346,N_3309);
and U7674 (N_7674,N_4448,N_5718);
xor U7675 (N_7675,N_5508,N_5975);
nor U7676 (N_7676,N_5519,N_4260);
or U7677 (N_7677,N_3213,N_3893);
and U7678 (N_7678,N_3957,N_4714);
nand U7679 (N_7679,N_5504,N_4569);
or U7680 (N_7680,N_5925,N_6071);
and U7681 (N_7681,N_3404,N_6008);
and U7682 (N_7682,N_5210,N_6180);
nand U7683 (N_7683,N_3736,N_4302);
and U7684 (N_7684,N_5472,N_6144);
nor U7685 (N_7685,N_5036,N_6214);
and U7686 (N_7686,N_5487,N_3916);
or U7687 (N_7687,N_4804,N_3587);
and U7688 (N_7688,N_5767,N_5120);
nand U7689 (N_7689,N_5581,N_4594);
or U7690 (N_7690,N_4883,N_5415);
nand U7691 (N_7691,N_5198,N_5313);
nand U7692 (N_7692,N_3779,N_5601);
xor U7693 (N_7693,N_5161,N_5877);
xnor U7694 (N_7694,N_3905,N_3433);
xnor U7695 (N_7695,N_3913,N_5552);
nand U7696 (N_7696,N_3715,N_5255);
and U7697 (N_7697,N_6238,N_4415);
nor U7698 (N_7698,N_5231,N_4493);
xor U7699 (N_7699,N_3690,N_3746);
xnor U7700 (N_7700,N_4622,N_5789);
and U7701 (N_7701,N_3221,N_4133);
and U7702 (N_7702,N_5410,N_4477);
xor U7703 (N_7703,N_6005,N_5590);
nand U7704 (N_7704,N_6034,N_4232);
or U7705 (N_7705,N_3364,N_5582);
or U7706 (N_7706,N_4328,N_4406);
and U7707 (N_7707,N_3436,N_5188);
or U7708 (N_7708,N_4991,N_5811);
nand U7709 (N_7709,N_4719,N_5428);
nor U7710 (N_7710,N_5378,N_5944);
or U7711 (N_7711,N_4132,N_4640);
nand U7712 (N_7712,N_5305,N_5923);
nand U7713 (N_7713,N_4288,N_4931);
nand U7714 (N_7714,N_3377,N_4139);
or U7715 (N_7715,N_3694,N_4512);
nor U7716 (N_7716,N_4676,N_6152);
xor U7717 (N_7717,N_3980,N_5816);
xor U7718 (N_7718,N_4323,N_5845);
nor U7719 (N_7719,N_4546,N_4509);
or U7720 (N_7720,N_5916,N_3672);
and U7721 (N_7721,N_4964,N_4796);
and U7722 (N_7722,N_4814,N_5645);
xnor U7723 (N_7723,N_3414,N_5285);
nand U7724 (N_7724,N_3614,N_4316);
xnor U7725 (N_7725,N_4468,N_6123);
or U7726 (N_7726,N_5249,N_5825);
or U7727 (N_7727,N_3792,N_4388);
nor U7728 (N_7728,N_5445,N_3380);
nand U7729 (N_7729,N_3469,N_4633);
and U7730 (N_7730,N_3167,N_3689);
or U7731 (N_7731,N_4649,N_4258);
nor U7732 (N_7732,N_5754,N_4867);
nor U7733 (N_7733,N_6151,N_3701);
and U7734 (N_7734,N_5643,N_5687);
and U7735 (N_7735,N_4586,N_6016);
and U7736 (N_7736,N_3944,N_6165);
nand U7737 (N_7737,N_3203,N_3342);
nor U7738 (N_7738,N_4453,N_5852);
and U7739 (N_7739,N_4833,N_6055);
and U7740 (N_7740,N_4383,N_5193);
or U7741 (N_7741,N_4836,N_6226);
nor U7742 (N_7742,N_5862,N_4036);
nand U7743 (N_7743,N_5768,N_4182);
xor U7744 (N_7744,N_4171,N_6107);
nor U7745 (N_7745,N_3422,N_3530);
nor U7746 (N_7746,N_3212,N_3482);
xor U7747 (N_7747,N_4580,N_5800);
xnor U7748 (N_7748,N_5090,N_4623);
and U7749 (N_7749,N_5003,N_5688);
and U7750 (N_7750,N_3633,N_4573);
or U7751 (N_7751,N_4444,N_3543);
xor U7752 (N_7752,N_3354,N_4752);
or U7753 (N_7753,N_3379,N_3330);
xnor U7754 (N_7754,N_5892,N_4387);
nand U7755 (N_7755,N_3805,N_4211);
xor U7756 (N_7756,N_5144,N_4126);
and U7757 (N_7757,N_4063,N_3966);
nor U7758 (N_7758,N_4708,N_5950);
nor U7759 (N_7759,N_4227,N_4598);
and U7760 (N_7760,N_3170,N_3970);
or U7761 (N_7761,N_4941,N_4634);
nand U7762 (N_7762,N_3621,N_4027);
or U7763 (N_7763,N_5640,N_3273);
xnor U7764 (N_7764,N_3401,N_4914);
nor U7765 (N_7765,N_4421,N_5576);
or U7766 (N_7766,N_3270,N_4174);
or U7767 (N_7767,N_4202,N_4203);
or U7768 (N_7768,N_3748,N_4428);
and U7769 (N_7769,N_3537,N_5400);
and U7770 (N_7770,N_3236,N_4590);
or U7771 (N_7771,N_3291,N_6089);
nand U7772 (N_7772,N_3616,N_3842);
or U7773 (N_7773,N_5598,N_4017);
and U7774 (N_7774,N_3837,N_4069);
xor U7775 (N_7775,N_3182,N_3228);
nand U7776 (N_7776,N_5273,N_4449);
or U7777 (N_7777,N_3682,N_5064);
or U7778 (N_7778,N_5619,N_4353);
nand U7779 (N_7779,N_5371,N_4846);
nand U7780 (N_7780,N_6237,N_5728);
or U7781 (N_7781,N_6204,N_3726);
xnor U7782 (N_7782,N_3533,N_3432);
nor U7783 (N_7783,N_5559,N_4729);
xor U7784 (N_7784,N_4206,N_3392);
or U7785 (N_7785,N_4520,N_3930);
or U7786 (N_7786,N_5105,N_3312);
nand U7787 (N_7787,N_5820,N_5238);
or U7788 (N_7788,N_3959,N_3594);
and U7789 (N_7789,N_6131,N_4619);
nor U7790 (N_7790,N_5373,N_6140);
and U7791 (N_7791,N_4459,N_3773);
or U7792 (N_7792,N_4890,N_4413);
nor U7793 (N_7793,N_5014,N_3318);
or U7794 (N_7794,N_5490,N_4271);
and U7795 (N_7795,N_4826,N_3429);
xnor U7796 (N_7796,N_3596,N_5208);
and U7797 (N_7797,N_5726,N_4011);
and U7798 (N_7798,N_4907,N_3699);
xnor U7799 (N_7799,N_5655,N_3744);
xor U7800 (N_7800,N_3383,N_3960);
xor U7801 (N_7801,N_3261,N_5318);
nand U7802 (N_7802,N_4023,N_4040);
nor U7803 (N_7803,N_4478,N_5702);
xor U7804 (N_7804,N_5139,N_4900);
nor U7805 (N_7805,N_4460,N_4375);
nand U7806 (N_7806,N_4432,N_4504);
xnor U7807 (N_7807,N_4639,N_3527);
and U7808 (N_7808,N_5388,N_4129);
xnor U7809 (N_7809,N_5657,N_3492);
nor U7810 (N_7810,N_5676,N_5366);
or U7811 (N_7811,N_4054,N_4946);
or U7812 (N_7812,N_5721,N_6049);
xnor U7813 (N_7813,N_4881,N_4284);
xor U7814 (N_7814,N_4345,N_5477);
xnor U7815 (N_7815,N_5513,N_4374);
or U7816 (N_7816,N_4024,N_3860);
nor U7817 (N_7817,N_4012,N_5707);
nand U7818 (N_7818,N_3881,N_3604);
nor U7819 (N_7819,N_4133,N_3498);
xor U7820 (N_7820,N_6097,N_4362);
and U7821 (N_7821,N_5305,N_5588);
and U7822 (N_7822,N_3650,N_3296);
and U7823 (N_7823,N_3228,N_4729);
nor U7824 (N_7824,N_3583,N_4485);
and U7825 (N_7825,N_4295,N_5474);
or U7826 (N_7826,N_5827,N_5719);
xnor U7827 (N_7827,N_5513,N_3799);
nor U7828 (N_7828,N_3615,N_3771);
or U7829 (N_7829,N_3286,N_3387);
xnor U7830 (N_7830,N_3589,N_5311);
xnor U7831 (N_7831,N_5486,N_5260);
nor U7832 (N_7832,N_3884,N_4854);
nor U7833 (N_7833,N_4909,N_3258);
and U7834 (N_7834,N_5894,N_6003);
nor U7835 (N_7835,N_4152,N_3512);
nor U7836 (N_7836,N_4650,N_3401);
nand U7837 (N_7837,N_4173,N_4779);
nor U7838 (N_7838,N_4431,N_4241);
xnor U7839 (N_7839,N_4639,N_5755);
and U7840 (N_7840,N_3445,N_5018);
and U7841 (N_7841,N_5619,N_4080);
or U7842 (N_7842,N_4757,N_4207);
nor U7843 (N_7843,N_3704,N_3685);
nor U7844 (N_7844,N_4866,N_5199);
or U7845 (N_7845,N_4820,N_4751);
and U7846 (N_7846,N_6186,N_5034);
nor U7847 (N_7847,N_3754,N_5027);
nand U7848 (N_7848,N_5842,N_3176);
nand U7849 (N_7849,N_5554,N_5941);
nand U7850 (N_7850,N_6146,N_3922);
and U7851 (N_7851,N_3481,N_5816);
nor U7852 (N_7852,N_5914,N_4546);
and U7853 (N_7853,N_4638,N_3617);
xor U7854 (N_7854,N_3615,N_4059);
nand U7855 (N_7855,N_3556,N_3595);
nor U7856 (N_7856,N_4285,N_3773);
nor U7857 (N_7857,N_3835,N_4422);
or U7858 (N_7858,N_5803,N_5000);
xor U7859 (N_7859,N_5185,N_3153);
nand U7860 (N_7860,N_3524,N_4326);
nand U7861 (N_7861,N_4843,N_3545);
and U7862 (N_7862,N_4591,N_3446);
or U7863 (N_7863,N_3620,N_5917);
nand U7864 (N_7864,N_3832,N_3616);
xnor U7865 (N_7865,N_4383,N_3409);
nor U7866 (N_7866,N_6242,N_3832);
nor U7867 (N_7867,N_4504,N_5086);
and U7868 (N_7868,N_5658,N_4275);
and U7869 (N_7869,N_4503,N_5648);
and U7870 (N_7870,N_3144,N_5259);
nand U7871 (N_7871,N_5455,N_5448);
nand U7872 (N_7872,N_4211,N_4357);
nor U7873 (N_7873,N_3969,N_5305);
or U7874 (N_7874,N_5044,N_3485);
nor U7875 (N_7875,N_6107,N_6144);
or U7876 (N_7876,N_5523,N_5866);
or U7877 (N_7877,N_5333,N_3180);
nand U7878 (N_7878,N_5212,N_4161);
xor U7879 (N_7879,N_4219,N_5901);
nor U7880 (N_7880,N_5677,N_4614);
nand U7881 (N_7881,N_4111,N_4527);
and U7882 (N_7882,N_4064,N_3373);
nand U7883 (N_7883,N_3318,N_5399);
nand U7884 (N_7884,N_4847,N_4170);
nor U7885 (N_7885,N_3602,N_5633);
nor U7886 (N_7886,N_4818,N_4724);
and U7887 (N_7887,N_3381,N_4003);
nand U7888 (N_7888,N_3943,N_3568);
xnor U7889 (N_7889,N_4252,N_5067);
and U7890 (N_7890,N_4092,N_3177);
nand U7891 (N_7891,N_3833,N_4548);
or U7892 (N_7892,N_5355,N_4528);
xnor U7893 (N_7893,N_3259,N_4004);
nand U7894 (N_7894,N_3884,N_4841);
xnor U7895 (N_7895,N_5329,N_3605);
xnor U7896 (N_7896,N_4161,N_3551);
or U7897 (N_7897,N_5704,N_5609);
nor U7898 (N_7898,N_5278,N_4806);
nand U7899 (N_7899,N_5314,N_4657);
xor U7900 (N_7900,N_5371,N_4785);
nand U7901 (N_7901,N_4454,N_4641);
or U7902 (N_7902,N_5929,N_4169);
xnor U7903 (N_7903,N_5186,N_5309);
nor U7904 (N_7904,N_5623,N_4596);
nor U7905 (N_7905,N_4593,N_4577);
xnor U7906 (N_7906,N_4268,N_6238);
xor U7907 (N_7907,N_4521,N_5316);
and U7908 (N_7908,N_6043,N_3808);
and U7909 (N_7909,N_3561,N_4124);
nor U7910 (N_7910,N_5386,N_3717);
or U7911 (N_7911,N_5052,N_3700);
nor U7912 (N_7912,N_4343,N_3545);
nor U7913 (N_7913,N_4930,N_4234);
or U7914 (N_7914,N_5019,N_4111);
nand U7915 (N_7915,N_4894,N_3486);
nand U7916 (N_7916,N_3584,N_3896);
nand U7917 (N_7917,N_3705,N_4611);
nor U7918 (N_7918,N_3667,N_4201);
nor U7919 (N_7919,N_3409,N_3883);
and U7920 (N_7920,N_5396,N_6071);
nand U7921 (N_7921,N_6078,N_4881);
nand U7922 (N_7922,N_4684,N_5500);
nor U7923 (N_7923,N_4784,N_5141);
or U7924 (N_7924,N_5123,N_5928);
nor U7925 (N_7925,N_3523,N_6110);
nor U7926 (N_7926,N_4080,N_4342);
or U7927 (N_7927,N_4711,N_3811);
and U7928 (N_7928,N_5378,N_5595);
and U7929 (N_7929,N_5703,N_3708);
nor U7930 (N_7930,N_5219,N_3936);
nand U7931 (N_7931,N_4815,N_6238);
nor U7932 (N_7932,N_3591,N_3615);
nand U7933 (N_7933,N_6036,N_4975);
or U7934 (N_7934,N_3779,N_4566);
nor U7935 (N_7935,N_3248,N_5896);
nand U7936 (N_7936,N_3459,N_4675);
nor U7937 (N_7937,N_5129,N_4437);
nor U7938 (N_7938,N_4070,N_3898);
nand U7939 (N_7939,N_5352,N_3729);
xor U7940 (N_7940,N_5838,N_4880);
nand U7941 (N_7941,N_5450,N_3676);
nor U7942 (N_7942,N_4841,N_5697);
nor U7943 (N_7943,N_4426,N_3426);
xnor U7944 (N_7944,N_4462,N_3320);
nor U7945 (N_7945,N_4288,N_5581);
nand U7946 (N_7946,N_4112,N_5203);
xnor U7947 (N_7947,N_4410,N_3715);
or U7948 (N_7948,N_4590,N_5405);
nand U7949 (N_7949,N_5398,N_4386);
nand U7950 (N_7950,N_6148,N_4936);
or U7951 (N_7951,N_5140,N_5436);
nand U7952 (N_7952,N_4739,N_6205);
or U7953 (N_7953,N_4608,N_3174);
xnor U7954 (N_7954,N_5344,N_5291);
nand U7955 (N_7955,N_3250,N_4072);
or U7956 (N_7956,N_6135,N_5750);
xor U7957 (N_7957,N_4585,N_5157);
nor U7958 (N_7958,N_5009,N_5200);
nand U7959 (N_7959,N_3742,N_3593);
nand U7960 (N_7960,N_3160,N_4534);
nand U7961 (N_7961,N_5467,N_4198);
xnor U7962 (N_7962,N_6238,N_3887);
nor U7963 (N_7963,N_5407,N_4322);
or U7964 (N_7964,N_3265,N_3175);
and U7965 (N_7965,N_3969,N_5773);
nand U7966 (N_7966,N_3488,N_3659);
or U7967 (N_7967,N_4087,N_5628);
or U7968 (N_7968,N_3679,N_4470);
nor U7969 (N_7969,N_4702,N_4617);
nand U7970 (N_7970,N_3869,N_4350);
nand U7971 (N_7971,N_4080,N_5159);
xnor U7972 (N_7972,N_3653,N_5392);
nand U7973 (N_7973,N_4140,N_5635);
nor U7974 (N_7974,N_5696,N_4478);
nor U7975 (N_7975,N_3313,N_6084);
xor U7976 (N_7976,N_5176,N_4425);
nand U7977 (N_7977,N_5466,N_3942);
and U7978 (N_7978,N_5624,N_6190);
nor U7979 (N_7979,N_5603,N_3721);
or U7980 (N_7980,N_4479,N_5259);
or U7981 (N_7981,N_4541,N_5838);
and U7982 (N_7982,N_5815,N_5141);
xnor U7983 (N_7983,N_5616,N_6055);
xor U7984 (N_7984,N_4493,N_5425);
or U7985 (N_7985,N_3246,N_5240);
nand U7986 (N_7986,N_3506,N_5449);
nand U7987 (N_7987,N_6034,N_4056);
and U7988 (N_7988,N_3522,N_5869);
or U7989 (N_7989,N_5588,N_5825);
and U7990 (N_7990,N_3624,N_4914);
or U7991 (N_7991,N_4902,N_5015);
or U7992 (N_7992,N_5977,N_5445);
xor U7993 (N_7993,N_3944,N_5193);
nor U7994 (N_7994,N_4925,N_3128);
xor U7995 (N_7995,N_5467,N_3497);
and U7996 (N_7996,N_5757,N_3454);
xor U7997 (N_7997,N_3627,N_5039);
nor U7998 (N_7998,N_5713,N_5335);
or U7999 (N_7999,N_4873,N_5661);
or U8000 (N_8000,N_3135,N_3617);
and U8001 (N_8001,N_3719,N_3470);
or U8002 (N_8002,N_6048,N_4493);
or U8003 (N_8003,N_3133,N_4509);
xor U8004 (N_8004,N_5609,N_3392);
xor U8005 (N_8005,N_4191,N_4103);
or U8006 (N_8006,N_4689,N_5517);
nor U8007 (N_8007,N_5404,N_5673);
nor U8008 (N_8008,N_6221,N_6170);
nor U8009 (N_8009,N_3730,N_5741);
and U8010 (N_8010,N_3955,N_5645);
or U8011 (N_8011,N_4596,N_5324);
and U8012 (N_8012,N_3998,N_5187);
and U8013 (N_8013,N_4921,N_3219);
nor U8014 (N_8014,N_5199,N_4664);
nand U8015 (N_8015,N_3419,N_4163);
nand U8016 (N_8016,N_6136,N_4992);
nor U8017 (N_8017,N_4970,N_3487);
xor U8018 (N_8018,N_5515,N_4158);
or U8019 (N_8019,N_5225,N_4821);
nor U8020 (N_8020,N_4190,N_5045);
nand U8021 (N_8021,N_4140,N_3659);
nor U8022 (N_8022,N_3662,N_5732);
nand U8023 (N_8023,N_5028,N_4022);
xor U8024 (N_8024,N_5180,N_3293);
and U8025 (N_8025,N_5196,N_4966);
or U8026 (N_8026,N_5038,N_5896);
xnor U8027 (N_8027,N_4870,N_3748);
or U8028 (N_8028,N_4053,N_3215);
nand U8029 (N_8029,N_5241,N_6062);
nand U8030 (N_8030,N_3902,N_3759);
xor U8031 (N_8031,N_5186,N_5206);
nor U8032 (N_8032,N_3306,N_5404);
nor U8033 (N_8033,N_4828,N_4191);
or U8034 (N_8034,N_5481,N_5553);
and U8035 (N_8035,N_5295,N_3192);
and U8036 (N_8036,N_4519,N_3440);
or U8037 (N_8037,N_5807,N_5177);
and U8038 (N_8038,N_3378,N_3777);
or U8039 (N_8039,N_5378,N_3452);
xor U8040 (N_8040,N_5550,N_4346);
nor U8041 (N_8041,N_4861,N_3497);
nand U8042 (N_8042,N_3405,N_4609);
and U8043 (N_8043,N_4707,N_4684);
nand U8044 (N_8044,N_5625,N_3629);
or U8045 (N_8045,N_3816,N_6238);
nor U8046 (N_8046,N_3212,N_4516);
and U8047 (N_8047,N_3567,N_3294);
xor U8048 (N_8048,N_5890,N_6184);
nor U8049 (N_8049,N_5420,N_4555);
nor U8050 (N_8050,N_6088,N_3609);
or U8051 (N_8051,N_4913,N_4999);
or U8052 (N_8052,N_3722,N_5979);
or U8053 (N_8053,N_3320,N_5132);
nand U8054 (N_8054,N_4588,N_4613);
and U8055 (N_8055,N_5620,N_3921);
xor U8056 (N_8056,N_4898,N_5907);
and U8057 (N_8057,N_3448,N_3753);
nand U8058 (N_8058,N_4400,N_4788);
or U8059 (N_8059,N_3634,N_4772);
nor U8060 (N_8060,N_3876,N_3964);
nand U8061 (N_8061,N_4379,N_4753);
xnor U8062 (N_8062,N_4271,N_3620);
and U8063 (N_8063,N_4846,N_3640);
nand U8064 (N_8064,N_3469,N_3326);
nand U8065 (N_8065,N_5711,N_5978);
and U8066 (N_8066,N_4897,N_5968);
nor U8067 (N_8067,N_3195,N_4779);
xnor U8068 (N_8068,N_4813,N_5149);
nor U8069 (N_8069,N_5689,N_3300);
or U8070 (N_8070,N_3473,N_3625);
and U8071 (N_8071,N_5038,N_6175);
nor U8072 (N_8072,N_3947,N_5638);
xor U8073 (N_8073,N_5608,N_5378);
nor U8074 (N_8074,N_3533,N_4173);
xnor U8075 (N_8075,N_4454,N_3917);
nand U8076 (N_8076,N_5422,N_5661);
nor U8077 (N_8077,N_3450,N_3663);
nand U8078 (N_8078,N_3933,N_3952);
nor U8079 (N_8079,N_3768,N_4253);
nand U8080 (N_8080,N_4317,N_5577);
or U8081 (N_8081,N_4299,N_3132);
or U8082 (N_8082,N_5483,N_3678);
and U8083 (N_8083,N_3856,N_5142);
or U8084 (N_8084,N_3683,N_3654);
xor U8085 (N_8085,N_4127,N_6093);
and U8086 (N_8086,N_6110,N_3229);
xnor U8087 (N_8087,N_3448,N_5632);
and U8088 (N_8088,N_4816,N_5231);
nand U8089 (N_8089,N_6175,N_4447);
xnor U8090 (N_8090,N_3826,N_3293);
and U8091 (N_8091,N_3437,N_5376);
nand U8092 (N_8092,N_3984,N_5726);
xnor U8093 (N_8093,N_5814,N_5030);
nand U8094 (N_8094,N_5303,N_3992);
and U8095 (N_8095,N_3896,N_4400);
or U8096 (N_8096,N_5411,N_5129);
nor U8097 (N_8097,N_4704,N_4174);
xnor U8098 (N_8098,N_4842,N_5125);
nand U8099 (N_8099,N_4894,N_6198);
nand U8100 (N_8100,N_3339,N_4001);
xor U8101 (N_8101,N_3472,N_3425);
nor U8102 (N_8102,N_5764,N_3509);
or U8103 (N_8103,N_4347,N_3348);
or U8104 (N_8104,N_4579,N_4539);
xor U8105 (N_8105,N_3576,N_5053);
nand U8106 (N_8106,N_5924,N_6021);
and U8107 (N_8107,N_3285,N_6111);
and U8108 (N_8108,N_3462,N_3303);
xor U8109 (N_8109,N_3289,N_6049);
and U8110 (N_8110,N_3835,N_3379);
nand U8111 (N_8111,N_5894,N_6082);
xor U8112 (N_8112,N_4442,N_4650);
nand U8113 (N_8113,N_5320,N_5590);
nand U8114 (N_8114,N_5129,N_4462);
nand U8115 (N_8115,N_3431,N_3362);
nor U8116 (N_8116,N_3588,N_5131);
and U8117 (N_8117,N_3265,N_3761);
and U8118 (N_8118,N_3260,N_4548);
and U8119 (N_8119,N_3634,N_3896);
nor U8120 (N_8120,N_3211,N_4994);
nand U8121 (N_8121,N_5595,N_3177);
nor U8122 (N_8122,N_5732,N_3661);
xor U8123 (N_8123,N_5275,N_6151);
nand U8124 (N_8124,N_3128,N_4283);
nand U8125 (N_8125,N_5278,N_6196);
or U8126 (N_8126,N_5845,N_5622);
or U8127 (N_8127,N_4096,N_5250);
or U8128 (N_8128,N_3865,N_4108);
xnor U8129 (N_8129,N_3921,N_3588);
xor U8130 (N_8130,N_4785,N_5012);
nor U8131 (N_8131,N_3955,N_4457);
and U8132 (N_8132,N_5523,N_5039);
nor U8133 (N_8133,N_4467,N_4000);
or U8134 (N_8134,N_5548,N_4743);
nand U8135 (N_8135,N_3979,N_5493);
nor U8136 (N_8136,N_3131,N_6197);
and U8137 (N_8137,N_5961,N_3829);
or U8138 (N_8138,N_4481,N_5150);
and U8139 (N_8139,N_4781,N_4651);
nor U8140 (N_8140,N_3957,N_4459);
and U8141 (N_8141,N_5577,N_6228);
or U8142 (N_8142,N_3406,N_6235);
and U8143 (N_8143,N_4988,N_3247);
and U8144 (N_8144,N_5192,N_3284);
xor U8145 (N_8145,N_3702,N_5743);
nand U8146 (N_8146,N_3500,N_4311);
and U8147 (N_8147,N_4167,N_3413);
nor U8148 (N_8148,N_5014,N_6153);
and U8149 (N_8149,N_3762,N_6185);
nand U8150 (N_8150,N_6104,N_6139);
xnor U8151 (N_8151,N_4097,N_3441);
nand U8152 (N_8152,N_4014,N_4108);
xnor U8153 (N_8153,N_3855,N_5887);
xor U8154 (N_8154,N_5404,N_5505);
nor U8155 (N_8155,N_3475,N_4866);
and U8156 (N_8156,N_4791,N_6234);
nor U8157 (N_8157,N_3916,N_5174);
nand U8158 (N_8158,N_3431,N_5891);
and U8159 (N_8159,N_4140,N_3257);
or U8160 (N_8160,N_3428,N_5169);
nand U8161 (N_8161,N_5796,N_3999);
nor U8162 (N_8162,N_3988,N_6179);
nand U8163 (N_8163,N_3532,N_5482);
nor U8164 (N_8164,N_6241,N_3316);
nor U8165 (N_8165,N_4572,N_6133);
nand U8166 (N_8166,N_3174,N_4895);
nand U8167 (N_8167,N_5543,N_3635);
or U8168 (N_8168,N_3362,N_5093);
nor U8169 (N_8169,N_4787,N_5385);
xor U8170 (N_8170,N_5518,N_4054);
nand U8171 (N_8171,N_3641,N_3701);
nand U8172 (N_8172,N_6208,N_3376);
and U8173 (N_8173,N_4155,N_3416);
xnor U8174 (N_8174,N_4652,N_4961);
nand U8175 (N_8175,N_5973,N_5653);
nor U8176 (N_8176,N_4826,N_4106);
nand U8177 (N_8177,N_5899,N_5840);
nor U8178 (N_8178,N_4297,N_5112);
xor U8179 (N_8179,N_5907,N_3181);
xnor U8180 (N_8180,N_4676,N_5380);
nand U8181 (N_8181,N_3739,N_3409);
xor U8182 (N_8182,N_5297,N_5634);
nand U8183 (N_8183,N_5203,N_4732);
nor U8184 (N_8184,N_5555,N_4505);
nor U8185 (N_8185,N_5208,N_4204);
nand U8186 (N_8186,N_4545,N_5191);
or U8187 (N_8187,N_5958,N_3427);
xnor U8188 (N_8188,N_4530,N_3758);
or U8189 (N_8189,N_5821,N_3592);
or U8190 (N_8190,N_6162,N_4998);
nand U8191 (N_8191,N_5546,N_4657);
xnor U8192 (N_8192,N_5966,N_4118);
or U8193 (N_8193,N_5218,N_5576);
and U8194 (N_8194,N_5088,N_6006);
or U8195 (N_8195,N_5739,N_3833);
nand U8196 (N_8196,N_3186,N_5091);
nand U8197 (N_8197,N_3503,N_5807);
and U8198 (N_8198,N_4721,N_4151);
xor U8199 (N_8199,N_4151,N_3342);
nor U8200 (N_8200,N_3690,N_3527);
nand U8201 (N_8201,N_4245,N_3446);
or U8202 (N_8202,N_5945,N_3890);
or U8203 (N_8203,N_4838,N_4522);
nor U8204 (N_8204,N_3534,N_4621);
and U8205 (N_8205,N_4352,N_5857);
xor U8206 (N_8206,N_3253,N_5334);
and U8207 (N_8207,N_4318,N_5633);
and U8208 (N_8208,N_4077,N_4367);
or U8209 (N_8209,N_4096,N_3272);
xor U8210 (N_8210,N_4206,N_4056);
nand U8211 (N_8211,N_4888,N_3269);
nand U8212 (N_8212,N_5275,N_4892);
nand U8213 (N_8213,N_5876,N_4838);
nand U8214 (N_8214,N_3607,N_4308);
and U8215 (N_8215,N_4763,N_3621);
nand U8216 (N_8216,N_3402,N_3247);
and U8217 (N_8217,N_5388,N_5763);
nand U8218 (N_8218,N_5828,N_5179);
xor U8219 (N_8219,N_5975,N_6244);
nand U8220 (N_8220,N_5469,N_3481);
nor U8221 (N_8221,N_4216,N_4361);
nor U8222 (N_8222,N_3501,N_4230);
nand U8223 (N_8223,N_4324,N_3322);
and U8224 (N_8224,N_6156,N_4086);
nor U8225 (N_8225,N_3852,N_3641);
nor U8226 (N_8226,N_3515,N_3762);
or U8227 (N_8227,N_5590,N_4339);
nor U8228 (N_8228,N_5607,N_3650);
nand U8229 (N_8229,N_3559,N_3182);
nor U8230 (N_8230,N_5274,N_4454);
xnor U8231 (N_8231,N_3742,N_5269);
or U8232 (N_8232,N_3558,N_4995);
and U8233 (N_8233,N_5524,N_3750);
and U8234 (N_8234,N_5985,N_5313);
or U8235 (N_8235,N_4472,N_5517);
nand U8236 (N_8236,N_3661,N_4809);
or U8237 (N_8237,N_5902,N_3304);
nor U8238 (N_8238,N_5702,N_6026);
nor U8239 (N_8239,N_3614,N_4352);
and U8240 (N_8240,N_3378,N_4412);
or U8241 (N_8241,N_3215,N_3642);
and U8242 (N_8242,N_5452,N_6203);
or U8243 (N_8243,N_3202,N_4053);
xnor U8244 (N_8244,N_4701,N_4105);
and U8245 (N_8245,N_5568,N_4180);
or U8246 (N_8246,N_3301,N_5962);
xnor U8247 (N_8247,N_4505,N_4219);
and U8248 (N_8248,N_3660,N_3563);
nand U8249 (N_8249,N_3558,N_6019);
or U8250 (N_8250,N_4287,N_5057);
xor U8251 (N_8251,N_6055,N_3873);
nor U8252 (N_8252,N_5291,N_4123);
xnor U8253 (N_8253,N_4630,N_4153);
nor U8254 (N_8254,N_5660,N_5151);
or U8255 (N_8255,N_5692,N_6221);
xor U8256 (N_8256,N_3276,N_4013);
and U8257 (N_8257,N_6059,N_5232);
and U8258 (N_8258,N_5769,N_5519);
nand U8259 (N_8259,N_3542,N_3265);
nand U8260 (N_8260,N_4149,N_5896);
nand U8261 (N_8261,N_3740,N_4898);
nor U8262 (N_8262,N_3547,N_3620);
xor U8263 (N_8263,N_5302,N_3155);
nand U8264 (N_8264,N_4001,N_4392);
nand U8265 (N_8265,N_4643,N_5127);
nor U8266 (N_8266,N_3496,N_5116);
xnor U8267 (N_8267,N_5177,N_5935);
nand U8268 (N_8268,N_3886,N_4357);
nand U8269 (N_8269,N_4744,N_3659);
or U8270 (N_8270,N_3916,N_3278);
xor U8271 (N_8271,N_3308,N_6020);
nand U8272 (N_8272,N_5949,N_3143);
nor U8273 (N_8273,N_3569,N_3937);
nand U8274 (N_8274,N_5110,N_5115);
nor U8275 (N_8275,N_4996,N_5793);
nand U8276 (N_8276,N_5374,N_3770);
nor U8277 (N_8277,N_5658,N_4064);
nor U8278 (N_8278,N_3929,N_4763);
nor U8279 (N_8279,N_6076,N_4737);
nand U8280 (N_8280,N_3528,N_3493);
nor U8281 (N_8281,N_4875,N_4804);
or U8282 (N_8282,N_5804,N_6241);
or U8283 (N_8283,N_3940,N_3860);
nor U8284 (N_8284,N_4428,N_5621);
and U8285 (N_8285,N_5373,N_6088);
xor U8286 (N_8286,N_4839,N_4602);
nand U8287 (N_8287,N_5935,N_5291);
nand U8288 (N_8288,N_3470,N_3557);
xor U8289 (N_8289,N_4039,N_5504);
and U8290 (N_8290,N_3532,N_5181);
nor U8291 (N_8291,N_5475,N_5272);
or U8292 (N_8292,N_3175,N_4057);
nor U8293 (N_8293,N_4023,N_4943);
nor U8294 (N_8294,N_4045,N_6085);
or U8295 (N_8295,N_3385,N_3565);
and U8296 (N_8296,N_4375,N_4507);
or U8297 (N_8297,N_3818,N_5658);
or U8298 (N_8298,N_3895,N_4204);
nor U8299 (N_8299,N_4243,N_5668);
nor U8300 (N_8300,N_5452,N_4145);
xnor U8301 (N_8301,N_6125,N_3766);
and U8302 (N_8302,N_3185,N_5142);
nor U8303 (N_8303,N_5768,N_3649);
and U8304 (N_8304,N_4474,N_5116);
and U8305 (N_8305,N_5219,N_6012);
nor U8306 (N_8306,N_5195,N_4678);
nor U8307 (N_8307,N_4261,N_4465);
or U8308 (N_8308,N_5203,N_3799);
nor U8309 (N_8309,N_3452,N_4950);
nor U8310 (N_8310,N_5658,N_3922);
nand U8311 (N_8311,N_5671,N_4430);
nand U8312 (N_8312,N_6229,N_4144);
and U8313 (N_8313,N_3263,N_3900);
and U8314 (N_8314,N_4904,N_3751);
or U8315 (N_8315,N_5426,N_5073);
and U8316 (N_8316,N_4534,N_4880);
nand U8317 (N_8317,N_6051,N_4668);
or U8318 (N_8318,N_6046,N_3822);
and U8319 (N_8319,N_6010,N_4986);
nor U8320 (N_8320,N_5218,N_5004);
or U8321 (N_8321,N_5446,N_5561);
nand U8322 (N_8322,N_5721,N_5903);
xor U8323 (N_8323,N_3446,N_4041);
nand U8324 (N_8324,N_5960,N_5851);
or U8325 (N_8325,N_3375,N_3659);
or U8326 (N_8326,N_5630,N_5322);
nand U8327 (N_8327,N_5872,N_4499);
and U8328 (N_8328,N_3436,N_5263);
nor U8329 (N_8329,N_4597,N_4860);
nor U8330 (N_8330,N_5860,N_3996);
and U8331 (N_8331,N_4132,N_5870);
and U8332 (N_8332,N_4069,N_5223);
nor U8333 (N_8333,N_3135,N_5808);
or U8334 (N_8334,N_6030,N_4767);
nor U8335 (N_8335,N_5451,N_6199);
and U8336 (N_8336,N_4167,N_5494);
and U8337 (N_8337,N_3658,N_3558);
or U8338 (N_8338,N_4700,N_4009);
xnor U8339 (N_8339,N_3512,N_4194);
nor U8340 (N_8340,N_5718,N_3356);
xnor U8341 (N_8341,N_4502,N_3655);
or U8342 (N_8342,N_5314,N_4661);
nand U8343 (N_8343,N_5501,N_4620);
nand U8344 (N_8344,N_5775,N_6183);
nor U8345 (N_8345,N_3154,N_4374);
nand U8346 (N_8346,N_3662,N_5435);
and U8347 (N_8347,N_4574,N_5923);
xnor U8348 (N_8348,N_4077,N_3929);
nand U8349 (N_8349,N_3448,N_5859);
or U8350 (N_8350,N_4403,N_3560);
and U8351 (N_8351,N_4525,N_4581);
xnor U8352 (N_8352,N_4236,N_6151);
or U8353 (N_8353,N_4330,N_5833);
nand U8354 (N_8354,N_5249,N_4301);
nand U8355 (N_8355,N_5526,N_3551);
and U8356 (N_8356,N_4172,N_4132);
nor U8357 (N_8357,N_5017,N_5038);
nand U8358 (N_8358,N_3375,N_3523);
xor U8359 (N_8359,N_3462,N_3239);
nand U8360 (N_8360,N_5927,N_5006);
nor U8361 (N_8361,N_3862,N_4242);
xor U8362 (N_8362,N_4991,N_5652);
nor U8363 (N_8363,N_3325,N_5027);
nand U8364 (N_8364,N_5449,N_5052);
nand U8365 (N_8365,N_5531,N_4002);
nor U8366 (N_8366,N_5673,N_6162);
nand U8367 (N_8367,N_3208,N_4554);
and U8368 (N_8368,N_6053,N_3183);
nand U8369 (N_8369,N_5447,N_5365);
nand U8370 (N_8370,N_6084,N_3930);
nor U8371 (N_8371,N_5383,N_5817);
or U8372 (N_8372,N_3668,N_6139);
and U8373 (N_8373,N_3615,N_4741);
nand U8374 (N_8374,N_5253,N_4317);
nor U8375 (N_8375,N_4386,N_4798);
and U8376 (N_8376,N_5578,N_3477);
nand U8377 (N_8377,N_4555,N_4493);
or U8378 (N_8378,N_4598,N_3421);
nor U8379 (N_8379,N_5651,N_4878);
nand U8380 (N_8380,N_5087,N_4245);
nand U8381 (N_8381,N_4823,N_4791);
and U8382 (N_8382,N_4321,N_5690);
or U8383 (N_8383,N_5025,N_4503);
or U8384 (N_8384,N_4119,N_5215);
and U8385 (N_8385,N_6032,N_6076);
and U8386 (N_8386,N_3613,N_4578);
xor U8387 (N_8387,N_5895,N_5604);
or U8388 (N_8388,N_5298,N_3241);
xor U8389 (N_8389,N_5677,N_4952);
nand U8390 (N_8390,N_3907,N_4725);
xnor U8391 (N_8391,N_5066,N_5124);
nor U8392 (N_8392,N_5501,N_5832);
or U8393 (N_8393,N_6181,N_5888);
nor U8394 (N_8394,N_5890,N_4049);
xnor U8395 (N_8395,N_5924,N_6079);
and U8396 (N_8396,N_5596,N_5449);
nand U8397 (N_8397,N_5773,N_5141);
and U8398 (N_8398,N_3512,N_4475);
and U8399 (N_8399,N_5599,N_3806);
and U8400 (N_8400,N_6164,N_4321);
and U8401 (N_8401,N_4281,N_4728);
and U8402 (N_8402,N_3233,N_5448);
nor U8403 (N_8403,N_5691,N_3559);
nand U8404 (N_8404,N_5645,N_4308);
and U8405 (N_8405,N_5048,N_4820);
nand U8406 (N_8406,N_6160,N_3693);
or U8407 (N_8407,N_5971,N_4878);
and U8408 (N_8408,N_3475,N_6021);
or U8409 (N_8409,N_4956,N_4245);
nand U8410 (N_8410,N_3510,N_5789);
or U8411 (N_8411,N_5476,N_4450);
xor U8412 (N_8412,N_6028,N_5009);
and U8413 (N_8413,N_3718,N_4295);
nor U8414 (N_8414,N_4785,N_4881);
or U8415 (N_8415,N_4430,N_5676);
nor U8416 (N_8416,N_5495,N_5040);
nor U8417 (N_8417,N_5503,N_5006);
nor U8418 (N_8418,N_5521,N_4861);
nand U8419 (N_8419,N_6134,N_4492);
nor U8420 (N_8420,N_4720,N_4273);
nand U8421 (N_8421,N_4438,N_3701);
nand U8422 (N_8422,N_4345,N_4042);
or U8423 (N_8423,N_5647,N_6189);
nand U8424 (N_8424,N_5575,N_6176);
xor U8425 (N_8425,N_3773,N_5228);
nor U8426 (N_8426,N_4201,N_4902);
or U8427 (N_8427,N_5328,N_5953);
nand U8428 (N_8428,N_5914,N_4406);
xnor U8429 (N_8429,N_5992,N_4912);
nor U8430 (N_8430,N_3564,N_3304);
nand U8431 (N_8431,N_4325,N_3212);
or U8432 (N_8432,N_5291,N_5405);
nor U8433 (N_8433,N_5699,N_3583);
or U8434 (N_8434,N_5822,N_4088);
nand U8435 (N_8435,N_3269,N_5112);
and U8436 (N_8436,N_4038,N_3225);
nand U8437 (N_8437,N_5014,N_5075);
nand U8438 (N_8438,N_3564,N_6175);
and U8439 (N_8439,N_5295,N_3264);
nor U8440 (N_8440,N_3725,N_3327);
nand U8441 (N_8441,N_4503,N_3360);
or U8442 (N_8442,N_6004,N_4619);
nor U8443 (N_8443,N_4805,N_5899);
xnor U8444 (N_8444,N_5260,N_3874);
nand U8445 (N_8445,N_5173,N_3465);
or U8446 (N_8446,N_4530,N_5518);
xor U8447 (N_8447,N_3957,N_4896);
and U8448 (N_8448,N_4386,N_3220);
and U8449 (N_8449,N_4098,N_6106);
nor U8450 (N_8450,N_4419,N_5584);
nor U8451 (N_8451,N_3138,N_3337);
nor U8452 (N_8452,N_5055,N_3793);
and U8453 (N_8453,N_3191,N_4043);
xnor U8454 (N_8454,N_4498,N_4980);
and U8455 (N_8455,N_4895,N_3258);
or U8456 (N_8456,N_3406,N_5152);
and U8457 (N_8457,N_4779,N_5181);
or U8458 (N_8458,N_4743,N_3495);
or U8459 (N_8459,N_4797,N_5032);
nand U8460 (N_8460,N_5736,N_6012);
or U8461 (N_8461,N_4718,N_4850);
nor U8462 (N_8462,N_5080,N_5620);
nor U8463 (N_8463,N_5923,N_3586);
or U8464 (N_8464,N_4528,N_4870);
nand U8465 (N_8465,N_5060,N_5992);
and U8466 (N_8466,N_5782,N_4440);
nor U8467 (N_8467,N_4747,N_3447);
xor U8468 (N_8468,N_5271,N_3364);
and U8469 (N_8469,N_3268,N_4437);
and U8470 (N_8470,N_4295,N_3962);
or U8471 (N_8471,N_5598,N_6003);
nand U8472 (N_8472,N_4151,N_3709);
and U8473 (N_8473,N_6123,N_5615);
xor U8474 (N_8474,N_5563,N_5139);
nand U8475 (N_8475,N_3399,N_4948);
nor U8476 (N_8476,N_3724,N_5028);
and U8477 (N_8477,N_5717,N_3959);
xnor U8478 (N_8478,N_3800,N_5607);
nand U8479 (N_8479,N_3444,N_6216);
xor U8480 (N_8480,N_5955,N_3559);
nand U8481 (N_8481,N_4875,N_5371);
xnor U8482 (N_8482,N_5320,N_3812);
nor U8483 (N_8483,N_5703,N_4656);
nand U8484 (N_8484,N_4936,N_3811);
nor U8485 (N_8485,N_4445,N_5727);
nand U8486 (N_8486,N_3508,N_6132);
and U8487 (N_8487,N_3801,N_4818);
or U8488 (N_8488,N_5823,N_5313);
xnor U8489 (N_8489,N_6096,N_5510);
or U8490 (N_8490,N_5706,N_5730);
nand U8491 (N_8491,N_4926,N_3577);
nand U8492 (N_8492,N_5667,N_4150);
or U8493 (N_8493,N_4751,N_4376);
or U8494 (N_8494,N_3259,N_3796);
and U8495 (N_8495,N_4428,N_4252);
or U8496 (N_8496,N_5370,N_4794);
or U8497 (N_8497,N_5387,N_5084);
xor U8498 (N_8498,N_4468,N_3523);
xor U8499 (N_8499,N_3617,N_3484);
and U8500 (N_8500,N_4112,N_4417);
and U8501 (N_8501,N_4553,N_4809);
nor U8502 (N_8502,N_6026,N_3400);
nor U8503 (N_8503,N_5387,N_3811);
nor U8504 (N_8504,N_5545,N_4208);
and U8505 (N_8505,N_5547,N_5457);
or U8506 (N_8506,N_3370,N_4745);
or U8507 (N_8507,N_5415,N_3189);
xor U8508 (N_8508,N_4455,N_5921);
and U8509 (N_8509,N_5033,N_6070);
nor U8510 (N_8510,N_3708,N_5667);
nor U8511 (N_8511,N_6155,N_5618);
and U8512 (N_8512,N_5405,N_4935);
xor U8513 (N_8513,N_4544,N_4601);
xor U8514 (N_8514,N_5984,N_5634);
nor U8515 (N_8515,N_4160,N_4553);
nand U8516 (N_8516,N_4405,N_5468);
nor U8517 (N_8517,N_6241,N_4776);
or U8518 (N_8518,N_4468,N_4253);
and U8519 (N_8519,N_5085,N_5324);
nand U8520 (N_8520,N_3161,N_4084);
nand U8521 (N_8521,N_3317,N_5649);
or U8522 (N_8522,N_4691,N_4236);
and U8523 (N_8523,N_4664,N_5349);
or U8524 (N_8524,N_5592,N_4192);
xor U8525 (N_8525,N_5137,N_5342);
nor U8526 (N_8526,N_3162,N_4306);
nand U8527 (N_8527,N_6119,N_3911);
xor U8528 (N_8528,N_5727,N_4550);
xnor U8529 (N_8529,N_3541,N_5544);
nand U8530 (N_8530,N_3364,N_5486);
xnor U8531 (N_8531,N_3757,N_6145);
nor U8532 (N_8532,N_3735,N_3993);
xnor U8533 (N_8533,N_3805,N_3830);
xnor U8534 (N_8534,N_5968,N_4743);
and U8535 (N_8535,N_5691,N_4518);
or U8536 (N_8536,N_3536,N_4193);
nor U8537 (N_8537,N_3130,N_3376);
xor U8538 (N_8538,N_4082,N_3998);
nand U8539 (N_8539,N_4936,N_4939);
nor U8540 (N_8540,N_5457,N_4759);
and U8541 (N_8541,N_3941,N_3299);
nor U8542 (N_8542,N_6203,N_4356);
and U8543 (N_8543,N_3268,N_4168);
nand U8544 (N_8544,N_5702,N_6050);
and U8545 (N_8545,N_4216,N_5189);
or U8546 (N_8546,N_6223,N_4459);
nor U8547 (N_8547,N_3527,N_4784);
nor U8548 (N_8548,N_3936,N_3662);
and U8549 (N_8549,N_3625,N_3555);
or U8550 (N_8550,N_5257,N_3230);
and U8551 (N_8551,N_4417,N_4069);
and U8552 (N_8552,N_3530,N_3415);
nor U8553 (N_8553,N_4928,N_6183);
xnor U8554 (N_8554,N_4352,N_3758);
xnor U8555 (N_8555,N_3338,N_4068);
nand U8556 (N_8556,N_4580,N_4452);
nor U8557 (N_8557,N_5324,N_4490);
nor U8558 (N_8558,N_3642,N_3216);
nor U8559 (N_8559,N_5220,N_5710);
nor U8560 (N_8560,N_3610,N_3893);
xor U8561 (N_8561,N_6220,N_5464);
nand U8562 (N_8562,N_4340,N_5366);
nor U8563 (N_8563,N_3395,N_4506);
xnor U8564 (N_8564,N_4692,N_3153);
nor U8565 (N_8565,N_4953,N_5302);
and U8566 (N_8566,N_3875,N_4768);
nand U8567 (N_8567,N_6209,N_3541);
nor U8568 (N_8568,N_4210,N_3547);
and U8569 (N_8569,N_5422,N_5857);
nor U8570 (N_8570,N_4257,N_3996);
xor U8571 (N_8571,N_6192,N_3142);
nor U8572 (N_8572,N_4035,N_3701);
and U8573 (N_8573,N_5871,N_3368);
nand U8574 (N_8574,N_3564,N_6118);
or U8575 (N_8575,N_5362,N_3940);
xor U8576 (N_8576,N_5708,N_5195);
nand U8577 (N_8577,N_3706,N_3893);
or U8578 (N_8578,N_6226,N_3154);
xnor U8579 (N_8579,N_3460,N_5049);
and U8580 (N_8580,N_4508,N_4775);
nor U8581 (N_8581,N_5992,N_4457);
nand U8582 (N_8582,N_5674,N_3404);
xor U8583 (N_8583,N_3466,N_5817);
nand U8584 (N_8584,N_5575,N_5625);
xnor U8585 (N_8585,N_3871,N_3887);
xor U8586 (N_8586,N_3651,N_4146);
nand U8587 (N_8587,N_5150,N_3551);
and U8588 (N_8588,N_4843,N_5157);
nand U8589 (N_8589,N_4973,N_5870);
nand U8590 (N_8590,N_3642,N_3246);
and U8591 (N_8591,N_5326,N_3245);
or U8592 (N_8592,N_5213,N_3632);
or U8593 (N_8593,N_5978,N_6075);
nor U8594 (N_8594,N_4160,N_4958);
or U8595 (N_8595,N_5511,N_5949);
nand U8596 (N_8596,N_5496,N_5888);
and U8597 (N_8597,N_5461,N_3637);
nand U8598 (N_8598,N_4081,N_6133);
nand U8599 (N_8599,N_4978,N_5229);
and U8600 (N_8600,N_4119,N_4102);
xor U8601 (N_8601,N_5599,N_5949);
and U8602 (N_8602,N_3859,N_4108);
xor U8603 (N_8603,N_3771,N_5726);
or U8604 (N_8604,N_4971,N_4870);
and U8605 (N_8605,N_3674,N_4232);
nor U8606 (N_8606,N_5094,N_3208);
xor U8607 (N_8607,N_4487,N_4948);
nand U8608 (N_8608,N_4940,N_4129);
nor U8609 (N_8609,N_6107,N_3500);
nand U8610 (N_8610,N_5323,N_4623);
or U8611 (N_8611,N_3417,N_4675);
xnor U8612 (N_8612,N_3964,N_5433);
xnor U8613 (N_8613,N_4210,N_4358);
nor U8614 (N_8614,N_5415,N_3284);
and U8615 (N_8615,N_3913,N_3272);
nand U8616 (N_8616,N_5968,N_3654);
and U8617 (N_8617,N_3997,N_4514);
nand U8618 (N_8618,N_5541,N_5085);
and U8619 (N_8619,N_6089,N_3913);
xor U8620 (N_8620,N_5410,N_5583);
or U8621 (N_8621,N_4392,N_4743);
or U8622 (N_8622,N_5404,N_6165);
or U8623 (N_8623,N_4926,N_4990);
nor U8624 (N_8624,N_5201,N_3453);
nand U8625 (N_8625,N_5309,N_5798);
xnor U8626 (N_8626,N_5744,N_4950);
and U8627 (N_8627,N_4449,N_3669);
and U8628 (N_8628,N_5671,N_5564);
or U8629 (N_8629,N_4421,N_3899);
nand U8630 (N_8630,N_3633,N_3690);
or U8631 (N_8631,N_5190,N_5071);
or U8632 (N_8632,N_3200,N_4685);
and U8633 (N_8633,N_3288,N_3502);
or U8634 (N_8634,N_4170,N_5567);
nor U8635 (N_8635,N_4431,N_4393);
and U8636 (N_8636,N_4905,N_5894);
and U8637 (N_8637,N_3133,N_4865);
and U8638 (N_8638,N_6215,N_5007);
or U8639 (N_8639,N_5844,N_4660);
xnor U8640 (N_8640,N_4199,N_3530);
xor U8641 (N_8641,N_5643,N_5436);
xor U8642 (N_8642,N_5197,N_3254);
and U8643 (N_8643,N_3607,N_4535);
nand U8644 (N_8644,N_4796,N_3475);
nor U8645 (N_8645,N_3353,N_4440);
or U8646 (N_8646,N_5657,N_4190);
nand U8647 (N_8647,N_5077,N_5279);
and U8648 (N_8648,N_4596,N_5964);
and U8649 (N_8649,N_5412,N_5760);
xnor U8650 (N_8650,N_4017,N_4088);
nand U8651 (N_8651,N_3232,N_5005);
nor U8652 (N_8652,N_3178,N_5787);
xnor U8653 (N_8653,N_6211,N_5542);
and U8654 (N_8654,N_3918,N_4396);
nor U8655 (N_8655,N_4963,N_6183);
and U8656 (N_8656,N_3679,N_5324);
nand U8657 (N_8657,N_4129,N_5533);
or U8658 (N_8658,N_5413,N_3965);
or U8659 (N_8659,N_4953,N_4565);
nand U8660 (N_8660,N_5364,N_3886);
nand U8661 (N_8661,N_5510,N_3301);
nor U8662 (N_8662,N_3949,N_5105);
nor U8663 (N_8663,N_5156,N_4316);
xor U8664 (N_8664,N_5759,N_3443);
or U8665 (N_8665,N_4510,N_4755);
nand U8666 (N_8666,N_3889,N_4743);
and U8667 (N_8667,N_5823,N_5592);
nor U8668 (N_8668,N_5603,N_5003);
nor U8669 (N_8669,N_3653,N_5621);
or U8670 (N_8670,N_4849,N_5902);
xor U8671 (N_8671,N_5940,N_3518);
and U8672 (N_8672,N_4650,N_4876);
nand U8673 (N_8673,N_5739,N_5421);
or U8674 (N_8674,N_3791,N_5269);
nand U8675 (N_8675,N_5547,N_6227);
and U8676 (N_8676,N_5599,N_3472);
nor U8677 (N_8677,N_5781,N_4718);
nor U8678 (N_8678,N_5971,N_5357);
xor U8679 (N_8679,N_5065,N_3706);
nand U8680 (N_8680,N_5838,N_4143);
nor U8681 (N_8681,N_5182,N_4049);
nor U8682 (N_8682,N_5080,N_3899);
nand U8683 (N_8683,N_3257,N_5261);
or U8684 (N_8684,N_3956,N_5744);
xor U8685 (N_8685,N_4407,N_5400);
nand U8686 (N_8686,N_4731,N_5803);
xnor U8687 (N_8687,N_3951,N_6181);
and U8688 (N_8688,N_3954,N_5504);
nor U8689 (N_8689,N_5967,N_4590);
or U8690 (N_8690,N_3302,N_4718);
xor U8691 (N_8691,N_3343,N_4584);
nor U8692 (N_8692,N_6052,N_4981);
and U8693 (N_8693,N_4531,N_3704);
or U8694 (N_8694,N_3683,N_3165);
nor U8695 (N_8695,N_4601,N_4952);
nand U8696 (N_8696,N_3240,N_5808);
nand U8697 (N_8697,N_3573,N_4523);
and U8698 (N_8698,N_4064,N_5158);
xor U8699 (N_8699,N_4941,N_6109);
nand U8700 (N_8700,N_5236,N_6100);
xor U8701 (N_8701,N_4839,N_4918);
nor U8702 (N_8702,N_5073,N_5550);
xnor U8703 (N_8703,N_4681,N_4111);
nand U8704 (N_8704,N_3741,N_5369);
or U8705 (N_8705,N_3482,N_3288);
or U8706 (N_8706,N_3322,N_4130);
nor U8707 (N_8707,N_4464,N_3136);
and U8708 (N_8708,N_3371,N_5807);
xnor U8709 (N_8709,N_6095,N_5407);
and U8710 (N_8710,N_3178,N_4248);
and U8711 (N_8711,N_3174,N_4906);
xnor U8712 (N_8712,N_3522,N_3711);
and U8713 (N_8713,N_3623,N_5349);
xor U8714 (N_8714,N_3209,N_3925);
nor U8715 (N_8715,N_5042,N_5423);
nand U8716 (N_8716,N_5473,N_5565);
nand U8717 (N_8717,N_3343,N_5413);
xor U8718 (N_8718,N_3227,N_5683);
or U8719 (N_8719,N_5522,N_5084);
and U8720 (N_8720,N_3798,N_5099);
or U8721 (N_8721,N_5351,N_5456);
and U8722 (N_8722,N_5406,N_6187);
and U8723 (N_8723,N_5232,N_4209);
nand U8724 (N_8724,N_4891,N_4509);
nand U8725 (N_8725,N_4866,N_6042);
xnor U8726 (N_8726,N_3236,N_6022);
xnor U8727 (N_8727,N_4238,N_4606);
nand U8728 (N_8728,N_3423,N_4623);
or U8729 (N_8729,N_4721,N_5851);
nor U8730 (N_8730,N_4645,N_3516);
nor U8731 (N_8731,N_6029,N_4152);
or U8732 (N_8732,N_4623,N_4938);
nor U8733 (N_8733,N_4788,N_5329);
nor U8734 (N_8734,N_5736,N_4691);
or U8735 (N_8735,N_3212,N_5642);
or U8736 (N_8736,N_3558,N_3413);
nor U8737 (N_8737,N_5581,N_4578);
and U8738 (N_8738,N_4102,N_6194);
or U8739 (N_8739,N_3677,N_5221);
xor U8740 (N_8740,N_4473,N_3593);
nor U8741 (N_8741,N_5064,N_4956);
nor U8742 (N_8742,N_5918,N_5504);
nor U8743 (N_8743,N_3287,N_4217);
nand U8744 (N_8744,N_5031,N_6114);
nor U8745 (N_8745,N_4918,N_5715);
nor U8746 (N_8746,N_6004,N_5322);
nand U8747 (N_8747,N_3493,N_3220);
nor U8748 (N_8748,N_5792,N_5171);
nor U8749 (N_8749,N_4682,N_3942);
or U8750 (N_8750,N_4782,N_5850);
or U8751 (N_8751,N_5002,N_5543);
and U8752 (N_8752,N_3573,N_5725);
or U8753 (N_8753,N_3929,N_3882);
and U8754 (N_8754,N_4144,N_3220);
nand U8755 (N_8755,N_3819,N_3954);
or U8756 (N_8756,N_3827,N_3992);
xnor U8757 (N_8757,N_5502,N_4607);
nor U8758 (N_8758,N_3784,N_3586);
or U8759 (N_8759,N_4211,N_6233);
and U8760 (N_8760,N_5354,N_5233);
nand U8761 (N_8761,N_3480,N_4675);
or U8762 (N_8762,N_4749,N_4664);
or U8763 (N_8763,N_5777,N_5136);
nor U8764 (N_8764,N_3416,N_3862);
nor U8765 (N_8765,N_3310,N_5829);
nand U8766 (N_8766,N_4271,N_3540);
or U8767 (N_8767,N_4933,N_4192);
and U8768 (N_8768,N_6077,N_3853);
nand U8769 (N_8769,N_4036,N_3859);
or U8770 (N_8770,N_5937,N_3763);
and U8771 (N_8771,N_5449,N_5551);
or U8772 (N_8772,N_6018,N_4834);
xor U8773 (N_8773,N_6242,N_4701);
nand U8774 (N_8774,N_6193,N_5468);
nand U8775 (N_8775,N_5003,N_4829);
nand U8776 (N_8776,N_3753,N_3652);
xnor U8777 (N_8777,N_5065,N_5507);
or U8778 (N_8778,N_3639,N_3724);
and U8779 (N_8779,N_5025,N_5768);
and U8780 (N_8780,N_4828,N_3452);
nor U8781 (N_8781,N_4101,N_4451);
nor U8782 (N_8782,N_6169,N_3227);
or U8783 (N_8783,N_6108,N_4543);
and U8784 (N_8784,N_5238,N_4851);
xor U8785 (N_8785,N_5929,N_4819);
and U8786 (N_8786,N_5175,N_4738);
nor U8787 (N_8787,N_4310,N_6060);
xnor U8788 (N_8788,N_5945,N_5348);
and U8789 (N_8789,N_3534,N_3700);
and U8790 (N_8790,N_5790,N_5434);
nor U8791 (N_8791,N_5308,N_3656);
or U8792 (N_8792,N_3859,N_4616);
nand U8793 (N_8793,N_4204,N_4332);
or U8794 (N_8794,N_4985,N_5444);
nand U8795 (N_8795,N_5801,N_4005);
nor U8796 (N_8796,N_5613,N_3167);
and U8797 (N_8797,N_5513,N_5455);
and U8798 (N_8798,N_5107,N_6016);
nand U8799 (N_8799,N_5812,N_4146);
nand U8800 (N_8800,N_4078,N_4924);
or U8801 (N_8801,N_5395,N_5240);
and U8802 (N_8802,N_3561,N_5742);
xor U8803 (N_8803,N_4801,N_5229);
xor U8804 (N_8804,N_3508,N_3394);
and U8805 (N_8805,N_5134,N_6164);
nand U8806 (N_8806,N_5094,N_4270);
nand U8807 (N_8807,N_4897,N_4896);
nor U8808 (N_8808,N_3687,N_3986);
nor U8809 (N_8809,N_5907,N_6162);
nor U8810 (N_8810,N_4300,N_5596);
nand U8811 (N_8811,N_4494,N_3329);
or U8812 (N_8812,N_4571,N_4915);
and U8813 (N_8813,N_4242,N_5480);
or U8814 (N_8814,N_3545,N_4745);
xor U8815 (N_8815,N_4792,N_3428);
and U8816 (N_8816,N_3237,N_5107);
nor U8817 (N_8817,N_5511,N_5691);
or U8818 (N_8818,N_4741,N_4594);
nor U8819 (N_8819,N_4916,N_3701);
or U8820 (N_8820,N_3697,N_3522);
nor U8821 (N_8821,N_4342,N_4225);
xor U8822 (N_8822,N_3232,N_3935);
nand U8823 (N_8823,N_5690,N_3792);
nor U8824 (N_8824,N_4031,N_4396);
xnor U8825 (N_8825,N_3413,N_5681);
and U8826 (N_8826,N_4073,N_3702);
xor U8827 (N_8827,N_5641,N_4344);
xor U8828 (N_8828,N_5423,N_6152);
nand U8829 (N_8829,N_4285,N_5426);
nand U8830 (N_8830,N_5452,N_5478);
nor U8831 (N_8831,N_4571,N_3372);
xor U8832 (N_8832,N_4176,N_3238);
nand U8833 (N_8833,N_4449,N_5814);
xnor U8834 (N_8834,N_3603,N_6175);
or U8835 (N_8835,N_4723,N_4769);
nand U8836 (N_8836,N_6010,N_5256);
xnor U8837 (N_8837,N_4796,N_4811);
xor U8838 (N_8838,N_3403,N_4136);
and U8839 (N_8839,N_4652,N_6233);
nand U8840 (N_8840,N_5918,N_4412);
nor U8841 (N_8841,N_5698,N_4687);
xnor U8842 (N_8842,N_4260,N_5855);
and U8843 (N_8843,N_3770,N_4804);
or U8844 (N_8844,N_3782,N_6044);
xor U8845 (N_8845,N_5668,N_3949);
or U8846 (N_8846,N_5925,N_4820);
and U8847 (N_8847,N_5087,N_5207);
or U8848 (N_8848,N_5534,N_5632);
or U8849 (N_8849,N_4959,N_4908);
and U8850 (N_8850,N_4547,N_4085);
and U8851 (N_8851,N_6246,N_4254);
or U8852 (N_8852,N_4276,N_4763);
nand U8853 (N_8853,N_3220,N_4197);
and U8854 (N_8854,N_5597,N_4947);
nor U8855 (N_8855,N_3265,N_4751);
and U8856 (N_8856,N_5171,N_3481);
and U8857 (N_8857,N_5074,N_3258);
nor U8858 (N_8858,N_3359,N_4755);
xor U8859 (N_8859,N_5052,N_4746);
nor U8860 (N_8860,N_5247,N_5900);
nand U8861 (N_8861,N_3237,N_4542);
xnor U8862 (N_8862,N_4237,N_3285);
and U8863 (N_8863,N_5215,N_4734);
nor U8864 (N_8864,N_4272,N_5902);
xnor U8865 (N_8865,N_4807,N_3465);
or U8866 (N_8866,N_3426,N_5038);
and U8867 (N_8867,N_3418,N_5338);
nor U8868 (N_8868,N_4031,N_3139);
nand U8869 (N_8869,N_5099,N_5046);
nor U8870 (N_8870,N_5200,N_3756);
nand U8871 (N_8871,N_3334,N_5509);
and U8872 (N_8872,N_5925,N_6229);
and U8873 (N_8873,N_5961,N_3174);
nand U8874 (N_8874,N_4584,N_4926);
nor U8875 (N_8875,N_6189,N_5698);
and U8876 (N_8876,N_3244,N_5254);
nor U8877 (N_8877,N_3476,N_4234);
nor U8878 (N_8878,N_5699,N_3663);
and U8879 (N_8879,N_3243,N_6232);
xnor U8880 (N_8880,N_4129,N_4543);
or U8881 (N_8881,N_3946,N_3595);
xnor U8882 (N_8882,N_4045,N_3535);
xor U8883 (N_8883,N_4349,N_5448);
xnor U8884 (N_8884,N_3557,N_4919);
nor U8885 (N_8885,N_5447,N_3125);
xnor U8886 (N_8886,N_5664,N_5016);
xnor U8887 (N_8887,N_4149,N_6058);
nor U8888 (N_8888,N_4505,N_4553);
xnor U8889 (N_8889,N_5477,N_5518);
and U8890 (N_8890,N_5151,N_4567);
nor U8891 (N_8891,N_5934,N_4332);
nor U8892 (N_8892,N_4676,N_6246);
nand U8893 (N_8893,N_4651,N_5126);
nor U8894 (N_8894,N_4715,N_4193);
xor U8895 (N_8895,N_3460,N_4471);
nor U8896 (N_8896,N_5452,N_6181);
xor U8897 (N_8897,N_4079,N_5303);
or U8898 (N_8898,N_3894,N_3530);
or U8899 (N_8899,N_5515,N_5783);
or U8900 (N_8900,N_4669,N_3271);
xor U8901 (N_8901,N_5759,N_4720);
nand U8902 (N_8902,N_4850,N_6139);
or U8903 (N_8903,N_3696,N_4266);
nand U8904 (N_8904,N_4832,N_3126);
and U8905 (N_8905,N_4916,N_5714);
and U8906 (N_8906,N_4303,N_3776);
nand U8907 (N_8907,N_5532,N_5135);
xnor U8908 (N_8908,N_3439,N_4576);
xnor U8909 (N_8909,N_3548,N_4812);
nand U8910 (N_8910,N_3561,N_5855);
or U8911 (N_8911,N_4124,N_3384);
or U8912 (N_8912,N_4403,N_4414);
nand U8913 (N_8913,N_3743,N_5707);
and U8914 (N_8914,N_6198,N_4360);
xor U8915 (N_8915,N_4666,N_6115);
or U8916 (N_8916,N_3487,N_3845);
nor U8917 (N_8917,N_3271,N_5501);
and U8918 (N_8918,N_3306,N_4601);
nor U8919 (N_8919,N_4182,N_3694);
nand U8920 (N_8920,N_4629,N_5641);
or U8921 (N_8921,N_4416,N_4011);
nand U8922 (N_8922,N_3226,N_4244);
nand U8923 (N_8923,N_5028,N_3343);
nor U8924 (N_8924,N_5170,N_5433);
nor U8925 (N_8925,N_5706,N_4280);
nor U8926 (N_8926,N_3612,N_4569);
nor U8927 (N_8927,N_3761,N_4294);
nand U8928 (N_8928,N_3476,N_5188);
nand U8929 (N_8929,N_3898,N_4455);
or U8930 (N_8930,N_3887,N_3574);
nor U8931 (N_8931,N_3149,N_5495);
or U8932 (N_8932,N_5923,N_4681);
and U8933 (N_8933,N_4494,N_5773);
xor U8934 (N_8934,N_3170,N_4952);
nand U8935 (N_8935,N_5073,N_3568);
nand U8936 (N_8936,N_4304,N_4675);
or U8937 (N_8937,N_3996,N_3335);
nor U8938 (N_8938,N_4458,N_5251);
xnor U8939 (N_8939,N_3296,N_4610);
or U8940 (N_8940,N_5903,N_3324);
nor U8941 (N_8941,N_4299,N_5070);
xor U8942 (N_8942,N_4361,N_6014);
and U8943 (N_8943,N_3983,N_5435);
or U8944 (N_8944,N_5505,N_3497);
xnor U8945 (N_8945,N_3725,N_4719);
nor U8946 (N_8946,N_3714,N_5670);
xnor U8947 (N_8947,N_6118,N_4275);
nor U8948 (N_8948,N_3315,N_5476);
and U8949 (N_8949,N_4042,N_3737);
nor U8950 (N_8950,N_3431,N_3214);
nor U8951 (N_8951,N_4223,N_4855);
nand U8952 (N_8952,N_5788,N_4445);
nor U8953 (N_8953,N_5765,N_3728);
and U8954 (N_8954,N_3139,N_5767);
nand U8955 (N_8955,N_5535,N_4761);
nor U8956 (N_8956,N_4651,N_5716);
xnor U8957 (N_8957,N_3273,N_4094);
xor U8958 (N_8958,N_4372,N_4466);
nand U8959 (N_8959,N_3812,N_5245);
nor U8960 (N_8960,N_5437,N_3646);
or U8961 (N_8961,N_3884,N_4216);
and U8962 (N_8962,N_4133,N_4311);
and U8963 (N_8963,N_5921,N_6147);
and U8964 (N_8964,N_3482,N_4837);
xor U8965 (N_8965,N_5579,N_4378);
nor U8966 (N_8966,N_5181,N_6062);
xor U8967 (N_8967,N_4650,N_4557);
nor U8968 (N_8968,N_4589,N_5472);
nand U8969 (N_8969,N_4404,N_4065);
nor U8970 (N_8970,N_5762,N_3757);
and U8971 (N_8971,N_4550,N_4571);
xnor U8972 (N_8972,N_5355,N_5004);
and U8973 (N_8973,N_5189,N_5356);
and U8974 (N_8974,N_3290,N_3373);
or U8975 (N_8975,N_3202,N_5672);
nor U8976 (N_8976,N_3683,N_6219);
xnor U8977 (N_8977,N_5215,N_4657);
nor U8978 (N_8978,N_5215,N_4254);
nor U8979 (N_8979,N_5381,N_6192);
and U8980 (N_8980,N_5876,N_4545);
nor U8981 (N_8981,N_4970,N_4932);
nand U8982 (N_8982,N_5674,N_6021);
xnor U8983 (N_8983,N_4911,N_5676);
nand U8984 (N_8984,N_5994,N_6079);
and U8985 (N_8985,N_3886,N_5904);
nor U8986 (N_8986,N_3565,N_4927);
nand U8987 (N_8987,N_3209,N_5073);
nor U8988 (N_8988,N_3997,N_4876);
or U8989 (N_8989,N_5392,N_4302);
nor U8990 (N_8990,N_5684,N_5724);
nand U8991 (N_8991,N_6067,N_4027);
nand U8992 (N_8992,N_5181,N_5550);
xnor U8993 (N_8993,N_4091,N_4276);
xor U8994 (N_8994,N_3231,N_5514);
nand U8995 (N_8995,N_3348,N_5003);
xnor U8996 (N_8996,N_4755,N_4130);
xnor U8997 (N_8997,N_5162,N_5768);
xor U8998 (N_8998,N_4258,N_6067);
and U8999 (N_8999,N_4875,N_5859);
nor U9000 (N_9000,N_5592,N_4517);
and U9001 (N_9001,N_6018,N_4304);
nor U9002 (N_9002,N_4570,N_5128);
or U9003 (N_9003,N_4022,N_4580);
and U9004 (N_9004,N_6240,N_6026);
or U9005 (N_9005,N_3691,N_5435);
and U9006 (N_9006,N_4410,N_5184);
nand U9007 (N_9007,N_4542,N_4492);
nor U9008 (N_9008,N_5047,N_5582);
nor U9009 (N_9009,N_4306,N_5358);
nand U9010 (N_9010,N_3908,N_4442);
xnor U9011 (N_9011,N_3225,N_5153);
and U9012 (N_9012,N_3431,N_5342);
or U9013 (N_9013,N_4630,N_6012);
and U9014 (N_9014,N_4112,N_3440);
xnor U9015 (N_9015,N_6235,N_3160);
nor U9016 (N_9016,N_3177,N_6115);
and U9017 (N_9017,N_4918,N_4676);
or U9018 (N_9018,N_3894,N_4492);
or U9019 (N_9019,N_5148,N_4530);
and U9020 (N_9020,N_3587,N_6231);
xnor U9021 (N_9021,N_3932,N_4939);
or U9022 (N_9022,N_5174,N_3978);
and U9023 (N_9023,N_5082,N_4395);
nor U9024 (N_9024,N_3717,N_3765);
nand U9025 (N_9025,N_3357,N_4604);
nand U9026 (N_9026,N_5032,N_5468);
nor U9027 (N_9027,N_3634,N_3678);
and U9028 (N_9028,N_3264,N_3453);
nand U9029 (N_9029,N_5418,N_5893);
xnor U9030 (N_9030,N_4748,N_4292);
xor U9031 (N_9031,N_3433,N_4261);
nor U9032 (N_9032,N_5422,N_4139);
and U9033 (N_9033,N_4913,N_6089);
xnor U9034 (N_9034,N_4201,N_4566);
nand U9035 (N_9035,N_5191,N_5768);
xnor U9036 (N_9036,N_3780,N_5253);
nand U9037 (N_9037,N_5952,N_5188);
nand U9038 (N_9038,N_6192,N_4699);
nand U9039 (N_9039,N_5589,N_3332);
nand U9040 (N_9040,N_4309,N_3269);
or U9041 (N_9041,N_3211,N_4684);
nor U9042 (N_9042,N_4780,N_5878);
xor U9043 (N_9043,N_5059,N_6217);
nand U9044 (N_9044,N_4369,N_5050);
xnor U9045 (N_9045,N_5462,N_4296);
nand U9046 (N_9046,N_3978,N_4070);
nor U9047 (N_9047,N_5790,N_4274);
nor U9048 (N_9048,N_4978,N_5230);
xnor U9049 (N_9049,N_4001,N_3275);
nor U9050 (N_9050,N_4849,N_3230);
xnor U9051 (N_9051,N_3286,N_3735);
xor U9052 (N_9052,N_5958,N_4230);
and U9053 (N_9053,N_5499,N_4068);
or U9054 (N_9054,N_3506,N_4717);
xor U9055 (N_9055,N_4302,N_3725);
nand U9056 (N_9056,N_4327,N_6118);
and U9057 (N_9057,N_6228,N_5309);
xor U9058 (N_9058,N_4319,N_5152);
and U9059 (N_9059,N_5305,N_4330);
nand U9060 (N_9060,N_4298,N_4017);
nor U9061 (N_9061,N_4486,N_3593);
xor U9062 (N_9062,N_5047,N_4258);
xnor U9063 (N_9063,N_6214,N_6191);
xnor U9064 (N_9064,N_3376,N_5789);
nor U9065 (N_9065,N_6167,N_3248);
nand U9066 (N_9066,N_5433,N_5409);
xor U9067 (N_9067,N_4068,N_5186);
xor U9068 (N_9068,N_5693,N_3364);
nand U9069 (N_9069,N_3723,N_4534);
and U9070 (N_9070,N_5696,N_4180);
xor U9071 (N_9071,N_3860,N_3881);
or U9072 (N_9072,N_6148,N_3692);
and U9073 (N_9073,N_6108,N_5267);
xnor U9074 (N_9074,N_4947,N_5633);
nand U9075 (N_9075,N_3970,N_3890);
xor U9076 (N_9076,N_3609,N_6129);
xnor U9077 (N_9077,N_5367,N_4721);
xnor U9078 (N_9078,N_3669,N_3257);
nand U9079 (N_9079,N_3587,N_4181);
nor U9080 (N_9080,N_3668,N_4179);
or U9081 (N_9081,N_4786,N_5365);
nor U9082 (N_9082,N_4682,N_5788);
xor U9083 (N_9083,N_3478,N_4775);
nand U9084 (N_9084,N_3870,N_5965);
xor U9085 (N_9085,N_3360,N_4604);
or U9086 (N_9086,N_5569,N_5201);
and U9087 (N_9087,N_4641,N_5378);
xor U9088 (N_9088,N_6043,N_3871);
xor U9089 (N_9089,N_4122,N_5911);
and U9090 (N_9090,N_4222,N_3856);
nor U9091 (N_9091,N_3343,N_3624);
nor U9092 (N_9092,N_5502,N_5852);
nor U9093 (N_9093,N_6217,N_6094);
or U9094 (N_9094,N_4416,N_5326);
and U9095 (N_9095,N_5943,N_5740);
nand U9096 (N_9096,N_5254,N_6018);
nor U9097 (N_9097,N_5121,N_4338);
and U9098 (N_9098,N_4845,N_5758);
and U9099 (N_9099,N_3228,N_4285);
and U9100 (N_9100,N_3891,N_6052);
and U9101 (N_9101,N_5425,N_5214);
and U9102 (N_9102,N_4703,N_4156);
nand U9103 (N_9103,N_5389,N_4202);
nor U9104 (N_9104,N_4839,N_3126);
or U9105 (N_9105,N_5013,N_3240);
nand U9106 (N_9106,N_4636,N_6151);
or U9107 (N_9107,N_5543,N_5326);
and U9108 (N_9108,N_5652,N_4111);
or U9109 (N_9109,N_5109,N_5651);
nor U9110 (N_9110,N_4380,N_5658);
nand U9111 (N_9111,N_4453,N_3747);
or U9112 (N_9112,N_4573,N_4523);
or U9113 (N_9113,N_5040,N_5596);
nor U9114 (N_9114,N_4425,N_5585);
nand U9115 (N_9115,N_5932,N_3589);
and U9116 (N_9116,N_4051,N_5184);
and U9117 (N_9117,N_5337,N_5795);
nor U9118 (N_9118,N_5607,N_5116);
or U9119 (N_9119,N_6024,N_4584);
nor U9120 (N_9120,N_3487,N_4120);
or U9121 (N_9121,N_4392,N_5290);
and U9122 (N_9122,N_5445,N_3540);
and U9123 (N_9123,N_3947,N_4274);
and U9124 (N_9124,N_4029,N_3990);
or U9125 (N_9125,N_3678,N_4940);
xnor U9126 (N_9126,N_3906,N_4098);
nor U9127 (N_9127,N_4079,N_4714);
nand U9128 (N_9128,N_4126,N_4156);
nand U9129 (N_9129,N_5714,N_4326);
xor U9130 (N_9130,N_4276,N_5386);
nor U9131 (N_9131,N_3657,N_6090);
nand U9132 (N_9132,N_4563,N_5426);
xor U9133 (N_9133,N_6025,N_4241);
and U9134 (N_9134,N_5980,N_3633);
xnor U9135 (N_9135,N_3733,N_6132);
or U9136 (N_9136,N_3390,N_3263);
and U9137 (N_9137,N_6015,N_4883);
nand U9138 (N_9138,N_4420,N_4302);
xor U9139 (N_9139,N_5081,N_4916);
nor U9140 (N_9140,N_3716,N_5280);
or U9141 (N_9141,N_3326,N_4588);
nor U9142 (N_9142,N_4003,N_3903);
xor U9143 (N_9143,N_3305,N_3811);
nor U9144 (N_9144,N_3958,N_3904);
xor U9145 (N_9145,N_5095,N_3191);
nor U9146 (N_9146,N_4482,N_6067);
or U9147 (N_9147,N_4787,N_5794);
nor U9148 (N_9148,N_5966,N_4007);
or U9149 (N_9149,N_4598,N_4975);
xnor U9150 (N_9150,N_6233,N_5582);
xor U9151 (N_9151,N_5960,N_6156);
or U9152 (N_9152,N_4723,N_4763);
nor U9153 (N_9153,N_3623,N_4073);
and U9154 (N_9154,N_5302,N_3380);
xor U9155 (N_9155,N_4241,N_3264);
xor U9156 (N_9156,N_6080,N_4846);
xor U9157 (N_9157,N_5081,N_4731);
nor U9158 (N_9158,N_4789,N_5744);
and U9159 (N_9159,N_4506,N_3244);
xor U9160 (N_9160,N_4430,N_3987);
xnor U9161 (N_9161,N_4332,N_3135);
and U9162 (N_9162,N_4938,N_4019);
nor U9163 (N_9163,N_5855,N_4519);
or U9164 (N_9164,N_5992,N_5431);
nor U9165 (N_9165,N_3664,N_3555);
and U9166 (N_9166,N_3150,N_4408);
nand U9167 (N_9167,N_4669,N_5639);
nand U9168 (N_9168,N_3616,N_4781);
or U9169 (N_9169,N_3825,N_3208);
nor U9170 (N_9170,N_5299,N_3745);
xnor U9171 (N_9171,N_5480,N_3477);
nor U9172 (N_9172,N_3457,N_3572);
nor U9173 (N_9173,N_5220,N_5896);
or U9174 (N_9174,N_5111,N_5473);
or U9175 (N_9175,N_5147,N_6196);
nor U9176 (N_9176,N_3758,N_5424);
and U9177 (N_9177,N_3153,N_3892);
or U9178 (N_9178,N_5793,N_3739);
xor U9179 (N_9179,N_5084,N_5037);
and U9180 (N_9180,N_4569,N_6083);
nand U9181 (N_9181,N_4247,N_3638);
and U9182 (N_9182,N_3150,N_4669);
nand U9183 (N_9183,N_4264,N_6111);
nand U9184 (N_9184,N_6153,N_3300);
and U9185 (N_9185,N_5851,N_5094);
or U9186 (N_9186,N_5444,N_5771);
or U9187 (N_9187,N_4228,N_5207);
xor U9188 (N_9188,N_5794,N_4418);
or U9189 (N_9189,N_3987,N_4954);
and U9190 (N_9190,N_5342,N_5907);
nor U9191 (N_9191,N_3413,N_5693);
nand U9192 (N_9192,N_5272,N_5218);
or U9193 (N_9193,N_5353,N_5208);
xor U9194 (N_9194,N_6101,N_5798);
xor U9195 (N_9195,N_4133,N_6178);
xnor U9196 (N_9196,N_5584,N_3677);
nor U9197 (N_9197,N_3885,N_6185);
nand U9198 (N_9198,N_3685,N_4458);
nor U9199 (N_9199,N_4796,N_4057);
nand U9200 (N_9200,N_4966,N_4587);
xnor U9201 (N_9201,N_5513,N_3969);
xnor U9202 (N_9202,N_6100,N_4166);
or U9203 (N_9203,N_4411,N_4812);
or U9204 (N_9204,N_4770,N_6197);
and U9205 (N_9205,N_4401,N_3663);
xor U9206 (N_9206,N_5702,N_6177);
and U9207 (N_9207,N_3870,N_4660);
nand U9208 (N_9208,N_6070,N_6006);
nor U9209 (N_9209,N_3263,N_3341);
nor U9210 (N_9210,N_3210,N_6135);
or U9211 (N_9211,N_4442,N_4802);
or U9212 (N_9212,N_5497,N_4571);
and U9213 (N_9213,N_3288,N_5576);
or U9214 (N_9214,N_5551,N_3578);
nand U9215 (N_9215,N_4878,N_4317);
nand U9216 (N_9216,N_3225,N_3539);
xnor U9217 (N_9217,N_3434,N_5258);
and U9218 (N_9218,N_6097,N_4038);
nor U9219 (N_9219,N_3925,N_3142);
or U9220 (N_9220,N_3426,N_3473);
xnor U9221 (N_9221,N_4583,N_5724);
nor U9222 (N_9222,N_3417,N_5901);
and U9223 (N_9223,N_3482,N_4976);
nand U9224 (N_9224,N_4085,N_3870);
xnor U9225 (N_9225,N_5284,N_3752);
nand U9226 (N_9226,N_3182,N_3235);
and U9227 (N_9227,N_3295,N_3962);
or U9228 (N_9228,N_6137,N_4407);
or U9229 (N_9229,N_4853,N_4856);
nand U9230 (N_9230,N_5103,N_3514);
xnor U9231 (N_9231,N_4688,N_3319);
nor U9232 (N_9232,N_5323,N_3268);
or U9233 (N_9233,N_5295,N_5420);
or U9234 (N_9234,N_4051,N_4057);
and U9235 (N_9235,N_4423,N_5078);
or U9236 (N_9236,N_5295,N_5155);
nand U9237 (N_9237,N_3332,N_4208);
nand U9238 (N_9238,N_3525,N_5277);
nor U9239 (N_9239,N_6147,N_3676);
and U9240 (N_9240,N_5242,N_5018);
or U9241 (N_9241,N_6217,N_5028);
nor U9242 (N_9242,N_3420,N_5739);
xnor U9243 (N_9243,N_5415,N_5255);
nand U9244 (N_9244,N_5504,N_4380);
nand U9245 (N_9245,N_5638,N_4948);
xor U9246 (N_9246,N_5819,N_5436);
xnor U9247 (N_9247,N_4668,N_5769);
xor U9248 (N_9248,N_3291,N_3414);
and U9249 (N_9249,N_5890,N_5983);
or U9250 (N_9250,N_3290,N_4260);
nor U9251 (N_9251,N_5949,N_5753);
nand U9252 (N_9252,N_3436,N_4481);
nor U9253 (N_9253,N_6091,N_5812);
and U9254 (N_9254,N_5445,N_5092);
and U9255 (N_9255,N_4909,N_5203);
xnor U9256 (N_9256,N_4073,N_3718);
xor U9257 (N_9257,N_3374,N_5334);
xor U9258 (N_9258,N_3496,N_4204);
nand U9259 (N_9259,N_5072,N_6107);
xor U9260 (N_9260,N_3499,N_3246);
or U9261 (N_9261,N_6164,N_5890);
and U9262 (N_9262,N_3855,N_4989);
nor U9263 (N_9263,N_3848,N_5371);
xor U9264 (N_9264,N_3449,N_4818);
and U9265 (N_9265,N_4262,N_5372);
xor U9266 (N_9266,N_4760,N_4884);
nor U9267 (N_9267,N_3422,N_4716);
or U9268 (N_9268,N_5289,N_5151);
nor U9269 (N_9269,N_4739,N_3868);
and U9270 (N_9270,N_4388,N_3947);
nor U9271 (N_9271,N_5534,N_3148);
and U9272 (N_9272,N_5576,N_3664);
xnor U9273 (N_9273,N_5713,N_4206);
xor U9274 (N_9274,N_4063,N_5618);
and U9275 (N_9275,N_3767,N_5769);
or U9276 (N_9276,N_4524,N_5311);
or U9277 (N_9277,N_6128,N_3698);
and U9278 (N_9278,N_3159,N_6021);
nand U9279 (N_9279,N_3150,N_3196);
and U9280 (N_9280,N_4314,N_6185);
and U9281 (N_9281,N_5035,N_6183);
nand U9282 (N_9282,N_4738,N_5028);
nand U9283 (N_9283,N_6109,N_5036);
and U9284 (N_9284,N_5672,N_4402);
xor U9285 (N_9285,N_4612,N_5432);
xor U9286 (N_9286,N_4592,N_3294);
and U9287 (N_9287,N_5314,N_5172);
or U9288 (N_9288,N_3900,N_4700);
or U9289 (N_9289,N_4464,N_4142);
nor U9290 (N_9290,N_5963,N_6129);
and U9291 (N_9291,N_5313,N_5240);
nor U9292 (N_9292,N_3199,N_4947);
xor U9293 (N_9293,N_5581,N_5214);
nand U9294 (N_9294,N_4857,N_6118);
xnor U9295 (N_9295,N_4454,N_5587);
xnor U9296 (N_9296,N_4949,N_5294);
nand U9297 (N_9297,N_4738,N_3993);
nand U9298 (N_9298,N_4296,N_3160);
or U9299 (N_9299,N_3319,N_3557);
xor U9300 (N_9300,N_4714,N_4779);
and U9301 (N_9301,N_3329,N_3206);
nand U9302 (N_9302,N_6062,N_4863);
nor U9303 (N_9303,N_3881,N_6093);
nand U9304 (N_9304,N_5284,N_4038);
nor U9305 (N_9305,N_4421,N_5677);
nand U9306 (N_9306,N_5976,N_4822);
and U9307 (N_9307,N_3214,N_4616);
nor U9308 (N_9308,N_5844,N_5517);
or U9309 (N_9309,N_5714,N_5962);
xnor U9310 (N_9310,N_3354,N_5442);
xnor U9311 (N_9311,N_4082,N_5380);
nor U9312 (N_9312,N_4497,N_4333);
xor U9313 (N_9313,N_4893,N_4861);
nor U9314 (N_9314,N_3285,N_3231);
xor U9315 (N_9315,N_6205,N_3150);
or U9316 (N_9316,N_5767,N_3586);
or U9317 (N_9317,N_5240,N_4091);
xor U9318 (N_9318,N_5073,N_4625);
and U9319 (N_9319,N_4180,N_3446);
xnor U9320 (N_9320,N_4235,N_4581);
xor U9321 (N_9321,N_4545,N_3309);
xnor U9322 (N_9322,N_4109,N_3728);
nor U9323 (N_9323,N_4934,N_5724);
or U9324 (N_9324,N_5461,N_5509);
nor U9325 (N_9325,N_6019,N_4837);
nand U9326 (N_9326,N_3372,N_4074);
nor U9327 (N_9327,N_4203,N_3572);
and U9328 (N_9328,N_6136,N_3453);
and U9329 (N_9329,N_5668,N_4368);
and U9330 (N_9330,N_3570,N_6182);
nand U9331 (N_9331,N_6088,N_3343);
or U9332 (N_9332,N_5398,N_4377);
nor U9333 (N_9333,N_5612,N_5647);
nand U9334 (N_9334,N_4098,N_5460);
and U9335 (N_9335,N_4610,N_5943);
xor U9336 (N_9336,N_6165,N_6063);
nor U9337 (N_9337,N_3530,N_5777);
and U9338 (N_9338,N_5200,N_4708);
or U9339 (N_9339,N_4176,N_4392);
or U9340 (N_9340,N_4198,N_3558);
and U9341 (N_9341,N_5754,N_5667);
and U9342 (N_9342,N_4463,N_4917);
nor U9343 (N_9343,N_3864,N_6073);
nor U9344 (N_9344,N_4318,N_6039);
nor U9345 (N_9345,N_4788,N_5821);
and U9346 (N_9346,N_3514,N_3198);
or U9347 (N_9347,N_4653,N_5871);
nor U9348 (N_9348,N_4654,N_5598);
nor U9349 (N_9349,N_4336,N_4523);
nand U9350 (N_9350,N_4291,N_4658);
and U9351 (N_9351,N_4416,N_5162);
xnor U9352 (N_9352,N_4128,N_4078);
xor U9353 (N_9353,N_5253,N_5463);
xor U9354 (N_9354,N_6067,N_3687);
and U9355 (N_9355,N_4506,N_5696);
xor U9356 (N_9356,N_5511,N_4942);
and U9357 (N_9357,N_4295,N_5355);
nor U9358 (N_9358,N_6188,N_3933);
or U9359 (N_9359,N_4342,N_5762);
nand U9360 (N_9360,N_6164,N_3270);
and U9361 (N_9361,N_3595,N_4236);
and U9362 (N_9362,N_3374,N_4167);
nor U9363 (N_9363,N_5360,N_5180);
nand U9364 (N_9364,N_4408,N_4417);
or U9365 (N_9365,N_3551,N_3265);
nor U9366 (N_9366,N_3645,N_3635);
xnor U9367 (N_9367,N_5468,N_4459);
and U9368 (N_9368,N_5217,N_5095);
and U9369 (N_9369,N_3455,N_5294);
and U9370 (N_9370,N_5703,N_3983);
or U9371 (N_9371,N_4031,N_3224);
nand U9372 (N_9372,N_4754,N_5152);
nor U9373 (N_9373,N_4104,N_3666);
or U9374 (N_9374,N_3404,N_4616);
nand U9375 (N_9375,N_6540,N_7812);
nor U9376 (N_9376,N_8742,N_8785);
and U9377 (N_9377,N_8285,N_7208);
or U9378 (N_9378,N_7556,N_6425);
or U9379 (N_9379,N_7927,N_7007);
and U9380 (N_9380,N_8160,N_8954);
nand U9381 (N_9381,N_8780,N_6824);
nand U9382 (N_9382,N_7575,N_7937);
and U9383 (N_9383,N_7380,N_7497);
and U9384 (N_9384,N_8173,N_8003);
xor U9385 (N_9385,N_7229,N_6317);
nor U9386 (N_9386,N_9187,N_8210);
xor U9387 (N_9387,N_8922,N_6850);
nor U9388 (N_9388,N_8429,N_7829);
nor U9389 (N_9389,N_8759,N_9205);
xor U9390 (N_9390,N_6823,N_6876);
nand U9391 (N_9391,N_7475,N_7421);
xnor U9392 (N_9392,N_9256,N_8907);
nor U9393 (N_9393,N_7234,N_9183);
nor U9394 (N_9394,N_8323,N_7018);
and U9395 (N_9395,N_8573,N_8821);
nor U9396 (N_9396,N_7981,N_6562);
xnor U9397 (N_9397,N_7117,N_6928);
and U9398 (N_9398,N_8225,N_8622);
nand U9399 (N_9399,N_8478,N_8257);
nor U9400 (N_9400,N_9363,N_7797);
and U9401 (N_9401,N_9270,N_6854);
nor U9402 (N_9402,N_7818,N_8050);
xnor U9403 (N_9403,N_7088,N_6874);
xnor U9404 (N_9404,N_8259,N_8949);
or U9405 (N_9405,N_6409,N_9352);
or U9406 (N_9406,N_8692,N_9282);
or U9407 (N_9407,N_6461,N_6713);
nor U9408 (N_9408,N_9218,N_8807);
and U9409 (N_9409,N_8871,N_8006);
and U9410 (N_9410,N_7305,N_6313);
nor U9411 (N_9411,N_8670,N_7557);
nor U9412 (N_9412,N_7591,N_8794);
nand U9413 (N_9413,N_7342,N_7307);
nor U9414 (N_9414,N_6894,N_8467);
nand U9415 (N_9415,N_9075,N_9334);
nand U9416 (N_9416,N_6256,N_9016);
and U9417 (N_9417,N_7989,N_8168);
xor U9418 (N_9418,N_9144,N_7075);
and U9419 (N_9419,N_6529,N_7677);
nor U9420 (N_9420,N_7185,N_7770);
and U9421 (N_9421,N_6655,N_7359);
nor U9422 (N_9422,N_6950,N_8343);
and U9423 (N_9423,N_7548,N_8081);
or U9424 (N_9424,N_6706,N_7984);
nand U9425 (N_9425,N_8613,N_8514);
and U9426 (N_9426,N_7217,N_8798);
or U9427 (N_9427,N_7531,N_8602);
xor U9428 (N_9428,N_6323,N_7791);
xor U9429 (N_9429,N_6347,N_9152);
nor U9430 (N_9430,N_9370,N_6653);
nand U9431 (N_9431,N_7175,N_6276);
nand U9432 (N_9432,N_6818,N_7616);
and U9433 (N_9433,N_9090,N_6756);
nor U9434 (N_9434,N_8576,N_9357);
and U9435 (N_9435,N_7333,N_7335);
and U9436 (N_9436,N_6644,N_8647);
or U9437 (N_9437,N_8087,N_7317);
xor U9438 (N_9438,N_8452,N_6384);
nand U9439 (N_9439,N_8543,N_7923);
nand U9440 (N_9440,N_9247,N_6433);
xnor U9441 (N_9441,N_6365,N_8362);
or U9442 (N_9442,N_6424,N_8273);
nor U9443 (N_9443,N_7733,N_7336);
nor U9444 (N_9444,N_6331,N_6572);
or U9445 (N_9445,N_7841,N_7426);
xnor U9446 (N_9446,N_8558,N_8062);
nand U9447 (N_9447,N_8611,N_7360);
nor U9448 (N_9448,N_7951,N_6666);
and U9449 (N_9449,N_8022,N_6481);
and U9450 (N_9450,N_8275,N_8769);
or U9451 (N_9451,N_7111,N_6863);
nand U9452 (N_9452,N_6661,N_8487);
or U9453 (N_9453,N_7119,N_8339);
xnor U9454 (N_9454,N_6807,N_6960);
xor U9455 (N_9455,N_7718,N_7169);
nor U9456 (N_9456,N_6813,N_8928);
xor U9457 (N_9457,N_8408,N_9306);
and U9458 (N_9458,N_8792,N_8412);
or U9459 (N_9459,N_6889,N_8474);
xnor U9460 (N_9460,N_8953,N_7022);
nor U9461 (N_9461,N_7938,N_7459);
xnor U9462 (N_9462,N_8265,N_8315);
and U9463 (N_9463,N_6916,N_8975);
xnor U9464 (N_9464,N_7914,N_9325);
and U9465 (N_9465,N_6286,N_6785);
or U9466 (N_9466,N_7936,N_7237);
nor U9467 (N_9467,N_7757,N_6257);
or U9468 (N_9468,N_7184,N_8032);
and U9469 (N_9469,N_9131,N_7982);
or U9470 (N_9470,N_9103,N_7104);
and U9471 (N_9471,N_7279,N_8182);
xor U9472 (N_9472,N_8040,N_6386);
and U9473 (N_9473,N_9177,N_7810);
xor U9474 (N_9474,N_9318,N_9176);
xor U9475 (N_9475,N_8970,N_6367);
and U9476 (N_9476,N_8974,N_8246);
nor U9477 (N_9477,N_6322,N_7775);
nand U9478 (N_9478,N_7940,N_6455);
or U9479 (N_9479,N_7407,N_6619);
xnor U9480 (N_9480,N_8189,N_8528);
nand U9481 (N_9481,N_7446,N_9319);
nand U9482 (N_9482,N_7203,N_8069);
xor U9483 (N_9483,N_6279,N_6768);
nand U9484 (N_9484,N_7862,N_8112);
or U9485 (N_9485,N_7058,N_7245);
nand U9486 (N_9486,N_6571,N_6511);
xor U9487 (N_9487,N_7034,N_9088);
xnor U9488 (N_9488,N_6849,N_8674);
and U9489 (N_9489,N_6566,N_7482);
and U9490 (N_9490,N_7507,N_7894);
xnor U9491 (N_9491,N_6370,N_8608);
nand U9492 (N_9492,N_7837,N_9155);
xnor U9493 (N_9493,N_9219,N_8817);
and U9494 (N_9494,N_9055,N_8936);
and U9495 (N_9495,N_8373,N_7855);
or U9496 (N_9496,N_8144,N_7723);
and U9497 (N_9497,N_8034,N_8092);
nand U9498 (N_9498,N_8178,N_8462);
xor U9499 (N_9499,N_9367,N_8646);
or U9500 (N_9500,N_6938,N_7593);
nand U9501 (N_9501,N_6265,N_9287);
xnor U9502 (N_9502,N_7023,N_8014);
nor U9503 (N_9503,N_9126,N_9265);
and U9504 (N_9504,N_8902,N_8722);
xnor U9505 (N_9505,N_8012,N_7006);
nor U9506 (N_9506,N_9244,N_8959);
nand U9507 (N_9507,N_9006,N_6293);
and U9508 (N_9508,N_7352,N_6261);
nor U9509 (N_9509,N_9173,N_7182);
xor U9510 (N_9510,N_6995,N_6701);
xnor U9511 (N_9511,N_7639,N_9138);
nor U9512 (N_9512,N_7172,N_7684);
nand U9513 (N_9513,N_6589,N_8167);
xor U9514 (N_9514,N_6883,N_6593);
nor U9515 (N_9515,N_7216,N_7919);
nand U9516 (N_9516,N_8303,N_7496);
and U9517 (N_9517,N_8741,N_6518);
xnor U9518 (N_9518,N_8848,N_8630);
nor U9519 (N_9519,N_7364,N_6548);
xor U9520 (N_9520,N_6498,N_7188);
nand U9521 (N_9521,N_8453,N_8378);
and U9522 (N_9522,N_7271,N_7662);
nor U9523 (N_9523,N_7734,N_8753);
and U9524 (N_9524,N_6525,N_6369);
nor U9525 (N_9525,N_6395,N_8276);
and U9526 (N_9526,N_8901,N_8399);
or U9527 (N_9527,N_8481,N_8326);
xnor U9528 (N_9528,N_7632,N_6591);
nor U9529 (N_9529,N_8620,N_7994);
nor U9530 (N_9530,N_6885,N_7236);
nand U9531 (N_9531,N_8296,N_8464);
or U9532 (N_9532,N_9013,N_6774);
and U9533 (N_9533,N_7410,N_7577);
nand U9534 (N_9534,N_8508,N_8786);
nand U9535 (N_9535,N_8708,N_7338);
xor U9536 (N_9536,N_8396,N_8480);
nor U9537 (N_9537,N_6787,N_6899);
or U9538 (N_9538,N_6345,N_7000);
nand U9539 (N_9539,N_8238,N_6586);
and U9540 (N_9540,N_7976,N_8852);
nand U9541 (N_9541,N_9057,N_8213);
nor U9542 (N_9542,N_9214,N_6830);
nand U9543 (N_9543,N_7053,N_7758);
and U9544 (N_9544,N_7641,N_6259);
and U9545 (N_9545,N_6764,N_6321);
and U9546 (N_9546,N_8477,N_9317);
nor U9547 (N_9547,N_8079,N_9121);
and U9548 (N_9548,N_9250,N_8150);
nand U9549 (N_9549,N_9077,N_7732);
nand U9550 (N_9550,N_6658,N_8074);
xor U9551 (N_9551,N_6329,N_6640);
xnor U9552 (N_9552,N_9246,N_7462);
xnor U9553 (N_9553,N_7563,N_8253);
and U9554 (N_9554,N_8590,N_6762);
xor U9555 (N_9555,N_8230,N_7154);
xnor U9556 (N_9556,N_6746,N_7189);
and U9557 (N_9557,N_7397,N_6716);
and U9558 (N_9558,N_6297,N_7030);
nand U9559 (N_9559,N_7167,N_8952);
xnor U9560 (N_9560,N_8194,N_7032);
nor U9561 (N_9561,N_6426,N_6614);
xor U9562 (N_9562,N_7724,N_8130);
xnor U9563 (N_9563,N_8512,N_8998);
or U9564 (N_9564,N_8124,N_6350);
or U9565 (N_9565,N_9175,N_8117);
nor U9566 (N_9566,N_7588,N_7500);
nor U9567 (N_9567,N_7151,N_6973);
xor U9568 (N_9568,N_7879,N_8675);
nand U9569 (N_9569,N_9066,N_7534);
or U9570 (N_9570,N_6444,N_9178);
xor U9571 (N_9571,N_8199,N_6942);
nand U9572 (N_9572,N_9046,N_6929);
or U9573 (N_9573,N_8271,N_8393);
xor U9574 (N_9574,N_7078,N_7766);
or U9575 (N_9575,N_6576,N_7089);
and U9576 (N_9576,N_7781,N_8007);
and U9577 (N_9577,N_6336,N_8663);
nand U9578 (N_9578,N_7622,N_6616);
and U9579 (N_9579,N_9172,N_9115);
xnor U9580 (N_9580,N_7223,N_6523);
xor U9581 (N_9581,N_8603,N_6503);
or U9582 (N_9582,N_7045,N_7915);
nor U9583 (N_9583,N_7280,N_9231);
nor U9584 (N_9584,N_6393,N_8874);
nor U9585 (N_9585,N_6599,N_6631);
nand U9586 (N_9586,N_6325,N_6887);
xor U9587 (N_9587,N_8290,N_7828);
and U9588 (N_9588,N_7396,N_8418);
or U9589 (N_9589,N_8231,N_7767);
and U9590 (N_9590,N_6451,N_8267);
and U9591 (N_9591,N_8697,N_6811);
or U9592 (N_9592,N_6366,N_7739);
nor U9593 (N_9593,N_8320,N_6659);
or U9594 (N_9594,N_7564,N_7458);
or U9595 (N_9595,N_6790,N_6837);
nand U9596 (N_9596,N_8456,N_8234);
nor U9597 (N_9597,N_7587,N_7845);
and U9598 (N_9598,N_8472,N_6656);
nand U9599 (N_9599,N_7099,N_6888);
or U9600 (N_9600,N_6684,N_8245);
nand U9601 (N_9601,N_6860,N_7884);
or U9602 (N_9602,N_7387,N_7549);
nand U9603 (N_9603,N_6996,N_8374);
nor U9604 (N_9604,N_6538,N_7453);
nand U9605 (N_9605,N_8447,N_7491);
or U9606 (N_9606,N_8333,N_8933);
or U9607 (N_9607,N_8135,N_6568);
nor U9608 (N_9608,N_6549,N_8395);
or U9609 (N_9609,N_9264,N_6534);
or U9610 (N_9610,N_9258,N_6550);
and U9611 (N_9611,N_8502,N_9081);
or U9612 (N_9612,N_8162,N_9369);
nand U9613 (N_9613,N_8621,N_9327);
xor U9614 (N_9614,N_7647,N_7819);
and U9615 (N_9615,N_7744,N_6886);
nand U9616 (N_9616,N_9185,N_7823);
xnor U9617 (N_9617,N_7634,N_9161);
nand U9618 (N_9618,N_6980,N_6903);
nand U9619 (N_9619,N_8664,N_6630);
nor U9620 (N_9620,N_9192,N_8357);
xor U9621 (N_9621,N_9109,N_7560);
nor U9622 (N_9622,N_8927,N_9149);
or U9623 (N_9623,N_9275,N_7833);
xor U9624 (N_9624,N_6625,N_7553);
nor U9625 (N_9625,N_8018,N_9373);
xor U9626 (N_9626,N_8826,N_6439);
nor U9627 (N_9627,N_8485,N_8428);
or U9628 (N_9628,N_7076,N_8658);
nor U9629 (N_9629,N_6705,N_7404);
xor U9630 (N_9630,N_8053,N_7153);
xor U9631 (N_9631,N_7749,N_7660);
nor U9632 (N_9632,N_6979,N_7431);
and U9633 (N_9633,N_8574,N_7599);
and U9634 (N_9634,N_7691,N_7952);
xnor U9635 (N_9635,N_8945,N_8437);
or U9636 (N_9636,N_6800,N_7096);
or U9637 (N_9637,N_6877,N_6453);
xnor U9638 (N_9638,N_6397,N_7572);
nor U9639 (N_9639,N_7121,N_8700);
or U9640 (N_9640,N_8235,N_6810);
or U9641 (N_9641,N_8145,N_6855);
nor U9642 (N_9642,N_9251,N_7048);
nor U9643 (N_9643,N_7895,N_6871);
xor U9644 (N_9644,N_8356,N_6825);
nand U9645 (N_9645,N_7206,N_7195);
xnor U9646 (N_9646,N_9353,N_9293);
nor U9647 (N_9647,N_8873,N_9076);
nor U9648 (N_9648,N_7002,N_7017);
nand U9649 (N_9649,N_7853,N_9132);
nor U9650 (N_9650,N_7093,N_7737);
and U9651 (N_9651,N_8990,N_6688);
and U9652 (N_9652,N_9344,N_6612);
nand U9653 (N_9653,N_6275,N_7191);
xor U9654 (N_9654,N_7283,N_9233);
xnor U9655 (N_9655,N_8579,N_8035);
nor U9656 (N_9656,N_6896,N_8017);
and U9657 (N_9657,N_7255,N_7896);
nand U9658 (N_9658,N_9022,N_6387);
or U9659 (N_9659,N_7753,N_6624);
nor U9660 (N_9660,N_6700,N_6760);
and U9661 (N_9661,N_7343,N_8442);
xnor U9662 (N_9662,N_7941,N_6808);
nand U9663 (N_9663,N_8232,N_8370);
or U9664 (N_9664,N_8745,N_7081);
xnor U9665 (N_9665,N_6971,N_8771);
and U9666 (N_9666,N_7149,N_8483);
or U9667 (N_9667,N_8187,N_8261);
nand U9668 (N_9668,N_8942,N_9245);
nand U9669 (N_9669,N_6668,N_8777);
xor U9670 (N_9670,N_7028,N_6697);
and U9671 (N_9671,N_7820,N_7264);
or U9672 (N_9672,N_8416,N_8385);
and U9673 (N_9673,N_6250,N_6274);
nand U9674 (N_9674,N_7629,N_9010);
xnor U9675 (N_9675,N_7947,N_7207);
and U9676 (N_9676,N_7106,N_8283);
nor U9677 (N_9677,N_8388,N_7621);
nor U9678 (N_9678,N_8736,N_7510);
and U9679 (N_9679,N_9106,N_8986);
nor U9680 (N_9680,N_6835,N_7289);
or U9681 (N_9681,N_8762,N_8256);
and U9682 (N_9682,N_8037,N_7950);
nor U9683 (N_9683,N_7246,N_7685);
nand U9684 (N_9684,N_7406,N_9285);
nand U9685 (N_9685,N_8772,N_9223);
nand U9686 (N_9686,N_7922,N_7826);
and U9687 (N_9687,N_7526,N_7346);
xor U9688 (N_9688,N_7728,N_7012);
nand U9689 (N_9689,N_6907,N_7388);
nor U9690 (N_9690,N_9048,N_7558);
xnor U9691 (N_9691,N_8033,N_9295);
and U9692 (N_9692,N_8489,N_8822);
or U9693 (N_9693,N_6420,N_8754);
nor U9694 (N_9694,N_7657,N_8376);
xor U9695 (N_9695,N_9328,N_8095);
and U9696 (N_9696,N_9360,N_8318);
xor U9697 (N_9697,N_6744,N_7354);
and U9698 (N_9698,N_8828,N_7416);
nand U9699 (N_9699,N_7573,N_8248);
or U9700 (N_9700,N_8799,N_8240);
and U9701 (N_9701,N_6710,N_8750);
xor U9702 (N_9702,N_8043,N_6598);
nand U9703 (N_9703,N_8728,N_7466);
or U9704 (N_9704,N_7463,N_8152);
xnor U9705 (N_9705,N_7490,N_8363);
or U9706 (N_9706,N_8170,N_6958);
xor U9707 (N_9707,N_8098,N_9292);
or U9708 (N_9708,N_6326,N_8638);
nand U9709 (N_9709,N_8364,N_8681);
and U9710 (N_9710,N_9056,N_9020);
and U9711 (N_9711,N_6474,N_7921);
and U9712 (N_9712,N_9217,N_8650);
or U9713 (N_9713,N_8526,N_7130);
and U9714 (N_9714,N_7681,N_8841);
xor U9715 (N_9715,N_9080,N_6278);
xnor U9716 (N_9716,N_6704,N_7334);
or U9717 (N_9717,N_7693,N_9366);
xnor U9718 (N_9718,N_7257,N_8522);
nor U9719 (N_9719,N_7384,N_6398);
nand U9720 (N_9720,N_8748,N_7225);
xor U9721 (N_9721,N_9084,N_8787);
nor U9722 (N_9722,N_6969,N_9329);
or U9723 (N_9723,N_6314,N_7221);
nand U9724 (N_9724,N_8895,N_8500);
nand U9725 (N_9725,N_8476,N_6934);
xnor U9726 (N_9726,N_7265,N_6375);
nor U9727 (N_9727,N_6922,N_7583);
nor U9728 (N_9728,N_8354,N_7393);
nor U9729 (N_9729,N_7747,N_8091);
xnor U9730 (N_9730,N_6743,N_7874);
and U9731 (N_9731,N_7964,N_7610);
nor U9732 (N_9732,N_7779,N_9310);
or U9733 (N_9733,N_6324,N_6949);
or U9734 (N_9734,N_6878,N_7975);
nor U9735 (N_9735,N_7210,N_7570);
and U9736 (N_9736,N_7301,N_8131);
nand U9737 (N_9737,N_7051,N_8570);
nand U9738 (N_9738,N_7442,N_8561);
or U9739 (N_9739,N_6530,N_6812);
nor U9740 (N_9740,N_7049,N_8301);
and U9741 (N_9741,N_8156,N_8969);
nor U9742 (N_9742,N_6993,N_7485);
nand U9743 (N_9743,N_6795,N_6493);
nand U9744 (N_9744,N_8604,N_8133);
nor U9745 (N_9745,N_8571,N_7834);
or U9746 (N_9746,N_8185,N_8097);
nand U9747 (N_9747,N_8084,N_6703);
or U9748 (N_9748,N_6287,N_7899);
xnor U9749 (N_9749,N_7316,N_8801);
nor U9750 (N_9750,N_6904,N_6406);
and U9751 (N_9751,N_6479,N_8045);
xnor U9752 (N_9752,N_7418,N_8864);
and U9753 (N_9753,N_7174,N_7569);
nand U9754 (N_9754,N_8312,N_8094);
and U9755 (N_9755,N_9201,N_7555);
nand U9756 (N_9756,N_6959,N_9294);
or U9757 (N_9757,N_6590,N_7486);
or U9758 (N_9758,N_8101,N_8859);
and U9759 (N_9759,N_7376,N_8734);
or U9760 (N_9760,N_8585,N_7918);
xor U9761 (N_9761,N_7772,N_6569);
xnor U9762 (N_9762,N_6567,N_8494);
xor U9763 (N_9763,N_7576,N_7495);
nand U9764 (N_9764,N_8831,N_6999);
and U9765 (N_9765,N_9316,N_8950);
nor U9766 (N_9766,N_6266,N_9014);
nand U9767 (N_9767,N_7107,N_8744);
nor U9768 (N_9768,N_9044,N_7965);
or U9769 (N_9769,N_7551,N_7778);
nand U9770 (N_9770,N_8843,N_7525);
nand U9771 (N_9771,N_8606,N_9261);
and U9772 (N_9772,N_7315,N_6608);
xor U9773 (N_9773,N_7072,N_8431);
nand U9774 (N_9774,N_8054,N_8937);
nand U9775 (N_9775,N_6427,N_7532);
and U9776 (N_9776,N_8346,N_7243);
or U9777 (N_9777,N_9082,N_6463);
xnor U9778 (N_9778,N_7150,N_8816);
or U9779 (N_9779,N_9129,N_8776);
nand U9780 (N_9780,N_7699,N_8071);
nor U9781 (N_9781,N_7103,N_7726);
nand U9782 (N_9782,N_6291,N_7679);
xnor U9783 (N_9783,N_8118,N_7859);
nand U9784 (N_9784,N_7717,N_9335);
and U9785 (N_9785,N_9089,N_7291);
and U9786 (N_9786,N_7671,N_8375);
xnor U9787 (N_9787,N_9093,N_9359);
nor U9788 (N_9788,N_8732,N_9211);
and U9789 (N_9789,N_8183,N_8177);
nand U9790 (N_9790,N_6584,N_7358);
or U9791 (N_9791,N_7754,N_8938);
nand U9792 (N_9792,N_8890,N_7197);
or U9793 (N_9793,N_6497,N_6510);
xor U9794 (N_9794,N_8932,N_8121);
or U9795 (N_9795,N_6660,N_8731);
nand U9796 (N_9796,N_9012,N_9311);
nor U9797 (N_9797,N_7559,N_7323);
nor U9798 (N_9798,N_6798,N_8000);
xnor U9799 (N_9799,N_6844,N_8419);
nor U9800 (N_9800,N_6648,N_9001);
and U9801 (N_9801,N_6376,N_6263);
and U9802 (N_9802,N_9030,N_7613);
and U9803 (N_9803,N_7186,N_7592);
nand U9804 (N_9804,N_7155,N_8504);
nand U9805 (N_9805,N_7383,N_7454);
or U9806 (N_9806,N_8212,N_6303);
or U9807 (N_9807,N_8501,N_6681);
xor U9808 (N_9808,N_7057,N_7437);
and U9809 (N_9809,N_8262,N_6680);
nor U9810 (N_9810,N_7906,N_7313);
nand U9811 (N_9811,N_8490,N_6306);
and U9812 (N_9812,N_7957,N_7931);
and U9813 (N_9813,N_8401,N_8336);
nand U9814 (N_9814,N_6385,N_6817);
xnor U9815 (N_9815,N_6604,N_6438);
and U9816 (N_9816,N_8906,N_7585);
and U9817 (N_9817,N_7815,N_6643);
xor U9818 (N_9818,N_7807,N_9284);
xor U9819 (N_9819,N_6595,N_7962);
and U9820 (N_9820,N_7856,N_7109);
and U9821 (N_9821,N_7444,N_8779);
nor U9822 (N_9822,N_6416,N_6283);
and U9823 (N_9823,N_6752,N_8155);
nand U9824 (N_9824,N_6780,N_9162);
xnor U9825 (N_9825,N_9002,N_7303);
or U9826 (N_9826,N_7768,N_8313);
xnor U9827 (N_9827,N_8812,N_7501);
or U9828 (N_9828,N_7005,N_9193);
and U9829 (N_9829,N_8207,N_7318);
xnor U9830 (N_9830,N_8729,N_8499);
and U9831 (N_9831,N_8833,N_8115);
xnor U9832 (N_9832,N_7494,N_6985);
or U9833 (N_9833,N_6953,N_6272);
nand U9834 (N_9834,N_8090,N_6609);
and U9835 (N_9835,N_8589,N_8694);
and U9836 (N_9836,N_6948,N_7902);
and U9837 (N_9837,N_6946,N_7678);
nor U9838 (N_9838,N_7042,N_7706);
nor U9839 (N_9839,N_7220,N_7201);
nand U9840 (N_9840,N_8025,N_6448);
xnor U9841 (N_9841,N_6729,N_7287);
or U9842 (N_9842,N_7039,N_7127);
and U9843 (N_9843,N_7235,N_7566);
and U9844 (N_9844,N_8962,N_8683);
nor U9845 (N_9845,N_8580,N_8402);
or U9846 (N_9846,N_8122,N_9122);
nand U9847 (N_9847,N_9221,N_6341);
or U9848 (N_9848,N_7653,N_9150);
nand U9849 (N_9849,N_7873,N_8048);
or U9850 (N_9850,N_7771,N_7978);
xnor U9851 (N_9851,N_6723,N_6831);
or U9852 (N_9852,N_7435,N_7441);
and U9853 (N_9853,N_7344,N_6515);
nor U9854 (N_9854,N_6429,N_7649);
xnor U9855 (N_9855,N_6867,N_9099);
and U9856 (N_9856,N_9314,N_8104);
xor U9857 (N_9857,N_6925,N_8876);
and U9858 (N_9858,N_8846,N_7209);
or U9859 (N_9859,N_8545,N_6758);
and U9860 (N_9860,N_6763,N_6601);
and U9861 (N_9861,N_7980,N_7755);
and U9862 (N_9862,N_8068,N_7471);
or U9863 (N_9863,N_6841,N_7312);
and U9864 (N_9864,N_7350,N_7973);
nand U9865 (N_9865,N_8739,N_8988);
xor U9866 (N_9866,N_9153,N_6260);
nand U9867 (N_9867,N_8915,N_9179);
xor U9868 (N_9868,N_8426,N_8699);
nand U9869 (N_9869,N_8908,N_7783);
nand U9870 (N_9870,N_6486,N_6547);
nor U9871 (N_9871,N_8879,N_7741);
nand U9872 (N_9872,N_8317,N_9184);
and U9873 (N_9873,N_6298,N_7420);
nor U9874 (N_9874,N_6622,N_8912);
and U9875 (N_9875,N_7509,N_7190);
nand U9876 (N_9876,N_6920,N_7498);
nand U9877 (N_9877,N_7131,N_9313);
or U9878 (N_9878,N_6937,N_9039);
nor U9879 (N_9879,N_7436,N_6718);
nor U9880 (N_9880,N_8436,N_7545);
xnor U9881 (N_9881,N_8353,N_8171);
nor U9882 (N_9882,N_7809,N_9073);
or U9883 (N_9883,N_6603,N_6513);
nand U9884 (N_9884,N_6805,N_8767);
and U9885 (N_9885,N_9362,N_7219);
or U9886 (N_9886,N_8557,N_8180);
nor U9887 (N_9887,N_8909,N_8976);
nor U9888 (N_9888,N_8190,N_7108);
nor U9889 (N_9889,N_8463,N_9085);
nor U9890 (N_9890,N_6759,N_9116);
xor U9891 (N_9891,N_7596,N_9368);
nor U9892 (N_9892,N_8714,N_7911);
or U9893 (N_9893,N_7063,N_6797);
nor U9894 (N_9894,N_9337,N_7959);
nor U9895 (N_9895,N_6742,N_8880);
xor U9896 (N_9896,N_6819,N_6469);
and U9897 (N_9897,N_7543,N_7055);
nand U9898 (N_9898,N_8241,N_7087);
nor U9899 (N_9899,N_7925,N_7008);
xor U9900 (N_9900,N_7403,N_8784);
xnor U9901 (N_9901,N_8051,N_7886);
or U9902 (N_9902,N_8836,N_7817);
and U9903 (N_9903,N_6694,N_8208);
xor U9904 (N_9904,N_6543,N_9083);
nand U9905 (N_9905,N_8960,N_8390);
xor U9906 (N_9906,N_9358,N_7395);
xor U9907 (N_9907,N_8002,N_8586);
xor U9908 (N_9908,N_7405,N_8800);
xor U9909 (N_9909,N_8148,N_8427);
xnor U9910 (N_9910,N_8279,N_7579);
nor U9911 (N_9911,N_8868,N_8947);
nor U9912 (N_9912,N_8023,N_8319);
or U9913 (N_9913,N_7547,N_7773);
xnor U9914 (N_9914,N_8233,N_6647);
and U9915 (N_9915,N_7550,N_6777);
and U9916 (N_9916,N_6685,N_7648);
and U9917 (N_9917,N_9031,N_7796);
nor U9918 (N_9918,N_8920,N_8367);
nand U9919 (N_9919,N_7930,N_8584);
nor U9920 (N_9920,N_8321,N_6380);
xor U9921 (N_9921,N_6459,N_8582);
or U9922 (N_9922,N_7293,N_7689);
nor U9923 (N_9923,N_6931,N_8804);
and U9924 (N_9924,N_8689,N_7183);
or U9925 (N_9925,N_6452,N_7399);
or U9926 (N_9926,N_7077,N_6754);
nor U9927 (N_9927,N_6255,N_9034);
nor U9928 (N_9928,N_6349,N_8342);
nand U9929 (N_9929,N_8305,N_6882);
and U9930 (N_9930,N_7605,N_8929);
nor U9931 (N_9931,N_8311,N_6457);
xnor U9932 (N_9932,N_6602,N_6845);
nor U9933 (N_9933,N_6400,N_7998);
nor U9934 (N_9934,N_7637,N_8575);
xnor U9935 (N_9935,N_7328,N_8637);
and U9936 (N_9936,N_7419,N_8515);
xnor U9937 (N_9937,N_6596,N_8387);
and U9938 (N_9938,N_7541,N_8001);
nand U9939 (N_9939,N_9069,N_9181);
or U9940 (N_9940,N_6717,N_8605);
xor U9941 (N_9941,N_9148,N_7266);
xnor U9942 (N_9942,N_8384,N_8181);
and U9943 (N_9943,N_6578,N_7574);
nor U9944 (N_9944,N_8061,N_8626);
xor U9945 (N_9945,N_8517,N_6727);
and U9946 (N_9946,N_8803,N_8013);
and U9947 (N_9947,N_6908,N_7615);
xnor U9948 (N_9948,N_7337,N_8143);
xnor U9949 (N_9949,N_8632,N_7881);
and U9950 (N_9950,N_8805,N_7031);
and U9951 (N_9951,N_6657,N_7004);
and U9952 (N_9952,N_8982,N_7663);
xnor U9953 (N_9953,N_9209,N_8835);
nor U9954 (N_9954,N_8866,N_8544);
or U9955 (N_9955,N_6806,N_6490);
or U9956 (N_9956,N_7891,N_8548);
xnor U9957 (N_9957,N_9257,N_8147);
or U9958 (N_9958,N_6417,N_6552);
xnor U9959 (N_9959,N_8039,N_6449);
nor U9960 (N_9960,N_7133,N_9333);
xor U9961 (N_9961,N_7562,N_7363);
or U9962 (N_9962,N_8691,N_7644);
and U9963 (N_9963,N_7468,N_8935);
nor U9964 (N_9964,N_9305,N_6564);
xnor U9965 (N_9965,N_7793,N_9304);
or U9966 (N_9966,N_7479,N_6911);
nor U9967 (N_9967,N_8191,N_7378);
or U9968 (N_9968,N_9255,N_6337);
nand U9969 (N_9969,N_8684,N_6652);
nor U9970 (N_9970,N_6769,N_7230);
nand U9971 (N_9971,N_6446,N_6747);
nor U9972 (N_9972,N_8713,N_7214);
xor U9973 (N_9973,N_6956,N_6682);
or U9974 (N_9974,N_9018,N_7517);
or U9975 (N_9975,N_6332,N_7898);
nor U9976 (N_9976,N_9240,N_8434);
nor U9977 (N_9977,N_6765,N_7277);
nand U9978 (N_9978,N_7869,N_8614);
xnor U9979 (N_9979,N_7400,N_7224);
xor U9980 (N_9980,N_7180,N_8957);
nand U9981 (N_9981,N_7366,N_6771);
or U9982 (N_9982,N_8562,N_7170);
xnor U9983 (N_9983,N_8563,N_7092);
xnor U9984 (N_9984,N_7371,N_8934);
xnor U9985 (N_9985,N_7162,N_6264);
nand U9986 (N_9986,N_7086,N_9101);
xnor U9987 (N_9987,N_7054,N_9151);
nand U9988 (N_9988,N_6898,N_8698);
nand U9989 (N_9989,N_8216,N_6940);
nor U9990 (N_9990,N_6741,N_7114);
nor U9991 (N_9991,N_8616,N_9198);
xnor U9992 (N_9992,N_9224,N_6441);
nand U9993 (N_9993,N_6477,N_7798);
nor U9994 (N_9994,N_8910,N_8665);
xnor U9995 (N_9995,N_9052,N_8196);
or U9996 (N_9996,N_7268,N_8594);
xor U9997 (N_9997,N_8764,N_6402);
and U9998 (N_9998,N_8671,N_7847);
or U9999 (N_9999,N_7339,N_7200);
or U10000 (N_10000,N_6307,N_8639);
nand U10001 (N_10001,N_6773,N_7503);
and U10002 (N_10002,N_7595,N_7251);
nand U10003 (N_10003,N_7580,N_7392);
and U10004 (N_10004,N_8161,N_7676);
xor U10005 (N_10005,N_6289,N_6311);
or U10006 (N_10006,N_7890,N_7161);
and U10007 (N_10007,N_8830,N_6900);
or U10008 (N_10008,N_6649,N_8349);
nor U10009 (N_10009,N_7913,N_6753);
nand U10010 (N_10010,N_6683,N_6494);
nor U10011 (N_10011,N_6554,N_7381);
nand U10012 (N_10012,N_9104,N_6674);
xnor U10013 (N_10013,N_9272,N_7799);
xor U10014 (N_10014,N_9253,N_8701);
nand U10015 (N_10015,N_9051,N_8093);
nor U10016 (N_10016,N_6440,N_7609);
or U10017 (N_10017,N_8471,N_8838);
nor U10018 (N_10018,N_8781,N_8503);
and U10019 (N_10019,N_8810,N_8865);
and U10020 (N_10020,N_6342,N_7966);
and U10021 (N_10021,N_8818,N_8334);
or U10022 (N_10022,N_8382,N_9123);
nor U10023 (N_10023,N_8878,N_8226);
nand U10024 (N_10024,N_8597,N_8855);
and U10025 (N_10025,N_6319,N_7666);
and U10026 (N_10026,N_9100,N_7138);
nand U10027 (N_10027,N_6693,N_8289);
or U10028 (N_10028,N_6915,N_8716);
or U10029 (N_10029,N_7270,N_8082);
nand U10030 (N_10030,N_7527,N_6989);
nand U10031 (N_10031,N_8298,N_7871);
nor U10032 (N_10032,N_7838,N_8710);
nand U10033 (N_10033,N_8175,N_7953);
nand U10034 (N_10034,N_8588,N_6597);
and U10035 (N_10035,N_8725,N_6610);
or U10036 (N_10036,N_9182,N_6615);
xor U10037 (N_10037,N_7060,N_6975);
and U10038 (N_10038,N_8656,N_7473);
and U10039 (N_10039,N_8218,N_8309);
xnor U10040 (N_10040,N_6553,N_6633);
or U10041 (N_10041,N_6388,N_8530);
and U10042 (N_10042,N_7969,N_8851);
and U10043 (N_10043,N_7298,N_7863);
and U10044 (N_10044,N_7763,N_8887);
nand U10045 (N_10045,N_6277,N_7370);
nand U10046 (N_10046,N_7674,N_6695);
nand U10047 (N_10047,N_8657,N_7524);
nor U10048 (N_10048,N_8862,N_6262);
nor U10049 (N_10049,N_9300,N_7619);
xor U10050 (N_10050,N_8223,N_8724);
nor U10051 (N_10051,N_7990,N_6301);
and U10052 (N_10052,N_7630,N_6981);
nand U10053 (N_10053,N_8344,N_6528);
nor U10054 (N_10054,N_8380,N_7205);
nand U10055 (N_10055,N_9220,N_7173);
and U10056 (N_10056,N_7607,N_7661);
nor U10057 (N_10057,N_8536,N_6767);
and U10058 (N_10058,N_6532,N_6944);
and U10059 (N_10059,N_9248,N_7907);
or U10060 (N_10060,N_9043,N_7062);
or U10061 (N_10061,N_8292,N_7105);
and U10062 (N_10062,N_7148,N_9134);
xnor U10063 (N_10063,N_7697,N_7253);
nor U10064 (N_10064,N_8711,N_7999);
nor U10065 (N_10065,N_7084,N_8397);
or U10066 (N_10066,N_9191,N_7286);
xor U10067 (N_10067,N_7083,N_6374);
nor U10068 (N_10068,N_6910,N_7288);
and U10069 (N_10069,N_7375,N_7033);
and U10070 (N_10070,N_7272,N_7704);
xnor U10071 (N_10071,N_8703,N_6565);
xor U10072 (N_10072,N_8527,N_6519);
and U10073 (N_10073,N_9307,N_7233);
nor U10074 (N_10074,N_7159,N_6628);
nor U10075 (N_10075,N_7518,N_8202);
xnor U10076 (N_10076,N_9354,N_6390);
nor U10077 (N_10077,N_8219,N_9035);
nand U10078 (N_10078,N_7261,N_6536);
xor U10079 (N_10079,N_7977,N_7882);
nor U10080 (N_10080,N_6502,N_8823);
xor U10081 (N_10081,N_8789,N_6581);
xor U10082 (N_10082,N_8892,N_8154);
or U10083 (N_10083,N_6853,N_7617);
nand U10084 (N_10084,N_8894,N_9137);
xnor U10085 (N_10085,N_8310,N_9062);
and U10086 (N_10086,N_7842,N_8391);
nand U10087 (N_10087,N_6379,N_6983);
and U10088 (N_10088,N_6719,N_7460);
or U10089 (N_10089,N_7228,N_6587);
and U10090 (N_10090,N_7983,N_8972);
nor U10091 (N_10091,N_9068,N_8111);
xor U10092 (N_10092,N_7512,N_8560);
nand U10093 (N_10093,N_8591,N_8565);
and U10094 (N_10094,N_9365,N_8795);
nor U10095 (N_10095,N_9267,N_8497);
xnor U10096 (N_10096,N_8020,N_6354);
nor U10097 (N_10097,N_6917,N_6924);
nor U10098 (N_10098,N_7451,N_8755);
and U10099 (N_10099,N_7581,N_6890);
or U10100 (N_10100,N_9237,N_9263);
nor U10101 (N_10101,N_7719,N_7589);
and U10102 (N_10102,N_7357,N_8718);
and U10103 (N_10103,N_6802,N_8829);
xnor U10104 (N_10104,N_8242,N_8981);
and U10105 (N_10105,N_7785,N_9338);
or U10106 (N_10106,N_7025,N_7263);
xnor U10107 (N_10107,N_7521,N_6611);
nor U10108 (N_10108,N_7912,N_9283);
nor U10109 (N_10109,N_8108,N_6932);
xnor U10110 (N_10110,N_7920,N_9324);
nand U10111 (N_10111,N_8433,N_7612);
xnor U10112 (N_10112,N_6761,N_7854);
and U10113 (N_10113,N_9059,N_7349);
or U10114 (N_10114,N_9297,N_8371);
nand U10115 (N_10115,N_7456,N_8631);
or U10116 (N_10116,N_8943,N_7571);
nand U10117 (N_10117,N_8046,N_8324);
and U10118 (N_10118,N_8752,N_6654);
nand U10119 (N_10119,N_9308,N_6299);
and U10120 (N_10120,N_8192,N_7852);
and U10121 (N_10121,N_7836,N_6383);
and U10122 (N_10122,N_6308,N_7887);
nand U10123 (N_10123,N_6373,N_9259);
xnor U10124 (N_10124,N_8404,N_7187);
or U10125 (N_10125,N_6282,N_8550);
and U10126 (N_10126,N_8559,N_7068);
xnor U10127 (N_10127,N_6789,N_7278);
xor U10128 (N_10128,N_8457,N_7604);
nand U10129 (N_10129,N_7046,N_9036);
or U10130 (N_10130,N_7445,N_8883);
nor U10131 (N_10131,N_8793,N_8930);
nand U10132 (N_10132,N_7536,N_7904);
nor U10133 (N_10133,N_8535,N_8856);
nor U10134 (N_10134,N_7059,N_8662);
nand U10135 (N_10135,N_9026,N_8641);
or U10136 (N_10136,N_9374,N_6353);
xnor U10137 (N_10137,N_8286,N_9028);
nand U10138 (N_10138,N_7163,N_6467);
nor U10139 (N_10139,N_8272,N_8400);
or U10140 (N_10140,N_9213,N_6731);
or U10141 (N_10141,N_8666,N_7274);
nand U10142 (N_10142,N_8524,N_9202);
xor U10143 (N_10143,N_8839,N_7248);
xor U10144 (N_10144,N_8475,N_6634);
and U10145 (N_10145,N_8819,N_8761);
and U10146 (N_10146,N_7825,N_7877);
nor U10147 (N_10147,N_7567,N_8540);
nand U10148 (N_10148,N_6304,N_6936);
or U10149 (N_10149,N_6394,N_6560);
and U10150 (N_10150,N_6378,N_7422);
xor U10151 (N_10151,N_6755,N_6318);
xnor U10152 (N_10152,N_8338,N_7014);
xor U10153 (N_10153,N_6781,N_6483);
nor U10154 (N_10154,N_9145,N_7168);
nand U10155 (N_10155,N_6642,N_6281);
nand U10156 (N_10156,N_8410,N_8847);
or U10157 (N_10157,N_7729,N_7425);
nor U10158 (N_10158,N_8599,N_7124);
nand U10159 (N_10159,N_6672,N_6858);
or U10160 (N_10160,N_7320,N_6698);
nor U10161 (N_10161,N_9011,N_9356);
nand U10162 (N_10162,N_9078,N_7750);
or U10163 (N_10163,N_8297,N_6507);
nor U10164 (N_10164,N_8749,N_7910);
and U10165 (N_10165,N_7627,N_8409);
nor U10166 (N_10166,N_8567,N_8653);
xnor U10167 (N_10167,N_8243,N_6820);
and U10168 (N_10168,N_8625,N_7394);
nor U10169 (N_10169,N_8454,N_7821);
xnor U10170 (N_10170,N_6921,N_8513);
and U10171 (N_10171,N_8209,N_6372);
xnor U10172 (N_10172,N_6456,N_7652);
xor U10173 (N_10173,N_8174,N_8158);
xor U10174 (N_10174,N_9190,N_7708);
xnor U10175 (N_10175,N_7198,N_8853);
nand U10176 (N_10176,N_8941,N_6865);
and U10177 (N_10177,N_6381,N_8005);
and U10178 (N_10178,N_7244,N_6846);
or U10179 (N_10179,N_6962,N_6933);
nor U10180 (N_10180,N_6558,N_9047);
and U10181 (N_10181,N_9041,N_9303);
nor U10182 (N_10182,N_6253,N_8723);
nor U10183 (N_10183,N_7368,N_7933);
xor U10184 (N_10184,N_7179,N_8142);
or U10185 (N_10185,N_9336,N_8963);
or U10186 (N_10186,N_8973,N_9208);
or U10187 (N_10187,N_9096,N_8989);
nor U10188 (N_10188,N_8126,N_8444);
nand U10189 (N_10189,N_8556,N_6645);
and U10190 (N_10190,N_7584,N_7669);
or U10191 (N_10191,N_7626,N_9215);
nand U10192 (N_10192,N_9114,N_7967);
nor U10193 (N_10193,N_6791,N_9322);
xnor U10194 (N_10194,N_6669,N_8533);
nand U10195 (N_10195,N_6517,N_8875);
nor U10196 (N_10196,N_7658,N_8619);
or U10197 (N_10197,N_7016,N_8123);
nor U10198 (N_10198,N_8331,N_6930);
or U10199 (N_10199,N_9021,N_8790);
and U10200 (N_10200,N_6363,N_7582);
nand U10201 (N_10201,N_6258,N_6505);
nor U10202 (N_10202,N_8900,N_7506);
xnor U10203 (N_10203,N_9112,N_8891);
nor U10204 (N_10204,N_9235,N_8308);
or U10205 (N_10205,N_8861,N_9299);
and U10206 (N_10206,N_7939,N_8352);
nand U10207 (N_10207,N_6403,N_7620);
nand U10208 (N_10208,N_6766,N_8473);
nor U10209 (N_10209,N_8541,N_8971);
xnor U10210 (N_10210,N_6535,N_6251);
or U10211 (N_10211,N_9033,N_7844);
xor U10212 (N_10212,N_7457,N_6296);
nor U10213 (N_10213,N_9227,N_7552);
and U10214 (N_10214,N_8076,N_6861);
nand U10215 (N_10215,N_8008,N_8651);
and U10216 (N_10216,N_7714,N_6522);
nor U10217 (N_10217,N_8863,N_7866);
xor U10218 (N_10218,N_6984,N_7811);
xnor U10219 (N_10219,N_8987,N_9280);
nor U10220 (N_10220,N_9019,N_7411);
xnor U10221 (N_10221,N_8643,N_9023);
nor U10222 (N_10222,N_6636,N_9107);
nand U10223 (N_10223,N_6667,N_6472);
nor U10224 (N_10224,N_8956,N_7867);
nand U10225 (N_10225,N_6864,N_7348);
and U10226 (N_10226,N_6784,N_6335);
nand U10227 (N_10227,N_7505,N_7254);
xnor U10228 (N_10228,N_7680,N_6926);
and U10229 (N_10229,N_7888,N_9351);
xnor U10230 (N_10230,N_6857,N_8629);
or U10231 (N_10231,N_6371,N_6405);
or U10232 (N_10232,N_8466,N_8469);
nand U10233 (N_10233,N_7667,N_7713);
nand U10234 (N_10234,N_6470,N_8146);
xor U10235 (N_10235,N_7705,N_7134);
or U10236 (N_10236,N_8488,N_7664);
or U10237 (N_10237,N_7211,N_6635);
nand U10238 (N_10238,N_8788,N_9119);
xor U10239 (N_10239,N_6651,N_9249);
xor U10240 (N_10240,N_8965,N_6852);
xor U10241 (N_10241,N_9323,N_8284);
nand U10242 (N_10242,N_7565,N_9160);
and U10243 (N_10243,N_6732,N_6712);
xor U10244 (N_10244,N_7192,N_8832);
and U10245 (N_10245,N_7743,N_6711);
and U10246 (N_10246,N_9053,N_8898);
nor U10247 (N_10247,N_8120,N_9207);
xor U10248 (N_10248,N_7492,N_7840);
and U10249 (N_10249,N_7600,N_7688);
nor U10250 (N_10250,N_7861,N_8669);
nor U10251 (N_10251,N_8041,N_6485);
nor U10252 (N_10252,N_7402,N_9060);
xnor U10253 (N_10253,N_8229,N_7472);
nand U10254 (N_10254,N_8015,N_7469);
or U10255 (N_10255,N_6735,N_6280);
and U10256 (N_10256,N_6750,N_8770);
and U10257 (N_10257,N_7929,N_8461);
nor U10258 (N_10258,N_6897,N_6952);
and U10259 (N_10259,N_7539,N_7935);
nand U10260 (N_10260,N_8307,N_6843);
xor U10261 (N_10261,N_8422,N_9125);
xnor U10262 (N_10262,N_7212,N_7765);
and U10263 (N_10263,N_8224,N_7777);
nor U10264 (N_10264,N_7157,N_8858);
nor U10265 (N_10265,N_7801,N_7240);
nand U10266 (N_10266,N_9171,N_6978);
and U10267 (N_10267,N_7258,N_8840);
and U10268 (N_10268,N_6623,N_9120);
xnor U10269 (N_10269,N_8206,N_7080);
nor U10270 (N_10270,N_8676,N_7439);
nand U10271 (N_10271,N_8028,N_6516);
nor U10272 (N_10272,N_7218,N_8294);
xor U10273 (N_10273,N_8166,N_8735);
nand U10274 (N_10274,N_9108,N_8114);
and U10275 (N_10275,N_6728,N_9200);
or U10276 (N_10276,N_9004,N_7858);
or U10277 (N_10277,N_6879,N_6679);
xor U10278 (N_10278,N_8583,N_8077);
or U10279 (N_10279,N_7434,N_9027);
nand U10280 (N_10280,N_6464,N_9350);
nand U10281 (N_10281,N_8029,N_7702);
and U10282 (N_10282,N_6357,N_6816);
or U10283 (N_10283,N_7814,N_8089);
and U10284 (N_10284,N_7332,N_8021);
and U10285 (N_10285,N_8138,N_7267);
nand U10286 (N_10286,N_7074,N_7736);
nor U10287 (N_10287,N_8268,N_7256);
nor U10288 (N_10288,N_7806,N_8893);
or U10289 (N_10289,N_7073,N_8715);
and U10290 (N_10290,N_8036,N_8139);
or U10291 (N_10291,N_8919,N_6436);
xnor U10292 (N_10292,N_8441,N_6726);
or U10293 (N_10293,N_7132,N_8824);
nor U10294 (N_10294,N_8249,N_9348);
nor U10295 (N_10295,N_7748,N_6458);
and U10296 (N_10296,N_6687,N_8566);
or U10297 (N_10297,N_6252,N_7284);
and U10298 (N_10298,N_7696,N_6368);
nand U10299 (N_10299,N_6714,N_6288);
and U10300 (N_10300,N_8392,N_7011);
xnor U10301 (N_10301,N_6875,N_7001);
nor U10302 (N_10302,N_8539,N_6945);
nand U10303 (N_10303,N_7839,N_8554);
nor U10304 (N_10304,N_7987,N_9347);
or U10305 (N_10305,N_7480,N_6715);
nand U10306 (N_10306,N_7356,N_8980);
or U10307 (N_10307,N_8886,N_8964);
nand U10308 (N_10308,N_8163,N_6339);
or U10309 (N_10309,N_8176,N_9142);
or U10310 (N_10310,N_9086,N_8727);
xnor U10311 (N_10311,N_7282,N_6893);
nor U10312 (N_10312,N_7135,N_7070);
xor U10313 (N_10313,N_9097,N_8065);
nor U10314 (N_10314,N_6389,N_6734);
xor U10315 (N_10315,N_7193,N_7934);
xor U10316 (N_10316,N_6617,N_6968);
or U10317 (N_10317,N_7449,N_7493);
xor U10318 (N_10318,N_7047,N_7438);
and U10319 (N_10319,N_7901,N_9007);
or U10320 (N_10320,N_8491,N_6833);
and U10321 (N_10321,N_8766,N_6982);
and U10322 (N_10322,N_6408,N_6738);
nand U10323 (N_10323,N_7003,N_7483);
xor U10324 (N_10324,N_7294,N_7618);
and U10325 (N_10325,N_8451,N_8587);
or U10326 (N_10326,N_6627,N_8277);
nand U10327 (N_10327,N_8200,N_8702);
nor U10328 (N_10328,N_7306,N_6585);
and U10329 (N_10329,N_6838,N_7995);
nand U10330 (N_10330,N_7948,N_6902);
nor U10331 (N_10331,N_8552,N_8931);
or U10332 (N_10332,N_9124,N_7297);
nor U10333 (N_10333,N_8073,N_8925);
nand U10334 (N_10334,N_6626,N_7740);
xnor U10335 (N_10335,N_6343,N_8010);
and U10336 (N_10336,N_9230,N_9025);
or U10337 (N_10337,N_8648,N_7171);
and U10338 (N_10338,N_8690,N_8368);
nor U10339 (N_10339,N_6702,N_7414);
nand U10340 (N_10340,N_6545,N_6862);
and U10341 (N_10341,N_7707,N_8197);
and U10342 (N_10342,N_7423,N_7636);
xor U10343 (N_10343,N_8870,N_8059);
xor U10344 (N_10344,N_7850,N_7362);
nand U10345 (N_10345,N_8783,N_8924);
nand U10346 (N_10346,N_7885,N_8860);
and U10347 (N_10347,N_8398,N_8760);
nand U10348 (N_10348,N_6504,N_6848);
xor U10349 (N_10349,N_7513,N_6641);
and U10350 (N_10350,N_7554,N_9074);
and U10351 (N_10351,N_7628,N_9277);
nor U10352 (N_10352,N_9296,N_8854);
or U10353 (N_10353,N_6460,N_9188);
or U10354 (N_10354,N_8659,N_8058);
nand U10355 (N_10355,N_8443,N_6445);
xor U10356 (N_10356,N_7009,N_7568);
nor U10357 (N_10357,N_8169,N_7712);
xnor U10358 (N_10358,N_8696,N_7325);
nor U10359 (N_10359,N_9330,N_7943);
nand U10360 (N_10360,N_6512,N_7429);
or U10361 (N_10361,N_8072,N_7730);
xnor U10362 (N_10362,N_8458,N_9009);
xor U10363 (N_10363,N_7516,N_8896);
and U10364 (N_10364,N_7642,N_7327);
nand U10365 (N_10365,N_7123,N_6707);
or U10366 (N_10366,N_6539,N_7027);
nor U10367 (N_10367,N_7752,N_7353);
and U10368 (N_10368,N_8578,N_9180);
nand U10369 (N_10369,N_7120,N_6847);
xor U10370 (N_10370,N_8047,N_6868);
or U10371 (N_10371,N_6770,N_7295);
and U10372 (N_10372,N_7262,N_6665);
and U10373 (N_10373,N_8492,N_7611);
or U10374 (N_10374,N_6396,N_8394);
and U10375 (N_10375,N_7113,N_8695);
nand U10376 (N_10376,N_8295,N_7204);
or U10377 (N_10377,N_7515,N_6961);
nand U10378 (N_10378,N_7355,N_8765);
nand U10379 (N_10379,N_7098,N_8926);
xnor U10380 (N_10380,N_7126,N_8768);
xnor U10381 (N_10381,N_6391,N_7946);
and U10382 (N_10382,N_9072,N_6822);
nor U10383 (N_10383,N_9238,N_8052);
xnor U10384 (N_10384,N_6663,N_7413);
xor U10385 (N_10385,N_7961,N_6814);
nand U10386 (N_10386,N_6991,N_6994);
xor U10387 (N_10387,N_7156,N_6360);
and U10388 (N_10388,N_6316,N_7710);
and U10389 (N_10389,N_8595,N_7695);
nor U10390 (N_10390,N_7478,N_6836);
xor U10391 (N_10391,N_6618,N_8287);
or U10392 (N_10392,N_9286,N_8172);
nand U10393 (N_10393,N_6295,N_7537);
nor U10394 (N_10394,N_8661,N_7594);
and U10395 (N_10395,N_7467,N_6976);
xnor U10396 (N_10396,N_7805,N_8814);
nor U10397 (N_10397,N_8542,N_7128);
nor U10398 (N_10398,N_8763,N_9061);
and U10399 (N_10399,N_7499,N_8198);
xnor U10400 (N_10400,N_7722,N_8406);
or U10401 (N_10401,N_8921,N_8274);
and U10402 (N_10402,N_8730,N_6488);
and U10403 (N_10403,N_7520,N_8961);
or U10404 (N_10404,N_7326,N_8940);
or U10405 (N_10405,N_7389,N_8551);
xor U10406 (N_10406,N_8260,N_8572);
xnor U10407 (N_10407,N_7683,N_8348);
nand U10408 (N_10408,N_9279,N_6721);
or U10409 (N_10409,N_6918,N_7102);
xnor U10410 (N_10410,N_9269,N_8519);
nand U10411 (N_10411,N_6639,N_7988);
or U10412 (N_10412,N_7260,N_7166);
and U10413 (N_10413,N_8215,N_7625);
nand U10414 (N_10414,N_6521,N_9092);
and U10415 (N_10415,N_8977,N_6588);
or U10416 (N_10416,N_9199,N_9168);
nor U10417 (N_10417,N_8815,N_9242);
nand U10418 (N_10418,N_8372,N_9166);
xor U10419 (N_10419,N_8827,N_8383);
nor U10420 (N_10420,N_8979,N_7876);
xor U10421 (N_10421,N_7095,N_7377);
or U10422 (N_10422,N_9371,N_7782);
or U10423 (N_10423,N_7700,N_7949);
and U10424 (N_10424,N_8270,N_7066);
and U10425 (N_10425,N_6965,N_9236);
or U10426 (N_10426,N_6607,N_7795);
nor U10427 (N_10427,N_9302,N_8511);
xor U10428 (N_10428,N_6606,N_6906);
nand U10429 (N_10429,N_8027,N_8341);
and U10430 (N_10430,N_6484,N_7308);
nor U10431 (N_10431,N_6414,N_7024);
and U10432 (N_10432,N_7774,N_7041);
xor U10433 (N_10433,N_8775,N_6533);
and U10434 (N_10434,N_8660,N_6870);
or U10435 (N_10435,N_6856,N_6582);
or U10436 (N_10436,N_8624,N_6799);
and U10437 (N_10437,N_7985,N_6579);
nand U10438 (N_10438,N_8119,N_7146);
or U10439 (N_10439,N_8293,N_7067);
or U10440 (N_10440,N_8239,N_8328);
nand U10441 (N_10441,N_8258,N_8999);
or U10442 (N_10442,N_7900,N_8291);
and U10443 (N_10443,N_6772,N_8905);
xor U10444 (N_10444,N_7720,N_6955);
nor U10445 (N_10445,N_6872,N_9260);
and U10446 (N_10446,N_7408,N_6583);
xor U10447 (N_10447,N_7535,N_7848);
nand U10448 (N_10448,N_9032,N_7310);
nor U10449 (N_10449,N_9174,N_6499);
or U10450 (N_10450,N_9312,N_8366);
or U10451 (N_10451,N_6537,N_8593);
xor U10452 (N_10452,N_7029,N_8598);
and U10453 (N_10453,N_8797,N_7374);
nand U10454 (N_10454,N_8042,N_8179);
nor U10455 (N_10455,N_6468,N_8968);
nor U10456 (N_10456,N_6594,N_7542);
xnor U10457 (N_10457,N_9345,N_7125);
nand U10458 (N_10458,N_7993,N_8688);
nor U10459 (N_10459,N_9038,N_6401);
and U10460 (N_10460,N_8680,N_6972);
and U10461 (N_10461,N_6699,N_9050);
nor U10462 (N_10462,N_6509,N_8904);
nor U10463 (N_10463,N_7974,N_8157);
nand U10464 (N_10464,N_7094,N_8088);
and U10465 (N_10465,N_8510,N_8030);
xnor U10466 (N_10466,N_6736,N_7176);
nand U10467 (N_10467,N_7252,N_8612);
nor U10468 (N_10468,N_6592,N_6471);
xnor U10469 (N_10469,N_6826,N_9226);
xor U10470 (N_10470,N_7514,N_6421);
or U10471 (N_10471,N_7954,N_8813);
nor U10472 (N_10472,N_8978,N_9164);
nor U10473 (N_10473,N_9222,N_8203);
nand U10474 (N_10474,N_8075,N_7231);
xnor U10475 (N_10475,N_8186,N_6334);
xor U10476 (N_10476,N_8110,N_6919);
xnor U10477 (N_10477,N_8151,N_9243);
nand U10478 (N_10478,N_8330,N_7141);
nand U10479 (N_10479,N_6794,N_8159);
and U10480 (N_10480,N_6432,N_8460);
xnor U10481 (N_10481,N_9102,N_8304);
or U10482 (N_10482,N_6546,N_6254);
or U10483 (N_10483,N_6302,N_6829);
and U10484 (N_10484,N_6575,N_6834);
and U10485 (N_10485,N_9229,N_8332);
and U10486 (N_10486,N_8532,N_7373);
nand U10487 (N_10487,N_8884,N_8165);
xor U10488 (N_10488,N_6466,N_7790);
xnor U10489 (N_10489,N_6412,N_6988);
and U10490 (N_10490,N_8100,N_6977);
nand U10491 (N_10491,N_6392,N_9070);
nor U10492 (N_10492,N_8984,N_8717);
or U10493 (N_10493,N_7052,N_8842);
xor U10494 (N_10494,N_9049,N_8078);
or U10495 (N_10495,N_6671,N_6362);
or U10496 (N_10496,N_6722,N_8470);
and U10497 (N_10497,N_8948,N_8264);
xnor U10498 (N_10498,N_7314,N_7751);
xor U10499 (N_10499,N_6620,N_8704);
and U10500 (N_10500,N_7742,N_6828);
xnor U10501 (N_10501,N_8026,N_6492);
or U10502 (N_10502,N_7650,N_8654);
and U10503 (N_10503,N_7249,N_6561);
or U10504 (N_10504,N_7038,N_9206);
or U10505 (N_10505,N_6793,N_7239);
xnor U10506 (N_10506,N_7504,N_8791);
and U10507 (N_10507,N_7488,N_8407);
nor U10508 (N_10508,N_8610,N_8278);
or U10509 (N_10509,N_7586,N_7832);
xnor U10510 (N_10510,N_9029,N_8538);
nor U10511 (N_10511,N_8778,N_6696);
xor U10512 (N_10512,N_8889,N_6407);
nand U10513 (N_10513,N_8555,N_6415);
xor U10514 (N_10514,N_7140,N_6284);
xor U10515 (N_10515,N_7036,N_8056);
xnor U10516 (N_10516,N_7533,N_9321);
nor U10517 (N_10517,N_7802,N_8350);
nand U10518 (N_10518,N_8857,N_7889);
nor U10519 (N_10519,N_7015,N_7924);
nor U10520 (N_10520,N_7021,N_8649);
nand U10521 (N_10521,N_7523,N_7956);
or U10522 (N_10522,N_8618,N_6435);
nor U10523 (N_10523,N_9241,N_9301);
nor U10524 (N_10524,N_9273,N_8636);
nor U10525 (N_10525,N_6312,N_6330);
and U10526 (N_10526,N_7780,N_6895);
nand U10527 (N_10527,N_8726,N_8581);
nand U10528 (N_10528,N_9186,N_7452);
and U10529 (N_10529,N_9087,N_7450);
nand U10530 (N_10530,N_8951,N_6577);
nand U10531 (N_10531,N_7643,N_9212);
nor U10532 (N_10532,N_8024,N_8531);
xor U10533 (N_10533,N_9147,N_6555);
xnor U10534 (N_10534,N_8254,N_6939);
xnor U10535 (N_10535,N_7764,N_7968);
and U10536 (N_10536,N_8991,N_8359);
and U10537 (N_10537,N_6442,N_6356);
or U10538 (N_10538,N_7129,N_8004);
or U10539 (N_10539,N_7226,N_7597);
and U10540 (N_10540,N_6692,N_7341);
and U10541 (N_10541,N_6646,N_8060);
nor U10542 (N_10542,N_6737,N_7606);
xor U10543 (N_10543,N_8897,N_6821);
nor U10544 (N_10544,N_7385,N_8136);
and U10545 (N_10545,N_7703,N_8432);
nand U10546 (N_10546,N_9158,N_9017);
and U10547 (N_10547,N_7540,N_8496);
nand U10548 (N_10548,N_6346,N_6832);
nand U10549 (N_10549,N_6783,N_7602);
or U10550 (N_10550,N_7321,N_9141);
xor U10551 (N_10551,N_7875,N_6869);
and U10552 (N_10552,N_6859,N_9000);
and U10553 (N_10553,N_8733,N_6267);
xor U10554 (N_10554,N_8737,N_8751);
and U10555 (N_10555,N_8439,N_8719);
nor U10556 (N_10556,N_7675,N_7892);
or U10557 (N_10557,N_6970,N_8756);
or U10558 (N_10558,N_8939,N_6842);
and U10559 (N_10559,N_6792,N_7118);
and U10560 (N_10560,N_7302,N_9133);
nor U10561 (N_10561,N_7232,N_7417);
xor U10562 (N_10562,N_7786,N_9203);
and U10563 (N_10563,N_8482,N_8381);
nor U10564 (N_10564,N_6866,N_9054);
or U10565 (N_10565,N_6544,N_8549);
nand U10566 (N_10566,N_8085,N_7476);
xnor U10567 (N_10567,N_6891,N_8153);
nor U10568 (N_10568,N_8435,N_6796);
and U10569 (N_10569,N_8705,N_8946);
and U10570 (N_10570,N_8424,N_7971);
or U10571 (N_10571,N_8221,N_7601);
and U10572 (N_10572,N_8706,N_7330);
and U10573 (N_10573,N_6678,N_6487);
nand U10574 (N_10574,N_7386,N_9146);
xnor U10575 (N_10575,N_7928,N_6344);
and U10576 (N_10576,N_7484,N_7958);
nand U10577 (N_10577,N_6454,N_7085);
nor U10578 (N_10578,N_8263,N_8377);
xor U10579 (N_10579,N_7044,N_8011);
nor U10580 (N_10580,N_8486,N_8128);
or U10581 (N_10581,N_7827,N_6786);
nand U10582 (N_10582,N_6677,N_8996);
and U10583 (N_10583,N_8888,N_6404);
and U10584 (N_10584,N_7290,N_6803);
nand U10585 (N_10585,N_7035,N_8102);
or U10586 (N_10586,N_9042,N_8420);
xor U10587 (N_10587,N_8652,N_7020);
and U10588 (N_10588,N_8132,N_7090);
xor U10589 (N_10589,N_7996,N_8985);
xor U10590 (N_10590,N_8459,N_8743);
nand U10591 (N_10591,N_9064,N_8425);
and U10592 (N_10592,N_6664,N_8534);
nand U10593 (N_10593,N_9127,N_9194);
xor U10594 (N_10594,N_9289,N_8450);
xor U10595 (N_10595,N_8302,N_7139);
or U10596 (N_10596,N_8314,N_8820);
nor U10597 (N_10597,N_9266,N_9095);
xor U10598 (N_10598,N_7440,N_8633);
and U10599 (N_10599,N_8067,N_7530);
xor U10600 (N_10600,N_8064,N_6268);
xor U10601 (N_10601,N_7903,N_8782);
nand U10602 (N_10602,N_7578,N_6778);
or U10603 (N_10603,N_7069,N_6473);
nand U10604 (N_10604,N_9278,N_8645);
xnor U10605 (N_10605,N_8634,N_7019);
nor U10606 (N_10606,N_9165,N_9128);
xnor U10607 (N_10607,N_6270,N_7275);
nand U10608 (N_10608,N_8709,N_8236);
and U10609 (N_10609,N_8627,N_8149);
nand U10610 (N_10610,N_8411,N_8806);
or U10611 (N_10611,N_6600,N_9065);
xnor U10612 (N_10612,N_7329,N_8080);
nor U10613 (N_10613,N_7430,N_7448);
nand U10614 (N_10614,N_6359,N_7972);
nand U10615 (N_10615,N_6637,N_7432);
or U10616 (N_10616,N_9331,N_7992);
and U10617 (N_10617,N_7698,N_8525);
and U10618 (N_10618,N_9290,N_8417);
nand U10619 (N_10619,N_9340,N_7561);
nor U10620 (N_10620,N_8635,N_8955);
xnor U10621 (N_10621,N_7849,N_7603);
nand U10622 (N_10622,N_7725,N_8044);
and U10623 (N_10623,N_8113,N_8063);
or U10624 (N_10624,N_8107,N_8423);
nor U10625 (N_10625,N_6873,N_9067);
and U10626 (N_10626,N_7633,N_7868);
nand U10627 (N_10627,N_7115,N_7789);
and U10628 (N_10628,N_8031,N_8217);
or U10629 (N_10629,N_7382,N_8916);
or U10630 (N_10630,N_8747,N_8438);
nand U10631 (N_10631,N_9071,N_7835);
nand U10632 (N_10632,N_6662,N_7917);
xor U10633 (N_10633,N_8329,N_6559);
or U10634 (N_10634,N_7808,N_8569);
xor U10635 (N_10635,N_6650,N_8105);
or U10636 (N_10636,N_9157,N_7590);
nor U10637 (N_10637,N_7746,N_6290);
and U10638 (N_10638,N_9094,N_9309);
xnor U10639 (N_10639,N_8617,N_6491);
nand U10640 (N_10640,N_7638,N_7870);
or U10641 (N_10641,N_8300,N_8903);
and U10642 (N_10642,N_8682,N_7756);
or U10643 (N_10643,N_8325,N_7433);
and U10644 (N_10644,N_6355,N_9197);
nand U10645 (N_10645,N_7942,N_9169);
nand U10646 (N_10646,N_6605,N_6300);
nor U10647 (N_10647,N_8687,N_9276);
and U10648 (N_10648,N_7079,N_6422);
nand U10649 (N_10649,N_7979,N_7259);
nand U10650 (N_10650,N_9239,N_6840);
xnor U10651 (N_10651,N_7883,N_8137);
or U10652 (N_10652,N_7788,N_8009);
xor U10653 (N_10653,N_6776,N_8992);
nand U10654 (N_10654,N_7242,N_7635);
and U10655 (N_10655,N_7489,N_6901);
or U10656 (N_10656,N_9117,N_7202);
nor U10657 (N_10657,N_8553,N_6629);
or U10658 (N_10658,N_6632,N_6437);
nand U10659 (N_10659,N_8337,N_9058);
nor U10660 (N_10660,N_7672,N_6418);
or U10661 (N_10661,N_6749,N_9139);
nor U10662 (N_10662,N_7963,N_9045);
xnor U10663 (N_10663,N_6740,N_7412);
or U10664 (N_10664,N_6328,N_6431);
and U10665 (N_10665,N_7502,N_8601);
nor U10666 (N_10666,N_9332,N_9361);
and U10667 (N_10667,N_7101,N_7716);
or U10668 (N_10668,N_7292,N_8609);
or U10669 (N_10669,N_9274,N_7646);
and U10670 (N_10670,N_7455,N_8414);
or U10671 (N_10671,N_8899,N_8355);
nand U10672 (N_10672,N_8430,N_8872);
nand U10673 (N_10673,N_7311,N_7955);
nand U10674 (N_10674,N_9288,N_7064);
nor U10675 (N_10675,N_8667,N_8642);
and U10676 (N_10676,N_8738,N_6892);
nand U10677 (N_10677,N_8693,N_8679);
xnor U10678 (N_10678,N_8193,N_6410);
nand U10679 (N_10679,N_7116,N_8347);
xnor U10680 (N_10680,N_7390,N_7215);
nand U10681 (N_10681,N_6364,N_8070);
nand U10682 (N_10682,N_8484,N_7145);
or U10683 (N_10683,N_6751,N_6500);
or U10684 (N_10684,N_9281,N_8211);
xnor U10685 (N_10685,N_7061,N_7178);
nor U10686 (N_10686,N_8678,N_7309);
xnor U10687 (N_10687,N_9079,N_6292);
nand U10688 (N_10688,N_6361,N_7361);
xor U10689 (N_10689,N_8712,N_8983);
and U10690 (N_10690,N_9355,N_8205);
nor U10691 (N_10691,N_7227,N_8914);
and U10692 (N_10692,N_8316,N_8335);
nand U10693 (N_10693,N_7711,N_8520);
nand U10694 (N_10694,N_7110,N_6686);
xnor U10695 (N_10695,N_6923,N_8468);
or U10696 (N_10696,N_6327,N_6542);
nor U10697 (N_10697,N_8440,N_6676);
and U10698 (N_10698,N_8228,N_7727);
nor U10699 (N_10699,N_7687,N_6462);
xnor U10700 (N_10700,N_8086,N_7347);
nor U10701 (N_10701,N_6508,N_6340);
and U10702 (N_10702,N_9005,N_8773);
or U10703 (N_10703,N_6527,N_8850);
or U10704 (N_10704,N_9195,N_7447);
and U10705 (N_10705,N_8299,N_8993);
and U10706 (N_10706,N_7991,N_8505);
xor U10707 (N_10707,N_7909,N_8918);
nand U10708 (N_10708,N_7709,N_6990);
nand U10709 (N_10709,N_9234,N_8600);
or U10710 (N_10710,N_7165,N_9326);
and U10711 (N_10711,N_6430,N_7656);
or U10712 (N_10712,N_8049,N_6447);
nand U10713 (N_10713,N_7247,N_6724);
nor U10714 (N_10714,N_9130,N_7645);
nand U10715 (N_10715,N_8997,N_7285);
or U10716 (N_10716,N_8288,N_6827);
or U10717 (N_10717,N_9252,N_7147);
and U10718 (N_10718,N_7043,N_8495);
and U10719 (N_10719,N_8758,N_8607);
nand U10720 (N_10720,N_6966,N_7196);
and U10721 (N_10721,N_6880,N_6310);
nor U10722 (N_10722,N_8413,N_6399);
xnor U10723 (N_10723,N_7427,N_7546);
or U10724 (N_10724,N_8369,N_7372);
xnor U10725 (N_10725,N_8994,N_8845);
nor U10726 (N_10726,N_8720,N_6951);
and U10727 (N_10727,N_6974,N_7071);
and U10728 (N_10728,N_8340,N_6638);
and U10729 (N_10729,N_7474,N_9154);
nor U10730 (N_10730,N_8386,N_8389);
xor U10731 (N_10731,N_9349,N_7365);
and U10732 (N_10732,N_6815,N_8740);
or U10733 (N_10733,N_9196,N_6556);
and U10734 (N_10734,N_9040,N_8686);
or U10735 (N_10735,N_7152,N_8644);
or U10736 (N_10736,N_6739,N_8913);
nand U10737 (N_10737,N_7668,N_9298);
nand U10738 (N_10738,N_6475,N_8195);
xor U10739 (N_10739,N_6285,N_8849);
nand U10740 (N_10740,N_7960,N_9110);
and U10741 (N_10741,N_8568,N_7670);
nor U10742 (N_10742,N_7144,N_8244);
nor U10743 (N_10743,N_6352,N_8529);
nor U10744 (N_10744,N_9339,N_7322);
nand U10745 (N_10745,N_6779,N_8498);
xor U10746 (N_10746,N_7831,N_8184);
nor U10747 (N_10747,N_7164,N_8250);
nand U10748 (N_10748,N_7897,N_8445);
xor U10749 (N_10749,N_7701,N_6914);
xor U10750 (N_10750,N_6689,N_8252);
nor U10751 (N_10751,N_9268,N_7137);
nand U10752 (N_10752,N_7470,N_7319);
or U10753 (N_10753,N_7846,N_7122);
and U10754 (N_10754,N_7158,N_6273);
or U10755 (N_10755,N_7843,N_6351);
xor U10756 (N_10756,N_7694,N_8881);
nor U10757 (N_10757,N_7800,N_7614);
and U10758 (N_10758,N_7761,N_7598);
and U10759 (N_10759,N_6809,N_7160);
nor U10760 (N_10760,N_7673,N_6382);
nand U10761 (N_10761,N_9135,N_6935);
xor U10762 (N_10762,N_7872,N_7735);
and U10763 (N_10763,N_6423,N_8351);
or U10764 (N_10764,N_7544,N_7401);
xnor U10765 (N_10765,N_7177,N_8796);
nand U10766 (N_10766,N_8967,N_8655);
and U10767 (N_10767,N_7464,N_6574);
or U10768 (N_10768,N_9008,N_8266);
xor U10769 (N_10769,N_6730,N_7398);
xor U10770 (N_10770,N_7624,N_7013);
nand U10771 (N_10771,N_6541,N_8623);
and U10772 (N_10772,N_7784,N_6851);
xnor U10773 (N_10773,N_7608,N_6524);
and U10774 (N_10774,N_8129,N_7065);
or U10775 (N_10775,N_8188,N_6673);
nand U10776 (N_10776,N_9003,N_7932);
nor U10777 (N_10777,N_8141,N_8577);
nand U10778 (N_10778,N_7487,N_6478);
nand U10779 (N_10779,N_6580,N_6480);
xor U10780 (N_10780,N_9346,N_7529);
xnor U10781 (N_10781,N_7908,N_7345);
nand U10782 (N_10782,N_6909,N_9113);
or U10783 (N_10783,N_8361,N_7864);
nor U10784 (N_10784,N_6963,N_9170);
nand U10785 (N_10785,N_7654,N_7631);
or U10786 (N_10786,N_8493,N_6271);
xor U10787 (N_10787,N_8615,N_7136);
nor U10788 (N_10788,N_6782,N_7379);
xnor U10789 (N_10789,N_9291,N_7519);
xnor U10790 (N_10790,N_8204,N_7822);
and U10791 (N_10791,N_8509,N_8811);
xnor U10792 (N_10792,N_7351,N_8923);
and U10793 (N_10793,N_9091,N_9159);
and U10794 (N_10794,N_7762,N_7461);
nand U10795 (N_10795,N_9015,N_8592);
xor U10796 (N_10796,N_6804,N_7538);
nor U10797 (N_10797,N_8220,N_7112);
xnor U10798 (N_10798,N_8546,N_7824);
xnor U10799 (N_10799,N_9143,N_8345);
nor U10800 (N_10800,N_7686,N_6526);
or U10801 (N_10801,N_7905,N_7769);
xnor U10802 (N_10802,N_8360,N_7528);
nor U10803 (N_10803,N_6670,N_7273);
and U10804 (N_10804,N_6333,N_7367);
or U10805 (N_10805,N_7997,N_8201);
nor U10806 (N_10806,N_9037,N_7787);
nand U10807 (N_10807,N_7428,N_8306);
and U10808 (N_10808,N_8564,N_6419);
nor U10809 (N_10809,N_8327,N_7181);
or U10810 (N_10810,N_7511,N_8449);
xnor U10811 (N_10811,N_7369,N_8083);
or U10812 (N_10812,N_6489,N_6801);
xnor U10813 (N_10813,N_7091,N_7443);
xor U10814 (N_10814,N_6745,N_7481);
and U10815 (N_10815,N_6675,N_6839);
nand U10816 (N_10816,N_7056,N_6358);
nor U10817 (N_10817,N_8521,N_6320);
or U10818 (N_10818,N_7804,N_7738);
and U10819 (N_10819,N_6927,N_6496);
nand U10820 (N_10820,N_6947,N_6294);
or U10821 (N_10821,N_6551,N_6434);
or U10822 (N_10822,N_7803,N_8269);
or U10823 (N_10823,N_7816,N_8672);
or U10824 (N_10824,N_8016,N_7299);
or U10825 (N_10825,N_6531,N_8237);
or U10826 (N_10826,N_6557,N_8944);
nor U10827 (N_10827,N_7415,N_8506);
xnor U10828 (N_10828,N_8877,N_8809);
nand U10829 (N_10829,N_6967,N_7324);
and U10830 (N_10830,N_6748,N_7916);
nand U10831 (N_10831,N_9342,N_8844);
nand U10832 (N_10832,N_7715,N_9024);
and U10833 (N_10833,N_8134,N_8640);
nor U10834 (N_10834,N_8222,N_6315);
xnor U10835 (N_10835,N_7926,N_8164);
nor U10836 (N_10836,N_9225,N_7281);
nand U10837 (N_10837,N_8995,N_6954);
xnor U10838 (N_10838,N_8673,N_7893);
nor U10839 (N_10839,N_8911,N_7477);
nand U10840 (N_10840,N_6905,N_7745);
or U10841 (N_10841,N_7508,N_7238);
and U10842 (N_10842,N_8518,N_8415);
xnor U10843 (N_10843,N_9341,N_8421);
nor U10844 (N_10844,N_8403,N_8808);
nor U10845 (N_10845,N_7222,N_7296);
nand U10846 (N_10846,N_9254,N_7241);
nor U10847 (N_10847,N_6338,N_6997);
and U10848 (N_10848,N_8099,N_8869);
and U10849 (N_10849,N_8677,N_6573);
and U10850 (N_10850,N_6377,N_7300);
xor U10851 (N_10851,N_8537,N_7050);
xor U10852 (N_10852,N_7794,N_7865);
nor U10853 (N_10853,N_8405,N_7944);
nor U10854 (N_10854,N_6269,N_6691);
nor U10855 (N_10855,N_7391,N_6709);
nand U10856 (N_10856,N_8507,N_9271);
or U10857 (N_10857,N_6998,N_9063);
nor U10858 (N_10858,N_7037,N_7759);
nand U10859 (N_10859,N_8251,N_9343);
xor U10860 (N_10860,N_8140,N_6690);
and U10861 (N_10861,N_6957,N_8479);
and U10862 (N_10862,N_7792,N_8523);
and U10863 (N_10863,N_8721,N_9315);
xnor U10864 (N_10864,N_7100,N_8668);
or U10865 (N_10865,N_8281,N_7465);
nor U10866 (N_10866,N_6465,N_7199);
nand U10867 (N_10867,N_6501,N_8516);
nor U10868 (N_10868,N_6305,N_9136);
xnor U10869 (N_10869,N_8116,N_6309);
and U10870 (N_10870,N_8358,N_6411);
nand U10871 (N_10871,N_9216,N_6613);
xor U10872 (N_10872,N_6987,N_7692);
nor U10873 (N_10873,N_7409,N_9320);
or U10874 (N_10874,N_6506,N_7304);
or U10875 (N_10875,N_9232,N_6476);
xnor U10876 (N_10876,N_8707,N_8109);
nand U10877 (N_10877,N_8958,N_9167);
xor U10878 (N_10878,N_6708,N_6725);
and U10879 (N_10879,N_7655,N_8455);
nand U10880 (N_10880,N_7269,N_6495);
nor U10881 (N_10881,N_7760,N_8280);
and U10882 (N_10882,N_9118,N_6884);
or U10883 (N_10883,N_6986,N_7690);
nand U10884 (N_10884,N_6941,N_7097);
or U10885 (N_10885,N_8379,N_6881);
nand U10886 (N_10886,N_8227,N_7143);
nor U10887 (N_10887,N_7082,N_8966);
or U10888 (N_10888,N_6964,N_7040);
and U10889 (N_10889,N_8057,N_9111);
nor U10890 (N_10890,N_8446,N_6733);
nor U10891 (N_10891,N_9204,N_8465);
xnor U10892 (N_10892,N_8255,N_8019);
and U10893 (N_10893,N_8628,N_8825);
nor U10894 (N_10894,N_6913,N_8802);
nor U10895 (N_10895,N_7640,N_7830);
and U10896 (N_10896,N_7276,N_7813);
and U10897 (N_10897,N_6482,N_7522);
and U10898 (N_10898,N_6428,N_6992);
nor U10899 (N_10899,N_8882,N_6413);
and U10900 (N_10900,N_8103,N_8066);
and U10901 (N_10901,N_8247,N_9156);
nand U10902 (N_10902,N_6621,N_8837);
nor U10903 (N_10903,N_9098,N_7682);
xor U10904 (N_10904,N_7623,N_6775);
nor U10905 (N_10905,N_7026,N_7651);
and U10906 (N_10906,N_7340,N_8106);
or U10907 (N_10907,N_7213,N_6757);
or U10908 (N_10908,N_8448,N_7731);
xnor U10909 (N_10909,N_9140,N_8757);
or U10910 (N_10910,N_8125,N_7331);
and U10911 (N_10911,N_9163,N_6720);
nor U10912 (N_10912,N_6348,N_6450);
or U10913 (N_10913,N_7721,N_9105);
nand U10914 (N_10914,N_8885,N_7857);
or U10915 (N_10915,N_7142,N_8365);
nand U10916 (N_10916,N_8917,N_9262);
nor U10917 (N_10917,N_8774,N_8867);
nand U10918 (N_10918,N_9189,N_9364);
and U10919 (N_10919,N_8746,N_9210);
nor U10920 (N_10920,N_7424,N_9228);
nand U10921 (N_10921,N_6788,N_8322);
nor U10922 (N_10922,N_7659,N_8055);
nand U10923 (N_10923,N_7194,N_8596);
or U10924 (N_10924,N_8547,N_6514);
nand U10925 (N_10925,N_6563,N_9372);
nand U10926 (N_10926,N_7860,N_7665);
and U10927 (N_10927,N_8038,N_6570);
nand U10928 (N_10928,N_7945,N_8834);
nand U10929 (N_10929,N_8214,N_7250);
nor U10930 (N_10930,N_8096,N_8685);
nand U10931 (N_10931,N_6943,N_6912);
and U10932 (N_10932,N_6443,N_7986);
nand U10933 (N_10933,N_7776,N_6520);
xor U10934 (N_10934,N_8282,N_7880);
and U10935 (N_10935,N_7970,N_7878);
nand U10936 (N_10936,N_7851,N_7010);
and U10937 (N_10937,N_8127,N_8807);
nor U10938 (N_10938,N_8348,N_7559);
xnor U10939 (N_10939,N_8616,N_6894);
nor U10940 (N_10940,N_7775,N_8087);
nor U10941 (N_10941,N_9092,N_8016);
nand U10942 (N_10942,N_6937,N_7834);
or U10943 (N_10943,N_6864,N_9138);
nand U10944 (N_10944,N_8349,N_7725);
nor U10945 (N_10945,N_7763,N_7906);
nand U10946 (N_10946,N_8861,N_9003);
and U10947 (N_10947,N_9196,N_6808);
and U10948 (N_10948,N_8485,N_8737);
or U10949 (N_10949,N_6523,N_7825);
nor U10950 (N_10950,N_7400,N_7118);
and U10951 (N_10951,N_8332,N_8645);
xor U10952 (N_10952,N_9231,N_8197);
nor U10953 (N_10953,N_6929,N_6312);
nand U10954 (N_10954,N_8078,N_7939);
nand U10955 (N_10955,N_6342,N_9092);
nand U10956 (N_10956,N_7571,N_7930);
xor U10957 (N_10957,N_7196,N_7226);
or U10958 (N_10958,N_9166,N_6454);
nor U10959 (N_10959,N_6840,N_8997);
nor U10960 (N_10960,N_8497,N_6292);
nor U10961 (N_10961,N_8479,N_7590);
nand U10962 (N_10962,N_8475,N_8560);
nor U10963 (N_10963,N_7272,N_7779);
or U10964 (N_10964,N_6356,N_8627);
and U10965 (N_10965,N_8070,N_8046);
nand U10966 (N_10966,N_6536,N_9074);
xor U10967 (N_10967,N_7258,N_7832);
or U10968 (N_10968,N_7553,N_7388);
nand U10969 (N_10969,N_8071,N_8277);
nor U10970 (N_10970,N_6409,N_6708);
or U10971 (N_10971,N_6919,N_6576);
nand U10972 (N_10972,N_6719,N_6376);
nand U10973 (N_10973,N_7549,N_8821);
nand U10974 (N_10974,N_6862,N_7241);
and U10975 (N_10975,N_8418,N_7276);
or U10976 (N_10976,N_7330,N_8746);
and U10977 (N_10977,N_6968,N_7210);
or U10978 (N_10978,N_8016,N_7097);
or U10979 (N_10979,N_9037,N_9297);
or U10980 (N_10980,N_6280,N_7898);
and U10981 (N_10981,N_6649,N_7413);
nor U10982 (N_10982,N_9181,N_7330);
or U10983 (N_10983,N_7304,N_8584);
xor U10984 (N_10984,N_6552,N_6953);
xnor U10985 (N_10985,N_7308,N_6357);
or U10986 (N_10986,N_6555,N_7282);
nor U10987 (N_10987,N_9199,N_9242);
nand U10988 (N_10988,N_6827,N_8321);
xor U10989 (N_10989,N_6942,N_7213);
nand U10990 (N_10990,N_8899,N_9122);
xnor U10991 (N_10991,N_7197,N_7896);
and U10992 (N_10992,N_7527,N_6622);
or U10993 (N_10993,N_7801,N_8702);
or U10994 (N_10994,N_8966,N_6502);
nor U10995 (N_10995,N_8899,N_7449);
xnor U10996 (N_10996,N_6838,N_8647);
nand U10997 (N_10997,N_6401,N_6391);
xor U10998 (N_10998,N_8656,N_6905);
and U10999 (N_10999,N_9292,N_8459);
and U11000 (N_11000,N_7932,N_8768);
xnor U11001 (N_11001,N_8875,N_7706);
nand U11002 (N_11002,N_9171,N_9042);
nor U11003 (N_11003,N_6298,N_6534);
and U11004 (N_11004,N_7477,N_8603);
or U11005 (N_11005,N_7900,N_7017);
xor U11006 (N_11006,N_9044,N_8567);
and U11007 (N_11007,N_8204,N_7613);
and U11008 (N_11008,N_9035,N_6722);
and U11009 (N_11009,N_6806,N_7656);
nor U11010 (N_11010,N_7846,N_9005);
and U11011 (N_11011,N_6679,N_9295);
xor U11012 (N_11012,N_6970,N_6808);
nand U11013 (N_11013,N_8785,N_6473);
or U11014 (N_11014,N_7123,N_9095);
or U11015 (N_11015,N_8854,N_7758);
nand U11016 (N_11016,N_6788,N_6386);
xor U11017 (N_11017,N_6596,N_6861);
or U11018 (N_11018,N_7476,N_8397);
nor U11019 (N_11019,N_7915,N_7262);
or U11020 (N_11020,N_8046,N_7081);
nor U11021 (N_11021,N_8517,N_8658);
and U11022 (N_11022,N_6462,N_6886);
nor U11023 (N_11023,N_7465,N_7844);
and U11024 (N_11024,N_7469,N_7380);
nand U11025 (N_11025,N_7112,N_6491);
and U11026 (N_11026,N_9262,N_7531);
or U11027 (N_11027,N_6783,N_7257);
nand U11028 (N_11028,N_7855,N_8252);
nand U11029 (N_11029,N_9181,N_8116);
xor U11030 (N_11030,N_6897,N_8491);
xor U11031 (N_11031,N_7323,N_7813);
and U11032 (N_11032,N_7027,N_9290);
xnor U11033 (N_11033,N_8780,N_7827);
xor U11034 (N_11034,N_8072,N_8092);
xnor U11035 (N_11035,N_6900,N_8580);
nand U11036 (N_11036,N_8011,N_7344);
nand U11037 (N_11037,N_8877,N_9054);
or U11038 (N_11038,N_7961,N_6767);
nand U11039 (N_11039,N_8839,N_6907);
or U11040 (N_11040,N_6949,N_6458);
nand U11041 (N_11041,N_7922,N_6727);
xor U11042 (N_11042,N_8656,N_8117);
nor U11043 (N_11043,N_8986,N_6484);
nand U11044 (N_11044,N_8128,N_6541);
nand U11045 (N_11045,N_8549,N_9028);
nand U11046 (N_11046,N_6713,N_6526);
and U11047 (N_11047,N_6738,N_8321);
or U11048 (N_11048,N_6878,N_8123);
nand U11049 (N_11049,N_6528,N_7525);
and U11050 (N_11050,N_6270,N_7930);
nor U11051 (N_11051,N_9007,N_8495);
nand U11052 (N_11052,N_7089,N_8697);
and U11053 (N_11053,N_8867,N_7777);
or U11054 (N_11054,N_9126,N_8664);
nand U11055 (N_11055,N_8344,N_7565);
nor U11056 (N_11056,N_6323,N_8588);
and U11057 (N_11057,N_7692,N_8672);
nor U11058 (N_11058,N_7929,N_6660);
nand U11059 (N_11059,N_8809,N_8299);
nor U11060 (N_11060,N_7550,N_8763);
xnor U11061 (N_11061,N_6353,N_9124);
nor U11062 (N_11062,N_8625,N_6965);
nand U11063 (N_11063,N_8634,N_6757);
xnor U11064 (N_11064,N_8227,N_6251);
and U11065 (N_11065,N_6924,N_8445);
nor U11066 (N_11066,N_7628,N_9358);
xnor U11067 (N_11067,N_6296,N_6431);
xor U11068 (N_11068,N_8326,N_7030);
and U11069 (N_11069,N_6707,N_8804);
nand U11070 (N_11070,N_8443,N_7307);
or U11071 (N_11071,N_8129,N_8018);
xnor U11072 (N_11072,N_8156,N_9097);
or U11073 (N_11073,N_9177,N_8011);
xor U11074 (N_11074,N_6683,N_8305);
nor U11075 (N_11075,N_8174,N_8213);
and U11076 (N_11076,N_8282,N_7110);
or U11077 (N_11077,N_6538,N_6437);
nand U11078 (N_11078,N_9270,N_7212);
xor U11079 (N_11079,N_8784,N_8900);
and U11080 (N_11080,N_6944,N_7689);
or U11081 (N_11081,N_9114,N_7997);
or U11082 (N_11082,N_8687,N_9287);
or U11083 (N_11083,N_7806,N_6712);
nor U11084 (N_11084,N_6308,N_7191);
and U11085 (N_11085,N_8766,N_6715);
nand U11086 (N_11086,N_8683,N_8968);
nor U11087 (N_11087,N_7560,N_9047);
or U11088 (N_11088,N_8092,N_8464);
nor U11089 (N_11089,N_6318,N_6634);
nor U11090 (N_11090,N_6819,N_6979);
and U11091 (N_11091,N_6315,N_7479);
or U11092 (N_11092,N_7828,N_9021);
or U11093 (N_11093,N_7116,N_6620);
and U11094 (N_11094,N_8632,N_7099);
nand U11095 (N_11095,N_8363,N_6724);
nand U11096 (N_11096,N_6331,N_8417);
xor U11097 (N_11097,N_7109,N_7974);
and U11098 (N_11098,N_8973,N_8328);
or U11099 (N_11099,N_7614,N_8833);
and U11100 (N_11100,N_7333,N_6913);
nand U11101 (N_11101,N_6909,N_8513);
xor U11102 (N_11102,N_8393,N_6308);
xnor U11103 (N_11103,N_7487,N_7944);
xor U11104 (N_11104,N_8028,N_7208);
nor U11105 (N_11105,N_7672,N_7524);
and U11106 (N_11106,N_8590,N_6313);
nand U11107 (N_11107,N_6429,N_7662);
nor U11108 (N_11108,N_6866,N_6280);
xnor U11109 (N_11109,N_6303,N_8568);
xnor U11110 (N_11110,N_8484,N_9143);
and U11111 (N_11111,N_8702,N_6265);
or U11112 (N_11112,N_6653,N_7853);
and U11113 (N_11113,N_6989,N_8266);
or U11114 (N_11114,N_7699,N_8611);
xor U11115 (N_11115,N_8852,N_9067);
and U11116 (N_11116,N_8741,N_9128);
nor U11117 (N_11117,N_7465,N_7892);
nand U11118 (N_11118,N_7986,N_8446);
xnor U11119 (N_11119,N_8298,N_8434);
xnor U11120 (N_11120,N_8106,N_7835);
or U11121 (N_11121,N_8370,N_6948);
xnor U11122 (N_11122,N_8922,N_8649);
and U11123 (N_11123,N_8081,N_7340);
nor U11124 (N_11124,N_7907,N_6570);
and U11125 (N_11125,N_7065,N_8601);
and U11126 (N_11126,N_9238,N_7636);
and U11127 (N_11127,N_8758,N_9348);
nand U11128 (N_11128,N_8872,N_6275);
or U11129 (N_11129,N_8668,N_7024);
or U11130 (N_11130,N_8443,N_7046);
or U11131 (N_11131,N_7596,N_8400);
nand U11132 (N_11132,N_7757,N_7566);
or U11133 (N_11133,N_6580,N_8384);
xor U11134 (N_11134,N_7822,N_7025);
nor U11135 (N_11135,N_8032,N_8919);
xnor U11136 (N_11136,N_8145,N_6784);
nand U11137 (N_11137,N_8877,N_8808);
nand U11138 (N_11138,N_6369,N_7968);
nand U11139 (N_11139,N_7780,N_7996);
nand U11140 (N_11140,N_8908,N_6839);
nand U11141 (N_11141,N_6657,N_8944);
xnor U11142 (N_11142,N_8818,N_8691);
nor U11143 (N_11143,N_7382,N_7026);
xnor U11144 (N_11144,N_8380,N_7259);
xnor U11145 (N_11145,N_6663,N_7730);
and U11146 (N_11146,N_8669,N_7958);
xor U11147 (N_11147,N_6419,N_6671);
or U11148 (N_11148,N_7533,N_6749);
xor U11149 (N_11149,N_8853,N_6601);
or U11150 (N_11150,N_8589,N_7246);
xnor U11151 (N_11151,N_6568,N_8703);
and U11152 (N_11152,N_8171,N_7644);
or U11153 (N_11153,N_9057,N_8726);
xor U11154 (N_11154,N_7768,N_6853);
nor U11155 (N_11155,N_8029,N_8500);
nand U11156 (N_11156,N_8777,N_8646);
xnor U11157 (N_11157,N_6271,N_9337);
and U11158 (N_11158,N_8039,N_7163);
nor U11159 (N_11159,N_6611,N_7544);
xnor U11160 (N_11160,N_7271,N_7528);
and U11161 (N_11161,N_6509,N_6680);
and U11162 (N_11162,N_6486,N_7232);
xor U11163 (N_11163,N_7746,N_7935);
nor U11164 (N_11164,N_7381,N_8991);
nand U11165 (N_11165,N_9287,N_7366);
xor U11166 (N_11166,N_6428,N_6357);
and U11167 (N_11167,N_6364,N_6291);
or U11168 (N_11168,N_7958,N_8284);
xnor U11169 (N_11169,N_7533,N_8101);
nand U11170 (N_11170,N_6870,N_7765);
and U11171 (N_11171,N_7356,N_9262);
or U11172 (N_11172,N_8501,N_8577);
xnor U11173 (N_11173,N_9143,N_8243);
nand U11174 (N_11174,N_8078,N_7124);
xnor U11175 (N_11175,N_7549,N_9251);
or U11176 (N_11176,N_7493,N_8299);
nand U11177 (N_11177,N_7639,N_6606);
or U11178 (N_11178,N_7554,N_8570);
nor U11179 (N_11179,N_7180,N_6461);
nand U11180 (N_11180,N_6821,N_9359);
xnor U11181 (N_11181,N_8852,N_8951);
xnor U11182 (N_11182,N_7100,N_6413);
or U11183 (N_11183,N_6957,N_7280);
nand U11184 (N_11184,N_6983,N_8602);
or U11185 (N_11185,N_8546,N_8359);
or U11186 (N_11186,N_8444,N_6704);
xnor U11187 (N_11187,N_6627,N_8738);
or U11188 (N_11188,N_7228,N_7376);
nand U11189 (N_11189,N_6718,N_6275);
and U11190 (N_11190,N_7819,N_8968);
and U11191 (N_11191,N_8036,N_8721);
nor U11192 (N_11192,N_8221,N_8986);
nand U11193 (N_11193,N_7876,N_9016);
nor U11194 (N_11194,N_7701,N_6858);
nand U11195 (N_11195,N_7409,N_6902);
xnor U11196 (N_11196,N_7252,N_7585);
or U11197 (N_11197,N_8361,N_8986);
nor U11198 (N_11198,N_6759,N_7105);
and U11199 (N_11199,N_7580,N_8489);
or U11200 (N_11200,N_7993,N_7840);
or U11201 (N_11201,N_6765,N_6737);
and U11202 (N_11202,N_6670,N_8309);
and U11203 (N_11203,N_7652,N_7746);
and U11204 (N_11204,N_8126,N_7079);
or U11205 (N_11205,N_8219,N_7592);
and U11206 (N_11206,N_9203,N_6519);
nor U11207 (N_11207,N_8386,N_7382);
xnor U11208 (N_11208,N_6337,N_8446);
xnor U11209 (N_11209,N_7360,N_6346);
xor U11210 (N_11210,N_6720,N_8950);
and U11211 (N_11211,N_7000,N_7660);
or U11212 (N_11212,N_7386,N_7511);
xnor U11213 (N_11213,N_7552,N_7764);
xnor U11214 (N_11214,N_8295,N_7781);
xnor U11215 (N_11215,N_6356,N_6355);
nor U11216 (N_11216,N_6830,N_6478);
nor U11217 (N_11217,N_8397,N_7775);
and U11218 (N_11218,N_8865,N_8433);
nand U11219 (N_11219,N_9189,N_7440);
and U11220 (N_11220,N_7965,N_8268);
nand U11221 (N_11221,N_7188,N_8696);
and U11222 (N_11222,N_6714,N_7130);
nor U11223 (N_11223,N_6370,N_8337);
nor U11224 (N_11224,N_7587,N_8369);
xnor U11225 (N_11225,N_7197,N_7102);
and U11226 (N_11226,N_6411,N_7161);
and U11227 (N_11227,N_8933,N_7665);
nor U11228 (N_11228,N_6440,N_8924);
or U11229 (N_11229,N_9167,N_7440);
nand U11230 (N_11230,N_6901,N_6542);
or U11231 (N_11231,N_6679,N_6489);
and U11232 (N_11232,N_9372,N_8636);
or U11233 (N_11233,N_6537,N_9003);
or U11234 (N_11234,N_7715,N_9363);
or U11235 (N_11235,N_9098,N_7828);
xor U11236 (N_11236,N_8415,N_9143);
nor U11237 (N_11237,N_7470,N_8748);
xor U11238 (N_11238,N_8516,N_8819);
and U11239 (N_11239,N_8267,N_6785);
and U11240 (N_11240,N_7613,N_8807);
xor U11241 (N_11241,N_6990,N_8289);
or U11242 (N_11242,N_7671,N_8556);
or U11243 (N_11243,N_8025,N_7962);
and U11244 (N_11244,N_7778,N_9042);
nor U11245 (N_11245,N_8775,N_6566);
xor U11246 (N_11246,N_8756,N_8349);
xor U11247 (N_11247,N_6776,N_7952);
and U11248 (N_11248,N_8960,N_7713);
or U11249 (N_11249,N_8885,N_6305);
xor U11250 (N_11250,N_8901,N_8226);
xnor U11251 (N_11251,N_6699,N_9055);
xnor U11252 (N_11252,N_6763,N_6879);
nor U11253 (N_11253,N_6987,N_6749);
nor U11254 (N_11254,N_6305,N_6748);
or U11255 (N_11255,N_8145,N_8650);
xor U11256 (N_11256,N_8781,N_7513);
nand U11257 (N_11257,N_7579,N_8878);
nor U11258 (N_11258,N_8741,N_8704);
and U11259 (N_11259,N_8829,N_9278);
or U11260 (N_11260,N_6587,N_9118);
nor U11261 (N_11261,N_9345,N_7800);
and U11262 (N_11262,N_8018,N_7029);
xor U11263 (N_11263,N_8285,N_7155);
and U11264 (N_11264,N_7749,N_6917);
xnor U11265 (N_11265,N_7905,N_7672);
nor U11266 (N_11266,N_7971,N_6320);
nor U11267 (N_11267,N_6955,N_6990);
nand U11268 (N_11268,N_8928,N_8226);
or U11269 (N_11269,N_9268,N_9161);
and U11270 (N_11270,N_8523,N_6462);
xor U11271 (N_11271,N_9344,N_8767);
xnor U11272 (N_11272,N_8581,N_7811);
nor U11273 (N_11273,N_6625,N_6577);
nand U11274 (N_11274,N_8361,N_8450);
nor U11275 (N_11275,N_7991,N_9199);
and U11276 (N_11276,N_7417,N_6689);
or U11277 (N_11277,N_6699,N_8810);
xnor U11278 (N_11278,N_7556,N_6321);
xor U11279 (N_11279,N_8645,N_7193);
or U11280 (N_11280,N_7835,N_8407);
xor U11281 (N_11281,N_7505,N_8670);
and U11282 (N_11282,N_6690,N_7043);
and U11283 (N_11283,N_8967,N_7822);
nand U11284 (N_11284,N_8717,N_8099);
nor U11285 (N_11285,N_7197,N_7805);
or U11286 (N_11286,N_7795,N_9038);
nor U11287 (N_11287,N_8640,N_8877);
nand U11288 (N_11288,N_8861,N_7178);
or U11289 (N_11289,N_9356,N_9094);
and U11290 (N_11290,N_6637,N_9051);
and U11291 (N_11291,N_9202,N_7104);
nor U11292 (N_11292,N_6590,N_8423);
nor U11293 (N_11293,N_7977,N_9295);
nor U11294 (N_11294,N_8808,N_8380);
nor U11295 (N_11295,N_8200,N_6312);
and U11296 (N_11296,N_7086,N_7177);
xor U11297 (N_11297,N_7501,N_7798);
or U11298 (N_11298,N_8351,N_8762);
or U11299 (N_11299,N_7854,N_6704);
or U11300 (N_11300,N_9012,N_7984);
and U11301 (N_11301,N_7826,N_8999);
or U11302 (N_11302,N_8082,N_8199);
nor U11303 (N_11303,N_8033,N_6839);
and U11304 (N_11304,N_8949,N_6895);
and U11305 (N_11305,N_7267,N_6679);
xor U11306 (N_11306,N_7284,N_7231);
and U11307 (N_11307,N_8317,N_8524);
nand U11308 (N_11308,N_8886,N_7325);
or U11309 (N_11309,N_8558,N_6331);
and U11310 (N_11310,N_7006,N_6624);
nor U11311 (N_11311,N_7370,N_6765);
nand U11312 (N_11312,N_7759,N_6907);
or U11313 (N_11313,N_7122,N_8841);
xnor U11314 (N_11314,N_7894,N_9281);
xnor U11315 (N_11315,N_8603,N_6494);
and U11316 (N_11316,N_8935,N_6373);
nor U11317 (N_11317,N_8809,N_7502);
xnor U11318 (N_11318,N_6848,N_8203);
nor U11319 (N_11319,N_7023,N_8011);
nor U11320 (N_11320,N_8807,N_6334);
nor U11321 (N_11321,N_9009,N_6274);
nand U11322 (N_11322,N_8721,N_7635);
xor U11323 (N_11323,N_7995,N_6548);
and U11324 (N_11324,N_6557,N_8456);
xor U11325 (N_11325,N_8803,N_9036);
and U11326 (N_11326,N_8815,N_6695);
xor U11327 (N_11327,N_7125,N_6835);
nand U11328 (N_11328,N_7685,N_6812);
nand U11329 (N_11329,N_7070,N_8242);
nor U11330 (N_11330,N_8774,N_7447);
xor U11331 (N_11331,N_8685,N_8687);
nand U11332 (N_11332,N_9203,N_7665);
nor U11333 (N_11333,N_9019,N_7722);
nand U11334 (N_11334,N_7288,N_7877);
xor U11335 (N_11335,N_7156,N_6892);
xor U11336 (N_11336,N_6622,N_6955);
nor U11337 (N_11337,N_7368,N_7833);
nand U11338 (N_11338,N_8662,N_9131);
nand U11339 (N_11339,N_6914,N_6533);
nor U11340 (N_11340,N_7917,N_7164);
or U11341 (N_11341,N_7832,N_8375);
and U11342 (N_11342,N_6604,N_7968);
nor U11343 (N_11343,N_8526,N_7372);
and U11344 (N_11344,N_6488,N_9160);
and U11345 (N_11345,N_8123,N_8722);
nor U11346 (N_11346,N_7551,N_9021);
or U11347 (N_11347,N_8056,N_8613);
and U11348 (N_11348,N_7800,N_8763);
nand U11349 (N_11349,N_8627,N_8953);
nor U11350 (N_11350,N_6948,N_8426);
xor U11351 (N_11351,N_9312,N_8139);
nand U11352 (N_11352,N_7426,N_6305);
xnor U11353 (N_11353,N_7665,N_6276);
nand U11354 (N_11354,N_8366,N_9186);
nor U11355 (N_11355,N_8503,N_7956);
and U11356 (N_11356,N_7703,N_7195);
nor U11357 (N_11357,N_8850,N_8910);
xor U11358 (N_11358,N_8709,N_6600);
nand U11359 (N_11359,N_6945,N_8427);
xor U11360 (N_11360,N_9221,N_6474);
nor U11361 (N_11361,N_6491,N_7650);
nand U11362 (N_11362,N_8211,N_7885);
and U11363 (N_11363,N_6422,N_7478);
or U11364 (N_11364,N_7215,N_8287);
or U11365 (N_11365,N_6840,N_6355);
xor U11366 (N_11366,N_8111,N_6439);
and U11367 (N_11367,N_8771,N_8564);
and U11368 (N_11368,N_7032,N_8078);
nor U11369 (N_11369,N_6897,N_7322);
or U11370 (N_11370,N_8429,N_8098);
nand U11371 (N_11371,N_8504,N_8903);
or U11372 (N_11372,N_8863,N_8590);
nor U11373 (N_11373,N_7161,N_7602);
or U11374 (N_11374,N_7506,N_7528);
nand U11375 (N_11375,N_8541,N_6645);
or U11376 (N_11376,N_9281,N_6323);
xnor U11377 (N_11377,N_8909,N_6849);
and U11378 (N_11378,N_8339,N_6959);
or U11379 (N_11379,N_8877,N_6988);
xnor U11380 (N_11380,N_8449,N_6631);
or U11381 (N_11381,N_8334,N_8367);
xor U11382 (N_11382,N_7744,N_7045);
xnor U11383 (N_11383,N_6859,N_7216);
xnor U11384 (N_11384,N_8446,N_7058);
and U11385 (N_11385,N_6602,N_8048);
nand U11386 (N_11386,N_8313,N_6900);
and U11387 (N_11387,N_9161,N_7700);
and U11388 (N_11388,N_7037,N_8216);
nand U11389 (N_11389,N_9198,N_9053);
xor U11390 (N_11390,N_9036,N_9142);
nand U11391 (N_11391,N_7017,N_6324);
nor U11392 (N_11392,N_6313,N_6761);
nor U11393 (N_11393,N_7129,N_7631);
or U11394 (N_11394,N_7959,N_8432);
and U11395 (N_11395,N_7187,N_7341);
xor U11396 (N_11396,N_8572,N_7085);
nand U11397 (N_11397,N_8403,N_7912);
xnor U11398 (N_11398,N_8703,N_6478);
nor U11399 (N_11399,N_9267,N_6413);
nor U11400 (N_11400,N_6405,N_6893);
xor U11401 (N_11401,N_7483,N_8182);
nand U11402 (N_11402,N_6461,N_8693);
or U11403 (N_11403,N_8629,N_9354);
xor U11404 (N_11404,N_8600,N_8113);
nor U11405 (N_11405,N_7741,N_9000);
and U11406 (N_11406,N_9267,N_6520);
or U11407 (N_11407,N_8951,N_8199);
and U11408 (N_11408,N_9168,N_6821);
nand U11409 (N_11409,N_6553,N_7963);
and U11410 (N_11410,N_6263,N_6908);
nand U11411 (N_11411,N_9337,N_8942);
xnor U11412 (N_11412,N_8405,N_6941);
nor U11413 (N_11413,N_6267,N_9065);
or U11414 (N_11414,N_8312,N_6983);
nand U11415 (N_11415,N_7100,N_9292);
or U11416 (N_11416,N_8212,N_7911);
nand U11417 (N_11417,N_8445,N_7100);
nor U11418 (N_11418,N_9039,N_8683);
xnor U11419 (N_11419,N_7713,N_9341);
nand U11420 (N_11420,N_6701,N_8466);
nand U11421 (N_11421,N_7118,N_7895);
nor U11422 (N_11422,N_7888,N_8824);
and U11423 (N_11423,N_7348,N_6571);
nand U11424 (N_11424,N_7435,N_7848);
nor U11425 (N_11425,N_6343,N_8367);
xnor U11426 (N_11426,N_9302,N_7702);
and U11427 (N_11427,N_9232,N_9356);
nand U11428 (N_11428,N_8676,N_6280);
nand U11429 (N_11429,N_8361,N_7287);
and U11430 (N_11430,N_8631,N_6879);
nand U11431 (N_11431,N_7996,N_8773);
and U11432 (N_11432,N_6393,N_7685);
xor U11433 (N_11433,N_8831,N_6473);
nand U11434 (N_11434,N_7666,N_6814);
and U11435 (N_11435,N_7324,N_6381);
xnor U11436 (N_11436,N_8213,N_8799);
and U11437 (N_11437,N_6576,N_7773);
nor U11438 (N_11438,N_7507,N_7542);
nor U11439 (N_11439,N_7402,N_6592);
nor U11440 (N_11440,N_7688,N_8526);
nor U11441 (N_11441,N_7923,N_8060);
nand U11442 (N_11442,N_6607,N_9159);
xor U11443 (N_11443,N_8248,N_8761);
and U11444 (N_11444,N_9079,N_8597);
or U11445 (N_11445,N_8700,N_7623);
nand U11446 (N_11446,N_6784,N_6800);
nor U11447 (N_11447,N_7545,N_6890);
xor U11448 (N_11448,N_7749,N_9186);
nand U11449 (N_11449,N_7352,N_6921);
or U11450 (N_11450,N_6436,N_8681);
nor U11451 (N_11451,N_6270,N_8029);
nand U11452 (N_11452,N_6709,N_7567);
nor U11453 (N_11453,N_8181,N_7770);
and U11454 (N_11454,N_7686,N_6590);
nor U11455 (N_11455,N_9003,N_7435);
or U11456 (N_11456,N_7272,N_7309);
nand U11457 (N_11457,N_8911,N_7999);
and U11458 (N_11458,N_7413,N_8482);
or U11459 (N_11459,N_7997,N_9348);
nand U11460 (N_11460,N_7500,N_6843);
and U11461 (N_11461,N_7996,N_9149);
or U11462 (N_11462,N_8900,N_7109);
nand U11463 (N_11463,N_6889,N_8080);
nor U11464 (N_11464,N_8457,N_7478);
and U11465 (N_11465,N_8378,N_7937);
nor U11466 (N_11466,N_8268,N_7118);
nor U11467 (N_11467,N_9340,N_7732);
nand U11468 (N_11468,N_9153,N_8017);
nand U11469 (N_11469,N_9215,N_6998);
xnor U11470 (N_11470,N_6939,N_7043);
xor U11471 (N_11471,N_9057,N_7444);
nor U11472 (N_11472,N_9174,N_7640);
and U11473 (N_11473,N_7913,N_6928);
nand U11474 (N_11474,N_7532,N_6949);
and U11475 (N_11475,N_6677,N_6462);
or U11476 (N_11476,N_8292,N_8982);
nand U11477 (N_11477,N_7061,N_7579);
nand U11478 (N_11478,N_6655,N_7198);
and U11479 (N_11479,N_8526,N_8765);
and U11480 (N_11480,N_6901,N_7729);
nand U11481 (N_11481,N_6662,N_7864);
and U11482 (N_11482,N_6843,N_7906);
nor U11483 (N_11483,N_6520,N_9081);
and U11484 (N_11484,N_7495,N_7442);
and U11485 (N_11485,N_8795,N_8260);
xnor U11486 (N_11486,N_9220,N_6910);
nand U11487 (N_11487,N_6578,N_8947);
xnor U11488 (N_11488,N_8315,N_7730);
and U11489 (N_11489,N_8034,N_7457);
or U11490 (N_11490,N_8501,N_8275);
nor U11491 (N_11491,N_6798,N_6548);
xor U11492 (N_11492,N_6897,N_7791);
or U11493 (N_11493,N_6847,N_8824);
xnor U11494 (N_11494,N_6645,N_6847);
nor U11495 (N_11495,N_8466,N_7259);
nand U11496 (N_11496,N_7036,N_7445);
xor U11497 (N_11497,N_7406,N_6485);
nand U11498 (N_11498,N_6389,N_7383);
nand U11499 (N_11499,N_8686,N_6751);
and U11500 (N_11500,N_6973,N_8703);
or U11501 (N_11501,N_7808,N_9079);
nand U11502 (N_11502,N_8408,N_7199);
nand U11503 (N_11503,N_9272,N_8452);
nor U11504 (N_11504,N_7380,N_6308);
or U11505 (N_11505,N_6685,N_8066);
and U11506 (N_11506,N_8765,N_9143);
nand U11507 (N_11507,N_8760,N_6348);
nand U11508 (N_11508,N_8246,N_9143);
and U11509 (N_11509,N_8328,N_9341);
and U11510 (N_11510,N_6695,N_7430);
and U11511 (N_11511,N_8660,N_9152);
nand U11512 (N_11512,N_7901,N_8570);
or U11513 (N_11513,N_7752,N_7344);
and U11514 (N_11514,N_6259,N_8397);
or U11515 (N_11515,N_6904,N_7947);
nand U11516 (N_11516,N_8917,N_7913);
nand U11517 (N_11517,N_7714,N_7803);
nor U11518 (N_11518,N_6848,N_8113);
xor U11519 (N_11519,N_7790,N_8853);
or U11520 (N_11520,N_8517,N_8151);
nor U11521 (N_11521,N_7541,N_7960);
xnor U11522 (N_11522,N_7879,N_6646);
nor U11523 (N_11523,N_6628,N_8683);
nand U11524 (N_11524,N_9251,N_7749);
or U11525 (N_11525,N_7328,N_7692);
xnor U11526 (N_11526,N_9067,N_8200);
and U11527 (N_11527,N_8824,N_6910);
xor U11528 (N_11528,N_6372,N_8032);
and U11529 (N_11529,N_8790,N_8915);
nand U11530 (N_11530,N_7069,N_7801);
nor U11531 (N_11531,N_7120,N_8334);
or U11532 (N_11532,N_7401,N_7768);
xnor U11533 (N_11533,N_7642,N_7700);
or U11534 (N_11534,N_8974,N_7632);
nand U11535 (N_11535,N_9123,N_8143);
and U11536 (N_11536,N_6687,N_6914);
nor U11537 (N_11537,N_6874,N_7075);
nand U11538 (N_11538,N_6418,N_8657);
or U11539 (N_11539,N_7244,N_7707);
or U11540 (N_11540,N_8261,N_9336);
xnor U11541 (N_11541,N_9059,N_8743);
nor U11542 (N_11542,N_7329,N_8890);
nand U11543 (N_11543,N_9094,N_8576);
or U11544 (N_11544,N_7830,N_7144);
or U11545 (N_11545,N_7691,N_6709);
xnor U11546 (N_11546,N_6886,N_8068);
or U11547 (N_11547,N_7954,N_7802);
nand U11548 (N_11548,N_8271,N_6939);
nand U11549 (N_11549,N_9306,N_7396);
nand U11550 (N_11550,N_6291,N_8395);
xor U11551 (N_11551,N_7612,N_8385);
and U11552 (N_11552,N_8605,N_9252);
or U11553 (N_11553,N_7895,N_6988);
nor U11554 (N_11554,N_8199,N_8602);
xnor U11555 (N_11555,N_7208,N_7470);
xnor U11556 (N_11556,N_8827,N_6705);
nand U11557 (N_11557,N_8345,N_7436);
and U11558 (N_11558,N_8543,N_7878);
xor U11559 (N_11559,N_8230,N_7892);
and U11560 (N_11560,N_8367,N_6522);
nand U11561 (N_11561,N_7366,N_7023);
nor U11562 (N_11562,N_6371,N_6693);
xor U11563 (N_11563,N_8546,N_8739);
and U11564 (N_11564,N_9202,N_9038);
xor U11565 (N_11565,N_9044,N_7075);
or U11566 (N_11566,N_7440,N_8904);
or U11567 (N_11567,N_7274,N_7929);
or U11568 (N_11568,N_8288,N_6601);
or U11569 (N_11569,N_8117,N_8336);
and U11570 (N_11570,N_7957,N_7204);
or U11571 (N_11571,N_8254,N_8189);
and U11572 (N_11572,N_6780,N_7753);
nor U11573 (N_11573,N_7318,N_8830);
nand U11574 (N_11574,N_8689,N_6287);
or U11575 (N_11575,N_6405,N_6793);
nand U11576 (N_11576,N_8396,N_8143);
or U11577 (N_11577,N_6741,N_8417);
and U11578 (N_11578,N_6418,N_6454);
or U11579 (N_11579,N_7689,N_7130);
or U11580 (N_11580,N_7968,N_7721);
and U11581 (N_11581,N_9052,N_8276);
nand U11582 (N_11582,N_7407,N_7945);
nand U11583 (N_11583,N_6491,N_7271);
or U11584 (N_11584,N_8897,N_7904);
and U11585 (N_11585,N_8320,N_8585);
xor U11586 (N_11586,N_6871,N_8943);
or U11587 (N_11587,N_9346,N_8478);
xor U11588 (N_11588,N_8135,N_7897);
nand U11589 (N_11589,N_8443,N_8717);
nor U11590 (N_11590,N_8009,N_6656);
nand U11591 (N_11591,N_6570,N_6643);
xnor U11592 (N_11592,N_7857,N_6838);
and U11593 (N_11593,N_6767,N_6509);
and U11594 (N_11594,N_9355,N_7989);
nand U11595 (N_11595,N_8485,N_6315);
and U11596 (N_11596,N_6438,N_8826);
xnor U11597 (N_11597,N_9109,N_8364);
nor U11598 (N_11598,N_8546,N_6820);
and U11599 (N_11599,N_7779,N_7083);
nand U11600 (N_11600,N_8275,N_7300);
and U11601 (N_11601,N_8932,N_7081);
xnor U11602 (N_11602,N_7364,N_8130);
nor U11603 (N_11603,N_7877,N_8633);
nand U11604 (N_11604,N_6780,N_9254);
xor U11605 (N_11605,N_7445,N_7955);
or U11606 (N_11606,N_7864,N_6608);
nor U11607 (N_11607,N_7435,N_7800);
and U11608 (N_11608,N_7959,N_9066);
nor U11609 (N_11609,N_8987,N_7895);
or U11610 (N_11610,N_6311,N_7489);
nand U11611 (N_11611,N_7609,N_7991);
nor U11612 (N_11612,N_8418,N_7220);
nand U11613 (N_11613,N_8199,N_8944);
nand U11614 (N_11614,N_8456,N_7470);
nand U11615 (N_11615,N_8307,N_7529);
and U11616 (N_11616,N_6534,N_9286);
nand U11617 (N_11617,N_6274,N_7312);
nand U11618 (N_11618,N_8317,N_6440);
xor U11619 (N_11619,N_6690,N_8842);
xnor U11620 (N_11620,N_7493,N_6889);
nand U11621 (N_11621,N_8768,N_7628);
or U11622 (N_11622,N_9084,N_7926);
or U11623 (N_11623,N_9263,N_6792);
or U11624 (N_11624,N_7325,N_6287);
nand U11625 (N_11625,N_8888,N_6522);
and U11626 (N_11626,N_7697,N_7900);
nor U11627 (N_11627,N_9309,N_6463);
nand U11628 (N_11628,N_7206,N_6720);
xnor U11629 (N_11629,N_8940,N_9071);
and U11630 (N_11630,N_8226,N_7536);
nor U11631 (N_11631,N_8959,N_6633);
or U11632 (N_11632,N_9017,N_9048);
nand U11633 (N_11633,N_6781,N_8986);
nor U11634 (N_11634,N_7344,N_8691);
and U11635 (N_11635,N_8747,N_8454);
and U11636 (N_11636,N_8556,N_7603);
nor U11637 (N_11637,N_8518,N_6595);
nor U11638 (N_11638,N_6252,N_7653);
nor U11639 (N_11639,N_7530,N_8863);
nand U11640 (N_11640,N_8166,N_9003);
or U11641 (N_11641,N_6911,N_7333);
nand U11642 (N_11642,N_8789,N_8890);
nand U11643 (N_11643,N_7894,N_8527);
xnor U11644 (N_11644,N_8769,N_6472);
nand U11645 (N_11645,N_9112,N_8770);
nor U11646 (N_11646,N_7385,N_8481);
or U11647 (N_11647,N_9188,N_6419);
xnor U11648 (N_11648,N_8775,N_7058);
and U11649 (N_11649,N_7930,N_9222);
nand U11650 (N_11650,N_7641,N_8042);
nand U11651 (N_11651,N_6477,N_9341);
nor U11652 (N_11652,N_8306,N_6801);
or U11653 (N_11653,N_7357,N_8630);
nor U11654 (N_11654,N_8691,N_6938);
and U11655 (N_11655,N_7025,N_7257);
nor U11656 (N_11656,N_9099,N_8230);
xor U11657 (N_11657,N_6487,N_8585);
and U11658 (N_11658,N_6405,N_6470);
xor U11659 (N_11659,N_7265,N_6437);
xnor U11660 (N_11660,N_9201,N_7661);
nor U11661 (N_11661,N_6335,N_6858);
and U11662 (N_11662,N_6370,N_8999);
xor U11663 (N_11663,N_8633,N_6895);
nand U11664 (N_11664,N_9306,N_9131);
xor U11665 (N_11665,N_6366,N_7277);
nor U11666 (N_11666,N_7984,N_7238);
and U11667 (N_11667,N_8008,N_7590);
xnor U11668 (N_11668,N_8274,N_6584);
or U11669 (N_11669,N_6690,N_8721);
or U11670 (N_11670,N_7777,N_9141);
and U11671 (N_11671,N_9153,N_7097);
nor U11672 (N_11672,N_8522,N_6930);
or U11673 (N_11673,N_6830,N_7863);
nand U11674 (N_11674,N_6421,N_8600);
or U11675 (N_11675,N_8485,N_6761);
xnor U11676 (N_11676,N_7158,N_8488);
or U11677 (N_11677,N_8415,N_6772);
or U11678 (N_11678,N_8742,N_7977);
or U11679 (N_11679,N_6495,N_7873);
nand U11680 (N_11680,N_9213,N_8147);
or U11681 (N_11681,N_8356,N_8625);
nor U11682 (N_11682,N_6436,N_6844);
xor U11683 (N_11683,N_8990,N_8430);
nand U11684 (N_11684,N_7578,N_6781);
or U11685 (N_11685,N_6712,N_6344);
nor U11686 (N_11686,N_7988,N_6402);
xor U11687 (N_11687,N_6411,N_7232);
xnor U11688 (N_11688,N_9155,N_7992);
xnor U11689 (N_11689,N_6530,N_7976);
nor U11690 (N_11690,N_8279,N_9356);
nor U11691 (N_11691,N_9346,N_8655);
and U11692 (N_11692,N_7663,N_6638);
or U11693 (N_11693,N_8884,N_8686);
xnor U11694 (N_11694,N_7324,N_8581);
nor U11695 (N_11695,N_9040,N_7252);
or U11696 (N_11696,N_6367,N_8905);
and U11697 (N_11697,N_8621,N_8199);
nand U11698 (N_11698,N_8626,N_8449);
nand U11699 (N_11699,N_7924,N_8155);
or U11700 (N_11700,N_7505,N_7250);
xnor U11701 (N_11701,N_8838,N_8752);
and U11702 (N_11702,N_6318,N_6371);
xnor U11703 (N_11703,N_9059,N_7751);
nand U11704 (N_11704,N_8517,N_8677);
and U11705 (N_11705,N_8339,N_6601);
xnor U11706 (N_11706,N_8345,N_6303);
and U11707 (N_11707,N_6650,N_7764);
nand U11708 (N_11708,N_7131,N_7485);
xnor U11709 (N_11709,N_6707,N_8034);
nor U11710 (N_11710,N_8980,N_8896);
nor U11711 (N_11711,N_7474,N_9047);
or U11712 (N_11712,N_8241,N_6602);
or U11713 (N_11713,N_7621,N_7380);
or U11714 (N_11714,N_6560,N_6294);
xor U11715 (N_11715,N_7560,N_8899);
nor U11716 (N_11716,N_8742,N_7745);
nand U11717 (N_11717,N_7663,N_7702);
xnor U11718 (N_11718,N_7116,N_7815);
xor U11719 (N_11719,N_7134,N_8546);
nand U11720 (N_11720,N_6270,N_8788);
or U11721 (N_11721,N_6435,N_6676);
nand U11722 (N_11722,N_8551,N_6292);
nand U11723 (N_11723,N_8401,N_9131);
and U11724 (N_11724,N_8081,N_8009);
xor U11725 (N_11725,N_8670,N_6922);
xnor U11726 (N_11726,N_7056,N_8904);
nand U11727 (N_11727,N_7382,N_7226);
nand U11728 (N_11728,N_7168,N_8478);
and U11729 (N_11729,N_7404,N_8330);
and U11730 (N_11730,N_8553,N_7930);
nor U11731 (N_11731,N_7377,N_6661);
or U11732 (N_11732,N_7051,N_7496);
xor U11733 (N_11733,N_6870,N_8372);
xor U11734 (N_11734,N_7228,N_8059);
xnor U11735 (N_11735,N_6305,N_7192);
and U11736 (N_11736,N_7210,N_9324);
and U11737 (N_11737,N_7794,N_9273);
xor U11738 (N_11738,N_8033,N_7444);
xor U11739 (N_11739,N_7783,N_7798);
nand U11740 (N_11740,N_7000,N_8305);
or U11741 (N_11741,N_6800,N_6829);
and U11742 (N_11742,N_8750,N_6389);
and U11743 (N_11743,N_7152,N_7467);
nand U11744 (N_11744,N_9002,N_8603);
nand U11745 (N_11745,N_7122,N_7516);
nand U11746 (N_11746,N_6853,N_7552);
xnor U11747 (N_11747,N_7017,N_6412);
nor U11748 (N_11748,N_8253,N_8033);
nand U11749 (N_11749,N_7771,N_8377);
or U11750 (N_11750,N_7928,N_7007);
xnor U11751 (N_11751,N_8612,N_7379);
or U11752 (N_11752,N_8233,N_7918);
and U11753 (N_11753,N_8973,N_7403);
nand U11754 (N_11754,N_8615,N_7477);
nand U11755 (N_11755,N_7777,N_7904);
nand U11756 (N_11756,N_8694,N_7959);
nor U11757 (N_11757,N_8605,N_9354);
xnor U11758 (N_11758,N_6564,N_9222);
and U11759 (N_11759,N_7348,N_6592);
or U11760 (N_11760,N_7613,N_8564);
or U11761 (N_11761,N_6581,N_8972);
nand U11762 (N_11762,N_8193,N_8355);
nand U11763 (N_11763,N_8611,N_7818);
nor U11764 (N_11764,N_7588,N_7114);
and U11765 (N_11765,N_9174,N_9038);
and U11766 (N_11766,N_7665,N_6350);
nand U11767 (N_11767,N_7152,N_7511);
and U11768 (N_11768,N_7717,N_7640);
and U11769 (N_11769,N_8271,N_8533);
nand U11770 (N_11770,N_7886,N_7304);
or U11771 (N_11771,N_7884,N_8838);
and U11772 (N_11772,N_9340,N_8460);
nand U11773 (N_11773,N_9047,N_8680);
or U11774 (N_11774,N_6279,N_7682);
or U11775 (N_11775,N_8598,N_6361);
or U11776 (N_11776,N_7122,N_8861);
and U11777 (N_11777,N_9156,N_7534);
nand U11778 (N_11778,N_7936,N_8629);
nand U11779 (N_11779,N_8053,N_8136);
xnor U11780 (N_11780,N_7974,N_7044);
and U11781 (N_11781,N_8860,N_8505);
and U11782 (N_11782,N_7848,N_8098);
xor U11783 (N_11783,N_7910,N_7843);
xnor U11784 (N_11784,N_7557,N_7204);
and U11785 (N_11785,N_7308,N_7526);
nor U11786 (N_11786,N_8815,N_7991);
nand U11787 (N_11787,N_8223,N_7404);
nor U11788 (N_11788,N_8729,N_8172);
nor U11789 (N_11789,N_8184,N_8453);
or U11790 (N_11790,N_9086,N_6651);
nand U11791 (N_11791,N_9091,N_7224);
nor U11792 (N_11792,N_6780,N_8529);
xnor U11793 (N_11793,N_8165,N_6485);
nor U11794 (N_11794,N_8387,N_7207);
or U11795 (N_11795,N_6774,N_7466);
or U11796 (N_11796,N_6406,N_8332);
and U11797 (N_11797,N_6999,N_8320);
nand U11798 (N_11798,N_8157,N_9013);
and U11799 (N_11799,N_7983,N_7465);
or U11800 (N_11800,N_7714,N_8468);
or U11801 (N_11801,N_6528,N_9281);
and U11802 (N_11802,N_6860,N_8056);
nand U11803 (N_11803,N_8317,N_6704);
and U11804 (N_11804,N_9271,N_8236);
nand U11805 (N_11805,N_6314,N_9334);
xor U11806 (N_11806,N_7957,N_8246);
or U11807 (N_11807,N_9343,N_7711);
nand U11808 (N_11808,N_8107,N_6577);
nand U11809 (N_11809,N_7378,N_6682);
xor U11810 (N_11810,N_6844,N_8376);
or U11811 (N_11811,N_8445,N_7990);
and U11812 (N_11812,N_8527,N_7835);
nand U11813 (N_11813,N_8526,N_7204);
or U11814 (N_11814,N_7075,N_9039);
and U11815 (N_11815,N_6577,N_9217);
or U11816 (N_11816,N_7863,N_7743);
or U11817 (N_11817,N_6686,N_8015);
nor U11818 (N_11818,N_7281,N_6567);
and U11819 (N_11819,N_6990,N_7482);
or U11820 (N_11820,N_8580,N_7754);
nor U11821 (N_11821,N_6919,N_6769);
xor U11822 (N_11822,N_7142,N_7514);
xor U11823 (N_11823,N_8822,N_6450);
and U11824 (N_11824,N_6435,N_6288);
nand U11825 (N_11825,N_9130,N_6282);
and U11826 (N_11826,N_7423,N_7379);
xnor U11827 (N_11827,N_6865,N_7117);
xor U11828 (N_11828,N_7246,N_7248);
nor U11829 (N_11829,N_6678,N_7453);
nand U11830 (N_11830,N_6493,N_8308);
xor U11831 (N_11831,N_6781,N_8343);
xnor U11832 (N_11832,N_8979,N_6270);
and U11833 (N_11833,N_9278,N_7786);
nor U11834 (N_11834,N_8261,N_8052);
nor U11835 (N_11835,N_6740,N_8553);
and U11836 (N_11836,N_7512,N_9234);
xnor U11837 (N_11837,N_8877,N_6498);
nand U11838 (N_11838,N_9167,N_8200);
nor U11839 (N_11839,N_7745,N_6728);
nand U11840 (N_11840,N_7044,N_8306);
xor U11841 (N_11841,N_7239,N_8183);
and U11842 (N_11842,N_8884,N_7469);
nand U11843 (N_11843,N_8782,N_6595);
nand U11844 (N_11844,N_7634,N_8832);
and U11845 (N_11845,N_6299,N_8944);
or U11846 (N_11846,N_6406,N_8543);
nor U11847 (N_11847,N_7706,N_6271);
and U11848 (N_11848,N_7564,N_7572);
nand U11849 (N_11849,N_8141,N_7168);
or U11850 (N_11850,N_6941,N_8288);
or U11851 (N_11851,N_8585,N_6363);
xor U11852 (N_11852,N_6601,N_8218);
and U11853 (N_11853,N_7917,N_8416);
and U11854 (N_11854,N_9227,N_7000);
or U11855 (N_11855,N_7793,N_9108);
and U11856 (N_11856,N_7552,N_7885);
and U11857 (N_11857,N_7346,N_7314);
and U11858 (N_11858,N_8563,N_7145);
xnor U11859 (N_11859,N_8769,N_7102);
and U11860 (N_11860,N_7075,N_7541);
or U11861 (N_11861,N_6301,N_7576);
nor U11862 (N_11862,N_9170,N_6586);
nor U11863 (N_11863,N_6395,N_7636);
xor U11864 (N_11864,N_7965,N_9199);
and U11865 (N_11865,N_8884,N_8648);
nor U11866 (N_11866,N_8960,N_6414);
and U11867 (N_11867,N_7969,N_9281);
nand U11868 (N_11868,N_7964,N_6516);
nor U11869 (N_11869,N_7046,N_6644);
or U11870 (N_11870,N_8075,N_8398);
and U11871 (N_11871,N_8832,N_7504);
and U11872 (N_11872,N_8746,N_7945);
xnor U11873 (N_11873,N_6888,N_8767);
xnor U11874 (N_11874,N_8423,N_6756);
nor U11875 (N_11875,N_7898,N_6934);
nor U11876 (N_11876,N_6698,N_7681);
nand U11877 (N_11877,N_7787,N_9326);
nand U11878 (N_11878,N_6781,N_8616);
nand U11879 (N_11879,N_8549,N_7717);
nor U11880 (N_11880,N_9156,N_7216);
or U11881 (N_11881,N_9280,N_9362);
nand U11882 (N_11882,N_8448,N_8718);
nand U11883 (N_11883,N_8048,N_6630);
xor U11884 (N_11884,N_8121,N_8260);
xor U11885 (N_11885,N_9256,N_6824);
and U11886 (N_11886,N_8971,N_8725);
or U11887 (N_11887,N_7214,N_8826);
xor U11888 (N_11888,N_8381,N_7829);
xnor U11889 (N_11889,N_6609,N_9032);
or U11890 (N_11890,N_7762,N_8946);
nand U11891 (N_11891,N_6985,N_8744);
nand U11892 (N_11892,N_8623,N_8466);
xor U11893 (N_11893,N_8238,N_8644);
and U11894 (N_11894,N_7068,N_6252);
nand U11895 (N_11895,N_9282,N_8972);
nor U11896 (N_11896,N_6953,N_6651);
and U11897 (N_11897,N_7298,N_9372);
nor U11898 (N_11898,N_7695,N_6634);
or U11899 (N_11899,N_7974,N_7771);
and U11900 (N_11900,N_7041,N_8262);
nand U11901 (N_11901,N_8945,N_6668);
nand U11902 (N_11902,N_8371,N_7885);
nand U11903 (N_11903,N_8469,N_6299);
or U11904 (N_11904,N_6620,N_7476);
xor U11905 (N_11905,N_6506,N_6866);
nand U11906 (N_11906,N_6288,N_8059);
nor U11907 (N_11907,N_7015,N_9299);
xor U11908 (N_11908,N_8269,N_8117);
and U11909 (N_11909,N_7806,N_8529);
nand U11910 (N_11910,N_8139,N_7894);
nand U11911 (N_11911,N_8485,N_6460);
and U11912 (N_11912,N_6673,N_6869);
xnor U11913 (N_11913,N_6339,N_7324);
xor U11914 (N_11914,N_9244,N_6602);
nand U11915 (N_11915,N_7903,N_7675);
xor U11916 (N_11916,N_9337,N_8198);
xor U11917 (N_11917,N_9046,N_6787);
or U11918 (N_11918,N_6405,N_8365);
xnor U11919 (N_11919,N_6688,N_6859);
and U11920 (N_11920,N_8888,N_6828);
or U11921 (N_11921,N_9179,N_7574);
nand U11922 (N_11922,N_7149,N_8940);
nor U11923 (N_11923,N_7919,N_8455);
and U11924 (N_11924,N_8232,N_9365);
or U11925 (N_11925,N_7559,N_8450);
and U11926 (N_11926,N_9359,N_9086);
xnor U11927 (N_11927,N_9341,N_6874);
or U11928 (N_11928,N_9055,N_9049);
nor U11929 (N_11929,N_7560,N_7531);
or U11930 (N_11930,N_7757,N_7702);
and U11931 (N_11931,N_7412,N_6345);
nand U11932 (N_11932,N_7476,N_7765);
nand U11933 (N_11933,N_6907,N_7832);
or U11934 (N_11934,N_8987,N_7694);
nor U11935 (N_11935,N_8054,N_6737);
or U11936 (N_11936,N_8050,N_6417);
and U11937 (N_11937,N_7422,N_7232);
nor U11938 (N_11938,N_8188,N_6710);
xnor U11939 (N_11939,N_8014,N_6535);
or U11940 (N_11940,N_9338,N_7352);
nand U11941 (N_11941,N_6814,N_8062);
xor U11942 (N_11942,N_8054,N_7356);
nand U11943 (N_11943,N_6810,N_7694);
and U11944 (N_11944,N_7751,N_9209);
and U11945 (N_11945,N_7159,N_6709);
xor U11946 (N_11946,N_7217,N_9035);
xnor U11947 (N_11947,N_8253,N_6463);
xor U11948 (N_11948,N_9171,N_6545);
nand U11949 (N_11949,N_7972,N_8472);
and U11950 (N_11950,N_6637,N_6830);
xor U11951 (N_11951,N_9252,N_8398);
nor U11952 (N_11952,N_6568,N_9163);
or U11953 (N_11953,N_7968,N_6373);
nor U11954 (N_11954,N_6792,N_7385);
and U11955 (N_11955,N_7742,N_9045);
nand U11956 (N_11956,N_8401,N_6381);
or U11957 (N_11957,N_7056,N_7084);
or U11958 (N_11958,N_7997,N_6334);
nand U11959 (N_11959,N_7759,N_8927);
xnor U11960 (N_11960,N_7230,N_7631);
nor U11961 (N_11961,N_9348,N_8595);
or U11962 (N_11962,N_8558,N_8912);
nor U11963 (N_11963,N_6636,N_8043);
xor U11964 (N_11964,N_7660,N_7306);
nand U11965 (N_11965,N_7313,N_6656);
nor U11966 (N_11966,N_6805,N_7915);
xnor U11967 (N_11967,N_7307,N_8879);
nand U11968 (N_11968,N_7544,N_7887);
and U11969 (N_11969,N_8870,N_6743);
nand U11970 (N_11970,N_7444,N_7442);
xnor U11971 (N_11971,N_7608,N_8796);
nor U11972 (N_11972,N_9161,N_6670);
xnor U11973 (N_11973,N_6350,N_6519);
or U11974 (N_11974,N_9371,N_8642);
xnor U11975 (N_11975,N_7114,N_6302);
or U11976 (N_11976,N_7615,N_8183);
nor U11977 (N_11977,N_9271,N_8198);
nor U11978 (N_11978,N_7475,N_6693);
xnor U11979 (N_11979,N_9305,N_8108);
and U11980 (N_11980,N_9019,N_6788);
and U11981 (N_11981,N_8753,N_8254);
nand U11982 (N_11982,N_7107,N_7174);
nor U11983 (N_11983,N_9181,N_7170);
or U11984 (N_11984,N_6662,N_6512);
nor U11985 (N_11985,N_6303,N_6966);
xnor U11986 (N_11986,N_6356,N_6598);
or U11987 (N_11987,N_7457,N_8930);
and U11988 (N_11988,N_8045,N_7642);
nand U11989 (N_11989,N_8547,N_6844);
xor U11990 (N_11990,N_8161,N_6592);
or U11991 (N_11991,N_6821,N_7684);
xnor U11992 (N_11992,N_6527,N_7044);
nor U11993 (N_11993,N_6890,N_8048);
nor U11994 (N_11994,N_7068,N_8048);
or U11995 (N_11995,N_8893,N_7697);
and U11996 (N_11996,N_6749,N_8387);
xor U11997 (N_11997,N_7698,N_6464);
xnor U11998 (N_11998,N_6386,N_8679);
and U11999 (N_11999,N_8811,N_6425);
or U12000 (N_12000,N_7771,N_8684);
nand U12001 (N_12001,N_7180,N_7073);
xor U12002 (N_12002,N_9010,N_7298);
and U12003 (N_12003,N_9165,N_8695);
and U12004 (N_12004,N_6425,N_8474);
xor U12005 (N_12005,N_7695,N_8225);
xnor U12006 (N_12006,N_8711,N_8926);
and U12007 (N_12007,N_8174,N_6812);
nand U12008 (N_12008,N_9306,N_8414);
xor U12009 (N_12009,N_7204,N_7935);
nand U12010 (N_12010,N_7002,N_6848);
or U12011 (N_12011,N_7173,N_7549);
nand U12012 (N_12012,N_9367,N_8567);
xor U12013 (N_12013,N_9203,N_7848);
nor U12014 (N_12014,N_9135,N_9070);
nor U12015 (N_12015,N_9176,N_6937);
or U12016 (N_12016,N_7818,N_7759);
or U12017 (N_12017,N_8660,N_8620);
xor U12018 (N_12018,N_8007,N_8714);
or U12019 (N_12019,N_8486,N_8535);
nand U12020 (N_12020,N_8167,N_9173);
nand U12021 (N_12021,N_8506,N_6467);
nand U12022 (N_12022,N_8082,N_6388);
and U12023 (N_12023,N_7291,N_6425);
nand U12024 (N_12024,N_6709,N_8674);
xnor U12025 (N_12025,N_8678,N_9112);
nand U12026 (N_12026,N_8721,N_8486);
or U12027 (N_12027,N_9274,N_6810);
nand U12028 (N_12028,N_7374,N_7021);
nor U12029 (N_12029,N_9232,N_6894);
or U12030 (N_12030,N_6902,N_7927);
nor U12031 (N_12031,N_8934,N_9209);
nor U12032 (N_12032,N_7283,N_6588);
and U12033 (N_12033,N_7894,N_8082);
xnor U12034 (N_12034,N_6484,N_7255);
nor U12035 (N_12035,N_8198,N_6533);
and U12036 (N_12036,N_8457,N_8799);
nor U12037 (N_12037,N_8269,N_7882);
nand U12038 (N_12038,N_7867,N_6468);
and U12039 (N_12039,N_6748,N_7457);
and U12040 (N_12040,N_7387,N_6946);
nor U12041 (N_12041,N_6387,N_8060);
xnor U12042 (N_12042,N_7668,N_7115);
xnor U12043 (N_12043,N_8915,N_8611);
and U12044 (N_12044,N_9160,N_6858);
nand U12045 (N_12045,N_8262,N_6472);
xnor U12046 (N_12046,N_7323,N_8311);
or U12047 (N_12047,N_6527,N_8319);
and U12048 (N_12048,N_6526,N_8916);
and U12049 (N_12049,N_9260,N_7032);
xor U12050 (N_12050,N_7352,N_9134);
nand U12051 (N_12051,N_7512,N_6840);
nor U12052 (N_12052,N_8185,N_7174);
nand U12053 (N_12053,N_7291,N_6465);
xnor U12054 (N_12054,N_7438,N_8902);
or U12055 (N_12055,N_8495,N_7938);
or U12056 (N_12056,N_7234,N_9316);
or U12057 (N_12057,N_8615,N_8144);
xnor U12058 (N_12058,N_8153,N_8163);
and U12059 (N_12059,N_9133,N_9153);
nor U12060 (N_12060,N_7280,N_8532);
xnor U12061 (N_12061,N_6607,N_8558);
nor U12062 (N_12062,N_7525,N_6904);
nand U12063 (N_12063,N_8728,N_8376);
nor U12064 (N_12064,N_9251,N_6897);
nand U12065 (N_12065,N_8688,N_7797);
or U12066 (N_12066,N_8696,N_7670);
or U12067 (N_12067,N_8218,N_6359);
nand U12068 (N_12068,N_8251,N_8739);
nand U12069 (N_12069,N_8340,N_7123);
nor U12070 (N_12070,N_7602,N_7490);
xor U12071 (N_12071,N_7081,N_9138);
xnor U12072 (N_12072,N_6268,N_7194);
or U12073 (N_12073,N_7696,N_6411);
or U12074 (N_12074,N_6855,N_8661);
nor U12075 (N_12075,N_6362,N_7729);
or U12076 (N_12076,N_7404,N_7739);
xnor U12077 (N_12077,N_7214,N_7929);
or U12078 (N_12078,N_6737,N_8015);
or U12079 (N_12079,N_7924,N_8104);
nor U12080 (N_12080,N_7607,N_8616);
nor U12081 (N_12081,N_7406,N_7678);
and U12082 (N_12082,N_6851,N_9120);
nand U12083 (N_12083,N_8576,N_8903);
and U12084 (N_12084,N_8816,N_7540);
nand U12085 (N_12085,N_7592,N_8208);
xor U12086 (N_12086,N_6494,N_7204);
nand U12087 (N_12087,N_8026,N_7613);
xnor U12088 (N_12088,N_6679,N_7224);
nor U12089 (N_12089,N_6634,N_7078);
nor U12090 (N_12090,N_7176,N_7586);
and U12091 (N_12091,N_7908,N_7084);
nand U12092 (N_12092,N_7364,N_8258);
or U12093 (N_12093,N_7275,N_7265);
and U12094 (N_12094,N_8113,N_8243);
or U12095 (N_12095,N_6729,N_8705);
nor U12096 (N_12096,N_7799,N_8137);
nand U12097 (N_12097,N_7829,N_8252);
xor U12098 (N_12098,N_6425,N_6635);
nor U12099 (N_12099,N_6921,N_8784);
nor U12100 (N_12100,N_7421,N_7939);
or U12101 (N_12101,N_8478,N_7669);
and U12102 (N_12102,N_8698,N_8351);
nor U12103 (N_12103,N_8082,N_7867);
nor U12104 (N_12104,N_6823,N_6529);
or U12105 (N_12105,N_8874,N_8096);
nand U12106 (N_12106,N_8349,N_6532);
or U12107 (N_12107,N_8132,N_7597);
nand U12108 (N_12108,N_7792,N_9041);
nand U12109 (N_12109,N_8709,N_8848);
xor U12110 (N_12110,N_7229,N_8257);
xnor U12111 (N_12111,N_7739,N_9245);
or U12112 (N_12112,N_6379,N_8528);
or U12113 (N_12113,N_6591,N_6788);
and U12114 (N_12114,N_6619,N_8152);
xnor U12115 (N_12115,N_7745,N_7964);
nor U12116 (N_12116,N_6361,N_9176);
nor U12117 (N_12117,N_8660,N_7511);
nand U12118 (N_12118,N_7218,N_6690);
nor U12119 (N_12119,N_8239,N_7686);
and U12120 (N_12120,N_8905,N_7188);
and U12121 (N_12121,N_8786,N_6765);
and U12122 (N_12122,N_8478,N_9106);
nand U12123 (N_12123,N_7485,N_7701);
nor U12124 (N_12124,N_6715,N_8691);
xor U12125 (N_12125,N_6654,N_6525);
xor U12126 (N_12126,N_8410,N_6709);
or U12127 (N_12127,N_7537,N_7345);
nand U12128 (N_12128,N_6341,N_7369);
xnor U12129 (N_12129,N_7607,N_7853);
or U12130 (N_12130,N_8423,N_8706);
and U12131 (N_12131,N_8617,N_9082);
and U12132 (N_12132,N_9189,N_7228);
nand U12133 (N_12133,N_8468,N_7823);
xor U12134 (N_12134,N_7645,N_7616);
xnor U12135 (N_12135,N_8062,N_6958);
xnor U12136 (N_12136,N_8698,N_7022);
nand U12137 (N_12137,N_8939,N_8943);
or U12138 (N_12138,N_7835,N_7258);
nand U12139 (N_12139,N_7382,N_8403);
and U12140 (N_12140,N_7421,N_6834);
xor U12141 (N_12141,N_6499,N_8153);
nand U12142 (N_12142,N_6469,N_6608);
and U12143 (N_12143,N_7716,N_6400);
or U12144 (N_12144,N_9184,N_7564);
or U12145 (N_12145,N_6987,N_6577);
and U12146 (N_12146,N_9157,N_7973);
or U12147 (N_12147,N_6541,N_8288);
nand U12148 (N_12148,N_8916,N_9193);
xor U12149 (N_12149,N_8922,N_7866);
and U12150 (N_12150,N_8738,N_6912);
and U12151 (N_12151,N_8863,N_6455);
nor U12152 (N_12152,N_7067,N_7506);
or U12153 (N_12153,N_8372,N_6714);
nand U12154 (N_12154,N_7689,N_7643);
or U12155 (N_12155,N_7928,N_6663);
nor U12156 (N_12156,N_8838,N_8776);
or U12157 (N_12157,N_9043,N_9365);
xor U12158 (N_12158,N_7173,N_8069);
nand U12159 (N_12159,N_9247,N_6686);
nand U12160 (N_12160,N_7918,N_8377);
xor U12161 (N_12161,N_7317,N_7578);
nand U12162 (N_12162,N_6644,N_7064);
nor U12163 (N_12163,N_8601,N_6684);
nand U12164 (N_12164,N_7413,N_6499);
nand U12165 (N_12165,N_7662,N_9091);
nor U12166 (N_12166,N_8254,N_7232);
and U12167 (N_12167,N_7289,N_8788);
xnor U12168 (N_12168,N_7225,N_8966);
or U12169 (N_12169,N_7559,N_7967);
nor U12170 (N_12170,N_7278,N_9268);
xnor U12171 (N_12171,N_7851,N_6980);
nand U12172 (N_12172,N_8352,N_6748);
xnor U12173 (N_12173,N_6561,N_9114);
or U12174 (N_12174,N_9256,N_6320);
and U12175 (N_12175,N_7265,N_7786);
nand U12176 (N_12176,N_6932,N_9323);
and U12177 (N_12177,N_8381,N_9333);
and U12178 (N_12178,N_6292,N_7588);
nand U12179 (N_12179,N_7087,N_8725);
or U12180 (N_12180,N_6720,N_7153);
and U12181 (N_12181,N_8301,N_7844);
or U12182 (N_12182,N_9354,N_6585);
or U12183 (N_12183,N_6549,N_8765);
nand U12184 (N_12184,N_7310,N_6261);
and U12185 (N_12185,N_7015,N_8265);
and U12186 (N_12186,N_6650,N_7890);
and U12187 (N_12187,N_6390,N_7158);
nor U12188 (N_12188,N_9075,N_7832);
nand U12189 (N_12189,N_7311,N_9165);
and U12190 (N_12190,N_9160,N_9122);
nor U12191 (N_12191,N_9064,N_8626);
or U12192 (N_12192,N_6728,N_7975);
nand U12193 (N_12193,N_7724,N_7389);
xor U12194 (N_12194,N_8028,N_8873);
nand U12195 (N_12195,N_7993,N_7568);
xnor U12196 (N_12196,N_9197,N_6474);
xor U12197 (N_12197,N_8924,N_8946);
nand U12198 (N_12198,N_8435,N_8406);
xor U12199 (N_12199,N_7155,N_7583);
xor U12200 (N_12200,N_6638,N_7240);
nor U12201 (N_12201,N_8499,N_6979);
nor U12202 (N_12202,N_9242,N_9160);
nand U12203 (N_12203,N_7817,N_9321);
nor U12204 (N_12204,N_9324,N_9105);
and U12205 (N_12205,N_7616,N_8674);
xnor U12206 (N_12206,N_8487,N_6659);
and U12207 (N_12207,N_8981,N_6702);
xnor U12208 (N_12208,N_7990,N_8345);
or U12209 (N_12209,N_6279,N_6694);
nor U12210 (N_12210,N_9204,N_6502);
xnor U12211 (N_12211,N_7790,N_7741);
nor U12212 (N_12212,N_8592,N_8024);
or U12213 (N_12213,N_7973,N_6644);
nand U12214 (N_12214,N_7311,N_8479);
nand U12215 (N_12215,N_9267,N_7226);
and U12216 (N_12216,N_7508,N_6683);
nand U12217 (N_12217,N_7043,N_6251);
nor U12218 (N_12218,N_8117,N_6370);
xor U12219 (N_12219,N_9020,N_9313);
and U12220 (N_12220,N_8990,N_9202);
nor U12221 (N_12221,N_7570,N_9002);
nand U12222 (N_12222,N_6714,N_9017);
and U12223 (N_12223,N_6710,N_7394);
nand U12224 (N_12224,N_7456,N_6341);
nand U12225 (N_12225,N_8558,N_9289);
nand U12226 (N_12226,N_9115,N_7169);
or U12227 (N_12227,N_7181,N_7843);
nand U12228 (N_12228,N_7288,N_9357);
or U12229 (N_12229,N_8143,N_7476);
nand U12230 (N_12230,N_7079,N_7541);
nand U12231 (N_12231,N_8385,N_7119);
nor U12232 (N_12232,N_6759,N_7365);
xnor U12233 (N_12233,N_7001,N_8531);
nor U12234 (N_12234,N_7202,N_6295);
xnor U12235 (N_12235,N_6576,N_8166);
nand U12236 (N_12236,N_8808,N_9158);
nand U12237 (N_12237,N_8998,N_6732);
nand U12238 (N_12238,N_7871,N_9141);
nand U12239 (N_12239,N_7501,N_8155);
or U12240 (N_12240,N_6313,N_8984);
xor U12241 (N_12241,N_7000,N_6560);
and U12242 (N_12242,N_7114,N_7315);
nor U12243 (N_12243,N_7043,N_8497);
nor U12244 (N_12244,N_6772,N_8126);
nor U12245 (N_12245,N_7329,N_8569);
nor U12246 (N_12246,N_9137,N_8242);
or U12247 (N_12247,N_8245,N_7280);
xnor U12248 (N_12248,N_8001,N_8778);
nor U12249 (N_12249,N_6513,N_8238);
xor U12250 (N_12250,N_7131,N_9230);
nand U12251 (N_12251,N_6767,N_8465);
xnor U12252 (N_12252,N_8078,N_8373);
nand U12253 (N_12253,N_7059,N_8347);
and U12254 (N_12254,N_7897,N_9102);
nand U12255 (N_12255,N_7979,N_8365);
nor U12256 (N_12256,N_7200,N_6478);
nand U12257 (N_12257,N_8269,N_9318);
nand U12258 (N_12258,N_6259,N_8917);
nand U12259 (N_12259,N_9177,N_7434);
nor U12260 (N_12260,N_6389,N_7114);
nand U12261 (N_12261,N_8569,N_6594);
and U12262 (N_12262,N_8347,N_7372);
xnor U12263 (N_12263,N_6579,N_9088);
xnor U12264 (N_12264,N_8179,N_8671);
or U12265 (N_12265,N_8351,N_6371);
nand U12266 (N_12266,N_6322,N_8740);
nand U12267 (N_12267,N_7101,N_8223);
nand U12268 (N_12268,N_9081,N_6588);
or U12269 (N_12269,N_8804,N_6308);
or U12270 (N_12270,N_6342,N_7211);
nand U12271 (N_12271,N_7661,N_7197);
or U12272 (N_12272,N_8072,N_7745);
xor U12273 (N_12273,N_8962,N_6855);
nand U12274 (N_12274,N_9161,N_9226);
nand U12275 (N_12275,N_7719,N_7932);
or U12276 (N_12276,N_8007,N_6899);
nand U12277 (N_12277,N_9254,N_7324);
or U12278 (N_12278,N_7273,N_9365);
xor U12279 (N_12279,N_8466,N_6939);
nor U12280 (N_12280,N_8365,N_8955);
and U12281 (N_12281,N_7402,N_8461);
xor U12282 (N_12282,N_9315,N_6331);
xnor U12283 (N_12283,N_8082,N_8980);
and U12284 (N_12284,N_7686,N_6618);
or U12285 (N_12285,N_6312,N_8275);
or U12286 (N_12286,N_7097,N_9103);
nor U12287 (N_12287,N_7951,N_7979);
or U12288 (N_12288,N_7858,N_8490);
and U12289 (N_12289,N_6294,N_7861);
or U12290 (N_12290,N_7109,N_7381);
or U12291 (N_12291,N_7274,N_7375);
or U12292 (N_12292,N_7103,N_7327);
xor U12293 (N_12293,N_7441,N_8062);
and U12294 (N_12294,N_8028,N_8391);
or U12295 (N_12295,N_6685,N_6378);
or U12296 (N_12296,N_9193,N_7372);
nor U12297 (N_12297,N_8351,N_9202);
nor U12298 (N_12298,N_8808,N_6821);
and U12299 (N_12299,N_8848,N_6571);
or U12300 (N_12300,N_8777,N_8994);
xnor U12301 (N_12301,N_9007,N_7322);
and U12302 (N_12302,N_8806,N_7141);
or U12303 (N_12303,N_8494,N_8156);
nor U12304 (N_12304,N_6648,N_6566);
xnor U12305 (N_12305,N_6845,N_8876);
nand U12306 (N_12306,N_8659,N_7419);
nor U12307 (N_12307,N_7203,N_8763);
nand U12308 (N_12308,N_9166,N_7179);
nor U12309 (N_12309,N_8724,N_9363);
nor U12310 (N_12310,N_8705,N_6365);
xor U12311 (N_12311,N_6398,N_8618);
and U12312 (N_12312,N_7343,N_6695);
xnor U12313 (N_12313,N_6995,N_8726);
nand U12314 (N_12314,N_7151,N_7607);
and U12315 (N_12315,N_7898,N_7047);
or U12316 (N_12316,N_7655,N_8592);
nand U12317 (N_12317,N_8072,N_6822);
nor U12318 (N_12318,N_7843,N_6306);
xor U12319 (N_12319,N_7078,N_9046);
xnor U12320 (N_12320,N_7302,N_6269);
or U12321 (N_12321,N_6377,N_6579);
xnor U12322 (N_12322,N_9047,N_9354);
and U12323 (N_12323,N_7707,N_8099);
xor U12324 (N_12324,N_7136,N_6704);
or U12325 (N_12325,N_6861,N_7319);
or U12326 (N_12326,N_6523,N_6377);
and U12327 (N_12327,N_6569,N_7166);
nor U12328 (N_12328,N_9083,N_8135);
and U12329 (N_12329,N_8026,N_6375);
xor U12330 (N_12330,N_9209,N_7681);
or U12331 (N_12331,N_6327,N_8429);
or U12332 (N_12332,N_8709,N_7749);
or U12333 (N_12333,N_7587,N_7596);
nor U12334 (N_12334,N_9304,N_7947);
and U12335 (N_12335,N_8669,N_7868);
and U12336 (N_12336,N_6310,N_6439);
or U12337 (N_12337,N_8948,N_8843);
nand U12338 (N_12338,N_6862,N_8646);
nand U12339 (N_12339,N_7295,N_8478);
xor U12340 (N_12340,N_9261,N_6279);
nand U12341 (N_12341,N_8940,N_8637);
and U12342 (N_12342,N_6295,N_9055);
nand U12343 (N_12343,N_8944,N_8925);
nand U12344 (N_12344,N_7270,N_7121);
or U12345 (N_12345,N_7698,N_8011);
or U12346 (N_12346,N_8300,N_9314);
xor U12347 (N_12347,N_8331,N_7812);
nor U12348 (N_12348,N_8022,N_8375);
nand U12349 (N_12349,N_7446,N_8947);
or U12350 (N_12350,N_8114,N_7762);
nor U12351 (N_12351,N_6563,N_8862);
and U12352 (N_12352,N_6905,N_7749);
xnor U12353 (N_12353,N_9363,N_8103);
nor U12354 (N_12354,N_9327,N_7271);
or U12355 (N_12355,N_7110,N_7941);
and U12356 (N_12356,N_6384,N_8912);
nor U12357 (N_12357,N_8885,N_6987);
and U12358 (N_12358,N_8117,N_8728);
and U12359 (N_12359,N_8848,N_8445);
or U12360 (N_12360,N_8794,N_6583);
and U12361 (N_12361,N_8402,N_6405);
and U12362 (N_12362,N_6941,N_8336);
nand U12363 (N_12363,N_7624,N_8479);
nor U12364 (N_12364,N_6731,N_9363);
nor U12365 (N_12365,N_8284,N_6272);
nand U12366 (N_12366,N_8587,N_8699);
xnor U12367 (N_12367,N_7808,N_6300);
or U12368 (N_12368,N_8264,N_7087);
or U12369 (N_12369,N_8718,N_6961);
nand U12370 (N_12370,N_7542,N_7980);
or U12371 (N_12371,N_6531,N_8477);
nor U12372 (N_12372,N_8458,N_8441);
xnor U12373 (N_12373,N_9057,N_6309);
nor U12374 (N_12374,N_8716,N_7924);
xor U12375 (N_12375,N_8583,N_7205);
nand U12376 (N_12376,N_6872,N_8369);
and U12377 (N_12377,N_8653,N_6347);
or U12378 (N_12378,N_6459,N_8531);
and U12379 (N_12379,N_7680,N_6713);
or U12380 (N_12380,N_9250,N_7337);
xor U12381 (N_12381,N_9240,N_8329);
xor U12382 (N_12382,N_7250,N_6788);
or U12383 (N_12383,N_7315,N_7111);
nor U12384 (N_12384,N_7066,N_6832);
xor U12385 (N_12385,N_7081,N_7941);
nand U12386 (N_12386,N_9068,N_7510);
or U12387 (N_12387,N_6372,N_7065);
and U12388 (N_12388,N_9130,N_8985);
nor U12389 (N_12389,N_6373,N_8532);
nand U12390 (N_12390,N_8545,N_8123);
and U12391 (N_12391,N_6737,N_7802);
and U12392 (N_12392,N_7504,N_7280);
or U12393 (N_12393,N_9193,N_8391);
nand U12394 (N_12394,N_7028,N_9018);
nand U12395 (N_12395,N_8496,N_7542);
nand U12396 (N_12396,N_7581,N_6326);
nand U12397 (N_12397,N_6576,N_7017);
or U12398 (N_12398,N_8126,N_8046);
xor U12399 (N_12399,N_8836,N_9362);
or U12400 (N_12400,N_6645,N_8841);
or U12401 (N_12401,N_8328,N_8451);
and U12402 (N_12402,N_9178,N_6362);
nand U12403 (N_12403,N_8040,N_6866);
nor U12404 (N_12404,N_7887,N_9178);
xnor U12405 (N_12405,N_6523,N_7062);
nor U12406 (N_12406,N_9036,N_8314);
or U12407 (N_12407,N_7389,N_8871);
nor U12408 (N_12408,N_8786,N_6293);
nor U12409 (N_12409,N_7918,N_7716);
or U12410 (N_12410,N_7950,N_6718);
or U12411 (N_12411,N_9260,N_8420);
nor U12412 (N_12412,N_9002,N_9166);
and U12413 (N_12413,N_6625,N_7866);
and U12414 (N_12414,N_8429,N_7214);
or U12415 (N_12415,N_7055,N_7427);
nand U12416 (N_12416,N_7330,N_8869);
and U12417 (N_12417,N_8154,N_6416);
or U12418 (N_12418,N_8046,N_7015);
nor U12419 (N_12419,N_8213,N_7250);
xor U12420 (N_12420,N_7236,N_6537);
xnor U12421 (N_12421,N_7570,N_8422);
or U12422 (N_12422,N_6879,N_9017);
or U12423 (N_12423,N_6369,N_6528);
and U12424 (N_12424,N_7984,N_7584);
nand U12425 (N_12425,N_6688,N_6951);
or U12426 (N_12426,N_7732,N_8869);
xnor U12427 (N_12427,N_8301,N_8704);
or U12428 (N_12428,N_7138,N_7498);
or U12429 (N_12429,N_9033,N_8774);
and U12430 (N_12430,N_6476,N_7299);
nor U12431 (N_12431,N_6374,N_9242);
xnor U12432 (N_12432,N_6282,N_9236);
and U12433 (N_12433,N_8523,N_6505);
nand U12434 (N_12434,N_7142,N_6831);
nand U12435 (N_12435,N_9110,N_7271);
nor U12436 (N_12436,N_6721,N_6487);
and U12437 (N_12437,N_9325,N_6320);
nor U12438 (N_12438,N_8919,N_8046);
nor U12439 (N_12439,N_8842,N_9330);
nor U12440 (N_12440,N_8531,N_8711);
nor U12441 (N_12441,N_9021,N_8970);
or U12442 (N_12442,N_7704,N_7148);
and U12443 (N_12443,N_8177,N_8784);
xnor U12444 (N_12444,N_6397,N_7646);
nand U12445 (N_12445,N_8877,N_8915);
nor U12446 (N_12446,N_8311,N_7711);
nand U12447 (N_12447,N_7529,N_7426);
or U12448 (N_12448,N_7480,N_8274);
and U12449 (N_12449,N_8567,N_9037);
nand U12450 (N_12450,N_7816,N_6768);
or U12451 (N_12451,N_7131,N_7081);
or U12452 (N_12452,N_8484,N_8754);
nand U12453 (N_12453,N_7824,N_8245);
nor U12454 (N_12454,N_7967,N_9102);
or U12455 (N_12455,N_8083,N_8557);
nand U12456 (N_12456,N_6382,N_8491);
or U12457 (N_12457,N_8706,N_8813);
or U12458 (N_12458,N_9212,N_9036);
nor U12459 (N_12459,N_6987,N_9146);
xor U12460 (N_12460,N_8735,N_9063);
nor U12461 (N_12461,N_7781,N_8843);
nand U12462 (N_12462,N_7113,N_6654);
nand U12463 (N_12463,N_7400,N_7085);
xnor U12464 (N_12464,N_6730,N_6883);
xnor U12465 (N_12465,N_8297,N_7145);
nand U12466 (N_12466,N_9001,N_7838);
xor U12467 (N_12467,N_8477,N_7754);
xnor U12468 (N_12468,N_8213,N_8754);
and U12469 (N_12469,N_7167,N_8508);
nor U12470 (N_12470,N_6623,N_8522);
and U12471 (N_12471,N_7992,N_8542);
nor U12472 (N_12472,N_8728,N_6276);
nor U12473 (N_12473,N_7340,N_7299);
and U12474 (N_12474,N_9083,N_6941);
nor U12475 (N_12475,N_8131,N_8598);
nand U12476 (N_12476,N_7986,N_6986);
xnor U12477 (N_12477,N_8210,N_7519);
nor U12478 (N_12478,N_6418,N_6776);
or U12479 (N_12479,N_8910,N_7047);
xnor U12480 (N_12480,N_6437,N_6467);
xor U12481 (N_12481,N_8372,N_8101);
xnor U12482 (N_12482,N_8423,N_6254);
xor U12483 (N_12483,N_8806,N_9297);
nor U12484 (N_12484,N_8421,N_8115);
xor U12485 (N_12485,N_8963,N_8115);
xor U12486 (N_12486,N_8333,N_6853);
nand U12487 (N_12487,N_8153,N_6430);
nor U12488 (N_12488,N_8661,N_7832);
xor U12489 (N_12489,N_8374,N_6493);
nand U12490 (N_12490,N_7555,N_6491);
nor U12491 (N_12491,N_8414,N_6402);
nand U12492 (N_12492,N_8470,N_8731);
xor U12493 (N_12493,N_6472,N_8982);
xnor U12494 (N_12494,N_7957,N_6905);
nor U12495 (N_12495,N_7143,N_6843);
and U12496 (N_12496,N_8457,N_8319);
xor U12497 (N_12497,N_7984,N_6312);
nand U12498 (N_12498,N_9318,N_7731);
and U12499 (N_12499,N_6573,N_7696);
and U12500 (N_12500,N_10682,N_10166);
nor U12501 (N_12501,N_11533,N_10948);
nand U12502 (N_12502,N_11904,N_10904);
or U12503 (N_12503,N_10847,N_12341);
nand U12504 (N_12504,N_9806,N_12346);
nand U12505 (N_12505,N_10506,N_9997);
and U12506 (N_12506,N_10479,N_10561);
or U12507 (N_12507,N_9897,N_12151);
and U12508 (N_12508,N_11009,N_11166);
nand U12509 (N_12509,N_9537,N_9440);
xnor U12510 (N_12510,N_11013,N_10358);
nand U12511 (N_12511,N_11513,N_12278);
nor U12512 (N_12512,N_9453,N_11095);
xor U12513 (N_12513,N_9596,N_11562);
nor U12514 (N_12514,N_11132,N_10516);
nor U12515 (N_12515,N_10229,N_9906);
nand U12516 (N_12516,N_10216,N_9526);
or U12517 (N_12517,N_12444,N_11658);
and U12518 (N_12518,N_11207,N_12314);
and U12519 (N_12519,N_12113,N_10626);
nor U12520 (N_12520,N_11493,N_11942);
xnor U12521 (N_12521,N_9552,N_12211);
xnor U12522 (N_12522,N_10616,N_10518);
nand U12523 (N_12523,N_12179,N_11148);
nand U12524 (N_12524,N_11229,N_12060);
and U12525 (N_12525,N_10504,N_11289);
and U12526 (N_12526,N_10599,N_10890);
xor U12527 (N_12527,N_11872,N_10167);
nor U12528 (N_12528,N_9990,N_11469);
nor U12529 (N_12529,N_9489,N_11483);
or U12530 (N_12530,N_9564,N_11999);
and U12531 (N_12531,N_12072,N_11110);
xor U12532 (N_12532,N_11609,N_10064);
nor U12533 (N_12533,N_11263,N_11097);
and U12534 (N_12534,N_11695,N_10586);
or U12535 (N_12535,N_9782,N_10238);
or U12536 (N_12536,N_11932,N_11138);
and U12537 (N_12537,N_9527,N_11425);
nor U12538 (N_12538,N_11142,N_11621);
and U12539 (N_12539,N_11988,N_11901);
nor U12540 (N_12540,N_9391,N_12339);
nand U12541 (N_12541,N_10542,N_11434);
nor U12542 (N_12542,N_11671,N_9483);
nor U12543 (N_12543,N_11508,N_10022);
xor U12544 (N_12544,N_11921,N_11010);
nand U12545 (N_12545,N_11213,N_12200);
nor U12546 (N_12546,N_10783,N_11446);
xnor U12547 (N_12547,N_9447,N_11729);
or U12548 (N_12548,N_11801,N_10720);
or U12549 (N_12549,N_12329,N_11778);
nor U12550 (N_12550,N_12269,N_11666);
xor U12551 (N_12551,N_9765,N_10149);
nand U12552 (N_12552,N_9849,N_11819);
nand U12553 (N_12553,N_12224,N_12401);
and U12554 (N_12554,N_9571,N_12023);
nor U12555 (N_12555,N_10255,N_12057);
or U12556 (N_12556,N_11254,N_10099);
nand U12557 (N_12557,N_9503,N_12459);
xor U12558 (N_12558,N_10631,N_10851);
nor U12559 (N_12559,N_12364,N_10295);
nor U12560 (N_12560,N_10877,N_9620);
or U12561 (N_12561,N_12216,N_9589);
or U12562 (N_12562,N_9567,N_12294);
nand U12563 (N_12563,N_11236,N_12220);
and U12564 (N_12564,N_11029,N_12315);
and U12565 (N_12565,N_10517,N_12494);
xor U12566 (N_12566,N_11141,N_11812);
or U12567 (N_12567,N_12458,N_10269);
or U12568 (N_12568,N_9962,N_11720);
and U12569 (N_12569,N_10939,N_12239);
and U12570 (N_12570,N_11985,N_11136);
nand U12571 (N_12571,N_12000,N_9455);
xnor U12572 (N_12572,N_12487,N_12370);
xor U12573 (N_12573,N_10246,N_10932);
or U12574 (N_12574,N_10310,N_12373);
or U12575 (N_12575,N_10670,N_10540);
or U12576 (N_12576,N_11690,N_10034);
and U12577 (N_12577,N_10854,N_10287);
or U12578 (N_12578,N_9928,N_11913);
and U12579 (N_12579,N_11147,N_11731);
and U12580 (N_12580,N_10133,N_12282);
xor U12581 (N_12581,N_11847,N_10672);
nand U12582 (N_12582,N_10780,N_11159);
and U12583 (N_12583,N_9973,N_11541);
nor U12584 (N_12584,N_12044,N_11089);
xnor U12585 (N_12585,N_11435,N_12413);
nand U12586 (N_12586,N_11899,N_9711);
nor U12587 (N_12587,N_12146,N_11455);
and U12588 (N_12588,N_10487,N_12311);
or U12589 (N_12589,N_9947,N_11206);
nand U12590 (N_12590,N_12367,N_11874);
or U12591 (N_12591,N_10334,N_11252);
and U12592 (N_12592,N_10837,N_11046);
nor U12593 (N_12593,N_12340,N_11968);
and U12594 (N_12594,N_9777,N_10488);
and U12595 (N_12595,N_12188,N_9511);
nand U12596 (N_12596,N_10136,N_12051);
nor U12597 (N_12597,N_11885,N_12041);
or U12598 (N_12598,N_11960,N_9734);
nor U12599 (N_12599,N_12244,N_10966);
xor U12600 (N_12600,N_9380,N_9456);
nor U12601 (N_12601,N_10318,N_12495);
or U12602 (N_12602,N_10155,N_10951);
and U12603 (N_12603,N_11194,N_9794);
nand U12604 (N_12604,N_11087,N_11193);
and U12605 (N_12605,N_10585,N_11426);
nand U12606 (N_12606,N_9866,N_9384);
nand U12607 (N_12607,N_11864,N_10933);
nand U12608 (N_12608,N_10129,N_11567);
nor U12609 (N_12609,N_10570,N_9914);
and U12610 (N_12610,N_11754,N_11056);
or U12611 (N_12611,N_12331,N_11271);
and U12612 (N_12612,N_9550,N_9429);
or U12613 (N_12613,N_10926,N_11100);
nand U12614 (N_12614,N_10914,N_10285);
nand U12615 (N_12615,N_11675,N_11176);
xor U12616 (N_12616,N_11982,N_12391);
nor U12617 (N_12617,N_12018,N_10895);
nand U12618 (N_12618,N_10581,N_11001);
and U12619 (N_12619,N_10541,N_11413);
nor U12620 (N_12620,N_12074,N_10613);
or U12621 (N_12621,N_9484,N_11634);
and U12622 (N_12622,N_9877,N_9898);
nor U12623 (N_12623,N_10326,N_9624);
nand U12624 (N_12624,N_9414,N_9814);
or U12625 (N_12625,N_10913,N_12428);
nand U12626 (N_12626,N_9604,N_10312);
nand U12627 (N_12627,N_9381,N_12131);
nor U12628 (N_12628,N_11727,N_10148);
nand U12629 (N_12629,N_12075,N_10249);
nor U12630 (N_12630,N_10401,N_11412);
nor U12631 (N_12631,N_10111,N_12109);
xnor U12632 (N_12632,N_10537,N_9843);
nand U12633 (N_12633,N_9802,N_10856);
nor U12634 (N_12634,N_9671,N_12248);
or U12635 (N_12635,N_9530,N_11613);
or U12636 (N_12636,N_10708,N_9965);
and U12637 (N_12637,N_12300,N_9666);
or U12638 (N_12638,N_12205,N_10547);
or U12639 (N_12639,N_12240,N_11118);
xnor U12640 (N_12640,N_11733,N_10562);
nor U12641 (N_12641,N_11403,N_9938);
or U12642 (N_12642,N_9387,N_11368);
xor U12643 (N_12643,N_10676,N_9570);
nor U12644 (N_12644,N_9848,N_10811);
nor U12645 (N_12645,N_11633,N_10972);
xor U12646 (N_12646,N_11339,N_12307);
or U12647 (N_12647,N_11386,N_11930);
or U12648 (N_12648,N_11694,N_9967);
xor U12649 (N_12649,N_11811,N_10885);
and U12650 (N_12650,N_11753,N_11381);
xor U12651 (N_12651,N_10481,N_11879);
xnor U12652 (N_12652,N_10241,N_9678);
and U12653 (N_12653,N_9916,N_10432);
nand U12654 (N_12654,N_9515,N_10798);
or U12655 (N_12655,N_11762,N_10795);
xor U12656 (N_12656,N_10378,N_11162);
nand U12657 (N_12657,N_10224,N_10715);
xnor U12658 (N_12658,N_11449,N_9879);
nor U12659 (N_12659,N_9749,N_11787);
or U12660 (N_12660,N_10359,N_10299);
nor U12661 (N_12661,N_11121,N_10640);
nor U12662 (N_12662,N_10164,N_9619);
or U12663 (N_12663,N_10649,N_10499);
nor U12664 (N_12664,N_10557,N_11342);
nand U12665 (N_12665,N_10362,N_11517);
and U12666 (N_12666,N_9707,N_10991);
nand U12667 (N_12667,N_11591,N_9547);
nand U12668 (N_12668,N_10744,N_9392);
nand U12669 (N_12669,N_10686,N_10364);
nor U12670 (N_12670,N_12005,N_10677);
nor U12671 (N_12671,N_10835,N_12422);
nor U12672 (N_12672,N_11718,N_11155);
nor U12673 (N_12673,N_9759,N_9867);
nand U12674 (N_12674,N_11126,N_9560);
xnor U12675 (N_12675,N_10793,N_11400);
or U12676 (N_12676,N_11250,N_12204);
or U12677 (N_12677,N_9412,N_9838);
and U12678 (N_12678,N_11068,N_11700);
nand U12679 (N_12679,N_10794,N_11572);
or U12680 (N_12680,N_10028,N_9776);
or U12681 (N_12681,N_11222,N_10577);
xnor U12682 (N_12682,N_10871,N_10098);
or U12683 (N_12683,N_12147,N_9493);
nand U12684 (N_12684,N_10371,N_9837);
or U12685 (N_12685,N_9651,N_11824);
nand U12686 (N_12686,N_10905,N_12283);
nand U12687 (N_12687,N_11215,N_10580);
nand U12688 (N_12688,N_11057,N_10700);
and U12689 (N_12689,N_11320,N_10220);
nand U12690 (N_12690,N_10694,N_9491);
and U12691 (N_12691,N_10170,N_11767);
xnor U12692 (N_12692,N_12049,N_11333);
nand U12693 (N_12693,N_10668,N_9390);
nor U12694 (N_12694,N_12402,N_10159);
and U12695 (N_12695,N_9949,N_9839);
nand U12696 (N_12696,N_10648,N_10600);
and U12697 (N_12697,N_11829,N_11061);
xnor U12698 (N_12698,N_10699,N_9855);
and U12699 (N_12699,N_9538,N_11372);
nand U12700 (N_12700,N_11310,N_9730);
nand U12701 (N_12701,N_10426,N_11177);
nor U12702 (N_12702,N_12484,N_11346);
nand U12703 (N_12703,N_11487,N_11067);
and U12704 (N_12704,N_11407,N_9846);
xor U12705 (N_12705,N_10734,N_12295);
xnor U12706 (N_12706,N_10495,N_11924);
and U12707 (N_12707,N_12380,N_9506);
and U12708 (N_12708,N_11771,N_10707);
nand U12709 (N_12709,N_12419,N_11563);
nand U12710 (N_12710,N_11037,N_12008);
xnor U12711 (N_12711,N_10883,N_10763);
nand U12712 (N_12712,N_9864,N_9542);
or U12713 (N_12713,N_10662,N_9791);
nor U12714 (N_12714,N_11915,N_10360);
nor U12715 (N_12715,N_12090,N_12384);
nand U12716 (N_12716,N_12214,N_10297);
or U12717 (N_12717,N_11270,N_11117);
nand U12718 (N_12718,N_12454,N_11374);
nor U12719 (N_12719,N_12160,N_9512);
nor U12720 (N_12720,N_9808,N_12359);
xor U12721 (N_12721,N_9932,N_10770);
nand U12722 (N_12722,N_9409,N_11676);
nand U12723 (N_12723,N_9544,N_9912);
nand U12724 (N_12724,N_11855,N_9425);
and U12725 (N_12725,N_10058,N_9675);
and U12726 (N_12726,N_11708,N_11882);
and U12727 (N_12727,N_9850,N_10532);
and U12728 (N_12728,N_12336,N_12446);
and U12729 (N_12729,N_12030,N_12395);
and U12730 (N_12730,N_9861,N_11317);
or U12731 (N_12731,N_11581,N_9813);
or U12732 (N_12732,N_11000,N_12376);
nand U12733 (N_12733,N_10912,N_12353);
nand U12734 (N_12734,N_9685,N_12493);
or U12735 (N_12735,N_10717,N_11789);
nand U12736 (N_12736,N_11728,N_11408);
nand U12737 (N_12737,N_12114,N_10633);
or U12738 (N_12738,N_9658,N_11402);
and U12739 (N_12739,N_9719,N_11935);
nor U12740 (N_12740,N_9972,N_10251);
nand U12741 (N_12741,N_11308,N_11463);
xnor U12742 (N_12742,N_10531,N_10329);
nor U12743 (N_12743,N_10317,N_11981);
nand U12744 (N_12744,N_9774,N_9466);
and U12745 (N_12745,N_11496,N_10878);
nor U12746 (N_12746,N_9878,N_10974);
nor U12747 (N_12747,N_9653,N_9956);
or U12748 (N_12748,N_10419,N_10582);
and U12749 (N_12749,N_11826,N_10845);
nand U12750 (N_12750,N_9643,N_12327);
and U12751 (N_12751,N_10211,N_9461);
nor U12752 (N_12752,N_9605,N_11448);
and U12753 (N_12753,N_10342,N_11040);
xor U12754 (N_12754,N_11940,N_9534);
and U12755 (N_12755,N_9918,N_9609);
xor U12756 (N_12756,N_9767,N_10529);
and U12757 (N_12757,N_11098,N_9545);
nand U12758 (N_12758,N_9395,N_10181);
nand U12759 (N_12759,N_11373,N_10874);
nor U12760 (N_12760,N_10592,N_10415);
nand U12761 (N_12761,N_12056,N_10869);
and U12762 (N_12762,N_11612,N_12496);
or U12763 (N_12763,N_11546,N_11741);
or U12764 (N_12764,N_11625,N_10923);
nand U12765 (N_12765,N_12318,N_9923);
xor U12766 (N_12766,N_10969,N_11258);
nor U12767 (N_12767,N_10071,N_10889);
and U12768 (N_12768,N_12426,N_11835);
or U12769 (N_12769,N_9939,N_12238);
nand U12770 (N_12770,N_10896,N_10387);
nand U12771 (N_12771,N_11417,N_9688);
nor U12772 (N_12772,N_11843,N_10400);
nor U12773 (N_12773,N_9684,N_12138);
and U12774 (N_12774,N_10458,N_11189);
or U12775 (N_12775,N_10897,N_12048);
nand U12776 (N_12776,N_10916,N_9479);
and U12777 (N_12777,N_12261,N_11848);
xnor U12778 (N_12778,N_9950,N_10283);
or U12779 (N_12779,N_9845,N_10799);
nor U12780 (N_12780,N_10866,N_10920);
xor U12781 (N_12781,N_11149,N_11890);
nor U12782 (N_12782,N_9665,N_11547);
nor U12783 (N_12783,N_9668,N_12483);
nor U12784 (N_12784,N_10293,N_9536);
nor U12785 (N_12785,N_10349,N_11041);
xnor U12786 (N_12786,N_11534,N_11655);
xor U12787 (N_12787,N_12045,N_9809);
nor U12788 (N_12788,N_9410,N_11451);
or U12789 (N_12789,N_9873,N_10921);
xor U12790 (N_12790,N_10803,N_11322);
nor U12791 (N_12791,N_9736,N_10703);
or U12792 (N_12792,N_11703,N_9630);
xor U12793 (N_12793,N_12177,N_10177);
nand U12794 (N_12794,N_10683,N_11929);
and U12795 (N_12795,N_9903,N_10842);
or U12796 (N_12796,N_10138,N_10453);
and U12797 (N_12797,N_11775,N_9513);
or U12798 (N_12798,N_9880,N_12040);
xor U12799 (N_12799,N_10990,N_12301);
nor U12800 (N_12800,N_11792,N_9687);
xor U12801 (N_12801,N_9573,N_12482);
nor U12802 (N_12802,N_11321,N_10705);
or U12803 (N_12803,N_12118,N_10375);
nor U12804 (N_12804,N_12396,N_10952);
and U12805 (N_12805,N_9424,N_12172);
and U12806 (N_12806,N_10369,N_9746);
xnor U12807 (N_12807,N_11522,N_12488);
xnor U12808 (N_12808,N_11641,N_11084);
xnor U12809 (N_12809,N_9647,N_11382);
nand U12810 (N_12810,N_10829,N_11687);
and U12811 (N_12811,N_12234,N_10637);
or U12812 (N_12812,N_11277,N_9648);
or U12813 (N_12813,N_10500,N_12328);
and U12814 (N_12814,N_10962,N_11376);
nand U12815 (N_12815,N_11759,N_10353);
nor U12816 (N_12816,N_11123,N_11026);
or U12817 (N_12817,N_11130,N_11049);
xnor U12818 (N_12818,N_12129,N_11114);
nor U12819 (N_12819,N_11033,N_12195);
and U12820 (N_12820,N_10596,N_11477);
nor U12821 (N_12821,N_10989,N_10088);
and U12822 (N_12822,N_10043,N_12120);
and U12823 (N_12823,N_11167,N_11273);
xor U12824 (N_12824,N_12297,N_12362);
nand U12825 (N_12825,N_11833,N_11268);
xnor U12826 (N_12826,N_11397,N_10525);
nor U12827 (N_12827,N_11598,N_10194);
nor U12828 (N_12828,N_11889,N_9403);
and U12829 (N_12829,N_11256,N_11652);
nor U12830 (N_12830,N_9936,N_9557);
and U12831 (N_12831,N_10828,N_10523);
xnor U12832 (N_12832,N_10711,N_9416);
and U12833 (N_12833,N_10258,N_11616);
nand U12834 (N_12834,N_11008,N_12447);
xor U12835 (N_12835,N_10519,N_11844);
and U12836 (N_12836,N_9881,N_10443);
nand U12837 (N_12837,N_9869,N_11638);
xnor U12838 (N_12838,N_10591,N_11636);
xnor U12839 (N_12839,N_10652,N_11518);
or U12840 (N_12840,N_9454,N_10186);
nand U12841 (N_12841,N_10767,N_11596);
xnor U12842 (N_12842,N_10406,N_10049);
nand U12843 (N_12843,N_10199,N_10328);
nor U12844 (N_12844,N_12187,N_12343);
xor U12845 (N_12845,N_12157,N_9716);
xor U12846 (N_12846,N_11818,N_9434);
nand U12847 (N_12847,N_11594,N_11583);
nor U12848 (N_12848,N_9631,N_10381);
nor U12849 (N_12849,N_12445,N_11232);
or U12850 (N_12850,N_11312,N_9486);
or U12851 (N_12851,N_9768,N_10993);
nand U12852 (N_12852,N_11674,N_10663);
nor U12853 (N_12853,N_11362,N_12251);
xnor U12854 (N_12854,N_12386,N_10865);
nand U12855 (N_12855,N_9704,N_12105);
and U12856 (N_12856,N_9994,N_11357);
nor U12857 (N_12857,N_10018,N_12246);
or U12858 (N_12858,N_10644,N_11152);
or U12859 (N_12859,N_12174,N_11306);
nor U12860 (N_12860,N_11610,N_9642);
xnor U12861 (N_12861,N_10171,N_11521);
xnor U12862 (N_12862,N_11444,N_12249);
nor U12863 (N_12863,N_12361,N_11686);
or U12864 (N_12864,N_9607,N_10096);
xnor U12865 (N_12865,N_9785,N_10690);
nand U12866 (N_12866,N_10918,N_9520);
xnor U12867 (N_12867,N_11863,N_9964);
xor U12868 (N_12868,N_10910,N_10698);
and U12869 (N_12869,N_10056,N_10279);
or U12870 (N_12870,N_9502,N_11253);
or U12871 (N_12871,N_11973,N_10257);
nor U12872 (N_12872,N_12097,N_9613);
nand U12873 (N_12873,N_9929,N_10183);
nor U12874 (N_12874,N_10104,N_9610);
nand U12875 (N_12875,N_10787,N_11315);
nor U12876 (N_12876,N_10968,N_9789);
and U12877 (N_12877,N_9840,N_11479);
nor U12878 (N_12878,N_9800,N_9832);
and U12879 (N_12879,N_11351,N_10976);
or U12880 (N_12880,N_9927,N_10745);
and U12881 (N_12881,N_11230,N_10272);
and U12882 (N_12882,N_11223,N_12107);
nand U12883 (N_12883,N_10041,N_11458);
or U12884 (N_12884,N_12134,N_11717);
or U12885 (N_12885,N_9807,N_9663);
nand U12886 (N_12886,N_10740,N_11936);
or U12887 (N_12887,N_11143,N_10389);
nor U12888 (N_12888,N_11044,N_12034);
nor U12889 (N_12889,N_9656,N_11119);
or U12890 (N_12890,N_9496,N_10669);
or U12891 (N_12891,N_9494,N_10901);
xnor U12892 (N_12892,N_11875,N_9485);
xor U12893 (N_12893,N_10758,N_9398);
nor U12894 (N_12894,N_10270,N_10908);
and U12895 (N_12895,N_9989,N_11466);
or U12896 (N_12896,N_12095,N_11489);
xnor U12897 (N_12897,N_10134,N_12203);
and U12898 (N_12898,N_9862,N_12207);
xor U12899 (N_12899,N_11345,N_11174);
nand U12900 (N_12900,N_11994,N_10309);
and U12901 (N_12901,N_10535,N_11643);
nor U12902 (N_12902,N_11943,N_11265);
or U12903 (N_12903,N_10737,N_10046);
xnor U12904 (N_12904,N_10298,N_9915);
xor U12905 (N_12905,N_10144,N_11313);
and U12906 (N_12906,N_11330,N_12433);
or U12907 (N_12907,N_11475,N_10373);
nor U12908 (N_12908,N_10943,N_10014);
and U12909 (N_12909,N_10641,N_12443);
xor U12910 (N_12910,N_9715,N_12465);
nor U12911 (N_12911,N_10583,N_10462);
xor U12912 (N_12912,N_10870,N_11172);
xor U12913 (N_12913,N_11359,N_12158);
and U12914 (N_12914,N_9554,N_10053);
nand U12915 (N_12915,N_11106,N_10555);
xor U12916 (N_12916,N_9692,N_9933);
or U12917 (N_12917,N_11760,N_11706);
and U12918 (N_12918,N_12022,N_11918);
nor U12919 (N_12919,N_12026,N_11030);
nor U12920 (N_12920,N_9854,N_9559);
xnor U12921 (N_12921,N_11269,N_10730);
nand U12922 (N_12922,N_10000,N_11623);
nand U12923 (N_12923,N_10286,N_11470);
or U12924 (N_12924,N_11977,N_11219);
nor U12925 (N_12925,N_11461,N_11881);
nor U12926 (N_12926,N_9468,N_11139);
nor U12927 (N_12927,N_11996,N_11076);
or U12928 (N_12928,N_10861,N_11845);
or U12929 (N_12929,N_11484,N_10634);
or U12930 (N_12930,N_10067,N_9993);
xnor U12931 (N_12931,N_11954,N_10944);
or U12932 (N_12932,N_11804,N_11646);
xor U12933 (N_12933,N_11335,N_11014);
and U12934 (N_12934,N_10755,N_9669);
or U12935 (N_12935,N_9522,N_11715);
xor U12936 (N_12936,N_10749,N_10628);
nand U12937 (N_12937,N_9652,N_11347);
and U12938 (N_12938,N_12007,N_10819);
or U12939 (N_12939,N_10760,N_9925);
nand U12940 (N_12940,N_11751,N_12012);
xnor U12941 (N_12941,N_12397,N_10185);
and U12942 (N_12942,N_11133,N_9644);
nand U12943 (N_12943,N_10496,N_12167);
xor U12944 (N_12944,N_10218,N_11737);
nor U12945 (N_12945,N_12135,N_11251);
nor U12946 (N_12946,N_10240,N_11669);
xor U12947 (N_12947,N_11334,N_12274);
nand U12948 (N_12948,N_11004,N_12043);
or U12949 (N_12949,N_10100,N_11202);
xnor U12950 (N_12950,N_10497,N_10556);
and U12951 (N_12951,N_9773,N_9885);
nand U12952 (N_12952,N_11048,N_11356);
or U12953 (N_12953,N_11301,N_11822);
nor U12954 (N_12954,N_10765,N_11916);
nand U12955 (N_12955,N_12451,N_10469);
xnor U12956 (N_12956,N_9408,N_10219);
and U12957 (N_12957,N_12276,N_12291);
and U12958 (N_12958,N_9578,N_11560);
and U12959 (N_12959,N_9421,N_10924);
or U12960 (N_12960,N_12096,N_10403);
xor U12961 (N_12961,N_11006,N_10174);
or U12962 (N_12962,N_12490,N_9805);
nor U12963 (N_12963,N_11525,N_12460);
xor U12964 (N_12964,N_12281,N_9830);
and U12965 (N_12965,N_10121,N_11590);
nand U12966 (N_12966,N_12178,N_10544);
xnor U12967 (N_12967,N_12102,N_11442);
and U12968 (N_12968,N_12025,N_11553);
and U12969 (N_12969,N_12310,N_12006);
xor U12970 (N_12970,N_10528,N_12024);
nor U12971 (N_12971,N_10746,N_10788);
or U12972 (N_12972,N_10137,N_12442);
and U12973 (N_12973,N_11965,N_11244);
or U12974 (N_12974,N_9476,N_12171);
nand U12975 (N_12975,N_12247,N_12093);
nand U12976 (N_12976,N_10815,N_11103);
or U12977 (N_12977,N_12308,N_9888);
nor U12978 (N_12978,N_11739,N_10612);
or U12979 (N_12979,N_10187,N_9533);
xnor U12980 (N_12980,N_12227,N_10033);
and U12981 (N_12981,N_11876,N_9397);
or U12982 (N_12982,N_10513,N_10435);
nor U12983 (N_12983,N_10135,N_12266);
nor U12984 (N_12984,N_12111,N_12132);
nand U12985 (N_12985,N_10475,N_11050);
and U12986 (N_12986,N_11503,N_10797);
and U12987 (N_12987,N_11548,N_12421);
nor U12988 (N_12988,N_12063,N_10474);
and U12989 (N_12989,N_10005,N_9612);
xnor U12990 (N_12990,N_12463,N_10550);
xnor U12991 (N_12991,N_10604,N_11938);
and U12992 (N_12992,N_11539,N_10434);
and U12993 (N_12993,N_9591,N_10017);
or U12994 (N_12994,N_10625,N_11724);
nand U12995 (N_12995,N_12130,N_10817);
xnor U12996 (N_12996,N_12152,N_11651);
nand U12997 (N_12997,N_10482,N_10691);
or U12998 (N_12998,N_10796,N_11235);
or U12999 (N_12999,N_11714,N_10304);
nor U13000 (N_13000,N_11624,N_11266);
nand U13001 (N_13001,N_10052,N_10998);
or U13002 (N_13002,N_11070,N_10665);
nand U13003 (N_13003,N_10491,N_11353);
xnor U13004 (N_13004,N_9811,N_11113);
nor U13005 (N_13005,N_11797,N_10446);
nor U13006 (N_13006,N_11107,N_12393);
xnor U13007 (N_13007,N_11239,N_11530);
or U13008 (N_13008,N_10769,N_9771);
nand U13009 (N_13009,N_10431,N_10684);
xnor U13010 (N_13010,N_11908,N_11264);
nor U13011 (N_13011,N_11919,N_11561);
and U13012 (N_13012,N_10554,N_11846);
or U13013 (N_13013,N_9420,N_11922);
xor U13014 (N_13014,N_9541,N_10200);
nand U13015 (N_13015,N_12252,N_12140);
and U13016 (N_13016,N_11214,N_10152);
xor U13017 (N_13017,N_9991,N_10671);
nand U13018 (N_13018,N_9875,N_10179);
xor U13019 (N_13019,N_11409,N_11319);
xor U13020 (N_13020,N_11111,N_11385);
nor U13021 (N_13021,N_11730,N_12080);
xor U13022 (N_13022,N_10456,N_10261);
nor U13023 (N_13023,N_11770,N_10473);
xnor U13024 (N_13024,N_10223,N_9543);
or U13025 (N_13025,N_11604,N_12498);
xnor U13026 (N_13026,N_12223,N_11538);
nor U13027 (N_13027,N_12312,N_10365);
nor U13028 (N_13028,N_11240,N_10574);
nor U13029 (N_13029,N_11071,N_9532);
nand U13030 (N_13030,N_11668,N_9735);
nor U13031 (N_13031,N_11657,N_11173);
xnor U13032 (N_13032,N_12110,N_11725);
and U13033 (N_13033,N_11810,N_9469);
or U13034 (N_13034,N_10726,N_12027);
or U13035 (N_13035,N_11197,N_10651);
or U13036 (N_13036,N_10996,N_11672);
nand U13037 (N_13037,N_11241,N_11839);
nand U13038 (N_13038,N_9695,N_11018);
nand U13039 (N_13039,N_10762,N_11744);
nor U13040 (N_13040,N_10485,N_12162);
or U13041 (N_13041,N_12144,N_12037);
or U13042 (N_13042,N_12321,N_9539);
xor U13043 (N_13043,N_10459,N_11888);
nor U13044 (N_13044,N_10810,N_11422);
nor U13045 (N_13045,N_10376,N_11157);
xor U13046 (N_13046,N_9863,N_10421);
or U13047 (N_13047,N_10316,N_12055);
xor U13048 (N_13048,N_10973,N_11894);
and U13049 (N_13049,N_9889,N_12356);
nor U13050 (N_13050,N_11761,N_12258);
xnor U13051 (N_13051,N_12084,N_11424);
nand U13052 (N_13052,N_10131,N_9480);
and U13053 (N_13053,N_9988,N_11688);
nand U13054 (N_13054,N_11506,N_10549);
nor U13055 (N_13055,N_11267,N_12383);
nand U13056 (N_13056,N_11275,N_11783);
and U13057 (N_13057,N_12337,N_9510);
nand U13058 (N_13058,N_10305,N_12485);
nand U13059 (N_13059,N_9957,N_12183);
xnor U13060 (N_13060,N_12382,N_11341);
and U13061 (N_13061,N_9518,N_9452);
or U13062 (N_13062,N_10109,N_11047);
nand U13063 (N_13063,N_9629,N_11987);
nor U13064 (N_13064,N_10050,N_11165);
nor U13065 (N_13065,N_12015,N_12330);
nand U13066 (N_13066,N_10278,N_10068);
nor U13067 (N_13067,N_12381,N_11116);
and U13068 (N_13068,N_12303,N_9579);
or U13069 (N_13069,N_10953,N_10922);
xnor U13070 (N_13070,N_11282,N_10277);
xor U13071 (N_13071,N_10428,N_10303);
and U13072 (N_13072,N_9601,N_11927);
and U13073 (N_13073,N_10059,N_11806);
nor U13074 (N_13074,N_11259,N_12020);
nor U13075 (N_13075,N_11016,N_9525);
nor U13076 (N_13076,N_12036,N_11027);
nor U13077 (N_13077,N_11827,N_11281);
or U13078 (N_13078,N_12032,N_11369);
xor U13079 (N_13079,N_11108,N_11573);
xnor U13080 (N_13080,N_11286,N_9951);
or U13081 (N_13081,N_11732,N_10985);
nand U13082 (N_13082,N_10569,N_11179);
nand U13083 (N_13083,N_10732,N_11870);
nor U13084 (N_13084,N_10863,N_12001);
nor U13085 (N_13085,N_10938,N_11970);
nand U13086 (N_13086,N_10775,N_10398);
xor U13087 (N_13087,N_10526,N_10397);
nor U13088 (N_13088,N_11343,N_11234);
nor U13089 (N_13089,N_11821,N_12115);
and U13090 (N_13090,N_10060,N_11631);
nand U13091 (N_13091,N_10029,N_11805);
and U13092 (N_13092,N_11294,N_9521);
nor U13093 (N_13093,N_10533,N_12455);
or U13094 (N_13094,N_11073,N_11278);
or U13095 (N_13095,N_11025,N_9761);
nand U13096 (N_13096,N_12375,N_9935);
and U13097 (N_13097,N_12125,N_12417);
xor U13098 (N_13098,N_9501,N_11944);
xor U13099 (N_13099,N_9592,N_11948);
xnor U13100 (N_13100,N_11665,N_10308);
and U13101 (N_13101,N_11360,N_9500);
nor U13102 (N_13102,N_11247,N_10761);
xnor U13103 (N_13103,N_10127,N_11431);
or U13104 (N_13104,N_12236,N_10221);
xor U13105 (N_13105,N_9531,N_10436);
xor U13106 (N_13106,N_10404,N_12450);
nor U13107 (N_13107,N_10178,N_11284);
and U13108 (N_13108,N_12159,N_10695);
xnor U13109 (N_13109,N_12322,N_11928);
nor U13110 (N_13110,N_11682,N_9529);
nor U13111 (N_13111,N_11420,N_11742);
and U13112 (N_13112,N_11091,N_10906);
nor U13113 (N_13113,N_9874,N_10716);
nand U13114 (N_13114,N_9729,N_10840);
nand U13115 (N_13115,N_11871,N_11492);
nand U13116 (N_13116,N_12379,N_11740);
nor U13117 (N_13117,N_10825,N_11632);
xor U13118 (N_13118,N_10675,N_9772);
and U13119 (N_13119,N_11907,N_9974);
nor U13120 (N_13120,N_9549,N_9676);
nand U13121 (N_13121,N_10667,N_9896);
nor U13122 (N_13122,N_10163,N_10975);
nor U13123 (N_13123,N_10915,N_11023);
nor U13124 (N_13124,N_9548,N_12441);
and U13125 (N_13125,N_10314,N_12182);
nor U13126 (N_13126,N_11681,N_12309);
nand U13127 (N_13127,N_12265,N_10407);
xnor U13128 (N_13128,N_11054,N_11860);
nand U13129 (N_13129,N_11834,N_9460);
nor U13130 (N_13130,N_10019,N_9718);
and U13131 (N_13131,N_11902,N_11072);
nor U13132 (N_13132,N_11305,N_10986);
xor U13133 (N_13133,N_12166,N_10422);
nand U13134 (N_13134,N_12121,N_10172);
or U13135 (N_13135,N_11683,N_9982);
nand U13136 (N_13136,N_11459,N_11710);
nor U13137 (N_13137,N_9645,N_12112);
xnor U13138 (N_13138,N_9999,N_10452);
and U13139 (N_13139,N_11823,N_11774);
xor U13140 (N_13140,N_11752,N_12264);
or U13141 (N_13141,N_10848,N_12042);
xnor U13142 (N_13142,N_12462,N_10011);
xnor U13143 (N_13143,N_10350,N_11637);
and U13144 (N_13144,N_11802,N_10981);
or U13145 (N_13145,N_11622,N_9427);
xnor U13146 (N_13146,N_10451,N_10250);
nand U13147 (N_13147,N_10467,N_11480);
nand U13148 (N_13148,N_10658,N_12409);
nand U13149 (N_13149,N_11858,N_10593);
nand U13150 (N_13150,N_11473,N_11237);
and U13151 (N_13151,N_10417,N_12335);
xnor U13152 (N_13152,N_10553,N_10374);
nor U13153 (N_13153,N_10493,N_10119);
xnor U13154 (N_13154,N_9985,N_11188);
or U13155 (N_13155,N_10444,N_10572);
nor U13156 (N_13156,N_12089,N_9975);
nor U13157 (N_13157,N_9900,N_11437);
and U13158 (N_13158,N_10191,N_10460);
nor U13159 (N_13159,N_12290,N_11595);
and U13160 (N_13160,N_10281,N_11605);
or U13161 (N_13161,N_11304,N_10026);
xnor U13162 (N_13162,N_12245,N_11125);
xor U13163 (N_13163,N_9740,N_11887);
nor U13164 (N_13164,N_9986,N_11800);
or U13165 (N_13165,N_11081,N_11905);
nand U13166 (N_13166,N_10151,N_10013);
nor U13167 (N_13167,N_10645,N_11628);
and U13168 (N_13168,N_12377,N_11660);
or U13169 (N_13169,N_11452,N_10900);
and U13170 (N_13170,N_10830,N_11036);
nand U13171 (N_13171,N_12344,N_9661);
nor U13172 (N_13172,N_11495,N_11791);
or U13173 (N_13173,N_11620,N_12087);
nand U13174 (N_13174,N_10855,N_9446);
xor U13175 (N_13175,N_10410,N_11296);
and U13176 (N_13176,N_10015,N_9732);
nand U13177 (N_13177,N_9742,N_12275);
and U13178 (N_13178,N_11516,N_10113);
or U13179 (N_13179,N_11884,N_11707);
nand U13180 (N_13180,N_12255,N_10370);
or U13181 (N_13181,N_11663,N_11895);
and U13182 (N_13182,N_12059,N_10887);
xnor U13183 (N_13183,N_10980,N_11586);
nor U13184 (N_13184,N_11363,N_12390);
or U13185 (N_13185,N_10692,N_12013);
and U13186 (N_13186,N_12101,N_10492);
nor U13187 (N_13187,N_10723,N_9611);
nor U13188 (N_13188,N_11716,N_9659);
xnor U13189 (N_13189,N_10074,N_12126);
nor U13190 (N_13190,N_10066,N_10805);
nor U13191 (N_13191,N_11365,N_11670);
xor U13192 (N_13192,N_11291,N_9959);
nand U13193 (N_13193,N_11565,N_12400);
xnor U13194 (N_13194,N_11187,N_10042);
nor U13195 (N_13195,N_10080,N_11993);
or U13196 (N_13196,N_11020,N_10917);
xor U13197 (N_13197,N_10610,N_12153);
or U13198 (N_13198,N_12163,N_9738);
or U13199 (N_13199,N_11276,N_11526);
and U13200 (N_13200,N_10853,N_10954);
nand U13201 (N_13201,N_11667,N_11648);
or U13202 (N_13202,N_10624,N_9708);
nand U13203 (N_13203,N_11227,N_10892);
nor U13204 (N_13204,N_11512,N_12123);
or U13205 (N_13205,N_11075,N_12260);
and U13206 (N_13206,N_12285,N_10153);
and U13207 (N_13207,N_11112,N_9917);
nor U13208 (N_13208,N_9475,N_10824);
or U13209 (N_13209,N_10831,N_10212);
and U13210 (N_13210,N_9741,N_11052);
nand U13211 (N_13211,N_9680,N_10266);
xor U13212 (N_13212,N_10841,N_9628);
and U13213 (N_13213,N_9382,N_10994);
nor U13214 (N_13214,N_12351,N_11105);
and U13215 (N_13215,N_12029,N_9868);
nand U13216 (N_13216,N_10490,N_12201);
nor U13217 (N_13217,N_9823,N_10731);
or U13218 (N_13218,N_12360,N_10789);
nand U13219 (N_13219,N_11523,N_11211);
nor U13220 (N_13220,N_9954,N_9835);
or U13221 (N_13221,N_10206,N_10468);
and U13222 (N_13222,N_11869,N_10320);
nand U13223 (N_13223,N_10253,N_12436);
and U13224 (N_13224,N_11969,N_12349);
and U13225 (N_13225,N_11205,N_11765);
and U13226 (N_13226,N_11185,N_11809);
nor U13227 (N_13227,N_9795,N_12127);
nand U13228 (N_13228,N_12438,N_11745);
and U13229 (N_13229,N_10367,N_10551);
nor U13230 (N_13230,N_10522,N_11959);
nand U13231 (N_13231,N_9509,N_9442);
or U13232 (N_13232,N_9396,N_10440);
xnor U13233 (N_13233,N_11140,N_10713);
and U13234 (N_13234,N_10725,N_11396);
or U13235 (N_13235,N_10175,N_9702);
and U13236 (N_13236,N_10085,N_9481);
nor U13237 (N_13237,N_9764,N_11427);
xor U13238 (N_13238,N_11853,N_12486);
and U13239 (N_13239,N_9717,N_10282);
or U13240 (N_13240,N_9516,N_10971);
xor U13241 (N_13241,N_11584,N_11974);
xnor U13242 (N_13242,N_12424,N_11963);
nand U13243 (N_13243,N_9576,N_11464);
nor U13244 (N_13244,N_10337,N_10202);
nand U13245 (N_13245,N_11747,N_11124);
nor U13246 (N_13246,N_11600,N_11005);
xnor U13247 (N_13247,N_11178,N_10233);
xor U13248 (N_13248,N_10498,N_10728);
nor U13249 (N_13249,N_10145,N_11536);
nand U13250 (N_13250,N_10030,N_11580);
or U13251 (N_13251,N_9842,N_9747);
nor U13252 (N_13252,N_10265,N_10198);
nor U13253 (N_13253,N_12180,N_10605);
and U13254 (N_13254,N_9422,N_11292);
nand U13255 (N_13255,N_12186,N_9448);
xor U13256 (N_13256,N_11896,N_11639);
xor U13257 (N_13257,N_10950,N_11171);
xor U13258 (N_13258,N_10630,N_12479);
and U13259 (N_13259,N_10324,N_9419);
and U13260 (N_13260,N_11364,N_10330);
xor U13261 (N_13261,N_11777,N_11478);
xor U13262 (N_13262,N_10666,N_10606);
xnor U13263 (N_13263,N_11062,N_11090);
xnor U13264 (N_13264,N_10899,N_10210);
xor U13265 (N_13265,N_12031,N_11257);
nand U13266 (N_13266,N_12173,N_12452);
nand U13267 (N_13267,N_10225,N_10168);
xnor U13268 (N_13268,N_11419,N_12423);
xnor U13269 (N_13269,N_10623,N_10092);
or U13270 (N_13270,N_9377,N_12213);
xnor U13271 (N_13271,N_9913,N_11704);
nand U13272 (N_13272,N_10785,N_11436);
nor U13273 (N_13273,N_9482,N_10442);
nor U13274 (N_13274,N_9890,N_9588);
xor U13275 (N_13275,N_11588,N_10274);
nor U13276 (N_13276,N_10372,N_9883);
xor U13277 (N_13277,N_10396,N_10832);
and U13278 (N_13278,N_12070,N_10609);
or U13279 (N_13279,N_12196,N_12448);
or U13280 (N_13280,N_11443,N_9540);
nand U13281 (N_13281,N_10445,N_10339);
or U13282 (N_13282,N_9664,N_11245);
and U13283 (N_13283,N_12439,N_12241);
nand U13284 (N_13284,N_12389,N_10259);
xor U13285 (N_13285,N_10879,N_11926);
nor U13286 (N_13286,N_9597,N_10608);
and U13287 (N_13287,N_10379,N_10047);
or U13288 (N_13288,N_10007,N_9723);
or U13289 (N_13289,N_9615,N_10930);
nor U13290 (N_13290,N_10987,N_10394);
nor U13291 (N_13291,N_9804,N_10927);
nand U13292 (N_13292,N_11693,N_11743);
or U13293 (N_13293,N_9546,N_11131);
nand U13294 (N_13294,N_10685,N_10196);
and U13295 (N_13295,N_11293,N_12194);
or U13296 (N_13296,N_10243,N_12100);
nand U13297 (N_13297,N_11209,N_10539);
or U13298 (N_13298,N_9443,N_10327);
and U13299 (N_13299,N_12306,N_11307);
xnor U13300 (N_13300,N_11158,N_11153);
nand U13301 (N_13301,N_11274,N_10486);
xnor U13302 (N_13302,N_12133,N_11196);
or U13303 (N_13303,N_10739,N_10276);
or U13304 (N_13304,N_10031,N_11080);
nor U13305 (N_13305,N_11279,N_10169);
and U13306 (N_13306,N_9649,N_11911);
or U13307 (N_13307,N_11995,N_11699);
nand U13308 (N_13308,N_10363,N_9998);
and U13309 (N_13309,N_11946,N_11979);
or U13310 (N_13310,N_9691,N_11183);
or U13311 (N_13311,N_11723,N_9733);
or U13312 (N_13312,N_9517,N_12304);
nand U13313 (N_13313,N_12067,N_12139);
and U13314 (N_13314,N_9886,N_11456);
or U13315 (N_13315,N_9763,N_12254);
nand U13316 (N_13316,N_11329,N_11311);
and U13317 (N_13317,N_10888,N_12432);
nand U13318 (N_13318,N_10480,N_10733);
or U13319 (N_13319,N_10721,N_11832);
or U13320 (N_13320,N_9902,N_12268);
and U13321 (N_13321,N_9786,N_9438);
nand U13322 (N_13322,N_10463,N_10418);
nor U13323 (N_13323,N_11722,N_11606);
nor U13324 (N_13324,N_10790,N_12288);
and U13325 (N_13325,N_9852,N_12038);
and U13326 (N_13326,N_11543,N_10507);
nand U13327 (N_13327,N_12481,N_12062);
and U13328 (N_13328,N_11482,N_10543);
xnor U13329 (N_13329,N_10108,N_10735);
and U13330 (N_13330,N_10348,N_10361);
xor U13331 (N_13331,N_11208,N_9432);
xnor U13332 (N_13332,N_9968,N_12394);
nor U13333 (N_13333,N_12033,N_11615);
nand U13334 (N_13334,N_11045,N_10383);
nor U13335 (N_13335,N_11028,N_11544);
nor U13336 (N_13336,N_11238,N_11297);
nor U13337 (N_13337,N_10627,N_9581);
nor U13338 (N_13338,N_10025,N_11144);
nand U13339 (N_13339,N_9921,N_11763);
nand U13340 (N_13340,N_10288,N_11465);
nor U13341 (N_13341,N_11430,N_10234);
nand U13342 (N_13342,N_10524,N_11577);
nand U13343 (N_13343,N_10380,N_12073);
nand U13344 (N_13344,N_12404,N_9977);
nand U13345 (N_13345,N_9725,N_9586);
xnor U13346 (N_13346,N_11410,N_11984);
or U13347 (N_13347,N_11991,N_9551);
and U13348 (N_13348,N_10838,N_11951);
or U13349 (N_13349,N_11868,N_12298);
nor U13350 (N_13350,N_10289,N_9504);
nand U13351 (N_13351,N_10118,N_11989);
xor U13352 (N_13352,N_9709,N_11680);
or U13353 (N_13353,N_10594,N_10439);
nand U13354 (N_13354,N_11937,N_11217);
nor U13355 (N_13355,N_10091,N_11619);
xor U13356 (N_13356,N_10806,N_10204);
or U13357 (N_13357,N_11735,N_11825);
xor U13358 (N_13358,N_9674,N_9981);
xor U13359 (N_13359,N_9758,N_9565);
nand U13360 (N_13360,N_10860,N_10368);
or U13361 (N_13361,N_11712,N_11514);
nand U13362 (N_13362,N_9599,N_10182);
nor U13363 (N_13363,N_11550,N_10027);
or U13364 (N_13364,N_11998,N_10940);
nor U13365 (N_13365,N_9721,N_11423);
and U13366 (N_13366,N_10142,N_11692);
and U13367 (N_13367,N_9820,N_9722);
nor U13368 (N_13368,N_11485,N_9608);
xnor U13369 (N_13369,N_11654,N_10301);
nand U13370 (N_13370,N_10294,N_11861);
nand U13371 (N_13371,N_10073,N_11405);
and U13372 (N_13372,N_10455,N_10928);
nand U13373 (N_13373,N_10809,N_10674);
xor U13374 (N_13374,N_11352,N_10751);
or U13375 (N_13375,N_10102,N_10345);
nand U13376 (N_13376,N_10438,N_11569);
nand U13377 (N_13377,N_11755,N_11099);
nor U13378 (N_13378,N_12313,N_11494);
and U13379 (N_13379,N_12491,N_9799);
nand U13380 (N_13380,N_9379,N_9473);
nand U13381 (N_13381,N_12324,N_9770);
and U13382 (N_13382,N_9757,N_10388);
and U13383 (N_13383,N_11170,N_10176);
nor U13384 (N_13384,N_12259,N_10814);
nand U13385 (N_13385,N_10489,N_10188);
xnor U13386 (N_13386,N_10464,N_10611);
or U13387 (N_13387,N_11490,N_10160);
and U13388 (N_13388,N_9693,N_10748);
xnor U13389 (N_13389,N_12145,N_10189);
nand U13390 (N_13390,N_9640,N_11137);
and U13391 (N_13391,N_9787,N_11758);
and U13392 (N_13392,N_10955,N_10642);
or U13393 (N_13393,N_10931,N_9478);
xor U13394 (N_13394,N_11182,N_11094);
nor U13395 (N_13395,N_10508,N_10323);
or U13396 (N_13396,N_10984,N_9946);
or U13397 (N_13397,N_10655,N_11085);
or U13398 (N_13398,N_10816,N_12467);
or U13399 (N_13399,N_11447,N_9884);
nor U13400 (N_13400,N_9574,N_11332);
or U13401 (N_13401,N_9829,N_10201);
xnor U13402 (N_13402,N_11324,N_9528);
nand U13403 (N_13403,N_11433,N_11127);
and U13404 (N_13404,N_9433,N_11380);
xnor U13405 (N_13405,N_11830,N_10821);
and U13406 (N_13406,N_12219,N_12017);
and U13407 (N_13407,N_11529,N_10872);
xor U13408 (N_13408,N_9562,N_12232);
nor U13409 (N_13409,N_12065,N_10140);
nand U13410 (N_13410,N_12430,N_11958);
nand U13411 (N_13411,N_10180,N_11034);
nand U13412 (N_13412,N_9617,N_9407);
nand U13413 (N_13413,N_10280,N_11817);
xnor U13414 (N_13414,N_12091,N_10222);
nor U13415 (N_13415,N_10184,N_11017);
or U13416 (N_13416,N_9922,N_10882);
nor U13417 (N_13417,N_12253,N_9969);
xor U13418 (N_13418,N_10083,N_9603);
and U13419 (N_13419,N_12098,N_10886);
or U13420 (N_13420,N_11328,N_10146);
xor U13421 (N_13421,N_12354,N_10264);
nand U13422 (N_13422,N_11186,N_11816);
nand U13423 (N_13423,N_9499,N_11705);
or U13424 (N_13424,N_12054,N_10722);
or U13425 (N_13425,N_12385,N_11201);
nor U13426 (N_13426,N_11210,N_11589);
xor U13427 (N_13427,N_12198,N_11807);
and U13428 (N_13428,N_10909,N_9828);
nor U13429 (N_13429,N_10450,N_9672);
nor U13430 (N_13430,N_9860,N_10567);
and U13431 (N_13431,N_9779,N_10433);
nand U13432 (N_13432,N_10313,N_12299);
xor U13433 (N_13433,N_12478,N_11857);
or U13434 (N_13434,N_10946,N_9706);
nand U13435 (N_13435,N_10273,N_11203);
nor U13436 (N_13436,N_12347,N_10141);
and U13437 (N_13437,N_10696,N_10800);
nand U13438 (N_13438,N_9474,N_11199);
nor U13439 (N_13439,N_10425,N_10538);
nor U13440 (N_13440,N_11285,N_10228);
and U13441 (N_13441,N_12237,N_11866);
nand U13442 (N_13442,N_11476,N_12415);
and U13443 (N_13443,N_11379,N_10964);
nand U13444 (N_13444,N_9689,N_11627);
or U13445 (N_13445,N_11401,N_9677);
nor U13446 (N_13446,N_11021,N_11820);
nand U13447 (N_13447,N_11039,N_11956);
nor U13448 (N_13448,N_9712,N_12357);
and U13449 (N_13449,N_11611,N_11618);
or U13450 (N_13450,N_9487,N_10941);
nand U13451 (N_13451,N_11910,N_10051);
nor U13452 (N_13452,N_11772,N_11997);
xnor U13453 (N_13453,N_12217,N_9681);
xor U13454 (N_13454,N_10601,N_11570);
nor U13455 (N_13455,N_10768,N_9386);
xor U13456 (N_13456,N_9464,N_10414);
nor U13457 (N_13457,N_11554,N_9934);
and U13458 (N_13458,N_10093,N_9955);
nand U13459 (N_13459,N_10678,N_12489);
nand U13460 (N_13460,N_12193,N_10090);
xnor U13461 (N_13461,N_12410,N_10239);
and U13462 (N_13462,N_9488,N_9492);
nor U13463 (N_13463,N_10045,N_11104);
nand U13464 (N_13464,N_12368,N_9497);
and U13465 (N_13465,N_10448,N_12185);
nand U13466 (N_13466,N_10568,N_12137);
xor U13467 (N_13467,N_10021,N_11702);
nor U13468 (N_13468,N_9892,N_9563);
xnor U13469 (N_13469,N_11053,N_9821);
and U13470 (N_13470,N_12372,N_11630);
xnor U13471 (N_13471,N_10902,N_9882);
nand U13472 (N_13472,N_10719,N_11659);
xor U13473 (N_13473,N_10441,N_10244);
nor U13474 (N_13474,N_9941,N_11371);
and U13475 (N_13475,N_10284,N_10827);
nor U13476 (N_13476,N_10530,N_9931);
xnor U13477 (N_13477,N_11395,N_12009);
or U13478 (N_13478,N_10689,N_9595);
and U13479 (N_13479,N_11537,N_12184);
nand U13480 (N_13480,N_10412,N_12010);
nor U13481 (N_13481,N_12420,N_10852);
or U13482 (N_13482,N_10503,N_9635);
xnor U13483 (N_13483,N_11290,N_10710);
nor U13484 (N_13484,N_10430,N_9701);
and U13485 (N_13485,N_12053,N_11865);
nor U13486 (N_13486,N_11642,N_9444);
and U13487 (N_13487,N_10843,N_12035);
or U13488 (N_13488,N_9944,N_12469);
and U13489 (N_13489,N_10578,N_9703);
nor U13490 (N_13490,N_12079,N_11077);
or U13491 (N_13491,N_11557,N_9602);
xnor U13492 (N_13492,N_11952,N_12270);
or U13493 (N_13493,N_11906,N_10661);
xnor U13494 (N_13494,N_10300,N_10907);
xnor U13495 (N_13495,N_10035,N_11007);
and U13496 (N_13496,N_11024,N_11325);
xor U13497 (N_13497,N_11603,N_11803);
nor U13498 (N_13498,N_9650,N_11909);
and U13499 (N_13499,N_11181,N_9780);
nor U13500 (N_13500,N_12019,N_12411);
nor U13501 (N_13501,N_9904,N_9841);
xor U13502 (N_13502,N_10036,N_9937);
or U13503 (N_13503,N_10548,N_9556);
xor U13504 (N_13504,N_9870,N_12243);
or U13505 (N_13505,N_11454,N_9660);
nand U13506 (N_13506,N_12345,N_9815);
xnor U13507 (N_13507,N_10271,N_10603);
nor U13508 (N_13508,N_12425,N_11318);
xor U13509 (N_13509,N_9788,N_10771);
or U13510 (N_13510,N_11387,N_10470);
and U13511 (N_13511,N_10709,N_9618);
and U13512 (N_13512,N_11813,N_11055);
xor U13513 (N_13513,N_11923,N_10935);
or U13514 (N_13514,N_10325,N_11486);
nor U13515 (N_13515,N_9945,N_12150);
nor U13516 (N_13516,N_11990,N_12003);
nor U13517 (N_13517,N_9930,N_11058);
nand U13518 (N_13518,N_10566,N_9926);
or U13519 (N_13519,N_12039,N_9430);
xor U13520 (N_13520,N_10701,N_12398);
nor U13521 (N_13521,N_11355,N_10743);
and U13522 (N_13522,N_10215,N_10629);
nor U13523 (N_13523,N_11218,N_9847);
or U13524 (N_13524,N_10729,N_10706);
nor U13525 (N_13525,N_10782,N_10089);
xor U13526 (N_13526,N_9519,N_10209);
xor U13527 (N_13527,N_11415,N_9524);
and U13528 (N_13528,N_10786,N_12412);
nor U13529 (N_13529,N_9459,N_11390);
nor U13530 (N_13530,N_12077,N_11491);
nand U13531 (N_13531,N_10128,N_10560);
nand U13532 (N_13532,N_10718,N_12333);
or U13533 (N_13533,N_10801,N_12088);
nor U13534 (N_13534,N_11184,N_9561);
or U13535 (N_13535,N_11168,N_9752);
and U13536 (N_13536,N_11344,N_9441);
nand U13537 (N_13537,N_11280,N_10413);
and U13538 (N_13538,N_11367,N_10402);
xnor U13539 (N_13539,N_11786,N_10589);
xnor U13540 (N_13540,N_10515,N_10411);
xor U13541 (N_13541,N_11391,N_11169);
nor U13542 (N_13542,N_10296,N_10192);
xnor U13543 (N_13543,N_10501,N_10366);
nor U13544 (N_13544,N_10679,N_10112);
nor U13545 (N_13545,N_12164,N_12284);
nor U13546 (N_13546,N_11361,N_11366);
xor U13547 (N_13547,N_11891,N_10023);
or U13548 (N_13548,N_9966,N_10822);
xnor U13549 (N_13549,N_11992,N_9436);
or U13550 (N_13550,N_10511,N_9983);
xor U13551 (N_13551,N_9639,N_10054);
and U13552 (N_13552,N_10621,N_9585);
xnor U13553 (N_13553,N_9696,N_11966);
xor U13554 (N_13554,N_10390,N_9389);
or U13555 (N_13555,N_11976,N_10833);
nand U13556 (N_13556,N_12128,N_11662);
nor U13557 (N_13557,N_10970,N_10254);
or U13558 (N_13558,N_12218,N_10126);
xor U13559 (N_13559,N_11326,N_11101);
or U13560 (N_13560,N_9445,N_12480);
xnor U13561 (N_13561,N_11945,N_12076);
nand U13562 (N_13562,N_10101,N_10237);
xor U13563 (N_13563,N_11673,N_10945);
or U13564 (N_13564,N_11593,N_9818);
nor U13565 (N_13565,N_11200,N_9810);
xnor U13566 (N_13566,N_11088,N_11527);
or U13567 (N_13567,N_10065,N_10750);
nand U13568 (N_13568,N_10903,N_10781);
xor U13569 (N_13569,N_9616,N_12464);
nand U13570 (N_13570,N_9853,N_11795);
nor U13571 (N_13571,N_10687,N_12403);
or U13572 (N_13572,N_9388,N_10999);
or U13573 (N_13573,N_11576,N_9958);
and U13574 (N_13574,N_9827,N_10764);
xnor U13575 (N_13575,N_12358,N_10106);
xnor U13576 (N_13576,N_11043,N_10607);
nor U13577 (N_13577,N_10105,N_10873);
or U13578 (N_13578,N_11331,N_11115);
and U13579 (N_13579,N_10868,N_11726);
nand U13580 (N_13580,N_9598,N_11790);
and U13581 (N_13581,N_11128,N_11011);
and U13582 (N_13582,N_9698,N_10346);
nor U13583 (N_13583,N_10116,N_11051);
and U13584 (N_13584,N_9580,N_11135);
nor U13585 (N_13585,N_11120,N_10846);
or U13586 (N_13586,N_11689,N_11592);
or U13587 (N_13587,N_12440,N_11416);
and U13588 (N_13588,N_11327,N_11348);
xor U13589 (N_13589,N_11782,N_12296);
nand U13590 (N_13590,N_12154,N_10039);
nor U13591 (N_13591,N_10997,N_10124);
and U13592 (N_13592,N_9727,N_10125);
and U13593 (N_13593,N_11134,N_10632);
xnor U13594 (N_13594,N_11949,N_11545);
or U13595 (N_13595,N_10614,N_9673);
nand U13596 (N_13596,N_10399,N_11468);
nor U13597 (N_13597,N_9670,N_11886);
nor U13598 (N_13598,N_9404,N_11784);
and U13599 (N_13599,N_9450,N_11501);
and U13600 (N_13600,N_11224,N_10357);
or U13601 (N_13601,N_9731,N_11019);
nand U13602 (N_13602,N_11261,N_9960);
xor U13603 (N_13603,N_12473,N_11933);
or U13604 (N_13604,N_10595,N_12142);
xnor U13605 (N_13605,N_9784,N_11532);
nand U13606 (N_13606,N_9402,N_11038);
and U13607 (N_13607,N_11204,N_10256);
nand U13608 (N_13608,N_10502,N_9793);
or U13609 (N_13609,N_11074,N_11260);
nor U13610 (N_13610,N_11287,N_12016);
nand U13611 (N_13611,N_11350,N_9411);
nor U13612 (N_13612,N_11650,N_9587);
nor U13613 (N_13613,N_10263,N_12206);
and U13614 (N_13614,N_10898,N_10157);
nor U13615 (N_13615,N_12471,N_10807);
nand U13616 (N_13616,N_12378,N_9783);
nand U13617 (N_13617,N_11851,N_10653);
xnor U13618 (N_13618,N_11925,N_11779);
nor U13619 (N_13619,N_11691,N_10117);
xor U13620 (N_13620,N_10232,N_11519);
or U13621 (N_13621,N_11877,N_11429);
xor U13622 (N_13622,N_11295,N_10063);
xnor U13623 (N_13623,N_11354,N_11102);
xor U13624 (N_13624,N_11849,N_10635);
xnor U13625 (N_13625,N_9699,N_11488);
or U13626 (N_13626,N_12064,N_11065);
nand U13627 (N_13627,N_11962,N_12271);
nand U13628 (N_13628,N_11957,N_10759);
xor U13629 (N_13629,N_11520,N_12169);
xor U13630 (N_13630,N_12338,N_10754);
or U13631 (N_13631,N_10527,N_12325);
xor U13632 (N_13632,N_9760,N_12267);
or U13633 (N_13633,N_11212,N_11507);
and U13634 (N_13634,N_11375,N_9905);
nor U13635 (N_13635,N_10245,N_10420);
or U13636 (N_13636,N_10636,N_12279);
nand U13637 (N_13637,N_10858,N_11559);
nand U13638 (N_13638,N_10075,N_12228);
xor U13639 (N_13639,N_11302,N_11129);
nor U13640 (N_13640,N_10355,N_10004);
nor U13641 (N_13641,N_10812,N_11228);
xor U13642 (N_13642,N_11582,N_10565);
nand U13643 (N_13643,N_9394,N_11815);
or U13644 (N_13644,N_9458,N_11323);
nor U13645 (N_13645,N_11035,N_9801);
nor U13646 (N_13646,N_12141,N_9457);
and U13647 (N_13647,N_11032,N_9714);
or U13648 (N_13648,N_10391,N_9498);
nand U13649 (N_13649,N_11500,N_10291);
nand U13650 (N_13650,N_11842,N_11063);
xnor U13651 (N_13651,N_10772,N_11836);
nand U13652 (N_13652,N_9753,N_12061);
or U13653 (N_13653,N_11551,N_11316);
or U13654 (N_13654,N_10536,N_10747);
nand U13655 (N_13655,N_10268,N_12472);
xnor U13656 (N_13656,N_9909,N_11384);
and U13657 (N_13657,N_12457,N_10429);
and U13658 (N_13658,N_11912,N_10963);
nand U13659 (N_13659,N_9385,N_10078);
nand U13660 (N_13660,N_10311,N_10978);
nor U13661 (N_13661,N_12014,N_10844);
nor U13662 (N_13662,N_10156,N_9984);
and U13663 (N_13663,N_10657,N_10290);
nand U13664 (N_13664,N_11164,N_10774);
or U13665 (N_13665,N_9523,N_9679);
or U13666 (N_13666,N_10752,N_11093);
and U13667 (N_13667,N_12071,N_9682);
or U13668 (N_13668,N_11216,N_10070);
xnor U13669 (N_13669,N_10107,N_10081);
or U13670 (N_13670,N_11656,N_9694);
and U13671 (N_13671,N_11756,N_9633);
xnor U13672 (N_13672,N_10510,N_10925);
nand U13673 (N_13673,N_11552,N_10576);
xor U13674 (N_13674,N_9490,N_12317);
nand U13675 (N_13675,N_10949,N_10395);
xnor U13676 (N_13676,N_12221,N_11878);
or U13677 (N_13677,N_11393,N_10802);
or U13678 (N_13678,N_12168,N_12170);
and U13679 (N_13679,N_10639,N_10808);
nor U13680 (N_13680,N_10333,N_10893);
or U13681 (N_13681,N_11854,N_11474);
or U13682 (N_13682,N_11579,N_10988);
nor U13683 (N_13683,N_10207,N_11558);
and U13684 (N_13684,N_11358,N_11950);
nor U13685 (N_13685,N_10659,N_11440);
or U13686 (N_13686,N_10009,N_9720);
nor U13687 (N_13687,N_10055,N_9816);
nand U13688 (N_13688,N_11644,N_10193);
or U13689 (N_13689,N_10688,N_10784);
and U13690 (N_13690,N_11394,N_9871);
nand U13691 (N_13691,N_10057,N_11498);
nor U13692 (N_13692,N_10983,N_9792);
nand U13693 (N_13693,N_11607,N_10563);
nor U13694 (N_13694,N_11082,N_11769);
nor U13695 (N_13695,N_10875,N_10103);
xnor U13696 (N_13696,N_12190,N_9558);
nor U13697 (N_13697,N_11064,N_12028);
and U13698 (N_13698,N_10876,N_11785);
and U13699 (N_13699,N_10130,N_9507);
nor U13700 (N_13700,N_9435,N_11457);
and U13701 (N_13701,N_12225,N_12058);
or U13702 (N_13702,N_11540,N_10584);
nand U13703 (N_13703,N_11971,N_11840);
nand U13704 (N_13704,N_11531,N_12435);
nand U13705 (N_13705,N_11411,N_11421);
and U13706 (N_13706,N_10638,N_11978);
or U13707 (N_13707,N_12094,N_10347);
xor U13708 (N_13708,N_12189,N_12222);
nand U13709 (N_13709,N_11768,N_10472);
nor U13710 (N_13710,N_11713,N_9575);
or U13711 (N_13711,N_10704,N_9907);
or U13712 (N_13712,N_10252,N_12407);
nand U13713 (N_13713,N_11220,N_12277);
nor U13714 (N_13714,N_10423,N_10162);
and U13715 (N_13715,N_12292,N_11776);
nor U13716 (N_13716,N_12319,N_9995);
nor U13717 (N_13717,N_11002,N_10937);
nor U13718 (N_13718,N_9876,N_11850);
nand U13719 (N_13719,N_11750,N_10849);
nor U13720 (N_13720,N_11059,N_9622);
or U13721 (N_13721,N_12021,N_9463);
xor U13722 (N_13722,N_11838,N_11629);
nor U13723 (N_13723,N_9751,N_9978);
and U13724 (N_13724,N_11060,N_11684);
nand U13725 (N_13725,N_11617,N_11719);
xnor U13726 (N_13726,N_10457,N_9683);
and U13727 (N_13727,N_10385,N_11575);
nor U13728 (N_13728,N_9423,N_9857);
or U13729 (N_13729,N_10427,N_10738);
nand U13730 (N_13730,N_11505,N_10319);
nor U13731 (N_13731,N_12499,N_9895);
nand U13732 (N_13732,N_10077,N_11568);
xnor U13733 (N_13733,N_11337,N_9971);
or U13734 (N_13734,N_9577,N_10120);
and U13735 (N_13735,N_9417,N_10934);
and U13736 (N_13736,N_10862,N_11298);
nand U13737 (N_13737,N_9901,N_10712);
nand U13738 (N_13738,N_11418,N_10062);
and U13739 (N_13739,N_12305,N_10929);
or U13740 (N_13740,N_10016,N_11649);
xnor U13741 (N_13741,N_10741,N_9553);
or U13742 (N_13742,N_10214,N_9439);
and U13743 (N_13743,N_9769,N_9375);
nor U13744 (N_13744,N_11814,N_9943);
or U13745 (N_13745,N_11299,N_9636);
or U13746 (N_13746,N_10344,N_12406);
xor U13747 (N_13747,N_11154,N_10115);
xor U13748 (N_13748,N_11574,N_12320);
nor U13749 (N_13749,N_10559,N_11249);
or U13750 (N_13750,N_12106,N_10405);
or U13751 (N_13751,N_10911,N_10356);
nand U13752 (N_13752,N_12492,N_12323);
nor U13753 (N_13753,N_9495,N_10477);
xor U13754 (N_13754,N_10037,N_11404);
and U13755 (N_13755,N_9910,N_9634);
or U13756 (N_13756,N_11749,N_11509);
or U13757 (N_13757,N_11180,N_9781);
xnor U13758 (N_13758,N_9614,N_9686);
nor U13759 (N_13759,N_11377,N_12453);
xor U13760 (N_13760,N_11504,N_9952);
xor U13761 (N_13761,N_11964,N_11564);
and U13762 (N_13762,N_10656,N_11192);
nor U13763 (N_13763,N_11499,N_11862);
nand U13764 (N_13764,N_12476,N_10024);
xor U13765 (N_13765,N_12399,N_11383);
nor U13766 (N_13766,N_12165,N_10857);
and U13767 (N_13767,N_12197,N_12355);
nand U13768 (N_13768,N_12233,N_9431);
nand U13769 (N_13769,N_10602,N_10505);
nand U13770 (N_13770,N_11897,N_12374);
nor U13771 (N_13771,N_11150,N_10960);
xnor U13772 (N_13772,N_11947,N_11428);
nor U13773 (N_13773,N_12143,N_10197);
xor U13774 (N_13774,N_12176,N_9465);
or U13775 (N_13775,N_11934,N_11190);
or U13776 (N_13776,N_11272,N_9851);
or U13777 (N_13777,N_10587,N_11920);
xnor U13778 (N_13778,N_10393,N_11764);
nor U13779 (N_13779,N_11079,N_10714);
nand U13780 (N_13780,N_11195,N_10132);
or U13781 (N_13781,N_10227,N_9401);
or U13782 (N_13782,N_10002,N_10377);
nor U13783 (N_13783,N_9426,N_9891);
nor U13784 (N_13784,N_10958,N_10236);
and U13785 (N_13785,N_9826,N_11983);
and U13786 (N_13786,N_12427,N_9724);
nand U13787 (N_13787,N_12348,N_11685);
and U13788 (N_13788,N_10048,N_9627);
xnor U13789 (N_13789,N_9654,N_10521);
and U13790 (N_13790,N_10514,N_9632);
xnor U13791 (N_13791,N_10465,N_12416);
and U13792 (N_13792,N_10248,N_11856);
nor U13793 (N_13793,N_10384,N_12280);
nor U13794 (N_13794,N_10742,N_11096);
nand U13795 (N_13795,N_10813,N_11939);
or U13796 (N_13796,N_12263,N_11602);
or U13797 (N_13797,N_9844,N_11151);
and U13798 (N_13798,N_12242,N_11794);
and U13799 (N_13799,N_10773,N_10087);
nand U13800 (N_13800,N_9775,N_10859);
or U13801 (N_13801,N_10020,N_10965);
nand U13802 (N_13802,N_10110,N_10340);
xnor U13803 (N_13803,N_10260,N_9790);
xnor U13804 (N_13804,N_11066,N_9467);
xnor U13805 (N_13805,N_11314,N_12199);
or U13806 (N_13806,N_10476,N_11696);
xnor U13807 (N_13807,N_10959,N_12155);
or U13808 (N_13808,N_10588,N_12108);
or U13809 (N_13809,N_11399,N_11635);
and U13810 (N_13810,N_11160,N_10006);
nand U13811 (N_13811,N_11467,N_12250);
nor U13812 (N_13812,N_10351,N_11163);
nand U13813 (N_13813,N_10512,N_10449);
or U13814 (N_13814,N_12082,N_10161);
nor U13815 (N_13815,N_11243,N_10977);
xor U13816 (N_13816,N_10804,N_10386);
nand U13817 (N_13817,N_12273,N_11083);
or U13818 (N_13818,N_10335,N_10697);
and U13819 (N_13819,N_9745,N_10466);
xor U13820 (N_13820,N_12117,N_11338);
nand U13821 (N_13821,N_9754,N_10217);
or U13822 (N_13822,N_11859,N_12136);
nand U13823 (N_13823,N_11462,N_11378);
nand U13824 (N_13824,N_11255,N_11773);
or U13825 (N_13825,N_10867,N_9728);
nand U13826 (N_13826,N_10995,N_10724);
nor U13827 (N_13827,N_9623,N_9940);
xnor U13828 (N_13828,N_10001,N_11757);
nor U13829 (N_13829,N_9378,N_11841);
nor U13830 (N_13830,N_10331,N_11161);
nand U13831 (N_13831,N_10979,N_12332);
nor U13832 (N_13832,N_9667,N_9566);
or U13833 (N_13833,N_10322,N_11225);
or U13834 (N_13834,N_9470,N_12004);
nor U13835 (N_13835,N_12104,N_12470);
nand U13836 (N_13836,N_9400,N_9762);
or U13837 (N_13837,N_12119,N_9697);
xnor U13838 (N_13838,N_12474,N_10673);
nand U13839 (N_13839,N_11578,N_10834);
and U13840 (N_13840,N_9590,N_9942);
xnor U13841 (N_13841,N_11042,N_11601);
or U13842 (N_13842,N_9963,N_10341);
and U13843 (N_13843,N_10509,N_10072);
and U13844 (N_13844,N_10352,N_9584);
xor U13845 (N_13845,N_10332,N_9700);
nor U13846 (N_13846,N_10660,N_12352);
and U13847 (N_13847,N_10424,N_10736);
xor U13848 (N_13848,N_12286,N_11453);
and U13849 (N_13849,N_9606,N_11900);
nand U13850 (N_13850,N_9568,N_9594);
and U13851 (N_13851,N_10681,N_11734);
nand U13852 (N_13852,N_10961,N_10230);
and U13853 (N_13853,N_9582,N_11221);
xor U13854 (N_13854,N_11701,N_9812);
and U13855 (N_13855,N_12363,N_10262);
nor U13856 (N_13856,N_9961,N_11524);
and U13857 (N_13857,N_12477,N_9413);
nand U13858 (N_13858,N_12468,N_11972);
nand U13859 (N_13859,N_11388,N_10494);
and U13860 (N_13860,N_11406,N_12408);
nand U13861 (N_13861,N_12293,N_10154);
xor U13862 (N_13862,N_9872,N_12212);
xor U13863 (N_13863,N_11914,N_10618);
nor U13864 (N_13864,N_9737,N_9535);
xnor U13865 (N_13865,N_11883,N_9798);
nor U13866 (N_13866,N_12092,N_10919);
nand U13867 (N_13867,N_10779,N_11799);
nor U13868 (N_13868,N_9858,N_10165);
and U13869 (N_13869,N_10076,N_11078);
nand U13870 (N_13870,N_9797,N_12226);
or U13871 (N_13871,N_12047,N_11961);
xnor U13872 (N_13872,N_11031,N_11828);
xnor U13873 (N_13873,N_11122,N_9819);
nand U13874 (N_13874,N_11709,N_11146);
nand U13875 (N_13875,N_12316,N_10757);
or U13876 (N_13876,N_12334,N_10590);
xnor U13877 (N_13877,N_9744,N_11953);
nand U13878 (N_13878,N_12434,N_12050);
nor U13879 (N_13879,N_11471,N_11198);
nor U13880 (N_13880,N_9662,N_10247);
nor U13881 (N_13881,N_12099,N_9824);
or U13882 (N_13882,N_10643,N_10095);
nor U13883 (N_13883,N_11015,N_11283);
nor U13884 (N_13884,N_11515,N_11571);
and U13885 (N_13885,N_12414,N_10650);
and U13886 (N_13886,N_12124,N_9713);
xor U13887 (N_13887,N_10382,N_10957);
or U13888 (N_13888,N_12369,N_9894);
and U13889 (N_13889,N_11640,N_11748);
xor U13890 (N_13890,N_10573,N_11661);
or U13891 (N_13891,N_11781,N_9948);
or U13892 (N_13892,N_10213,N_11145);
nand U13893 (N_13893,N_11898,N_10321);
xnor U13894 (N_13894,N_11246,N_12052);
nand U13895 (N_13895,N_9778,N_10343);
xnor U13896 (N_13896,N_12192,N_9987);
nor U13897 (N_13897,N_10546,N_11903);
nand U13898 (N_13898,N_10654,N_10982);
and U13899 (N_13899,N_12456,N_11156);
and U13900 (N_13900,N_9569,N_11679);
nor U13901 (N_13901,N_11472,N_12497);
and U13902 (N_13902,N_10267,N_12078);
and U13903 (N_13903,N_10936,N_10575);
xor U13904 (N_13904,N_9831,N_10571);
xnor U13905 (N_13905,N_11831,N_10947);
nor U13906 (N_13906,N_9621,N_9705);
nor U13907 (N_13907,N_9748,N_10461);
and U13908 (N_13908,N_11746,N_9836);
xor U13909 (N_13909,N_11873,N_9893);
nand U13910 (N_13910,N_10597,N_10818);
nor U13911 (N_13911,N_9833,N_11597);
nor U13912 (N_13912,N_11798,N_12431);
or U13913 (N_13913,N_9739,N_9399);
nor U13914 (N_13914,N_10114,N_12122);
nor U13915 (N_13915,N_12388,N_12475);
nor U13916 (N_13916,N_10727,N_10622);
xnor U13917 (N_13917,N_10545,N_10756);
nor U13918 (N_13918,N_12229,N_9976);
and U13919 (N_13919,N_10302,N_12086);
xor U13920 (N_13920,N_11766,N_10956);
nand U13921 (N_13921,N_10040,N_10079);
nand U13922 (N_13922,N_11542,N_10069);
nor U13923 (N_13923,N_10884,N_9766);
and U13924 (N_13924,N_10680,N_11226);
xor U13925 (N_13925,N_9393,N_11697);
or U13926 (N_13926,N_10231,N_11441);
nor U13927 (N_13927,N_11698,N_10408);
nand U13928 (N_13928,N_12461,N_10454);
nand U13929 (N_13929,N_11626,N_12405);
xnor U13930 (N_13930,N_10664,N_10615);
nor U13931 (N_13931,N_9803,N_9472);
or U13932 (N_13932,N_10864,N_9383);
xor U13933 (N_13933,N_10942,N_12156);
xor U13934 (N_13934,N_9996,N_10242);
xor U13935 (N_13935,N_9625,N_12161);
nand U13936 (N_13936,N_12257,N_11678);
or U13937 (N_13937,N_12069,N_10777);
nand U13938 (N_13938,N_9593,N_11980);
xnor U13939 (N_13939,N_10084,N_12371);
xor U13940 (N_13940,N_11608,N_10617);
xnor U13941 (N_13941,N_11780,N_11510);
xnor U13942 (N_13942,N_12103,N_10992);
xnor U13943 (N_13943,N_9462,N_12208);
or U13944 (N_13944,N_12116,N_10336);
xor U13945 (N_13945,N_11645,N_10292);
and U13946 (N_13946,N_12046,N_10392);
nor U13947 (N_13947,N_12202,N_9555);
and U13948 (N_13948,N_9471,N_12429);
or U13949 (N_13949,N_10203,N_12418);
nor U13950 (N_13950,N_11392,N_10484);
xnor U13951 (N_13951,N_10778,N_12342);
nand U13952 (N_13952,N_9646,N_9415);
and U13953 (N_13953,N_10306,N_10839);
xnor U13954 (N_13954,N_11917,N_10173);
xor U13955 (N_13955,N_11242,N_9376);
xnor U13956 (N_13956,N_9911,N_9756);
or U13957 (N_13957,N_10082,N_12081);
or U13958 (N_13958,N_11389,N_10307);
nor U13959 (N_13959,N_11262,N_10437);
and U13960 (N_13960,N_10558,N_10147);
nor U13961 (N_13961,N_10123,N_11880);
or U13962 (N_13962,N_10032,N_11349);
or U13963 (N_13963,N_11336,N_11012);
or U13964 (N_13964,N_10208,N_10097);
nand U13965 (N_13965,N_12148,N_11092);
nor U13966 (N_13966,N_9992,N_9979);
or U13967 (N_13967,N_12011,N_10008);
and U13968 (N_13968,N_11086,N_12287);
and U13969 (N_13969,N_9449,N_9750);
nand U13970 (N_13970,N_12002,N_11438);
xnor U13971 (N_13971,N_9859,N_11340);
nand U13972 (N_13972,N_10836,N_12210);
or U13973 (N_13973,N_12466,N_12230);
xnor U13974 (N_13974,N_9887,N_9583);
nor U13975 (N_13975,N_11653,N_10647);
or U13976 (N_13976,N_9755,N_11502);
or U13977 (N_13977,N_11893,N_11022);
xnor U13978 (N_13978,N_10094,N_11788);
nand U13979 (N_13979,N_12289,N_12262);
xor U13980 (N_13980,N_9908,N_10792);
xor U13981 (N_13981,N_10139,N_11233);
or U13982 (N_13982,N_12231,N_11793);
nor U13983 (N_13983,N_11566,N_12387);
or U13984 (N_13984,N_9626,N_11549);
nand U13985 (N_13985,N_9710,N_12209);
or U13986 (N_13986,N_10012,N_9817);
nor U13987 (N_13987,N_10776,N_10823);
nand U13988 (N_13988,N_12181,N_12350);
nor U13989 (N_13989,N_9514,N_10235);
and U13990 (N_13990,N_11432,N_10850);
or U13991 (N_13991,N_10478,N_9980);
nand U13992 (N_13992,N_9477,N_10471);
or U13993 (N_13993,N_11796,N_10226);
nor U13994 (N_13994,N_12085,N_11892);
nand U13995 (N_13995,N_9834,N_11231);
or U13996 (N_13996,N_11248,N_12326);
xor U13997 (N_13997,N_11711,N_11191);
or U13998 (N_13998,N_9418,N_11647);
xnor U13999 (N_13999,N_12083,N_10766);
and U14000 (N_14000,N_9641,N_12302);
and U14001 (N_14001,N_11585,N_11398);
nand U14002 (N_14002,N_11587,N_11439);
nor U14003 (N_14003,N_10620,N_9865);
nand U14004 (N_14004,N_11808,N_11528);
and U14005 (N_14005,N_11664,N_10195);
nor U14006 (N_14006,N_10891,N_10894);
nor U14007 (N_14007,N_9743,N_10205);
or U14008 (N_14008,N_11837,N_10354);
nand U14009 (N_14009,N_11955,N_11736);
xor U14010 (N_14010,N_9825,N_9657);
nor U14011 (N_14011,N_10881,N_9919);
nor U14012 (N_14012,N_10416,N_11069);
and U14013 (N_14013,N_10579,N_9924);
or U14014 (N_14014,N_11370,N_11303);
or U14015 (N_14015,N_11975,N_9856);
xnor U14016 (N_14016,N_11109,N_12365);
and U14017 (N_14017,N_10791,N_9655);
and U14018 (N_14018,N_10646,N_11175);
xnor U14019 (N_14019,N_9405,N_11556);
xor U14020 (N_14020,N_10753,N_12235);
or U14021 (N_14021,N_10150,N_11445);
and U14022 (N_14022,N_9726,N_10564);
or U14023 (N_14023,N_10044,N_10190);
nor U14024 (N_14024,N_11599,N_10447);
or U14025 (N_14025,N_9437,N_10826);
or U14026 (N_14026,N_11931,N_10003);
xor U14027 (N_14027,N_12272,N_10820);
and U14028 (N_14028,N_11481,N_9600);
and U14029 (N_14029,N_10702,N_9451);
or U14030 (N_14030,N_9428,N_11721);
xnor U14031 (N_14031,N_12175,N_11614);
nand U14032 (N_14032,N_9796,N_12256);
or U14033 (N_14033,N_12392,N_11867);
and U14034 (N_14034,N_10552,N_11309);
nand U14035 (N_14035,N_10338,N_10483);
xnor U14036 (N_14036,N_10534,N_11300);
or U14037 (N_14037,N_11288,N_11941);
nor U14038 (N_14038,N_11460,N_11852);
nor U14039 (N_14039,N_12449,N_9638);
nand U14040 (N_14040,N_12191,N_9505);
or U14041 (N_14041,N_9690,N_12149);
xnor U14042 (N_14042,N_9572,N_10315);
and U14043 (N_14043,N_10010,N_9953);
and U14044 (N_14044,N_10038,N_11497);
nand U14045 (N_14045,N_12066,N_9899);
nand U14046 (N_14046,N_9920,N_11986);
nor U14047 (N_14047,N_9508,N_10619);
nor U14048 (N_14048,N_10086,N_10409);
nor U14049 (N_14049,N_10598,N_11414);
xnor U14050 (N_14050,N_10693,N_11555);
or U14051 (N_14051,N_11677,N_12366);
or U14052 (N_14052,N_12068,N_11967);
xnor U14053 (N_14053,N_10880,N_10061);
or U14054 (N_14054,N_9406,N_10122);
or U14055 (N_14055,N_12437,N_9637);
xor U14056 (N_14056,N_10158,N_10520);
nor U14057 (N_14057,N_9970,N_9822);
nor U14058 (N_14058,N_10967,N_10143);
or U14059 (N_14059,N_10275,N_11003);
nor U14060 (N_14060,N_11511,N_11535);
and U14061 (N_14061,N_11450,N_11738);
xor U14062 (N_14062,N_12215,N_10361);
nand U14063 (N_14063,N_11757,N_10693);
nor U14064 (N_14064,N_11554,N_11179);
nand U14065 (N_14065,N_10637,N_9415);
or U14066 (N_14066,N_10036,N_12187);
xnor U14067 (N_14067,N_11226,N_10900);
and U14068 (N_14068,N_10963,N_11161);
nor U14069 (N_14069,N_11366,N_11442);
nand U14070 (N_14070,N_11703,N_10973);
nand U14071 (N_14071,N_11934,N_12419);
nand U14072 (N_14072,N_11655,N_10838);
xor U14073 (N_14073,N_9659,N_11434);
nor U14074 (N_14074,N_12403,N_10348);
nor U14075 (N_14075,N_10173,N_9927);
or U14076 (N_14076,N_10392,N_9999);
nand U14077 (N_14077,N_10996,N_10897);
nand U14078 (N_14078,N_11497,N_9418);
and U14079 (N_14079,N_11699,N_10655);
or U14080 (N_14080,N_11704,N_10759);
nor U14081 (N_14081,N_9560,N_9668);
xor U14082 (N_14082,N_9444,N_9455);
and U14083 (N_14083,N_11350,N_9816);
or U14084 (N_14084,N_9835,N_11489);
xnor U14085 (N_14085,N_11860,N_10638);
and U14086 (N_14086,N_12086,N_9995);
and U14087 (N_14087,N_9704,N_12093);
and U14088 (N_14088,N_10143,N_9525);
and U14089 (N_14089,N_10891,N_10960);
or U14090 (N_14090,N_9783,N_10511);
xor U14091 (N_14091,N_10105,N_10419);
or U14092 (N_14092,N_11819,N_10310);
xor U14093 (N_14093,N_11345,N_9506);
xnor U14094 (N_14094,N_12256,N_12173);
and U14095 (N_14095,N_11008,N_11882);
and U14096 (N_14096,N_10103,N_12456);
nor U14097 (N_14097,N_12448,N_9821);
and U14098 (N_14098,N_11344,N_11593);
or U14099 (N_14099,N_9497,N_10346);
xor U14100 (N_14100,N_9738,N_11012);
nor U14101 (N_14101,N_12022,N_12436);
xor U14102 (N_14102,N_11893,N_12194);
nor U14103 (N_14103,N_12251,N_9920);
nor U14104 (N_14104,N_11783,N_12365);
xnor U14105 (N_14105,N_11971,N_11294);
nand U14106 (N_14106,N_11394,N_10919);
or U14107 (N_14107,N_11901,N_12069);
and U14108 (N_14108,N_10116,N_11015);
nor U14109 (N_14109,N_9852,N_9402);
or U14110 (N_14110,N_11686,N_10438);
xor U14111 (N_14111,N_10392,N_10587);
nor U14112 (N_14112,N_10482,N_10081);
nand U14113 (N_14113,N_11288,N_12015);
xnor U14114 (N_14114,N_11391,N_10924);
and U14115 (N_14115,N_10430,N_10577);
nand U14116 (N_14116,N_10657,N_11792);
nand U14117 (N_14117,N_11666,N_12489);
and U14118 (N_14118,N_11705,N_10833);
xnor U14119 (N_14119,N_10100,N_10522);
and U14120 (N_14120,N_11473,N_10890);
nand U14121 (N_14121,N_10914,N_9530);
nor U14122 (N_14122,N_12478,N_9977);
xnor U14123 (N_14123,N_11431,N_11094);
or U14124 (N_14124,N_10482,N_11620);
nand U14125 (N_14125,N_11532,N_9700);
xor U14126 (N_14126,N_11273,N_9455);
or U14127 (N_14127,N_10969,N_10687);
nor U14128 (N_14128,N_10613,N_10833);
or U14129 (N_14129,N_10894,N_10908);
xor U14130 (N_14130,N_11730,N_10480);
nor U14131 (N_14131,N_10240,N_9486);
and U14132 (N_14132,N_10557,N_12445);
nor U14133 (N_14133,N_10642,N_9452);
nand U14134 (N_14134,N_10584,N_11346);
xor U14135 (N_14135,N_11480,N_10791);
and U14136 (N_14136,N_11276,N_11643);
nor U14137 (N_14137,N_11676,N_11076);
or U14138 (N_14138,N_11571,N_11332);
nand U14139 (N_14139,N_9837,N_11668);
or U14140 (N_14140,N_11246,N_9565);
nor U14141 (N_14141,N_12345,N_12001);
nand U14142 (N_14142,N_10330,N_9641);
xor U14143 (N_14143,N_10491,N_10262);
nor U14144 (N_14144,N_11787,N_10476);
and U14145 (N_14145,N_11596,N_11516);
and U14146 (N_14146,N_10195,N_9448);
nor U14147 (N_14147,N_12185,N_10593);
nor U14148 (N_14148,N_12366,N_10584);
and U14149 (N_14149,N_11274,N_11412);
xnor U14150 (N_14150,N_11464,N_9528);
nand U14151 (N_14151,N_10164,N_10764);
nand U14152 (N_14152,N_10901,N_10841);
nand U14153 (N_14153,N_11316,N_10081);
xnor U14154 (N_14154,N_11413,N_9632);
or U14155 (N_14155,N_10792,N_11830);
and U14156 (N_14156,N_9675,N_9943);
nor U14157 (N_14157,N_12308,N_10453);
nand U14158 (N_14158,N_12399,N_11843);
nor U14159 (N_14159,N_10330,N_12169);
xor U14160 (N_14160,N_11937,N_11268);
nor U14161 (N_14161,N_10732,N_9908);
xor U14162 (N_14162,N_11955,N_9872);
xor U14163 (N_14163,N_10631,N_10354);
nor U14164 (N_14164,N_10137,N_10752);
nand U14165 (N_14165,N_11497,N_11165);
nand U14166 (N_14166,N_9997,N_10623);
xnor U14167 (N_14167,N_12418,N_9496);
or U14168 (N_14168,N_12308,N_11943);
xnor U14169 (N_14169,N_9427,N_10937);
xnor U14170 (N_14170,N_9479,N_10912);
xnor U14171 (N_14171,N_9659,N_11129);
nor U14172 (N_14172,N_10512,N_10527);
nor U14173 (N_14173,N_12266,N_9445);
nor U14174 (N_14174,N_11638,N_12031);
nand U14175 (N_14175,N_11737,N_10988);
xor U14176 (N_14176,N_11598,N_11570);
or U14177 (N_14177,N_10560,N_9713);
nand U14178 (N_14178,N_10652,N_9630);
nor U14179 (N_14179,N_10167,N_10627);
or U14180 (N_14180,N_11821,N_10729);
or U14181 (N_14181,N_11728,N_9894);
nand U14182 (N_14182,N_10945,N_11632);
xor U14183 (N_14183,N_9499,N_12038);
or U14184 (N_14184,N_11363,N_11721);
and U14185 (N_14185,N_9400,N_10943);
xor U14186 (N_14186,N_11067,N_9897);
xor U14187 (N_14187,N_12362,N_11551);
xnor U14188 (N_14188,N_9406,N_12308);
and U14189 (N_14189,N_10478,N_11299);
xor U14190 (N_14190,N_9626,N_10079);
nand U14191 (N_14191,N_9646,N_10335);
or U14192 (N_14192,N_10387,N_10118);
xor U14193 (N_14193,N_10312,N_10708);
or U14194 (N_14194,N_11515,N_11356);
xnor U14195 (N_14195,N_11717,N_10173);
and U14196 (N_14196,N_9433,N_10286);
and U14197 (N_14197,N_11460,N_12084);
nand U14198 (N_14198,N_9761,N_9467);
and U14199 (N_14199,N_12264,N_12109);
nand U14200 (N_14200,N_12052,N_12302);
nor U14201 (N_14201,N_11734,N_10775);
xor U14202 (N_14202,N_10001,N_9656);
nand U14203 (N_14203,N_9465,N_10613);
xor U14204 (N_14204,N_11047,N_10526);
or U14205 (N_14205,N_10395,N_12478);
nor U14206 (N_14206,N_11994,N_9841);
or U14207 (N_14207,N_10132,N_11910);
or U14208 (N_14208,N_12390,N_10433);
nor U14209 (N_14209,N_10653,N_11053);
or U14210 (N_14210,N_12094,N_11618);
nand U14211 (N_14211,N_10002,N_11655);
xor U14212 (N_14212,N_11568,N_10761);
xnor U14213 (N_14213,N_12110,N_10621);
and U14214 (N_14214,N_11735,N_9442);
xor U14215 (N_14215,N_11996,N_9606);
nor U14216 (N_14216,N_9801,N_12433);
xnor U14217 (N_14217,N_9920,N_12446);
and U14218 (N_14218,N_11010,N_10010);
nor U14219 (N_14219,N_10094,N_11857);
nand U14220 (N_14220,N_9566,N_12014);
nand U14221 (N_14221,N_10057,N_10465);
nor U14222 (N_14222,N_10284,N_11438);
xor U14223 (N_14223,N_9576,N_10731);
and U14224 (N_14224,N_12398,N_10872);
nor U14225 (N_14225,N_9690,N_10220);
or U14226 (N_14226,N_10066,N_11681);
xnor U14227 (N_14227,N_10737,N_12319);
or U14228 (N_14228,N_9421,N_9599);
nand U14229 (N_14229,N_11105,N_12305);
and U14230 (N_14230,N_11656,N_9760);
xnor U14231 (N_14231,N_10545,N_10711);
xor U14232 (N_14232,N_9745,N_10415);
xor U14233 (N_14233,N_12292,N_11530);
and U14234 (N_14234,N_10662,N_11923);
and U14235 (N_14235,N_11224,N_11810);
nand U14236 (N_14236,N_10436,N_11204);
and U14237 (N_14237,N_9885,N_11711);
nand U14238 (N_14238,N_11811,N_10419);
and U14239 (N_14239,N_11409,N_10830);
or U14240 (N_14240,N_10880,N_12318);
nand U14241 (N_14241,N_11105,N_10479);
or U14242 (N_14242,N_9778,N_11694);
xor U14243 (N_14243,N_9485,N_10419);
xnor U14244 (N_14244,N_9422,N_12372);
nand U14245 (N_14245,N_11262,N_11932);
nor U14246 (N_14246,N_10349,N_12152);
nor U14247 (N_14247,N_9604,N_10232);
xor U14248 (N_14248,N_12131,N_11568);
xnor U14249 (N_14249,N_9929,N_9973);
nor U14250 (N_14250,N_10773,N_10167);
or U14251 (N_14251,N_10978,N_10793);
or U14252 (N_14252,N_9941,N_11443);
xnor U14253 (N_14253,N_9724,N_11741);
or U14254 (N_14254,N_9440,N_9705);
nor U14255 (N_14255,N_12384,N_11168);
nor U14256 (N_14256,N_9486,N_12222);
nand U14257 (N_14257,N_10298,N_12274);
and U14258 (N_14258,N_11154,N_10557);
xor U14259 (N_14259,N_9723,N_11875);
nand U14260 (N_14260,N_10011,N_10295);
nor U14261 (N_14261,N_10448,N_10333);
nand U14262 (N_14262,N_9982,N_9841);
nor U14263 (N_14263,N_10996,N_10023);
and U14264 (N_14264,N_10127,N_10410);
nand U14265 (N_14265,N_9942,N_12230);
xnor U14266 (N_14266,N_11388,N_11652);
nor U14267 (N_14267,N_11322,N_11501);
nor U14268 (N_14268,N_11293,N_11602);
or U14269 (N_14269,N_10094,N_10378);
xor U14270 (N_14270,N_9566,N_11376);
xnor U14271 (N_14271,N_9789,N_12360);
xor U14272 (N_14272,N_11241,N_11987);
or U14273 (N_14273,N_9628,N_12044);
and U14274 (N_14274,N_10048,N_9422);
nor U14275 (N_14275,N_10189,N_12373);
nand U14276 (N_14276,N_11648,N_12225);
and U14277 (N_14277,N_11296,N_9443);
and U14278 (N_14278,N_11963,N_10887);
xnor U14279 (N_14279,N_11077,N_10215);
nor U14280 (N_14280,N_9804,N_10235);
and U14281 (N_14281,N_9847,N_11563);
or U14282 (N_14282,N_11877,N_10712);
nor U14283 (N_14283,N_10713,N_11712);
or U14284 (N_14284,N_10784,N_12182);
nor U14285 (N_14285,N_10395,N_11635);
xnor U14286 (N_14286,N_11945,N_10707);
nand U14287 (N_14287,N_10369,N_11037);
nand U14288 (N_14288,N_9437,N_11029);
nor U14289 (N_14289,N_10111,N_11603);
nor U14290 (N_14290,N_11359,N_10186);
xnor U14291 (N_14291,N_10959,N_9837);
xnor U14292 (N_14292,N_9558,N_12237);
nand U14293 (N_14293,N_9868,N_11201);
xnor U14294 (N_14294,N_11613,N_11012);
nand U14295 (N_14295,N_11354,N_10919);
or U14296 (N_14296,N_10238,N_11132);
or U14297 (N_14297,N_11335,N_10294);
nor U14298 (N_14298,N_10095,N_10233);
or U14299 (N_14299,N_9676,N_11401);
nor U14300 (N_14300,N_9889,N_10828);
or U14301 (N_14301,N_10484,N_10015);
and U14302 (N_14302,N_11648,N_9608);
nor U14303 (N_14303,N_11029,N_10530);
nand U14304 (N_14304,N_10911,N_9423);
nor U14305 (N_14305,N_10020,N_11888);
xnor U14306 (N_14306,N_11116,N_10651);
or U14307 (N_14307,N_12126,N_10837);
nand U14308 (N_14308,N_12090,N_12116);
nand U14309 (N_14309,N_12417,N_12300);
nor U14310 (N_14310,N_9900,N_12167);
nand U14311 (N_14311,N_11696,N_12093);
and U14312 (N_14312,N_10911,N_10001);
xnor U14313 (N_14313,N_10666,N_10830);
nor U14314 (N_14314,N_12080,N_10093);
xor U14315 (N_14315,N_10167,N_11887);
and U14316 (N_14316,N_10638,N_11151);
nand U14317 (N_14317,N_10162,N_9579);
xor U14318 (N_14318,N_9964,N_10780);
nand U14319 (N_14319,N_11357,N_11263);
nand U14320 (N_14320,N_9568,N_11872);
nor U14321 (N_14321,N_11164,N_11592);
xnor U14322 (N_14322,N_9681,N_9469);
and U14323 (N_14323,N_11197,N_9528);
xnor U14324 (N_14324,N_9543,N_12493);
or U14325 (N_14325,N_9595,N_12399);
or U14326 (N_14326,N_10324,N_9383);
or U14327 (N_14327,N_11535,N_10659);
or U14328 (N_14328,N_9580,N_11937);
and U14329 (N_14329,N_9616,N_11558);
nor U14330 (N_14330,N_11248,N_11641);
and U14331 (N_14331,N_9684,N_11560);
xor U14332 (N_14332,N_10101,N_11708);
nand U14333 (N_14333,N_10747,N_11159);
nor U14334 (N_14334,N_11164,N_12195);
nand U14335 (N_14335,N_10424,N_11979);
xor U14336 (N_14336,N_9475,N_11974);
or U14337 (N_14337,N_9405,N_10499);
xor U14338 (N_14338,N_9789,N_12124);
and U14339 (N_14339,N_9475,N_10238);
or U14340 (N_14340,N_11137,N_11774);
and U14341 (N_14341,N_11500,N_9857);
nand U14342 (N_14342,N_9519,N_12248);
xor U14343 (N_14343,N_12342,N_11269);
nand U14344 (N_14344,N_12335,N_9760);
nor U14345 (N_14345,N_12397,N_11767);
xnor U14346 (N_14346,N_12410,N_11790);
and U14347 (N_14347,N_11273,N_11551);
nand U14348 (N_14348,N_11768,N_11470);
xor U14349 (N_14349,N_11480,N_10169);
or U14350 (N_14350,N_11143,N_9916);
xor U14351 (N_14351,N_11276,N_10455);
nand U14352 (N_14352,N_10940,N_9407);
or U14353 (N_14353,N_11803,N_9778);
xnor U14354 (N_14354,N_11730,N_12475);
nand U14355 (N_14355,N_9633,N_12293);
nor U14356 (N_14356,N_11673,N_10259);
and U14357 (N_14357,N_9406,N_10494);
xnor U14358 (N_14358,N_12231,N_11029);
or U14359 (N_14359,N_9472,N_11880);
nor U14360 (N_14360,N_10207,N_9933);
xor U14361 (N_14361,N_10116,N_11531);
or U14362 (N_14362,N_11201,N_10001);
xnor U14363 (N_14363,N_12067,N_12239);
and U14364 (N_14364,N_12194,N_9449);
or U14365 (N_14365,N_9495,N_10184);
nand U14366 (N_14366,N_9727,N_10296);
nand U14367 (N_14367,N_11542,N_11322);
or U14368 (N_14368,N_12437,N_9625);
and U14369 (N_14369,N_10431,N_12124);
nor U14370 (N_14370,N_11392,N_10412);
nand U14371 (N_14371,N_10144,N_12142);
or U14372 (N_14372,N_10657,N_10206);
xnor U14373 (N_14373,N_10193,N_12370);
xor U14374 (N_14374,N_12443,N_10966);
nand U14375 (N_14375,N_12340,N_11316);
and U14376 (N_14376,N_11531,N_10031);
or U14377 (N_14377,N_11076,N_10558);
nor U14378 (N_14378,N_12378,N_9790);
nor U14379 (N_14379,N_12009,N_12302);
and U14380 (N_14380,N_9860,N_11315);
and U14381 (N_14381,N_11300,N_10551);
or U14382 (N_14382,N_10356,N_12057);
xor U14383 (N_14383,N_10717,N_12005);
or U14384 (N_14384,N_11565,N_11959);
nand U14385 (N_14385,N_10339,N_10351);
xor U14386 (N_14386,N_11728,N_9428);
xnor U14387 (N_14387,N_11462,N_10956);
and U14388 (N_14388,N_11738,N_11311);
nor U14389 (N_14389,N_12253,N_12251);
nor U14390 (N_14390,N_12344,N_9695);
nor U14391 (N_14391,N_9508,N_9708);
nor U14392 (N_14392,N_10631,N_10923);
and U14393 (N_14393,N_10221,N_11720);
xnor U14394 (N_14394,N_10444,N_10993);
and U14395 (N_14395,N_10342,N_10901);
xnor U14396 (N_14396,N_10561,N_10588);
or U14397 (N_14397,N_11649,N_11761);
nand U14398 (N_14398,N_11860,N_12460);
and U14399 (N_14399,N_11274,N_10820);
or U14400 (N_14400,N_11622,N_12255);
or U14401 (N_14401,N_11599,N_10893);
nand U14402 (N_14402,N_12464,N_11008);
or U14403 (N_14403,N_11877,N_11739);
nor U14404 (N_14404,N_12332,N_11594);
xor U14405 (N_14405,N_12051,N_10194);
xor U14406 (N_14406,N_10923,N_10264);
nor U14407 (N_14407,N_9609,N_11497);
and U14408 (N_14408,N_9561,N_12116);
xor U14409 (N_14409,N_12490,N_10184);
and U14410 (N_14410,N_9565,N_11733);
xnor U14411 (N_14411,N_9916,N_12028);
or U14412 (N_14412,N_10981,N_12416);
and U14413 (N_14413,N_9768,N_9387);
nand U14414 (N_14414,N_10702,N_11578);
xnor U14415 (N_14415,N_10835,N_11568);
nand U14416 (N_14416,N_12123,N_12344);
nor U14417 (N_14417,N_12335,N_11104);
nor U14418 (N_14418,N_9627,N_9487);
and U14419 (N_14419,N_11647,N_10260);
xnor U14420 (N_14420,N_10265,N_11408);
xor U14421 (N_14421,N_12346,N_11503);
nor U14422 (N_14422,N_10029,N_11447);
xor U14423 (N_14423,N_10591,N_11667);
nor U14424 (N_14424,N_11807,N_10374);
and U14425 (N_14425,N_11057,N_11236);
xnor U14426 (N_14426,N_12405,N_11382);
or U14427 (N_14427,N_10648,N_11769);
nand U14428 (N_14428,N_11727,N_10092);
or U14429 (N_14429,N_9502,N_10947);
xnor U14430 (N_14430,N_12204,N_10566);
xnor U14431 (N_14431,N_11450,N_12238);
nor U14432 (N_14432,N_12081,N_10078);
xor U14433 (N_14433,N_9440,N_9583);
xnor U14434 (N_14434,N_11767,N_10628);
xor U14435 (N_14435,N_10571,N_11738);
nand U14436 (N_14436,N_11741,N_10510);
nor U14437 (N_14437,N_10499,N_9552);
nand U14438 (N_14438,N_10729,N_11775);
xor U14439 (N_14439,N_10201,N_10973);
or U14440 (N_14440,N_9470,N_11985);
and U14441 (N_14441,N_10784,N_11621);
nor U14442 (N_14442,N_10722,N_10974);
and U14443 (N_14443,N_12096,N_9600);
xnor U14444 (N_14444,N_9436,N_9399);
nor U14445 (N_14445,N_11930,N_11730);
nor U14446 (N_14446,N_9761,N_10797);
or U14447 (N_14447,N_11307,N_9909);
nor U14448 (N_14448,N_12353,N_9977);
and U14449 (N_14449,N_9438,N_11646);
xnor U14450 (N_14450,N_11691,N_10696);
xor U14451 (N_14451,N_12002,N_11610);
nor U14452 (N_14452,N_10404,N_12196);
nor U14453 (N_14453,N_10294,N_10023);
nand U14454 (N_14454,N_12109,N_12426);
and U14455 (N_14455,N_9904,N_10774);
nor U14456 (N_14456,N_10857,N_10370);
xnor U14457 (N_14457,N_12100,N_9878);
nor U14458 (N_14458,N_9463,N_10163);
or U14459 (N_14459,N_10721,N_11031);
xor U14460 (N_14460,N_10413,N_11261);
or U14461 (N_14461,N_12171,N_10937);
nand U14462 (N_14462,N_11766,N_9578);
nand U14463 (N_14463,N_10438,N_12451);
or U14464 (N_14464,N_11988,N_11181);
or U14465 (N_14465,N_11215,N_10491);
xnor U14466 (N_14466,N_12359,N_12009);
nor U14467 (N_14467,N_11754,N_11547);
nand U14468 (N_14468,N_10159,N_12263);
and U14469 (N_14469,N_9640,N_12231);
or U14470 (N_14470,N_9773,N_10032);
and U14471 (N_14471,N_10210,N_12189);
and U14472 (N_14472,N_9886,N_10959);
and U14473 (N_14473,N_11090,N_12149);
and U14474 (N_14474,N_10138,N_9752);
xnor U14475 (N_14475,N_10540,N_10597);
xor U14476 (N_14476,N_12436,N_10002);
or U14477 (N_14477,N_10418,N_10093);
nand U14478 (N_14478,N_10247,N_11316);
nand U14479 (N_14479,N_10198,N_11785);
and U14480 (N_14480,N_11630,N_11019);
or U14481 (N_14481,N_11112,N_10854);
nand U14482 (N_14482,N_12224,N_12333);
nand U14483 (N_14483,N_10002,N_11582);
xnor U14484 (N_14484,N_9478,N_10788);
and U14485 (N_14485,N_9602,N_11511);
xor U14486 (N_14486,N_11443,N_9526);
xnor U14487 (N_14487,N_12131,N_9907);
nand U14488 (N_14488,N_11263,N_9844);
nand U14489 (N_14489,N_10555,N_10969);
and U14490 (N_14490,N_11702,N_10993);
nor U14491 (N_14491,N_11206,N_11728);
or U14492 (N_14492,N_10769,N_11792);
and U14493 (N_14493,N_10535,N_11648);
xor U14494 (N_14494,N_11985,N_11488);
or U14495 (N_14495,N_11801,N_10838);
nor U14496 (N_14496,N_10586,N_12051);
nor U14497 (N_14497,N_10086,N_9964);
nand U14498 (N_14498,N_10556,N_10222);
and U14499 (N_14499,N_12053,N_10687);
xor U14500 (N_14500,N_10941,N_11381);
nand U14501 (N_14501,N_11579,N_11599);
xor U14502 (N_14502,N_10336,N_11314);
or U14503 (N_14503,N_9613,N_11050);
and U14504 (N_14504,N_11245,N_9503);
or U14505 (N_14505,N_9703,N_9377);
nand U14506 (N_14506,N_9546,N_11512);
and U14507 (N_14507,N_12178,N_9587);
or U14508 (N_14508,N_9964,N_11916);
nor U14509 (N_14509,N_11194,N_11286);
or U14510 (N_14510,N_11996,N_11900);
nor U14511 (N_14511,N_10935,N_10477);
nor U14512 (N_14512,N_9952,N_10135);
xnor U14513 (N_14513,N_10846,N_11928);
nor U14514 (N_14514,N_10746,N_10906);
or U14515 (N_14515,N_11646,N_10789);
nor U14516 (N_14516,N_10000,N_9658);
nor U14517 (N_14517,N_11389,N_11209);
xor U14518 (N_14518,N_10041,N_11377);
nor U14519 (N_14519,N_10465,N_10318);
or U14520 (N_14520,N_11969,N_11496);
nor U14521 (N_14521,N_10379,N_12128);
xnor U14522 (N_14522,N_10342,N_10892);
nor U14523 (N_14523,N_10040,N_10662);
nor U14524 (N_14524,N_9610,N_12144);
and U14525 (N_14525,N_11558,N_11829);
nor U14526 (N_14526,N_12278,N_10790);
nor U14527 (N_14527,N_10129,N_11228);
nand U14528 (N_14528,N_10211,N_10678);
nand U14529 (N_14529,N_10738,N_11250);
or U14530 (N_14530,N_9830,N_12064);
or U14531 (N_14531,N_10577,N_12094);
or U14532 (N_14532,N_11827,N_9911);
xor U14533 (N_14533,N_10511,N_11989);
nor U14534 (N_14534,N_9582,N_12383);
or U14535 (N_14535,N_11007,N_12366);
and U14536 (N_14536,N_11364,N_10869);
nand U14537 (N_14537,N_11286,N_10309);
xnor U14538 (N_14538,N_10471,N_11335);
and U14539 (N_14539,N_11121,N_10472);
xor U14540 (N_14540,N_11383,N_9426);
nand U14541 (N_14541,N_9518,N_12411);
nand U14542 (N_14542,N_10179,N_12333);
nand U14543 (N_14543,N_11111,N_10854);
nor U14544 (N_14544,N_9709,N_11610);
nor U14545 (N_14545,N_9380,N_12132);
xor U14546 (N_14546,N_9555,N_12286);
or U14547 (N_14547,N_11954,N_10213);
xnor U14548 (N_14548,N_10420,N_11006);
xor U14549 (N_14549,N_12479,N_10510);
nor U14550 (N_14550,N_11776,N_10670);
nor U14551 (N_14551,N_10364,N_9543);
xor U14552 (N_14552,N_12023,N_10364);
and U14553 (N_14553,N_10877,N_10301);
xor U14554 (N_14554,N_10292,N_10389);
nor U14555 (N_14555,N_10760,N_10228);
xnor U14556 (N_14556,N_10360,N_10922);
xnor U14557 (N_14557,N_9605,N_12019);
nand U14558 (N_14558,N_10674,N_11499);
or U14559 (N_14559,N_9579,N_10978);
xnor U14560 (N_14560,N_11821,N_12217);
and U14561 (N_14561,N_10320,N_10513);
or U14562 (N_14562,N_10344,N_10877);
nor U14563 (N_14563,N_10037,N_9474);
nor U14564 (N_14564,N_10192,N_11617);
and U14565 (N_14565,N_10055,N_11475);
nand U14566 (N_14566,N_11930,N_9405);
nand U14567 (N_14567,N_9765,N_10267);
nand U14568 (N_14568,N_11707,N_11965);
nor U14569 (N_14569,N_11749,N_10913);
xnor U14570 (N_14570,N_11098,N_11622);
nor U14571 (N_14571,N_9962,N_10238);
or U14572 (N_14572,N_12196,N_9636);
or U14573 (N_14573,N_10694,N_12178);
nor U14574 (N_14574,N_12214,N_10655);
or U14575 (N_14575,N_12333,N_11198);
xor U14576 (N_14576,N_11383,N_10614);
or U14577 (N_14577,N_11415,N_9678);
xor U14578 (N_14578,N_11025,N_9728);
nor U14579 (N_14579,N_11236,N_11836);
nor U14580 (N_14580,N_10553,N_10155);
nor U14581 (N_14581,N_11932,N_10479);
and U14582 (N_14582,N_10400,N_12298);
nor U14583 (N_14583,N_10751,N_12142);
nand U14584 (N_14584,N_10698,N_11271);
nor U14585 (N_14585,N_9555,N_11338);
or U14586 (N_14586,N_10726,N_11258);
and U14587 (N_14587,N_12043,N_11767);
and U14588 (N_14588,N_12132,N_10720);
nand U14589 (N_14589,N_12044,N_10614);
or U14590 (N_14590,N_9945,N_11579);
nand U14591 (N_14591,N_9416,N_12150);
xnor U14592 (N_14592,N_10089,N_9767);
nor U14593 (N_14593,N_10035,N_11229);
or U14594 (N_14594,N_12356,N_9604);
or U14595 (N_14595,N_12454,N_9835);
and U14596 (N_14596,N_10441,N_11740);
or U14597 (N_14597,N_9936,N_11899);
nand U14598 (N_14598,N_10737,N_10657);
xor U14599 (N_14599,N_11246,N_9406);
or U14600 (N_14600,N_11591,N_11489);
nand U14601 (N_14601,N_9425,N_11405);
and U14602 (N_14602,N_12056,N_10524);
nand U14603 (N_14603,N_9924,N_11632);
and U14604 (N_14604,N_11467,N_12327);
nand U14605 (N_14605,N_10008,N_11761);
or U14606 (N_14606,N_10209,N_9611);
nand U14607 (N_14607,N_12496,N_11611);
nand U14608 (N_14608,N_9979,N_12055);
or U14609 (N_14609,N_9449,N_10447);
xor U14610 (N_14610,N_11935,N_12224);
nor U14611 (N_14611,N_11758,N_11368);
nand U14612 (N_14612,N_10149,N_12383);
or U14613 (N_14613,N_9458,N_9713);
xnor U14614 (N_14614,N_12119,N_11654);
or U14615 (N_14615,N_12228,N_10649);
xor U14616 (N_14616,N_11647,N_10174);
xnor U14617 (N_14617,N_11113,N_12037);
and U14618 (N_14618,N_12284,N_10551);
nor U14619 (N_14619,N_11832,N_11290);
and U14620 (N_14620,N_12324,N_10661);
nor U14621 (N_14621,N_10861,N_12098);
and U14622 (N_14622,N_10389,N_11669);
xor U14623 (N_14623,N_11343,N_9694);
nand U14624 (N_14624,N_11095,N_11244);
and U14625 (N_14625,N_12330,N_10299);
xor U14626 (N_14626,N_12143,N_10148);
xor U14627 (N_14627,N_11728,N_9567);
nor U14628 (N_14628,N_11587,N_12050);
or U14629 (N_14629,N_9405,N_11536);
or U14630 (N_14630,N_10329,N_10807);
or U14631 (N_14631,N_9975,N_11780);
nor U14632 (N_14632,N_10128,N_9889);
or U14633 (N_14633,N_9929,N_11598);
nor U14634 (N_14634,N_10611,N_11551);
nand U14635 (N_14635,N_10893,N_12014);
nand U14636 (N_14636,N_9748,N_10691);
xor U14637 (N_14637,N_12392,N_11009);
and U14638 (N_14638,N_10695,N_9831);
xor U14639 (N_14639,N_9425,N_10940);
or U14640 (N_14640,N_9969,N_10019);
nor U14641 (N_14641,N_12452,N_12498);
and U14642 (N_14642,N_11945,N_11682);
nor U14643 (N_14643,N_12100,N_11595);
nand U14644 (N_14644,N_11051,N_11263);
xor U14645 (N_14645,N_10312,N_9564);
xnor U14646 (N_14646,N_11216,N_10683);
nand U14647 (N_14647,N_10745,N_9697);
and U14648 (N_14648,N_9413,N_9758);
and U14649 (N_14649,N_12304,N_10635);
xor U14650 (N_14650,N_10282,N_10515);
or U14651 (N_14651,N_10543,N_10641);
nand U14652 (N_14652,N_10658,N_10549);
nor U14653 (N_14653,N_10240,N_9641);
or U14654 (N_14654,N_11508,N_10547);
xor U14655 (N_14655,N_10177,N_11555);
and U14656 (N_14656,N_11706,N_12200);
xnor U14657 (N_14657,N_9471,N_11597);
nor U14658 (N_14658,N_10305,N_9526);
nand U14659 (N_14659,N_9854,N_12000);
nand U14660 (N_14660,N_12452,N_10623);
or U14661 (N_14661,N_10357,N_11606);
and U14662 (N_14662,N_11308,N_10458);
nand U14663 (N_14663,N_10435,N_12117);
nand U14664 (N_14664,N_12122,N_12234);
and U14665 (N_14665,N_9421,N_10527);
xnor U14666 (N_14666,N_10478,N_12467);
xnor U14667 (N_14667,N_10572,N_12481);
or U14668 (N_14668,N_12271,N_10913);
nand U14669 (N_14669,N_11381,N_9430);
or U14670 (N_14670,N_12128,N_9992);
and U14671 (N_14671,N_12101,N_9853);
or U14672 (N_14672,N_10062,N_9699);
nand U14673 (N_14673,N_9808,N_11117);
xor U14674 (N_14674,N_12188,N_11883);
nor U14675 (N_14675,N_12047,N_10528);
xor U14676 (N_14676,N_10017,N_11696);
nor U14677 (N_14677,N_9761,N_12126);
nand U14678 (N_14678,N_10610,N_9977);
xor U14679 (N_14679,N_10505,N_12287);
xor U14680 (N_14680,N_12011,N_9907);
nand U14681 (N_14681,N_12308,N_10517);
and U14682 (N_14682,N_10249,N_10165);
or U14683 (N_14683,N_9599,N_12476);
nand U14684 (N_14684,N_11253,N_10471);
or U14685 (N_14685,N_9411,N_11750);
xnor U14686 (N_14686,N_10017,N_10412);
xnor U14687 (N_14687,N_11051,N_10708);
and U14688 (N_14688,N_11153,N_10724);
nand U14689 (N_14689,N_10118,N_12147);
or U14690 (N_14690,N_12091,N_10264);
and U14691 (N_14691,N_9843,N_10935);
or U14692 (N_14692,N_11966,N_10204);
nor U14693 (N_14693,N_11831,N_11415);
nor U14694 (N_14694,N_11759,N_10405);
and U14695 (N_14695,N_9868,N_11314);
or U14696 (N_14696,N_10891,N_12217);
or U14697 (N_14697,N_10652,N_10811);
and U14698 (N_14698,N_9923,N_10572);
nand U14699 (N_14699,N_10242,N_12341);
or U14700 (N_14700,N_9715,N_12103);
or U14701 (N_14701,N_11113,N_10004);
nor U14702 (N_14702,N_9443,N_10288);
nand U14703 (N_14703,N_11147,N_9614);
nor U14704 (N_14704,N_10992,N_10600);
or U14705 (N_14705,N_11001,N_10392);
and U14706 (N_14706,N_9983,N_10447);
or U14707 (N_14707,N_10241,N_9661);
nand U14708 (N_14708,N_10137,N_10281);
nand U14709 (N_14709,N_11657,N_10316);
xnor U14710 (N_14710,N_12411,N_11111);
xor U14711 (N_14711,N_9472,N_12024);
nand U14712 (N_14712,N_9692,N_12395);
xor U14713 (N_14713,N_12454,N_10971);
nand U14714 (N_14714,N_9397,N_11457);
or U14715 (N_14715,N_10021,N_10631);
nand U14716 (N_14716,N_10900,N_10044);
and U14717 (N_14717,N_11625,N_12285);
nand U14718 (N_14718,N_10178,N_10791);
or U14719 (N_14719,N_11388,N_9818);
nand U14720 (N_14720,N_11416,N_11195);
or U14721 (N_14721,N_10016,N_11703);
xor U14722 (N_14722,N_11071,N_11619);
xor U14723 (N_14723,N_9685,N_10914);
xnor U14724 (N_14724,N_10689,N_12403);
nor U14725 (N_14725,N_9786,N_11881);
and U14726 (N_14726,N_10896,N_10399);
xnor U14727 (N_14727,N_9837,N_9473);
xnor U14728 (N_14728,N_10022,N_10747);
nand U14729 (N_14729,N_10438,N_12039);
and U14730 (N_14730,N_11485,N_9375);
nor U14731 (N_14731,N_10438,N_10167);
or U14732 (N_14732,N_11506,N_10472);
nand U14733 (N_14733,N_9753,N_9437);
nor U14734 (N_14734,N_11918,N_10384);
nor U14735 (N_14735,N_10671,N_11212);
xor U14736 (N_14736,N_10419,N_12270);
nand U14737 (N_14737,N_10845,N_9924);
or U14738 (N_14738,N_11561,N_10879);
nor U14739 (N_14739,N_10471,N_10126);
or U14740 (N_14740,N_10507,N_9524);
nor U14741 (N_14741,N_12003,N_11601);
xor U14742 (N_14742,N_10409,N_10978);
nor U14743 (N_14743,N_10580,N_9887);
xor U14744 (N_14744,N_11380,N_11800);
nor U14745 (N_14745,N_9430,N_10246);
and U14746 (N_14746,N_10916,N_12108);
and U14747 (N_14747,N_12155,N_9504);
and U14748 (N_14748,N_11827,N_9586);
nand U14749 (N_14749,N_10700,N_10318);
nand U14750 (N_14750,N_9717,N_9470);
or U14751 (N_14751,N_10940,N_12194);
and U14752 (N_14752,N_10238,N_10205);
and U14753 (N_14753,N_12021,N_10705);
and U14754 (N_14754,N_12390,N_10334);
nor U14755 (N_14755,N_9735,N_10927);
nand U14756 (N_14756,N_11881,N_12122);
nor U14757 (N_14757,N_9906,N_10979);
xor U14758 (N_14758,N_10147,N_9846);
nand U14759 (N_14759,N_12250,N_11252);
nor U14760 (N_14760,N_12012,N_10835);
xnor U14761 (N_14761,N_11088,N_11217);
nand U14762 (N_14762,N_11006,N_11675);
or U14763 (N_14763,N_11873,N_11018);
nand U14764 (N_14764,N_11306,N_10359);
xor U14765 (N_14765,N_9998,N_11782);
and U14766 (N_14766,N_9701,N_11099);
nand U14767 (N_14767,N_9634,N_11518);
nand U14768 (N_14768,N_11321,N_12307);
or U14769 (N_14769,N_11423,N_11424);
and U14770 (N_14770,N_9564,N_10427);
or U14771 (N_14771,N_10023,N_10731);
nor U14772 (N_14772,N_12200,N_10656);
or U14773 (N_14773,N_11088,N_10011);
xor U14774 (N_14774,N_9594,N_11616);
nand U14775 (N_14775,N_10417,N_11496);
nor U14776 (N_14776,N_10085,N_10530);
xor U14777 (N_14777,N_10830,N_10571);
nand U14778 (N_14778,N_12182,N_10175);
xnor U14779 (N_14779,N_11180,N_12134);
nand U14780 (N_14780,N_9758,N_12311);
nand U14781 (N_14781,N_11496,N_12487);
and U14782 (N_14782,N_10383,N_11367);
xor U14783 (N_14783,N_10429,N_10076);
nand U14784 (N_14784,N_10018,N_10418);
nand U14785 (N_14785,N_10335,N_9755);
nor U14786 (N_14786,N_11888,N_11412);
nor U14787 (N_14787,N_12452,N_11339);
and U14788 (N_14788,N_10666,N_10083);
or U14789 (N_14789,N_11529,N_9840);
nand U14790 (N_14790,N_11463,N_9558);
xor U14791 (N_14791,N_11514,N_9573);
xor U14792 (N_14792,N_9452,N_11147);
and U14793 (N_14793,N_11326,N_11961);
or U14794 (N_14794,N_11462,N_9557);
nand U14795 (N_14795,N_11853,N_12319);
nor U14796 (N_14796,N_11718,N_10001);
or U14797 (N_14797,N_11324,N_10777);
or U14798 (N_14798,N_11427,N_10325);
or U14799 (N_14799,N_10468,N_12301);
xnor U14800 (N_14800,N_10352,N_10057);
nor U14801 (N_14801,N_12008,N_10460);
nor U14802 (N_14802,N_11935,N_12045);
nor U14803 (N_14803,N_11147,N_9801);
xor U14804 (N_14804,N_10935,N_9865);
and U14805 (N_14805,N_11074,N_11386);
nor U14806 (N_14806,N_11336,N_12286);
nor U14807 (N_14807,N_12386,N_9381);
xor U14808 (N_14808,N_11213,N_9685);
nor U14809 (N_14809,N_10060,N_9680);
and U14810 (N_14810,N_12296,N_9467);
and U14811 (N_14811,N_12037,N_10457);
xor U14812 (N_14812,N_12318,N_11077);
and U14813 (N_14813,N_12407,N_11402);
xor U14814 (N_14814,N_10758,N_12100);
nand U14815 (N_14815,N_10438,N_11725);
nor U14816 (N_14816,N_10506,N_11125);
and U14817 (N_14817,N_10210,N_11925);
nand U14818 (N_14818,N_12307,N_11477);
xnor U14819 (N_14819,N_9497,N_11249);
and U14820 (N_14820,N_10461,N_9614);
nor U14821 (N_14821,N_10667,N_11979);
nor U14822 (N_14822,N_10512,N_11344);
and U14823 (N_14823,N_10350,N_9757);
nand U14824 (N_14824,N_12367,N_12000);
xor U14825 (N_14825,N_11972,N_9382);
and U14826 (N_14826,N_10218,N_12335);
xnor U14827 (N_14827,N_9871,N_12102);
and U14828 (N_14828,N_10441,N_10484);
and U14829 (N_14829,N_12092,N_12376);
nor U14830 (N_14830,N_11565,N_10783);
nor U14831 (N_14831,N_12407,N_9670);
nand U14832 (N_14832,N_10118,N_11205);
or U14833 (N_14833,N_11236,N_10174);
nand U14834 (N_14834,N_11668,N_12218);
nand U14835 (N_14835,N_10199,N_9727);
nor U14836 (N_14836,N_11671,N_10489);
xor U14837 (N_14837,N_9837,N_10758);
xnor U14838 (N_14838,N_11439,N_11204);
and U14839 (N_14839,N_9979,N_10500);
nand U14840 (N_14840,N_10463,N_11505);
nand U14841 (N_14841,N_10754,N_9923);
nor U14842 (N_14842,N_9722,N_12038);
and U14843 (N_14843,N_9774,N_9789);
nor U14844 (N_14844,N_10487,N_10105);
and U14845 (N_14845,N_12067,N_10082);
xnor U14846 (N_14846,N_12137,N_11066);
and U14847 (N_14847,N_10592,N_10632);
xnor U14848 (N_14848,N_12172,N_11846);
and U14849 (N_14849,N_9514,N_11133);
nand U14850 (N_14850,N_9776,N_10616);
and U14851 (N_14851,N_11319,N_11217);
xnor U14852 (N_14852,N_10351,N_11991);
and U14853 (N_14853,N_9929,N_11399);
nand U14854 (N_14854,N_9721,N_10631);
or U14855 (N_14855,N_12036,N_10934);
nor U14856 (N_14856,N_11345,N_12132);
nor U14857 (N_14857,N_9965,N_10781);
or U14858 (N_14858,N_10925,N_12069);
nand U14859 (N_14859,N_11295,N_11237);
nor U14860 (N_14860,N_10825,N_10238);
xnor U14861 (N_14861,N_10530,N_10403);
or U14862 (N_14862,N_11769,N_11781);
and U14863 (N_14863,N_11137,N_12281);
nand U14864 (N_14864,N_12316,N_11291);
nand U14865 (N_14865,N_10123,N_9954);
or U14866 (N_14866,N_10126,N_10517);
nand U14867 (N_14867,N_10017,N_11380);
nand U14868 (N_14868,N_11741,N_10195);
xnor U14869 (N_14869,N_11251,N_9378);
and U14870 (N_14870,N_9657,N_9446);
nand U14871 (N_14871,N_12032,N_12458);
and U14872 (N_14872,N_12310,N_10533);
or U14873 (N_14873,N_11495,N_10763);
nand U14874 (N_14874,N_9674,N_9740);
xor U14875 (N_14875,N_10374,N_11395);
nor U14876 (N_14876,N_12314,N_12322);
xnor U14877 (N_14877,N_10938,N_11713);
xor U14878 (N_14878,N_11334,N_12398);
nor U14879 (N_14879,N_10478,N_10371);
nand U14880 (N_14880,N_9505,N_9560);
or U14881 (N_14881,N_12049,N_11596);
and U14882 (N_14882,N_10276,N_11938);
and U14883 (N_14883,N_9377,N_12424);
nor U14884 (N_14884,N_10015,N_9508);
nor U14885 (N_14885,N_11601,N_10100);
nand U14886 (N_14886,N_10140,N_11719);
nand U14887 (N_14887,N_9422,N_9424);
or U14888 (N_14888,N_10599,N_10045);
xnor U14889 (N_14889,N_9609,N_9384);
or U14890 (N_14890,N_11485,N_10029);
nand U14891 (N_14891,N_10580,N_10236);
nor U14892 (N_14892,N_10572,N_11339);
or U14893 (N_14893,N_12465,N_10468);
xnor U14894 (N_14894,N_10382,N_10905);
or U14895 (N_14895,N_11435,N_10594);
xnor U14896 (N_14896,N_11913,N_10754);
nand U14897 (N_14897,N_12215,N_11731);
and U14898 (N_14898,N_10940,N_10183);
nand U14899 (N_14899,N_10875,N_9850);
xor U14900 (N_14900,N_11092,N_11843);
nand U14901 (N_14901,N_12168,N_11691);
and U14902 (N_14902,N_12353,N_9449);
and U14903 (N_14903,N_10078,N_10255);
or U14904 (N_14904,N_10883,N_10099);
nand U14905 (N_14905,N_10024,N_10803);
nor U14906 (N_14906,N_10186,N_9509);
nor U14907 (N_14907,N_10840,N_11419);
nor U14908 (N_14908,N_11468,N_10098);
nand U14909 (N_14909,N_10164,N_10055);
and U14910 (N_14910,N_9526,N_11180);
and U14911 (N_14911,N_9900,N_11944);
or U14912 (N_14912,N_9410,N_11112);
or U14913 (N_14913,N_12253,N_10388);
nor U14914 (N_14914,N_11081,N_10829);
nand U14915 (N_14915,N_11554,N_9644);
xor U14916 (N_14916,N_12128,N_11103);
nand U14917 (N_14917,N_9570,N_11157);
nand U14918 (N_14918,N_10389,N_10316);
xor U14919 (N_14919,N_9841,N_11816);
nor U14920 (N_14920,N_9967,N_10561);
nor U14921 (N_14921,N_9704,N_9974);
nor U14922 (N_14922,N_10289,N_11306);
and U14923 (N_14923,N_9705,N_10032);
and U14924 (N_14924,N_9682,N_10924);
nor U14925 (N_14925,N_9976,N_11423);
and U14926 (N_14926,N_11805,N_11675);
and U14927 (N_14927,N_11139,N_11194);
nor U14928 (N_14928,N_9383,N_10442);
or U14929 (N_14929,N_9646,N_9418);
xor U14930 (N_14930,N_12106,N_12265);
or U14931 (N_14931,N_10010,N_11954);
nand U14932 (N_14932,N_9549,N_10409);
and U14933 (N_14933,N_10364,N_11754);
nand U14934 (N_14934,N_11670,N_10670);
and U14935 (N_14935,N_11682,N_10124);
or U14936 (N_14936,N_10958,N_10492);
nand U14937 (N_14937,N_9584,N_11197);
xor U14938 (N_14938,N_11502,N_11137);
and U14939 (N_14939,N_11932,N_11280);
nor U14940 (N_14940,N_11831,N_11827);
xor U14941 (N_14941,N_11122,N_12481);
xor U14942 (N_14942,N_9980,N_12110);
nor U14943 (N_14943,N_12113,N_10249);
nand U14944 (N_14944,N_10896,N_10320);
nand U14945 (N_14945,N_9670,N_10528);
xor U14946 (N_14946,N_11954,N_9525);
xnor U14947 (N_14947,N_10329,N_9444);
nor U14948 (N_14948,N_10074,N_10605);
and U14949 (N_14949,N_12181,N_11527);
nand U14950 (N_14950,N_10756,N_12197);
xor U14951 (N_14951,N_12016,N_10148);
and U14952 (N_14952,N_12262,N_11234);
xnor U14953 (N_14953,N_10958,N_9650);
nor U14954 (N_14954,N_10938,N_10853);
or U14955 (N_14955,N_9946,N_9421);
and U14956 (N_14956,N_11912,N_10766);
or U14957 (N_14957,N_9692,N_9966);
nand U14958 (N_14958,N_12199,N_12302);
nor U14959 (N_14959,N_12418,N_12349);
xor U14960 (N_14960,N_10028,N_12221);
or U14961 (N_14961,N_10950,N_9434);
nand U14962 (N_14962,N_10830,N_10861);
and U14963 (N_14963,N_12082,N_9722);
or U14964 (N_14964,N_10517,N_9524);
or U14965 (N_14965,N_12402,N_11928);
or U14966 (N_14966,N_11193,N_10841);
and U14967 (N_14967,N_9932,N_11472);
xor U14968 (N_14968,N_10710,N_11576);
nor U14969 (N_14969,N_9426,N_10267);
and U14970 (N_14970,N_11903,N_10536);
nor U14971 (N_14971,N_10938,N_11901);
nor U14972 (N_14972,N_11675,N_9566);
nor U14973 (N_14973,N_10046,N_12241);
xor U14974 (N_14974,N_11122,N_11571);
and U14975 (N_14975,N_12013,N_9472);
nand U14976 (N_14976,N_10679,N_9758);
and U14977 (N_14977,N_10717,N_9766);
xnor U14978 (N_14978,N_11342,N_11761);
nor U14979 (N_14979,N_11872,N_9379);
xor U14980 (N_14980,N_12209,N_10180);
nand U14981 (N_14981,N_9614,N_11255);
or U14982 (N_14982,N_11657,N_11738);
and U14983 (N_14983,N_11964,N_10468);
xnor U14984 (N_14984,N_10808,N_10355);
xnor U14985 (N_14985,N_12153,N_12349);
or U14986 (N_14986,N_11598,N_9404);
xnor U14987 (N_14987,N_10203,N_11251);
and U14988 (N_14988,N_11827,N_11480);
or U14989 (N_14989,N_9878,N_10600);
and U14990 (N_14990,N_9640,N_9807);
and U14991 (N_14991,N_11312,N_11180);
nand U14992 (N_14992,N_11155,N_10340);
or U14993 (N_14993,N_9943,N_10063);
nand U14994 (N_14994,N_9808,N_12077);
xnor U14995 (N_14995,N_12003,N_12314);
nor U14996 (N_14996,N_12177,N_11704);
nor U14997 (N_14997,N_12339,N_10945);
nand U14998 (N_14998,N_12371,N_12082);
xnor U14999 (N_14999,N_9937,N_10340);
xor U15000 (N_15000,N_12360,N_9902);
and U15001 (N_15001,N_11294,N_10104);
and U15002 (N_15002,N_10453,N_12001);
and U15003 (N_15003,N_10694,N_10631);
nor U15004 (N_15004,N_11255,N_11490);
xnor U15005 (N_15005,N_11991,N_9954);
nor U15006 (N_15006,N_10217,N_10819);
xnor U15007 (N_15007,N_10316,N_10356);
or U15008 (N_15008,N_12250,N_11510);
xor U15009 (N_15009,N_11944,N_9713);
or U15010 (N_15010,N_10746,N_10347);
nor U15011 (N_15011,N_12393,N_11213);
xor U15012 (N_15012,N_10545,N_12060);
nand U15013 (N_15013,N_11396,N_10559);
nor U15014 (N_15014,N_12179,N_11809);
and U15015 (N_15015,N_10314,N_10422);
nor U15016 (N_15016,N_12111,N_12266);
and U15017 (N_15017,N_10333,N_11207);
xor U15018 (N_15018,N_10361,N_9993);
xor U15019 (N_15019,N_10914,N_12449);
nor U15020 (N_15020,N_11782,N_11754);
xnor U15021 (N_15021,N_10954,N_11659);
xnor U15022 (N_15022,N_11760,N_11695);
nand U15023 (N_15023,N_9824,N_12025);
or U15024 (N_15024,N_10163,N_11457);
nand U15025 (N_15025,N_9968,N_10956);
xnor U15026 (N_15026,N_10392,N_9942);
and U15027 (N_15027,N_12377,N_12288);
or U15028 (N_15028,N_12167,N_12445);
nand U15029 (N_15029,N_10005,N_10176);
and U15030 (N_15030,N_11395,N_11604);
nor U15031 (N_15031,N_10268,N_10549);
or U15032 (N_15032,N_11997,N_10894);
nand U15033 (N_15033,N_10581,N_12340);
nand U15034 (N_15034,N_9961,N_10855);
xnor U15035 (N_15035,N_11909,N_9975);
xnor U15036 (N_15036,N_11547,N_12227);
and U15037 (N_15037,N_11529,N_9534);
nor U15038 (N_15038,N_12263,N_9396);
nand U15039 (N_15039,N_9906,N_11356);
nor U15040 (N_15040,N_9709,N_10423);
nor U15041 (N_15041,N_12188,N_10674);
and U15042 (N_15042,N_11015,N_9456);
or U15043 (N_15043,N_10455,N_9705);
nand U15044 (N_15044,N_10019,N_9837);
nor U15045 (N_15045,N_11323,N_12322);
xnor U15046 (N_15046,N_9908,N_12379);
and U15047 (N_15047,N_12108,N_9740);
nor U15048 (N_15048,N_9580,N_11030);
and U15049 (N_15049,N_11726,N_11559);
xnor U15050 (N_15050,N_11862,N_12180);
nor U15051 (N_15051,N_9441,N_9901);
and U15052 (N_15052,N_12025,N_9781);
nor U15053 (N_15053,N_9672,N_11035);
xor U15054 (N_15054,N_10996,N_11815);
or U15055 (N_15055,N_10714,N_9476);
or U15056 (N_15056,N_11385,N_10840);
nor U15057 (N_15057,N_12068,N_11260);
nor U15058 (N_15058,N_10237,N_10641);
nand U15059 (N_15059,N_11349,N_10924);
or U15060 (N_15060,N_10098,N_11898);
or U15061 (N_15061,N_11944,N_10237);
nor U15062 (N_15062,N_9829,N_10553);
nor U15063 (N_15063,N_10298,N_10677);
or U15064 (N_15064,N_10507,N_10146);
and U15065 (N_15065,N_11177,N_10216);
nand U15066 (N_15066,N_9532,N_10378);
nand U15067 (N_15067,N_11083,N_11281);
xnor U15068 (N_15068,N_10466,N_11555);
nor U15069 (N_15069,N_11769,N_10995);
or U15070 (N_15070,N_11509,N_10179);
nor U15071 (N_15071,N_9736,N_11936);
nand U15072 (N_15072,N_9770,N_10077);
and U15073 (N_15073,N_9605,N_10224);
and U15074 (N_15074,N_10536,N_11009);
and U15075 (N_15075,N_10290,N_10084);
xnor U15076 (N_15076,N_11166,N_10992);
nand U15077 (N_15077,N_12299,N_10307);
xor U15078 (N_15078,N_9775,N_10105);
xor U15079 (N_15079,N_10919,N_12357);
nand U15080 (N_15080,N_12308,N_9814);
nand U15081 (N_15081,N_10272,N_10302);
and U15082 (N_15082,N_10147,N_9877);
nor U15083 (N_15083,N_12147,N_11235);
nor U15084 (N_15084,N_11027,N_11897);
xnor U15085 (N_15085,N_12338,N_10530);
nand U15086 (N_15086,N_12182,N_11862);
nand U15087 (N_15087,N_11285,N_12279);
nand U15088 (N_15088,N_11391,N_9377);
nor U15089 (N_15089,N_11913,N_10104);
nor U15090 (N_15090,N_11307,N_10149);
nand U15091 (N_15091,N_10335,N_11051);
or U15092 (N_15092,N_10785,N_12324);
nor U15093 (N_15093,N_9496,N_11808);
xor U15094 (N_15094,N_12279,N_12031);
xnor U15095 (N_15095,N_10875,N_10780);
or U15096 (N_15096,N_9737,N_12047);
xor U15097 (N_15097,N_9460,N_12169);
or U15098 (N_15098,N_10198,N_11729);
or U15099 (N_15099,N_10876,N_10038);
nand U15100 (N_15100,N_10577,N_10863);
and U15101 (N_15101,N_10483,N_11707);
xnor U15102 (N_15102,N_9444,N_11189);
and U15103 (N_15103,N_10655,N_10236);
nand U15104 (N_15104,N_9859,N_10918);
xor U15105 (N_15105,N_11651,N_10997);
and U15106 (N_15106,N_12220,N_11200);
xor U15107 (N_15107,N_11635,N_10304);
xnor U15108 (N_15108,N_10007,N_10633);
nor U15109 (N_15109,N_10350,N_11648);
or U15110 (N_15110,N_11424,N_11830);
and U15111 (N_15111,N_10499,N_10823);
nand U15112 (N_15112,N_10627,N_9938);
xnor U15113 (N_15113,N_10234,N_11865);
nand U15114 (N_15114,N_11230,N_10830);
or U15115 (N_15115,N_9829,N_12103);
or U15116 (N_15116,N_12280,N_9649);
nand U15117 (N_15117,N_10461,N_10665);
nor U15118 (N_15118,N_11168,N_9399);
xnor U15119 (N_15119,N_11911,N_12028);
or U15120 (N_15120,N_11840,N_11468);
xnor U15121 (N_15121,N_9848,N_12144);
xor U15122 (N_15122,N_12090,N_12066);
or U15123 (N_15123,N_9552,N_9452);
and U15124 (N_15124,N_9539,N_12164);
and U15125 (N_15125,N_10850,N_9927);
nand U15126 (N_15126,N_9670,N_10771);
and U15127 (N_15127,N_11359,N_12227);
nor U15128 (N_15128,N_9885,N_10411);
and U15129 (N_15129,N_11885,N_10428);
xnor U15130 (N_15130,N_9510,N_10251);
nand U15131 (N_15131,N_12056,N_12390);
nand U15132 (N_15132,N_9599,N_10203);
or U15133 (N_15133,N_10520,N_11389);
or U15134 (N_15134,N_9477,N_11795);
xor U15135 (N_15135,N_10725,N_12404);
and U15136 (N_15136,N_10660,N_9627);
xor U15137 (N_15137,N_10171,N_9905);
nand U15138 (N_15138,N_12473,N_10853);
xnor U15139 (N_15139,N_12345,N_11277);
xnor U15140 (N_15140,N_10603,N_10062);
or U15141 (N_15141,N_12348,N_10700);
or U15142 (N_15142,N_11528,N_11755);
nand U15143 (N_15143,N_10023,N_9408);
or U15144 (N_15144,N_9932,N_10489);
nand U15145 (N_15145,N_12455,N_9447);
or U15146 (N_15146,N_10449,N_12301);
nor U15147 (N_15147,N_9487,N_11400);
and U15148 (N_15148,N_12060,N_11797);
nor U15149 (N_15149,N_10721,N_11331);
or U15150 (N_15150,N_9842,N_10248);
xor U15151 (N_15151,N_11645,N_12429);
or U15152 (N_15152,N_10108,N_9899);
nor U15153 (N_15153,N_10596,N_10536);
nor U15154 (N_15154,N_10137,N_12114);
nand U15155 (N_15155,N_12328,N_10807);
xor U15156 (N_15156,N_10678,N_10591);
and U15157 (N_15157,N_11811,N_10630);
nand U15158 (N_15158,N_12096,N_10122);
nand U15159 (N_15159,N_10205,N_10601);
or U15160 (N_15160,N_10859,N_11963);
nor U15161 (N_15161,N_10829,N_10992);
nor U15162 (N_15162,N_10422,N_12330);
or U15163 (N_15163,N_11150,N_12201);
nand U15164 (N_15164,N_10170,N_9553);
or U15165 (N_15165,N_11855,N_9471);
nand U15166 (N_15166,N_11435,N_10572);
nand U15167 (N_15167,N_11484,N_11260);
and U15168 (N_15168,N_10906,N_11593);
or U15169 (N_15169,N_10233,N_9731);
and U15170 (N_15170,N_11538,N_12092);
nand U15171 (N_15171,N_11916,N_11018);
and U15172 (N_15172,N_10309,N_11853);
nand U15173 (N_15173,N_10377,N_11669);
or U15174 (N_15174,N_11205,N_11956);
xor U15175 (N_15175,N_11494,N_9694);
and U15176 (N_15176,N_12458,N_10430);
xnor U15177 (N_15177,N_12403,N_11382);
nor U15178 (N_15178,N_10641,N_11682);
xor U15179 (N_15179,N_12410,N_9535);
xor U15180 (N_15180,N_11447,N_9788);
and U15181 (N_15181,N_12066,N_9532);
nand U15182 (N_15182,N_11366,N_11454);
xnor U15183 (N_15183,N_11139,N_11932);
nor U15184 (N_15184,N_11650,N_9625);
and U15185 (N_15185,N_9539,N_10216);
nand U15186 (N_15186,N_10724,N_10783);
nor U15187 (N_15187,N_10719,N_12403);
nor U15188 (N_15188,N_11570,N_12469);
or U15189 (N_15189,N_11191,N_12332);
nor U15190 (N_15190,N_10577,N_10770);
nand U15191 (N_15191,N_12143,N_11436);
or U15192 (N_15192,N_11678,N_10867);
and U15193 (N_15193,N_11433,N_9419);
and U15194 (N_15194,N_9664,N_11929);
xnor U15195 (N_15195,N_11384,N_11432);
or U15196 (N_15196,N_11124,N_10040);
nor U15197 (N_15197,N_11266,N_11293);
or U15198 (N_15198,N_11858,N_11924);
xnor U15199 (N_15199,N_12485,N_11846);
nand U15200 (N_15200,N_9691,N_10512);
or U15201 (N_15201,N_11718,N_11724);
and U15202 (N_15202,N_11496,N_11555);
xnor U15203 (N_15203,N_9917,N_10809);
nor U15204 (N_15204,N_10163,N_11557);
xor U15205 (N_15205,N_11635,N_10669);
nand U15206 (N_15206,N_10915,N_11366);
or U15207 (N_15207,N_10119,N_9733);
nand U15208 (N_15208,N_10723,N_12215);
or U15209 (N_15209,N_10429,N_11337);
or U15210 (N_15210,N_9791,N_10166);
or U15211 (N_15211,N_11313,N_10790);
and U15212 (N_15212,N_10589,N_11051);
and U15213 (N_15213,N_9490,N_12400);
nand U15214 (N_15214,N_10998,N_11685);
xor U15215 (N_15215,N_11241,N_11035);
or U15216 (N_15216,N_11865,N_10690);
xor U15217 (N_15217,N_10637,N_12242);
xor U15218 (N_15218,N_10102,N_10230);
xnor U15219 (N_15219,N_11126,N_12451);
xor U15220 (N_15220,N_10307,N_11377);
xnor U15221 (N_15221,N_10437,N_12233);
or U15222 (N_15222,N_10079,N_10911);
xor U15223 (N_15223,N_11779,N_9728);
nand U15224 (N_15224,N_10812,N_11089);
nor U15225 (N_15225,N_11856,N_11570);
nor U15226 (N_15226,N_12341,N_9581);
and U15227 (N_15227,N_10480,N_12064);
xnor U15228 (N_15228,N_11550,N_11402);
or U15229 (N_15229,N_9995,N_9788);
xnor U15230 (N_15230,N_10320,N_12210);
or U15231 (N_15231,N_11691,N_10437);
or U15232 (N_15232,N_10833,N_9520);
nand U15233 (N_15233,N_10364,N_12298);
nor U15234 (N_15234,N_10634,N_11169);
or U15235 (N_15235,N_12142,N_12175);
xnor U15236 (N_15236,N_11950,N_10376);
xor U15237 (N_15237,N_12433,N_10725);
nor U15238 (N_15238,N_9415,N_11608);
xnor U15239 (N_15239,N_11828,N_11276);
and U15240 (N_15240,N_11810,N_11178);
and U15241 (N_15241,N_11188,N_9835);
and U15242 (N_15242,N_11918,N_10267);
and U15243 (N_15243,N_9404,N_10496);
and U15244 (N_15244,N_11758,N_10288);
or U15245 (N_15245,N_10759,N_10542);
or U15246 (N_15246,N_10447,N_10187);
nor U15247 (N_15247,N_11476,N_11533);
nor U15248 (N_15248,N_10062,N_9829);
nor U15249 (N_15249,N_9697,N_11541);
xor U15250 (N_15250,N_12351,N_10127);
and U15251 (N_15251,N_10436,N_10528);
and U15252 (N_15252,N_9567,N_11602);
xor U15253 (N_15253,N_10662,N_11113);
or U15254 (N_15254,N_9778,N_11124);
and U15255 (N_15255,N_9439,N_9937);
or U15256 (N_15256,N_9910,N_11048);
and U15257 (N_15257,N_10371,N_10985);
or U15258 (N_15258,N_9555,N_12409);
xor U15259 (N_15259,N_9756,N_9910);
xor U15260 (N_15260,N_11429,N_12450);
and U15261 (N_15261,N_9854,N_10119);
or U15262 (N_15262,N_9420,N_10079);
nand U15263 (N_15263,N_11987,N_9657);
nand U15264 (N_15264,N_12160,N_9479);
nor U15265 (N_15265,N_12243,N_12417);
nand U15266 (N_15266,N_9614,N_11581);
xor U15267 (N_15267,N_11128,N_11820);
or U15268 (N_15268,N_9480,N_9655);
or U15269 (N_15269,N_11597,N_11260);
and U15270 (N_15270,N_11840,N_11143);
nor U15271 (N_15271,N_10601,N_12160);
or U15272 (N_15272,N_12358,N_11378);
nand U15273 (N_15273,N_10286,N_9422);
nand U15274 (N_15274,N_9898,N_12052);
xnor U15275 (N_15275,N_12051,N_10053);
and U15276 (N_15276,N_11378,N_12072);
and U15277 (N_15277,N_12427,N_12049);
xor U15278 (N_15278,N_11289,N_10071);
and U15279 (N_15279,N_10991,N_9483);
and U15280 (N_15280,N_12377,N_11282);
nor U15281 (N_15281,N_11512,N_10530);
or U15282 (N_15282,N_11042,N_12274);
xor U15283 (N_15283,N_9701,N_12291);
nand U15284 (N_15284,N_12264,N_10107);
and U15285 (N_15285,N_11607,N_10587);
xnor U15286 (N_15286,N_9863,N_11054);
nor U15287 (N_15287,N_10218,N_9556);
nor U15288 (N_15288,N_9532,N_11251);
nor U15289 (N_15289,N_11985,N_9803);
or U15290 (N_15290,N_10871,N_9941);
nor U15291 (N_15291,N_10277,N_12152);
xnor U15292 (N_15292,N_9529,N_10372);
nor U15293 (N_15293,N_9686,N_11978);
xnor U15294 (N_15294,N_10773,N_11705);
nand U15295 (N_15295,N_9467,N_10844);
or U15296 (N_15296,N_11376,N_10887);
nor U15297 (N_15297,N_12306,N_11827);
nand U15298 (N_15298,N_10435,N_11425);
and U15299 (N_15299,N_10134,N_9809);
nand U15300 (N_15300,N_9852,N_9690);
xor U15301 (N_15301,N_10642,N_11469);
xnor U15302 (N_15302,N_12016,N_11797);
nor U15303 (N_15303,N_12062,N_10457);
or U15304 (N_15304,N_10495,N_11607);
nor U15305 (N_15305,N_10760,N_10379);
xor U15306 (N_15306,N_12330,N_10688);
xnor U15307 (N_15307,N_12091,N_11014);
nor U15308 (N_15308,N_9854,N_11869);
nor U15309 (N_15309,N_12358,N_10474);
xor U15310 (N_15310,N_11357,N_12462);
nor U15311 (N_15311,N_12174,N_9947);
xnor U15312 (N_15312,N_12347,N_10192);
or U15313 (N_15313,N_10825,N_10852);
xor U15314 (N_15314,N_10228,N_10892);
nor U15315 (N_15315,N_12018,N_9735);
nor U15316 (N_15316,N_12370,N_12296);
nand U15317 (N_15317,N_12486,N_9637);
and U15318 (N_15318,N_10210,N_9657);
xor U15319 (N_15319,N_9918,N_12136);
or U15320 (N_15320,N_11488,N_12031);
nand U15321 (N_15321,N_9914,N_10156);
or U15322 (N_15322,N_9479,N_11996);
nor U15323 (N_15323,N_11998,N_11952);
and U15324 (N_15324,N_11212,N_9531);
or U15325 (N_15325,N_10310,N_12315);
nor U15326 (N_15326,N_11563,N_12326);
nor U15327 (N_15327,N_9768,N_9848);
xor U15328 (N_15328,N_10795,N_10322);
and U15329 (N_15329,N_12120,N_11076);
nand U15330 (N_15330,N_10464,N_10538);
nand U15331 (N_15331,N_9607,N_11946);
and U15332 (N_15332,N_10276,N_12301);
nor U15333 (N_15333,N_11718,N_11703);
nor U15334 (N_15334,N_11971,N_9927);
xor U15335 (N_15335,N_9443,N_9600);
xor U15336 (N_15336,N_9831,N_10059);
nand U15337 (N_15337,N_11218,N_11578);
and U15338 (N_15338,N_11170,N_10188);
xnor U15339 (N_15339,N_12399,N_10127);
nor U15340 (N_15340,N_9517,N_12090);
and U15341 (N_15341,N_11254,N_12404);
xor U15342 (N_15342,N_11272,N_11554);
nor U15343 (N_15343,N_9378,N_11346);
nand U15344 (N_15344,N_10102,N_10353);
xor U15345 (N_15345,N_10853,N_9914);
xnor U15346 (N_15346,N_10156,N_10377);
nor U15347 (N_15347,N_12125,N_11238);
or U15348 (N_15348,N_10082,N_10553);
xnor U15349 (N_15349,N_10857,N_11296);
xnor U15350 (N_15350,N_10317,N_10746);
or U15351 (N_15351,N_11394,N_10725);
nor U15352 (N_15352,N_9926,N_9605);
nor U15353 (N_15353,N_10567,N_9804);
nand U15354 (N_15354,N_11090,N_12269);
nor U15355 (N_15355,N_11278,N_9820);
xor U15356 (N_15356,N_9789,N_11873);
xor U15357 (N_15357,N_10213,N_11794);
nand U15358 (N_15358,N_9778,N_12361);
and U15359 (N_15359,N_11566,N_10585);
xnor U15360 (N_15360,N_9735,N_11670);
and U15361 (N_15361,N_11185,N_10433);
nand U15362 (N_15362,N_10902,N_10537);
nand U15363 (N_15363,N_11761,N_11459);
xor U15364 (N_15364,N_11189,N_11229);
xor U15365 (N_15365,N_11209,N_10833);
xor U15366 (N_15366,N_11591,N_11149);
and U15367 (N_15367,N_11108,N_11532);
and U15368 (N_15368,N_10949,N_11421);
nor U15369 (N_15369,N_9841,N_11130);
nor U15370 (N_15370,N_11085,N_10666);
or U15371 (N_15371,N_10281,N_10939);
xnor U15372 (N_15372,N_12286,N_11018);
xor U15373 (N_15373,N_11006,N_11698);
nor U15374 (N_15374,N_10892,N_10316);
nand U15375 (N_15375,N_11786,N_10455);
and U15376 (N_15376,N_9458,N_12038);
nor U15377 (N_15377,N_10234,N_11801);
and U15378 (N_15378,N_10950,N_9566);
or U15379 (N_15379,N_10586,N_12003);
xor U15380 (N_15380,N_10395,N_9501);
nor U15381 (N_15381,N_9637,N_12145);
or U15382 (N_15382,N_11406,N_11899);
xor U15383 (N_15383,N_10331,N_11008);
and U15384 (N_15384,N_12232,N_11434);
nand U15385 (N_15385,N_11256,N_10996);
xnor U15386 (N_15386,N_11849,N_11012);
nand U15387 (N_15387,N_9439,N_12484);
xnor U15388 (N_15388,N_12232,N_12154);
xnor U15389 (N_15389,N_9422,N_11978);
nor U15390 (N_15390,N_11959,N_10310);
nor U15391 (N_15391,N_10844,N_12245);
or U15392 (N_15392,N_9792,N_10282);
nor U15393 (N_15393,N_11860,N_12130);
nand U15394 (N_15394,N_11934,N_10897);
and U15395 (N_15395,N_10478,N_9540);
nor U15396 (N_15396,N_12035,N_10473);
and U15397 (N_15397,N_11145,N_10553);
xnor U15398 (N_15398,N_9697,N_12311);
and U15399 (N_15399,N_10408,N_9680);
nand U15400 (N_15400,N_12479,N_9877);
xnor U15401 (N_15401,N_10789,N_12399);
xor U15402 (N_15402,N_11142,N_9852);
or U15403 (N_15403,N_10244,N_11711);
xnor U15404 (N_15404,N_12371,N_11777);
or U15405 (N_15405,N_11324,N_11741);
or U15406 (N_15406,N_9424,N_9592);
xor U15407 (N_15407,N_11845,N_9665);
xnor U15408 (N_15408,N_9866,N_10213);
nand U15409 (N_15409,N_11444,N_12112);
nor U15410 (N_15410,N_10717,N_12456);
nand U15411 (N_15411,N_9961,N_11356);
nor U15412 (N_15412,N_11941,N_12032);
or U15413 (N_15413,N_11686,N_12205);
nor U15414 (N_15414,N_11154,N_11426);
xnor U15415 (N_15415,N_11408,N_12455);
nand U15416 (N_15416,N_9381,N_12171);
nor U15417 (N_15417,N_11716,N_11072);
and U15418 (N_15418,N_10583,N_12457);
xor U15419 (N_15419,N_11720,N_11473);
nor U15420 (N_15420,N_11652,N_12380);
xnor U15421 (N_15421,N_11864,N_11401);
and U15422 (N_15422,N_10211,N_12274);
nor U15423 (N_15423,N_9686,N_10653);
or U15424 (N_15424,N_12447,N_9393);
nor U15425 (N_15425,N_10699,N_9598);
nor U15426 (N_15426,N_9882,N_12362);
xnor U15427 (N_15427,N_12186,N_10279);
xor U15428 (N_15428,N_12184,N_11869);
xor U15429 (N_15429,N_11082,N_11151);
nand U15430 (N_15430,N_9944,N_10716);
xor U15431 (N_15431,N_10225,N_11955);
and U15432 (N_15432,N_12031,N_11026);
xor U15433 (N_15433,N_12164,N_10433);
or U15434 (N_15434,N_12338,N_9637);
nand U15435 (N_15435,N_10528,N_10562);
nand U15436 (N_15436,N_11290,N_11517);
or U15437 (N_15437,N_11531,N_12275);
or U15438 (N_15438,N_11177,N_9432);
nor U15439 (N_15439,N_12446,N_11334);
or U15440 (N_15440,N_9933,N_10268);
and U15441 (N_15441,N_10480,N_11485);
xor U15442 (N_15442,N_10399,N_9503);
nand U15443 (N_15443,N_11135,N_12187);
and U15444 (N_15444,N_10414,N_10641);
nand U15445 (N_15445,N_10266,N_12486);
or U15446 (N_15446,N_9527,N_9453);
and U15447 (N_15447,N_9589,N_9410);
nor U15448 (N_15448,N_12422,N_10645);
nand U15449 (N_15449,N_12225,N_10405);
nor U15450 (N_15450,N_11158,N_12003);
nand U15451 (N_15451,N_10639,N_9466);
xnor U15452 (N_15452,N_10852,N_12289);
nand U15453 (N_15453,N_9754,N_10569);
xnor U15454 (N_15454,N_11501,N_9838);
xnor U15455 (N_15455,N_12264,N_9498);
nand U15456 (N_15456,N_9695,N_9980);
xor U15457 (N_15457,N_11069,N_12227);
nor U15458 (N_15458,N_10954,N_11844);
xor U15459 (N_15459,N_10646,N_10592);
nor U15460 (N_15460,N_10058,N_9534);
nand U15461 (N_15461,N_9810,N_10281);
or U15462 (N_15462,N_12047,N_12442);
nor U15463 (N_15463,N_11960,N_10487);
xor U15464 (N_15464,N_12312,N_12196);
or U15465 (N_15465,N_9764,N_10962);
or U15466 (N_15466,N_11458,N_9606);
nor U15467 (N_15467,N_11865,N_10462);
xor U15468 (N_15468,N_10417,N_9997);
xor U15469 (N_15469,N_11613,N_10049);
or U15470 (N_15470,N_9747,N_10673);
or U15471 (N_15471,N_9702,N_12475);
nand U15472 (N_15472,N_10045,N_12059);
nand U15473 (N_15473,N_10198,N_12380);
nor U15474 (N_15474,N_9407,N_12141);
and U15475 (N_15475,N_11391,N_10226);
nor U15476 (N_15476,N_11841,N_11292);
nand U15477 (N_15477,N_10113,N_10559);
and U15478 (N_15478,N_11201,N_9618);
nor U15479 (N_15479,N_9965,N_11010);
and U15480 (N_15480,N_9404,N_10018);
nor U15481 (N_15481,N_9751,N_11835);
or U15482 (N_15482,N_10698,N_11185);
and U15483 (N_15483,N_11748,N_11971);
or U15484 (N_15484,N_9624,N_9854);
nand U15485 (N_15485,N_12327,N_11914);
nor U15486 (N_15486,N_12304,N_9510);
nor U15487 (N_15487,N_9483,N_9467);
nand U15488 (N_15488,N_12495,N_11565);
nor U15489 (N_15489,N_12376,N_11341);
nand U15490 (N_15490,N_9987,N_9712);
and U15491 (N_15491,N_11729,N_11100);
or U15492 (N_15492,N_9760,N_10457);
nand U15493 (N_15493,N_10869,N_12323);
or U15494 (N_15494,N_10645,N_12476);
xnor U15495 (N_15495,N_11336,N_9538);
and U15496 (N_15496,N_10037,N_11435);
nor U15497 (N_15497,N_10730,N_12346);
nand U15498 (N_15498,N_11494,N_12165);
nor U15499 (N_15499,N_9789,N_11121);
nand U15500 (N_15500,N_11574,N_10271);
or U15501 (N_15501,N_12498,N_12031);
or U15502 (N_15502,N_10213,N_12141);
nand U15503 (N_15503,N_10561,N_9652);
nor U15504 (N_15504,N_11565,N_12223);
or U15505 (N_15505,N_9869,N_9866);
nand U15506 (N_15506,N_12137,N_11494);
and U15507 (N_15507,N_11671,N_9720);
xor U15508 (N_15508,N_10711,N_9586);
xnor U15509 (N_15509,N_12290,N_9524);
and U15510 (N_15510,N_11054,N_11578);
and U15511 (N_15511,N_12009,N_10607);
nor U15512 (N_15512,N_10738,N_10392);
or U15513 (N_15513,N_10241,N_10339);
xor U15514 (N_15514,N_10040,N_11633);
xor U15515 (N_15515,N_9736,N_10071);
or U15516 (N_15516,N_10602,N_11046);
and U15517 (N_15517,N_10532,N_11409);
and U15518 (N_15518,N_10594,N_12318);
xor U15519 (N_15519,N_10475,N_9562);
or U15520 (N_15520,N_9709,N_12021);
nand U15521 (N_15521,N_10098,N_12457);
and U15522 (N_15522,N_11394,N_11593);
xor U15523 (N_15523,N_10817,N_9552);
nand U15524 (N_15524,N_10153,N_11669);
xor U15525 (N_15525,N_11992,N_9903);
or U15526 (N_15526,N_9597,N_10665);
nor U15527 (N_15527,N_11075,N_10155);
and U15528 (N_15528,N_9432,N_10351);
and U15529 (N_15529,N_11098,N_10018);
nand U15530 (N_15530,N_10375,N_12198);
nand U15531 (N_15531,N_10677,N_12054);
nor U15532 (N_15532,N_12317,N_11528);
xor U15533 (N_15533,N_11189,N_9979);
nor U15534 (N_15534,N_9376,N_12243);
nand U15535 (N_15535,N_11838,N_11527);
or U15536 (N_15536,N_12303,N_9730);
and U15537 (N_15537,N_9404,N_9566);
and U15538 (N_15538,N_9418,N_12158);
or U15539 (N_15539,N_9835,N_12036);
and U15540 (N_15540,N_11219,N_12231);
and U15541 (N_15541,N_10977,N_11103);
nand U15542 (N_15542,N_9746,N_12150);
nand U15543 (N_15543,N_9426,N_9753);
and U15544 (N_15544,N_12033,N_11577);
nand U15545 (N_15545,N_10934,N_10599);
and U15546 (N_15546,N_10754,N_12088);
and U15547 (N_15547,N_9979,N_10255);
nand U15548 (N_15548,N_9456,N_9924);
or U15549 (N_15549,N_11431,N_9427);
or U15550 (N_15550,N_10463,N_11928);
and U15551 (N_15551,N_10738,N_10498);
xor U15552 (N_15552,N_9892,N_10176);
or U15553 (N_15553,N_10134,N_9463);
nand U15554 (N_15554,N_9747,N_9931);
nor U15555 (N_15555,N_12139,N_10905);
nor U15556 (N_15556,N_10624,N_10050);
and U15557 (N_15557,N_11617,N_11832);
nand U15558 (N_15558,N_10151,N_12021);
nand U15559 (N_15559,N_12490,N_9425);
xor U15560 (N_15560,N_9687,N_10920);
nor U15561 (N_15561,N_12395,N_11713);
xnor U15562 (N_15562,N_10116,N_10354);
xor U15563 (N_15563,N_10545,N_11353);
or U15564 (N_15564,N_11818,N_10018);
xor U15565 (N_15565,N_12487,N_10331);
and U15566 (N_15566,N_10017,N_10580);
and U15567 (N_15567,N_10030,N_10447);
and U15568 (N_15568,N_9870,N_11001);
and U15569 (N_15569,N_12021,N_9910);
xnor U15570 (N_15570,N_10226,N_9805);
xor U15571 (N_15571,N_10380,N_11591);
nand U15572 (N_15572,N_12163,N_11368);
nor U15573 (N_15573,N_12111,N_11779);
nor U15574 (N_15574,N_12423,N_11448);
and U15575 (N_15575,N_9544,N_9414);
nand U15576 (N_15576,N_11010,N_9638);
and U15577 (N_15577,N_12029,N_11701);
and U15578 (N_15578,N_11089,N_11482);
nor U15579 (N_15579,N_9539,N_10827);
nor U15580 (N_15580,N_11930,N_10499);
or U15581 (N_15581,N_11242,N_12362);
nor U15582 (N_15582,N_12033,N_9643);
and U15583 (N_15583,N_12019,N_12366);
or U15584 (N_15584,N_10100,N_10101);
or U15585 (N_15585,N_9724,N_9933);
xnor U15586 (N_15586,N_9553,N_10351);
nand U15587 (N_15587,N_9686,N_9679);
xor U15588 (N_15588,N_10425,N_12156);
xnor U15589 (N_15589,N_11151,N_11902);
xor U15590 (N_15590,N_10311,N_11467);
xnor U15591 (N_15591,N_10513,N_10558);
nand U15592 (N_15592,N_9625,N_11612);
or U15593 (N_15593,N_10129,N_11283);
nand U15594 (N_15594,N_9508,N_11556);
or U15595 (N_15595,N_11927,N_9963);
or U15596 (N_15596,N_10068,N_11086);
nand U15597 (N_15597,N_12117,N_11094);
nand U15598 (N_15598,N_10818,N_11822);
or U15599 (N_15599,N_12061,N_10304);
xnor U15600 (N_15600,N_11358,N_11203);
or U15601 (N_15601,N_9588,N_11384);
xnor U15602 (N_15602,N_12276,N_11546);
nor U15603 (N_15603,N_11653,N_12428);
or U15604 (N_15604,N_11479,N_9702);
and U15605 (N_15605,N_12121,N_9540);
and U15606 (N_15606,N_10446,N_9586);
nand U15607 (N_15607,N_9734,N_9446);
nand U15608 (N_15608,N_10239,N_11061);
nor U15609 (N_15609,N_9744,N_11455);
or U15610 (N_15610,N_10704,N_11391);
xnor U15611 (N_15611,N_10253,N_9580);
xnor U15612 (N_15612,N_11433,N_10879);
nor U15613 (N_15613,N_11955,N_11166);
or U15614 (N_15614,N_9798,N_10642);
and U15615 (N_15615,N_12451,N_12400);
and U15616 (N_15616,N_11074,N_10700);
nor U15617 (N_15617,N_10021,N_9399);
or U15618 (N_15618,N_11444,N_10527);
nor U15619 (N_15619,N_11723,N_12343);
xnor U15620 (N_15620,N_11347,N_12054);
and U15621 (N_15621,N_10948,N_9895);
nor U15622 (N_15622,N_12144,N_10527);
or U15623 (N_15623,N_11005,N_11768);
nand U15624 (N_15624,N_10767,N_11779);
nand U15625 (N_15625,N_14408,N_15238);
nand U15626 (N_15626,N_14194,N_12929);
and U15627 (N_15627,N_12547,N_13760);
and U15628 (N_15628,N_14288,N_14210);
or U15629 (N_15629,N_12764,N_12718);
or U15630 (N_15630,N_14416,N_15278);
nor U15631 (N_15631,N_13077,N_14629);
nor U15632 (N_15632,N_15540,N_14640);
or U15633 (N_15633,N_15539,N_15242);
nand U15634 (N_15634,N_13218,N_14552);
nor U15635 (N_15635,N_13086,N_14948);
nand U15636 (N_15636,N_15223,N_15180);
nor U15637 (N_15637,N_13147,N_13192);
nand U15638 (N_15638,N_13657,N_13102);
and U15639 (N_15639,N_13775,N_14699);
or U15640 (N_15640,N_14915,N_14690);
xor U15641 (N_15641,N_15460,N_15397);
or U15642 (N_15642,N_13071,N_15040);
nor U15643 (N_15643,N_14113,N_14365);
nand U15644 (N_15644,N_14589,N_13438);
nand U15645 (N_15645,N_14145,N_13090);
or U15646 (N_15646,N_14134,N_14614);
and U15647 (N_15647,N_13982,N_14587);
or U15648 (N_15648,N_13095,N_14601);
and U15649 (N_15649,N_13936,N_12670);
and U15650 (N_15650,N_15500,N_13836);
xor U15651 (N_15651,N_12696,N_12559);
xnor U15652 (N_15652,N_12549,N_14506);
nor U15653 (N_15653,N_13774,N_14532);
or U15654 (N_15654,N_14485,N_12554);
nor U15655 (N_15655,N_15232,N_14004);
and U15656 (N_15656,N_12912,N_13377);
or U15657 (N_15657,N_15075,N_14637);
and U15658 (N_15658,N_13143,N_15128);
and U15659 (N_15659,N_12780,N_13296);
nor U15660 (N_15660,N_12980,N_14765);
nor U15661 (N_15661,N_15410,N_15213);
and U15662 (N_15662,N_12822,N_14177);
xor U15663 (N_15663,N_14292,N_15623);
nand U15664 (N_15664,N_15588,N_14569);
xor U15665 (N_15665,N_14498,N_13957);
or U15666 (N_15666,N_13313,N_12686);
xor U15667 (N_15667,N_15022,N_13809);
nand U15668 (N_15668,N_15271,N_15217);
or U15669 (N_15669,N_14588,N_14738);
and U15670 (N_15670,N_12689,N_13683);
nand U15671 (N_15671,N_14716,N_14800);
or U15672 (N_15672,N_15027,N_13883);
and U15673 (N_15673,N_13257,N_13167);
xor U15674 (N_15674,N_14493,N_14153);
xnor U15675 (N_15675,N_13796,N_15338);
and U15676 (N_15676,N_14985,N_15381);
nand U15677 (N_15677,N_13433,N_15455);
or U15678 (N_15678,N_14154,N_12662);
xnor U15679 (N_15679,N_12934,N_12707);
or U15680 (N_15680,N_14271,N_14734);
and U15681 (N_15681,N_15331,N_12719);
and U15682 (N_15682,N_12658,N_12527);
xnor U15683 (N_15683,N_13491,N_14127);
nor U15684 (N_15684,N_13868,N_13819);
nand U15685 (N_15685,N_13104,N_14516);
or U15686 (N_15686,N_12902,N_13069);
and U15687 (N_15687,N_13097,N_13413);
nand U15688 (N_15688,N_14576,N_15045);
nand U15689 (N_15689,N_12983,N_13004);
nand U15690 (N_15690,N_14471,N_15544);
xnor U15691 (N_15691,N_14624,N_15442);
nor U15692 (N_15692,N_12959,N_13894);
or U15693 (N_15693,N_13552,N_14842);
and U15694 (N_15694,N_14306,N_14163);
and U15695 (N_15695,N_14970,N_14804);
xnor U15696 (N_15696,N_13101,N_13988);
nand U15697 (N_15697,N_14266,N_14044);
and U15698 (N_15698,N_15082,N_14360);
and U15699 (N_15699,N_15193,N_13272);
or U15700 (N_15700,N_13470,N_13591);
and U15701 (N_15701,N_14902,N_14321);
or U15702 (N_15702,N_15345,N_14853);
and U15703 (N_15703,N_13050,N_12898);
nand U15704 (N_15704,N_14940,N_12779);
nor U15705 (N_15705,N_13509,N_13314);
or U15706 (N_15706,N_14421,N_14062);
xnor U15707 (N_15707,N_14592,N_15302);
or U15708 (N_15708,N_13790,N_14191);
nor U15709 (N_15709,N_12743,N_14870);
nand U15710 (N_15710,N_15587,N_13535);
and U15711 (N_15711,N_13892,N_14770);
nor U15712 (N_15712,N_13932,N_15101);
and U15713 (N_15713,N_14814,N_12885);
nand U15714 (N_15714,N_15535,N_15608);
and U15715 (N_15715,N_14504,N_14726);
or U15716 (N_15716,N_14079,N_14967);
xnor U15717 (N_15717,N_14147,N_12888);
nor U15718 (N_15718,N_12704,N_12682);
and U15719 (N_15719,N_13083,N_14984);
xnor U15720 (N_15720,N_14497,N_14295);
xnor U15721 (N_15721,N_12678,N_14168);
and U15722 (N_15722,N_14730,N_12768);
nor U15723 (N_15723,N_12500,N_13288);
and U15724 (N_15724,N_13079,N_14833);
nor U15725 (N_15725,N_13975,N_12796);
and U15726 (N_15726,N_13755,N_14742);
or U15727 (N_15727,N_15194,N_13389);
xnor U15728 (N_15728,N_14867,N_12951);
nor U15729 (N_15729,N_15253,N_12544);
or U15730 (N_15730,N_14054,N_15077);
xor U15731 (N_15731,N_14415,N_12785);
nand U15732 (N_15732,N_12803,N_14381);
and U15733 (N_15733,N_13538,N_13772);
nand U15734 (N_15734,N_12633,N_12841);
xor U15735 (N_15735,N_13539,N_15118);
and U15736 (N_15736,N_14761,N_14012);
nor U15737 (N_15737,N_14228,N_14863);
nand U15738 (N_15738,N_13447,N_13091);
and U15739 (N_15739,N_12680,N_13204);
xor U15740 (N_15740,N_13264,N_13831);
nand U15741 (N_15741,N_12711,N_13939);
xor U15742 (N_15742,N_12932,N_13494);
nor U15743 (N_15743,N_14141,N_14227);
nor U15744 (N_15744,N_14521,N_13019);
nor U15745 (N_15745,N_12714,N_15435);
nor U15746 (N_15746,N_13574,N_15255);
and U15747 (N_15747,N_14192,N_12879);
xnor U15748 (N_15748,N_13888,N_14911);
nand U15749 (N_15749,N_15208,N_15273);
xnor U15750 (N_15750,N_13034,N_15571);
xor U15751 (N_15751,N_12660,N_13958);
nand U15752 (N_15752,N_13385,N_15536);
xor U15753 (N_15753,N_14159,N_13265);
xnor U15754 (N_15754,N_14565,N_15138);
nor U15755 (N_15755,N_13219,N_13979);
nor U15756 (N_15756,N_14267,N_13795);
or U15757 (N_15757,N_14435,N_14423);
nor U15758 (N_15758,N_15497,N_14320);
nor U15759 (N_15759,N_14489,N_14884);
and U15760 (N_15760,N_15337,N_14274);
nand U15761 (N_15761,N_15252,N_13676);
or U15762 (N_15762,N_13542,N_12863);
xnor U15763 (N_15763,N_15034,N_13611);
xor U15764 (N_15764,N_14420,N_12757);
xnor U15765 (N_15765,N_12823,N_15579);
and U15766 (N_15766,N_12792,N_12608);
nor U15767 (N_15767,N_14546,N_14083);
or U15768 (N_15768,N_13467,N_14347);
nor U15769 (N_15769,N_14344,N_14965);
nand U15770 (N_15770,N_13905,N_12669);
xnor U15771 (N_15771,N_13697,N_13812);
and U15772 (N_15772,N_13808,N_14816);
nor U15773 (N_15773,N_15141,N_14829);
or U15774 (N_15774,N_14590,N_13189);
xor U15775 (N_15775,N_14836,N_13827);
and U15776 (N_15776,N_13837,N_12816);
xnor U15777 (N_15777,N_14541,N_14304);
nand U15778 (N_15778,N_15339,N_15062);
and U15779 (N_15779,N_13974,N_15283);
nand U15780 (N_15780,N_13287,N_12521);
and U15781 (N_15781,N_15009,N_14317);
and U15782 (N_15782,N_13210,N_13155);
and U15783 (N_15783,N_13881,N_12926);
and U15784 (N_15784,N_14411,N_14830);
or U15785 (N_15785,N_13785,N_14865);
and U15786 (N_15786,N_13127,N_13263);
or U15787 (N_15787,N_13021,N_15327);
or U15788 (N_15788,N_13465,N_13511);
xor U15789 (N_15789,N_14939,N_14710);
or U15790 (N_15790,N_14468,N_15069);
nand U15791 (N_15791,N_14400,N_13153);
and U15792 (N_15792,N_15063,N_15306);
or U15793 (N_15793,N_15490,N_14956);
or U15794 (N_15794,N_13064,N_13724);
nand U15795 (N_15795,N_15513,N_13858);
and U15796 (N_15796,N_14473,N_14069);
or U15797 (N_15797,N_15143,N_15079);
nand U15798 (N_15798,N_13334,N_13586);
nor U15799 (N_15799,N_15085,N_13184);
and U15800 (N_15800,N_13158,N_13233);
xor U15801 (N_15801,N_13451,N_14050);
nor U15802 (N_15802,N_13955,N_13931);
or U15803 (N_15803,N_13556,N_13874);
xor U15804 (N_15804,N_14034,N_14018);
or U15805 (N_15805,N_13637,N_14312);
xor U15806 (N_15806,N_14989,N_14561);
nor U15807 (N_15807,N_13782,N_15043);
xor U15808 (N_15808,N_12784,N_14483);
or U15809 (N_15809,N_14839,N_13066);
xor U15810 (N_15810,N_14622,N_12817);
xnor U15811 (N_15811,N_14449,N_13386);
xnor U15812 (N_15812,N_14551,N_14136);
nor U15813 (N_15813,N_14263,N_14701);
or U15814 (N_15814,N_14739,N_14394);
nor U15815 (N_15815,N_13661,N_14037);
or U15816 (N_15816,N_14005,N_14443);
xor U15817 (N_15817,N_13185,N_13146);
nand U15818 (N_15818,N_12690,N_12966);
xor U15819 (N_15819,N_13216,N_14242);
nor U15820 (N_15820,N_14262,N_14482);
or U15821 (N_15821,N_15323,N_15239);
or U15822 (N_15822,N_13047,N_12578);
or U15823 (N_15823,N_14847,N_15542);
xor U15824 (N_15824,N_14611,N_12679);
xnor U15825 (N_15825,N_13387,N_14375);
xnor U15826 (N_15826,N_12519,N_13853);
xnor U15827 (N_15827,N_12828,N_14427);
and U15828 (N_15828,N_15474,N_13113);
nor U15829 (N_15829,N_14111,N_14619);
or U15830 (N_15830,N_15491,N_14457);
nor U15831 (N_15831,N_15090,N_12742);
or U15832 (N_15832,N_14605,N_13654);
and U15833 (N_15833,N_15452,N_12575);
and U15834 (N_15834,N_14882,N_14533);
and U15835 (N_15835,N_15350,N_14883);
nor U15836 (N_15836,N_15117,N_12988);
nand U15837 (N_15837,N_12835,N_12505);
xnor U15838 (N_15838,N_14960,N_15219);
xor U15839 (N_15839,N_13407,N_12552);
nand U15840 (N_15840,N_15624,N_13706);
nor U15841 (N_15841,N_12514,N_14469);
or U15842 (N_15842,N_14142,N_14821);
and U15843 (N_15843,N_14923,N_15523);
nor U15844 (N_15844,N_13701,N_15550);
or U15845 (N_15845,N_14291,N_14796);
nand U15846 (N_15846,N_15095,N_13609);
nand U15847 (N_15847,N_14221,N_14968);
and U15848 (N_15848,N_14664,N_13350);
and U15849 (N_15849,N_13440,N_12981);
xor U15850 (N_15850,N_13597,N_15249);
nor U15851 (N_15851,N_14934,N_15318);
nor U15852 (N_15852,N_12591,N_13846);
xor U15853 (N_15853,N_13890,N_15394);
xnor U15854 (N_15854,N_15458,N_14009);
or U15855 (N_15855,N_13716,N_14244);
nand U15856 (N_15856,N_13373,N_15260);
and U15857 (N_15857,N_14746,N_14299);
and U15858 (N_15858,N_14980,N_14852);
or U15859 (N_15859,N_14966,N_13945);
xnor U15860 (N_15860,N_13012,N_13545);
or U15861 (N_15861,N_13128,N_14452);
nor U15862 (N_15862,N_12917,N_12513);
xor U15863 (N_15863,N_13285,N_14309);
nand U15864 (N_15864,N_12586,N_15241);
xor U15865 (N_15865,N_13321,N_13032);
or U15866 (N_15866,N_14580,N_13277);
xnor U15867 (N_15867,N_12761,N_14214);
nor U15868 (N_15868,N_12577,N_13567);
xor U15869 (N_15869,N_14799,N_12830);
nand U15870 (N_15870,N_14338,N_12756);
nor U15871 (N_15871,N_12977,N_15604);
nor U15872 (N_15872,N_13388,N_15356);
or U15873 (N_15873,N_15307,N_13948);
and U15874 (N_15874,N_15083,N_13307);
xnor U15875 (N_15875,N_13633,N_15231);
nor U15876 (N_15876,N_14217,N_14310);
xnor U15877 (N_15877,N_12772,N_15052);
xnor U15878 (N_15878,N_15177,N_14876);
nand U15879 (N_15879,N_13000,N_15284);
or U15880 (N_15880,N_14208,N_12727);
xnor U15881 (N_15881,N_14524,N_13481);
or U15882 (N_15882,N_13170,N_13860);
nor U15883 (N_15883,N_14771,N_13767);
or U15884 (N_15884,N_15317,N_12890);
xor U15885 (N_15885,N_15501,N_15261);
nor U15886 (N_15886,N_13540,N_15355);
nand U15887 (N_15887,N_14155,N_13698);
nor U15888 (N_15888,N_14950,N_15372);
xor U15889 (N_15889,N_15233,N_14308);
nor U15890 (N_15890,N_13286,N_14118);
nand U15891 (N_15891,N_13190,N_14526);
and U15892 (N_15892,N_12845,N_15256);
nor U15893 (N_15893,N_13517,N_12661);
nand U15894 (N_15894,N_14249,N_14490);
nand U15895 (N_15895,N_12877,N_14602);
nand U15896 (N_15896,N_12821,N_15153);
nand U15897 (N_15897,N_13327,N_13937);
and U15898 (N_15898,N_14021,N_15609);
or U15899 (N_15899,N_15152,N_14325);
or U15900 (N_15900,N_13275,N_14709);
and U15901 (N_15901,N_14754,N_13548);
xor U15902 (N_15902,N_14279,N_14927);
or U15903 (N_15903,N_13457,N_14802);
nor U15904 (N_15904,N_14314,N_13878);
xnor U15905 (N_15905,N_14877,N_12611);
nor U15906 (N_15906,N_12589,N_14405);
xnor U15907 (N_15907,N_15157,N_14260);
and U15908 (N_15908,N_14182,N_14463);
xnor U15909 (N_15909,N_14092,N_14837);
or U15910 (N_15910,N_14439,N_15598);
xor U15911 (N_15911,N_13106,N_13282);
or U15912 (N_15912,N_12558,N_15582);
nor U15913 (N_15913,N_14795,N_13675);
nand U15914 (N_15914,N_15567,N_14744);
xnor U15915 (N_15915,N_13619,N_13986);
nor U15916 (N_15916,N_13520,N_13518);
and U15917 (N_15917,N_14049,N_13052);
and U15918 (N_15918,N_15602,N_13799);
nand U15919 (N_15919,N_12543,N_15057);
nand U15920 (N_15920,N_14947,N_14315);
nand U15921 (N_15921,N_13682,N_15597);
or U15922 (N_15922,N_15329,N_14207);
or U15923 (N_15923,N_13737,N_12753);
xnor U15924 (N_15924,N_13429,N_15420);
nor U15925 (N_15925,N_15246,N_14313);
nand U15926 (N_15926,N_12524,N_13728);
nand U15927 (N_15927,N_12506,N_15421);
xor U15928 (N_15928,N_14760,N_14362);
nor U15929 (N_15929,N_13815,N_14047);
nor U15930 (N_15930,N_14977,N_13717);
nor U15931 (N_15931,N_13507,N_12992);
or U15932 (N_15932,N_14071,N_13869);
xnor U15933 (N_15933,N_14848,N_12688);
nand U15934 (N_15934,N_15585,N_14704);
or U15935 (N_15935,N_14674,N_14132);
xnor U15936 (N_15936,N_13311,N_13412);
nand U15937 (N_15937,N_13182,N_13022);
xor U15938 (N_15938,N_13033,N_14456);
and U15939 (N_15939,N_12581,N_15134);
and U15940 (N_15940,N_15558,N_15080);
xnor U15941 (N_15941,N_12539,N_14817);
nor U15942 (N_15942,N_12954,N_14016);
and U15943 (N_15943,N_14641,N_13803);
xnor U15944 (N_15944,N_14003,N_13152);
nand U15945 (N_15945,N_15019,N_13254);
nand U15946 (N_15946,N_14385,N_12636);
nand U15947 (N_15947,N_13991,N_13844);
xor U15948 (N_15948,N_14146,N_15320);
nand U15949 (N_15949,N_14918,N_14696);
or U15950 (N_15950,N_15175,N_12755);
and U15951 (N_15951,N_14662,N_15006);
and U15952 (N_15952,N_12928,N_13604);
and U15953 (N_15953,N_13178,N_14444);
xnor U15954 (N_15954,N_13764,N_14820);
or U15955 (N_15955,N_15370,N_12778);
nand U15956 (N_15956,N_15228,N_14232);
nor U15957 (N_15957,N_13001,N_13685);
xnor U15958 (N_15958,N_13217,N_13773);
nand U15959 (N_15959,N_13075,N_14577);
xnor U15960 (N_15960,N_15416,N_13765);
and U15961 (N_15961,N_14236,N_14555);
nor U15962 (N_15962,N_15144,N_12815);
and U15963 (N_15963,N_13593,N_12553);
or U15964 (N_15964,N_14247,N_15594);
xor U15965 (N_15965,N_12797,N_15171);
xnor U15966 (N_15966,N_12911,N_13797);
nor U15967 (N_15967,N_14975,N_12995);
nand U15968 (N_15968,N_13136,N_14697);
nand U15969 (N_15969,N_12886,N_13602);
nor U15970 (N_15970,N_15349,N_13258);
or U15971 (N_15971,N_14174,N_13512);
nand U15972 (N_15972,N_13476,N_13195);
xnor U15973 (N_15973,N_14706,N_14370);
xnor U15974 (N_15974,N_13145,N_15191);
xnor U15975 (N_15975,N_15211,N_14660);
nand U15976 (N_15976,N_12621,N_13072);
xnor U15977 (N_15977,N_14831,N_13201);
nand U15978 (N_15978,N_15116,N_13891);
and U15979 (N_15979,N_13255,N_14575);
or U15980 (N_15980,N_15396,N_12813);
nor U15981 (N_15981,N_13293,N_13503);
nor U15982 (N_15982,N_14097,N_13436);
or U15983 (N_15983,N_13897,N_12710);
xnor U15984 (N_15984,N_14212,N_15369);
nor U15985 (N_15985,N_13967,N_14594);
and U15986 (N_15986,N_12674,N_15467);
or U15987 (N_15987,N_15036,N_12987);
xnor U15988 (N_15988,N_13270,N_12991);
and U15989 (N_15989,N_14307,N_12601);
or U15990 (N_15990,N_12716,N_13383);
nor U15991 (N_15991,N_14250,N_13847);
xor U15992 (N_15992,N_13839,N_13581);
or U15993 (N_15993,N_15244,N_15408);
nor U15994 (N_15994,N_14530,N_13915);
xor U15995 (N_15995,N_13780,N_13197);
nand U15996 (N_15996,N_13622,N_12783);
nor U15997 (N_15997,N_13641,N_13405);
xnor U15998 (N_15998,N_12872,N_14296);
xor U15999 (N_15999,N_13365,N_12915);
xnor U16000 (N_16000,N_13235,N_12791);
xor U16001 (N_16001,N_14535,N_13213);
or U16002 (N_16002,N_13669,N_12804);
or U16003 (N_16003,N_13078,N_13461);
or U16004 (N_16004,N_13908,N_15070);
and U16005 (N_16005,N_14901,N_13014);
nand U16006 (N_16006,N_12744,N_13911);
nor U16007 (N_16007,N_12944,N_14711);
or U16008 (N_16008,N_12656,N_14909);
or U16009 (N_16009,N_14890,N_14265);
and U16010 (N_16010,N_12556,N_13667);
xor U16011 (N_16011,N_12747,N_12535);
and U16012 (N_16012,N_14149,N_14366);
or U16013 (N_16013,N_15115,N_14636);
xnor U16014 (N_16014,N_13393,N_15093);
nand U16015 (N_16015,N_14545,N_12883);
nand U16016 (N_16016,N_13849,N_14114);
and U16017 (N_16017,N_14283,N_12542);
xnor U16018 (N_16018,N_13743,N_14324);
nor U16019 (N_16019,N_12760,N_14121);
and U16020 (N_16020,N_14982,N_13699);
nand U16021 (N_16021,N_14585,N_12758);
and U16022 (N_16022,N_15114,N_12833);
or U16023 (N_16023,N_15142,N_14202);
or U16024 (N_16024,N_12593,N_14183);
nand U16025 (N_16025,N_13262,N_13444);
xnor U16026 (N_16026,N_15398,N_15301);
xnor U16027 (N_16027,N_13044,N_13065);
xor U16028 (N_16028,N_13183,N_14951);
xnor U16029 (N_16029,N_13524,N_13221);
xnor U16030 (N_16030,N_13759,N_13073);
and U16031 (N_16031,N_15367,N_13627);
nand U16032 (N_16032,N_14567,N_14426);
nor U16033 (N_16033,N_13893,N_14864);
and U16034 (N_16034,N_15049,N_15313);
xor U16035 (N_16035,N_12520,N_12606);
xnor U16036 (N_16036,N_13016,N_13851);
nor U16037 (N_16037,N_12994,N_13666);
or U16038 (N_16038,N_15105,N_12950);
nor U16039 (N_16039,N_15299,N_14251);
nor U16040 (N_16040,N_15517,N_14101);
xor U16041 (N_16041,N_13990,N_13960);
nor U16042 (N_16042,N_13696,N_14936);
nand U16043 (N_16043,N_12846,N_13976);
nor U16044 (N_16044,N_14666,N_12597);
and U16045 (N_16045,N_15276,N_15326);
and U16046 (N_16046,N_13267,N_14393);
or U16047 (N_16047,N_15123,N_15449);
xnor U16048 (N_16048,N_15433,N_12720);
nand U16049 (N_16049,N_12837,N_13151);
or U16050 (N_16050,N_14190,N_14649);
xnor U16051 (N_16051,N_15110,N_14737);
or U16052 (N_16052,N_15426,N_14733);
nor U16053 (N_16053,N_13123,N_14732);
or U16054 (N_16054,N_13713,N_13459);
xor U16055 (N_16055,N_15524,N_12630);
nand U16056 (N_16056,N_13921,N_14195);
nor U16057 (N_16057,N_13303,N_14527);
nand U16058 (N_16058,N_13292,N_14756);
and U16059 (N_16059,N_14792,N_15166);
nor U16060 (N_16060,N_13300,N_14178);
nor U16061 (N_16061,N_14091,N_15346);
xnor U16062 (N_16062,N_12693,N_13872);
or U16063 (N_16063,N_13043,N_15472);
nand U16064 (N_16064,N_13906,N_13362);
nand U16065 (N_16065,N_15492,N_15584);
and U16066 (N_16066,N_13416,N_12598);
and U16067 (N_16067,N_14402,N_15546);
nand U16068 (N_16068,N_14794,N_14287);
nand U16069 (N_16069,N_14834,N_13726);
or U16070 (N_16070,N_14053,N_13532);
and U16071 (N_16071,N_14246,N_15126);
nor U16072 (N_16072,N_13269,N_14782);
xor U16073 (N_16073,N_15133,N_14368);
or U16074 (N_16074,N_14032,N_15324);
nand U16075 (N_16075,N_14618,N_13150);
nor U16076 (N_16076,N_14124,N_13884);
or U16077 (N_16077,N_12839,N_15081);
nand U16078 (N_16078,N_14692,N_13228);
or U16079 (N_16079,N_13903,N_15615);
nand U16080 (N_16080,N_15427,N_15391);
nand U16081 (N_16081,N_15188,N_15525);
nor U16082 (N_16082,N_14987,N_14056);
or U16083 (N_16083,N_13966,N_15248);
nand U16084 (N_16084,N_12771,N_13568);
or U16085 (N_16085,N_12919,N_13242);
or U16086 (N_16086,N_13875,N_14775);
xor U16087 (N_16087,N_14596,N_13935);
and U16088 (N_16088,N_13169,N_15227);
nor U16089 (N_16089,N_14872,N_12762);
nor U16090 (N_16090,N_13754,N_13186);
or U16091 (N_16091,N_13294,N_13087);
xnor U16092 (N_16092,N_12584,N_15573);
xor U16093 (N_16093,N_14825,N_13650);
xor U16094 (N_16094,N_13687,N_13252);
or U16095 (N_16095,N_15607,N_14081);
or U16096 (N_16096,N_14382,N_13530);
nand U16097 (N_16097,N_12708,N_12574);
or U16098 (N_16098,N_15147,N_12805);
nand U16099 (N_16099,N_13900,N_12924);
nor U16100 (N_16100,N_14736,N_14333);
xnor U16101 (N_16101,N_14187,N_14805);
and U16102 (N_16102,N_14511,N_14945);
and U16103 (N_16103,N_14978,N_14031);
or U16104 (N_16104,N_15380,N_14215);
xnor U16105 (N_16105,N_13733,N_15414);
or U16106 (N_16106,N_13238,N_12857);
or U16107 (N_16107,N_12767,N_15366);
xor U16108 (N_16108,N_15173,N_13695);
or U16109 (N_16109,N_15444,N_12852);
and U16110 (N_16110,N_14904,N_14643);
or U16111 (N_16111,N_13505,N_13702);
nor U16112 (N_16112,N_12789,N_14022);
or U16113 (N_16113,N_15343,N_13046);
and U16114 (N_16114,N_15042,N_14453);
nor U16115 (N_16115,N_14639,N_14170);
nand U16116 (N_16116,N_13980,N_15028);
or U16117 (N_16117,N_12930,N_14562);
nor U16118 (N_16118,N_14017,N_12641);
xor U16119 (N_16119,N_12990,N_13866);
or U16120 (N_16120,N_13279,N_15392);
or U16121 (N_16121,N_13817,N_13317);
xnor U16122 (N_16122,N_13859,N_14454);
nor U16123 (N_16123,N_15510,N_13600);
xnor U16124 (N_16124,N_14684,N_12751);
and U16125 (N_16125,N_14522,N_14598);
and U16126 (N_16126,N_13801,N_13925);
nand U16127 (N_16127,N_14128,N_13901);
nand U16128 (N_16128,N_14560,N_13363);
xnor U16129 (N_16129,N_14813,N_13561);
nand U16130 (N_16130,N_12861,N_12665);
nand U16131 (N_16131,N_12610,N_15548);
and U16132 (N_16132,N_14789,N_13432);
or U16133 (N_16133,N_12961,N_13062);
or U16134 (N_16134,N_13660,N_14897);
xnor U16135 (N_16135,N_14748,N_15088);
or U16136 (N_16136,N_13784,N_13770);
or U16137 (N_16137,N_12996,N_14259);
and U16138 (N_16138,N_13610,N_12536);
nand U16139 (N_16139,N_15590,N_12946);
nor U16140 (N_16140,N_12976,N_14241);
xor U16141 (N_16141,N_14824,N_14554);
nor U16142 (N_16142,N_15487,N_13919);
xnor U16143 (N_16143,N_14334,N_15100);
nor U16144 (N_16144,N_14396,N_15178);
nor U16145 (N_16145,N_12570,N_13536);
nor U16146 (N_16146,N_14230,N_13741);
nand U16147 (N_16147,N_12501,N_13441);
or U16148 (N_16148,N_13329,N_13284);
and U16149 (N_16149,N_15515,N_14838);
xor U16150 (N_16150,N_13606,N_14773);
xnor U16151 (N_16151,N_12619,N_12856);
nor U16152 (N_16152,N_14278,N_14665);
xor U16153 (N_16153,N_13640,N_15431);
and U16154 (N_16154,N_13564,N_14675);
and U16155 (N_16155,N_15038,N_13477);
nor U16156 (N_16156,N_14774,N_14896);
nand U16157 (N_16157,N_15432,N_12899);
nand U16158 (N_16158,N_12529,N_12967);
nor U16159 (N_16159,N_12668,N_15310);
or U16160 (N_16160,N_12712,N_13229);
nor U16161 (N_16161,N_15176,N_13163);
or U16162 (N_16162,N_13588,N_14494);
nor U16163 (N_16163,N_15150,N_13502);
nand U16164 (N_16164,N_13351,N_14566);
xnor U16165 (N_16165,N_14478,N_14510);
and U16166 (N_16166,N_14095,N_13251);
and U16167 (N_16167,N_14714,N_12516);
and U16168 (N_16168,N_15059,N_15557);
xor U16169 (N_16169,N_12522,N_13756);
and U16170 (N_16170,N_14339,N_15013);
xnor U16171 (N_16171,N_13096,N_15204);
and U16172 (N_16172,N_12998,N_13177);
nor U16173 (N_16173,N_15247,N_13763);
nand U16174 (N_16174,N_14889,N_14350);
xnor U16175 (N_16175,N_13541,N_13359);
nand U16176 (N_16176,N_14203,N_13941);
and U16177 (N_16177,N_15503,N_14752);
or U16178 (N_16178,N_15574,N_13449);
nor U16179 (N_16179,N_14390,N_15132);
or U16180 (N_16180,N_13577,N_12733);
nor U16181 (N_16181,N_14264,N_14328);
xnor U16182 (N_16182,N_13969,N_13787);
and U16183 (N_16183,N_13008,N_14518);
nor U16184 (N_16184,N_15321,N_14949);
or U16185 (N_16185,N_14272,N_14544);
nor U16186 (N_16186,N_13721,N_13142);
nor U16187 (N_16187,N_13744,N_14143);
xnor U16188 (N_16188,N_14105,N_12603);
or U16189 (N_16189,N_14731,N_13620);
and U16190 (N_16190,N_13450,N_13566);
nor U16191 (N_16191,N_12732,N_14353);
nor U16192 (N_16192,N_12853,N_14926);
nand U16193 (N_16193,N_12602,N_12623);
nor U16194 (N_16194,N_15401,N_12615);
or U16195 (N_16195,N_14414,N_14181);
xnor U16196 (N_16196,N_14373,N_12869);
xor U16197 (N_16197,N_12515,N_15296);
nand U16198 (N_16198,N_13356,N_13578);
nand U16199 (N_16199,N_14959,N_15439);
nand U16200 (N_16200,N_13769,N_14574);
and U16201 (N_16201,N_14015,N_14440);
nand U16202 (N_16202,N_15120,N_13475);
or U16203 (N_16203,N_12798,N_15254);
or U16204 (N_16204,N_15111,N_13688);
xnor U16205 (N_16205,N_14503,N_15413);
xnor U16206 (N_16206,N_13735,N_12832);
and U16207 (N_16207,N_14708,N_14403);
and U16208 (N_16208,N_15312,N_15230);
nand U16209 (N_16209,N_15289,N_12681);
xnor U16210 (N_16210,N_14916,N_13983);
nand U16211 (N_16211,N_13584,N_15620);
xnor U16212 (N_16212,N_13731,N_15182);
and U16213 (N_16213,N_15450,N_14395);
or U16214 (N_16214,N_15017,N_14668);
or U16215 (N_16215,N_12538,N_15051);
nand U16216 (N_16216,N_14609,N_13041);
or U16217 (N_16217,N_12907,N_14631);
nor U16218 (N_16218,N_15288,N_13777);
nand U16219 (N_16219,N_15024,N_14455);
xnor U16220 (N_16220,N_12881,N_13378);
nor U16221 (N_16221,N_12896,N_13323);
nand U16222 (N_16222,N_14011,N_12786);
and U16223 (N_16223,N_13039,N_15565);
nor U16224 (N_16224,N_13206,N_15225);
or U16225 (N_16225,N_13295,N_14109);
or U16226 (N_16226,N_13401,N_15371);
nand U16227 (N_16227,N_13813,N_12507);
nor U16228 (N_16228,N_15071,N_12969);
nor U16229 (N_16229,N_13017,N_13998);
xor U16230 (N_16230,N_14981,N_14499);
and U16231 (N_16231,N_14401,N_14222);
or U16232 (N_16232,N_13367,N_15164);
or U16233 (N_16233,N_13122,N_13304);
and U16234 (N_16234,N_13571,N_14961);
nor U16235 (N_16235,N_13308,N_13482);
xnor U16236 (N_16236,N_13369,N_12525);
nand U16237 (N_16237,N_13333,N_14372);
and U16238 (N_16238,N_13729,N_14327);
nand U16239 (N_16239,N_13319,N_12599);
nor U16240 (N_16240,N_13842,N_13302);
nand U16241 (N_16241,N_13330,N_13704);
xor U16242 (N_16242,N_15112,N_13821);
nor U16243 (N_16243,N_12974,N_14786);
or U16244 (N_16244,N_15376,N_14924);
nor U16245 (N_16245,N_13337,N_13956);
nor U16246 (N_16246,N_13642,N_14068);
and U16247 (N_16247,N_12867,N_15554);
or U16248 (N_16248,N_15453,N_12699);
or U16249 (N_16249,N_13495,N_12626);
xnor U16250 (N_16250,N_15281,N_15507);
or U16251 (N_16251,N_15465,N_13719);
xnor U16252 (N_16252,N_14933,N_15290);
and U16253 (N_16253,N_15566,N_13557);
and U16254 (N_16254,N_13615,N_13036);
and U16255 (N_16255,N_12721,N_13331);
nor U16256 (N_16256,N_13997,N_13139);
or U16257 (N_16257,N_14479,N_14108);
or U16258 (N_16258,N_15183,N_13519);
nand U16259 (N_16259,N_13950,N_13852);
nor U16260 (N_16260,N_14311,N_14698);
nor U16261 (N_16261,N_13651,N_13025);
nand U16262 (N_16262,N_12504,N_14361);
nand U16263 (N_16263,N_14094,N_14991);
or U16264 (N_16264,N_13472,N_12814);
and U16265 (N_16265,N_14862,N_13156);
and U16266 (N_16266,N_13483,N_12582);
nand U16267 (N_16267,N_14983,N_15030);
and U16268 (N_16268,N_14712,N_13510);
nor U16269 (N_16269,N_15541,N_14486);
nand U16270 (N_16270,N_15170,N_14277);
xor U16271 (N_16271,N_12534,N_15122);
and U16272 (N_16272,N_13371,N_12639);
nand U16273 (N_16273,N_13212,N_14150);
nor U16274 (N_16274,N_15026,N_13486);
or U16275 (N_16275,N_12923,N_15333);
and U16276 (N_16276,N_13200,N_13281);
xor U16277 (N_16277,N_13121,N_15032);
or U16278 (N_16278,N_14286,N_14162);
nor U16279 (N_16279,N_13103,N_12622);
nor U16280 (N_16280,N_13161,N_14467);
nor U16281 (N_16281,N_12637,N_15151);
xnor U16282 (N_16282,N_14656,N_13045);
xnor U16283 (N_16283,N_14039,N_15613);
or U16284 (N_16284,N_13924,N_13993);
nor U16285 (N_16285,N_15291,N_12583);
xnor U16286 (N_16286,N_12842,N_15207);
xnor U16287 (N_16287,N_15197,N_13250);
or U16288 (N_16288,N_12701,N_13496);
and U16289 (N_16289,N_13886,N_15186);
nand U16290 (N_16290,N_13403,N_14089);
nand U16291 (N_16291,N_13962,N_15417);
nand U16292 (N_16292,N_14899,N_14495);
xnor U16293 (N_16293,N_13484,N_15352);
nand U16294 (N_16294,N_12579,N_14571);
nand U16295 (N_16295,N_12940,N_13690);
nor U16296 (N_16296,N_14705,N_13411);
or U16297 (N_16297,N_14156,N_12557);
xnor U16298 (N_16298,N_13092,N_15121);
nor U16299 (N_16299,N_12748,N_13463);
xor U16300 (N_16300,N_13968,N_14107);
or U16301 (N_16301,N_14944,N_13783);
nor U16302 (N_16302,N_14219,N_14099);
nand U16303 (N_16303,N_15384,N_15086);
or U16304 (N_16304,N_15534,N_13234);
nand U16305 (N_16305,N_13544,N_14201);
and U16306 (N_16306,N_13372,N_14112);
xnor U16307 (N_16307,N_13076,N_12700);
and U16308 (N_16308,N_14085,N_15212);
or U16309 (N_16309,N_12906,N_14090);
or U16310 (N_16310,N_13368,N_14874);
nor U16311 (N_16311,N_15545,N_15084);
and U16312 (N_16312,N_14226,N_13778);
and U16313 (N_16313,N_14663,N_13445);
and U16314 (N_16314,N_14866,N_14906);
nor U16315 (N_16315,N_14106,N_15375);
or U16316 (N_16316,N_14102,N_14189);
xnor U16317 (N_16317,N_13082,N_12864);
or U16318 (N_16318,N_13776,N_12564);
nand U16319 (N_16319,N_14061,N_13658);
or U16320 (N_16320,N_14597,N_12949);
nand U16321 (N_16321,N_12971,N_13987);
nor U16322 (N_16322,N_13616,N_13703);
and U16323 (N_16323,N_13710,N_13247);
nand U16324 (N_16324,N_15102,N_13670);
nand U16325 (N_16325,N_15240,N_15218);
or U16326 (N_16326,N_12939,N_14052);
or U16327 (N_16327,N_14531,N_12576);
or U16328 (N_16328,N_15363,N_14084);
nand U16329 (N_16329,N_12972,N_15559);
xnor U16330 (N_16330,N_13896,N_14507);
nand U16331 (N_16331,N_15187,N_13802);
or U16332 (N_16332,N_15098,N_15033);
and U16333 (N_16333,N_14235,N_12963);
nor U16334 (N_16334,N_15511,N_15564);
xnor U16335 (N_16335,N_13446,N_12838);
xor U16336 (N_16336,N_15002,N_15357);
xor U16337 (N_16337,N_13549,N_15470);
and U16338 (N_16338,N_15091,N_14826);
xnor U16339 (N_16339,N_15440,N_15160);
and U16340 (N_16340,N_14845,N_13972);
and U16341 (N_16341,N_13180,N_12809);
xnor U16342 (N_16342,N_13248,N_13026);
nor U16343 (N_16343,N_14986,N_12843);
xnor U16344 (N_16344,N_14646,N_14254);
xor U16345 (N_16345,N_12826,N_13318);
nand U16346 (N_16346,N_14604,N_13126);
xor U16347 (N_16347,N_13766,N_13938);
nand U16348 (N_16348,N_14667,N_13397);
nor U16349 (N_16349,N_15053,N_14476);
or U16350 (N_16350,N_15322,N_15179);
nor U16351 (N_16351,N_13558,N_14812);
or U16352 (N_16352,N_14298,N_14319);
nor U16353 (N_16353,N_13125,N_15527);
nand U16354 (N_16354,N_12765,N_15309);
xor U16355 (N_16355,N_12945,N_14351);
xor U16356 (N_16356,N_15466,N_15347);
nor U16357 (N_16357,N_13328,N_12858);
nand U16358 (N_16358,N_14900,N_14957);
or U16359 (N_16359,N_13452,N_13632);
nor U16360 (N_16360,N_12652,N_14819);
nand U16361 (N_16361,N_14908,N_12955);
nand U16362 (N_16362,N_14268,N_12794);
or U16363 (N_16363,N_13256,N_13454);
xor U16364 (N_16364,N_14481,N_14231);
nand U16365 (N_16365,N_13347,N_13811);
xor U16366 (N_16366,N_14707,N_15495);
or U16367 (N_16367,N_12870,N_13479);
and U16368 (N_16368,N_15617,N_12871);
or U16369 (N_16369,N_13135,N_12692);
xnor U16370 (N_16370,N_14648,N_13711);
nor U16371 (N_16371,N_15258,N_14445);
nor U16372 (N_16372,N_13138,N_13768);
and U16373 (N_16373,N_15016,N_15488);
nand U16374 (N_16374,N_12938,N_14023);
and U16375 (N_16375,N_13458,N_13715);
and U16376 (N_16376,N_14500,N_14735);
xor U16377 (N_16377,N_12812,N_14337);
xor U16378 (N_16378,N_12512,N_12618);
or U16379 (N_16379,N_12715,N_15499);
nand U16380 (N_16380,N_15459,N_15591);
and U16381 (N_16381,N_13060,N_15131);
nand U16382 (N_16382,N_14257,N_13879);
and U16383 (N_16383,N_14240,N_15113);
xor U16384 (N_16384,N_12655,N_13618);
and U16385 (N_16385,N_12595,N_14502);
and U16386 (N_16386,N_15263,N_14657);
or U16387 (N_16387,N_13824,N_14205);
xor U16388 (N_16388,N_14135,N_14930);
xnor U16389 (N_16389,N_15060,N_15578);
or U16390 (N_16390,N_12752,N_13322);
nor U16391 (N_16391,N_15275,N_15430);
and U16392 (N_16392,N_13917,N_13400);
nor U16393 (N_16393,N_13392,N_15229);
xnor U16394 (N_16394,N_13643,N_13188);
xor U16395 (N_16395,N_14176,N_12646);
nand U16396 (N_16396,N_14827,N_14879);
and U16397 (N_16397,N_15158,N_14534);
nand U16398 (N_16398,N_15262,N_15563);
nor U16399 (N_16399,N_12986,N_14341);
xnor U16400 (N_16400,N_13244,N_13603);
xnor U16401 (N_16401,N_12572,N_14809);
xor U16402 (N_16402,N_15050,N_15316);
or U16403 (N_16403,N_14284,N_13382);
nor U16404 (N_16404,N_13198,N_14419);
xnor U16405 (N_16405,N_13291,N_14464);
xor U16406 (N_16406,N_13010,N_13628);
or U16407 (N_16407,N_15023,N_13582);
and U16408 (N_16408,N_14990,N_14974);
and U16409 (N_16409,N_15386,N_15344);
or U16410 (N_16410,N_14305,N_13550);
and U16411 (N_16411,N_13358,N_13063);
nor U16412 (N_16412,N_12766,N_12893);
nand U16413 (N_16413,N_13455,N_14856);
and U16414 (N_16414,N_14840,N_14683);
xnor U16415 (N_16415,N_12787,N_13978);
nand U16416 (N_16416,N_14407,N_12677);
nor U16417 (N_16417,N_14871,N_15282);
nand U16418 (N_16418,N_14543,N_15438);
or U16419 (N_16419,N_13944,N_14846);
xor U16420 (N_16420,N_14129,N_13129);
and U16421 (N_16421,N_14059,N_13533);
or U16422 (N_16422,N_15280,N_13099);
nor U16423 (N_16423,N_12904,N_12518);
or U16424 (N_16424,N_14891,N_13224);
nand U16425 (N_16425,N_15037,N_15405);
nor U16426 (N_16426,N_12818,N_14780);
and U16427 (N_16427,N_12617,N_12965);
and U16428 (N_16428,N_13638,N_13992);
nand U16429 (N_16429,N_13579,N_12759);
or U16430 (N_16430,N_14694,N_13435);
or U16431 (N_16431,N_13422,N_14689);
or U16432 (N_16432,N_13048,N_13694);
xor U16433 (N_16433,N_14878,N_13410);
and U16434 (N_16434,N_14460,N_14432);
nor U16435 (N_16435,N_12648,N_13243);
or U16436 (N_16436,N_15167,N_14033);
xnor U16437 (N_16437,N_14673,N_12573);
nand U16438 (N_16438,N_14912,N_15146);
xor U16439 (N_16439,N_13614,N_15595);
xnor U16440 (N_16440,N_13364,N_13833);
and U16441 (N_16441,N_15514,N_12730);
xor U16442 (N_16442,N_15149,N_13996);
nor U16443 (N_16443,N_13723,N_15039);
xor U16444 (N_16444,N_15508,N_12717);
or U16445 (N_16445,N_14627,N_13531);
and U16446 (N_16446,N_12585,N_13882);
nor U16447 (N_16447,N_13943,N_14647);
xnor U16448 (N_16448,N_15139,N_14253);
or U16449 (N_16449,N_13623,N_14019);
or U16450 (N_16450,N_14808,N_13268);
and U16451 (N_16451,N_14855,N_14519);
xor U16452 (N_16452,N_13761,N_12657);
and U16453 (N_16453,N_15311,N_12975);
or U16454 (N_16454,N_15300,N_14332);
or U16455 (N_16455,N_14148,N_13825);
or U16456 (N_16456,N_14412,N_13516);
nand U16457 (N_16457,N_15315,N_13838);
nor U16458 (N_16458,N_12897,N_12625);
nor U16459 (N_16459,N_12824,N_12776);
or U16460 (N_16460,N_15169,N_15097);
nor U16461 (N_16461,N_14243,N_14512);
xnor U16462 (N_16462,N_15058,N_15475);
or U16463 (N_16463,N_14931,N_13088);
or U16464 (N_16464,N_15441,N_13959);
xor U16465 (N_16465,N_13738,N_15593);
and U16466 (N_16466,N_12675,N_14757);
nor U16467 (N_16467,N_14399,N_14179);
and U16468 (N_16468,N_13061,N_13753);
or U16469 (N_16469,N_13027,N_13404);
nor U16470 (N_16470,N_14801,N_15094);
or U16471 (N_16471,N_13345,N_14331);
nand U16472 (N_16472,N_14952,N_15304);
nand U16473 (N_16473,N_14650,N_15206);
nand U16474 (N_16474,N_14514,N_15549);
xor U16475 (N_16475,N_12825,N_13240);
or U16476 (N_16476,N_14173,N_14741);
xor U16477 (N_16477,N_15528,N_13231);
and U16478 (N_16478,N_14224,N_13116);
nor U16479 (N_16479,N_12698,N_15292);
nand U16480 (N_16480,N_14509,N_13488);
nand U16481 (N_16481,N_14942,N_13074);
and U16482 (N_16482,N_14655,N_12802);
nor U16483 (N_16483,N_15576,N_13672);
and U16484 (N_16484,N_13793,N_14632);
and U16485 (N_16485,N_15429,N_13647);
xor U16486 (N_16486,N_15520,N_15205);
nor U16487 (N_16487,N_15189,N_13118);
nand U16488 (N_16488,N_13834,N_14932);
nor U16489 (N_16489,N_15572,N_14430);
xnor U16490 (N_16490,N_14406,N_14994);
xnor U16491 (N_16491,N_12957,N_14029);
and U16492 (N_16492,N_13569,N_13850);
nor U16493 (N_16493,N_14027,N_13873);
or U16494 (N_16494,N_14077,N_14859);
and U16495 (N_16495,N_13140,N_13297);
xor U16496 (N_16496,N_14564,N_13923);
or U16497 (N_16497,N_13490,N_14921);
and U16498 (N_16498,N_12854,N_13984);
nor U16499 (N_16499,N_13771,N_14976);
or U16500 (N_16500,N_13829,N_12775);
and U16501 (N_16501,N_14180,N_13070);
nor U16502 (N_16502,N_13942,N_15104);
xnor U16503 (N_16503,N_14055,N_14060);
and U16504 (N_16504,N_14484,N_14058);
and U16505 (N_16505,N_15319,N_14844);
xor U16506 (N_16506,N_14658,N_13493);
xor U16507 (N_16507,N_12642,N_13339);
nor U16508 (N_16508,N_15519,N_14335);
nand U16509 (N_16509,N_14861,N_15583);
and U16510 (N_16510,N_15004,N_14893);
xnor U16511 (N_16511,N_13006,N_13973);
or U16512 (N_16512,N_12724,N_12964);
and U16513 (N_16513,N_13420,N_14326);
or U16514 (N_16514,N_12840,N_14480);
and U16515 (N_16515,N_14579,N_14225);
nor U16516 (N_16516,N_15512,N_14849);
xor U16517 (N_16517,N_13662,N_15018);
or U16518 (N_16518,N_14747,N_13587);
or U16519 (N_16519,N_13338,N_12937);
nor U16520 (N_16520,N_14769,N_15502);
nor U16521 (N_16521,N_15044,N_15325);
and U16522 (N_16522,N_15163,N_14024);
nor U16523 (N_16523,N_14001,N_12532);
and U16524 (N_16524,N_13462,N_15156);
and U16525 (N_16525,N_14130,N_13336);
or U16526 (N_16526,N_13818,N_13665);
nand U16527 (N_16527,N_14216,N_15378);
nand U16528 (N_16528,N_14922,N_13414);
and U16529 (N_16529,N_13278,N_15025);
nor U16530 (N_16530,N_13940,N_15106);
and U16531 (N_16531,N_15388,N_14359);
or U16532 (N_16532,N_12530,N_14573);
nand U16533 (N_16533,N_14357,N_14087);
and U16534 (N_16534,N_14488,N_14276);
nor U16535 (N_16535,N_12985,N_13202);
nor U16536 (N_16536,N_13226,N_13236);
xor U16537 (N_16537,N_13266,N_12878);
xor U16538 (N_16538,N_15154,N_13260);
and U16539 (N_16539,N_15010,N_14417);
or U16540 (N_16540,N_14437,N_12909);
and U16541 (N_16541,N_14057,N_15422);
xnor U16542 (N_16542,N_14157,N_13583);
nand U16543 (N_16543,N_15135,N_13332);
nor U16544 (N_16544,N_13276,N_15600);
and U16545 (N_16545,N_13885,N_14371);
or U16546 (N_16546,N_15235,N_15103);
or U16547 (N_16547,N_13601,N_14886);
nor U16548 (N_16548,N_13421,N_14626);
nand U16549 (N_16549,N_12643,N_14777);
nand U16550 (N_16550,N_15361,N_14659);
nand U16551 (N_16551,N_14508,N_15155);
or U16552 (N_16552,N_14294,N_15618);
and U16553 (N_16553,N_14165,N_14434);
or U16554 (N_16554,N_14717,N_12605);
xnor U16555 (N_16555,N_14465,N_15308);
nand U16556 (N_16556,N_13035,N_13473);
xor U16557 (N_16557,N_12953,N_14556);
nand U16558 (N_16558,N_14078,N_14233);
xnor U16559 (N_16559,N_15127,N_13525);
xor U16560 (N_16560,N_12705,N_13590);
nand U16561 (N_16561,N_13730,N_13196);
or U16562 (N_16562,N_13112,N_15616);
and U16563 (N_16563,N_15483,N_13119);
or U16564 (N_16564,N_12691,N_15270);
or U16565 (N_16565,N_14881,N_12650);
and U16566 (N_16566,N_12592,N_14119);
and U16567 (N_16567,N_14929,N_12873);
xnor U16568 (N_16568,N_15172,N_14380);
and U16569 (N_16569,N_13863,N_13058);
nor U16570 (N_16570,N_14073,N_13555);
nor U16571 (N_16571,N_12627,N_12587);
xnor U16572 (N_16572,N_15348,N_12695);
and U16573 (N_16573,N_15124,N_13909);
xor U16574 (N_16574,N_13830,N_12910);
nand U16575 (N_16575,N_14835,N_14751);
xnor U16576 (N_16576,N_15328,N_15614);
or U16577 (N_16577,N_13273,N_12891);
nand U16578 (N_16578,N_15020,N_15448);
nor U16579 (N_16579,N_14046,N_15407);
xnor U16580 (N_16580,N_14140,N_13024);
nor U16581 (N_16581,N_12770,N_14164);
xnor U16582 (N_16582,N_13162,N_13137);
and U16583 (N_16583,N_15592,N_12943);
xor U16584 (N_16584,N_13521,N_13375);
xor U16585 (N_16585,N_15473,N_15259);
nor U16586 (N_16586,N_13762,N_14783);
nor U16587 (N_16587,N_13120,N_15505);
nand U16588 (N_16588,N_13649,N_15061);
and U16589 (N_16589,N_13030,N_13453);
nor U16590 (N_16590,N_13309,N_14988);
nand U16591 (N_16591,N_12616,N_14248);
or U16592 (N_16592,N_12624,N_15365);
xor U16593 (N_16593,N_13406,N_12892);
nor U16594 (N_16594,N_12887,N_15457);
xor U16595 (N_16595,N_13592,N_14223);
nor U16596 (N_16596,N_14387,N_14762);
or U16597 (N_16597,N_13428,N_14729);
or U16598 (N_16598,N_13398,N_12941);
nor U16599 (N_16599,N_12736,N_14798);
and U16600 (N_16600,N_12635,N_15463);
and U16601 (N_16601,N_15522,N_13173);
nand U16602 (N_16602,N_15293,N_13865);
nand U16603 (N_16603,N_14211,N_15353);
and U16604 (N_16604,N_15264,N_13904);
xor U16605 (N_16605,N_12827,N_15257);
nor U16606 (N_16606,N_15202,N_15606);
xnor U16607 (N_16607,N_12550,N_13366);
and U16608 (N_16608,N_14791,N_13098);
or U16609 (N_16609,N_13916,N_13191);
or U16610 (N_16610,N_15569,N_14755);
xnor U16611 (N_16611,N_13325,N_12851);
or U16612 (N_16612,N_15390,N_12526);
or U16613 (N_16613,N_14110,N_12517);
and U16614 (N_16614,N_15532,N_15434);
nand U16615 (N_16615,N_15265,N_13504);
nand U16616 (N_16616,N_14677,N_13513);
nor U16617 (N_16617,N_13617,N_15330);
nand U16618 (N_16618,N_15234,N_13835);
nor U16619 (N_16619,N_14120,N_12612);
and U16620 (N_16620,N_15340,N_14725);
nand U16621 (N_16621,N_13630,N_13537);
or U16622 (N_16622,N_13864,N_14678);
and U16623 (N_16623,N_15251,N_13107);
xnor U16624 (N_16624,N_14026,N_12984);
xor U16625 (N_16625,N_13674,N_12568);
and U16626 (N_16626,N_12884,N_12860);
nand U16627 (N_16627,N_15373,N_12596);
and U16628 (N_16628,N_13573,N_13205);
or U16629 (N_16629,N_15418,N_12970);
nor U16630 (N_16630,N_15055,N_12725);
and U16631 (N_16631,N_13971,N_14887);
nand U16632 (N_16632,N_12865,N_12978);
or U16633 (N_16633,N_13902,N_13274);
nor U16634 (N_16634,N_15054,N_13949);
xor U16635 (N_16635,N_14229,N_13348);
or U16636 (N_16636,N_15174,N_13652);
xor U16637 (N_16637,N_14204,N_14785);
nor U16638 (N_16638,N_15368,N_15015);
xor U16639 (N_16639,N_13306,N_15612);
xor U16640 (N_16640,N_13807,N_14832);
or U16641 (N_16641,N_14466,N_14343);
nand U16642 (N_16642,N_15469,N_14570);
nor U16643 (N_16643,N_13469,N_14252);
or U16644 (N_16644,N_13038,N_12831);
nand U16645 (N_16645,N_14472,N_13340);
nand U16646 (N_16646,N_14035,N_13845);
xor U16647 (N_16647,N_14133,N_12722);
and U16648 (N_16648,N_13166,N_14529);
nor U16649 (N_16649,N_15437,N_13492);
nand U16650 (N_16650,N_13750,N_15531);
nand U16651 (N_16651,N_15570,N_13599);
and U16652 (N_16652,N_15445,N_13854);
and U16653 (N_16653,N_14860,N_12952);
xor U16654 (N_16654,N_13246,N_13572);
nand U16655 (N_16655,N_14413,N_12697);
nand U16656 (N_16656,N_14188,N_12551);
xor U16657 (N_16657,N_13700,N_13108);
nand U16658 (N_16658,N_14888,N_13752);
nor U16659 (N_16659,N_13927,N_15046);
nor U16660 (N_16660,N_15236,N_13895);
xnor U16661 (N_16661,N_13725,N_12880);
nand U16662 (N_16662,N_14972,N_13280);
or U16663 (N_16663,N_12781,N_12645);
and U16664 (N_16664,N_15509,N_14002);
nand U16665 (N_16665,N_14653,N_14013);
xnor U16666 (N_16666,N_14913,N_15404);
nand U16667 (N_16667,N_12999,N_12894);
xnor U16668 (N_16668,N_15185,N_13164);
nor U16669 (N_16669,N_14122,N_14894);
nor U16670 (N_16670,N_15342,N_14538);
nor U16671 (N_16671,N_14520,N_12836);
nand U16672 (N_16672,N_13011,N_13781);
or U16673 (N_16673,N_13918,N_12807);
nor U16674 (N_16674,N_14703,N_14558);
and U16675 (N_16675,N_15014,N_12849);
or U16676 (N_16676,N_13631,N_13862);
or U16677 (N_16677,N_13456,N_13051);
xor U16678 (N_16678,N_13644,N_13357);
or U16679 (N_16679,N_14342,N_13856);
nand U16680 (N_16680,N_13460,N_14822);
nor U16681 (N_16681,N_14790,N_13067);
nor U16682 (N_16682,N_14377,N_15468);
and U16683 (N_16683,N_14651,N_14451);
nor U16684 (N_16684,N_15589,N_12683);
nor U16685 (N_16685,N_14778,N_13748);
xor U16686 (N_16686,N_13746,N_14086);
nor U16687 (N_16687,N_12763,N_15516);
nor U16688 (N_16688,N_15551,N_13430);
nand U16689 (N_16689,N_14955,N_12844);
or U16690 (N_16690,N_14329,N_12703);
or U16691 (N_16691,N_14384,N_14184);
or U16692 (N_16692,N_14167,N_12540);
or U16693 (N_16693,N_13168,N_12806);
or U16694 (N_16694,N_12834,N_14779);
nand U16695 (N_16695,N_12927,N_14563);
nor U16696 (N_16696,N_12604,N_15130);
or U16697 (N_16697,N_12889,N_12667);
nand U16698 (N_16698,N_12628,N_12702);
and U16699 (N_16699,N_12855,N_13117);
nor U16700 (N_16700,N_15066,N_13179);
xor U16701 (N_16701,N_15446,N_13312);
and U16702 (N_16702,N_14935,N_14374);
xor U16703 (N_16703,N_13209,N_13396);
nor U16704 (N_16704,N_13408,N_13722);
or U16705 (N_16705,N_13732,N_13352);
nor U16706 (N_16706,N_13963,N_13059);
nor U16707 (N_16707,N_13560,N_14642);
nor U16708 (N_16708,N_13608,N_13970);
nand U16709 (N_16709,N_12729,N_13261);
xnor U16710 (N_16710,N_13843,N_15530);
nor U16711 (N_16711,N_14446,N_15462);
and U16712 (N_16712,N_14828,N_13487);
or U16713 (N_16713,N_14245,N_14261);
nand U16714 (N_16714,N_13553,N_14993);
and U16715 (N_16715,N_13912,N_14258);
nand U16716 (N_16716,N_12925,N_14548);
or U16717 (N_16717,N_15504,N_14297);
xnor U16718 (N_16718,N_15412,N_12993);
and U16719 (N_16719,N_14442,N_14687);
xnor U16720 (N_16720,N_14358,N_12741);
nor U16721 (N_16721,N_14051,N_13394);
nor U16722 (N_16722,N_12659,N_14386);
and U16723 (N_16723,N_15021,N_15279);
or U16724 (N_16724,N_13646,N_13576);
xor U16725 (N_16725,N_13301,N_13645);
xor U16726 (N_16726,N_14613,N_14958);
xor U16727 (N_16727,N_15305,N_12565);
xnor U16728 (N_16728,N_14525,N_13739);
xnor U16729 (N_16729,N_13877,N_13779);
or U16730 (N_16730,N_13720,N_13898);
nor U16731 (N_16731,N_15336,N_15161);
xnor U16732 (N_16732,N_13515,N_12649);
and U16733 (N_16733,N_14397,N_15109);
and U16734 (N_16734,N_12956,N_15266);
xor U16735 (N_16735,N_15272,N_13816);
nor U16736 (N_16736,N_13418,N_12749);
and U16737 (N_16737,N_13514,N_14348);
xor U16738 (N_16738,N_15489,N_13977);
and U16739 (N_16739,N_13227,N_15399);
xnor U16740 (N_16740,N_13349,N_13360);
nor U16741 (N_16741,N_13316,N_15041);
or U16742 (N_16742,N_13343,N_14591);
or U16743 (N_16743,N_14461,N_15089);
and U16744 (N_16744,N_13374,N_13907);
nor U16745 (N_16745,N_13320,N_14686);
xor U16746 (N_16746,N_14303,N_14953);
xnor U16747 (N_16747,N_13961,N_13040);
xnor U16748 (N_16748,N_13335,N_15547);
nand U16749 (N_16749,N_13353,N_13381);
and U16750 (N_16750,N_15243,N_13023);
and U16751 (N_16751,N_13523,N_12726);
or U16752 (N_16752,N_15203,N_13057);
nor U16753 (N_16753,N_15556,N_12935);
nor U16754 (N_16754,N_13341,N_13175);
nor U16755 (N_16755,N_14356,N_13671);
nand U16756 (N_16756,N_12916,N_14066);
nor U16757 (N_16757,N_14160,N_13466);
or U16758 (N_16758,N_12962,N_14652);
nand U16759 (N_16759,N_12947,N_14841);
nor U16760 (N_16760,N_12510,N_13054);
xor U16761 (N_16761,N_13994,N_14787);
nor U16762 (N_16762,N_13434,N_13934);
xnor U16763 (N_16763,N_15506,N_13415);
or U16764 (N_16764,N_12790,N_14428);
or U16765 (N_16765,N_13298,N_14772);
nand U16766 (N_16766,N_14123,N_15484);
nor U16767 (N_16767,N_14450,N_13789);
nand U16768 (N_16768,N_14364,N_14557);
and U16769 (N_16769,N_13709,N_14910);
nand U16770 (N_16770,N_13354,N_15603);
xnor U16771 (N_16771,N_13546,N_13718);
xnor U16772 (N_16772,N_13913,N_15395);
or U16773 (N_16773,N_13791,N_13681);
xnor U16774 (N_16774,N_12644,N_13727);
or U16775 (N_16775,N_13131,N_14766);
nor U16776 (N_16776,N_14547,N_15406);
nor U16777 (N_16777,N_13290,N_15245);
nor U16778 (N_16778,N_14749,N_13130);
xnor U16779 (N_16779,N_13736,N_13823);
or U16780 (N_16780,N_13691,N_14447);
nor U16781 (N_16781,N_13376,N_13594);
xor U16782 (N_16782,N_14125,N_14151);
or U16783 (N_16783,N_14962,N_14048);
and U16784 (N_16784,N_15577,N_14115);
nor U16785 (N_16785,N_12788,N_13575);
nor U16786 (N_16786,N_12566,N_14969);
or U16787 (N_16787,N_12918,N_13423);
xor U16788 (N_16788,N_15447,N_12942);
or U16789 (N_16789,N_15419,N_12653);
or U16790 (N_16790,N_13478,N_13310);
xnor U16791 (N_16791,N_13230,N_13522);
xor U16792 (N_16792,N_14040,N_13080);
or U16793 (N_16793,N_15074,N_13015);
and U16794 (N_16794,N_12546,N_15221);
xor U16795 (N_16795,N_14169,N_14020);
or U16796 (N_16796,N_13981,N_12634);
and U16797 (N_16797,N_14065,N_13132);
xor U16798 (N_16798,N_15274,N_13355);
nor U16799 (N_16799,N_12982,N_13526);
nand U16800 (N_16800,N_15580,N_14080);
nand U16801 (N_16801,N_12528,N_14964);
and U16802 (N_16802,N_12734,N_13342);
and U16803 (N_16803,N_14290,N_14578);
and U16804 (N_16804,N_14285,N_15622);
or U16805 (N_16805,N_12914,N_14137);
nor U16806 (N_16806,N_12773,N_13607);
nand U16807 (N_16807,N_13239,N_14369);
nand U16808 (N_16808,N_14006,N_14606);
xnor U16809 (N_16809,N_13686,N_14971);
xnor U16810 (N_16810,N_13426,N_14728);
and U16811 (N_16811,N_14603,N_13857);
or U16812 (N_16812,N_13160,N_13111);
nand U16813 (N_16813,N_13249,N_14196);
nor U16814 (N_16814,N_15181,N_14869);
nor U16815 (N_16815,N_14920,N_15294);
nand U16816 (N_16816,N_15415,N_15409);
nand U16817 (N_16817,N_13037,N_15383);
and U16818 (N_16818,N_14280,N_14363);
and U16819 (N_16819,N_14487,N_14172);
nor U16820 (N_16820,N_13933,N_13222);
or U16821 (N_16821,N_12664,N_14234);
or U16822 (N_16822,N_13928,N_15099);
and U16823 (N_16823,N_14470,N_14793);
xnor U16824 (N_16824,N_12614,N_14392);
and U16825 (N_16825,N_13110,N_13187);
nand U16826 (N_16826,N_14517,N_12545);
xnor U16827 (N_16827,N_14459,N_12638);
nor U16828 (N_16828,N_12819,N_13899);
nand U16829 (N_16829,N_13870,N_14166);
or U16830 (N_16830,N_14850,N_13299);
xor U16831 (N_16831,N_12895,N_14750);
and U16832 (N_16832,N_13305,N_15476);
and U16833 (N_16833,N_13081,N_12663);
and U16834 (N_16834,N_14851,N_15382);
and U16835 (N_16835,N_15267,N_12511);
nand U16836 (N_16836,N_12746,N_13489);
or U16837 (N_16837,N_14917,N_12997);
and U16838 (N_16838,N_14998,N_13964);
xnor U16839 (N_16839,N_15073,N_15518);
or U16840 (N_16840,N_14992,N_14695);
and U16841 (N_16841,N_12740,N_13105);
or U16842 (N_16842,N_13814,N_15137);
nand U16843 (N_16843,N_13157,N_15423);
nand U16844 (N_16844,N_13554,N_14715);
or U16845 (N_16845,N_14700,N_15198);
or U16846 (N_16846,N_15335,N_15003);
nand U16847 (N_16847,N_14615,N_13951);
and U16848 (N_16848,N_15537,N_13920);
and U16849 (N_16849,N_14740,N_13508);
or U16850 (N_16850,N_14788,N_12654);
nand U16851 (N_16851,N_14501,N_15605);
nor U16852 (N_16852,N_15402,N_14685);
xnor U16853 (N_16853,N_14448,N_15314);
and U16854 (N_16854,N_14810,N_12920);
and U16855 (N_16855,N_12569,N_14070);
nor U16856 (N_16856,N_15374,N_13626);
and U16857 (N_16857,N_13464,N_14293);
or U16858 (N_16858,N_13055,N_14161);
nor U16859 (N_16859,N_12672,N_15586);
xnor U16860 (N_16860,N_13344,N_13018);
xor U16861 (N_16861,N_15454,N_13237);
nand U16862 (N_16862,N_14346,N_14718);
nand U16863 (N_16863,N_15389,N_13880);
or U16864 (N_16864,N_13094,N_14719);
nand U16865 (N_16865,N_14763,N_14193);
xor U16866 (N_16866,N_15360,N_14074);
nor U16867 (N_16867,N_14349,N_14745);
or U16868 (N_16868,N_13208,N_14103);
or U16869 (N_16869,N_13914,N_13806);
or U16870 (N_16870,N_15478,N_13283);
and U16871 (N_16871,N_12687,N_14104);
nor U16872 (N_16872,N_14523,N_14075);
xor U16873 (N_16873,N_15443,N_14028);
nor U16874 (N_16874,N_13562,N_13624);
and U16875 (N_16875,N_14995,N_12739);
nor U16876 (N_16876,N_14880,N_15072);
nand U16877 (N_16877,N_13379,N_14138);
xor U16878 (N_16878,N_15005,N_13635);
or U16879 (N_16879,N_14340,N_14634);
nor U16880 (N_16880,N_13712,N_14175);
xor U16881 (N_16881,N_15411,N_14943);
xnor U16882 (N_16882,N_15200,N_14776);
nor U16883 (N_16883,N_13585,N_13840);
and U16884 (N_16884,N_15596,N_13663);
xor U16885 (N_16885,N_12859,N_14903);
nand U16886 (N_16886,N_12882,N_12948);
nor U16887 (N_16887,N_14418,N_14892);
and U16888 (N_16888,N_12671,N_13211);
xor U16889 (N_16889,N_13171,N_12745);
nand U16890 (N_16890,N_14797,N_12933);
nand U16891 (N_16891,N_13241,N_14635);
and U16892 (N_16892,N_14425,N_14954);
nand U16893 (N_16893,N_12868,N_15159);
nor U16894 (N_16894,N_13402,N_13144);
nor U16895 (N_16895,N_14158,N_13995);
or U16896 (N_16896,N_15220,N_13485);
nor U16897 (N_16897,N_12632,N_12800);
or U16898 (N_16898,N_12571,N_12631);
xor U16899 (N_16899,N_14670,N_15601);
nand U16900 (N_16900,N_14723,N_15007);
nor U16901 (N_16901,N_15162,N_12921);
or U16902 (N_16902,N_13100,N_13855);
nor U16903 (N_16903,N_14528,N_14682);
xor U16904 (N_16904,N_12706,N_13134);
nand U16905 (N_16905,N_12640,N_14088);
or U16906 (N_16906,N_12900,N_12769);
xor U16907 (N_16907,N_14691,N_14572);
and U16908 (N_16908,N_15526,N_12541);
nor U16909 (N_16909,N_14581,N_13926);
nor U16910 (N_16910,N_13953,N_14727);
nand U16911 (N_16911,N_13625,N_14474);
xor U16912 (N_16912,N_14654,N_14391);
and U16913 (N_16913,N_15498,N_15464);
or U16914 (N_16914,N_13947,N_14599);
nand U16915 (N_16915,N_15482,N_15196);
nand U16916 (N_16916,N_13742,N_13580);
nand U16917 (N_16917,N_12968,N_15400);
nand U16918 (N_16918,N_13946,N_13794);
or U16919 (N_16919,N_15136,N_15358);
or U16920 (N_16920,N_14007,N_13786);
nor U16921 (N_16921,N_13114,N_15226);
or U16922 (N_16922,N_12799,N_15297);
xor U16923 (N_16923,N_14355,N_12684);
and U16924 (N_16924,N_13154,N_13798);
xor U16925 (N_16925,N_13543,N_15268);
xor U16926 (N_16926,N_15385,N_12811);
nand U16927 (N_16927,N_15209,N_13053);
nand U16928 (N_16928,N_14582,N_13636);
or U16929 (N_16929,N_14818,N_14096);
xnor U16930 (N_16930,N_13629,N_15269);
or U16931 (N_16931,N_14724,N_14669);
xnor U16932 (N_16932,N_13999,N_14152);
nand U16933 (N_16933,N_13253,N_14559);
xor U16934 (N_16934,N_14595,N_14676);
nor U16935 (N_16935,N_14336,N_14041);
xor U16936 (N_16936,N_15562,N_14764);
xor U16937 (N_16937,N_12509,N_12694);
xor U16938 (N_16938,N_15210,N_15610);
nand U16939 (N_16939,N_15129,N_12613);
or U16940 (N_16940,N_12676,N_14213);
xor U16941 (N_16941,N_14743,N_14593);
and U16942 (N_16942,N_15393,N_13758);
nand U16943 (N_16943,N_15480,N_15295);
or U16944 (N_16944,N_15332,N_14186);
nor U16945 (N_16945,N_14722,N_14721);
and U16946 (N_16946,N_14610,N_13810);
xor U16947 (N_16947,N_15298,N_14082);
and U16948 (N_16948,N_15379,N_14781);
nand U16949 (N_16949,N_13417,N_15619);
xnor U16950 (N_16950,N_14281,N_14713);
and U16951 (N_16951,N_13612,N_12908);
nor U16952 (N_16952,N_14436,N_14378);
nor U16953 (N_16953,N_14680,N_14515);
nand U16954 (N_16954,N_12901,N_14409);
or U16955 (N_16955,N_14858,N_13474);
xnor U16956 (N_16956,N_13841,N_12738);
and U16957 (N_16957,N_14438,N_12737);
xnor U16958 (N_16958,N_15107,N_15486);
nand U16959 (N_16959,N_14398,N_15611);
nand U16960 (N_16960,N_12874,N_14823);
nor U16961 (N_16961,N_13395,N_15533);
nand U16962 (N_16962,N_14600,N_14458);
xnor U16963 (N_16963,N_13005,N_12607);
xnor U16964 (N_16964,N_13437,N_13871);
xor U16965 (N_16965,N_15148,N_13820);
and U16966 (N_16966,N_15277,N_14672);
nand U16967 (N_16967,N_13380,N_14422);
or U16968 (N_16968,N_14282,N_14389);
nor U16969 (N_16969,N_15056,N_14857);
and U16970 (N_16970,N_14645,N_13409);
and U16971 (N_16971,N_14496,N_14410);
nor U16972 (N_16972,N_13232,N_14875);
and U16973 (N_16973,N_13031,N_13826);
xor U16974 (N_16974,N_13648,N_14671);
or U16975 (N_16975,N_13165,N_13193);
or U16976 (N_16976,N_13124,N_13176);
nor U16977 (N_16977,N_12931,N_12647);
nor U16978 (N_16978,N_13876,N_14540);
or U16979 (N_16979,N_15216,N_14539);
nand U16980 (N_16980,N_14505,N_15451);
nand U16981 (N_16981,N_15354,N_14064);
nor U16982 (N_16982,N_12503,N_12750);
nor U16983 (N_16983,N_13595,N_14302);
and U16984 (N_16984,N_14491,N_14907);
nor U16985 (N_16985,N_13708,N_12523);
or U16986 (N_16986,N_12666,N_13596);
nand U16987 (N_16987,N_14885,N_14275);
and U16988 (N_16988,N_15387,N_13324);
nor U16989 (N_16989,N_15250,N_12600);
nor U16990 (N_16990,N_15334,N_13133);
and U16991 (N_16991,N_14868,N_13007);
nand U16992 (N_16992,N_14537,N_14914);
or U16993 (N_16993,N_13598,N_13399);
xor U16994 (N_16994,N_12903,N_15076);
or U16995 (N_16995,N_14553,N_14681);
xor U16996 (N_16996,N_14806,N_12629);
nor U16997 (N_16997,N_13468,N_15362);
or U16998 (N_16998,N_14941,N_13613);
nand U16999 (N_16999,N_13673,N_14843);
and U17000 (N_17000,N_13148,N_13149);
nand U17001 (N_17001,N_15285,N_12922);
or U17002 (N_17002,N_13214,N_13788);
and U17003 (N_17003,N_15000,N_13207);
nand U17004 (N_17004,N_12531,N_14126);
nor U17005 (N_17005,N_13271,N_14607);
or U17006 (N_17006,N_14536,N_15599);
or U17007 (N_17007,N_15286,N_14429);
nor U17008 (N_17008,N_15494,N_14815);
or U17009 (N_17009,N_15008,N_12609);
xnor U17010 (N_17010,N_12850,N_14919);
nand U17011 (N_17011,N_14759,N_14475);
nor U17012 (N_17012,N_14042,N_13570);
and U17013 (N_17013,N_14720,N_13013);
xor U17014 (N_17014,N_14144,N_13028);
and U17015 (N_17015,N_15035,N_12808);
nor U17016 (N_17016,N_15553,N_14623);
and U17017 (N_17017,N_15287,N_12728);
nand U17018 (N_17018,N_13734,N_15199);
nand U17019 (N_17019,N_15012,N_14185);
or U17020 (N_17020,N_14354,N_14963);
or U17021 (N_17021,N_14379,N_14768);
xor U17022 (N_17022,N_13439,N_15201);
nand U17023 (N_17023,N_15456,N_13245);
xor U17024 (N_17024,N_13223,N_13551);
or U17025 (N_17025,N_14433,N_13656);
or U17026 (N_17026,N_14688,N_13930);
xnor U17027 (N_17027,N_14404,N_13705);
xnor U17028 (N_17028,N_13828,N_13751);
xnor U17029 (N_17029,N_13425,N_12594);
or U17030 (N_17030,N_14612,N_14218);
nand U17031 (N_17031,N_15377,N_14269);
nor U17032 (N_17032,N_13141,N_14702);
nor U17033 (N_17033,N_14116,N_14270);
or U17034 (N_17034,N_14255,N_15555);
xor U17035 (N_17035,N_15214,N_13805);
nor U17036 (N_17036,N_13605,N_14289);
or U17037 (N_17037,N_12973,N_13693);
or U17038 (N_17038,N_13664,N_14462);
or U17039 (N_17039,N_12913,N_13889);
xor U17040 (N_17040,N_14045,N_14784);
nand U17041 (N_17041,N_14811,N_13501);
xnor U17042 (N_17042,N_13714,N_14117);
or U17043 (N_17043,N_12561,N_14979);
or U17044 (N_17044,N_15428,N_13315);
nor U17045 (N_17045,N_15568,N_12754);
nor U17046 (N_17046,N_12793,N_12848);
nand U17047 (N_17047,N_13747,N_12580);
xor U17048 (N_17048,N_15168,N_13259);
xor U17049 (N_17049,N_12562,N_13084);
or U17050 (N_17050,N_13020,N_12847);
and U17051 (N_17051,N_15493,N_13527);
and U17052 (N_17052,N_13529,N_15215);
or U17053 (N_17053,N_13634,N_14630);
xnor U17054 (N_17054,N_15481,N_12829);
xnor U17055 (N_17055,N_15222,N_15496);
or U17056 (N_17056,N_12979,N_14093);
nor U17057 (N_17057,N_13172,N_12533);
nor U17058 (N_17058,N_14198,N_15471);
or U17059 (N_17059,N_14583,N_13194);
and U17060 (N_17060,N_13361,N_13174);
nor U17061 (N_17061,N_12820,N_14043);
nand U17062 (N_17062,N_12876,N_14999);
xor U17063 (N_17063,N_14209,N_12862);
xor U17064 (N_17064,N_13678,N_12567);
or U17065 (N_17065,N_14388,N_13679);
nand U17066 (N_17066,N_14895,N_15065);
nor U17067 (N_17067,N_13049,N_14803);
nand U17068 (N_17068,N_13563,N_15145);
nand U17069 (N_17069,N_14220,N_15303);
and U17070 (N_17070,N_13639,N_14568);
or U17071 (N_17071,N_15125,N_15561);
or U17072 (N_17072,N_15560,N_12537);
nor U17073 (N_17073,N_15543,N_14383);
or U17074 (N_17074,N_13471,N_15087);
xor U17075 (N_17075,N_14620,N_15403);
xnor U17076 (N_17076,N_13534,N_14367);
xor U17077 (N_17077,N_14928,N_12958);
or U17078 (N_17078,N_14072,N_12723);
and U17079 (N_17079,N_13922,N_13887);
xnor U17080 (N_17080,N_14973,N_14586);
nor U17081 (N_17081,N_13528,N_14938);
and U17082 (N_17082,N_12590,N_14898);
nor U17083 (N_17083,N_14036,N_14542);
and U17084 (N_17084,N_15621,N_13085);
nor U17085 (N_17085,N_13822,N_14621);
nor U17086 (N_17086,N_14171,N_15364);
nand U17087 (N_17087,N_15461,N_14067);
xor U17088 (N_17088,N_13042,N_12548);
and U17089 (N_17089,N_15479,N_15425);
xor U17090 (N_17090,N_15068,N_13867);
and U17091 (N_17091,N_14206,N_15184);
xnor U17092 (N_17092,N_13419,N_12502);
nand U17093 (N_17093,N_14000,N_15341);
nor U17094 (N_17094,N_14345,N_12588);
or U17095 (N_17095,N_13109,N_15031);
or U17096 (N_17096,N_13589,N_12875);
xnor U17097 (N_17097,N_13159,N_13621);
nor U17098 (N_17098,N_13499,N_13692);
xnor U17099 (N_17099,N_13910,N_12555);
nor U17100 (N_17100,N_12620,N_15359);
or U17101 (N_17101,N_14758,N_15485);
or U17102 (N_17102,N_12508,N_12795);
or U17103 (N_17103,N_15538,N_13003);
and U17104 (N_17104,N_14492,N_13689);
xor U17105 (N_17105,N_13965,N_13390);
and U17106 (N_17106,N_14301,N_13199);
nor U17107 (N_17107,N_13480,N_13497);
nand U17108 (N_17108,N_14644,N_15581);
nor U17109 (N_17109,N_15237,N_13653);
nor U17110 (N_17110,N_14352,N_13115);
and U17111 (N_17111,N_14014,N_12905);
or U17112 (N_17112,N_13848,N_14997);
nand U17113 (N_17113,N_14197,N_13443);
xor U17114 (N_17114,N_13424,N_14323);
nor U17115 (N_17115,N_13370,N_15521);
nand U17116 (N_17116,N_14513,N_14063);
nor U17117 (N_17117,N_15195,N_12782);
nor U17118 (N_17118,N_14237,N_13952);
and U17119 (N_17119,N_14330,N_14608);
nand U17120 (N_17120,N_15351,N_13326);
or U17121 (N_17121,N_15067,N_14100);
nand U17122 (N_17122,N_13800,N_13757);
nand U17123 (N_17123,N_14424,N_13707);
nor U17124 (N_17124,N_12673,N_14025);
nor U17125 (N_17125,N_14753,N_12810);
xnor U17126 (N_17126,N_14076,N_15140);
or U17127 (N_17127,N_13792,N_12731);
nor U17128 (N_17128,N_14238,N_12777);
nand U17129 (N_17129,N_14925,N_15424);
nor U17130 (N_17130,N_14300,N_14098);
nand U17131 (N_17131,N_14256,N_13559);
xnor U17132 (N_17132,N_15078,N_14273);
xnor U17133 (N_17133,N_14010,N_13391);
and U17134 (N_17134,N_13954,N_15224);
or U17135 (N_17135,N_15108,N_15047);
nor U17136 (N_17136,N_13009,N_14008);
or U17137 (N_17137,N_14693,N_15011);
nor U17138 (N_17138,N_13431,N_13056);
or U17139 (N_17139,N_15029,N_12866);
nand U17140 (N_17140,N_14617,N_12989);
xnor U17141 (N_17141,N_15190,N_15064);
and U17142 (N_17142,N_13498,N_14584);
or U17143 (N_17143,N_13680,N_14239);
or U17144 (N_17144,N_13745,N_12735);
nor U17145 (N_17145,N_13448,N_13506);
nor U17146 (N_17146,N_13659,N_13684);
nor U17147 (N_17147,N_14679,N_15552);
or U17148 (N_17148,N_13677,N_13565);
or U17149 (N_17149,N_13002,N_14431);
xor U17150 (N_17150,N_13384,N_15436);
or U17151 (N_17151,N_12709,N_14139);
nand U17152 (N_17152,N_13740,N_13089);
nand U17153 (N_17153,N_13225,N_13989);
and U17154 (N_17154,N_13832,N_15477);
and U17155 (N_17155,N_14376,N_13442);
or U17156 (N_17156,N_13749,N_15048);
and U17157 (N_17157,N_14767,N_15001);
xnor U17158 (N_17158,N_15529,N_13668);
xor U17159 (N_17159,N_12936,N_14549);
nor U17160 (N_17160,N_14946,N_15119);
or U17161 (N_17161,N_13346,N_14550);
nor U17162 (N_17162,N_12685,N_14038);
nor U17163 (N_17163,N_14873,N_13181);
and U17164 (N_17164,N_15575,N_14030);
or U17165 (N_17165,N_13220,N_14807);
or U17166 (N_17166,N_14625,N_13655);
and U17167 (N_17167,N_12960,N_13861);
and U17168 (N_17168,N_15096,N_14131);
nand U17169 (N_17169,N_13215,N_14616);
nand U17170 (N_17170,N_14318,N_15192);
xnor U17171 (N_17171,N_12651,N_14905);
nand U17172 (N_17172,N_14322,N_14937);
xor U17173 (N_17173,N_15165,N_14199);
and U17174 (N_17174,N_14996,N_13804);
xor U17175 (N_17175,N_14661,N_13547);
and U17176 (N_17176,N_15092,N_14477);
or U17177 (N_17177,N_12563,N_13427);
and U17178 (N_17178,N_12801,N_13929);
nand U17179 (N_17179,N_13985,N_13029);
and U17180 (N_17180,N_14200,N_13068);
nor U17181 (N_17181,N_14633,N_14441);
nand U17182 (N_17182,N_14854,N_13203);
or U17183 (N_17183,N_12560,N_14638);
or U17184 (N_17184,N_13093,N_13500);
or U17185 (N_17185,N_13289,N_14316);
and U17186 (N_17186,N_12774,N_14628);
or U17187 (N_17187,N_12713,N_14832);
nand U17188 (N_17188,N_14658,N_15223);
and U17189 (N_17189,N_15199,N_13897);
nor U17190 (N_17190,N_13674,N_12974);
or U17191 (N_17191,N_13720,N_14796);
or U17192 (N_17192,N_13883,N_15501);
nand U17193 (N_17193,N_13564,N_15128);
or U17194 (N_17194,N_14734,N_13555);
xnor U17195 (N_17195,N_14332,N_15124);
or U17196 (N_17196,N_12968,N_14345);
xor U17197 (N_17197,N_13022,N_14549);
nor U17198 (N_17198,N_14889,N_13620);
nor U17199 (N_17199,N_13130,N_13014);
nand U17200 (N_17200,N_12972,N_15494);
nor U17201 (N_17201,N_12672,N_14765);
xor U17202 (N_17202,N_13885,N_14703);
nand U17203 (N_17203,N_13847,N_15412);
or U17204 (N_17204,N_13600,N_12858);
and U17205 (N_17205,N_12846,N_12542);
or U17206 (N_17206,N_12909,N_14482);
and U17207 (N_17207,N_13504,N_13371);
nand U17208 (N_17208,N_13129,N_14257);
xor U17209 (N_17209,N_14802,N_15170);
or U17210 (N_17210,N_14186,N_13805);
nand U17211 (N_17211,N_12712,N_14496);
xnor U17212 (N_17212,N_15330,N_13880);
or U17213 (N_17213,N_13860,N_12694);
nor U17214 (N_17214,N_13736,N_15498);
nand U17215 (N_17215,N_14196,N_13111);
and U17216 (N_17216,N_14503,N_13872);
and U17217 (N_17217,N_13439,N_15344);
xnor U17218 (N_17218,N_14360,N_15134);
nand U17219 (N_17219,N_15447,N_15091);
and U17220 (N_17220,N_14782,N_14116);
or U17221 (N_17221,N_14605,N_14579);
nor U17222 (N_17222,N_14934,N_13002);
or U17223 (N_17223,N_14475,N_14001);
xor U17224 (N_17224,N_13714,N_14294);
nand U17225 (N_17225,N_12721,N_14366);
nand U17226 (N_17226,N_15302,N_13719);
or U17227 (N_17227,N_14820,N_13193);
and U17228 (N_17228,N_14951,N_12630);
nand U17229 (N_17229,N_12514,N_14554);
nand U17230 (N_17230,N_12577,N_15476);
nand U17231 (N_17231,N_12729,N_15273);
or U17232 (N_17232,N_14228,N_14643);
nor U17233 (N_17233,N_13301,N_14577);
nor U17234 (N_17234,N_13333,N_13290);
and U17235 (N_17235,N_13399,N_14082);
nor U17236 (N_17236,N_13969,N_15542);
nor U17237 (N_17237,N_15574,N_14423);
nand U17238 (N_17238,N_13609,N_15344);
and U17239 (N_17239,N_12691,N_13032);
and U17240 (N_17240,N_13408,N_15493);
nor U17241 (N_17241,N_13256,N_14367);
and U17242 (N_17242,N_12624,N_15492);
nand U17243 (N_17243,N_14286,N_15302);
or U17244 (N_17244,N_14977,N_12820);
nor U17245 (N_17245,N_13487,N_13014);
or U17246 (N_17246,N_15242,N_15076);
xor U17247 (N_17247,N_15599,N_13510);
and U17248 (N_17248,N_14578,N_15208);
and U17249 (N_17249,N_15492,N_14225);
and U17250 (N_17250,N_14728,N_15250);
nor U17251 (N_17251,N_15569,N_13572);
or U17252 (N_17252,N_13524,N_15297);
nand U17253 (N_17253,N_12848,N_13674);
nor U17254 (N_17254,N_13973,N_13722);
or U17255 (N_17255,N_15168,N_14460);
nand U17256 (N_17256,N_14234,N_12826);
and U17257 (N_17257,N_12570,N_13906);
xnor U17258 (N_17258,N_15504,N_14398);
and U17259 (N_17259,N_14131,N_13908);
nand U17260 (N_17260,N_13516,N_14913);
or U17261 (N_17261,N_13540,N_14713);
nor U17262 (N_17262,N_13261,N_13723);
and U17263 (N_17263,N_15032,N_12656);
nor U17264 (N_17264,N_13574,N_14199);
xor U17265 (N_17265,N_14542,N_12671);
or U17266 (N_17266,N_14921,N_14813);
or U17267 (N_17267,N_14031,N_12881);
or U17268 (N_17268,N_12519,N_13180);
nand U17269 (N_17269,N_13862,N_12883);
xnor U17270 (N_17270,N_14276,N_14709);
nand U17271 (N_17271,N_13930,N_14256);
nand U17272 (N_17272,N_13309,N_14582);
xor U17273 (N_17273,N_14120,N_14208);
nand U17274 (N_17274,N_15591,N_13295);
and U17275 (N_17275,N_14019,N_14105);
and U17276 (N_17276,N_14728,N_15110);
and U17277 (N_17277,N_15041,N_15562);
nor U17278 (N_17278,N_15433,N_15273);
nor U17279 (N_17279,N_13290,N_12552);
xnor U17280 (N_17280,N_15483,N_13451);
xor U17281 (N_17281,N_14497,N_12518);
xor U17282 (N_17282,N_13258,N_13604);
and U17283 (N_17283,N_13271,N_14968);
nor U17284 (N_17284,N_13061,N_13393);
or U17285 (N_17285,N_13978,N_14923);
and U17286 (N_17286,N_13790,N_14331);
xor U17287 (N_17287,N_13883,N_13225);
and U17288 (N_17288,N_14740,N_13202);
nand U17289 (N_17289,N_12607,N_14721);
and U17290 (N_17290,N_15395,N_15221);
nor U17291 (N_17291,N_13598,N_13005);
nor U17292 (N_17292,N_14696,N_15164);
or U17293 (N_17293,N_12631,N_12552);
and U17294 (N_17294,N_15572,N_15483);
xor U17295 (N_17295,N_12881,N_14362);
nor U17296 (N_17296,N_14356,N_12699);
and U17297 (N_17297,N_14146,N_14677);
and U17298 (N_17298,N_14792,N_14188);
or U17299 (N_17299,N_14887,N_15384);
nand U17300 (N_17300,N_13851,N_13457);
nor U17301 (N_17301,N_14834,N_12546);
and U17302 (N_17302,N_13887,N_15218);
nor U17303 (N_17303,N_13498,N_15462);
nor U17304 (N_17304,N_15372,N_15442);
nor U17305 (N_17305,N_13233,N_12871);
xor U17306 (N_17306,N_14398,N_15241);
nor U17307 (N_17307,N_13993,N_13011);
nor U17308 (N_17308,N_13982,N_14172);
nand U17309 (N_17309,N_12627,N_15374);
and U17310 (N_17310,N_12971,N_15545);
xor U17311 (N_17311,N_14037,N_13608);
or U17312 (N_17312,N_14800,N_13242);
nand U17313 (N_17313,N_15315,N_13134);
nand U17314 (N_17314,N_15222,N_12815);
nand U17315 (N_17315,N_15548,N_13140);
and U17316 (N_17316,N_14400,N_15621);
nor U17317 (N_17317,N_13071,N_13554);
and U17318 (N_17318,N_12652,N_14710);
xor U17319 (N_17319,N_14876,N_13124);
nand U17320 (N_17320,N_13063,N_14790);
nand U17321 (N_17321,N_12632,N_13505);
or U17322 (N_17322,N_12758,N_14436);
and U17323 (N_17323,N_14081,N_12802);
xnor U17324 (N_17324,N_15305,N_13802);
nor U17325 (N_17325,N_12544,N_14787);
and U17326 (N_17326,N_12612,N_12879);
or U17327 (N_17327,N_15613,N_15010);
xor U17328 (N_17328,N_14350,N_13458);
xnor U17329 (N_17329,N_14783,N_15448);
and U17330 (N_17330,N_14441,N_13787);
nor U17331 (N_17331,N_15328,N_13703);
and U17332 (N_17332,N_14264,N_12967);
nand U17333 (N_17333,N_15570,N_14990);
nor U17334 (N_17334,N_12589,N_13611);
nor U17335 (N_17335,N_14880,N_14338);
nand U17336 (N_17336,N_13910,N_12776);
or U17337 (N_17337,N_13797,N_14133);
or U17338 (N_17338,N_14730,N_13249);
nor U17339 (N_17339,N_15249,N_14375);
or U17340 (N_17340,N_13300,N_12820);
nand U17341 (N_17341,N_12866,N_14471);
xor U17342 (N_17342,N_14629,N_15461);
nand U17343 (N_17343,N_15456,N_15135);
and U17344 (N_17344,N_13170,N_13677);
xnor U17345 (N_17345,N_15452,N_13025);
xor U17346 (N_17346,N_14285,N_13817);
nor U17347 (N_17347,N_12713,N_15175);
or U17348 (N_17348,N_15202,N_14987);
xor U17349 (N_17349,N_14014,N_15609);
xnor U17350 (N_17350,N_15432,N_14348);
nand U17351 (N_17351,N_14708,N_15168);
nand U17352 (N_17352,N_14502,N_13507);
xor U17353 (N_17353,N_13539,N_13162);
or U17354 (N_17354,N_14220,N_15259);
xor U17355 (N_17355,N_15503,N_13262);
nand U17356 (N_17356,N_14857,N_13924);
and U17357 (N_17357,N_14923,N_15571);
and U17358 (N_17358,N_12797,N_15312);
xor U17359 (N_17359,N_15509,N_15515);
nor U17360 (N_17360,N_14706,N_13729);
and U17361 (N_17361,N_15264,N_13199);
xor U17362 (N_17362,N_15623,N_14477);
nand U17363 (N_17363,N_12801,N_14490);
xor U17364 (N_17364,N_12723,N_15517);
or U17365 (N_17365,N_12735,N_13699);
and U17366 (N_17366,N_14346,N_14440);
xor U17367 (N_17367,N_13828,N_15099);
nand U17368 (N_17368,N_13737,N_14398);
xnor U17369 (N_17369,N_15616,N_15301);
or U17370 (N_17370,N_13404,N_13007);
and U17371 (N_17371,N_15552,N_14958);
nor U17372 (N_17372,N_15386,N_13408);
nand U17373 (N_17373,N_13779,N_14285);
nor U17374 (N_17374,N_13208,N_15231);
xor U17375 (N_17375,N_13104,N_14607);
and U17376 (N_17376,N_12669,N_13989);
nor U17377 (N_17377,N_13697,N_15062);
or U17378 (N_17378,N_13732,N_13046);
nand U17379 (N_17379,N_12901,N_13895);
xnor U17380 (N_17380,N_14611,N_14651);
or U17381 (N_17381,N_14123,N_13039);
or U17382 (N_17382,N_12592,N_14483);
and U17383 (N_17383,N_14810,N_13984);
and U17384 (N_17384,N_13721,N_14127);
nor U17385 (N_17385,N_15315,N_12629);
or U17386 (N_17386,N_12713,N_14846);
nand U17387 (N_17387,N_14123,N_13090);
nand U17388 (N_17388,N_13164,N_13953);
or U17389 (N_17389,N_15032,N_13099);
xor U17390 (N_17390,N_12758,N_14325);
nand U17391 (N_17391,N_13174,N_13492);
or U17392 (N_17392,N_13141,N_12787);
nor U17393 (N_17393,N_12761,N_12767);
nand U17394 (N_17394,N_13417,N_13573);
xnor U17395 (N_17395,N_13942,N_12642);
and U17396 (N_17396,N_15439,N_12729);
xnor U17397 (N_17397,N_13557,N_14751);
nor U17398 (N_17398,N_12889,N_13828);
nand U17399 (N_17399,N_13268,N_14154);
and U17400 (N_17400,N_14013,N_14135);
and U17401 (N_17401,N_14578,N_14515);
and U17402 (N_17402,N_13716,N_13610);
nor U17403 (N_17403,N_12655,N_14150);
nand U17404 (N_17404,N_12583,N_15415);
or U17405 (N_17405,N_14409,N_14979);
or U17406 (N_17406,N_12959,N_15266);
nand U17407 (N_17407,N_14205,N_14929);
and U17408 (N_17408,N_12756,N_15130);
and U17409 (N_17409,N_13001,N_14157);
and U17410 (N_17410,N_14482,N_12735);
or U17411 (N_17411,N_15129,N_12565);
and U17412 (N_17412,N_12765,N_12883);
nor U17413 (N_17413,N_14508,N_13487);
nand U17414 (N_17414,N_14649,N_13862);
nand U17415 (N_17415,N_14710,N_12559);
xnor U17416 (N_17416,N_13679,N_14613);
nor U17417 (N_17417,N_12893,N_15349);
and U17418 (N_17418,N_13022,N_13641);
nor U17419 (N_17419,N_15349,N_14417);
and U17420 (N_17420,N_13451,N_15289);
nand U17421 (N_17421,N_13638,N_14259);
nor U17422 (N_17422,N_12600,N_15481);
or U17423 (N_17423,N_14552,N_15506);
nand U17424 (N_17424,N_14913,N_13013);
xor U17425 (N_17425,N_14253,N_14715);
and U17426 (N_17426,N_12861,N_13198);
and U17427 (N_17427,N_14099,N_15155);
and U17428 (N_17428,N_13527,N_12726);
nand U17429 (N_17429,N_15310,N_14647);
nand U17430 (N_17430,N_13472,N_12572);
and U17431 (N_17431,N_13029,N_14346);
xor U17432 (N_17432,N_13050,N_14203);
and U17433 (N_17433,N_15177,N_13703);
nand U17434 (N_17434,N_14512,N_14166);
xnor U17435 (N_17435,N_13881,N_12551);
and U17436 (N_17436,N_13822,N_14773);
or U17437 (N_17437,N_13433,N_13158);
or U17438 (N_17438,N_14694,N_14623);
or U17439 (N_17439,N_12605,N_13309);
nor U17440 (N_17440,N_15609,N_14871);
xor U17441 (N_17441,N_14231,N_13948);
nand U17442 (N_17442,N_13276,N_15230);
and U17443 (N_17443,N_13408,N_13465);
or U17444 (N_17444,N_15479,N_12985);
nand U17445 (N_17445,N_15001,N_15594);
or U17446 (N_17446,N_15555,N_14905);
nand U17447 (N_17447,N_13898,N_15607);
nand U17448 (N_17448,N_12827,N_12811);
or U17449 (N_17449,N_15413,N_12611);
xor U17450 (N_17450,N_15414,N_15049);
nand U17451 (N_17451,N_14290,N_14207);
nand U17452 (N_17452,N_15540,N_12876);
nand U17453 (N_17453,N_15090,N_13166);
nand U17454 (N_17454,N_12755,N_14416);
nand U17455 (N_17455,N_14036,N_14061);
nor U17456 (N_17456,N_12739,N_13588);
and U17457 (N_17457,N_13543,N_14040);
xnor U17458 (N_17458,N_13690,N_14470);
nand U17459 (N_17459,N_12739,N_13986);
or U17460 (N_17460,N_14664,N_12869);
and U17461 (N_17461,N_15455,N_13472);
nand U17462 (N_17462,N_12758,N_14723);
or U17463 (N_17463,N_15482,N_13934);
xnor U17464 (N_17464,N_13872,N_13721);
or U17465 (N_17465,N_13176,N_15530);
xnor U17466 (N_17466,N_13214,N_14149);
nor U17467 (N_17467,N_13732,N_14702);
and U17468 (N_17468,N_14757,N_14709);
nand U17469 (N_17469,N_13833,N_14995);
or U17470 (N_17470,N_14447,N_13039);
nor U17471 (N_17471,N_13335,N_13033);
and U17472 (N_17472,N_13236,N_13495);
nor U17473 (N_17473,N_12557,N_14784);
nand U17474 (N_17474,N_12633,N_15217);
or U17475 (N_17475,N_14466,N_15160);
xor U17476 (N_17476,N_13928,N_13882);
xor U17477 (N_17477,N_13560,N_14625);
xnor U17478 (N_17478,N_15332,N_15388);
or U17479 (N_17479,N_14392,N_15358);
nand U17480 (N_17480,N_15577,N_13826);
and U17481 (N_17481,N_13736,N_13950);
and U17482 (N_17482,N_12671,N_13833);
or U17483 (N_17483,N_14132,N_13715);
xor U17484 (N_17484,N_15083,N_14053);
nand U17485 (N_17485,N_15555,N_14489);
xnor U17486 (N_17486,N_12697,N_15033);
and U17487 (N_17487,N_12887,N_13412);
nor U17488 (N_17488,N_12743,N_14713);
or U17489 (N_17489,N_14855,N_12886);
nor U17490 (N_17490,N_12863,N_13944);
or U17491 (N_17491,N_13570,N_13664);
nand U17492 (N_17492,N_15491,N_13018);
nor U17493 (N_17493,N_12561,N_15249);
nand U17494 (N_17494,N_14343,N_12953);
xnor U17495 (N_17495,N_12752,N_14459);
xnor U17496 (N_17496,N_14419,N_13025);
and U17497 (N_17497,N_15329,N_13119);
xnor U17498 (N_17498,N_13712,N_14373);
and U17499 (N_17499,N_15472,N_15243);
or U17500 (N_17500,N_14386,N_12736);
xnor U17501 (N_17501,N_14545,N_12768);
nand U17502 (N_17502,N_13496,N_12535);
and U17503 (N_17503,N_13201,N_13426);
or U17504 (N_17504,N_12648,N_12977);
nand U17505 (N_17505,N_14455,N_13993);
nand U17506 (N_17506,N_15349,N_13578);
xor U17507 (N_17507,N_15243,N_12748);
nand U17508 (N_17508,N_13503,N_14113);
and U17509 (N_17509,N_14474,N_14820);
and U17510 (N_17510,N_14407,N_13112);
and U17511 (N_17511,N_13821,N_13691);
xor U17512 (N_17512,N_15460,N_15330);
and U17513 (N_17513,N_13265,N_13744);
and U17514 (N_17514,N_14242,N_14722);
xnor U17515 (N_17515,N_13888,N_12944);
nor U17516 (N_17516,N_12966,N_13319);
xor U17517 (N_17517,N_15139,N_14281);
and U17518 (N_17518,N_14268,N_13476);
or U17519 (N_17519,N_13886,N_14596);
nand U17520 (N_17520,N_14541,N_15115);
or U17521 (N_17521,N_14411,N_13726);
or U17522 (N_17522,N_12648,N_14235);
nor U17523 (N_17523,N_13582,N_13991);
and U17524 (N_17524,N_12688,N_13140);
nor U17525 (N_17525,N_14342,N_15005);
nor U17526 (N_17526,N_12567,N_13837);
xnor U17527 (N_17527,N_14412,N_13750);
or U17528 (N_17528,N_15337,N_13054);
nand U17529 (N_17529,N_13691,N_12783);
xor U17530 (N_17530,N_14903,N_14505);
nor U17531 (N_17531,N_12667,N_12992);
nand U17532 (N_17532,N_15572,N_14749);
or U17533 (N_17533,N_13999,N_13796);
nand U17534 (N_17534,N_12657,N_15298);
nor U17535 (N_17535,N_13846,N_14429);
nor U17536 (N_17536,N_14065,N_14657);
nor U17537 (N_17537,N_14666,N_14353);
nor U17538 (N_17538,N_13369,N_12949);
nor U17539 (N_17539,N_13842,N_13640);
or U17540 (N_17540,N_13096,N_13915);
nand U17541 (N_17541,N_13654,N_12701);
nand U17542 (N_17542,N_14959,N_13406);
nor U17543 (N_17543,N_15057,N_14422);
xor U17544 (N_17544,N_14816,N_14831);
and U17545 (N_17545,N_14903,N_15344);
and U17546 (N_17546,N_14577,N_15333);
xor U17547 (N_17547,N_13340,N_12612);
and U17548 (N_17548,N_13141,N_12934);
xnor U17549 (N_17549,N_13765,N_14577);
xor U17550 (N_17550,N_14555,N_15035);
xor U17551 (N_17551,N_12503,N_13693);
nand U17552 (N_17552,N_13792,N_12725);
nor U17553 (N_17553,N_15062,N_14806);
nand U17554 (N_17554,N_14514,N_14250);
nand U17555 (N_17555,N_13176,N_13282);
xor U17556 (N_17556,N_12844,N_13548);
and U17557 (N_17557,N_15357,N_13863);
nor U17558 (N_17558,N_15194,N_13921);
nor U17559 (N_17559,N_15132,N_14530);
and U17560 (N_17560,N_13515,N_14728);
nor U17561 (N_17561,N_14545,N_13860);
and U17562 (N_17562,N_14935,N_15008);
nand U17563 (N_17563,N_13246,N_14157);
nor U17564 (N_17564,N_15286,N_14461);
xor U17565 (N_17565,N_14402,N_13586);
and U17566 (N_17566,N_13829,N_13873);
and U17567 (N_17567,N_15618,N_14185);
or U17568 (N_17568,N_15024,N_12689);
or U17569 (N_17569,N_14997,N_13201);
nand U17570 (N_17570,N_14144,N_13034);
nor U17571 (N_17571,N_15159,N_13525);
nand U17572 (N_17572,N_13827,N_14613);
and U17573 (N_17573,N_12515,N_13462);
xor U17574 (N_17574,N_13256,N_14649);
nor U17575 (N_17575,N_15319,N_14920);
or U17576 (N_17576,N_13940,N_14697);
and U17577 (N_17577,N_14726,N_12744);
or U17578 (N_17578,N_12987,N_13213);
or U17579 (N_17579,N_15214,N_12726);
and U17580 (N_17580,N_14402,N_14410);
xnor U17581 (N_17581,N_13958,N_13872);
or U17582 (N_17582,N_13734,N_13110);
or U17583 (N_17583,N_14978,N_12810);
xnor U17584 (N_17584,N_15223,N_13896);
and U17585 (N_17585,N_15184,N_13348);
xnor U17586 (N_17586,N_12829,N_13799);
and U17587 (N_17587,N_14122,N_15468);
xor U17588 (N_17588,N_12898,N_13205);
and U17589 (N_17589,N_12904,N_12750);
and U17590 (N_17590,N_15044,N_14985);
nor U17591 (N_17591,N_12748,N_13025);
and U17592 (N_17592,N_13518,N_13474);
nand U17593 (N_17593,N_13110,N_15266);
nor U17594 (N_17594,N_14033,N_12591);
or U17595 (N_17595,N_13986,N_12715);
and U17596 (N_17596,N_14948,N_14861);
xor U17597 (N_17597,N_13388,N_12852);
nor U17598 (N_17598,N_14564,N_14612);
xnor U17599 (N_17599,N_14982,N_14508);
xor U17600 (N_17600,N_14408,N_12952);
nor U17601 (N_17601,N_15038,N_14794);
nor U17602 (N_17602,N_14697,N_12557);
and U17603 (N_17603,N_13466,N_14827);
or U17604 (N_17604,N_14802,N_14496);
or U17605 (N_17605,N_14783,N_13245);
xnor U17606 (N_17606,N_14874,N_14554);
or U17607 (N_17607,N_13607,N_13887);
nand U17608 (N_17608,N_15193,N_14103);
xor U17609 (N_17609,N_14847,N_13237);
xnor U17610 (N_17610,N_14481,N_13190);
xor U17611 (N_17611,N_14861,N_14028);
xnor U17612 (N_17612,N_14828,N_15100);
nor U17613 (N_17613,N_15277,N_15542);
nand U17614 (N_17614,N_13095,N_14082);
nand U17615 (N_17615,N_15142,N_15024);
xnor U17616 (N_17616,N_12843,N_14423);
and U17617 (N_17617,N_15484,N_14342);
xor U17618 (N_17618,N_13095,N_15228);
nor U17619 (N_17619,N_13029,N_12853);
and U17620 (N_17620,N_15567,N_14418);
xor U17621 (N_17621,N_13985,N_12744);
nand U17622 (N_17622,N_15538,N_13311);
and U17623 (N_17623,N_13033,N_13863);
or U17624 (N_17624,N_13570,N_13382);
or U17625 (N_17625,N_13006,N_15108);
or U17626 (N_17626,N_13737,N_13128);
and U17627 (N_17627,N_13357,N_12701);
nand U17628 (N_17628,N_13573,N_15268);
nand U17629 (N_17629,N_12639,N_14149);
nand U17630 (N_17630,N_15430,N_14942);
or U17631 (N_17631,N_13740,N_13547);
or U17632 (N_17632,N_12608,N_14870);
nand U17633 (N_17633,N_12513,N_13083);
or U17634 (N_17634,N_14848,N_12893);
nand U17635 (N_17635,N_14471,N_13889);
xor U17636 (N_17636,N_14403,N_14159);
nand U17637 (N_17637,N_14448,N_13127);
and U17638 (N_17638,N_15404,N_14768);
and U17639 (N_17639,N_13984,N_12801);
or U17640 (N_17640,N_13438,N_13128);
xnor U17641 (N_17641,N_12763,N_14157);
xor U17642 (N_17642,N_12683,N_13544);
nand U17643 (N_17643,N_12912,N_14781);
nor U17644 (N_17644,N_14078,N_14806);
or U17645 (N_17645,N_14938,N_12764);
and U17646 (N_17646,N_13877,N_14040);
nor U17647 (N_17647,N_14438,N_15127);
or U17648 (N_17648,N_13130,N_12921);
and U17649 (N_17649,N_13102,N_14553);
nand U17650 (N_17650,N_12895,N_15547);
or U17651 (N_17651,N_15442,N_12777);
nor U17652 (N_17652,N_15240,N_12995);
xor U17653 (N_17653,N_14495,N_15120);
nand U17654 (N_17654,N_15340,N_14480);
and U17655 (N_17655,N_13025,N_15004);
and U17656 (N_17656,N_13843,N_13588);
xor U17657 (N_17657,N_14821,N_15449);
or U17658 (N_17658,N_13932,N_14129);
nor U17659 (N_17659,N_15399,N_14136);
and U17660 (N_17660,N_12596,N_14025);
nor U17661 (N_17661,N_13217,N_15485);
and U17662 (N_17662,N_13608,N_14326);
xnor U17663 (N_17663,N_14654,N_14095);
and U17664 (N_17664,N_14820,N_13762);
nor U17665 (N_17665,N_12699,N_13840);
nand U17666 (N_17666,N_13732,N_14926);
nor U17667 (N_17667,N_12896,N_13335);
nand U17668 (N_17668,N_12997,N_14592);
and U17669 (N_17669,N_13607,N_14607);
nand U17670 (N_17670,N_12699,N_15050);
nor U17671 (N_17671,N_13700,N_13919);
or U17672 (N_17672,N_12844,N_12533);
and U17673 (N_17673,N_13549,N_12995);
nor U17674 (N_17674,N_14949,N_13491);
xnor U17675 (N_17675,N_14584,N_15583);
and U17676 (N_17676,N_12720,N_13062);
nand U17677 (N_17677,N_14573,N_14078);
and U17678 (N_17678,N_14879,N_14150);
or U17679 (N_17679,N_13362,N_12676);
nand U17680 (N_17680,N_14338,N_13482);
xnor U17681 (N_17681,N_12898,N_13793);
and U17682 (N_17682,N_14864,N_13500);
nand U17683 (N_17683,N_15003,N_13892);
nor U17684 (N_17684,N_12809,N_14877);
nor U17685 (N_17685,N_13611,N_13267);
nand U17686 (N_17686,N_13029,N_15523);
and U17687 (N_17687,N_13624,N_12821);
xor U17688 (N_17688,N_13354,N_14013);
and U17689 (N_17689,N_14445,N_13284);
xnor U17690 (N_17690,N_14288,N_13358);
or U17691 (N_17691,N_12923,N_15302);
nor U17692 (N_17692,N_13639,N_12672);
nor U17693 (N_17693,N_14778,N_12599);
nand U17694 (N_17694,N_13667,N_14133);
xor U17695 (N_17695,N_13658,N_15386);
or U17696 (N_17696,N_14382,N_13782);
and U17697 (N_17697,N_15137,N_12509);
or U17698 (N_17698,N_12661,N_13360);
or U17699 (N_17699,N_12848,N_15048);
and U17700 (N_17700,N_13935,N_14632);
nor U17701 (N_17701,N_13830,N_14391);
xnor U17702 (N_17702,N_14318,N_13390);
and U17703 (N_17703,N_12813,N_12602);
xor U17704 (N_17704,N_14554,N_15054);
and U17705 (N_17705,N_13272,N_14118);
nand U17706 (N_17706,N_14161,N_13180);
nand U17707 (N_17707,N_15607,N_14348);
nor U17708 (N_17708,N_13875,N_15520);
or U17709 (N_17709,N_13602,N_13266);
nand U17710 (N_17710,N_14192,N_14506);
nor U17711 (N_17711,N_14316,N_15508);
xnor U17712 (N_17712,N_13203,N_14326);
xor U17713 (N_17713,N_13546,N_12637);
xor U17714 (N_17714,N_13127,N_12710);
or U17715 (N_17715,N_14936,N_13126);
or U17716 (N_17716,N_14513,N_15223);
and U17717 (N_17717,N_15512,N_14597);
nor U17718 (N_17718,N_13511,N_13038);
and U17719 (N_17719,N_15409,N_14893);
xor U17720 (N_17720,N_14296,N_13455);
or U17721 (N_17721,N_13270,N_13741);
xor U17722 (N_17722,N_12813,N_14180);
nor U17723 (N_17723,N_12595,N_13530);
nand U17724 (N_17724,N_15113,N_14847);
nor U17725 (N_17725,N_14329,N_13614);
nor U17726 (N_17726,N_14909,N_14574);
nand U17727 (N_17727,N_14132,N_13088);
and U17728 (N_17728,N_14206,N_12554);
nand U17729 (N_17729,N_12760,N_14114);
nor U17730 (N_17730,N_14823,N_14699);
or U17731 (N_17731,N_14948,N_12696);
and U17732 (N_17732,N_12804,N_12632);
or U17733 (N_17733,N_14182,N_14179);
nor U17734 (N_17734,N_12532,N_14670);
nand U17735 (N_17735,N_15497,N_15002);
and U17736 (N_17736,N_12676,N_15536);
nor U17737 (N_17737,N_13717,N_13426);
xor U17738 (N_17738,N_13503,N_12691);
nor U17739 (N_17739,N_14815,N_14848);
and U17740 (N_17740,N_13252,N_14375);
or U17741 (N_17741,N_13997,N_15131);
nand U17742 (N_17742,N_12566,N_15199);
nor U17743 (N_17743,N_15216,N_14210);
nand U17744 (N_17744,N_15234,N_14921);
and U17745 (N_17745,N_14126,N_14885);
xor U17746 (N_17746,N_12678,N_13219);
or U17747 (N_17747,N_15425,N_14499);
nor U17748 (N_17748,N_14358,N_13144);
nor U17749 (N_17749,N_12994,N_13474);
and U17750 (N_17750,N_15196,N_14711);
or U17751 (N_17751,N_13426,N_13134);
nand U17752 (N_17752,N_12762,N_15158);
xnor U17753 (N_17753,N_15198,N_13757);
and U17754 (N_17754,N_13889,N_12611);
and U17755 (N_17755,N_13754,N_14922);
nor U17756 (N_17756,N_13343,N_14450);
xnor U17757 (N_17757,N_14957,N_13018);
nor U17758 (N_17758,N_12549,N_13789);
and U17759 (N_17759,N_13285,N_14578);
or U17760 (N_17760,N_14752,N_12854);
or U17761 (N_17761,N_13137,N_13825);
and U17762 (N_17762,N_12909,N_14925);
nand U17763 (N_17763,N_13845,N_12998);
nor U17764 (N_17764,N_12796,N_15132);
nor U17765 (N_17765,N_15374,N_12609);
xnor U17766 (N_17766,N_14443,N_14541);
and U17767 (N_17767,N_13871,N_14287);
nand U17768 (N_17768,N_14080,N_12821);
and U17769 (N_17769,N_13500,N_14342);
and U17770 (N_17770,N_15300,N_14696);
nand U17771 (N_17771,N_14675,N_15169);
and U17772 (N_17772,N_15308,N_14972);
nor U17773 (N_17773,N_13055,N_14871);
nand U17774 (N_17774,N_15095,N_13044);
nand U17775 (N_17775,N_13501,N_14738);
or U17776 (N_17776,N_12941,N_15047);
xnor U17777 (N_17777,N_13967,N_12627);
xnor U17778 (N_17778,N_13321,N_14725);
xor U17779 (N_17779,N_14473,N_13557);
nor U17780 (N_17780,N_14776,N_14462);
xor U17781 (N_17781,N_14110,N_15170);
nor U17782 (N_17782,N_14485,N_14953);
nand U17783 (N_17783,N_12938,N_15499);
xnor U17784 (N_17784,N_14822,N_13692);
xor U17785 (N_17785,N_14862,N_13398);
and U17786 (N_17786,N_12656,N_12913);
nand U17787 (N_17787,N_12924,N_13329);
nor U17788 (N_17788,N_13171,N_12990);
xor U17789 (N_17789,N_14275,N_13318);
and U17790 (N_17790,N_15570,N_13924);
nand U17791 (N_17791,N_14475,N_14141);
nand U17792 (N_17792,N_13462,N_15016);
or U17793 (N_17793,N_14609,N_12854);
or U17794 (N_17794,N_13722,N_13685);
and U17795 (N_17795,N_13738,N_14106);
nor U17796 (N_17796,N_13993,N_14450);
and U17797 (N_17797,N_14713,N_14752);
nand U17798 (N_17798,N_13378,N_14926);
and U17799 (N_17799,N_13112,N_15614);
nand U17800 (N_17800,N_14522,N_13618);
nor U17801 (N_17801,N_13554,N_15346);
nor U17802 (N_17802,N_15355,N_14397);
nand U17803 (N_17803,N_14957,N_14939);
nand U17804 (N_17804,N_14385,N_14780);
nand U17805 (N_17805,N_14565,N_15075);
or U17806 (N_17806,N_15089,N_13055);
nand U17807 (N_17807,N_14687,N_15552);
xor U17808 (N_17808,N_12560,N_13516);
nor U17809 (N_17809,N_15240,N_15059);
or U17810 (N_17810,N_12635,N_13291);
nand U17811 (N_17811,N_14707,N_15357);
xnor U17812 (N_17812,N_13649,N_12791);
or U17813 (N_17813,N_12661,N_13809);
xor U17814 (N_17814,N_14680,N_14879);
nand U17815 (N_17815,N_15415,N_15474);
nand U17816 (N_17816,N_13090,N_14532);
and U17817 (N_17817,N_14896,N_15070);
and U17818 (N_17818,N_12537,N_14441);
nor U17819 (N_17819,N_13119,N_13450);
and U17820 (N_17820,N_12821,N_15567);
nor U17821 (N_17821,N_13817,N_12662);
and U17822 (N_17822,N_13359,N_12845);
nor U17823 (N_17823,N_13255,N_14543);
nor U17824 (N_17824,N_14631,N_14043);
nand U17825 (N_17825,N_14827,N_15033);
nand U17826 (N_17826,N_15518,N_14753);
and U17827 (N_17827,N_15430,N_13855);
and U17828 (N_17828,N_14803,N_15578);
xor U17829 (N_17829,N_15431,N_14060);
and U17830 (N_17830,N_13672,N_14006);
nand U17831 (N_17831,N_15456,N_13972);
or U17832 (N_17832,N_14886,N_15079);
xnor U17833 (N_17833,N_15267,N_12776);
nor U17834 (N_17834,N_13260,N_15174);
xnor U17835 (N_17835,N_12739,N_13004);
nand U17836 (N_17836,N_15047,N_13485);
nor U17837 (N_17837,N_14693,N_14432);
xor U17838 (N_17838,N_12911,N_12951);
or U17839 (N_17839,N_13952,N_13163);
nand U17840 (N_17840,N_14797,N_13126);
nand U17841 (N_17841,N_14044,N_13589);
nor U17842 (N_17842,N_13745,N_15316);
xor U17843 (N_17843,N_13005,N_15165);
nand U17844 (N_17844,N_12554,N_12904);
xnor U17845 (N_17845,N_13287,N_13447);
xor U17846 (N_17846,N_13501,N_14333);
xnor U17847 (N_17847,N_15484,N_13604);
or U17848 (N_17848,N_12873,N_13344);
or U17849 (N_17849,N_13061,N_13045);
xor U17850 (N_17850,N_12595,N_15486);
or U17851 (N_17851,N_13311,N_14484);
nand U17852 (N_17852,N_13584,N_12866);
or U17853 (N_17853,N_12783,N_13274);
and U17854 (N_17854,N_15466,N_14177);
xnor U17855 (N_17855,N_12788,N_14526);
nand U17856 (N_17856,N_15048,N_13856);
and U17857 (N_17857,N_15537,N_13049);
and U17858 (N_17858,N_12755,N_15190);
xor U17859 (N_17859,N_12536,N_15561);
nand U17860 (N_17860,N_12823,N_14234);
or U17861 (N_17861,N_13049,N_13786);
nor U17862 (N_17862,N_13680,N_14918);
or U17863 (N_17863,N_14463,N_15029);
nand U17864 (N_17864,N_13436,N_15528);
nand U17865 (N_17865,N_13941,N_12678);
and U17866 (N_17866,N_14805,N_14947);
or U17867 (N_17867,N_12644,N_15331);
or U17868 (N_17868,N_13302,N_15136);
and U17869 (N_17869,N_15506,N_14525);
and U17870 (N_17870,N_13248,N_12843);
nor U17871 (N_17871,N_13096,N_13565);
and U17872 (N_17872,N_13582,N_14832);
and U17873 (N_17873,N_15323,N_14004);
nand U17874 (N_17874,N_15264,N_14645);
or U17875 (N_17875,N_15573,N_12842);
and U17876 (N_17876,N_13778,N_12983);
nor U17877 (N_17877,N_15469,N_13993);
or U17878 (N_17878,N_12797,N_15136);
or U17879 (N_17879,N_15528,N_14937);
and U17880 (N_17880,N_15129,N_13052);
nor U17881 (N_17881,N_12846,N_13608);
nor U17882 (N_17882,N_14331,N_14537);
xor U17883 (N_17883,N_15462,N_13801);
or U17884 (N_17884,N_15418,N_13740);
nand U17885 (N_17885,N_13053,N_13770);
or U17886 (N_17886,N_15290,N_14186);
and U17887 (N_17887,N_14312,N_15577);
xnor U17888 (N_17888,N_12671,N_13036);
and U17889 (N_17889,N_15084,N_13152);
and U17890 (N_17890,N_13748,N_13901);
and U17891 (N_17891,N_13998,N_14402);
nor U17892 (N_17892,N_14297,N_13337);
nor U17893 (N_17893,N_13628,N_14693);
nand U17894 (N_17894,N_13941,N_15611);
nand U17895 (N_17895,N_15528,N_13990);
nand U17896 (N_17896,N_13875,N_14245);
xor U17897 (N_17897,N_12618,N_14150);
nand U17898 (N_17898,N_15452,N_13453);
or U17899 (N_17899,N_15580,N_13245);
and U17900 (N_17900,N_12765,N_13538);
nor U17901 (N_17901,N_12637,N_13524);
nand U17902 (N_17902,N_14086,N_15298);
xor U17903 (N_17903,N_13813,N_13816);
nor U17904 (N_17904,N_14077,N_13754);
or U17905 (N_17905,N_12840,N_13988);
nor U17906 (N_17906,N_15534,N_15085);
and U17907 (N_17907,N_13180,N_14719);
nand U17908 (N_17908,N_14813,N_13667);
xnor U17909 (N_17909,N_13615,N_13728);
xor U17910 (N_17910,N_12646,N_13909);
or U17911 (N_17911,N_14889,N_12652);
nand U17912 (N_17912,N_13482,N_14373);
nor U17913 (N_17913,N_14507,N_15030);
and U17914 (N_17914,N_14964,N_14428);
and U17915 (N_17915,N_14259,N_13507);
nor U17916 (N_17916,N_13707,N_13698);
and U17917 (N_17917,N_15529,N_14458);
or U17918 (N_17918,N_13709,N_12656);
or U17919 (N_17919,N_12916,N_15252);
nand U17920 (N_17920,N_14881,N_13580);
and U17921 (N_17921,N_13200,N_15320);
nand U17922 (N_17922,N_13699,N_13143);
xnor U17923 (N_17923,N_13634,N_13373);
and U17924 (N_17924,N_13350,N_14973);
xnor U17925 (N_17925,N_13532,N_12835);
xor U17926 (N_17926,N_14727,N_14635);
nor U17927 (N_17927,N_14080,N_13828);
and U17928 (N_17928,N_14700,N_12952);
xor U17929 (N_17929,N_13267,N_13338);
nor U17930 (N_17930,N_13742,N_13062);
nand U17931 (N_17931,N_15563,N_12521);
and U17932 (N_17932,N_15012,N_12820);
xnor U17933 (N_17933,N_15571,N_12724);
nand U17934 (N_17934,N_13579,N_15466);
nand U17935 (N_17935,N_12789,N_12648);
nor U17936 (N_17936,N_13854,N_13528);
nor U17937 (N_17937,N_15029,N_14609);
nand U17938 (N_17938,N_14491,N_12603);
or U17939 (N_17939,N_12779,N_13071);
nand U17940 (N_17940,N_13385,N_13073);
and U17941 (N_17941,N_15600,N_14724);
and U17942 (N_17942,N_15058,N_14549);
nor U17943 (N_17943,N_13442,N_14796);
nor U17944 (N_17944,N_12806,N_14992);
nor U17945 (N_17945,N_13595,N_13334);
and U17946 (N_17946,N_13529,N_15305);
and U17947 (N_17947,N_14192,N_14587);
and U17948 (N_17948,N_14543,N_12635);
xor U17949 (N_17949,N_13803,N_14409);
xor U17950 (N_17950,N_14164,N_12663);
nand U17951 (N_17951,N_12769,N_14567);
or U17952 (N_17952,N_13213,N_15049);
and U17953 (N_17953,N_13450,N_14868);
xnor U17954 (N_17954,N_15256,N_14168);
nor U17955 (N_17955,N_12701,N_14015);
nor U17956 (N_17956,N_12544,N_14249);
nand U17957 (N_17957,N_15234,N_13264);
xor U17958 (N_17958,N_13063,N_14822);
xnor U17959 (N_17959,N_13034,N_15373);
or U17960 (N_17960,N_13824,N_13956);
xor U17961 (N_17961,N_15196,N_14649);
or U17962 (N_17962,N_15037,N_15143);
and U17963 (N_17963,N_15039,N_15576);
xor U17964 (N_17964,N_14174,N_15224);
xnor U17965 (N_17965,N_12598,N_13894);
or U17966 (N_17966,N_13849,N_14979);
or U17967 (N_17967,N_12840,N_12738);
xor U17968 (N_17968,N_13709,N_13632);
or U17969 (N_17969,N_12548,N_13421);
xor U17970 (N_17970,N_12627,N_12976);
and U17971 (N_17971,N_13840,N_14897);
and U17972 (N_17972,N_15324,N_13697);
nand U17973 (N_17973,N_12857,N_14744);
and U17974 (N_17974,N_14870,N_13474);
and U17975 (N_17975,N_13183,N_12870);
xor U17976 (N_17976,N_15194,N_15147);
xor U17977 (N_17977,N_15269,N_13180);
or U17978 (N_17978,N_13310,N_15586);
xor U17979 (N_17979,N_13651,N_14392);
nand U17980 (N_17980,N_13770,N_14031);
xnor U17981 (N_17981,N_12849,N_15465);
xor U17982 (N_17982,N_13442,N_15043);
xor U17983 (N_17983,N_15458,N_14721);
nand U17984 (N_17984,N_14843,N_14528);
nor U17985 (N_17985,N_15230,N_15197);
nor U17986 (N_17986,N_14800,N_15546);
nor U17987 (N_17987,N_14627,N_13787);
and U17988 (N_17988,N_14282,N_13943);
or U17989 (N_17989,N_13369,N_14994);
and U17990 (N_17990,N_15131,N_12569);
nand U17991 (N_17991,N_12938,N_14183);
nor U17992 (N_17992,N_14721,N_14809);
and U17993 (N_17993,N_14349,N_14796);
and U17994 (N_17994,N_15205,N_14530);
nor U17995 (N_17995,N_15188,N_12850);
nor U17996 (N_17996,N_12709,N_13486);
nand U17997 (N_17997,N_13452,N_14535);
nor U17998 (N_17998,N_14506,N_13567);
and U17999 (N_17999,N_12981,N_15001);
and U18000 (N_18000,N_12969,N_15280);
and U18001 (N_18001,N_14220,N_15004);
xor U18002 (N_18002,N_14650,N_13905);
nor U18003 (N_18003,N_15547,N_13706);
xor U18004 (N_18004,N_12776,N_15458);
and U18005 (N_18005,N_14491,N_15233);
or U18006 (N_18006,N_13794,N_12654);
nand U18007 (N_18007,N_14014,N_12937);
nor U18008 (N_18008,N_12590,N_13947);
or U18009 (N_18009,N_15219,N_14374);
nand U18010 (N_18010,N_13651,N_15097);
nand U18011 (N_18011,N_14357,N_14396);
nand U18012 (N_18012,N_12878,N_15480);
and U18013 (N_18013,N_15292,N_13702);
or U18014 (N_18014,N_13477,N_12825);
xnor U18015 (N_18015,N_12633,N_14216);
nand U18016 (N_18016,N_12861,N_14604);
nand U18017 (N_18017,N_15261,N_15493);
xnor U18018 (N_18018,N_14438,N_13523);
xor U18019 (N_18019,N_12761,N_13421);
nor U18020 (N_18020,N_12704,N_15461);
nor U18021 (N_18021,N_14277,N_13895);
nand U18022 (N_18022,N_12558,N_13028);
nor U18023 (N_18023,N_14045,N_15517);
nor U18024 (N_18024,N_13443,N_15424);
and U18025 (N_18025,N_13849,N_15157);
nand U18026 (N_18026,N_15336,N_14164);
or U18027 (N_18027,N_13500,N_12917);
nand U18028 (N_18028,N_15613,N_15168);
xor U18029 (N_18029,N_15406,N_13597);
nand U18030 (N_18030,N_15587,N_14994);
and U18031 (N_18031,N_13694,N_15034);
nand U18032 (N_18032,N_14525,N_12921);
or U18033 (N_18033,N_14936,N_15010);
nand U18034 (N_18034,N_12858,N_14973);
or U18035 (N_18035,N_15543,N_13519);
xor U18036 (N_18036,N_12668,N_14057);
xor U18037 (N_18037,N_15393,N_13239);
and U18038 (N_18038,N_13498,N_12631);
nand U18039 (N_18039,N_15270,N_15485);
and U18040 (N_18040,N_13907,N_12963);
nor U18041 (N_18041,N_14057,N_15396);
xor U18042 (N_18042,N_15294,N_13128);
and U18043 (N_18043,N_14919,N_13854);
nor U18044 (N_18044,N_14973,N_14894);
and U18045 (N_18045,N_13530,N_12694);
or U18046 (N_18046,N_13581,N_15053);
nor U18047 (N_18047,N_15453,N_12869);
nor U18048 (N_18048,N_13855,N_15363);
xnor U18049 (N_18049,N_13102,N_14994);
and U18050 (N_18050,N_13622,N_14998);
xor U18051 (N_18051,N_12930,N_14516);
nor U18052 (N_18052,N_14236,N_15423);
and U18053 (N_18053,N_13127,N_15249);
nor U18054 (N_18054,N_13753,N_14140);
nor U18055 (N_18055,N_14187,N_14154);
nand U18056 (N_18056,N_12617,N_13446);
nor U18057 (N_18057,N_13970,N_12634);
or U18058 (N_18058,N_13797,N_15425);
or U18059 (N_18059,N_14107,N_14178);
nand U18060 (N_18060,N_13164,N_13076);
or U18061 (N_18061,N_13801,N_12561);
xor U18062 (N_18062,N_14112,N_13520);
and U18063 (N_18063,N_14468,N_15071);
xor U18064 (N_18064,N_12751,N_15025);
nor U18065 (N_18065,N_12535,N_12863);
and U18066 (N_18066,N_15489,N_12606);
nor U18067 (N_18067,N_14877,N_13839);
and U18068 (N_18068,N_12819,N_15209);
xnor U18069 (N_18069,N_12928,N_13062);
or U18070 (N_18070,N_13855,N_15138);
nand U18071 (N_18071,N_12847,N_14811);
nor U18072 (N_18072,N_12505,N_12603);
xnor U18073 (N_18073,N_14768,N_12775);
nand U18074 (N_18074,N_14873,N_13480);
nor U18075 (N_18075,N_12536,N_12790);
nand U18076 (N_18076,N_12853,N_14074);
xnor U18077 (N_18077,N_13406,N_14645);
or U18078 (N_18078,N_15281,N_14112);
and U18079 (N_18079,N_13506,N_14017);
or U18080 (N_18080,N_13093,N_14207);
xnor U18081 (N_18081,N_14683,N_14051);
nand U18082 (N_18082,N_14796,N_12833);
and U18083 (N_18083,N_14698,N_15185);
and U18084 (N_18084,N_14700,N_13074);
or U18085 (N_18085,N_13899,N_13245);
nand U18086 (N_18086,N_13741,N_15450);
and U18087 (N_18087,N_14145,N_14919);
nor U18088 (N_18088,N_14171,N_15280);
and U18089 (N_18089,N_14382,N_14313);
or U18090 (N_18090,N_13699,N_15544);
and U18091 (N_18091,N_15450,N_13720);
or U18092 (N_18092,N_14424,N_14925);
nor U18093 (N_18093,N_14536,N_13889);
and U18094 (N_18094,N_14107,N_14852);
or U18095 (N_18095,N_15443,N_12567);
nor U18096 (N_18096,N_14322,N_14790);
nand U18097 (N_18097,N_14144,N_12769);
or U18098 (N_18098,N_13884,N_13020);
nand U18099 (N_18099,N_12933,N_14008);
nor U18100 (N_18100,N_14381,N_14964);
nand U18101 (N_18101,N_15122,N_13647);
or U18102 (N_18102,N_13569,N_14577);
nand U18103 (N_18103,N_13671,N_13319);
xor U18104 (N_18104,N_14535,N_14913);
nand U18105 (N_18105,N_14131,N_14861);
nor U18106 (N_18106,N_13126,N_13990);
xor U18107 (N_18107,N_15391,N_13593);
and U18108 (N_18108,N_15199,N_13660);
and U18109 (N_18109,N_12589,N_12961);
and U18110 (N_18110,N_14041,N_12998);
and U18111 (N_18111,N_15229,N_12955);
and U18112 (N_18112,N_13672,N_15000);
and U18113 (N_18113,N_14142,N_15411);
nor U18114 (N_18114,N_14906,N_12572);
or U18115 (N_18115,N_13388,N_14687);
nor U18116 (N_18116,N_14861,N_12744);
and U18117 (N_18117,N_12559,N_12726);
or U18118 (N_18118,N_12711,N_15040);
xnor U18119 (N_18119,N_13355,N_15206);
and U18120 (N_18120,N_15306,N_14211);
nor U18121 (N_18121,N_13956,N_15526);
nor U18122 (N_18122,N_12736,N_14020);
or U18123 (N_18123,N_15395,N_14788);
nand U18124 (N_18124,N_14797,N_14880);
nor U18125 (N_18125,N_14347,N_12869);
xor U18126 (N_18126,N_15147,N_14347);
and U18127 (N_18127,N_14730,N_13955);
nor U18128 (N_18128,N_13706,N_14225);
xor U18129 (N_18129,N_13635,N_13377);
nand U18130 (N_18130,N_15037,N_12920);
or U18131 (N_18131,N_14862,N_15324);
and U18132 (N_18132,N_13904,N_13027);
or U18133 (N_18133,N_13976,N_14978);
nor U18134 (N_18134,N_14209,N_15429);
nor U18135 (N_18135,N_13665,N_13543);
nor U18136 (N_18136,N_14415,N_13036);
or U18137 (N_18137,N_15028,N_14019);
xor U18138 (N_18138,N_15205,N_14166);
nor U18139 (N_18139,N_12943,N_13048);
and U18140 (N_18140,N_13789,N_13097);
xnor U18141 (N_18141,N_13988,N_13588);
xor U18142 (N_18142,N_14773,N_14659);
nand U18143 (N_18143,N_14985,N_12868);
xnor U18144 (N_18144,N_12578,N_13755);
nor U18145 (N_18145,N_14799,N_12686);
or U18146 (N_18146,N_14133,N_15384);
nor U18147 (N_18147,N_12784,N_14166);
nor U18148 (N_18148,N_13134,N_15541);
nor U18149 (N_18149,N_15065,N_13919);
or U18150 (N_18150,N_13612,N_12675);
nor U18151 (N_18151,N_12608,N_14548);
or U18152 (N_18152,N_15143,N_13536);
and U18153 (N_18153,N_15574,N_13574);
nand U18154 (N_18154,N_13866,N_15326);
nor U18155 (N_18155,N_14283,N_12767);
xor U18156 (N_18156,N_14161,N_15562);
nand U18157 (N_18157,N_13956,N_12927);
nor U18158 (N_18158,N_14024,N_13776);
and U18159 (N_18159,N_13052,N_15511);
and U18160 (N_18160,N_12698,N_13954);
nor U18161 (N_18161,N_14224,N_13319);
nand U18162 (N_18162,N_14138,N_14139);
nor U18163 (N_18163,N_13116,N_13132);
nor U18164 (N_18164,N_14112,N_14384);
xnor U18165 (N_18165,N_14904,N_14172);
and U18166 (N_18166,N_13672,N_15524);
nor U18167 (N_18167,N_14066,N_14456);
nor U18168 (N_18168,N_14614,N_13766);
nand U18169 (N_18169,N_15431,N_14722);
nand U18170 (N_18170,N_15464,N_15003);
or U18171 (N_18171,N_13456,N_13009);
nand U18172 (N_18172,N_14504,N_12709);
nand U18173 (N_18173,N_13489,N_14206);
xnor U18174 (N_18174,N_15231,N_13107);
nor U18175 (N_18175,N_15615,N_13809);
nand U18176 (N_18176,N_13781,N_12974);
xor U18177 (N_18177,N_13360,N_15038);
nand U18178 (N_18178,N_12922,N_14260);
nand U18179 (N_18179,N_13442,N_14988);
nand U18180 (N_18180,N_14000,N_12806);
or U18181 (N_18181,N_15245,N_14263);
and U18182 (N_18182,N_15230,N_14797);
and U18183 (N_18183,N_13905,N_14408);
nand U18184 (N_18184,N_14775,N_12803);
nor U18185 (N_18185,N_13961,N_14750);
nand U18186 (N_18186,N_13704,N_14720);
xnor U18187 (N_18187,N_15618,N_15380);
nor U18188 (N_18188,N_13465,N_13519);
and U18189 (N_18189,N_15392,N_13616);
nor U18190 (N_18190,N_13520,N_15022);
nand U18191 (N_18191,N_12885,N_15505);
nor U18192 (N_18192,N_14103,N_13117);
nand U18193 (N_18193,N_12789,N_13296);
and U18194 (N_18194,N_15624,N_14333);
and U18195 (N_18195,N_13655,N_13066);
xnor U18196 (N_18196,N_15055,N_14436);
xnor U18197 (N_18197,N_14592,N_14135);
and U18198 (N_18198,N_14838,N_15202);
or U18199 (N_18199,N_12899,N_14493);
nor U18200 (N_18200,N_13356,N_13283);
or U18201 (N_18201,N_12655,N_12602);
nand U18202 (N_18202,N_14080,N_14244);
nor U18203 (N_18203,N_12766,N_14487);
nor U18204 (N_18204,N_12818,N_14778);
nor U18205 (N_18205,N_13274,N_14158);
xor U18206 (N_18206,N_14261,N_12777);
nand U18207 (N_18207,N_13013,N_15246);
and U18208 (N_18208,N_15319,N_15594);
xnor U18209 (N_18209,N_12596,N_13813);
and U18210 (N_18210,N_13100,N_13922);
xnor U18211 (N_18211,N_13531,N_12829);
or U18212 (N_18212,N_15220,N_13927);
xor U18213 (N_18213,N_13231,N_12615);
nand U18214 (N_18214,N_15612,N_14658);
nand U18215 (N_18215,N_15571,N_15413);
nor U18216 (N_18216,N_15298,N_14442);
xnor U18217 (N_18217,N_15293,N_13891);
xor U18218 (N_18218,N_14089,N_14409);
and U18219 (N_18219,N_12951,N_13851);
and U18220 (N_18220,N_14712,N_14682);
and U18221 (N_18221,N_12539,N_12511);
nor U18222 (N_18222,N_13227,N_13355);
and U18223 (N_18223,N_14205,N_15465);
nor U18224 (N_18224,N_14372,N_12613);
and U18225 (N_18225,N_14235,N_12910);
nand U18226 (N_18226,N_14067,N_14751);
or U18227 (N_18227,N_13025,N_14496);
xnor U18228 (N_18228,N_13552,N_14859);
and U18229 (N_18229,N_14291,N_13839);
or U18230 (N_18230,N_12958,N_14986);
nor U18231 (N_18231,N_12665,N_14474);
or U18232 (N_18232,N_13529,N_13036);
xnor U18233 (N_18233,N_14363,N_14969);
nand U18234 (N_18234,N_15372,N_15120);
xor U18235 (N_18235,N_13773,N_14924);
nor U18236 (N_18236,N_14927,N_14237);
and U18237 (N_18237,N_13230,N_12622);
xnor U18238 (N_18238,N_14297,N_14416);
or U18239 (N_18239,N_12651,N_13682);
nor U18240 (N_18240,N_15287,N_14486);
nand U18241 (N_18241,N_12707,N_15321);
xnor U18242 (N_18242,N_13502,N_14380);
or U18243 (N_18243,N_14810,N_12650);
and U18244 (N_18244,N_13416,N_13466);
or U18245 (N_18245,N_12769,N_13689);
or U18246 (N_18246,N_14379,N_14860);
or U18247 (N_18247,N_12814,N_14744);
nor U18248 (N_18248,N_12958,N_12785);
nor U18249 (N_18249,N_12512,N_15180);
and U18250 (N_18250,N_12616,N_13909);
nor U18251 (N_18251,N_15004,N_15290);
or U18252 (N_18252,N_14266,N_15198);
and U18253 (N_18253,N_15251,N_12891);
or U18254 (N_18254,N_13481,N_14911);
and U18255 (N_18255,N_14378,N_15483);
nor U18256 (N_18256,N_14737,N_14046);
xor U18257 (N_18257,N_14823,N_13784);
nand U18258 (N_18258,N_13633,N_14753);
nor U18259 (N_18259,N_13226,N_13980);
or U18260 (N_18260,N_14673,N_14152);
nor U18261 (N_18261,N_15441,N_13021);
xor U18262 (N_18262,N_15591,N_13988);
or U18263 (N_18263,N_12626,N_14496);
nor U18264 (N_18264,N_13701,N_14735);
and U18265 (N_18265,N_15086,N_13431);
xor U18266 (N_18266,N_13722,N_12672);
nor U18267 (N_18267,N_14952,N_14060);
and U18268 (N_18268,N_13708,N_13050);
and U18269 (N_18269,N_13495,N_14209);
or U18270 (N_18270,N_14898,N_13514);
or U18271 (N_18271,N_14633,N_12992);
and U18272 (N_18272,N_13138,N_15173);
nand U18273 (N_18273,N_15121,N_13774);
nand U18274 (N_18274,N_13338,N_14214);
nand U18275 (N_18275,N_13169,N_13542);
or U18276 (N_18276,N_15028,N_14864);
or U18277 (N_18277,N_14790,N_13870);
nor U18278 (N_18278,N_14438,N_15130);
nand U18279 (N_18279,N_14066,N_13957);
xor U18280 (N_18280,N_13481,N_14405);
nor U18281 (N_18281,N_14894,N_12643);
or U18282 (N_18282,N_12674,N_13477);
nor U18283 (N_18283,N_13603,N_12919);
nand U18284 (N_18284,N_14163,N_13393);
nand U18285 (N_18285,N_14931,N_13599);
nor U18286 (N_18286,N_13603,N_14586);
xnor U18287 (N_18287,N_13687,N_15262);
and U18288 (N_18288,N_14408,N_15304);
and U18289 (N_18289,N_14954,N_14264);
and U18290 (N_18290,N_13356,N_14040);
and U18291 (N_18291,N_13564,N_12830);
and U18292 (N_18292,N_13072,N_13062);
and U18293 (N_18293,N_13556,N_15257);
xor U18294 (N_18294,N_13918,N_15378);
nor U18295 (N_18295,N_13527,N_12731);
or U18296 (N_18296,N_15153,N_12808);
xor U18297 (N_18297,N_15528,N_14734);
nand U18298 (N_18298,N_13090,N_14510);
nor U18299 (N_18299,N_13611,N_13081);
xnor U18300 (N_18300,N_13121,N_13510);
nor U18301 (N_18301,N_13665,N_15186);
and U18302 (N_18302,N_15436,N_15221);
nand U18303 (N_18303,N_13051,N_13354);
or U18304 (N_18304,N_13946,N_14164);
nor U18305 (N_18305,N_13517,N_14420);
nor U18306 (N_18306,N_12854,N_14432);
xor U18307 (N_18307,N_15156,N_12738);
nor U18308 (N_18308,N_12686,N_12748);
and U18309 (N_18309,N_12689,N_15342);
or U18310 (N_18310,N_15593,N_14337);
and U18311 (N_18311,N_13015,N_13097);
nand U18312 (N_18312,N_14299,N_14059);
or U18313 (N_18313,N_14388,N_14911);
nor U18314 (N_18314,N_12917,N_15113);
nor U18315 (N_18315,N_14130,N_13397);
or U18316 (N_18316,N_15251,N_13586);
or U18317 (N_18317,N_15252,N_15255);
or U18318 (N_18318,N_14263,N_12662);
nor U18319 (N_18319,N_13987,N_14315);
or U18320 (N_18320,N_12620,N_13897);
nand U18321 (N_18321,N_15211,N_13248);
nand U18322 (N_18322,N_15409,N_15014);
and U18323 (N_18323,N_15527,N_14729);
or U18324 (N_18324,N_15510,N_13232);
and U18325 (N_18325,N_14752,N_14502);
or U18326 (N_18326,N_13604,N_14007);
nand U18327 (N_18327,N_15503,N_13289);
nor U18328 (N_18328,N_14904,N_13019);
xnor U18329 (N_18329,N_14427,N_15464);
or U18330 (N_18330,N_14695,N_13278);
nor U18331 (N_18331,N_13336,N_12560);
or U18332 (N_18332,N_13497,N_15472);
or U18333 (N_18333,N_15247,N_14325);
and U18334 (N_18334,N_15078,N_14577);
nand U18335 (N_18335,N_13340,N_15545);
and U18336 (N_18336,N_13692,N_14704);
nand U18337 (N_18337,N_13088,N_12962);
xnor U18338 (N_18338,N_12507,N_15574);
and U18339 (N_18339,N_15253,N_12840);
or U18340 (N_18340,N_14830,N_13748);
xnor U18341 (N_18341,N_14687,N_12709);
xor U18342 (N_18342,N_13094,N_13411);
nand U18343 (N_18343,N_12537,N_13704);
and U18344 (N_18344,N_15096,N_14400);
xnor U18345 (N_18345,N_13761,N_15304);
xor U18346 (N_18346,N_14850,N_15585);
xor U18347 (N_18347,N_14430,N_14049);
nor U18348 (N_18348,N_12832,N_12613);
xor U18349 (N_18349,N_13082,N_13486);
nand U18350 (N_18350,N_13326,N_14379);
xor U18351 (N_18351,N_15051,N_14022);
or U18352 (N_18352,N_13187,N_14010);
or U18353 (N_18353,N_13844,N_15045);
nand U18354 (N_18354,N_12762,N_13766);
or U18355 (N_18355,N_15290,N_14778);
and U18356 (N_18356,N_15603,N_13655);
or U18357 (N_18357,N_12905,N_14756);
or U18358 (N_18358,N_13084,N_15485);
or U18359 (N_18359,N_13727,N_14123);
or U18360 (N_18360,N_15136,N_14446);
nor U18361 (N_18361,N_13089,N_12546);
xnor U18362 (N_18362,N_13250,N_13147);
and U18363 (N_18363,N_14293,N_14528);
nor U18364 (N_18364,N_14807,N_15021);
and U18365 (N_18365,N_13559,N_14895);
and U18366 (N_18366,N_12920,N_14228);
xor U18367 (N_18367,N_14972,N_13443);
or U18368 (N_18368,N_13211,N_14696);
nand U18369 (N_18369,N_13380,N_14828);
and U18370 (N_18370,N_14624,N_14219);
or U18371 (N_18371,N_14945,N_15018);
and U18372 (N_18372,N_14711,N_15585);
nor U18373 (N_18373,N_13923,N_14791);
nand U18374 (N_18374,N_12729,N_12684);
and U18375 (N_18375,N_13683,N_14466);
and U18376 (N_18376,N_12993,N_14024);
or U18377 (N_18377,N_13848,N_14620);
xnor U18378 (N_18378,N_13355,N_14077);
xor U18379 (N_18379,N_13444,N_12562);
or U18380 (N_18380,N_13016,N_14627);
or U18381 (N_18381,N_14780,N_13265);
nor U18382 (N_18382,N_12791,N_12814);
and U18383 (N_18383,N_14752,N_12763);
and U18384 (N_18384,N_12692,N_13601);
xor U18385 (N_18385,N_12899,N_14436);
and U18386 (N_18386,N_15018,N_14466);
nor U18387 (N_18387,N_12752,N_13841);
and U18388 (N_18388,N_14562,N_13881);
nor U18389 (N_18389,N_13562,N_14527);
xor U18390 (N_18390,N_13726,N_14592);
nor U18391 (N_18391,N_15378,N_15413);
xnor U18392 (N_18392,N_14260,N_13968);
or U18393 (N_18393,N_13974,N_15081);
nand U18394 (N_18394,N_13203,N_14246);
nor U18395 (N_18395,N_15311,N_13460);
nor U18396 (N_18396,N_14863,N_12995);
xor U18397 (N_18397,N_14599,N_13825);
or U18398 (N_18398,N_13102,N_13156);
xor U18399 (N_18399,N_12966,N_13508);
and U18400 (N_18400,N_12538,N_13571);
xnor U18401 (N_18401,N_13254,N_12928);
nor U18402 (N_18402,N_15418,N_14159);
xnor U18403 (N_18403,N_12997,N_13831);
xor U18404 (N_18404,N_14751,N_14038);
nor U18405 (N_18405,N_13899,N_12730);
and U18406 (N_18406,N_15472,N_14515);
nand U18407 (N_18407,N_15422,N_14382);
nor U18408 (N_18408,N_15435,N_14574);
nand U18409 (N_18409,N_15119,N_13915);
xor U18410 (N_18410,N_14786,N_14645);
nand U18411 (N_18411,N_15149,N_14339);
xnor U18412 (N_18412,N_14484,N_14359);
xor U18413 (N_18413,N_15460,N_13439);
xor U18414 (N_18414,N_12661,N_13882);
nand U18415 (N_18415,N_13298,N_13135);
and U18416 (N_18416,N_12961,N_14240);
nand U18417 (N_18417,N_13967,N_14507);
nand U18418 (N_18418,N_12814,N_14463);
nor U18419 (N_18419,N_15259,N_14390);
nor U18420 (N_18420,N_14647,N_12615);
nand U18421 (N_18421,N_14499,N_14629);
xnor U18422 (N_18422,N_13511,N_14934);
and U18423 (N_18423,N_13017,N_13248);
or U18424 (N_18424,N_14959,N_13260);
or U18425 (N_18425,N_14027,N_13328);
nor U18426 (N_18426,N_14263,N_12998);
and U18427 (N_18427,N_13443,N_13544);
xor U18428 (N_18428,N_12691,N_15251);
xor U18429 (N_18429,N_14557,N_15309);
xnor U18430 (N_18430,N_13843,N_15169);
or U18431 (N_18431,N_15158,N_14591);
nand U18432 (N_18432,N_15395,N_12789);
nand U18433 (N_18433,N_13114,N_12736);
or U18434 (N_18434,N_13494,N_13203);
nand U18435 (N_18435,N_13522,N_14752);
and U18436 (N_18436,N_14233,N_14553);
or U18437 (N_18437,N_13303,N_12961);
nand U18438 (N_18438,N_14820,N_15071);
xor U18439 (N_18439,N_15550,N_14241);
nor U18440 (N_18440,N_14519,N_14717);
nor U18441 (N_18441,N_15370,N_14750);
nor U18442 (N_18442,N_15062,N_13420);
nor U18443 (N_18443,N_13992,N_12731);
and U18444 (N_18444,N_14417,N_12748);
nor U18445 (N_18445,N_15482,N_13412);
and U18446 (N_18446,N_12541,N_13957);
or U18447 (N_18447,N_15073,N_14630);
and U18448 (N_18448,N_12948,N_12810);
or U18449 (N_18449,N_12517,N_15081);
and U18450 (N_18450,N_14967,N_14905);
nand U18451 (N_18451,N_12507,N_12886);
nand U18452 (N_18452,N_13087,N_14299);
and U18453 (N_18453,N_14301,N_14272);
nor U18454 (N_18454,N_14709,N_14973);
nand U18455 (N_18455,N_12650,N_13609);
or U18456 (N_18456,N_13654,N_13800);
nand U18457 (N_18457,N_14812,N_15419);
nor U18458 (N_18458,N_14748,N_12725);
xnor U18459 (N_18459,N_14854,N_15345);
or U18460 (N_18460,N_12604,N_14915);
and U18461 (N_18461,N_12563,N_14449);
or U18462 (N_18462,N_14460,N_13434);
or U18463 (N_18463,N_13795,N_13032);
nor U18464 (N_18464,N_15026,N_14949);
nand U18465 (N_18465,N_12813,N_13031);
nor U18466 (N_18466,N_14118,N_12517);
or U18467 (N_18467,N_14044,N_14113);
or U18468 (N_18468,N_15240,N_13231);
nand U18469 (N_18469,N_14062,N_14942);
xnor U18470 (N_18470,N_14176,N_15083);
nor U18471 (N_18471,N_14817,N_15248);
xor U18472 (N_18472,N_14666,N_15157);
nor U18473 (N_18473,N_14557,N_14896);
and U18474 (N_18474,N_14407,N_13162);
nand U18475 (N_18475,N_15439,N_15213);
nand U18476 (N_18476,N_13614,N_13030);
nand U18477 (N_18477,N_15205,N_15462);
xnor U18478 (N_18478,N_13086,N_15459);
or U18479 (N_18479,N_13867,N_15504);
and U18480 (N_18480,N_14392,N_14568);
xor U18481 (N_18481,N_12940,N_13035);
nand U18482 (N_18482,N_12601,N_13042);
nand U18483 (N_18483,N_13683,N_14334);
xor U18484 (N_18484,N_14686,N_13132);
and U18485 (N_18485,N_15346,N_14996);
xor U18486 (N_18486,N_15214,N_15607);
nand U18487 (N_18487,N_15237,N_13176);
xor U18488 (N_18488,N_15013,N_13726);
xor U18489 (N_18489,N_12605,N_15492);
xor U18490 (N_18490,N_14801,N_13604);
nor U18491 (N_18491,N_15503,N_15433);
nor U18492 (N_18492,N_14974,N_15428);
and U18493 (N_18493,N_15080,N_15338);
nand U18494 (N_18494,N_15309,N_14132);
or U18495 (N_18495,N_14124,N_14992);
xnor U18496 (N_18496,N_14677,N_13966);
nor U18497 (N_18497,N_15154,N_15586);
nand U18498 (N_18498,N_12644,N_14708);
or U18499 (N_18499,N_12616,N_13158);
and U18500 (N_18500,N_13505,N_13184);
nor U18501 (N_18501,N_15221,N_14983);
xor U18502 (N_18502,N_14437,N_13462);
and U18503 (N_18503,N_14602,N_14363);
or U18504 (N_18504,N_14835,N_13827);
and U18505 (N_18505,N_12800,N_13001);
and U18506 (N_18506,N_14109,N_13633);
and U18507 (N_18507,N_14437,N_15429);
xor U18508 (N_18508,N_13842,N_12730);
and U18509 (N_18509,N_13406,N_14764);
and U18510 (N_18510,N_14528,N_14933);
nand U18511 (N_18511,N_12965,N_14460);
and U18512 (N_18512,N_12852,N_14291);
or U18513 (N_18513,N_14120,N_13641);
nand U18514 (N_18514,N_14407,N_13209);
and U18515 (N_18515,N_14250,N_14950);
and U18516 (N_18516,N_13992,N_14743);
or U18517 (N_18517,N_12514,N_12706);
xor U18518 (N_18518,N_15557,N_13152);
xnor U18519 (N_18519,N_12544,N_14771);
nor U18520 (N_18520,N_15517,N_14739);
and U18521 (N_18521,N_13201,N_15581);
and U18522 (N_18522,N_13652,N_14246);
nand U18523 (N_18523,N_13628,N_12653);
nor U18524 (N_18524,N_14383,N_13073);
or U18525 (N_18525,N_12689,N_13826);
or U18526 (N_18526,N_12572,N_15488);
and U18527 (N_18527,N_14506,N_13426);
and U18528 (N_18528,N_12918,N_14981);
nand U18529 (N_18529,N_14817,N_14604);
or U18530 (N_18530,N_14963,N_15467);
or U18531 (N_18531,N_15542,N_13320);
xor U18532 (N_18532,N_13792,N_15327);
and U18533 (N_18533,N_14476,N_14673);
and U18534 (N_18534,N_14985,N_14472);
or U18535 (N_18535,N_14914,N_13324);
nand U18536 (N_18536,N_14233,N_13868);
and U18537 (N_18537,N_12682,N_15135);
xor U18538 (N_18538,N_12630,N_12652);
xnor U18539 (N_18539,N_14269,N_13691);
nor U18540 (N_18540,N_12756,N_12909);
xor U18541 (N_18541,N_14130,N_12888);
nor U18542 (N_18542,N_13625,N_14012);
and U18543 (N_18543,N_12714,N_13132);
xor U18544 (N_18544,N_13354,N_14075);
and U18545 (N_18545,N_14394,N_13927);
nand U18546 (N_18546,N_13200,N_14379);
or U18547 (N_18547,N_13761,N_12934);
xnor U18548 (N_18548,N_13693,N_13463);
xnor U18549 (N_18549,N_12929,N_13510);
xnor U18550 (N_18550,N_14797,N_14237);
and U18551 (N_18551,N_14970,N_12869);
nand U18552 (N_18552,N_14595,N_13546);
nand U18553 (N_18553,N_14738,N_12621);
nor U18554 (N_18554,N_14358,N_13355);
or U18555 (N_18555,N_13496,N_13997);
nand U18556 (N_18556,N_15075,N_15394);
or U18557 (N_18557,N_14872,N_14296);
xnor U18558 (N_18558,N_13317,N_14291);
xor U18559 (N_18559,N_13313,N_14615);
nand U18560 (N_18560,N_14568,N_13695);
nor U18561 (N_18561,N_14724,N_14483);
xnor U18562 (N_18562,N_14964,N_12914);
or U18563 (N_18563,N_13620,N_14218);
or U18564 (N_18564,N_12981,N_12641);
nor U18565 (N_18565,N_12881,N_14695);
nor U18566 (N_18566,N_13562,N_14716);
nand U18567 (N_18567,N_12852,N_14565);
nand U18568 (N_18568,N_15298,N_12605);
or U18569 (N_18569,N_14922,N_14630);
nand U18570 (N_18570,N_15585,N_14422);
nand U18571 (N_18571,N_15077,N_13915);
or U18572 (N_18572,N_13953,N_15616);
or U18573 (N_18573,N_15200,N_12503);
nor U18574 (N_18574,N_15346,N_13277);
xor U18575 (N_18575,N_13118,N_15308);
nand U18576 (N_18576,N_15057,N_13177);
nand U18577 (N_18577,N_15031,N_14279);
nor U18578 (N_18578,N_15288,N_13898);
and U18579 (N_18579,N_14776,N_15100);
nor U18580 (N_18580,N_13936,N_13609);
nand U18581 (N_18581,N_14728,N_15057);
nor U18582 (N_18582,N_14199,N_12600);
and U18583 (N_18583,N_12859,N_15438);
and U18584 (N_18584,N_12549,N_12557);
nor U18585 (N_18585,N_12556,N_14884);
nand U18586 (N_18586,N_13213,N_14587);
nand U18587 (N_18587,N_14609,N_14243);
and U18588 (N_18588,N_15017,N_15034);
and U18589 (N_18589,N_12677,N_14137);
nand U18590 (N_18590,N_15021,N_13369);
xnor U18591 (N_18591,N_12920,N_13926);
xnor U18592 (N_18592,N_13658,N_12782);
xnor U18593 (N_18593,N_14031,N_15295);
or U18594 (N_18594,N_13891,N_15430);
nand U18595 (N_18595,N_15211,N_13926);
nor U18596 (N_18596,N_13949,N_13216);
nor U18597 (N_18597,N_13209,N_12885);
and U18598 (N_18598,N_14706,N_13552);
nor U18599 (N_18599,N_15543,N_15587);
or U18600 (N_18600,N_15164,N_12953);
nor U18601 (N_18601,N_12775,N_13338);
nand U18602 (N_18602,N_13203,N_13833);
nand U18603 (N_18603,N_13408,N_14553);
and U18604 (N_18604,N_14895,N_14044);
nand U18605 (N_18605,N_14042,N_12543);
nor U18606 (N_18606,N_13910,N_13162);
nor U18607 (N_18607,N_14489,N_15411);
nand U18608 (N_18608,N_13634,N_15074);
nand U18609 (N_18609,N_12933,N_15531);
and U18610 (N_18610,N_14662,N_13624);
nand U18611 (N_18611,N_14081,N_13673);
nand U18612 (N_18612,N_15605,N_13969);
nand U18613 (N_18613,N_13704,N_14917);
and U18614 (N_18614,N_15301,N_13685);
or U18615 (N_18615,N_13731,N_13285);
xor U18616 (N_18616,N_14043,N_13023);
xnor U18617 (N_18617,N_12685,N_14720);
xnor U18618 (N_18618,N_13848,N_14931);
nor U18619 (N_18619,N_15131,N_14417);
nand U18620 (N_18620,N_15173,N_13673);
or U18621 (N_18621,N_13658,N_15504);
or U18622 (N_18622,N_15117,N_13645);
nor U18623 (N_18623,N_13517,N_13978);
xnor U18624 (N_18624,N_13345,N_13923);
or U18625 (N_18625,N_13448,N_14787);
and U18626 (N_18626,N_13822,N_13721);
nor U18627 (N_18627,N_14005,N_15319);
nor U18628 (N_18628,N_14837,N_12977);
or U18629 (N_18629,N_12508,N_15589);
xor U18630 (N_18630,N_13550,N_13958);
xor U18631 (N_18631,N_13596,N_14441);
nor U18632 (N_18632,N_15004,N_14288);
and U18633 (N_18633,N_15582,N_14133);
nand U18634 (N_18634,N_15372,N_14501);
xor U18635 (N_18635,N_13312,N_15309);
and U18636 (N_18636,N_13693,N_14572);
nand U18637 (N_18637,N_14354,N_14553);
nand U18638 (N_18638,N_14924,N_13822);
xnor U18639 (N_18639,N_12936,N_14179);
nor U18640 (N_18640,N_12708,N_13261);
and U18641 (N_18641,N_12695,N_15002);
nor U18642 (N_18642,N_13289,N_13220);
xor U18643 (N_18643,N_15198,N_15408);
or U18644 (N_18644,N_13190,N_13710);
xnor U18645 (N_18645,N_13522,N_13245);
and U18646 (N_18646,N_14138,N_12978);
nand U18647 (N_18647,N_13626,N_14089);
or U18648 (N_18648,N_14481,N_13165);
and U18649 (N_18649,N_12588,N_15318);
nor U18650 (N_18650,N_13477,N_12527);
xnor U18651 (N_18651,N_14417,N_14215);
or U18652 (N_18652,N_14900,N_14366);
xor U18653 (N_18653,N_13308,N_14784);
nor U18654 (N_18654,N_13293,N_14215);
nor U18655 (N_18655,N_14136,N_14156);
xor U18656 (N_18656,N_12751,N_13153);
and U18657 (N_18657,N_12802,N_14807);
nor U18658 (N_18658,N_13805,N_14998);
or U18659 (N_18659,N_12542,N_14645);
nand U18660 (N_18660,N_14357,N_14496);
or U18661 (N_18661,N_12898,N_13000);
nand U18662 (N_18662,N_15313,N_13492);
nor U18663 (N_18663,N_14672,N_12744);
or U18664 (N_18664,N_14770,N_14461);
xor U18665 (N_18665,N_14759,N_14948);
and U18666 (N_18666,N_12646,N_14000);
and U18667 (N_18667,N_15000,N_13539);
and U18668 (N_18668,N_14676,N_14362);
nand U18669 (N_18669,N_13927,N_14968);
xor U18670 (N_18670,N_12988,N_14469);
and U18671 (N_18671,N_13073,N_13965);
and U18672 (N_18672,N_12576,N_14411);
xor U18673 (N_18673,N_13825,N_14457);
nand U18674 (N_18674,N_13958,N_15075);
or U18675 (N_18675,N_15247,N_13027);
and U18676 (N_18676,N_15376,N_14188);
or U18677 (N_18677,N_15225,N_15009);
nand U18678 (N_18678,N_14289,N_15053);
or U18679 (N_18679,N_13900,N_12620);
or U18680 (N_18680,N_12943,N_13617);
xnor U18681 (N_18681,N_14837,N_15129);
nor U18682 (N_18682,N_15139,N_13937);
nand U18683 (N_18683,N_13091,N_14292);
nand U18684 (N_18684,N_12698,N_13667);
nand U18685 (N_18685,N_14496,N_13378);
nor U18686 (N_18686,N_13555,N_15467);
nand U18687 (N_18687,N_13780,N_15422);
nor U18688 (N_18688,N_13189,N_12732);
and U18689 (N_18689,N_13832,N_15231);
xor U18690 (N_18690,N_14070,N_14812);
nor U18691 (N_18691,N_12534,N_14351);
nand U18692 (N_18692,N_13410,N_14657);
nor U18693 (N_18693,N_14510,N_14010);
and U18694 (N_18694,N_15408,N_14778);
nor U18695 (N_18695,N_14300,N_12512);
and U18696 (N_18696,N_12983,N_14478);
or U18697 (N_18697,N_14669,N_15331);
xor U18698 (N_18698,N_12709,N_13864);
xor U18699 (N_18699,N_13174,N_13491);
nor U18700 (N_18700,N_13172,N_14055);
or U18701 (N_18701,N_13835,N_12847);
nor U18702 (N_18702,N_12802,N_15429);
nor U18703 (N_18703,N_12603,N_12862);
nor U18704 (N_18704,N_12932,N_14435);
or U18705 (N_18705,N_15514,N_13137);
and U18706 (N_18706,N_13523,N_13787);
and U18707 (N_18707,N_13205,N_14582);
xor U18708 (N_18708,N_14296,N_13802);
xor U18709 (N_18709,N_14749,N_12824);
nor U18710 (N_18710,N_15525,N_15337);
xnor U18711 (N_18711,N_13847,N_14181);
and U18712 (N_18712,N_14970,N_14991);
nor U18713 (N_18713,N_15490,N_14161);
or U18714 (N_18714,N_14261,N_14123);
nand U18715 (N_18715,N_15251,N_15315);
nor U18716 (N_18716,N_14104,N_12809);
xnor U18717 (N_18717,N_14420,N_14156);
and U18718 (N_18718,N_12905,N_14107);
or U18719 (N_18719,N_14077,N_13727);
xor U18720 (N_18720,N_12736,N_13066);
and U18721 (N_18721,N_13827,N_14524);
nor U18722 (N_18722,N_15109,N_14559);
or U18723 (N_18723,N_14452,N_15338);
xnor U18724 (N_18724,N_13509,N_15086);
and U18725 (N_18725,N_12874,N_14565);
or U18726 (N_18726,N_14871,N_12731);
nor U18727 (N_18727,N_14864,N_13358);
nor U18728 (N_18728,N_15210,N_14599);
and U18729 (N_18729,N_14484,N_15466);
nor U18730 (N_18730,N_14607,N_13219);
nand U18731 (N_18731,N_14102,N_13237);
or U18732 (N_18732,N_13699,N_12721);
nand U18733 (N_18733,N_13735,N_14277);
and U18734 (N_18734,N_13665,N_14436);
or U18735 (N_18735,N_13517,N_13746);
xor U18736 (N_18736,N_13795,N_15418);
nand U18737 (N_18737,N_14617,N_14414);
nor U18738 (N_18738,N_13775,N_15340);
or U18739 (N_18739,N_12863,N_15135);
or U18740 (N_18740,N_12863,N_14244);
or U18741 (N_18741,N_12525,N_13294);
nor U18742 (N_18742,N_14162,N_14783);
nor U18743 (N_18743,N_13388,N_13027);
nand U18744 (N_18744,N_15608,N_15534);
or U18745 (N_18745,N_13743,N_15091);
or U18746 (N_18746,N_13141,N_15181);
nand U18747 (N_18747,N_14210,N_13799);
or U18748 (N_18748,N_15581,N_13060);
or U18749 (N_18749,N_13619,N_13279);
nand U18750 (N_18750,N_17826,N_17702);
nor U18751 (N_18751,N_16364,N_17788);
nor U18752 (N_18752,N_17723,N_16876);
or U18753 (N_18753,N_18418,N_16167);
and U18754 (N_18754,N_17738,N_16136);
or U18755 (N_18755,N_16893,N_15984);
and U18756 (N_18756,N_17841,N_16896);
xnor U18757 (N_18757,N_18312,N_16683);
nand U18758 (N_18758,N_17111,N_18195);
nor U18759 (N_18759,N_18506,N_15677);
or U18760 (N_18760,N_16731,N_16520);
xor U18761 (N_18761,N_16321,N_16479);
and U18762 (N_18762,N_17924,N_18318);
xor U18763 (N_18763,N_17072,N_18460);
nor U18764 (N_18764,N_17762,N_17995);
nand U18765 (N_18765,N_18438,N_17878);
and U18766 (N_18766,N_15747,N_18550);
nor U18767 (N_18767,N_16574,N_18415);
or U18768 (N_18768,N_18134,N_17750);
nand U18769 (N_18769,N_16898,N_18124);
nor U18770 (N_18770,N_17090,N_15988);
nor U18771 (N_18771,N_15830,N_16719);
nor U18772 (N_18772,N_16642,N_17716);
nand U18773 (N_18773,N_15741,N_18160);
xnor U18774 (N_18774,N_18332,N_18034);
or U18775 (N_18775,N_17401,N_18427);
xor U18776 (N_18776,N_16818,N_17134);
nor U18777 (N_18777,N_18327,N_17761);
nor U18778 (N_18778,N_16656,N_16016);
and U18779 (N_18779,N_15778,N_15683);
nand U18780 (N_18780,N_18029,N_18717);
nand U18781 (N_18781,N_16560,N_17264);
and U18782 (N_18782,N_16394,N_17317);
and U18783 (N_18783,N_16229,N_16933);
or U18784 (N_18784,N_17547,N_15963);
and U18785 (N_18785,N_17619,N_17038);
and U18786 (N_18786,N_18739,N_16852);
nand U18787 (N_18787,N_17412,N_18540);
xnor U18788 (N_18788,N_17026,N_18403);
nor U18789 (N_18789,N_16668,N_18191);
nor U18790 (N_18790,N_18702,N_17999);
or U18791 (N_18791,N_18388,N_16911);
nand U18792 (N_18792,N_18494,N_18263);
nand U18793 (N_18793,N_17964,N_17435);
nor U18794 (N_18794,N_15889,N_16410);
xor U18795 (N_18795,N_17551,N_17586);
or U18796 (N_18796,N_18436,N_18586);
and U18797 (N_18797,N_18012,N_17621);
nand U18798 (N_18798,N_16363,N_17543);
or U18799 (N_18799,N_17942,N_17955);
xor U18800 (N_18800,N_18073,N_16640);
and U18801 (N_18801,N_16472,N_15994);
and U18802 (N_18802,N_16102,N_18638);
nor U18803 (N_18803,N_17147,N_17060);
nand U18804 (N_18804,N_17468,N_18355);
nor U18805 (N_18805,N_18626,N_18059);
nand U18806 (N_18806,N_18202,N_17260);
and U18807 (N_18807,N_16908,N_17291);
nor U18808 (N_18808,N_17105,N_16807);
xor U18809 (N_18809,N_15877,N_15651);
nand U18810 (N_18810,N_16711,N_18306);
and U18811 (N_18811,N_16793,N_18634);
nand U18812 (N_18812,N_18534,N_18447);
nor U18813 (N_18813,N_16279,N_16502);
xor U18814 (N_18814,N_16559,N_17023);
and U18815 (N_18815,N_17922,N_17312);
nand U18816 (N_18816,N_17350,N_16270);
and U18817 (N_18817,N_16414,N_16493);
xor U18818 (N_18818,N_16018,N_18023);
or U18819 (N_18819,N_16643,N_17968);
nand U18820 (N_18820,N_16679,N_17570);
nor U18821 (N_18821,N_17882,N_16401);
xor U18822 (N_18822,N_16716,N_17909);
or U18823 (N_18823,N_17362,N_18591);
nand U18824 (N_18824,N_17216,N_18210);
nor U18825 (N_18825,N_17220,N_16914);
and U18826 (N_18826,N_17737,N_17657);
or U18827 (N_18827,N_16889,N_15645);
and U18828 (N_18828,N_16151,N_17289);
xnor U18829 (N_18829,N_16391,N_15855);
or U18830 (N_18830,N_17033,N_18461);
nor U18831 (N_18831,N_18641,N_16236);
nor U18832 (N_18832,N_17479,N_18685);
and U18833 (N_18833,N_16607,N_17717);
nor U18834 (N_18834,N_16968,N_16262);
and U18835 (N_18835,N_18176,N_17509);
nor U18836 (N_18836,N_16116,N_17607);
and U18837 (N_18837,N_18265,N_17673);
nor U18838 (N_18838,N_16326,N_15972);
or U18839 (N_18839,N_17608,N_16393);
nor U18840 (N_18840,N_18645,N_17976);
xor U18841 (N_18841,N_17648,N_15705);
or U18842 (N_18842,N_18162,N_16068);
xnor U18843 (N_18843,N_16517,N_15679);
xnor U18844 (N_18844,N_16282,N_15827);
nand U18845 (N_18845,N_17918,N_17348);
nand U18846 (N_18846,N_17649,N_17035);
and U18847 (N_18847,N_16745,N_18511);
and U18848 (N_18848,N_16095,N_15635);
or U18849 (N_18849,N_16214,N_16000);
and U18850 (N_18850,N_15694,N_15706);
xor U18851 (N_18851,N_17087,N_17425);
nand U18852 (N_18852,N_16781,N_16885);
and U18853 (N_18853,N_17981,N_18605);
nor U18854 (N_18854,N_17150,N_16727);
or U18855 (N_18855,N_16863,N_18635);
xnor U18856 (N_18856,N_16274,N_18393);
or U18857 (N_18857,N_16623,N_16589);
nand U18858 (N_18858,N_16961,N_17028);
or U18859 (N_18859,N_17246,N_16915);
xor U18860 (N_18860,N_18189,N_17498);
and U18861 (N_18861,N_17514,N_18678);
or U18862 (N_18862,N_17130,N_18343);
nor U18863 (N_18863,N_16402,N_17789);
or U18864 (N_18864,N_17001,N_18182);
nand U18865 (N_18865,N_18246,N_17945);
xnor U18866 (N_18866,N_16572,N_17893);
xnor U18867 (N_18867,N_18551,N_15886);
nor U18868 (N_18868,N_18425,N_16513);
nor U18869 (N_18869,N_18524,N_18688);
xor U18870 (N_18870,N_16843,N_16121);
xor U18871 (N_18871,N_16484,N_17987);
and U18872 (N_18872,N_15717,N_16604);
or U18873 (N_18873,N_17700,N_15755);
and U18874 (N_18874,N_18276,N_18479);
nor U18875 (N_18875,N_16421,N_16465);
nor U18876 (N_18876,N_15760,N_18649);
and U18877 (N_18877,N_18336,N_15836);
xor U18878 (N_18878,N_18086,N_17639);
or U18879 (N_18879,N_16239,N_16312);
or U18880 (N_18880,N_17019,N_16169);
and U18881 (N_18881,N_17424,N_16883);
xor U18882 (N_18882,N_17402,N_17617);
or U18883 (N_18883,N_16768,N_16750);
nand U18884 (N_18884,N_17475,N_15633);
nor U18885 (N_18885,N_15932,N_16432);
nand U18886 (N_18886,N_18274,N_15793);
or U18887 (N_18887,N_16669,N_17140);
and U18888 (N_18888,N_16746,N_16222);
or U18889 (N_18889,N_16844,N_18240);
xnor U18890 (N_18890,N_16228,N_17437);
xnor U18891 (N_18891,N_18552,N_17807);
or U18892 (N_18892,N_15891,N_17597);
and U18893 (N_18893,N_17025,N_16712);
or U18894 (N_18894,N_16037,N_16667);
or U18895 (N_18895,N_15869,N_18266);
and U18896 (N_18896,N_15680,N_16868);
or U18897 (N_18897,N_17017,N_18422);
nor U18898 (N_18898,N_16329,N_16995);
nor U18899 (N_18899,N_18308,N_17109);
xnor U18900 (N_18900,N_17040,N_17734);
xor U18901 (N_18901,N_18619,N_18219);
or U18902 (N_18902,N_18749,N_16980);
nor U18903 (N_18903,N_16390,N_17502);
nand U18904 (N_18904,N_16475,N_16760);
or U18905 (N_18905,N_18572,N_17940);
xnor U18906 (N_18906,N_15930,N_17281);
xor U18907 (N_18907,N_17912,N_16370);
nand U18908 (N_18908,N_17870,N_15941);
nor U18909 (N_18909,N_17201,N_18283);
nor U18910 (N_18910,N_15713,N_18163);
xnor U18911 (N_18911,N_15867,N_15900);
or U18912 (N_18912,N_16455,N_16543);
nand U18913 (N_18913,N_16459,N_18187);
and U18914 (N_18914,N_17011,N_15632);
or U18915 (N_18915,N_16259,N_17780);
and U18916 (N_18916,N_16869,N_18109);
nand U18917 (N_18917,N_16713,N_18245);
nand U18918 (N_18918,N_16237,N_17856);
nand U18919 (N_18919,N_16563,N_18106);
and U18920 (N_18920,N_16585,N_17373);
nand U18921 (N_18921,N_15859,N_16386);
nor U18922 (N_18922,N_18510,N_18734);
or U18923 (N_18923,N_18295,N_16693);
nand U18924 (N_18924,N_16248,N_18247);
xor U18925 (N_18925,N_16235,N_16346);
and U18926 (N_18926,N_17338,N_15879);
nor U18927 (N_18927,N_17352,N_15821);
or U18928 (N_18928,N_15749,N_15929);
nor U18929 (N_18929,N_16144,N_18065);
or U18930 (N_18930,N_16655,N_15654);
nand U18931 (N_18931,N_17499,N_16447);
xnor U18932 (N_18932,N_18742,N_15668);
xnor U18933 (N_18933,N_18133,N_17611);
and U18934 (N_18934,N_16216,N_17443);
nor U18935 (N_18935,N_16568,N_17899);
and U18936 (N_18936,N_18321,N_17655);
nand U18937 (N_18937,N_15686,N_15776);
or U18938 (N_18938,N_16650,N_17767);
nand U18939 (N_18939,N_17320,N_16878);
xor U18940 (N_18940,N_17549,N_16593);
or U18941 (N_18941,N_16184,N_15710);
or U18942 (N_18942,N_16641,N_17839);
and U18943 (N_18943,N_17745,N_18320);
xor U18944 (N_18944,N_16545,N_17451);
nand U18945 (N_18945,N_17828,N_18459);
nand U18946 (N_18946,N_18451,N_16498);
and U18947 (N_18947,N_17796,N_16612);
nand U18948 (N_18948,N_17292,N_15959);
xnor U18949 (N_18949,N_16610,N_17645);
nand U18950 (N_18950,N_16096,N_17198);
or U18951 (N_18951,N_16115,N_17076);
nand U18952 (N_18952,N_16174,N_15866);
nand U18953 (N_18953,N_17966,N_15913);
nand U18954 (N_18954,N_16483,N_17624);
or U18955 (N_18955,N_17152,N_16054);
and U18956 (N_18956,N_17178,N_18608);
nor U18957 (N_18957,N_15657,N_17861);
nand U18958 (N_18958,N_16306,N_18537);
nand U18959 (N_18959,N_15814,N_17715);
or U18960 (N_18960,N_17697,N_16118);
xor U18961 (N_18961,N_15802,N_16273);
nand U18962 (N_18962,N_18177,N_17548);
nor U18963 (N_18963,N_16130,N_16232);
xnor U18964 (N_18964,N_16419,N_18025);
nand U18965 (N_18965,N_17018,N_17578);
nor U18966 (N_18966,N_17824,N_16219);
or U18967 (N_18967,N_16891,N_17363);
or U18968 (N_18968,N_18428,N_18583);
and U18969 (N_18969,N_16895,N_16862);
xnor U18970 (N_18970,N_17869,N_16240);
xnor U18971 (N_18971,N_18179,N_17895);
xnor U18972 (N_18972,N_17851,N_18170);
xnor U18973 (N_18973,N_18502,N_16617);
nor U18974 (N_18974,N_16153,N_18450);
nand U18975 (N_18975,N_15810,N_15777);
nor U18976 (N_18976,N_17815,N_16110);
and U18977 (N_18977,N_18121,N_18030);
or U18978 (N_18978,N_15643,N_15779);
nand U18979 (N_18979,N_17757,N_16435);
nand U18980 (N_18980,N_18514,N_15722);
xnor U18981 (N_18981,N_17786,N_17431);
nor U18982 (N_18982,N_16725,N_18458);
nand U18983 (N_18983,N_17795,N_17167);
xor U18984 (N_18984,N_16085,N_17068);
xor U18985 (N_18985,N_18692,N_18464);
nand U18986 (N_18986,N_18492,N_16743);
and U18987 (N_18987,N_15895,N_17950);
nor U18988 (N_18988,N_15832,N_18720);
or U18989 (N_18989,N_17302,N_16556);
nor U18990 (N_18990,N_15730,N_17519);
nand U18991 (N_18991,N_16766,N_17127);
nand U18992 (N_18992,N_17539,N_15767);
and U18993 (N_18993,N_16361,N_16978);
and U18994 (N_18994,N_17599,N_15945);
nand U18995 (N_18995,N_17002,N_16139);
or U18996 (N_18996,N_17810,N_16382);
nand U18997 (N_18997,N_15809,N_15897);
nand U18998 (N_18998,N_16485,N_15907);
xor U18999 (N_18999,N_18171,N_17265);
nor U19000 (N_19000,N_17573,N_17961);
nand U19001 (N_19001,N_17095,N_16503);
xnor U19002 (N_19002,N_18212,N_17483);
and U19003 (N_19003,N_17565,N_15798);
or U19004 (N_19004,N_17615,N_17055);
nand U19005 (N_19005,N_17074,N_17531);
or U19006 (N_19006,N_17158,N_16998);
xor U19007 (N_19007,N_16443,N_16129);
or U19008 (N_19008,N_17943,N_18259);
nor U19009 (N_19009,N_16367,N_16417);
nand U19010 (N_19010,N_15919,N_16246);
or U19011 (N_19011,N_15999,N_17188);
and U19012 (N_19012,N_16645,N_16927);
xnor U19013 (N_19013,N_17347,N_15758);
nor U19014 (N_19014,N_17934,N_16358);
or U19015 (N_19015,N_15831,N_15634);
nand U19016 (N_19016,N_17914,N_18079);
and U19017 (N_19017,N_16708,N_16758);
nor U19018 (N_19018,N_15927,N_16302);
nand U19019 (N_19019,N_16072,N_16652);
nand U19020 (N_19020,N_17800,N_17142);
and U19021 (N_19021,N_15852,N_15974);
nand U19022 (N_19022,N_16964,N_18440);
nand U19023 (N_19023,N_18330,N_15762);
nand U19024 (N_19024,N_17058,N_16904);
nor U19025 (N_19025,N_18365,N_16431);
nand U19026 (N_19026,N_16910,N_18014);
nand U19027 (N_19027,N_18011,N_16280);
or U19028 (N_19028,N_16819,N_15716);
or U19029 (N_19029,N_17387,N_16829);
nand U19030 (N_19030,N_18527,N_17874);
and U19031 (N_19031,N_17679,N_18413);
nor U19032 (N_19032,N_16681,N_17891);
xor U19033 (N_19033,N_17181,N_18253);
nor U19034 (N_19034,N_16464,N_17064);
or U19035 (N_19035,N_18396,N_18571);
or U19036 (N_19036,N_17620,N_16586);
nor U19037 (N_19037,N_18594,N_16981);
or U19038 (N_19038,N_17277,N_18130);
and U19039 (N_19039,N_17637,N_18334);
or U19040 (N_19040,N_15922,N_16500);
nand U19041 (N_19041,N_16264,N_16848);
xor U19042 (N_19042,N_15688,N_15726);
and U19043 (N_19043,N_16395,N_16353);
nand U19044 (N_19044,N_16244,N_16297);
and U19045 (N_19045,N_18556,N_17664);
nor U19046 (N_19046,N_15640,N_16965);
xor U19047 (N_19047,N_16182,N_17034);
nand U19048 (N_19048,N_16303,N_17449);
xor U19049 (N_19049,N_16266,N_18693);
xor U19050 (N_19050,N_16113,N_15936);
xnor U19051 (N_19051,N_18603,N_18217);
or U19052 (N_19052,N_16813,N_16057);
or U19053 (N_19053,N_16835,N_16654);
or U19054 (N_19054,N_16373,N_18703);
xnor U19055 (N_19055,N_17677,N_16252);
and U19056 (N_19056,N_15955,N_16744);
nand U19057 (N_19057,N_16909,N_15977);
xor U19058 (N_19058,N_17252,N_18562);
xor U19059 (N_19059,N_18483,N_18260);
nand U19060 (N_19060,N_17385,N_18713);
nor U19061 (N_19061,N_17916,N_18710);
and U19062 (N_19062,N_18254,N_15638);
xnor U19063 (N_19063,N_17360,N_17335);
or U19064 (N_19064,N_17174,N_16079);
or U19065 (N_19065,N_18395,N_16810);
and U19066 (N_19066,N_16546,N_18015);
xor U19067 (N_19067,N_15976,N_15757);
xor U19068 (N_19068,N_17180,N_18357);
xnor U19069 (N_19069,N_17778,N_16374);
nor U19070 (N_19070,N_17144,N_17052);
xnor U19071 (N_19071,N_15813,N_16555);
xor U19072 (N_19072,N_15973,N_16518);
and U19073 (N_19073,N_18612,N_17334);
nand U19074 (N_19074,N_16529,N_17472);
and U19075 (N_19075,N_18663,N_17423);
xor U19076 (N_19076,N_18003,N_16991);
or U19077 (N_19077,N_18452,N_16164);
xor U19078 (N_19078,N_16434,N_15971);
nand U19079 (N_19079,N_17571,N_16659);
or U19080 (N_19080,N_17980,N_17609);
and U19081 (N_19081,N_17020,N_17651);
or U19082 (N_19082,N_17491,N_17092);
nand U19083 (N_19083,N_17836,N_18252);
nor U19084 (N_19084,N_16344,N_15650);
nand U19085 (N_19085,N_18640,N_16166);
xor U19086 (N_19086,N_17656,N_17868);
nor U19087 (N_19087,N_18190,N_17748);
nand U19088 (N_19088,N_16736,N_15829);
nand U19089 (N_19089,N_18430,N_16257);
xnor U19090 (N_19090,N_17821,N_17353);
nand U19091 (N_19091,N_16437,N_18261);
xnor U19092 (N_19092,N_18093,N_16770);
nor U19093 (N_19093,N_15873,N_17772);
nand U19094 (N_19094,N_18657,N_17618);
xnor U19095 (N_19095,N_17652,N_18414);
and U19096 (N_19096,N_17889,N_17930);
nor U19097 (N_19097,N_16782,N_15826);
or U19098 (N_19098,N_17217,N_18206);
nand U19099 (N_19099,N_17379,N_15735);
nor U19100 (N_19100,N_18486,N_17638);
nand U19101 (N_19101,N_16338,N_16777);
or U19102 (N_19102,N_15804,N_18397);
nor U19103 (N_19103,N_17230,N_17151);
or U19104 (N_19104,N_18662,N_17080);
or U19105 (N_19105,N_15625,N_16026);
xnor U19106 (N_19106,N_18083,N_16952);
and U19107 (N_19107,N_16564,N_18522);
nand U19108 (N_19108,N_17773,N_17414);
nor U19109 (N_19109,N_17952,N_17721);
and U19110 (N_19110,N_18225,N_17478);
nor U19111 (N_19111,N_16597,N_18238);
and U19112 (N_19112,N_16943,N_16613);
and U19113 (N_19113,N_16722,N_18362);
xnor U19114 (N_19114,N_16403,N_15950);
nand U19115 (N_19115,N_16696,N_18467);
nor U19116 (N_19116,N_18204,N_18021);
or U19117 (N_19117,N_15815,N_16396);
or U19118 (N_19118,N_18158,N_16124);
or U19119 (N_19119,N_15641,N_17753);
nor U19120 (N_19120,N_16140,N_17149);
and U19121 (N_19121,N_16408,N_16567);
xor U19122 (N_19122,N_17654,N_16028);
and U19123 (N_19123,N_15816,N_16019);
and U19124 (N_19124,N_18075,N_16931);
or U19125 (N_19125,N_15989,N_16734);
xor U19126 (N_19126,N_18383,N_16138);
or U19127 (N_19127,N_15653,N_18690);
or U19128 (N_19128,N_17703,N_15925);
nand U19129 (N_19129,N_17305,N_17865);
xnor U19130 (N_19130,N_17643,N_16993);
xor U19131 (N_19131,N_17915,N_16576);
and U19132 (N_19132,N_16089,N_18682);
xnor U19133 (N_19133,N_16425,N_17106);
nand U19134 (N_19134,N_16428,N_17207);
nand U19135 (N_19135,N_18542,N_17097);
xor U19136 (N_19136,N_16853,N_15631);
and U19137 (N_19137,N_18363,N_16786);
nand U19138 (N_19138,N_18076,N_18456);
and U19139 (N_19139,N_18315,N_16921);
and U19140 (N_19140,N_17481,N_15981);
or U19141 (N_19141,N_16263,N_16510);
nand U19142 (N_19142,N_16587,N_16206);
or U19143 (N_19143,N_16569,N_18544);
xnor U19144 (N_19144,N_16605,N_16788);
and U19145 (N_19145,N_15731,N_17537);
and U19146 (N_19146,N_17452,N_16724);
xor U19147 (N_19147,N_17453,N_16491);
and U19148 (N_19148,N_16951,N_17726);
and U19149 (N_19149,N_16918,N_17273);
nor U19150 (N_19150,N_18419,N_17794);
nand U19151 (N_19151,N_18251,N_17534);
or U19152 (N_19152,N_17120,N_18331);
xor U19153 (N_19153,N_16323,N_17860);
and U19154 (N_19154,N_18227,N_17577);
nor U19155 (N_19155,N_18304,N_15878);
or U19156 (N_19156,N_16762,N_16453);
and U19157 (N_19157,N_17085,N_18244);
and U19158 (N_19158,N_18490,N_16709);
xnor U19159 (N_19159,N_16354,N_16789);
nand U19160 (N_19160,N_16155,N_17495);
nand U19161 (N_19161,N_16997,N_18264);
xnor U19162 (N_19162,N_17262,N_18672);
nor U19163 (N_19163,N_17727,N_17683);
and U19164 (N_19164,N_17525,N_17770);
xor U19165 (N_19165,N_16371,N_16193);
xnor U19166 (N_19166,N_17706,N_17016);
nor U19167 (N_19167,N_17225,N_17696);
or U19168 (N_19168,N_16600,N_18126);
and U19169 (N_19169,N_16482,N_17634);
nand U19170 (N_19170,N_17971,N_17459);
or U19171 (N_19171,N_17200,N_15808);
or U19172 (N_19172,N_16183,N_16397);
and U19173 (N_19173,N_16226,N_15753);
xnor U19174 (N_19174,N_17078,N_15629);
and U19175 (N_19175,N_17689,N_15872);
xor U19176 (N_19176,N_17014,N_16439);
nand U19177 (N_19177,N_16454,N_16633);
nor U19178 (N_19178,N_18378,N_17880);
xnor U19179 (N_19179,N_17128,N_18463);
and U19180 (N_19180,N_17606,N_16937);
nor U19181 (N_19181,N_16767,N_16778);
and U19182 (N_19182,N_16119,N_18390);
xnor U19183 (N_19183,N_18153,N_17107);
nor U19184 (N_19184,N_16917,N_16553);
nand U19185 (N_19185,N_16084,N_17368);
nand U19186 (N_19186,N_17329,N_15956);
nand U19187 (N_19187,N_17659,N_17248);
nand U19188 (N_19188,N_16180,N_18590);
and U19189 (N_19189,N_17744,N_17194);
nand U19190 (N_19190,N_15910,N_15868);
nand U19191 (N_19191,N_16598,N_17015);
nor U19192 (N_19192,N_18684,N_16637);
nor U19193 (N_19193,N_17251,N_17859);
and U19194 (N_19194,N_16224,N_16143);
or U19195 (N_19195,N_17650,N_15765);
and U19196 (N_19196,N_18557,N_17122);
nand U19197 (N_19197,N_18437,N_18701);
xor U19198 (N_19198,N_18385,N_17195);
nor U19199 (N_19199,N_17269,N_16177);
nor U19200 (N_19200,N_16372,N_17285);
nand U19201 (N_19201,N_16456,N_17059);
nand U19202 (N_19202,N_16753,N_17141);
or U19203 (N_19203,N_17642,N_16957);
xor U19204 (N_19204,N_18518,N_15661);
nand U19205 (N_19205,N_17199,N_16653);
nand U19206 (N_19206,N_16627,N_16218);
nand U19207 (N_19207,N_16859,N_17872);
nand U19208 (N_19208,N_15708,N_18576);
or U19209 (N_19209,N_16197,N_18558);
nor U19210 (N_19210,N_17440,N_17990);
nor U19211 (N_19211,N_17843,N_16359);
nor U19212 (N_19212,N_16254,N_16635);
nand U19213 (N_19213,N_17210,N_16833);
xnor U19214 (N_19214,N_17678,N_18616);
or U19215 (N_19215,N_18407,N_15630);
nand U19216 (N_19216,N_15699,N_17300);
or U19217 (N_19217,N_16387,N_18356);
or U19218 (N_19218,N_15899,N_17049);
or U19219 (N_19219,N_15880,N_18444);
and U19220 (N_19220,N_18348,N_18653);
or U19221 (N_19221,N_17633,N_17829);
or U19222 (N_19222,N_18411,N_17675);
or U19223 (N_19223,N_17082,N_17827);
and U19224 (N_19224,N_16369,N_16191);
or U19225 (N_19225,N_18368,N_15796);
and U19226 (N_19226,N_16804,N_17250);
or U19227 (N_19227,N_18148,N_16301);
nand U19228 (N_19228,N_17792,N_15949);
xnor U19229 (N_19229,N_18392,N_18746);
or U19230 (N_19230,N_17729,N_16533);
nor U19231 (N_19231,N_16168,N_18166);
nand U19232 (N_19232,N_16021,N_16570);
or U19233 (N_19233,N_16058,N_15920);
nand U19234 (N_19234,N_17803,N_17900);
or U19235 (N_19235,N_17148,N_15754);
and U19236 (N_19236,N_17693,N_16541);
nand U19237 (N_19237,N_16832,N_16540);
and U19238 (N_19238,N_17948,N_15664);
and U19239 (N_19239,N_16514,N_17173);
or U19240 (N_19240,N_16692,N_17584);
and U19241 (N_19241,N_17243,N_17061);
nand U19242 (N_19242,N_17503,N_17755);
and U19243 (N_19243,N_18724,N_16606);
nor U19244 (N_19244,N_17600,N_16599);
nor U19245 (N_19245,N_17944,N_16106);
and U19246 (N_19246,N_17876,N_17351);
nand U19247 (N_19247,N_15906,N_15684);
nor U19248 (N_19248,N_18092,N_17844);
nor U19249 (N_19249,N_17388,N_16225);
nand U19250 (N_19250,N_17314,N_15719);
and U19251 (N_19251,N_17906,N_17904);
or U19252 (N_19252,N_18143,N_17834);
and U19253 (N_19253,N_15658,N_17086);
nor U19254 (N_19254,N_18664,N_17699);
and U19255 (N_19255,N_15805,N_18194);
xor U19256 (N_19256,N_16573,N_18373);
and U19257 (N_19257,N_16412,N_18301);
nor U19258 (N_19258,N_17817,N_17496);
nor U19259 (N_19259,N_16433,N_17647);
or U19260 (N_19260,N_18267,N_17129);
nand U19261 (N_19261,N_16362,N_18068);
xnor U19262 (N_19262,N_16196,N_17227);
and U19263 (N_19263,N_17469,N_16912);
xor U19264 (N_19264,N_16945,N_15933);
nor U19265 (N_19265,N_16710,N_17954);
nor U19266 (N_19266,N_16688,N_17073);
nand U19267 (N_19267,N_17886,N_16705);
nor U19268 (N_19268,N_17367,N_17456);
and U19269 (N_19269,N_18582,N_17439);
and U19270 (N_19270,N_18637,N_18528);
and U19271 (N_19271,N_17572,N_18051);
nor U19272 (N_19272,N_18446,N_18350);
and U19273 (N_19273,N_16020,N_17759);
xor U19274 (N_19274,N_17067,N_17233);
nand U19275 (N_19275,N_18229,N_16960);
or U19276 (N_19276,N_16043,N_16967);
or U19277 (N_19277,N_17177,N_16411);
xnor U19278 (N_19278,N_18449,N_15691);
nor U19279 (N_19279,N_17598,N_16318);
or U19280 (N_19280,N_18050,N_16671);
nor U19281 (N_19281,N_17413,N_16983);
or U19282 (N_19282,N_16448,N_17663);
xor U19283 (N_19283,N_18658,N_17298);
xnor U19284 (N_19284,N_16086,N_16595);
nand U19285 (N_19285,N_17371,N_16093);
and U19286 (N_19286,N_16537,N_18080);
xnor U19287 (N_19287,N_16004,N_18269);
xor U19288 (N_19288,N_16837,N_16827);
xnor U19289 (N_19289,N_17115,N_18366);
and U19290 (N_19290,N_16111,N_16165);
nor U19291 (N_19291,N_16160,N_18516);
and U19292 (N_19292,N_17937,N_17411);
and U19293 (N_19293,N_16689,N_18328);
or U19294 (N_19294,N_17546,N_17159);
xor U19295 (N_19295,N_18401,N_18213);
nand U19296 (N_19296,N_16081,N_16948);
and U19297 (N_19297,N_16256,N_15700);
and U19298 (N_19298,N_18201,N_16336);
nor U19299 (N_19299,N_16125,N_16581);
or U19300 (N_19300,N_18491,N_15985);
or U19301 (N_19301,N_16790,N_16060);
nor U19302 (N_19302,N_16249,N_18472);
nor U19303 (N_19303,N_18729,N_15946);
nand U19304 (N_19304,N_18135,N_17361);
and U19305 (N_19305,N_15892,N_17933);
nor U19306 (N_19306,N_17705,N_17286);
nand U19307 (N_19307,N_15828,N_16739);
nand U19308 (N_19308,N_16825,N_18017);
xnor U19309 (N_19309,N_18082,N_16839);
and U19310 (N_19310,N_17008,N_18453);
nand U19311 (N_19311,N_16065,N_18505);
xnor U19312 (N_19312,N_17467,N_18305);
or U19313 (N_19313,N_18358,N_18747);
or U19314 (N_19314,N_18705,N_17777);
xnor U19315 (N_19315,N_16012,N_16926);
or U19316 (N_19316,N_17027,N_17741);
and U19317 (N_19317,N_17206,N_16808);
nor U19318 (N_19318,N_17885,N_18655);
xor U19319 (N_19319,N_17113,N_18399);
xor U19320 (N_19320,N_15953,N_16011);
nand U19321 (N_19321,N_16854,N_16098);
nor U19322 (N_19322,N_16156,N_18500);
nor U19323 (N_19323,N_15665,N_16409);
nand U19324 (N_19324,N_17321,N_16399);
nand U19325 (N_19325,N_17172,N_16649);
or U19326 (N_19326,N_16154,N_16792);
and U19327 (N_19327,N_18154,N_16014);
or U19328 (N_19328,N_15662,N_16117);
or U19329 (N_19329,N_16071,N_18714);
nand U19330 (N_19330,N_15698,N_16773);
xnor U19331 (N_19331,N_17022,N_15853);
nand U19332 (N_19332,N_18055,N_17235);
and U19333 (N_19333,N_17377,N_16526);
and U19334 (N_19334,N_18044,N_17797);
or U19335 (N_19335,N_15928,N_16319);
or U19336 (N_19336,N_16732,N_16356);
nand U19337 (N_19337,N_17396,N_17879);
and U19338 (N_19338,N_17462,N_16398);
and U19339 (N_19339,N_18730,N_16077);
xor U19340 (N_19340,N_16523,N_18319);
and U19341 (N_19341,N_17395,N_17290);
xor U19342 (N_19342,N_16210,N_16657);
and U19343 (N_19343,N_16720,N_18181);
and U19344 (N_19344,N_17667,N_17374);
nand U19345 (N_19345,N_16986,N_18062);
and U19346 (N_19346,N_15871,N_18732);
and U19347 (N_19347,N_18149,N_17186);
and U19348 (N_19348,N_16406,N_17581);
or U19349 (N_19349,N_17062,N_17114);
nand U19350 (N_19350,N_15750,N_15885);
nor U19351 (N_19351,N_18642,N_17613);
nor U19352 (N_19352,N_17820,N_17877);
xnor U19353 (N_19353,N_18131,N_17108);
xor U19354 (N_19354,N_18043,N_18435);
and U19355 (N_19355,N_16186,N_16310);
nand U19356 (N_19356,N_16806,N_17641);
or U19357 (N_19357,N_18666,N_16188);
nand U19358 (N_19358,N_17470,N_15770);
nor U19359 (N_19359,N_15942,N_17466);
and U19360 (N_19360,N_17687,N_18627);
xor U19361 (N_19361,N_17610,N_17690);
and U19362 (N_19362,N_17189,N_18644);
nand U19363 (N_19363,N_16881,N_17063);
nor U19364 (N_19364,N_17998,N_16953);
or U19365 (N_19365,N_16330,N_17187);
nand U19366 (N_19366,N_18207,N_16471);
or U19367 (N_19367,N_18167,N_17962);
and U19368 (N_19368,N_17110,N_15898);
or U19369 (N_19369,N_18499,N_16938);
nor U19370 (N_19370,N_18371,N_17994);
xnor U19371 (N_19371,N_17383,N_17037);
or U19372 (N_19372,N_16954,N_17967);
and U19373 (N_19373,N_16048,N_18578);
or U19374 (N_19374,N_18024,N_16247);
or U19375 (N_19375,N_17400,N_18027);
xor U19376 (N_19376,N_18628,N_18683);
nor U19377 (N_19377,N_17604,N_16234);
nor U19378 (N_19378,N_17709,N_17562);
nand U19379 (N_19379,N_16803,N_17763);
and U19380 (N_19380,N_16440,N_17735);
or U19381 (N_19381,N_15952,N_17722);
nor U19382 (N_19382,N_17579,N_16161);
nor U19383 (N_19383,N_15948,N_16664);
and U19384 (N_19384,N_16561,N_17626);
and U19385 (N_19385,N_16622,N_16624);
nand U19386 (N_19386,N_18335,N_15714);
nand U19387 (N_19387,N_17508,N_17211);
and U19388 (N_19388,N_15794,N_18631);
nor U19389 (N_19389,N_16094,N_17328);
xnor U19390 (N_19390,N_18369,N_15783);
nand U19391 (N_19391,N_18727,N_15784);
or U19392 (N_19392,N_18144,N_16052);
nand U19393 (N_19393,N_16384,N_16067);
nand U19394 (N_19394,N_16939,N_18741);
and U19395 (N_19395,N_17595,N_16673);
xnor U19396 (N_19396,N_17517,N_16714);
nor U19397 (N_19397,N_15962,N_17365);
and U19398 (N_19398,N_16101,N_18344);
xor U19399 (N_19399,N_18237,N_18049);
nand U19400 (N_19400,N_17589,N_17871);
xnor U19401 (N_19401,N_17685,N_16871);
nor U19402 (N_19402,N_16422,N_16504);
and U19403 (N_19403,N_18735,N_17771);
nor U19404 (N_19404,N_17244,N_16780);
xnor U19405 (N_19405,N_17021,N_17561);
nand U19406 (N_19406,N_18429,N_18271);
and U19407 (N_19407,N_16864,N_16628);
xnor U19408 (N_19408,N_17887,N_18047);
nor U19409 (N_19409,N_16126,N_17858);
or U19410 (N_19410,N_16776,N_17331);
xnor U19411 (N_19411,N_15991,N_17297);
and U19412 (N_19412,N_17941,N_18375);
and U19413 (N_19413,N_17830,N_17775);
and U19414 (N_19414,N_18299,N_18743);
xor U19415 (N_19415,N_18119,N_17345);
nor U19416 (N_19416,N_17972,N_17309);
xnor U19417 (N_19417,N_17131,N_16571);
or U19418 (N_19418,N_16293,N_18367);
or U19419 (N_19419,N_15642,N_16579);
nor U19420 (N_19420,N_16053,N_16035);
xor U19421 (N_19421,N_17714,N_16083);
nand U19422 (N_19422,N_16947,N_17989);
or U19423 (N_19423,N_16036,N_16665);
xnor U19424 (N_19424,N_16499,N_17484);
and U19425 (N_19425,N_18533,N_17724);
nand U19426 (N_19426,N_18535,N_16047);
nand U19427 (N_19427,N_16858,N_16304);
or U19428 (N_19428,N_16337,N_18323);
and U19429 (N_19429,N_17894,N_17963);
xnor U19430 (N_19430,N_17319,N_18748);
or U19431 (N_19431,N_16278,N_17644);
or U19432 (N_19432,N_16087,N_18477);
and U19433 (N_19433,N_18620,N_18338);
or U19434 (N_19434,N_16879,N_18156);
xnor U19435 (N_19435,N_17736,N_16929);
or U19436 (N_19436,N_17669,N_17516);
or U19437 (N_19437,N_18432,N_18374);
nor U19438 (N_19438,N_17223,N_17168);
nand U19439 (N_19439,N_18096,N_16761);
or U19440 (N_19440,N_18513,N_16255);
nor U19441 (N_19441,N_17263,N_18337);
and U19442 (N_19442,N_17280,N_16870);
xor U19443 (N_19443,N_16040,N_18009);
xor U19444 (N_19444,N_16486,N_15782);
nor U19445 (N_19445,N_18676,N_17593);
nand U19446 (N_19446,N_17357,N_16342);
or U19447 (N_19447,N_18455,N_18412);
and U19448 (N_19448,N_17071,N_18007);
nor U19449 (N_19449,N_15882,N_15720);
nand U19450 (N_19450,N_18708,N_16481);
and U19451 (N_19451,N_16001,N_18208);
xor U19452 (N_19452,N_16480,N_15655);
nand U19453 (N_19453,N_17162,N_18005);
and U19454 (N_19454,N_16056,N_16441);
xor U19455 (N_19455,N_17682,N_18512);
nand U19456 (N_19456,N_16349,N_17668);
xor U19457 (N_19457,N_17804,N_17370);
or U19458 (N_19458,N_16756,N_16730);
or U19459 (N_19459,N_17179,N_17196);
xor U19460 (N_19460,N_15840,N_18013);
xnor U19461 (N_19461,N_18570,N_15711);
or U19462 (N_19462,N_16488,N_17240);
and U19463 (N_19463,N_18120,N_17234);
xor U19464 (N_19464,N_17614,N_17428);
xor U19465 (N_19465,N_15786,N_16701);
nor U19466 (N_19466,N_17204,N_18740);
nor U19467 (N_19467,N_16063,N_17996);
nand U19468 (N_19468,N_18697,N_18173);
or U19469 (N_19469,N_15672,N_18040);
xnor U19470 (N_19470,N_15801,N_17982);
nor U19471 (N_19471,N_18698,N_18707);
xnor U19472 (N_19472,N_15666,N_16888);
and U19473 (N_19473,N_17327,N_15893);
nor U19474 (N_19474,N_16307,N_18509);
xor U19475 (N_19475,N_17698,N_17304);
or U19476 (N_19476,N_16830,N_15835);
nand U19477 (N_19477,N_17203,N_15964);
xor U19478 (N_19478,N_17631,N_17118);
nand U19479 (N_19479,N_18370,N_17661);
xor U19480 (N_19480,N_16305,N_16192);
nor U19481 (N_19481,N_17190,N_17523);
xnor U19482 (N_19482,N_18292,N_16314);
xor U19483 (N_19483,N_16751,N_15792);
nand U19484 (N_19484,N_15939,N_15785);
or U19485 (N_19485,N_17536,N_18175);
nand U19486 (N_19486,N_17461,N_17533);
nand U19487 (N_19487,N_17433,N_16894);
or U19488 (N_19488,N_18039,N_18289);
xnor U19489 (N_19489,N_15669,N_16666);
or U19490 (N_19490,N_16271,N_18584);
and U19491 (N_19491,N_15903,N_18072);
xor U19492 (N_19492,N_17084,N_16509);
or U19493 (N_19493,N_17849,N_18630);
xor U19494 (N_19494,N_16109,N_18656);
nor U19495 (N_19495,N_18497,N_15844);
xnor U19496 (N_19496,N_16963,N_16860);
nor U19497 (N_19497,N_18716,N_16544);
and U19498 (N_19498,N_16979,N_18585);
or U19499 (N_19499,N_17791,N_17494);
nand U19500 (N_19500,N_17936,N_17378);
and U19501 (N_19501,N_18745,N_17896);
or U19502 (N_19502,N_17294,N_16771);
nor U19503 (N_19503,N_18632,N_18361);
nor U19504 (N_19504,N_18224,N_16051);
nand U19505 (N_19505,N_18000,N_15969);
or U19506 (N_19506,N_16846,N_17296);
xor U19507 (N_19507,N_16333,N_17926);
and U19508 (N_19508,N_16010,N_16973);
nand U19509 (N_19509,N_16882,N_17339);
nor U19510 (N_19510,N_17733,N_17783);
nand U19511 (N_19511,N_16385,N_17500);
xnor U19512 (N_19512,N_16340,N_18196);
nand U19513 (N_19513,N_16251,N_17184);
and U19514 (N_19514,N_18185,N_17507);
and U19515 (N_19515,N_17145,N_15732);
nor U19516 (N_19516,N_18670,N_16389);
nand U19517 (N_19517,N_16824,N_17254);
nor U19518 (N_19518,N_16836,N_17492);
and U19519 (N_19519,N_17566,N_16327);
nand U19520 (N_19520,N_17801,N_16042);
or U19521 (N_19521,N_17161,N_17231);
nor U19522 (N_19522,N_17039,N_16325);
nand U19523 (N_19523,N_18737,N_17532);
and U19524 (N_19524,N_18574,N_16250);
or U19525 (N_19525,N_16258,N_16033);
xor U19526 (N_19526,N_15850,N_15769);
xor U19527 (N_19527,N_17256,N_16783);
nand U19528 (N_19528,N_18617,N_17694);
nand U19529 (N_19529,N_17983,N_17742);
and U19530 (N_19530,N_17047,N_18089);
or U19531 (N_19531,N_16286,N_17299);
nand U19532 (N_19532,N_16718,N_17057);
xor U19533 (N_19533,N_18526,N_17261);
xor U19534 (N_19534,N_16516,N_16515);
or U19535 (N_19535,N_16703,N_17044);
xor U19536 (N_19536,N_18132,N_18699);
or U19537 (N_19537,N_17557,N_17446);
nand U19538 (N_19538,N_16950,N_16388);
and U19539 (N_19539,N_16212,N_16469);
and U19540 (N_19540,N_17432,N_17544);
xor U19541 (N_19541,N_18643,N_18046);
nor U19542 (N_19542,N_18112,N_17825);
and U19543 (N_19543,N_17501,N_18232);
nand U19544 (N_19544,N_15693,N_18138);
nand U19545 (N_19545,N_17308,N_15675);
xor U19546 (N_19546,N_16764,N_18476);
nand U19547 (N_19547,N_18462,N_17487);
nor U19548 (N_19548,N_15659,N_18151);
nor U19549 (N_19549,N_16317,N_17382);
and U19550 (N_19550,N_17066,N_17069);
or U19551 (N_19551,N_16204,N_18016);
or U19552 (N_19552,N_15862,N_15743);
and U19553 (N_19553,N_16122,N_18115);
nand U19554 (N_19554,N_16069,N_17725);
or U19555 (N_19555,N_17707,N_17903);
xnor U19556 (N_19556,N_16243,N_16413);
xnor U19557 (N_19557,N_16070,N_17458);
nand U19558 (N_19558,N_17070,N_16242);
nand U19559 (N_19559,N_15627,N_17665);
or U19560 (N_19560,N_17245,N_18045);
and U19561 (N_19561,N_16884,N_16566);
nor U19562 (N_19562,N_18549,N_15674);
nor U19563 (N_19563,N_17182,N_15670);
xnor U19564 (N_19564,N_18704,N_16674);
and U19565 (N_19565,N_16506,N_16900);
or U19566 (N_19566,N_17538,N_18316);
and U19567 (N_19567,N_16091,N_18161);
or U19568 (N_19568,N_17088,N_16834);
nand U19569 (N_19569,N_17282,N_15812);
nor U19570 (N_19570,N_17576,N_16463);
xor U19571 (N_19571,N_17776,N_16763);
nand U19572 (N_19572,N_18592,N_15917);
xnor U19573 (N_19573,N_16670,N_17442);
or U19574 (N_19574,N_17818,N_15756);
xor U19575 (N_19575,N_15915,N_18481);
xor U19576 (N_19576,N_18575,N_18382);
or U19577 (N_19577,N_16857,N_17864);
or U19578 (N_19578,N_16988,N_16733);
xnor U19579 (N_19579,N_17853,N_18278);
and U19580 (N_19580,N_16064,N_18031);
nand U19581 (N_19581,N_16611,N_17628);
xnor U19582 (N_19582,N_16474,N_17582);
or U19583 (N_19583,N_16691,N_16602);
and U19584 (N_19584,N_16097,N_17713);
nor U19585 (N_19585,N_15807,N_16352);
or U19586 (N_19586,N_18493,N_17552);
nor U19587 (N_19587,N_16287,N_15825);
and U19588 (N_19588,N_18104,N_16535);
xor U19589 (N_19589,N_16420,N_18680);
or U19590 (N_19590,N_17146,N_16851);
nor U19591 (N_19591,N_16976,N_16936);
or U19592 (N_19592,N_16845,N_17806);
nor U19593 (N_19593,N_18689,N_18587);
or U19594 (N_19594,N_15967,N_16039);
or U19595 (N_19595,N_16694,N_17104);
nand U19596 (N_19596,N_18297,N_17793);
xnor U19597 (N_19597,N_16742,N_18116);
xnor U19598 (N_19598,N_17041,N_18482);
and U19599 (N_19599,N_15771,N_16350);
or U19600 (N_19600,N_16288,N_15663);
xor U19601 (N_19601,N_17752,N_17143);
xnor U19602 (N_19602,N_17119,N_16355);
or U19603 (N_19603,N_17512,N_15884);
and U19604 (N_19604,N_16496,N_18281);
and U19605 (N_19605,N_15854,N_17306);
nor U19606 (N_19606,N_18300,N_17855);
or U19607 (N_19607,N_16201,N_18648);
or U19608 (N_19608,N_18174,N_16632);
or U19609 (N_19609,N_16195,N_17731);
and U19610 (N_19610,N_18424,N_17408);
nand U19611 (N_19611,N_17493,N_17096);
xnor U19612 (N_19612,N_18063,N_16822);
and U19613 (N_19613,N_16376,N_16146);
xor U19614 (N_19614,N_16436,N_17154);
or U19615 (N_19615,N_18223,N_15921);
xnor U19616 (N_19616,N_18380,N_17278);
nand U19617 (N_19617,N_18032,N_16285);
nand U19618 (N_19618,N_15997,N_17505);
and U19619 (N_19619,N_16661,N_17330);
or U19620 (N_19620,N_17875,N_18387);
xnor U19621 (N_19621,N_16932,N_15875);
xor U19622 (N_19622,N_17956,N_15839);
and U19623 (N_19623,N_18545,N_16940);
or U19624 (N_19624,N_16697,N_18052);
nand U19625 (N_19625,N_18111,N_16609);
nor U19626 (N_19626,N_15724,N_15865);
and U19627 (N_19627,N_16639,N_16817);
nor U19628 (N_19628,N_16024,N_16294);
xor U19629 (N_19629,N_15744,N_18468);
or U19630 (N_19630,N_16123,N_16038);
xnor U19631 (N_19631,N_16508,N_16539);
nor U19632 (N_19632,N_16577,N_16404);
xor U19633 (N_19633,N_17126,N_16728);
xor U19634 (N_19634,N_17460,N_17588);
nand U19635 (N_19635,N_15646,N_16542);
or U19636 (N_19636,N_15781,N_17958);
xor U19637 (N_19637,N_17065,N_17054);
or U19638 (N_19638,N_16241,N_15966);
and U19639 (N_19639,N_16253,N_17947);
nor U19640 (N_19640,N_15811,N_16647);
nor U19641 (N_19641,N_16008,N_16737);
nor U19642 (N_19642,N_17692,N_16322);
or U19643 (N_19643,N_15733,N_17091);
xor U19644 (N_19644,N_15628,N_16217);
or U19645 (N_19645,N_17921,N_16076);
or U19646 (N_19646,N_16132,N_18523);
and U19647 (N_19647,N_17953,N_16687);
nand U19648 (N_19648,N_17323,N_17545);
or U19649 (N_19649,N_17268,N_15704);
nor U19650 (N_19650,N_16663,N_16552);
or U19651 (N_19651,N_16849,N_18606);
xor U19652 (N_19652,N_16582,N_16227);
or U19653 (N_19653,N_17212,N_16027);
nand U19654 (N_19654,N_18147,N_16044);
nand U19655 (N_19655,N_16801,N_17226);
nand U19656 (N_19656,N_18561,N_16230);
nand U19657 (N_19657,N_17224,N_17768);
and U19658 (N_19658,N_16575,N_17811);
or U19659 (N_19659,N_16855,N_16261);
or U19660 (N_19660,N_18006,N_17311);
nand U19661 (N_19661,N_18114,N_16658);
nor U19662 (N_19662,N_17553,N_18394);
nor U19663 (N_19663,N_15687,N_18398);
nor U19664 (N_19664,N_15689,N_18110);
and U19665 (N_19665,N_16009,N_16041);
nor U19666 (N_19666,N_17823,N_16706);
or U19667 (N_19667,N_16774,N_17192);
and U19668 (N_19668,N_16892,N_18026);
nand U19669 (N_19669,N_18478,N_18661);
and U19670 (N_19670,N_16357,N_17612);
nand U19671 (N_19671,N_18618,N_18203);
and U19672 (N_19672,N_16551,N_17288);
and U19673 (N_19673,N_16994,N_16461);
nor U19674 (N_19674,N_16797,N_17480);
xor U19675 (N_19675,N_18102,N_16334);
xor U19676 (N_19676,N_16614,N_15938);
or U19677 (N_19677,N_15676,N_17436);
xor U19678 (N_19678,N_17170,N_18101);
nand U19679 (N_19679,N_18205,N_15861);
and U19680 (N_19680,N_17366,N_16494);
and U19681 (N_19681,N_18262,N_17814);
xor U19682 (N_19682,N_15718,N_15648);
nor U19683 (N_19683,N_17185,N_15970);
xnor U19684 (N_19684,N_16313,N_15819);
nand U19685 (N_19685,N_16890,N_16202);
and U19686 (N_19686,N_15834,N_17518);
nor U19687 (N_19687,N_16175,N_17482);
nand U19688 (N_19688,N_17751,N_16366);
xnor U19689 (N_19689,N_16935,N_17310);
or U19690 (N_19690,N_16631,N_17929);
nand U19691 (N_19691,N_18569,N_18277);
xor U19692 (N_19692,N_16532,N_16831);
or U19693 (N_19693,N_17005,N_17012);
and U19694 (N_19694,N_16149,N_18035);
or U19695 (N_19695,N_18381,N_18573);
xnor U19696 (N_19696,N_18193,N_17010);
nand U19697 (N_19697,N_17564,N_15738);
nand U19698 (N_19698,N_18665,N_18667);
and U19699 (N_19699,N_16172,N_18433);
and U19700 (N_19700,N_15681,N_16548);
and U19701 (N_19701,N_17583,N_18674);
and U19702 (N_19702,N_18726,N_18353);
or U19703 (N_19703,N_16620,N_18159);
nor U19704 (N_19704,N_17625,N_17528);
nor U19705 (N_19705,N_18081,N_17602);
and U19706 (N_19706,N_15846,N_15944);
xor U19707 (N_19707,N_16368,N_17325);
or U19708 (N_19708,N_16189,N_17024);
nor U19709 (N_19709,N_15721,N_17477);
nand U19710 (N_19710,N_16176,N_17550);
xor U19711 (N_19711,N_16867,N_18287);
or U19712 (N_19712,N_16816,N_16157);
or U19713 (N_19713,N_18360,N_16626);
nand U19714 (N_19714,N_18445,N_18070);
nand U19715 (N_19715,N_18498,N_17077);
nand U19716 (N_19716,N_18199,N_16906);
and U19717 (N_19717,N_17464,N_17782);
xor U19718 (N_19718,N_17951,N_16208);
nor U19719 (N_19719,N_17993,N_18744);
nand U19720 (N_19720,N_15797,N_17653);
or U19721 (N_19721,N_18736,N_18474);
xnor U19722 (N_19722,N_16785,N_15914);
nor U19723 (N_19723,N_18695,N_16949);
and U19724 (N_19724,N_17209,N_15702);
xor U19725 (N_19725,N_18728,N_16442);
xnor U19726 (N_19726,N_15857,N_16073);
nand U19727 (N_19727,N_18673,N_15736);
and U19728 (N_19728,N_16025,N_18094);
nand U19729 (N_19729,N_17985,N_18400);
and U19730 (N_19730,N_17988,N_15685);
nand U19731 (N_19731,N_17000,N_18568);
xor U19732 (N_19732,N_16120,N_16791);
nand U19733 (N_19733,N_18484,N_17473);
nor U19734 (N_19734,N_18077,N_17042);
nand U19735 (N_19735,N_16203,N_15723);
nand U19736 (N_19736,N_16992,N_16821);
and U19737 (N_19737,N_18431,N_18507);
or U19738 (N_19738,N_17594,N_17276);
xor U19739 (N_19739,N_17555,N_15975);
nor U19740 (N_19740,N_18496,N_16899);
nor U19741 (N_19741,N_17622,N_16444);
nand U19742 (N_19742,N_18091,N_17816);
nand U19743 (N_19743,N_17798,N_16090);
or U19744 (N_19744,N_18563,N_15739);
or U19745 (N_19745,N_17883,N_17949);
xor U19746 (N_19746,N_18508,N_18053);
and U19747 (N_19747,N_17045,N_15842);
and U19748 (N_19748,N_15695,N_18671);
nand U19749 (N_19749,N_16380,N_15911);
nand U19750 (N_19750,N_16467,N_18614);
xor U19751 (N_19751,N_16608,N_17228);
nor U19752 (N_19752,N_16128,N_16678);
nand U19753 (N_19753,N_18351,N_17342);
nand U19754 (N_19754,N_16339,N_17463);
or U19755 (N_19755,N_17931,N_17728);
nor U19756 (N_19756,N_18409,N_18184);
nor U19757 (N_19757,N_15881,N_17236);
or U19758 (N_19758,N_18625,N_18426);
nor U19759 (N_19759,N_16591,N_16695);
xor U19760 (N_19760,N_17979,N_16487);
xor U19761 (N_19761,N_18107,N_17009);
nand U19762 (N_19762,N_17403,N_15795);
xnor U19763 (N_19763,N_16215,N_16648);
and U19764 (N_19764,N_18633,N_16159);
and U19765 (N_19765,N_18293,N_18218);
or U19766 (N_19766,N_17157,N_18503);
xnor U19767 (N_19767,N_16100,N_18346);
xnor U19768 (N_19768,N_18298,N_18566);
and U19769 (N_19769,N_16531,N_18249);
or U19770 (N_19770,N_18341,N_17785);
xor U19771 (N_19771,N_15800,N_17506);
nand U19772 (N_19772,N_15979,N_18530);
xor U19773 (N_19773,N_18311,N_16826);
nor U19774 (N_19774,N_17407,N_17790);
nand U19775 (N_19775,N_18303,N_16820);
nor U19776 (N_19776,N_17574,N_17765);
or U19777 (N_19777,N_16114,N_18529);
and U19778 (N_19778,N_15924,N_17081);
xor U19779 (N_19779,N_18242,N_17917);
or U19780 (N_19780,N_17902,N_17191);
xnor U19781 (N_19781,N_18723,N_16796);
and U19782 (N_19782,N_18349,N_17781);
or U19783 (N_19783,N_15715,N_18694);
nand U19784 (N_19784,N_17392,N_18127);
or U19785 (N_19785,N_17427,N_18228);
nor U19786 (N_19786,N_16179,N_15772);
or U19787 (N_19787,N_16971,N_17701);
or U19788 (N_19788,N_16928,N_16185);
nand U19789 (N_19789,N_15822,N_18243);
nand U19790 (N_19790,N_18543,N_17939);
nand U19791 (N_19791,N_16596,N_16275);
nand U19792 (N_19792,N_17333,N_15951);
xor U19793 (N_19793,N_15787,N_16787);
or U19794 (N_19794,N_16220,N_17671);
and U19795 (N_19795,N_16536,N_16430);
xor U19796 (N_19796,N_16377,N_18711);
xor U19797 (N_19797,N_18377,N_18333);
or U19798 (N_19798,N_18078,N_17831);
xor U19799 (N_19799,N_18098,N_16934);
or U19800 (N_19800,N_15707,N_16429);
or U19801 (N_19801,N_17799,N_17504);
and U19802 (N_19802,N_18183,N_18454);
nand U19803 (N_19803,N_17984,N_18391);
or U19804 (N_19804,N_16924,N_16805);
nand U19805 (N_19805,N_15918,N_17476);
and U19806 (N_19806,N_17603,N_17166);
xnor U19807 (N_19807,N_18565,N_17666);
xnor U19808 (N_19808,N_17580,N_17708);
or U19809 (N_19809,N_18639,N_17629);
and U19810 (N_19810,N_17336,N_18372);
xnor U19811 (N_19811,N_16729,N_17524);
and U19812 (N_19812,N_16495,N_17386);
or U19813 (N_19813,N_16209,N_16944);
and U19814 (N_19814,N_16977,N_17832);
and U19815 (N_19815,N_16717,N_17324);
and U19816 (N_19816,N_18042,N_16309);
and U19817 (N_19817,N_16618,N_18597);
or U19818 (N_19818,N_18125,N_18652);
nand U19819 (N_19819,N_16558,N_17416);
and U19820 (N_19820,N_15940,N_16901);
or U19821 (N_19821,N_16341,N_16903);
or U19822 (N_19822,N_15763,N_18231);
or U19823 (N_19823,N_15934,N_17837);
xnor U19824 (N_19824,N_17249,N_16281);
or U19825 (N_19825,N_17747,N_18469);
nor U19826 (N_19826,N_18686,N_18041);
or U19827 (N_19827,N_18290,N_16741);
nor U19828 (N_19828,N_16534,N_17556);
or U19829 (N_19829,N_16913,N_18589);
nor U19830 (N_19830,N_16625,N_17630);
nor U19831 (N_19831,N_17410,N_18064);
nand U19832 (N_19832,N_18105,N_16171);
nand U19833 (N_19833,N_18439,N_18019);
and U19834 (N_19834,N_16872,N_17712);
or U19835 (N_19835,N_17169,N_17419);
or U19836 (N_19836,N_17965,N_16823);
xor U19837 (N_19837,N_18157,N_18291);
nand U19838 (N_19838,N_16765,N_17691);
xor U19839 (N_19839,N_15775,N_17585);
xor U19840 (N_19840,N_16426,N_18004);
nand U19841 (N_19841,N_15843,N_16320);
nand U19842 (N_19842,N_18647,N_16880);
nor U19843 (N_19843,N_17938,N_16989);
xnor U19844 (N_19844,N_16137,N_18473);
xnor U19845 (N_19845,N_17520,N_16062);
xor U19846 (N_19846,N_16446,N_16017);
or U19847 (N_19847,N_18056,N_16985);
nand U19848 (N_19848,N_18519,N_18410);
xor U19849 (N_19849,N_17927,N_16549);
xor U19850 (N_19850,N_17754,N_15740);
nand U19851 (N_19851,N_15671,N_18417);
nand U19852 (N_19852,N_18434,N_16505);
nand U19853 (N_19853,N_18309,N_16375);
and U19854 (N_19854,N_16061,N_16704);
nor U19855 (N_19855,N_18317,N_16152);
and U19856 (N_19856,N_17526,N_18018);
nand U19857 (N_19857,N_17672,N_15965);
nor U19858 (N_19858,N_17591,N_17563);
xnor U19859 (N_19859,N_18057,N_15848);
nand U19860 (N_19860,N_16772,N_16972);
nor U19861 (N_19861,N_15729,N_17089);
and U19862 (N_19862,N_15728,N_15851);
nand U19863 (N_19863,N_17138,N_17541);
or U19864 (N_19864,N_17704,N_16749);
nor U19865 (N_19865,N_18197,N_16887);
nand U19866 (N_19866,N_17632,N_16400);
and U19867 (N_19867,N_17784,N_17222);
nand U19868 (N_19868,N_15626,N_17394);
xnor U19869 (N_19869,N_17406,N_16562);
or U19870 (N_19870,N_16295,N_17959);
nand U19871 (N_19871,N_18718,N_16181);
and U19872 (N_19872,N_16970,N_15864);
nor U19873 (N_19873,N_18379,N_15682);
xnor U19874 (N_19874,N_18200,N_15993);
nand U19875 (N_19875,N_15947,N_16748);
or U19876 (N_19876,N_16594,N_17218);
or U19877 (N_19877,N_17135,N_17344);
and U19878 (N_19878,N_17910,N_16584);
nand U19879 (N_19879,N_18129,N_15961);
and U19880 (N_19880,N_15734,N_17590);
and U19881 (N_19881,N_17376,N_16757);
nor U19882 (N_19882,N_18141,N_16006);
or U19883 (N_19883,N_17711,N_15902);
xor U19884 (N_19884,N_18342,N_17710);
nor U19885 (N_19885,N_18280,N_16987);
nand U19886 (N_19886,N_17340,N_18001);
or U19887 (N_19887,N_18485,N_16296);
nor U19888 (N_19888,N_17587,N_17287);
nand U19889 (N_19889,N_18465,N_17838);
or U19890 (N_19890,N_16424,N_17053);
and U19891 (N_19891,N_18646,N_17974);
or U19892 (N_19892,N_16755,N_15943);
and U19893 (N_19893,N_15637,N_18307);
or U19894 (N_19894,N_16328,N_17862);
nor U19895 (N_19895,N_17102,N_15712);
or U19896 (N_19896,N_18443,N_16002);
xor U19897 (N_19897,N_17718,N_15876);
or U19898 (N_19898,N_16205,N_16798);
or U19899 (N_19899,N_15978,N_17051);
or U19900 (N_19900,N_18488,N_15995);
and U19901 (N_19901,N_16416,N_18475);
nand U19902 (N_19902,N_16996,N_18654);
or U19903 (N_19903,N_18234,N_16690);
xor U19904 (N_19904,N_17175,N_17448);
nor U19905 (N_19905,N_16769,N_17802);
nand U19906 (N_19906,N_17274,N_18408);
nand U19907 (N_19907,N_17346,N_16802);
xnor U19908 (N_19908,N_15690,N_18169);
nand U19909 (N_19909,N_16231,N_15894);
nor U19910 (N_19910,N_16311,N_18384);
and U19911 (N_19911,N_17241,N_15656);
and U19912 (N_19912,N_15818,N_18296);
xor U19913 (N_19913,N_18036,N_16415);
nand U19914 (N_19914,N_15845,N_17372);
nor U19915 (N_19915,N_16902,N_18404);
and U19916 (N_19916,N_18020,N_18209);
nand U19917 (N_19917,N_18359,N_16528);
and U19918 (N_19918,N_17756,N_16519);
or U19919 (N_19919,N_18501,N_17391);
nand U19920 (N_19920,N_17393,N_17835);
nor U19921 (N_19921,N_18164,N_15887);
nor U19922 (N_19922,N_17213,N_17369);
or U19923 (N_19923,N_16754,N_17221);
nor U19924 (N_19924,N_18691,N_17389);
nand U19925 (N_19925,N_17766,N_16603);
nor U19926 (N_19926,N_18405,N_18364);
nor U19927 (N_19927,N_16660,N_17833);
or U19928 (N_19928,N_17973,N_15837);
or U19929 (N_19929,N_18406,N_16477);
and U19930 (N_19930,N_18215,N_16315);
or U19931 (N_19931,N_18214,N_16211);
nor U19932 (N_19932,N_17031,N_18108);
xnor U19933 (N_19933,N_17969,N_16147);
or U19934 (N_19934,N_16501,N_16365);
nand U19935 (N_19935,N_15803,N_18037);
nor U19936 (N_19936,N_18066,N_17919);
xnor U19937 (N_19937,N_17928,N_17214);
nor U19938 (N_19938,N_15935,N_16347);
xnor U19939 (N_19939,N_16108,N_15774);
nor U19940 (N_19940,N_17380,N_18288);
xor U19941 (N_19941,N_18487,N_17497);
xor U19942 (N_19942,N_17430,N_18155);
and U19943 (N_19943,N_18470,N_15858);
nor U19944 (N_19944,N_18123,N_18386);
and U19945 (N_19945,N_16360,N_17740);
nand U19946 (N_19946,N_16925,N_18623);
and U19947 (N_19947,N_17911,N_17857);
nand U19948 (N_19948,N_17819,N_17746);
and U19949 (N_19949,N_17769,N_18257);
nand U19950 (N_19950,N_18054,N_17978);
or U19951 (N_19951,N_16378,N_15856);
xor U19952 (N_19952,N_17779,N_17255);
and U19953 (N_19953,N_16814,N_16292);
and U19954 (N_19954,N_15982,N_17358);
nor U19955 (N_19955,N_18139,N_16747);
and U19956 (N_19956,N_16490,N_17854);
and U19957 (N_19957,N_17004,N_17270);
xor U19958 (N_19958,N_16800,N_18255);
nor U19959 (N_19959,N_18604,N_18668);
nand U19960 (N_19960,N_15987,N_17421);
nor U19961 (N_19961,N_18554,N_18539);
nor U19962 (N_19962,N_16134,N_17133);
or U19963 (N_19963,N_15751,N_16847);
and U19964 (N_19964,N_16588,N_17764);
nand U19965 (N_19965,N_15847,N_17332);
and U19966 (N_19966,N_16990,N_16088);
xnor U19967 (N_19967,N_15725,N_18547);
and U19968 (N_19968,N_18084,N_17354);
nand U19969 (N_19969,N_15745,N_17890);
and U19970 (N_19970,N_18128,N_18599);
nand U19971 (N_19971,N_15908,N_16685);
or U19972 (N_19972,N_16331,N_17429);
nand U19973 (N_19973,N_17171,N_17153);
nor U19974 (N_19974,N_17686,N_17840);
nor U19975 (N_19975,N_16511,N_17991);
or U19976 (N_19976,N_18220,N_17259);
xor U19977 (N_19977,N_18216,N_17117);
nand U19978 (N_19978,N_18352,N_18118);
nand U19979 (N_19979,N_16187,N_16268);
and U19980 (N_19980,N_18058,N_16638);
nor U19981 (N_19981,N_16809,N_15841);
xnor U19982 (N_19982,N_16351,N_16828);
xor U19983 (N_19983,N_17418,N_17013);
and U19984 (N_19984,N_17417,N_18504);
xor U19985 (N_19985,N_18152,N_18448);
nor U19986 (N_19986,N_17375,N_18282);
or U19987 (N_19987,N_18211,N_15727);
nor U19988 (N_19988,N_18596,N_15983);
and U19989 (N_19989,N_18113,N_16811);
xnor U19990 (N_19990,N_16163,N_16462);
nand U19991 (N_19991,N_17486,N_15833);
and U19992 (N_19992,N_17123,N_16458);
nand U19993 (N_19993,N_18389,N_18268);
xnor U19994 (N_19994,N_17897,N_17760);
and U19995 (N_19995,N_17239,N_15874);
and U19996 (N_19996,N_16265,N_18239);
or U19997 (N_19997,N_16269,N_18284);
xor U19998 (N_19998,N_16476,N_16530);
or U19999 (N_19999,N_17075,N_17132);
nand U20000 (N_20000,N_18272,N_17957);
nand U20001 (N_20001,N_18258,N_17303);
and U20002 (N_20002,N_18150,N_16905);
or U20003 (N_20003,N_16726,N_16045);
nor U20004 (N_20004,N_16651,N_16343);
nand U20005 (N_20005,N_17381,N_18226);
or U20006 (N_20006,N_17219,N_15696);
or U20007 (N_20007,N_17946,N_17575);
or U20008 (N_20008,N_17670,N_15998);
xnor U20009 (N_20009,N_17326,N_17420);
xnor U20010 (N_20010,N_17970,N_16348);
nor U20011 (N_20011,N_16955,N_18532);
nor U20012 (N_20012,N_18517,N_16866);
xnor U20013 (N_20013,N_18061,N_16923);
nor U20014 (N_20014,N_17684,N_17932);
nor U20015 (N_20015,N_15980,N_15649);
nor U20016 (N_20016,N_17313,N_16392);
and U20017 (N_20017,N_18279,N_17322);
or U20018 (N_20018,N_15788,N_16875);
xnor U20019 (N_20019,N_16457,N_15912);
nand U20020 (N_20020,N_15647,N_18615);
nand U20021 (N_20021,N_18721,N_16276);
or U20022 (N_20022,N_17881,N_17356);
nor U20023 (N_20023,N_15761,N_15791);
and U20024 (N_20024,N_16946,N_16721);
or U20025 (N_20025,N_16916,N_16445);
and U20026 (N_20026,N_16238,N_17271);
or U20027 (N_20027,N_15909,N_16059);
nor U20028 (N_20028,N_16592,N_17489);
and U20029 (N_20029,N_15890,N_16583);
nor U20030 (N_20030,N_17488,N_17540);
nor U20031 (N_20031,N_18270,N_17415);
nor U20032 (N_20032,N_16450,N_18420);
and U20033 (N_20033,N_16680,N_17183);
xnor U20034 (N_20034,N_16066,N_16799);
nand U20035 (N_20035,N_17923,N_18521);
or U20036 (N_20036,N_16877,N_18712);
nor U20037 (N_20037,N_18564,N_16621);
nand U20038 (N_20038,N_15692,N_16554);
or U20039 (N_20039,N_17850,N_15931);
xor U20040 (N_20040,N_16698,N_18038);
or U20041 (N_20041,N_18495,N_18347);
nand U20042 (N_20042,N_18567,N_16699);
xnor U20043 (N_20043,N_18085,N_18651);
nand U20044 (N_20044,N_17513,N_16489);
xnor U20045 (N_20045,N_16840,N_15968);
and U20046 (N_20046,N_17193,N_17139);
nand U20047 (N_20047,N_16260,N_17124);
or U20048 (N_20048,N_16740,N_16738);
xor U20049 (N_20049,N_16150,N_18613);
nor U20050 (N_20050,N_16345,N_16005);
and U20051 (N_20051,N_18601,N_17349);
nand U20052 (N_20052,N_17730,N_18402);
xnor U20053 (N_20053,N_17205,N_18580);
xor U20054 (N_20054,N_17515,N_17847);
nor U20055 (N_20055,N_17079,N_16003);
nor U20056 (N_20056,N_16332,N_18087);
nand U20057 (N_20057,N_17341,N_18286);
or U20058 (N_20058,N_16013,N_17238);
and U20059 (N_20059,N_16007,N_17316);
and U20060 (N_20060,N_17103,N_18122);
nor U20061 (N_20061,N_15703,N_16492);
nor U20062 (N_20062,N_15888,N_17275);
or U20063 (N_20063,N_17098,N_16521);
and U20064 (N_20064,N_15958,N_16030);
xor U20065 (N_20065,N_17592,N_17560);
and U20066 (N_20066,N_16999,N_16451);
or U20067 (N_20067,N_16795,N_17121);
xor U20068 (N_20068,N_18421,N_16283);
xnor U20069 (N_20069,N_16676,N_18097);
and U20070 (N_20070,N_17635,N_16162);
or U20071 (N_20071,N_15644,N_17359);
or U20072 (N_20072,N_16922,N_17623);
nand U20073 (N_20073,N_18275,N_18709);
nor U20074 (N_20074,N_18559,N_16507);
or U20075 (N_20075,N_18525,N_15905);
nand U20076 (N_20076,N_18142,N_16046);
xor U20077 (N_20077,N_18339,N_16565);
nand U20078 (N_20078,N_16850,N_17920);
xor U20079 (N_20079,N_15697,N_15768);
nand U20080 (N_20080,N_18146,N_17434);
xor U20081 (N_20081,N_18248,N_18725);
xnor U20082 (N_20082,N_17680,N_18719);
or U20083 (N_20083,N_17913,N_15849);
nand U20084 (N_20084,N_16200,N_17535);
and U20085 (N_20085,N_17867,N_18329);
nor U20086 (N_20086,N_16316,N_17530);
or U20087 (N_20087,N_15652,N_16700);
xor U20088 (N_20088,N_16427,N_16470);
nand U20089 (N_20089,N_17813,N_17006);
or U20090 (N_20090,N_17892,N_17445);
xor U20091 (N_20091,N_18546,N_18067);
nor U20092 (N_20092,N_17056,N_17719);
or U20093 (N_20093,N_15667,N_17805);
nor U20094 (N_20094,N_16779,N_15883);
xor U20095 (N_20095,N_17083,N_17046);
xnor U20096 (N_20096,N_17674,N_17176);
or U20097 (N_20097,N_18579,N_18345);
xnor U20098 (N_20098,N_16677,N_18100);
nor U20099 (N_20099,N_16272,N_18022);
nor U20100 (N_20100,N_17845,N_17099);
nor U20101 (N_20101,N_15742,N_16919);
xor U20102 (N_20102,N_18095,N_17450);
nor U20103 (N_20103,N_17567,N_16127);
nand U20104 (N_20104,N_17197,N_16170);
nor U20105 (N_20105,N_18636,N_17093);
and U20106 (N_20106,N_16524,N_16145);
or U20107 (N_20107,N_16550,N_18136);
or U20108 (N_20108,N_16630,N_17007);
xnor U20109 (N_20109,N_17485,N_18233);
nand U20110 (N_20110,N_15764,N_16958);
nand U20111 (N_20111,N_16198,N_18733);
and U20112 (N_20112,N_15996,N_16752);
nand U20113 (N_20113,N_17925,N_17229);
and U20114 (N_20114,N_18188,N_18442);
or U20115 (N_20115,N_15759,N_17975);
nand U20116 (N_20116,N_16050,N_17997);
nor U20117 (N_20117,N_17559,N_17695);
xnor U20118 (N_20118,N_15992,N_17471);
and U20119 (N_20119,N_17960,N_17884);
nor U20120 (N_20120,N_18192,N_18180);
or U20121 (N_20121,N_16715,N_17542);
xor U20122 (N_20122,N_16473,N_16897);
and U20123 (N_20123,N_16379,N_17720);
xor U20124 (N_20124,N_17616,N_16873);
and U20125 (N_20125,N_17258,N_17232);
or U20126 (N_20126,N_17101,N_18222);
xor U20127 (N_20127,N_16907,N_16707);
xnor U20128 (N_20128,N_18679,N_18145);
or U20129 (N_20129,N_17404,N_15926);
nor U20130 (N_20130,N_16616,N_16974);
or U20131 (N_20131,N_16178,N_18354);
nand U20132 (N_20132,N_18457,N_17426);
nand U20133 (N_20133,N_16034,N_15990);
xor U20134 (N_20134,N_16080,N_16580);
xor U20135 (N_20135,N_18660,N_16969);
or U20136 (N_20136,N_16959,N_16223);
xnor U20137 (N_20137,N_17474,N_17681);
and U20138 (N_20138,N_16449,N_18609);
xnor U20139 (N_20139,N_16107,N_16794);
or U20140 (N_20140,N_17438,N_16418);
xor U20141 (N_20141,N_17447,N_18588);
nand U20142 (N_20142,N_16233,N_17043);
nor U20143 (N_20143,N_16104,N_17568);
nand U20144 (N_20144,N_18610,N_17558);
nand U20145 (N_20145,N_15901,N_18687);
nand U20146 (N_20146,N_18531,N_16842);
nor U20147 (N_20147,N_15986,N_16131);
nor U20148 (N_20148,N_17409,N_17050);
xnor U20149 (N_20149,N_17888,N_18294);
nand U20150 (N_20150,N_17510,N_15752);
xor U20151 (N_20151,N_18677,N_17905);
nand U20152 (N_20152,N_17808,N_17399);
nand U20153 (N_20153,N_17522,N_17521);
xor U20154 (N_20154,N_16289,N_16092);
and U20155 (N_20155,N_18598,N_17873);
xor U20156 (N_20156,N_17739,N_16662);
or U20157 (N_20157,N_17390,N_17554);
nor U20158 (N_20158,N_15817,N_18235);
nand U20159 (N_20159,N_16841,N_16245);
nand U20160 (N_20160,N_16525,N_15957);
and U20161 (N_20161,N_17986,N_17908);
xnor U20162 (N_20162,N_17812,N_16133);
xor U20163 (N_20163,N_17662,N_17398);
and U20164 (N_20164,N_17100,N_17267);
nor U20165 (N_20165,N_16672,N_17155);
and U20166 (N_20166,N_17660,N_18560);
xnor U20167 (N_20167,N_18416,N_15916);
and U20168 (N_20168,N_16522,N_17457);
and U20169 (N_20169,N_18621,N_16082);
nand U20170 (N_20170,N_16308,N_17852);
or U20171 (N_20171,N_17003,N_18541);
nand U20172 (N_20172,N_16557,N_17774);
xnor U20173 (N_20173,N_17569,N_15789);
nor U20174 (N_20174,N_18028,N_16956);
xnor U20175 (N_20175,N_17846,N_17749);
or U20176 (N_20176,N_17048,N_16103);
or U20177 (N_20177,N_17295,N_17422);
nand U20178 (N_20178,N_16199,N_16460);
nor U20179 (N_20179,N_17112,N_15806);
and U20180 (N_20180,N_17601,N_15748);
and U20181 (N_20181,N_15773,N_16031);
nand U20182 (N_20182,N_18548,N_16735);
nor U20183 (N_20183,N_16335,N_18140);
or U20184 (N_20184,N_18033,N_18520);
nand U20185 (N_20185,N_17977,N_17455);
or U20186 (N_20186,N_15709,N_15960);
nand U20187 (N_20187,N_17992,N_15823);
and U20188 (N_20188,N_16815,N_18002);
nor U20189 (N_20189,N_17907,N_15678);
nand U20190 (N_20190,N_16497,N_16135);
nor U20191 (N_20191,N_16675,N_16590);
or U20192 (N_20192,N_15701,N_18722);
or U20193 (N_20193,N_17283,N_17094);
nor U20194 (N_20194,N_18285,N_18593);
nor U20195 (N_20195,N_18577,N_18326);
or U20196 (N_20196,N_17315,N_18624);
or U20197 (N_20197,N_16298,N_15673);
nor U20198 (N_20198,N_16684,N_16686);
xnor U20199 (N_20199,N_16646,N_16538);
and U20200 (N_20200,N_17125,N_16075);
xnor U20201 (N_20201,N_16784,N_16578);
nand U20202 (N_20202,N_17809,N_18060);
nand U20203 (N_20203,N_15766,N_16466);
and U20204 (N_20204,N_16644,N_18595);
and U20205 (N_20205,N_18650,N_17384);
and U20206 (N_20206,N_16142,N_18236);
or U20207 (N_20207,N_17266,N_16775);
and U20208 (N_20208,N_17036,N_16601);
xor U20209 (N_20209,N_18099,N_18696);
nand U20210 (N_20210,N_18090,N_17627);
nor U20211 (N_20211,N_18010,N_16324);
nand U20212 (N_20212,N_18441,N_16975);
xnor U20213 (N_20213,N_18489,N_16629);
nand U20214 (N_20214,N_17364,N_17658);
nor U20215 (N_20215,N_17866,N_16941);
xnor U20216 (N_20216,N_18250,N_16148);
nor U20217 (N_20217,N_17441,N_17743);
xor U20218 (N_20218,N_16032,N_17279);
and U20219 (N_20219,N_18178,N_18607);
nor U20220 (N_20220,N_16190,N_16074);
nor U20221 (N_20221,N_18553,N_16920);
and U20222 (N_20222,N_16982,N_16984);
nor U20223 (N_20223,N_18273,N_17156);
nor U20224 (N_20224,N_18466,N_18731);
nor U20225 (N_20225,N_18715,N_17397);
nor U20226 (N_20226,N_15896,N_18515);
and U20227 (N_20227,N_18071,N_17527);
or U20228 (N_20228,N_15790,N_16158);
or U20229 (N_20229,N_17337,N_16112);
or U20230 (N_20230,N_16290,N_17646);
nand U20231 (N_20231,N_16861,N_15660);
xnor U20232 (N_20232,N_18313,N_18137);
xnor U20233 (N_20233,N_16029,N_17208);
xor U20234 (N_20234,N_18310,N_16512);
nand U20235 (N_20235,N_16105,N_17863);
nand U20236 (N_20236,N_16615,N_18700);
or U20237 (N_20237,N_15904,N_16838);
and U20238 (N_20238,N_17901,N_17511);
and U20239 (N_20239,N_18675,N_17732);
nand U20240 (N_20240,N_16452,N_17253);
or U20241 (N_20241,N_16207,N_16682);
and U20242 (N_20242,N_16049,N_16383);
nand U20243 (N_20243,N_16702,N_18738);
xor U20244 (N_20244,N_17030,N_17490);
and U20245 (N_20245,N_15923,N_16405);
nor U20246 (N_20246,N_16078,N_17163);
xor U20247 (N_20247,N_16812,N_18600);
xor U20248 (N_20248,N_17301,N_16194);
nand U20249 (N_20249,N_17842,N_18241);
nor U20250 (N_20250,N_18706,N_18198);
and U20251 (N_20251,N_18088,N_17596);
nor U20252 (N_20252,N_18340,N_16299);
or U20253 (N_20253,N_16962,N_18659);
and U20254 (N_20254,N_15780,N_17242);
or U20255 (N_20255,N_17136,N_17215);
and U20256 (N_20256,N_17307,N_17787);
or U20257 (N_20257,N_15863,N_15737);
xnor U20258 (N_20258,N_16886,N_17640);
nand U20259 (N_20259,N_16478,N_16468);
and U20260 (N_20260,N_17465,N_16284);
and U20261 (N_20261,N_16300,N_18322);
and U20262 (N_20262,N_16022,N_16213);
and U20263 (N_20263,N_17257,N_18681);
xor U20264 (N_20264,N_18629,N_16759);
nor U20265 (N_20265,N_16015,N_18376);
and U20266 (N_20266,N_17935,N_15636);
or U20267 (N_20267,N_15870,N_18230);
or U20268 (N_20268,N_16865,N_17116);
and U20269 (N_20269,N_18536,N_18423);
xor U20270 (N_20270,N_16942,N_18471);
or U20271 (N_20271,N_17605,N_15639);
nand U20272 (N_20272,N_18314,N_17454);
and U20273 (N_20273,N_17137,N_17164);
nor U20274 (N_20274,N_17676,N_17202);
or U20275 (N_20275,N_16055,N_16856);
nor U20276 (N_20276,N_16277,N_16438);
nor U20277 (N_20277,N_17898,N_16636);
nor U20278 (N_20278,N_16423,N_16966);
or U20279 (N_20279,N_16173,N_18480);
nor U20280 (N_20280,N_16619,N_15746);
nand U20281 (N_20281,N_17688,N_16381);
or U20282 (N_20282,N_17636,N_18117);
xnor U20283 (N_20283,N_18256,N_16547);
xor U20284 (N_20284,N_16141,N_18324);
nand U20285 (N_20285,N_17284,N_15824);
and U20286 (N_20286,N_18302,N_18221);
and U20287 (N_20287,N_18008,N_18611);
nand U20288 (N_20288,N_16723,N_17758);
and U20289 (N_20289,N_17444,N_15838);
and U20290 (N_20290,N_17029,N_18074);
and U20291 (N_20291,N_18165,N_17032);
or U20292 (N_20292,N_18669,N_15954);
and U20293 (N_20293,N_18325,N_18172);
xor U20294 (N_20294,N_18602,N_18168);
or U20295 (N_20295,N_18555,N_17343);
nand U20296 (N_20296,N_15820,N_16930);
nor U20297 (N_20297,N_17405,N_16874);
xnor U20298 (N_20298,N_15937,N_17247);
nand U20299 (N_20299,N_15799,N_17355);
or U20300 (N_20300,N_16221,N_16099);
xor U20301 (N_20301,N_17318,N_17822);
nor U20302 (N_20302,N_17165,N_18186);
nor U20303 (N_20303,N_16407,N_18069);
nand U20304 (N_20304,N_17272,N_18048);
nor U20305 (N_20305,N_18622,N_18103);
xor U20306 (N_20306,N_16291,N_16023);
and U20307 (N_20307,N_16527,N_17529);
and U20308 (N_20308,N_17160,N_17237);
or U20309 (N_20309,N_17848,N_17293);
nor U20310 (N_20310,N_15860,N_18581);
nand U20311 (N_20311,N_18538,N_16634);
nor U20312 (N_20312,N_16267,N_18732);
nand U20313 (N_20313,N_16357,N_15748);
nor U20314 (N_20314,N_17333,N_16899);
nand U20315 (N_20315,N_16820,N_17835);
and U20316 (N_20316,N_17158,N_18262);
nor U20317 (N_20317,N_18296,N_16196);
and U20318 (N_20318,N_16526,N_17067);
and U20319 (N_20319,N_16103,N_15811);
nor U20320 (N_20320,N_17394,N_17159);
and U20321 (N_20321,N_17652,N_16213);
or U20322 (N_20322,N_17665,N_17966);
nand U20323 (N_20323,N_16122,N_16593);
nor U20324 (N_20324,N_15991,N_16306);
nor U20325 (N_20325,N_18357,N_17807);
xnor U20326 (N_20326,N_18092,N_18729);
or U20327 (N_20327,N_18160,N_16294);
nand U20328 (N_20328,N_15958,N_16739);
or U20329 (N_20329,N_16319,N_17344);
xnor U20330 (N_20330,N_18207,N_17782);
or U20331 (N_20331,N_18417,N_17852);
xnor U20332 (N_20332,N_16071,N_17069);
nand U20333 (N_20333,N_17326,N_17250);
xnor U20334 (N_20334,N_18156,N_17046);
and U20335 (N_20335,N_17281,N_16869);
nor U20336 (N_20336,N_16863,N_17586);
nor U20337 (N_20337,N_18062,N_17068);
nand U20338 (N_20338,N_17629,N_17943);
xor U20339 (N_20339,N_15839,N_16479);
nor U20340 (N_20340,N_17432,N_18711);
and U20341 (N_20341,N_15891,N_17910);
or U20342 (N_20342,N_17598,N_17916);
or U20343 (N_20343,N_18636,N_18185);
or U20344 (N_20344,N_17176,N_17252);
and U20345 (N_20345,N_16775,N_17114);
nor U20346 (N_20346,N_16518,N_16529);
nor U20347 (N_20347,N_17154,N_16423);
or U20348 (N_20348,N_16138,N_16803);
nand U20349 (N_20349,N_15874,N_17864);
or U20350 (N_20350,N_17445,N_18158);
or U20351 (N_20351,N_16579,N_16074);
and U20352 (N_20352,N_16658,N_18396);
nand U20353 (N_20353,N_16607,N_16691);
xnor U20354 (N_20354,N_17746,N_16446);
nor U20355 (N_20355,N_17784,N_17805);
xnor U20356 (N_20356,N_16072,N_16974);
and U20357 (N_20357,N_16031,N_18463);
xnor U20358 (N_20358,N_15936,N_16592);
nand U20359 (N_20359,N_15669,N_16974);
and U20360 (N_20360,N_16279,N_16004);
xor U20361 (N_20361,N_16622,N_16634);
or U20362 (N_20362,N_18451,N_17856);
nand U20363 (N_20363,N_15938,N_15949);
or U20364 (N_20364,N_18171,N_16465);
or U20365 (N_20365,N_16157,N_15813);
nand U20366 (N_20366,N_18017,N_18498);
and U20367 (N_20367,N_17127,N_18209);
nor U20368 (N_20368,N_17652,N_16882);
and U20369 (N_20369,N_17459,N_16584);
and U20370 (N_20370,N_17103,N_18079);
nor U20371 (N_20371,N_16740,N_16858);
nor U20372 (N_20372,N_16271,N_16336);
xor U20373 (N_20373,N_18568,N_18505);
and U20374 (N_20374,N_16844,N_18442);
and U20375 (N_20375,N_17267,N_17563);
or U20376 (N_20376,N_15911,N_17331);
nand U20377 (N_20377,N_18137,N_17006);
nand U20378 (N_20378,N_16909,N_17811);
xnor U20379 (N_20379,N_16128,N_17475);
xor U20380 (N_20380,N_18317,N_18177);
nand U20381 (N_20381,N_17777,N_18556);
nand U20382 (N_20382,N_18340,N_18367);
or U20383 (N_20383,N_18359,N_15861);
nand U20384 (N_20384,N_18675,N_16173);
and U20385 (N_20385,N_16281,N_16491);
nand U20386 (N_20386,N_15883,N_18275);
xnor U20387 (N_20387,N_16840,N_18112);
and U20388 (N_20388,N_17343,N_16861);
nor U20389 (N_20389,N_15638,N_17260);
xnor U20390 (N_20390,N_16885,N_17501);
and U20391 (N_20391,N_18547,N_18696);
nand U20392 (N_20392,N_16144,N_17502);
xnor U20393 (N_20393,N_16190,N_18090);
nand U20394 (N_20394,N_17848,N_18160);
xnor U20395 (N_20395,N_18553,N_18627);
nor U20396 (N_20396,N_17212,N_18741);
nand U20397 (N_20397,N_16612,N_17323);
or U20398 (N_20398,N_17986,N_18706);
or U20399 (N_20399,N_17129,N_15630);
nand U20400 (N_20400,N_18744,N_18414);
or U20401 (N_20401,N_18015,N_17401);
xnor U20402 (N_20402,N_16751,N_18140);
xnor U20403 (N_20403,N_15793,N_18094);
xnor U20404 (N_20404,N_17561,N_17958);
nand U20405 (N_20405,N_18575,N_17515);
xor U20406 (N_20406,N_17218,N_16575);
nor U20407 (N_20407,N_16440,N_15897);
nand U20408 (N_20408,N_16006,N_17711);
and U20409 (N_20409,N_18634,N_17128);
or U20410 (N_20410,N_16814,N_17910);
or U20411 (N_20411,N_17108,N_18486);
xnor U20412 (N_20412,N_17734,N_17468);
nand U20413 (N_20413,N_16277,N_16287);
xor U20414 (N_20414,N_15834,N_17257);
xor U20415 (N_20415,N_15893,N_17412);
nor U20416 (N_20416,N_17653,N_16317);
or U20417 (N_20417,N_16232,N_16939);
nand U20418 (N_20418,N_18532,N_17255);
and U20419 (N_20419,N_16957,N_16386);
xor U20420 (N_20420,N_18579,N_17805);
or U20421 (N_20421,N_17293,N_17433);
nor U20422 (N_20422,N_17108,N_15730);
nand U20423 (N_20423,N_17852,N_17791);
or U20424 (N_20424,N_16379,N_17817);
xnor U20425 (N_20425,N_17879,N_15956);
xor U20426 (N_20426,N_18565,N_16930);
nand U20427 (N_20427,N_17487,N_17397);
nor U20428 (N_20428,N_17280,N_17858);
nor U20429 (N_20429,N_16451,N_16113);
nand U20430 (N_20430,N_16522,N_17261);
or U20431 (N_20431,N_15683,N_16926);
nand U20432 (N_20432,N_17161,N_16026);
nand U20433 (N_20433,N_16234,N_18596);
nor U20434 (N_20434,N_17342,N_15746);
nor U20435 (N_20435,N_18101,N_18742);
and U20436 (N_20436,N_17457,N_18531);
xnor U20437 (N_20437,N_18411,N_18040);
or U20438 (N_20438,N_16847,N_16561);
or U20439 (N_20439,N_16373,N_17065);
nor U20440 (N_20440,N_15818,N_15953);
and U20441 (N_20441,N_16237,N_15955);
nand U20442 (N_20442,N_16794,N_17538);
nand U20443 (N_20443,N_17650,N_16652);
nor U20444 (N_20444,N_16642,N_16788);
or U20445 (N_20445,N_18316,N_16671);
and U20446 (N_20446,N_15940,N_17691);
nor U20447 (N_20447,N_18486,N_17857);
nor U20448 (N_20448,N_17398,N_18311);
and U20449 (N_20449,N_16334,N_16188);
nand U20450 (N_20450,N_17429,N_16918);
and U20451 (N_20451,N_17722,N_17134);
nor U20452 (N_20452,N_17125,N_17183);
nor U20453 (N_20453,N_16006,N_18183);
nor U20454 (N_20454,N_18477,N_16025);
and U20455 (N_20455,N_18454,N_15840);
nand U20456 (N_20456,N_17456,N_15933);
nor U20457 (N_20457,N_18450,N_17056);
or U20458 (N_20458,N_15759,N_16448);
xnor U20459 (N_20459,N_16355,N_18365);
nor U20460 (N_20460,N_16423,N_16707);
nor U20461 (N_20461,N_17690,N_15961);
nand U20462 (N_20462,N_17850,N_16276);
nand U20463 (N_20463,N_18563,N_16641);
nand U20464 (N_20464,N_17252,N_16067);
nor U20465 (N_20465,N_17505,N_18299);
or U20466 (N_20466,N_17767,N_16678);
nand U20467 (N_20467,N_17579,N_16022);
xnor U20468 (N_20468,N_15625,N_18355);
nand U20469 (N_20469,N_16707,N_16823);
and U20470 (N_20470,N_18274,N_18179);
and U20471 (N_20471,N_17706,N_17100);
xnor U20472 (N_20472,N_16237,N_17641);
xnor U20473 (N_20473,N_16176,N_17660);
xnor U20474 (N_20474,N_17842,N_16621);
or U20475 (N_20475,N_17114,N_17185);
and U20476 (N_20476,N_17175,N_16953);
nor U20477 (N_20477,N_16794,N_17842);
nand U20478 (N_20478,N_18135,N_17319);
nand U20479 (N_20479,N_18271,N_17570);
and U20480 (N_20480,N_18126,N_18700);
nor U20481 (N_20481,N_15848,N_16650);
and U20482 (N_20482,N_17816,N_16251);
and U20483 (N_20483,N_16709,N_17988);
and U20484 (N_20484,N_18334,N_16924);
and U20485 (N_20485,N_16050,N_17191);
and U20486 (N_20486,N_16233,N_16387);
and U20487 (N_20487,N_16055,N_18005);
nor U20488 (N_20488,N_16660,N_18055);
or U20489 (N_20489,N_17475,N_15816);
and U20490 (N_20490,N_17064,N_17896);
xor U20491 (N_20491,N_16185,N_17005);
or U20492 (N_20492,N_18454,N_15843);
nor U20493 (N_20493,N_16776,N_16619);
or U20494 (N_20494,N_17512,N_16207);
nor U20495 (N_20495,N_18538,N_16236);
nand U20496 (N_20496,N_16488,N_17554);
or U20497 (N_20497,N_16057,N_16303);
or U20498 (N_20498,N_16865,N_16161);
nor U20499 (N_20499,N_18009,N_17267);
xnor U20500 (N_20500,N_15895,N_16426);
nor U20501 (N_20501,N_18400,N_17247);
xor U20502 (N_20502,N_15840,N_15867);
nor U20503 (N_20503,N_17036,N_16529);
xnor U20504 (N_20504,N_16752,N_15884);
nand U20505 (N_20505,N_18669,N_16221);
nand U20506 (N_20506,N_18399,N_17947);
or U20507 (N_20507,N_15788,N_18259);
xnor U20508 (N_20508,N_16219,N_16800);
and U20509 (N_20509,N_15769,N_15951);
or U20510 (N_20510,N_16871,N_16331);
nand U20511 (N_20511,N_17365,N_18583);
xnor U20512 (N_20512,N_17124,N_16194);
and U20513 (N_20513,N_17606,N_16632);
xor U20514 (N_20514,N_16166,N_16820);
xor U20515 (N_20515,N_16340,N_17528);
nand U20516 (N_20516,N_18685,N_18016);
and U20517 (N_20517,N_17608,N_18096);
or U20518 (N_20518,N_17203,N_15978);
nand U20519 (N_20519,N_18293,N_15696);
or U20520 (N_20520,N_16374,N_15933);
nand U20521 (N_20521,N_18077,N_16891);
nand U20522 (N_20522,N_17683,N_16667);
nor U20523 (N_20523,N_16134,N_18399);
and U20524 (N_20524,N_18171,N_17901);
xnor U20525 (N_20525,N_18654,N_17541);
or U20526 (N_20526,N_16220,N_17549);
or U20527 (N_20527,N_18521,N_16985);
or U20528 (N_20528,N_16674,N_16261);
nand U20529 (N_20529,N_18497,N_16438);
xor U20530 (N_20530,N_18557,N_18165);
and U20531 (N_20531,N_17181,N_15813);
or U20532 (N_20532,N_15879,N_18471);
nor U20533 (N_20533,N_16348,N_18518);
xor U20534 (N_20534,N_16234,N_18208);
nand U20535 (N_20535,N_17822,N_18175);
or U20536 (N_20536,N_17765,N_16101);
nand U20537 (N_20537,N_17609,N_16414);
or U20538 (N_20538,N_17497,N_17160);
xor U20539 (N_20539,N_16869,N_18216);
xor U20540 (N_20540,N_18161,N_15864);
or U20541 (N_20541,N_17045,N_18451);
xor U20542 (N_20542,N_17540,N_18485);
and U20543 (N_20543,N_18390,N_17815);
xor U20544 (N_20544,N_18373,N_16003);
nor U20545 (N_20545,N_17082,N_18466);
nand U20546 (N_20546,N_16031,N_15880);
nor U20547 (N_20547,N_18092,N_17714);
nand U20548 (N_20548,N_15807,N_16692);
or U20549 (N_20549,N_16250,N_17971);
nand U20550 (N_20550,N_16905,N_17062);
xor U20551 (N_20551,N_16796,N_18469);
nor U20552 (N_20552,N_17244,N_16795);
nand U20553 (N_20553,N_17730,N_16471);
and U20554 (N_20554,N_16980,N_16528);
xnor U20555 (N_20555,N_17036,N_15696);
nand U20556 (N_20556,N_18041,N_16292);
nor U20557 (N_20557,N_16650,N_16506);
nand U20558 (N_20558,N_18398,N_17029);
and U20559 (N_20559,N_17931,N_15897);
and U20560 (N_20560,N_16714,N_17727);
xor U20561 (N_20561,N_16698,N_17833);
nor U20562 (N_20562,N_18001,N_16547);
and U20563 (N_20563,N_17335,N_18475);
xor U20564 (N_20564,N_17660,N_16837);
or U20565 (N_20565,N_15692,N_18418);
nor U20566 (N_20566,N_18661,N_18113);
and U20567 (N_20567,N_18458,N_16620);
and U20568 (N_20568,N_15988,N_16635);
nor U20569 (N_20569,N_18607,N_15966);
nand U20570 (N_20570,N_16843,N_18588);
xnor U20571 (N_20571,N_15938,N_17355);
nor U20572 (N_20572,N_16073,N_18498);
nand U20573 (N_20573,N_17564,N_17487);
nand U20574 (N_20574,N_16879,N_17554);
nor U20575 (N_20575,N_17929,N_17278);
and U20576 (N_20576,N_15883,N_16854);
or U20577 (N_20577,N_17951,N_17685);
nand U20578 (N_20578,N_17635,N_18747);
nor U20579 (N_20579,N_18222,N_15833);
nor U20580 (N_20580,N_17200,N_18693);
nand U20581 (N_20581,N_17929,N_18504);
nand U20582 (N_20582,N_18168,N_18603);
and U20583 (N_20583,N_16819,N_18675);
or U20584 (N_20584,N_16304,N_15868);
nor U20585 (N_20585,N_17142,N_18047);
nor U20586 (N_20586,N_15794,N_17532);
or U20587 (N_20587,N_16366,N_17908);
nand U20588 (N_20588,N_17154,N_16966);
or U20589 (N_20589,N_17789,N_15886);
and U20590 (N_20590,N_17458,N_18502);
xor U20591 (N_20591,N_18173,N_16157);
and U20592 (N_20592,N_18686,N_15991);
nor U20593 (N_20593,N_16155,N_17637);
nand U20594 (N_20594,N_16348,N_16234);
nor U20595 (N_20595,N_16138,N_17764);
nand U20596 (N_20596,N_17202,N_15636);
and U20597 (N_20597,N_18358,N_17625);
xor U20598 (N_20598,N_18307,N_16874);
xnor U20599 (N_20599,N_15870,N_16195);
nand U20600 (N_20600,N_17150,N_16191);
or U20601 (N_20601,N_18069,N_17028);
nand U20602 (N_20602,N_17295,N_15901);
or U20603 (N_20603,N_17587,N_15986);
nand U20604 (N_20604,N_16225,N_16128);
or U20605 (N_20605,N_17850,N_18351);
xor U20606 (N_20606,N_16481,N_17691);
xor U20607 (N_20607,N_15891,N_17558);
nand U20608 (N_20608,N_17483,N_17292);
and U20609 (N_20609,N_16347,N_16099);
xor U20610 (N_20610,N_17836,N_17204);
nand U20611 (N_20611,N_18187,N_18478);
and U20612 (N_20612,N_17116,N_16274);
xor U20613 (N_20613,N_16984,N_17376);
nor U20614 (N_20614,N_15635,N_18603);
and U20615 (N_20615,N_17025,N_17288);
nor U20616 (N_20616,N_16689,N_15898);
and U20617 (N_20617,N_16200,N_17024);
and U20618 (N_20618,N_16947,N_17300);
or U20619 (N_20619,N_18718,N_17262);
xor U20620 (N_20620,N_16355,N_16818);
or U20621 (N_20621,N_16034,N_16420);
nand U20622 (N_20622,N_18637,N_18488);
nand U20623 (N_20623,N_16421,N_18494);
xor U20624 (N_20624,N_17373,N_18628);
or U20625 (N_20625,N_15911,N_15632);
nand U20626 (N_20626,N_17752,N_16289);
nor U20627 (N_20627,N_18380,N_17874);
nor U20628 (N_20628,N_18075,N_17314);
or U20629 (N_20629,N_18295,N_16730);
or U20630 (N_20630,N_16369,N_15632);
nor U20631 (N_20631,N_15680,N_17542);
xor U20632 (N_20632,N_18308,N_17957);
or U20633 (N_20633,N_16469,N_16095);
or U20634 (N_20634,N_18597,N_17595);
nor U20635 (N_20635,N_16650,N_16089);
or U20636 (N_20636,N_15670,N_17572);
and U20637 (N_20637,N_17927,N_18358);
and U20638 (N_20638,N_17751,N_17764);
and U20639 (N_20639,N_18314,N_15726);
xnor U20640 (N_20640,N_17634,N_17639);
xnor U20641 (N_20641,N_16957,N_18158);
nor U20642 (N_20642,N_18287,N_16656);
and U20643 (N_20643,N_15906,N_16387);
and U20644 (N_20644,N_17457,N_16649);
and U20645 (N_20645,N_16507,N_17023);
and U20646 (N_20646,N_17224,N_17491);
nand U20647 (N_20647,N_17424,N_17467);
nand U20648 (N_20648,N_17971,N_16443);
nand U20649 (N_20649,N_17996,N_17947);
nor U20650 (N_20650,N_16075,N_16872);
xnor U20651 (N_20651,N_17440,N_17841);
or U20652 (N_20652,N_16319,N_17142);
nand U20653 (N_20653,N_15968,N_18546);
or U20654 (N_20654,N_18643,N_15813);
or U20655 (N_20655,N_16143,N_17080);
xor U20656 (N_20656,N_18181,N_16778);
or U20657 (N_20657,N_17533,N_16821);
nor U20658 (N_20658,N_16471,N_17334);
nand U20659 (N_20659,N_18276,N_18192);
and U20660 (N_20660,N_16825,N_16473);
nor U20661 (N_20661,N_16262,N_17015);
and U20662 (N_20662,N_17433,N_16087);
and U20663 (N_20663,N_17870,N_18311);
and U20664 (N_20664,N_15941,N_16243);
xnor U20665 (N_20665,N_16802,N_18149);
nor U20666 (N_20666,N_16966,N_16990);
xnor U20667 (N_20667,N_16498,N_16623);
and U20668 (N_20668,N_18417,N_18655);
xor U20669 (N_20669,N_18690,N_17577);
nor U20670 (N_20670,N_18296,N_17023);
and U20671 (N_20671,N_18695,N_17895);
or U20672 (N_20672,N_16659,N_18276);
nor U20673 (N_20673,N_18686,N_17995);
xnor U20674 (N_20674,N_16906,N_16599);
nand U20675 (N_20675,N_18625,N_17252);
xor U20676 (N_20676,N_18524,N_16034);
or U20677 (N_20677,N_15776,N_17321);
xor U20678 (N_20678,N_18452,N_18321);
nor U20679 (N_20679,N_16247,N_16491);
xor U20680 (N_20680,N_16790,N_17664);
or U20681 (N_20681,N_17821,N_15876);
and U20682 (N_20682,N_18455,N_18719);
nand U20683 (N_20683,N_15815,N_17620);
nor U20684 (N_20684,N_16485,N_16427);
nor U20685 (N_20685,N_15907,N_15771);
nand U20686 (N_20686,N_17906,N_18437);
xor U20687 (N_20687,N_17773,N_17819);
xnor U20688 (N_20688,N_18285,N_16492);
or U20689 (N_20689,N_17948,N_16611);
or U20690 (N_20690,N_16853,N_17063);
and U20691 (N_20691,N_15774,N_15841);
nor U20692 (N_20692,N_16729,N_17133);
and U20693 (N_20693,N_17769,N_16527);
nor U20694 (N_20694,N_18541,N_17709);
nor U20695 (N_20695,N_17615,N_17363);
nand U20696 (N_20696,N_18528,N_16437);
or U20697 (N_20697,N_16061,N_17481);
nand U20698 (N_20698,N_18640,N_16672);
xor U20699 (N_20699,N_18168,N_16405);
nand U20700 (N_20700,N_17060,N_15747);
nor U20701 (N_20701,N_15768,N_16673);
xor U20702 (N_20702,N_16990,N_17827);
and U20703 (N_20703,N_17726,N_16217);
and U20704 (N_20704,N_16943,N_15857);
xnor U20705 (N_20705,N_18281,N_16238);
and U20706 (N_20706,N_18727,N_17114);
xor U20707 (N_20707,N_18182,N_17703);
and U20708 (N_20708,N_17367,N_17998);
or U20709 (N_20709,N_16220,N_16769);
or U20710 (N_20710,N_17872,N_16396);
xor U20711 (N_20711,N_15789,N_18186);
xnor U20712 (N_20712,N_17464,N_18446);
xnor U20713 (N_20713,N_16787,N_17598);
and U20714 (N_20714,N_16121,N_15666);
and U20715 (N_20715,N_17512,N_15907);
xnor U20716 (N_20716,N_17843,N_16162);
xnor U20717 (N_20717,N_16432,N_16595);
nor U20718 (N_20718,N_18287,N_16185);
or U20719 (N_20719,N_17425,N_18631);
nor U20720 (N_20720,N_15952,N_15974);
nor U20721 (N_20721,N_17631,N_16658);
and U20722 (N_20722,N_17309,N_17616);
or U20723 (N_20723,N_17159,N_17568);
and U20724 (N_20724,N_16470,N_16755);
nor U20725 (N_20725,N_16459,N_15694);
or U20726 (N_20726,N_17267,N_16096);
xor U20727 (N_20727,N_18459,N_18006);
or U20728 (N_20728,N_17952,N_18464);
nand U20729 (N_20729,N_17173,N_15630);
nor U20730 (N_20730,N_15672,N_17803);
nor U20731 (N_20731,N_17008,N_17490);
nand U20732 (N_20732,N_18033,N_17074);
and U20733 (N_20733,N_16653,N_18097);
xnor U20734 (N_20734,N_18559,N_16052);
nand U20735 (N_20735,N_16695,N_17709);
or U20736 (N_20736,N_16416,N_18014);
or U20737 (N_20737,N_17418,N_17679);
or U20738 (N_20738,N_16072,N_15864);
or U20739 (N_20739,N_16230,N_16746);
or U20740 (N_20740,N_17361,N_15747);
and U20741 (N_20741,N_15777,N_18037);
and U20742 (N_20742,N_17331,N_16219);
and U20743 (N_20743,N_17883,N_17230);
nor U20744 (N_20744,N_17184,N_18605);
and U20745 (N_20745,N_16871,N_18258);
nor U20746 (N_20746,N_17072,N_17615);
nor U20747 (N_20747,N_16675,N_15678);
or U20748 (N_20748,N_17943,N_16403);
and U20749 (N_20749,N_15754,N_17565);
nand U20750 (N_20750,N_18732,N_17084);
or U20751 (N_20751,N_16517,N_15915);
or U20752 (N_20752,N_16729,N_18694);
or U20753 (N_20753,N_16070,N_18029);
nor U20754 (N_20754,N_18281,N_16736);
nor U20755 (N_20755,N_16760,N_18507);
nand U20756 (N_20756,N_18547,N_17502);
nor U20757 (N_20757,N_18749,N_17386);
nand U20758 (N_20758,N_16195,N_18296);
and U20759 (N_20759,N_18012,N_18489);
nor U20760 (N_20760,N_16433,N_17023);
or U20761 (N_20761,N_17842,N_18679);
nor U20762 (N_20762,N_16643,N_16453);
and U20763 (N_20763,N_18301,N_16242);
nand U20764 (N_20764,N_16936,N_16358);
or U20765 (N_20765,N_18112,N_17336);
or U20766 (N_20766,N_17238,N_15963);
nor U20767 (N_20767,N_18173,N_16671);
or U20768 (N_20768,N_16768,N_17145);
or U20769 (N_20769,N_15806,N_17139);
xnor U20770 (N_20770,N_18437,N_18722);
nor U20771 (N_20771,N_16580,N_18074);
and U20772 (N_20772,N_17844,N_16541);
xnor U20773 (N_20773,N_17531,N_17341);
xnor U20774 (N_20774,N_15942,N_16887);
nand U20775 (N_20775,N_17881,N_15863);
nand U20776 (N_20776,N_18708,N_18721);
nand U20777 (N_20777,N_18307,N_16253);
and U20778 (N_20778,N_17559,N_17344);
xor U20779 (N_20779,N_15825,N_16737);
and U20780 (N_20780,N_18181,N_18213);
and U20781 (N_20781,N_17603,N_17899);
or U20782 (N_20782,N_15871,N_17962);
and U20783 (N_20783,N_18634,N_17751);
xnor U20784 (N_20784,N_17645,N_18745);
nand U20785 (N_20785,N_18007,N_17591);
xnor U20786 (N_20786,N_16043,N_18740);
xnor U20787 (N_20787,N_18037,N_16869);
xor U20788 (N_20788,N_18403,N_16918);
or U20789 (N_20789,N_16528,N_17065);
or U20790 (N_20790,N_15732,N_16811);
xor U20791 (N_20791,N_17268,N_15869);
nand U20792 (N_20792,N_16900,N_16100);
nor U20793 (N_20793,N_16020,N_18011);
and U20794 (N_20794,N_17842,N_16087);
xor U20795 (N_20795,N_17398,N_16284);
nand U20796 (N_20796,N_18461,N_16419);
nor U20797 (N_20797,N_18285,N_16398);
and U20798 (N_20798,N_18417,N_18249);
nand U20799 (N_20799,N_16301,N_17094);
nor U20800 (N_20800,N_17370,N_15710);
or U20801 (N_20801,N_15932,N_17001);
and U20802 (N_20802,N_18714,N_18523);
nor U20803 (N_20803,N_17147,N_18241);
nand U20804 (N_20804,N_16475,N_18349);
or U20805 (N_20805,N_16160,N_18587);
xnor U20806 (N_20806,N_17821,N_17612);
xor U20807 (N_20807,N_17158,N_16694);
nor U20808 (N_20808,N_16292,N_17920);
or U20809 (N_20809,N_17065,N_18478);
or U20810 (N_20810,N_17788,N_18096);
and U20811 (N_20811,N_17983,N_16353);
nor U20812 (N_20812,N_17809,N_18551);
nor U20813 (N_20813,N_16330,N_18000);
and U20814 (N_20814,N_17940,N_17318);
nor U20815 (N_20815,N_18694,N_16736);
nand U20816 (N_20816,N_17904,N_16923);
and U20817 (N_20817,N_16784,N_16351);
nand U20818 (N_20818,N_16192,N_16794);
and U20819 (N_20819,N_18115,N_17575);
nor U20820 (N_20820,N_17695,N_16853);
and U20821 (N_20821,N_18119,N_15676);
and U20822 (N_20822,N_17518,N_16326);
xnor U20823 (N_20823,N_16967,N_18218);
xor U20824 (N_20824,N_18560,N_17756);
and U20825 (N_20825,N_18244,N_16278);
or U20826 (N_20826,N_16522,N_16990);
xnor U20827 (N_20827,N_17872,N_16312);
or U20828 (N_20828,N_15719,N_16912);
or U20829 (N_20829,N_17937,N_17987);
nor U20830 (N_20830,N_16666,N_18178);
nand U20831 (N_20831,N_15998,N_17835);
and U20832 (N_20832,N_18296,N_16813);
nand U20833 (N_20833,N_15771,N_17301);
or U20834 (N_20834,N_15994,N_16867);
and U20835 (N_20835,N_17047,N_16949);
xnor U20836 (N_20836,N_17308,N_17675);
and U20837 (N_20837,N_18414,N_18582);
nor U20838 (N_20838,N_15737,N_17224);
and U20839 (N_20839,N_18485,N_17159);
nor U20840 (N_20840,N_17561,N_18478);
xor U20841 (N_20841,N_17756,N_18691);
xnor U20842 (N_20842,N_18185,N_15779);
and U20843 (N_20843,N_17078,N_15924);
and U20844 (N_20844,N_16014,N_17337);
nor U20845 (N_20845,N_18576,N_17874);
nand U20846 (N_20846,N_18150,N_17913);
or U20847 (N_20847,N_16837,N_16940);
or U20848 (N_20848,N_17969,N_18625);
nor U20849 (N_20849,N_17425,N_18106);
and U20850 (N_20850,N_17414,N_15832);
xor U20851 (N_20851,N_18683,N_16679);
and U20852 (N_20852,N_18261,N_16655);
or U20853 (N_20853,N_17954,N_16037);
nand U20854 (N_20854,N_15840,N_16415);
nand U20855 (N_20855,N_17781,N_15730);
nand U20856 (N_20856,N_16384,N_18097);
or U20857 (N_20857,N_15986,N_15931);
nand U20858 (N_20858,N_17890,N_16506);
nor U20859 (N_20859,N_15635,N_18699);
nand U20860 (N_20860,N_15690,N_17796);
nand U20861 (N_20861,N_17310,N_17109);
and U20862 (N_20862,N_18748,N_18385);
or U20863 (N_20863,N_17629,N_18630);
nor U20864 (N_20864,N_18442,N_16189);
or U20865 (N_20865,N_15789,N_17890);
or U20866 (N_20866,N_15822,N_16361);
or U20867 (N_20867,N_16156,N_18124);
or U20868 (N_20868,N_17058,N_17577);
xor U20869 (N_20869,N_15912,N_16335);
or U20870 (N_20870,N_18240,N_17340);
xor U20871 (N_20871,N_17095,N_15963);
nand U20872 (N_20872,N_17177,N_17026);
nor U20873 (N_20873,N_17430,N_15899);
or U20874 (N_20874,N_15986,N_18234);
or U20875 (N_20875,N_17771,N_16564);
nor U20876 (N_20876,N_15794,N_16321);
or U20877 (N_20877,N_15680,N_15815);
and U20878 (N_20878,N_16569,N_17846);
nand U20879 (N_20879,N_18645,N_16711);
nor U20880 (N_20880,N_18454,N_18121);
nor U20881 (N_20881,N_16351,N_16407);
xor U20882 (N_20882,N_16730,N_16881);
or U20883 (N_20883,N_17136,N_18163);
and U20884 (N_20884,N_16919,N_16629);
xor U20885 (N_20885,N_18656,N_15938);
nor U20886 (N_20886,N_18271,N_17137);
or U20887 (N_20887,N_18037,N_15860);
xor U20888 (N_20888,N_18299,N_17976);
and U20889 (N_20889,N_15913,N_18700);
xnor U20890 (N_20890,N_15932,N_16844);
xnor U20891 (N_20891,N_16029,N_16346);
and U20892 (N_20892,N_18694,N_17055);
and U20893 (N_20893,N_17796,N_18708);
nor U20894 (N_20894,N_17657,N_17021);
xnor U20895 (N_20895,N_17772,N_17715);
nor U20896 (N_20896,N_16789,N_16988);
xor U20897 (N_20897,N_18013,N_17600);
or U20898 (N_20898,N_18623,N_17791);
or U20899 (N_20899,N_16394,N_18028);
nor U20900 (N_20900,N_17515,N_18167);
xnor U20901 (N_20901,N_17732,N_15907);
and U20902 (N_20902,N_15750,N_17963);
and U20903 (N_20903,N_17472,N_18169);
nor U20904 (N_20904,N_17219,N_18631);
nand U20905 (N_20905,N_15766,N_17822);
xnor U20906 (N_20906,N_17667,N_17934);
or U20907 (N_20907,N_17224,N_17781);
and U20908 (N_20908,N_17974,N_18345);
xor U20909 (N_20909,N_18358,N_18642);
and U20910 (N_20910,N_16581,N_18127);
xor U20911 (N_20911,N_15646,N_17927);
nand U20912 (N_20912,N_17075,N_18636);
nand U20913 (N_20913,N_17195,N_16480);
or U20914 (N_20914,N_18095,N_17196);
or U20915 (N_20915,N_17088,N_18218);
or U20916 (N_20916,N_15965,N_17923);
or U20917 (N_20917,N_16114,N_18304);
nand U20918 (N_20918,N_16233,N_17419);
xnor U20919 (N_20919,N_16371,N_17202);
nor U20920 (N_20920,N_16263,N_16531);
and U20921 (N_20921,N_17164,N_16159);
nor U20922 (N_20922,N_15656,N_17298);
and U20923 (N_20923,N_17154,N_18361);
and U20924 (N_20924,N_18687,N_18565);
or U20925 (N_20925,N_18478,N_17562);
nand U20926 (N_20926,N_18365,N_16352);
xnor U20927 (N_20927,N_16325,N_16051);
nand U20928 (N_20928,N_18588,N_17310);
xor U20929 (N_20929,N_17686,N_17318);
xnor U20930 (N_20930,N_16722,N_18455);
nand U20931 (N_20931,N_16468,N_17909);
xnor U20932 (N_20932,N_17435,N_18717);
and U20933 (N_20933,N_16531,N_15904);
or U20934 (N_20934,N_15857,N_15779);
or U20935 (N_20935,N_18189,N_18029);
or U20936 (N_20936,N_15641,N_15642);
xnor U20937 (N_20937,N_17400,N_16781);
nor U20938 (N_20938,N_16722,N_16468);
and U20939 (N_20939,N_15743,N_16513);
nand U20940 (N_20940,N_18077,N_18009);
or U20941 (N_20941,N_17700,N_15793);
nand U20942 (N_20942,N_17143,N_17573);
xor U20943 (N_20943,N_18014,N_16495);
nand U20944 (N_20944,N_16241,N_17541);
or U20945 (N_20945,N_17579,N_17789);
xor U20946 (N_20946,N_16643,N_15739);
and U20947 (N_20947,N_17652,N_16021);
nor U20948 (N_20948,N_16402,N_16981);
nor U20949 (N_20949,N_16807,N_17175);
or U20950 (N_20950,N_16559,N_17481);
xor U20951 (N_20951,N_16510,N_18610);
and U20952 (N_20952,N_17775,N_18539);
nand U20953 (N_20953,N_15738,N_17987);
xnor U20954 (N_20954,N_17171,N_16731);
and U20955 (N_20955,N_17069,N_16124);
nor U20956 (N_20956,N_15754,N_15985);
xor U20957 (N_20957,N_18311,N_18601);
or U20958 (N_20958,N_17124,N_16809);
nor U20959 (N_20959,N_16889,N_17146);
xnor U20960 (N_20960,N_16852,N_15747);
or U20961 (N_20961,N_18636,N_17723);
or U20962 (N_20962,N_17529,N_18203);
nand U20963 (N_20963,N_15864,N_16437);
nor U20964 (N_20964,N_18525,N_17612);
nor U20965 (N_20965,N_16651,N_16982);
nor U20966 (N_20966,N_17380,N_15781);
and U20967 (N_20967,N_15856,N_16885);
nand U20968 (N_20968,N_17661,N_18340);
xnor U20969 (N_20969,N_17602,N_16417);
and U20970 (N_20970,N_18564,N_16876);
nor U20971 (N_20971,N_16908,N_15797);
xor U20972 (N_20972,N_17664,N_16936);
xor U20973 (N_20973,N_18544,N_17812);
and U20974 (N_20974,N_17351,N_18128);
or U20975 (N_20975,N_18557,N_15803);
xor U20976 (N_20976,N_15984,N_15719);
or U20977 (N_20977,N_15954,N_18157);
xor U20978 (N_20978,N_16031,N_18517);
and U20979 (N_20979,N_16353,N_16021);
and U20980 (N_20980,N_17310,N_18038);
nor U20981 (N_20981,N_16893,N_17110);
and U20982 (N_20982,N_17270,N_17115);
nand U20983 (N_20983,N_17266,N_17537);
xnor U20984 (N_20984,N_16012,N_16117);
xor U20985 (N_20985,N_16025,N_18118);
xor U20986 (N_20986,N_18133,N_18015);
xor U20987 (N_20987,N_16730,N_16573);
nor U20988 (N_20988,N_16399,N_18332);
xor U20989 (N_20989,N_16211,N_17980);
or U20990 (N_20990,N_18319,N_15786);
nand U20991 (N_20991,N_16967,N_17538);
or U20992 (N_20992,N_15872,N_16757);
nor U20993 (N_20993,N_18251,N_17663);
and U20994 (N_20994,N_16157,N_16092);
nor U20995 (N_20995,N_16725,N_16868);
nor U20996 (N_20996,N_17714,N_16442);
nand U20997 (N_20997,N_16340,N_15956);
nor U20998 (N_20998,N_15755,N_18160);
nor U20999 (N_20999,N_17148,N_17759);
or U21000 (N_21000,N_16227,N_17958);
nor U21001 (N_21001,N_16417,N_17589);
nand U21002 (N_21002,N_15851,N_17359);
nor U21003 (N_21003,N_17164,N_17924);
or U21004 (N_21004,N_15782,N_17356);
nor U21005 (N_21005,N_16291,N_15909);
and U21006 (N_21006,N_17691,N_18685);
or U21007 (N_21007,N_16169,N_15800);
nor U21008 (N_21008,N_18676,N_17709);
xnor U21009 (N_21009,N_16754,N_15891);
nor U21010 (N_21010,N_17146,N_17062);
nand U21011 (N_21011,N_18519,N_16652);
nand U21012 (N_21012,N_18618,N_16823);
xnor U21013 (N_21013,N_17146,N_16961);
or U21014 (N_21014,N_16534,N_16776);
nand U21015 (N_21015,N_17836,N_15912);
nand U21016 (N_21016,N_15783,N_18609);
nand U21017 (N_21017,N_17318,N_15874);
nand U21018 (N_21018,N_18548,N_17878);
xnor U21019 (N_21019,N_17980,N_17820);
nor U21020 (N_21020,N_17459,N_16861);
or U21021 (N_21021,N_16600,N_17724);
and U21022 (N_21022,N_18646,N_17553);
nand U21023 (N_21023,N_16577,N_16282);
nand U21024 (N_21024,N_18663,N_16557);
nor U21025 (N_21025,N_16090,N_17460);
xnor U21026 (N_21026,N_17209,N_18342);
nand U21027 (N_21027,N_17911,N_17485);
and U21028 (N_21028,N_16366,N_15639);
xnor U21029 (N_21029,N_17931,N_16133);
nand U21030 (N_21030,N_15825,N_16630);
and U21031 (N_21031,N_16488,N_15752);
nand U21032 (N_21032,N_18450,N_15693);
nand U21033 (N_21033,N_18227,N_15913);
and U21034 (N_21034,N_18343,N_16212);
nand U21035 (N_21035,N_17279,N_15885);
nor U21036 (N_21036,N_15639,N_15659);
nand U21037 (N_21037,N_17370,N_18425);
and U21038 (N_21038,N_17846,N_17321);
nor U21039 (N_21039,N_17208,N_16911);
nor U21040 (N_21040,N_18609,N_17699);
xnor U21041 (N_21041,N_18521,N_15812);
nand U21042 (N_21042,N_17774,N_18416);
xor U21043 (N_21043,N_16858,N_18215);
xnor U21044 (N_21044,N_17976,N_16290);
nor U21045 (N_21045,N_17468,N_17201);
nor U21046 (N_21046,N_17893,N_17344);
xor U21047 (N_21047,N_17019,N_17236);
or U21048 (N_21048,N_17082,N_18519);
and U21049 (N_21049,N_17023,N_16237);
nand U21050 (N_21050,N_16557,N_18558);
nor U21051 (N_21051,N_16140,N_17777);
nand U21052 (N_21052,N_16347,N_18232);
nand U21053 (N_21053,N_16110,N_17941);
or U21054 (N_21054,N_18312,N_17532);
nand U21055 (N_21055,N_16605,N_16140);
and U21056 (N_21056,N_17147,N_17001);
nor U21057 (N_21057,N_18197,N_16414);
xnor U21058 (N_21058,N_18332,N_17320);
xnor U21059 (N_21059,N_16169,N_16412);
and U21060 (N_21060,N_18479,N_17119);
and U21061 (N_21061,N_17094,N_17959);
xor U21062 (N_21062,N_18643,N_16068);
or U21063 (N_21063,N_17975,N_18535);
and U21064 (N_21064,N_17378,N_15785);
nand U21065 (N_21065,N_18061,N_16944);
nor U21066 (N_21066,N_17167,N_16738);
and U21067 (N_21067,N_16541,N_15942);
xnor U21068 (N_21068,N_16450,N_15708);
or U21069 (N_21069,N_18288,N_18103);
nand U21070 (N_21070,N_18477,N_17699);
or U21071 (N_21071,N_17540,N_15951);
or U21072 (N_21072,N_16224,N_18498);
nand U21073 (N_21073,N_16811,N_16656);
and U21074 (N_21074,N_16836,N_17696);
and U21075 (N_21075,N_16579,N_17645);
or U21076 (N_21076,N_16645,N_17956);
or U21077 (N_21077,N_17900,N_16900);
nand U21078 (N_21078,N_16590,N_17407);
or U21079 (N_21079,N_16736,N_17701);
nor U21080 (N_21080,N_18697,N_15756);
nand U21081 (N_21081,N_17944,N_17402);
xnor U21082 (N_21082,N_16256,N_16749);
or U21083 (N_21083,N_16480,N_16059);
xor U21084 (N_21084,N_17040,N_17558);
and U21085 (N_21085,N_18345,N_15795);
or U21086 (N_21086,N_15963,N_16667);
xor U21087 (N_21087,N_18740,N_16283);
and U21088 (N_21088,N_16052,N_16160);
nor U21089 (N_21089,N_15639,N_16193);
nor U21090 (N_21090,N_18264,N_18419);
and U21091 (N_21091,N_16944,N_16466);
nand U21092 (N_21092,N_17201,N_16685);
nor U21093 (N_21093,N_17757,N_16219);
xor U21094 (N_21094,N_18589,N_18695);
xnor U21095 (N_21095,N_17942,N_17720);
and U21096 (N_21096,N_16291,N_16137);
xor U21097 (N_21097,N_15910,N_15786);
nand U21098 (N_21098,N_18027,N_18226);
xor U21099 (N_21099,N_17924,N_17537);
nor U21100 (N_21100,N_17344,N_17920);
nand U21101 (N_21101,N_16021,N_15772);
or U21102 (N_21102,N_18574,N_17958);
and U21103 (N_21103,N_17523,N_17157);
nand U21104 (N_21104,N_17550,N_16507);
nor U21105 (N_21105,N_17859,N_18530);
xnor U21106 (N_21106,N_16204,N_17373);
nand U21107 (N_21107,N_16997,N_16995);
or U21108 (N_21108,N_17779,N_17411);
and U21109 (N_21109,N_16120,N_15837);
nand U21110 (N_21110,N_16114,N_17836);
nor U21111 (N_21111,N_17779,N_16400);
xor U21112 (N_21112,N_18419,N_16628);
or U21113 (N_21113,N_18260,N_18610);
xnor U21114 (N_21114,N_16864,N_15637);
nor U21115 (N_21115,N_15697,N_18255);
nor U21116 (N_21116,N_15653,N_15630);
xnor U21117 (N_21117,N_18679,N_17038);
nor U21118 (N_21118,N_15970,N_18027);
nand U21119 (N_21119,N_18441,N_17373);
or U21120 (N_21120,N_15717,N_17455);
or U21121 (N_21121,N_15949,N_18125);
nand U21122 (N_21122,N_16100,N_15687);
xnor U21123 (N_21123,N_18743,N_17868);
nor U21124 (N_21124,N_16442,N_16661);
xnor U21125 (N_21125,N_17201,N_16730);
or U21126 (N_21126,N_17712,N_16639);
nand U21127 (N_21127,N_16459,N_17714);
and U21128 (N_21128,N_18460,N_16775);
and U21129 (N_21129,N_18582,N_18540);
and U21130 (N_21130,N_17972,N_17007);
xnor U21131 (N_21131,N_16976,N_16883);
xnor U21132 (N_21132,N_15654,N_17869);
nor U21133 (N_21133,N_17461,N_18324);
and U21134 (N_21134,N_15896,N_17180);
nand U21135 (N_21135,N_16402,N_17828);
nand U21136 (N_21136,N_16581,N_18360);
nand U21137 (N_21137,N_17022,N_18112);
nor U21138 (N_21138,N_17768,N_18504);
nor U21139 (N_21139,N_16075,N_16424);
xnor U21140 (N_21140,N_18492,N_16497);
nor U21141 (N_21141,N_17373,N_16279);
nand U21142 (N_21142,N_16878,N_15645);
or U21143 (N_21143,N_16890,N_16309);
xnor U21144 (N_21144,N_17928,N_16834);
nor U21145 (N_21145,N_17803,N_17041);
or U21146 (N_21146,N_16084,N_18142);
xnor U21147 (N_21147,N_17513,N_16597);
and U21148 (N_21148,N_17100,N_16363);
nor U21149 (N_21149,N_16569,N_17638);
and U21150 (N_21150,N_16125,N_16098);
nand U21151 (N_21151,N_16583,N_17452);
and U21152 (N_21152,N_18583,N_16033);
and U21153 (N_21153,N_18173,N_15715);
nand U21154 (N_21154,N_15809,N_17858);
xor U21155 (N_21155,N_17088,N_17115);
or U21156 (N_21156,N_16250,N_16410);
nand U21157 (N_21157,N_16681,N_17513);
or U21158 (N_21158,N_18158,N_17407);
or U21159 (N_21159,N_18075,N_16104);
xor U21160 (N_21160,N_18213,N_17519);
and U21161 (N_21161,N_16706,N_16074);
nand U21162 (N_21162,N_15650,N_18043);
and U21163 (N_21163,N_17433,N_18220);
nor U21164 (N_21164,N_16318,N_16484);
or U21165 (N_21165,N_16227,N_15993);
xor U21166 (N_21166,N_17897,N_17459);
and U21167 (N_21167,N_16171,N_16308);
nor U21168 (N_21168,N_16432,N_18308);
nor U21169 (N_21169,N_16248,N_16483);
and U21170 (N_21170,N_18166,N_18302);
xor U21171 (N_21171,N_17400,N_18618);
and U21172 (N_21172,N_18378,N_17492);
xnor U21173 (N_21173,N_16075,N_17234);
and U21174 (N_21174,N_17166,N_18639);
xor U21175 (N_21175,N_17585,N_15723);
xnor U21176 (N_21176,N_15873,N_18691);
and U21177 (N_21177,N_16259,N_16060);
nand U21178 (N_21178,N_18103,N_16140);
or U21179 (N_21179,N_17700,N_17062);
nand U21180 (N_21180,N_16622,N_18407);
or U21181 (N_21181,N_16343,N_17545);
nand U21182 (N_21182,N_17991,N_15829);
or U21183 (N_21183,N_17722,N_15908);
xor U21184 (N_21184,N_18284,N_16673);
xnor U21185 (N_21185,N_17097,N_16859);
nand U21186 (N_21186,N_15974,N_16390);
and U21187 (N_21187,N_16188,N_18602);
or U21188 (N_21188,N_16029,N_16769);
nand U21189 (N_21189,N_16621,N_16246);
nand U21190 (N_21190,N_17404,N_17368);
nand U21191 (N_21191,N_17225,N_15654);
and U21192 (N_21192,N_17987,N_17300);
nor U21193 (N_21193,N_16020,N_17329);
nand U21194 (N_21194,N_16585,N_16891);
or U21195 (N_21195,N_16951,N_16568);
and U21196 (N_21196,N_16514,N_18621);
or U21197 (N_21197,N_17916,N_15971);
nand U21198 (N_21198,N_15631,N_17758);
nand U21199 (N_21199,N_16020,N_15758);
xnor U21200 (N_21200,N_17805,N_17041);
nand U21201 (N_21201,N_18263,N_16366);
nor U21202 (N_21202,N_16568,N_18650);
nand U21203 (N_21203,N_15704,N_15964);
and U21204 (N_21204,N_16354,N_18131);
and U21205 (N_21205,N_18563,N_18024);
nand U21206 (N_21206,N_18276,N_17518);
nand U21207 (N_21207,N_16498,N_17599);
xnor U21208 (N_21208,N_17599,N_17019);
nand U21209 (N_21209,N_18193,N_15991);
xnor U21210 (N_21210,N_15832,N_17752);
xnor U21211 (N_21211,N_17373,N_15873);
or U21212 (N_21212,N_17343,N_16621);
and U21213 (N_21213,N_16255,N_18486);
and U21214 (N_21214,N_16468,N_17637);
and U21215 (N_21215,N_17283,N_17959);
nor U21216 (N_21216,N_18116,N_16021);
or U21217 (N_21217,N_16159,N_18671);
nor U21218 (N_21218,N_17794,N_16444);
and U21219 (N_21219,N_17519,N_16515);
nand U21220 (N_21220,N_16380,N_15782);
nand U21221 (N_21221,N_17554,N_16737);
and U21222 (N_21222,N_18297,N_18535);
and U21223 (N_21223,N_18511,N_17816);
nor U21224 (N_21224,N_16119,N_16737);
nand U21225 (N_21225,N_16821,N_16517);
nor U21226 (N_21226,N_18176,N_16180);
nand U21227 (N_21227,N_17210,N_18390);
nor U21228 (N_21228,N_16035,N_16466);
or U21229 (N_21229,N_18632,N_16132);
xnor U21230 (N_21230,N_17198,N_16999);
and U21231 (N_21231,N_15772,N_17127);
xnor U21232 (N_21232,N_17459,N_18077);
xnor U21233 (N_21233,N_16817,N_18247);
nor U21234 (N_21234,N_16762,N_15998);
nand U21235 (N_21235,N_17036,N_17706);
xor U21236 (N_21236,N_16009,N_16695);
nand U21237 (N_21237,N_16568,N_18409);
nor U21238 (N_21238,N_17375,N_16940);
nand U21239 (N_21239,N_18083,N_16709);
nand U21240 (N_21240,N_15962,N_17482);
nor U21241 (N_21241,N_17463,N_17630);
xnor U21242 (N_21242,N_15802,N_18611);
xnor U21243 (N_21243,N_18476,N_16824);
xor U21244 (N_21244,N_18600,N_17999);
xnor U21245 (N_21245,N_18643,N_17825);
xor U21246 (N_21246,N_18268,N_18126);
and U21247 (N_21247,N_17296,N_18446);
nand U21248 (N_21248,N_18588,N_16422);
or U21249 (N_21249,N_18672,N_16323);
or U21250 (N_21250,N_16413,N_18354);
nor U21251 (N_21251,N_17238,N_18066);
and U21252 (N_21252,N_17213,N_15740);
and U21253 (N_21253,N_17184,N_18748);
and U21254 (N_21254,N_18689,N_17997);
nor U21255 (N_21255,N_16472,N_18704);
or U21256 (N_21256,N_17544,N_17164);
xor U21257 (N_21257,N_18391,N_18691);
nor U21258 (N_21258,N_17888,N_17603);
nand U21259 (N_21259,N_18284,N_16514);
nor U21260 (N_21260,N_16807,N_15897);
and U21261 (N_21261,N_17545,N_18638);
or U21262 (N_21262,N_18385,N_17591);
xor U21263 (N_21263,N_15845,N_15753);
and U21264 (N_21264,N_17785,N_17116);
or U21265 (N_21265,N_16581,N_17160);
nor U21266 (N_21266,N_17269,N_17707);
xor U21267 (N_21267,N_15834,N_17331);
xor U21268 (N_21268,N_18383,N_17576);
or U21269 (N_21269,N_18214,N_16865);
nand U21270 (N_21270,N_18654,N_18171);
nor U21271 (N_21271,N_17165,N_18627);
xor U21272 (N_21272,N_18423,N_17014);
nand U21273 (N_21273,N_16323,N_16818);
and U21274 (N_21274,N_16936,N_16520);
or U21275 (N_21275,N_15925,N_18420);
and U21276 (N_21276,N_17205,N_15701);
or U21277 (N_21277,N_16358,N_17207);
xnor U21278 (N_21278,N_18515,N_17962);
xnor U21279 (N_21279,N_17876,N_15806);
xor U21280 (N_21280,N_17878,N_18741);
xor U21281 (N_21281,N_17240,N_18213);
nor U21282 (N_21282,N_18406,N_17651);
or U21283 (N_21283,N_15923,N_16976);
nor U21284 (N_21284,N_16089,N_16005);
nand U21285 (N_21285,N_16446,N_18488);
nor U21286 (N_21286,N_16358,N_16014);
and U21287 (N_21287,N_17365,N_17596);
nor U21288 (N_21288,N_16319,N_16566);
and U21289 (N_21289,N_17502,N_15788);
nor U21290 (N_21290,N_17413,N_17591);
nor U21291 (N_21291,N_17001,N_17623);
xor U21292 (N_21292,N_17190,N_17168);
xor U21293 (N_21293,N_17341,N_17897);
xor U21294 (N_21294,N_15923,N_16579);
or U21295 (N_21295,N_18673,N_17207);
xor U21296 (N_21296,N_16115,N_17384);
or U21297 (N_21297,N_16411,N_16061);
nor U21298 (N_21298,N_17482,N_18685);
or U21299 (N_21299,N_18392,N_16577);
xor U21300 (N_21300,N_17834,N_18656);
or U21301 (N_21301,N_18290,N_17546);
nand U21302 (N_21302,N_18152,N_16875);
or U21303 (N_21303,N_16932,N_18600);
nor U21304 (N_21304,N_16974,N_17193);
and U21305 (N_21305,N_16161,N_17584);
or U21306 (N_21306,N_18631,N_18709);
and U21307 (N_21307,N_16376,N_15941);
or U21308 (N_21308,N_18370,N_18692);
and U21309 (N_21309,N_18140,N_18614);
and U21310 (N_21310,N_17589,N_17694);
nand U21311 (N_21311,N_17807,N_16353);
and U21312 (N_21312,N_18430,N_18481);
xor U21313 (N_21313,N_15789,N_16805);
xor U21314 (N_21314,N_16771,N_18176);
nand U21315 (N_21315,N_16231,N_17055);
nor U21316 (N_21316,N_16412,N_16286);
or U21317 (N_21317,N_17953,N_17418);
nor U21318 (N_21318,N_16273,N_17522);
nand U21319 (N_21319,N_17615,N_18584);
and U21320 (N_21320,N_17837,N_18158);
or U21321 (N_21321,N_16461,N_16044);
xnor U21322 (N_21322,N_15745,N_18351);
or U21323 (N_21323,N_18475,N_18423);
and U21324 (N_21324,N_16052,N_17265);
or U21325 (N_21325,N_16611,N_18012);
and U21326 (N_21326,N_16912,N_17944);
or U21327 (N_21327,N_15972,N_18661);
nor U21328 (N_21328,N_18477,N_17080);
nor U21329 (N_21329,N_17129,N_17403);
or U21330 (N_21330,N_16178,N_16033);
or U21331 (N_21331,N_18154,N_16350);
or U21332 (N_21332,N_17918,N_18185);
xor U21333 (N_21333,N_16546,N_18433);
and U21334 (N_21334,N_16517,N_15628);
xor U21335 (N_21335,N_17578,N_17607);
xor U21336 (N_21336,N_17532,N_17637);
xnor U21337 (N_21337,N_18401,N_16987);
nand U21338 (N_21338,N_18112,N_17869);
or U21339 (N_21339,N_16113,N_18202);
and U21340 (N_21340,N_18262,N_16164);
or U21341 (N_21341,N_17168,N_17590);
or U21342 (N_21342,N_15972,N_18142);
nand U21343 (N_21343,N_17289,N_16676);
xnor U21344 (N_21344,N_18307,N_15630);
or U21345 (N_21345,N_17411,N_17131);
and U21346 (N_21346,N_15732,N_18357);
nor U21347 (N_21347,N_18530,N_18475);
nand U21348 (N_21348,N_16713,N_17616);
nand U21349 (N_21349,N_15779,N_17206);
nor U21350 (N_21350,N_18033,N_15852);
nand U21351 (N_21351,N_17810,N_17032);
xor U21352 (N_21352,N_16266,N_15802);
nor U21353 (N_21353,N_17997,N_15665);
xnor U21354 (N_21354,N_15761,N_16425);
nand U21355 (N_21355,N_16357,N_18263);
nor U21356 (N_21356,N_16098,N_17441);
xor U21357 (N_21357,N_16739,N_17058);
xnor U21358 (N_21358,N_16624,N_17140);
nor U21359 (N_21359,N_17761,N_17038);
nand U21360 (N_21360,N_15672,N_16878);
or U21361 (N_21361,N_17278,N_18724);
xnor U21362 (N_21362,N_18447,N_18233);
xor U21363 (N_21363,N_15879,N_18364);
xnor U21364 (N_21364,N_16772,N_17146);
or U21365 (N_21365,N_18407,N_16038);
and U21366 (N_21366,N_17484,N_17358);
nor U21367 (N_21367,N_17112,N_15862);
nor U21368 (N_21368,N_17533,N_15910);
xnor U21369 (N_21369,N_17758,N_17044);
or U21370 (N_21370,N_17251,N_17445);
or U21371 (N_21371,N_16122,N_16295);
or U21372 (N_21372,N_18505,N_16368);
nand U21373 (N_21373,N_17857,N_15675);
xor U21374 (N_21374,N_16033,N_17416);
and U21375 (N_21375,N_18228,N_15983);
nand U21376 (N_21376,N_17865,N_16368);
or U21377 (N_21377,N_18190,N_16778);
xor U21378 (N_21378,N_16752,N_15964);
and U21379 (N_21379,N_17585,N_16959);
xnor U21380 (N_21380,N_17984,N_17726);
nor U21381 (N_21381,N_16384,N_16998);
nor U21382 (N_21382,N_18235,N_18558);
nor U21383 (N_21383,N_17478,N_17837);
or U21384 (N_21384,N_18573,N_16149);
or U21385 (N_21385,N_17248,N_16888);
nand U21386 (N_21386,N_16105,N_17900);
xor U21387 (N_21387,N_17425,N_16241);
xnor U21388 (N_21388,N_15759,N_15991);
nand U21389 (N_21389,N_16570,N_16060);
and U21390 (N_21390,N_16218,N_16999);
or U21391 (N_21391,N_17008,N_16570);
xnor U21392 (N_21392,N_16924,N_16732);
nand U21393 (N_21393,N_17814,N_17671);
nor U21394 (N_21394,N_16153,N_18178);
nand U21395 (N_21395,N_17641,N_18739);
nand U21396 (N_21396,N_17602,N_17129);
xnor U21397 (N_21397,N_17204,N_17737);
and U21398 (N_21398,N_16025,N_16331);
xor U21399 (N_21399,N_17947,N_15788);
xor U21400 (N_21400,N_16308,N_17120);
nor U21401 (N_21401,N_17923,N_15779);
nand U21402 (N_21402,N_16748,N_18332);
xnor U21403 (N_21403,N_18482,N_17347);
nand U21404 (N_21404,N_17000,N_17458);
xor U21405 (N_21405,N_17638,N_17913);
and U21406 (N_21406,N_15701,N_16835);
and U21407 (N_21407,N_18339,N_17614);
xor U21408 (N_21408,N_17050,N_17172);
xnor U21409 (N_21409,N_18047,N_17429);
nand U21410 (N_21410,N_15652,N_16366);
nor U21411 (N_21411,N_17996,N_16667);
nor U21412 (N_21412,N_15900,N_17220);
nand U21413 (N_21413,N_16208,N_17562);
nand U21414 (N_21414,N_16604,N_16814);
or U21415 (N_21415,N_16115,N_18559);
or U21416 (N_21416,N_17727,N_17856);
or U21417 (N_21417,N_17704,N_18309);
nand U21418 (N_21418,N_18178,N_16204);
xor U21419 (N_21419,N_16858,N_18595);
nand U21420 (N_21420,N_17578,N_17860);
and U21421 (N_21421,N_16298,N_16439);
xnor U21422 (N_21422,N_17210,N_16373);
nor U21423 (N_21423,N_18521,N_15789);
nor U21424 (N_21424,N_18025,N_17797);
xor U21425 (N_21425,N_17954,N_16084);
xor U21426 (N_21426,N_16455,N_15890);
nand U21427 (N_21427,N_18326,N_16444);
nor U21428 (N_21428,N_18100,N_16593);
nand U21429 (N_21429,N_18102,N_17931);
nor U21430 (N_21430,N_17154,N_17772);
and U21431 (N_21431,N_15754,N_18376);
and U21432 (N_21432,N_18259,N_16692);
xor U21433 (N_21433,N_16753,N_16189);
and U21434 (N_21434,N_18314,N_16095);
nor U21435 (N_21435,N_15659,N_18093);
xor U21436 (N_21436,N_16550,N_16790);
nor U21437 (N_21437,N_16799,N_16429);
or U21438 (N_21438,N_17833,N_17812);
and U21439 (N_21439,N_16626,N_17162);
and U21440 (N_21440,N_16277,N_16391);
xnor U21441 (N_21441,N_15886,N_17227);
and U21442 (N_21442,N_16729,N_17549);
or U21443 (N_21443,N_16457,N_18051);
xnor U21444 (N_21444,N_16927,N_18256);
nand U21445 (N_21445,N_17507,N_15674);
and U21446 (N_21446,N_16636,N_18028);
nor U21447 (N_21447,N_17758,N_16063);
and U21448 (N_21448,N_17849,N_16434);
nor U21449 (N_21449,N_16076,N_16523);
nor U21450 (N_21450,N_17028,N_17505);
and U21451 (N_21451,N_18623,N_16894);
or U21452 (N_21452,N_16061,N_17987);
nor U21453 (N_21453,N_16344,N_18365);
or U21454 (N_21454,N_16508,N_15812);
nand U21455 (N_21455,N_16111,N_16145);
nor U21456 (N_21456,N_18339,N_16752);
or U21457 (N_21457,N_17143,N_18266);
xor U21458 (N_21458,N_18687,N_16322);
nor U21459 (N_21459,N_16591,N_16181);
and U21460 (N_21460,N_17887,N_18434);
and U21461 (N_21461,N_17259,N_17254);
nand U21462 (N_21462,N_16627,N_16601);
xor U21463 (N_21463,N_17159,N_15788);
nand U21464 (N_21464,N_18314,N_15777);
xor U21465 (N_21465,N_17372,N_17156);
and U21466 (N_21466,N_17624,N_17454);
and U21467 (N_21467,N_16161,N_15850);
nor U21468 (N_21468,N_17226,N_18201);
or U21469 (N_21469,N_17983,N_17416);
nand U21470 (N_21470,N_16583,N_17857);
and U21471 (N_21471,N_17372,N_18408);
or U21472 (N_21472,N_15831,N_15972);
nand U21473 (N_21473,N_17818,N_15735);
xor U21474 (N_21474,N_17133,N_18596);
nand U21475 (N_21475,N_17472,N_17844);
or U21476 (N_21476,N_15916,N_16923);
or U21477 (N_21477,N_16847,N_18320);
or U21478 (N_21478,N_17051,N_18741);
or U21479 (N_21479,N_17324,N_17141);
nand U21480 (N_21480,N_16877,N_16573);
or U21481 (N_21481,N_18083,N_16685);
and U21482 (N_21482,N_16291,N_18322);
and U21483 (N_21483,N_18583,N_15861);
nor U21484 (N_21484,N_18039,N_15913);
xnor U21485 (N_21485,N_17268,N_16849);
or U21486 (N_21486,N_18738,N_18551);
nand U21487 (N_21487,N_17904,N_17788);
nand U21488 (N_21488,N_17274,N_16641);
nor U21489 (N_21489,N_17952,N_18374);
xor U21490 (N_21490,N_17071,N_17856);
and U21491 (N_21491,N_16696,N_18587);
and U21492 (N_21492,N_17013,N_17829);
or U21493 (N_21493,N_18222,N_16833);
and U21494 (N_21494,N_17771,N_18435);
and U21495 (N_21495,N_16213,N_16223);
and U21496 (N_21496,N_17892,N_16305);
or U21497 (N_21497,N_18512,N_18459);
and U21498 (N_21498,N_16750,N_18108);
and U21499 (N_21499,N_15625,N_17916);
nor U21500 (N_21500,N_17540,N_16512);
and U21501 (N_21501,N_18578,N_15859);
nor U21502 (N_21502,N_18006,N_17639);
and U21503 (N_21503,N_18737,N_17106);
or U21504 (N_21504,N_15796,N_16685);
nand U21505 (N_21505,N_18124,N_16015);
xnor U21506 (N_21506,N_16996,N_16987);
or U21507 (N_21507,N_17227,N_17731);
or U21508 (N_21508,N_17833,N_18484);
nand U21509 (N_21509,N_17249,N_16003);
nand U21510 (N_21510,N_17246,N_16184);
or U21511 (N_21511,N_18321,N_18072);
nor U21512 (N_21512,N_18117,N_16983);
nand U21513 (N_21513,N_18236,N_16515);
nand U21514 (N_21514,N_15702,N_18262);
or U21515 (N_21515,N_16205,N_17220);
nand U21516 (N_21516,N_17072,N_15997);
nand U21517 (N_21517,N_15868,N_17973);
or U21518 (N_21518,N_17004,N_18583);
or U21519 (N_21519,N_16754,N_18678);
xor U21520 (N_21520,N_16783,N_18405);
and U21521 (N_21521,N_17826,N_17335);
nor U21522 (N_21522,N_18671,N_17819);
xor U21523 (N_21523,N_16770,N_17313);
or U21524 (N_21524,N_18176,N_16629);
and U21525 (N_21525,N_17712,N_16484);
nand U21526 (N_21526,N_18730,N_16940);
nand U21527 (N_21527,N_15681,N_17622);
and U21528 (N_21528,N_18024,N_16992);
and U21529 (N_21529,N_17905,N_16027);
xnor U21530 (N_21530,N_16614,N_16844);
nor U21531 (N_21531,N_15744,N_17962);
or U21532 (N_21532,N_17661,N_16373);
xor U21533 (N_21533,N_16985,N_15895);
nand U21534 (N_21534,N_18243,N_16780);
or U21535 (N_21535,N_17916,N_15795);
and U21536 (N_21536,N_17836,N_17076);
xor U21537 (N_21537,N_17010,N_17784);
nor U21538 (N_21538,N_16499,N_16818);
xnor U21539 (N_21539,N_18160,N_17161);
xor U21540 (N_21540,N_17653,N_16023);
nand U21541 (N_21541,N_18352,N_16302);
nand U21542 (N_21542,N_18461,N_17842);
nand U21543 (N_21543,N_17487,N_16145);
and U21544 (N_21544,N_17167,N_18391);
and U21545 (N_21545,N_18654,N_16941);
nor U21546 (N_21546,N_17329,N_16303);
or U21547 (N_21547,N_16559,N_18347);
or U21548 (N_21548,N_16773,N_17982);
nand U21549 (N_21549,N_15704,N_17608);
and U21550 (N_21550,N_18235,N_17645);
nor U21551 (N_21551,N_15986,N_17375);
nand U21552 (N_21552,N_18405,N_16611);
and U21553 (N_21553,N_16910,N_17823);
and U21554 (N_21554,N_18620,N_17881);
or U21555 (N_21555,N_16233,N_18103);
or U21556 (N_21556,N_18630,N_17704);
nand U21557 (N_21557,N_16130,N_16458);
or U21558 (N_21558,N_18456,N_16095);
nor U21559 (N_21559,N_17811,N_17846);
xnor U21560 (N_21560,N_15771,N_16181);
or U21561 (N_21561,N_18619,N_17117);
nor U21562 (N_21562,N_15941,N_18424);
and U21563 (N_21563,N_16183,N_18675);
nor U21564 (N_21564,N_17467,N_16279);
nor U21565 (N_21565,N_17127,N_17573);
and U21566 (N_21566,N_17916,N_18661);
or U21567 (N_21567,N_15894,N_17141);
xnor U21568 (N_21568,N_15673,N_16390);
and U21569 (N_21569,N_16204,N_16155);
nand U21570 (N_21570,N_18128,N_16813);
nor U21571 (N_21571,N_17868,N_17402);
or U21572 (N_21572,N_16774,N_17233);
xor U21573 (N_21573,N_17573,N_17449);
xnor U21574 (N_21574,N_17123,N_16980);
nor U21575 (N_21575,N_16504,N_18247);
nor U21576 (N_21576,N_18130,N_16789);
nand U21577 (N_21577,N_17043,N_17570);
xor U21578 (N_21578,N_17000,N_16031);
and U21579 (N_21579,N_17804,N_18307);
xnor U21580 (N_21580,N_16392,N_17115);
or U21581 (N_21581,N_15858,N_15986);
nor U21582 (N_21582,N_15802,N_18522);
nand U21583 (N_21583,N_17831,N_17077);
or U21584 (N_21584,N_16300,N_16217);
xor U21585 (N_21585,N_17875,N_18232);
or U21586 (N_21586,N_18462,N_17213);
nor U21587 (N_21587,N_16857,N_16255);
and U21588 (N_21588,N_17970,N_17571);
xor U21589 (N_21589,N_17106,N_16262);
xor U21590 (N_21590,N_16217,N_16936);
nand U21591 (N_21591,N_18031,N_16378);
and U21592 (N_21592,N_17203,N_18035);
nor U21593 (N_21593,N_17736,N_16161);
or U21594 (N_21594,N_18303,N_18331);
or U21595 (N_21595,N_17217,N_17559);
and U21596 (N_21596,N_15873,N_18301);
and U21597 (N_21597,N_15708,N_18730);
xnor U21598 (N_21598,N_17510,N_16801);
and U21599 (N_21599,N_17208,N_18510);
nor U21600 (N_21600,N_16457,N_16729);
xnor U21601 (N_21601,N_16932,N_17001);
nand U21602 (N_21602,N_15702,N_15966);
nand U21603 (N_21603,N_18534,N_16336);
nor U21604 (N_21604,N_16080,N_17270);
and U21605 (N_21605,N_17321,N_17200);
or U21606 (N_21606,N_17383,N_17653);
nor U21607 (N_21607,N_16104,N_16409);
nand U21608 (N_21608,N_15637,N_17398);
nand U21609 (N_21609,N_16264,N_16900);
nor U21610 (N_21610,N_18249,N_17881);
xnor U21611 (N_21611,N_16338,N_18041);
xor U21612 (N_21612,N_16316,N_18161);
nor U21613 (N_21613,N_18026,N_16014);
and U21614 (N_21614,N_18658,N_16996);
or U21615 (N_21615,N_17885,N_16473);
nor U21616 (N_21616,N_16727,N_17785);
and U21617 (N_21617,N_15850,N_17778);
and U21618 (N_21618,N_17385,N_15745);
or U21619 (N_21619,N_16809,N_16759);
nand U21620 (N_21620,N_17553,N_16294);
nor U21621 (N_21621,N_17352,N_16791);
nor U21622 (N_21622,N_15966,N_18676);
or U21623 (N_21623,N_16027,N_17833);
and U21624 (N_21624,N_17698,N_16894);
or U21625 (N_21625,N_17809,N_17712);
nor U21626 (N_21626,N_17816,N_17359);
nand U21627 (N_21627,N_18189,N_17644);
nor U21628 (N_21628,N_16570,N_18081);
nor U21629 (N_21629,N_16147,N_16399);
nor U21630 (N_21630,N_17480,N_15628);
and U21631 (N_21631,N_15697,N_18622);
xnor U21632 (N_21632,N_18745,N_18133);
or U21633 (N_21633,N_18530,N_16223);
xor U21634 (N_21634,N_16029,N_17776);
or U21635 (N_21635,N_17057,N_17528);
or U21636 (N_21636,N_16247,N_15979);
xor U21637 (N_21637,N_17933,N_16786);
and U21638 (N_21638,N_17658,N_16632);
nand U21639 (N_21639,N_18414,N_17971);
nor U21640 (N_21640,N_18093,N_17388);
xnor U21641 (N_21641,N_17572,N_16117);
xnor U21642 (N_21642,N_17270,N_16872);
nor U21643 (N_21643,N_17448,N_16129);
nand U21644 (N_21644,N_16691,N_16363);
xor U21645 (N_21645,N_18074,N_16790);
xnor U21646 (N_21646,N_18031,N_16095);
nor U21647 (N_21647,N_17910,N_17761);
nor U21648 (N_21648,N_17352,N_18575);
xor U21649 (N_21649,N_16433,N_16406);
or U21650 (N_21650,N_18441,N_18286);
nand U21651 (N_21651,N_18334,N_17543);
xnor U21652 (N_21652,N_18455,N_18597);
nor U21653 (N_21653,N_16424,N_17494);
or U21654 (N_21654,N_17657,N_16701);
and U21655 (N_21655,N_18465,N_17912);
and U21656 (N_21656,N_17233,N_18590);
nand U21657 (N_21657,N_16693,N_18558);
or U21658 (N_21658,N_15833,N_16787);
nand U21659 (N_21659,N_17000,N_16838);
or U21660 (N_21660,N_16232,N_18131);
and U21661 (N_21661,N_18393,N_15970);
nor U21662 (N_21662,N_16664,N_16326);
or U21663 (N_21663,N_16780,N_16658);
and U21664 (N_21664,N_17487,N_17595);
nor U21665 (N_21665,N_17666,N_17009);
xnor U21666 (N_21666,N_16472,N_16736);
and U21667 (N_21667,N_16097,N_16315);
nand U21668 (N_21668,N_17206,N_15653);
nor U21669 (N_21669,N_16692,N_18014);
xnor U21670 (N_21670,N_16880,N_16435);
nor U21671 (N_21671,N_17398,N_16058);
or U21672 (N_21672,N_15825,N_16157);
and U21673 (N_21673,N_16640,N_15890);
nand U21674 (N_21674,N_17701,N_17308);
xor U21675 (N_21675,N_16964,N_17529);
nor U21676 (N_21676,N_18134,N_16952);
nor U21677 (N_21677,N_17541,N_18463);
xor U21678 (N_21678,N_16508,N_16592);
xnor U21679 (N_21679,N_17907,N_16982);
nand U21680 (N_21680,N_15747,N_17428);
and U21681 (N_21681,N_17847,N_18343);
or U21682 (N_21682,N_17195,N_15995);
nor U21683 (N_21683,N_17156,N_16578);
nand U21684 (N_21684,N_18370,N_16084);
and U21685 (N_21685,N_15892,N_18540);
or U21686 (N_21686,N_15700,N_16296);
or U21687 (N_21687,N_16173,N_17849);
nand U21688 (N_21688,N_16620,N_18014);
or U21689 (N_21689,N_15662,N_17206);
xnor U21690 (N_21690,N_18303,N_15829);
or U21691 (N_21691,N_18651,N_17449);
nor U21692 (N_21692,N_15654,N_17451);
or U21693 (N_21693,N_18513,N_16209);
or U21694 (N_21694,N_18012,N_16043);
xor U21695 (N_21695,N_18469,N_18496);
and U21696 (N_21696,N_18229,N_18033);
and U21697 (N_21697,N_16478,N_17615);
xor U21698 (N_21698,N_15630,N_17446);
xor U21699 (N_21699,N_16988,N_18301);
nor U21700 (N_21700,N_18222,N_16850);
xor U21701 (N_21701,N_17540,N_18047);
and U21702 (N_21702,N_18309,N_15649);
nand U21703 (N_21703,N_18365,N_16520);
nor U21704 (N_21704,N_16884,N_16398);
and U21705 (N_21705,N_18416,N_18342);
and U21706 (N_21706,N_16288,N_17874);
and U21707 (N_21707,N_17030,N_16296);
and U21708 (N_21708,N_17316,N_17352);
nor U21709 (N_21709,N_18121,N_17464);
and U21710 (N_21710,N_15680,N_16719);
nor U21711 (N_21711,N_16092,N_17000);
nand U21712 (N_21712,N_17588,N_18483);
xor U21713 (N_21713,N_15962,N_18276);
or U21714 (N_21714,N_17884,N_18569);
and U21715 (N_21715,N_18655,N_17138);
nand U21716 (N_21716,N_18423,N_18288);
or U21717 (N_21717,N_18695,N_18444);
xor U21718 (N_21718,N_18472,N_18407);
nand U21719 (N_21719,N_17114,N_16845);
nor U21720 (N_21720,N_15914,N_17931);
xnor U21721 (N_21721,N_17770,N_16474);
xnor U21722 (N_21722,N_18254,N_16859);
xor U21723 (N_21723,N_17531,N_18028);
or U21724 (N_21724,N_17336,N_16054);
or U21725 (N_21725,N_16986,N_16571);
nand U21726 (N_21726,N_18166,N_16981);
nand U21727 (N_21727,N_18706,N_17307);
nor U21728 (N_21728,N_17589,N_17690);
or U21729 (N_21729,N_18581,N_17738);
nand U21730 (N_21730,N_17951,N_18659);
or U21731 (N_21731,N_16988,N_17930);
nor U21732 (N_21732,N_17360,N_16704);
or U21733 (N_21733,N_16242,N_16365);
and U21734 (N_21734,N_17400,N_17466);
and U21735 (N_21735,N_16703,N_18385);
nor U21736 (N_21736,N_17912,N_16921);
nand U21737 (N_21737,N_15852,N_16847);
and U21738 (N_21738,N_18483,N_16212);
xnor U21739 (N_21739,N_16282,N_17500);
nand U21740 (N_21740,N_17660,N_16019);
nand U21741 (N_21741,N_16568,N_18010);
or U21742 (N_21742,N_17003,N_18043);
nor U21743 (N_21743,N_18330,N_17688);
or U21744 (N_21744,N_17994,N_16860);
nand U21745 (N_21745,N_16241,N_16882);
nor U21746 (N_21746,N_15686,N_15898);
nor U21747 (N_21747,N_15807,N_15855);
nand U21748 (N_21748,N_17164,N_16596);
or U21749 (N_21749,N_17363,N_15798);
nor U21750 (N_21750,N_17309,N_17866);
xor U21751 (N_21751,N_16211,N_15707);
and U21752 (N_21752,N_16817,N_16219);
and U21753 (N_21753,N_16075,N_16213);
xnor U21754 (N_21754,N_16554,N_17786);
nor U21755 (N_21755,N_18583,N_18190);
and U21756 (N_21756,N_17311,N_17661);
nand U21757 (N_21757,N_15698,N_16049);
or U21758 (N_21758,N_18101,N_17943);
nand U21759 (N_21759,N_16585,N_15716);
and U21760 (N_21760,N_16676,N_18183);
and U21761 (N_21761,N_16352,N_16872);
and U21762 (N_21762,N_16413,N_16296);
nor U21763 (N_21763,N_16777,N_18046);
and U21764 (N_21764,N_16489,N_18721);
xnor U21765 (N_21765,N_17921,N_17145);
and U21766 (N_21766,N_18702,N_17784);
nand U21767 (N_21767,N_18297,N_17461);
or U21768 (N_21768,N_18313,N_16296);
xor U21769 (N_21769,N_17494,N_17260);
nor U21770 (N_21770,N_18011,N_18421);
nor U21771 (N_21771,N_16050,N_16228);
nand U21772 (N_21772,N_17805,N_15845);
or U21773 (N_21773,N_16437,N_18379);
and U21774 (N_21774,N_16683,N_15917);
or U21775 (N_21775,N_16881,N_16045);
nand U21776 (N_21776,N_16357,N_16401);
and U21777 (N_21777,N_18239,N_16340);
or U21778 (N_21778,N_16091,N_18362);
nor U21779 (N_21779,N_17135,N_18040);
nand U21780 (N_21780,N_16172,N_17282);
and U21781 (N_21781,N_17854,N_17543);
or U21782 (N_21782,N_16608,N_15636);
nor U21783 (N_21783,N_16678,N_18109);
or U21784 (N_21784,N_18014,N_16772);
or U21785 (N_21785,N_17943,N_15793);
or U21786 (N_21786,N_17195,N_17491);
nor U21787 (N_21787,N_16531,N_18007);
or U21788 (N_21788,N_16448,N_15655);
nand U21789 (N_21789,N_18332,N_17439);
nand U21790 (N_21790,N_16145,N_16690);
xnor U21791 (N_21791,N_16753,N_18186);
nand U21792 (N_21792,N_18077,N_17881);
xnor U21793 (N_21793,N_16842,N_18525);
or U21794 (N_21794,N_17045,N_16381);
xnor U21795 (N_21795,N_16121,N_18411);
nand U21796 (N_21796,N_17843,N_15690);
or U21797 (N_21797,N_18578,N_18174);
or U21798 (N_21798,N_16739,N_15719);
or U21799 (N_21799,N_16016,N_16934);
nor U21800 (N_21800,N_18140,N_18123);
or U21801 (N_21801,N_17779,N_18113);
nand U21802 (N_21802,N_16497,N_15673);
nor U21803 (N_21803,N_18715,N_16203);
or U21804 (N_21804,N_17805,N_17583);
nand U21805 (N_21805,N_17767,N_17611);
and U21806 (N_21806,N_18707,N_17909);
xor U21807 (N_21807,N_17161,N_16773);
nor U21808 (N_21808,N_17671,N_15720);
nand U21809 (N_21809,N_16602,N_17229);
xnor U21810 (N_21810,N_16465,N_16755);
and U21811 (N_21811,N_17087,N_18017);
nor U21812 (N_21812,N_15708,N_18697);
or U21813 (N_21813,N_17346,N_17365);
nor U21814 (N_21814,N_18499,N_18093);
nor U21815 (N_21815,N_15840,N_16524);
or U21816 (N_21816,N_15859,N_18655);
or U21817 (N_21817,N_18575,N_15627);
nand U21818 (N_21818,N_17728,N_15639);
nand U21819 (N_21819,N_17959,N_17556);
or U21820 (N_21820,N_18196,N_17232);
xnor U21821 (N_21821,N_17295,N_16658);
nand U21822 (N_21822,N_17548,N_16480);
nand U21823 (N_21823,N_18744,N_17391);
nor U21824 (N_21824,N_17001,N_18250);
nor U21825 (N_21825,N_16725,N_17828);
xor U21826 (N_21826,N_17095,N_16183);
and U21827 (N_21827,N_18548,N_15987);
nor U21828 (N_21828,N_17027,N_16863);
and U21829 (N_21829,N_16601,N_16784);
and U21830 (N_21830,N_15861,N_15738);
nand U21831 (N_21831,N_16537,N_16030);
or U21832 (N_21832,N_16652,N_18410);
xor U21833 (N_21833,N_18155,N_17008);
or U21834 (N_21834,N_18114,N_17779);
or U21835 (N_21835,N_18191,N_16913);
nand U21836 (N_21836,N_17970,N_15818);
nand U21837 (N_21837,N_17765,N_18269);
or U21838 (N_21838,N_16893,N_18297);
or U21839 (N_21839,N_16340,N_15921);
nor U21840 (N_21840,N_17142,N_16091);
or U21841 (N_21841,N_16778,N_17599);
xor U21842 (N_21842,N_17603,N_18351);
xnor U21843 (N_21843,N_16694,N_18029);
and U21844 (N_21844,N_16603,N_16610);
nor U21845 (N_21845,N_15737,N_16859);
nor U21846 (N_21846,N_17060,N_16912);
or U21847 (N_21847,N_18008,N_16969);
and U21848 (N_21848,N_16122,N_17835);
and U21849 (N_21849,N_17618,N_18535);
or U21850 (N_21850,N_18298,N_15893);
xor U21851 (N_21851,N_16134,N_17221);
or U21852 (N_21852,N_17049,N_17063);
and U21853 (N_21853,N_17282,N_18046);
or U21854 (N_21854,N_17602,N_17385);
xnor U21855 (N_21855,N_18094,N_18336);
or U21856 (N_21856,N_17124,N_18467);
nand U21857 (N_21857,N_18123,N_16011);
xor U21858 (N_21858,N_17126,N_16328);
or U21859 (N_21859,N_15898,N_16487);
or U21860 (N_21860,N_17940,N_18169);
or U21861 (N_21861,N_17255,N_16262);
nor U21862 (N_21862,N_17726,N_17077);
xor U21863 (N_21863,N_15919,N_17575);
xor U21864 (N_21864,N_16575,N_15710);
and U21865 (N_21865,N_17142,N_17772);
or U21866 (N_21866,N_18399,N_17139);
nand U21867 (N_21867,N_17092,N_17377);
and U21868 (N_21868,N_17293,N_17347);
and U21869 (N_21869,N_16384,N_17835);
xnor U21870 (N_21870,N_16936,N_16086);
and U21871 (N_21871,N_16938,N_16221);
nor U21872 (N_21872,N_18556,N_17148);
nand U21873 (N_21873,N_17890,N_18175);
nor U21874 (N_21874,N_15994,N_17546);
or U21875 (N_21875,N_19431,N_19148);
nor U21876 (N_21876,N_19281,N_21814);
nor U21877 (N_21877,N_19364,N_20217);
nand U21878 (N_21878,N_21229,N_20244);
nor U21879 (N_21879,N_19865,N_20147);
nand U21880 (N_21880,N_21401,N_18988);
nand U21881 (N_21881,N_19673,N_19903);
nand U21882 (N_21882,N_19217,N_19860);
and U21883 (N_21883,N_20569,N_21178);
and U21884 (N_21884,N_19773,N_19243);
xnor U21885 (N_21885,N_20196,N_20105);
and U21886 (N_21886,N_18956,N_20616);
nand U21887 (N_21887,N_20568,N_20353);
nor U21888 (N_21888,N_19782,N_21614);
nand U21889 (N_21889,N_21687,N_21249);
or U21890 (N_21890,N_19192,N_20931);
nor U21891 (N_21891,N_19664,N_21426);
nand U21892 (N_21892,N_21787,N_19048);
or U21893 (N_21893,N_19471,N_20175);
or U21894 (N_21894,N_19415,N_20608);
xnor U21895 (N_21895,N_18957,N_18796);
or U21896 (N_21896,N_20272,N_21655);
nor U21897 (N_21897,N_19232,N_20613);
or U21898 (N_21898,N_20752,N_20121);
nor U21899 (N_21899,N_20500,N_18824);
nand U21900 (N_21900,N_20982,N_19653);
xor U21901 (N_21901,N_19271,N_19660);
xnor U21902 (N_21902,N_19485,N_19985);
nand U21903 (N_21903,N_19374,N_18839);
nand U21904 (N_21904,N_19967,N_21350);
nor U21905 (N_21905,N_20660,N_20909);
nand U21906 (N_21906,N_19642,N_21721);
nor U21907 (N_21907,N_20502,N_21524);
xnor U21908 (N_21908,N_21000,N_20089);
nand U21909 (N_21909,N_18897,N_19173);
xnor U21910 (N_21910,N_21520,N_20872);
and U21911 (N_21911,N_21035,N_20580);
and U21912 (N_21912,N_21549,N_20544);
nor U21913 (N_21913,N_19868,N_19762);
xnor U21914 (N_21914,N_19002,N_19120);
xor U21915 (N_21915,N_19283,N_20925);
nand U21916 (N_21916,N_20883,N_19227);
nor U21917 (N_21917,N_19538,N_21729);
and U21918 (N_21918,N_19358,N_18834);
or U21919 (N_21919,N_20065,N_21441);
xnor U21920 (N_21920,N_21718,N_20042);
xnor U21921 (N_21921,N_21352,N_21454);
or U21922 (N_21922,N_21416,N_20493);
nand U21923 (N_21923,N_19141,N_21231);
or U21924 (N_21924,N_20920,N_21665);
and U21925 (N_21925,N_20261,N_20832);
nor U21926 (N_21926,N_19931,N_19486);
or U21927 (N_21927,N_21255,N_18948);
nor U21928 (N_21928,N_19180,N_20142);
and U21929 (N_21929,N_20685,N_19615);
and U21930 (N_21930,N_21689,N_20160);
or U21931 (N_21931,N_21131,N_19666);
and U21932 (N_21932,N_21601,N_18856);
and U21933 (N_21933,N_21408,N_20820);
or U21934 (N_21934,N_19757,N_20784);
and U21935 (N_21935,N_19610,N_19396);
and U21936 (N_21936,N_20860,N_19453);
nor U21937 (N_21937,N_19166,N_18754);
nand U21938 (N_21938,N_21589,N_21769);
nor U21939 (N_21939,N_21287,N_18833);
and U21940 (N_21940,N_20997,N_19869);
nand U21941 (N_21941,N_19977,N_19592);
nor U21942 (N_21942,N_21590,N_21515);
and U21943 (N_21943,N_20370,N_20366);
nor U21944 (N_21944,N_19548,N_19044);
and U21945 (N_21945,N_19008,N_21006);
nand U21946 (N_21946,N_19984,N_20032);
and U21947 (N_21947,N_18898,N_19297);
and U21948 (N_21948,N_21027,N_18823);
nand U21949 (N_21949,N_20734,N_20642);
nor U21950 (N_21950,N_21099,N_21470);
and U21951 (N_21951,N_20672,N_20283);
nor U21952 (N_21952,N_20797,N_20178);
nand U21953 (N_21953,N_20495,N_19159);
and U21954 (N_21954,N_20840,N_19814);
or U21955 (N_21955,N_20480,N_19327);
nor U21956 (N_21956,N_18764,N_19612);
or U21957 (N_21957,N_20403,N_19355);
xor U21958 (N_21958,N_20474,N_19573);
xor U21959 (N_21959,N_19688,N_21015);
or U21960 (N_21960,N_21760,N_20712);
xnor U21961 (N_21961,N_18879,N_19668);
nor U21962 (N_21962,N_19140,N_21646);
or U21963 (N_21963,N_18950,N_21239);
or U21964 (N_21964,N_20892,N_18973);
xnor U21965 (N_21965,N_21855,N_21652);
nor U21966 (N_21966,N_20164,N_19606);
xor U21967 (N_21967,N_20870,N_20582);
xor U21968 (N_21968,N_18811,N_20700);
xor U21969 (N_21969,N_20950,N_19200);
or U21970 (N_21970,N_20649,N_20946);
or U21971 (N_21971,N_20037,N_19975);
xor U21972 (N_21972,N_20114,N_20043);
nor U21973 (N_21973,N_18835,N_21831);
nor U21974 (N_21974,N_20018,N_18975);
and U21975 (N_21975,N_19412,N_20652);
nor U21976 (N_21976,N_19797,N_21024);
xor U21977 (N_21977,N_21845,N_20522);
xor U21978 (N_21978,N_19378,N_19702);
and U21979 (N_21979,N_20809,N_18809);
and U21980 (N_21980,N_20967,N_18875);
or U21981 (N_21981,N_21253,N_20251);
nand U21982 (N_21982,N_19813,N_19963);
nor U21983 (N_21983,N_20205,N_20187);
and U21984 (N_21984,N_19562,N_19220);
nand U21985 (N_21985,N_19216,N_21840);
nand U21986 (N_21986,N_21355,N_21193);
and U21987 (N_21987,N_19542,N_19081);
and U21988 (N_21988,N_20288,N_20282);
and U21989 (N_21989,N_20262,N_20351);
and U21990 (N_21990,N_20773,N_19543);
and U21991 (N_21991,N_19098,N_20932);
or U21992 (N_21992,N_18935,N_20512);
and U21993 (N_21993,N_18813,N_19475);
or U21994 (N_21994,N_19717,N_19265);
nand U21995 (N_21995,N_18970,N_21750);
nor U21996 (N_21996,N_19085,N_21538);
nor U21997 (N_21997,N_21450,N_21080);
nand U21998 (N_21998,N_21620,N_20449);
nand U21999 (N_21999,N_20496,N_20629);
and U22000 (N_22000,N_20395,N_21474);
nand U22001 (N_22001,N_19272,N_20168);
or U22002 (N_22002,N_21442,N_19071);
or U22003 (N_22003,N_21272,N_21376);
xnor U22004 (N_22004,N_19713,N_20782);
and U22005 (N_22005,N_21838,N_19026);
xor U22006 (N_22006,N_18972,N_18954);
or U22007 (N_22007,N_21622,N_20384);
and U22008 (N_22008,N_18877,N_20003);
nand U22009 (N_22009,N_21326,N_19608);
nand U22010 (N_22010,N_20202,N_19480);
nand U22011 (N_22011,N_21862,N_21354);
nand U22012 (N_22012,N_20772,N_19988);
nor U22013 (N_22013,N_20647,N_19135);
nor U22014 (N_22014,N_21132,N_21499);
or U22015 (N_22015,N_21521,N_19231);
and U22016 (N_22016,N_21864,N_20890);
nand U22017 (N_22017,N_20881,N_21171);
and U22018 (N_22018,N_19215,N_18774);
xor U22019 (N_22019,N_19494,N_20362);
or U22020 (N_22020,N_20115,N_19254);
nand U22021 (N_22021,N_18960,N_21854);
nor U22022 (N_22022,N_20999,N_19059);
xnor U22023 (N_22023,N_19171,N_21714);
and U22024 (N_22024,N_20419,N_21172);
and U22025 (N_22025,N_21502,N_19082);
xnor U22026 (N_22026,N_20668,N_21294);
and U22027 (N_22027,N_20763,N_21090);
nand U22028 (N_22028,N_19518,N_19458);
nand U22029 (N_22029,N_20800,N_20238);
xor U22030 (N_22030,N_21105,N_21215);
xor U22031 (N_22031,N_20451,N_19925);
xor U22032 (N_22032,N_20343,N_20866);
nor U22033 (N_22033,N_18800,N_21835);
nand U22034 (N_22034,N_20492,N_19291);
and U22035 (N_22035,N_21429,N_19448);
or U22036 (N_22036,N_19435,N_19090);
nor U22037 (N_22037,N_19658,N_20225);
or U22038 (N_22038,N_19095,N_21785);
xnor U22039 (N_22039,N_19029,N_21706);
nor U22040 (N_22040,N_19206,N_18989);
or U22041 (N_22041,N_20180,N_21508);
or U22042 (N_22042,N_19398,N_19899);
nand U22043 (N_22043,N_21740,N_18807);
or U22044 (N_22044,N_19174,N_20711);
or U22045 (N_22045,N_20659,N_20898);
nor U22046 (N_22046,N_19182,N_20124);
nand U22047 (N_22047,N_21136,N_19692);
xnor U22048 (N_22048,N_21728,N_21274);
xor U22049 (N_22049,N_18886,N_20356);
and U22050 (N_22050,N_21813,N_21017);
or U22051 (N_22051,N_20688,N_19411);
nor U22052 (N_22052,N_19758,N_20011);
xor U22053 (N_22053,N_19003,N_20686);
or U22054 (N_22054,N_19484,N_19623);
or U22055 (N_22055,N_19835,N_20913);
xor U22056 (N_22056,N_20638,N_19761);
nand U22057 (N_22057,N_21043,N_21378);
or U22058 (N_22058,N_19292,N_19622);
and U22059 (N_22059,N_20783,N_20645);
xnor U22060 (N_22060,N_19995,N_19845);
nor U22061 (N_22061,N_18795,N_19332);
or U22062 (N_22062,N_20031,N_20602);
and U22063 (N_22063,N_20123,N_20905);
and U22064 (N_22064,N_20585,N_20656);
xor U22065 (N_22065,N_21564,N_21459);
or U22066 (N_22066,N_20100,N_21276);
nor U22067 (N_22067,N_18887,N_21501);
and U22068 (N_22068,N_20557,N_21347);
nand U22069 (N_22069,N_21784,N_21368);
and U22070 (N_22070,N_19674,N_21110);
nand U22071 (N_22071,N_18936,N_21517);
or U22072 (N_22072,N_20298,N_19567);
or U22073 (N_22073,N_19466,N_19482);
or U22074 (N_22074,N_21138,N_20744);
nand U22075 (N_22075,N_19418,N_20745);
or U22076 (N_22076,N_20437,N_19338);
xor U22077 (N_22077,N_19205,N_19022);
or U22078 (N_22078,N_21660,N_19062);
nor U22079 (N_22079,N_20604,N_19337);
nor U22080 (N_22080,N_19820,N_18844);
nand U22081 (N_22081,N_21361,N_18915);
nand U22082 (N_22082,N_19894,N_19862);
and U22083 (N_22083,N_19645,N_21561);
nor U22084 (N_22084,N_18995,N_20690);
xnor U22085 (N_22085,N_19444,N_19497);
or U22086 (N_22086,N_18863,N_21505);
nor U22087 (N_22087,N_20367,N_20578);
nand U22088 (N_22088,N_20072,N_20781);
nor U22089 (N_22089,N_20141,N_19744);
or U22090 (N_22090,N_19054,N_18781);
or U22091 (N_22091,N_19756,N_21794);
nor U22092 (N_22092,N_19441,N_20786);
nand U22093 (N_22093,N_20012,N_19724);
and U22094 (N_22094,N_21093,N_20228);
nand U22095 (N_22095,N_21619,N_21270);
or U22096 (N_22096,N_19170,N_20066);
or U22097 (N_22097,N_20731,N_19311);
nor U22098 (N_22098,N_20286,N_19460);
nand U22099 (N_22099,N_21310,N_19052);
xor U22100 (N_22100,N_19787,N_19703);
or U22101 (N_22101,N_18968,N_21039);
xnor U22102 (N_22102,N_19523,N_21316);
nand U22103 (N_22103,N_20850,N_20938);
or U22104 (N_22104,N_21303,N_19936);
and U22105 (N_22105,N_19406,N_21317);
nor U22106 (N_22106,N_21763,N_21325);
and U22107 (N_22107,N_19130,N_18902);
nand U22108 (N_22108,N_21166,N_18914);
or U22109 (N_22109,N_20348,N_19712);
nand U22110 (N_22110,N_19720,N_19604);
or U22111 (N_22111,N_20060,N_21424);
nand U22112 (N_22112,N_21009,N_20607);
or U22113 (N_22113,N_21573,N_20308);
xnor U22114 (N_22114,N_21220,N_20099);
xor U22115 (N_22115,N_20958,N_19155);
and U22116 (N_22116,N_20617,N_20696);
nand U22117 (N_22117,N_21174,N_19055);
xnor U22118 (N_22118,N_21681,N_21673);
and U22119 (N_22119,N_20681,N_20092);
or U22120 (N_22120,N_21440,N_21636);
or U22121 (N_22121,N_21663,N_21307);
or U22122 (N_22122,N_18949,N_21062);
or U22123 (N_22123,N_19509,N_20865);
nor U22124 (N_22124,N_19986,N_18930);
and U22125 (N_22125,N_20992,N_21243);
nand U22126 (N_22126,N_21569,N_20829);
or U22127 (N_22127,N_20603,N_21155);
and U22128 (N_22128,N_21273,N_19873);
or U22129 (N_22129,N_19331,N_20839);
or U22130 (N_22130,N_21106,N_20529);
or U22131 (N_22131,N_19267,N_19815);
nor U22132 (N_22132,N_20955,N_21349);
or U22133 (N_22133,N_20177,N_18852);
or U22134 (N_22134,N_20676,N_21667);
and U22135 (N_22135,N_20498,N_20666);
xnor U22136 (N_22136,N_21758,N_20886);
nor U22137 (N_22137,N_20118,N_21392);
xor U22138 (N_22138,N_19617,N_20837);
nor U22139 (N_22139,N_20363,N_20127);
and U22140 (N_22140,N_21168,N_20424);
and U22141 (N_22141,N_19840,N_20094);
or U22142 (N_22142,N_21338,N_21510);
xnor U22143 (N_22143,N_19909,N_21327);
xnor U22144 (N_22144,N_19763,N_21697);
xor U22145 (N_22145,N_20133,N_19288);
nor U22146 (N_22146,N_20624,N_20713);
or U22147 (N_22147,N_20742,N_21045);
xor U22148 (N_22148,N_19016,N_19990);
nor U22149 (N_22149,N_20143,N_19438);
or U22150 (N_22150,N_21185,N_21853);
nor U22151 (N_22151,N_21603,N_20365);
nor U22152 (N_22152,N_20691,N_19107);
and U22153 (N_22153,N_21135,N_21852);
nor U22154 (N_22154,N_19593,N_20709);
or U22155 (N_22155,N_20338,N_20754);
xor U22156 (N_22156,N_19121,N_20640);
or U22157 (N_22157,N_20942,N_18773);
xnor U22158 (N_22158,N_21001,N_20464);
nor U22159 (N_22159,N_19228,N_19144);
or U22160 (N_22160,N_19529,N_19348);
or U22161 (N_22161,N_20076,N_20211);
or U22162 (N_22162,N_20537,N_21363);
xnor U22163 (N_22163,N_19099,N_19427);
or U22164 (N_22164,N_21716,N_21702);
xnor U22165 (N_22165,N_19179,N_20306);
xor U22166 (N_22166,N_20350,N_21544);
or U22167 (N_22167,N_20488,N_19067);
xnor U22168 (N_22168,N_20015,N_21690);
xor U22169 (N_22169,N_20761,N_21115);
nor U22170 (N_22170,N_20780,N_21382);
and U22171 (N_22171,N_19390,N_21638);
nor U22172 (N_22172,N_21246,N_20923);
xnor U22173 (N_22173,N_19326,N_21358);
nor U22174 (N_22174,N_20132,N_20408);
nand U22175 (N_22175,N_20226,N_19759);
or U22176 (N_22176,N_20316,N_21701);
and U22177 (N_22177,N_21066,N_18880);
xor U22178 (N_22178,N_20867,N_19851);
or U22179 (N_22179,N_19040,N_21183);
nand U22180 (N_22180,N_19580,N_20802);
or U22181 (N_22181,N_21519,N_19006);
and U22182 (N_22182,N_20478,N_20268);
or U22183 (N_22183,N_19321,N_20893);
xnor U22184 (N_22184,N_21318,N_20239);
nand U22185 (N_22185,N_19305,N_21869);
or U22186 (N_22186,N_21822,N_20858);
or U22187 (N_22187,N_20884,N_21114);
and U22188 (N_22188,N_19589,N_20518);
or U22189 (N_22189,N_20441,N_19786);
nand U22190 (N_22190,N_20969,N_21799);
xnor U22191 (N_22191,N_20915,N_20394);
xor U22192 (N_22192,N_19676,N_19690);
nor U22193 (N_22193,N_20399,N_20233);
or U22194 (N_22194,N_21733,N_19245);
nor U22195 (N_22195,N_20000,N_19964);
nor U22196 (N_22196,N_20007,N_20311);
and U22197 (N_22197,N_18923,N_21753);
or U22198 (N_22198,N_19564,N_19613);
nand U22199 (N_22199,N_21288,N_19599);
and U22200 (N_22200,N_20271,N_19657);
and U22201 (N_22201,N_19208,N_20293);
and U22202 (N_22202,N_21731,N_21863);
nor U22203 (N_22203,N_18867,N_21216);
and U22204 (N_22204,N_20790,N_20130);
nand U22205 (N_22205,N_19858,N_21497);
or U22206 (N_22206,N_19609,N_19276);
or U22207 (N_22207,N_19824,N_21471);
or U22208 (N_22208,N_19994,N_19878);
xor U22209 (N_22209,N_19298,N_19591);
and U22210 (N_22210,N_19145,N_20949);
xnor U22211 (N_22211,N_19452,N_20022);
nand U22212 (N_22212,N_21010,N_19353);
xnor U22213 (N_22213,N_21798,N_21577);
or U22214 (N_22214,N_21257,N_20948);
xnor U22215 (N_22215,N_21531,N_19222);
nand U22216 (N_22216,N_20896,N_19571);
nand U22217 (N_22217,N_21371,N_21334);
nor U22218 (N_22218,N_21518,N_21545);
or U22219 (N_22219,N_20004,N_19855);
nor U22220 (N_22220,N_21348,N_19915);
nor U22221 (N_22221,N_19900,N_19684);
xor U22222 (N_22222,N_19100,N_21460);
and U22223 (N_22223,N_19956,N_20423);
xnor U22224 (N_22224,N_21723,N_19036);
nand U22225 (N_22225,N_21195,N_20542);
nand U22226 (N_22226,N_21608,N_20944);
and U22227 (N_22227,N_19508,N_20067);
nor U22228 (N_22228,N_20521,N_19998);
xnor U22229 (N_22229,N_19204,N_21872);
nand U22230 (N_22230,N_20814,N_21268);
or U22231 (N_22231,N_19236,N_19705);
xor U22232 (N_22232,N_21260,N_21643);
xor U22233 (N_22233,N_19264,N_20803);
xnor U22234 (N_22234,N_20392,N_20373);
and U22235 (N_22235,N_18778,N_19675);
nand U22236 (N_22236,N_19117,N_19038);
or U22237 (N_22237,N_21653,N_21801);
or U22238 (N_22238,N_18944,N_20369);
nand U22239 (N_22239,N_19183,N_21439);
nand U22240 (N_22240,N_21411,N_21611);
or U22241 (N_22241,N_18827,N_20903);
or U22242 (N_22242,N_20764,N_21568);
nor U22243 (N_22243,N_19000,N_21679);
and U22244 (N_22244,N_21202,N_19395);
nor U22245 (N_22245,N_21594,N_20794);
nand U22246 (N_22246,N_21205,N_20247);
xnor U22247 (N_22247,N_19957,N_21430);
and U22248 (N_22248,N_20965,N_21005);
nor U22249 (N_22249,N_21744,N_20937);
or U22250 (N_22250,N_21212,N_20325);
nand U22251 (N_22251,N_20220,N_21817);
and U22252 (N_22252,N_21337,N_20033);
and U22253 (N_22253,N_20223,N_19282);
nand U22254 (N_22254,N_21790,N_20064);
xor U22255 (N_22255,N_20834,N_21781);
nand U22256 (N_22256,N_20471,N_19659);
nand U22257 (N_22257,N_21096,N_20219);
nand U22258 (N_22258,N_19974,N_21865);
nor U22259 (N_22259,N_20103,N_19636);
nand U22260 (N_22260,N_18789,N_21369);
nand U22261 (N_22261,N_21719,N_21811);
xor U22262 (N_22262,N_19978,N_20654);
nand U22263 (N_22263,N_20467,N_19747);
nand U22264 (N_22264,N_21383,N_19537);
nand U22265 (N_22265,N_20341,N_20571);
nor U22266 (N_22266,N_18945,N_21776);
xnor U22267 (N_22267,N_19723,N_21063);
and U22268 (N_22268,N_20400,N_21150);
and U22269 (N_22269,N_20976,N_21765);
and U22270 (N_22270,N_21617,N_18772);
nand U22271 (N_22271,N_21026,N_21820);
and U22272 (N_22272,N_20534,N_18775);
and U22273 (N_22273,N_21391,N_19133);
nor U22274 (N_22274,N_20303,N_21175);
xnor U22275 (N_22275,N_19630,N_19914);
nor U22276 (N_22276,N_20145,N_19916);
nand U22277 (N_22277,N_20911,N_19234);
nand U22278 (N_22278,N_19001,N_19825);
or U22279 (N_22279,N_20766,N_20549);
and U22280 (N_22280,N_21446,N_20515);
xor U22281 (N_22281,N_21192,N_21423);
or U22282 (N_22282,N_19483,N_21658);
xor U22283 (N_22283,N_21486,N_19057);
or U22284 (N_22284,N_19652,N_19350);
nor U22285 (N_22285,N_18986,N_20470);
and U22286 (N_22286,N_20572,N_19633);
and U22287 (N_22287,N_21057,N_20090);
and U22288 (N_22288,N_19698,N_21016);
nor U22289 (N_22289,N_20725,N_19760);
or U22290 (N_22290,N_21214,N_19197);
and U22291 (N_22291,N_19695,N_19410);
xnor U22292 (N_22292,N_19437,N_21584);
or U22293 (N_22293,N_21064,N_21842);
and U22294 (N_22294,N_21144,N_20129);
nor U22295 (N_22295,N_20664,N_21217);
and U22296 (N_22296,N_19575,N_18885);
nand U22297 (N_22297,N_21805,N_21693);
and U22298 (N_22298,N_21433,N_19118);
or U22299 (N_22299,N_21311,N_19422);
nor U22300 (N_22300,N_19965,N_20346);
or U22301 (N_22301,N_21049,N_19149);
xor U22302 (N_22302,N_21598,N_19011);
nand U22303 (N_22303,N_20533,N_18984);
nand U22304 (N_22304,N_21251,N_21299);
nor U22305 (N_22305,N_20816,N_20382);
nand U22306 (N_22306,N_19290,N_18907);
or U22307 (N_22307,N_20035,N_21755);
xor U22308 (N_22308,N_19740,N_19469);
and U22309 (N_22309,N_20039,N_19678);
nor U22310 (N_22310,N_20447,N_20564);
xor U22311 (N_22311,N_20391,N_19320);
xnor U22312 (N_22312,N_19046,N_20425);
nor U22313 (N_22313,N_21588,N_20721);
or U22314 (N_22314,N_18974,N_21657);
and U22315 (N_22315,N_21370,N_21803);
nor U22316 (N_22316,N_21301,N_19969);
nor U22317 (N_22317,N_20016,N_18872);
nor U22318 (N_22318,N_18771,N_19745);
or U22319 (N_22319,N_19211,N_20631);
xor U22320 (N_22320,N_21271,N_19999);
and U22321 (N_22321,N_20151,N_21686);
or U22322 (N_22322,N_19876,N_19459);
nor U22323 (N_22323,N_19072,N_19446);
nand U22324 (N_22324,N_19788,N_18874);
or U22325 (N_22325,N_19365,N_20560);
xor U22326 (N_22326,N_21668,N_20815);
and U22327 (N_22327,N_19273,N_19382);
or U22328 (N_22328,N_21621,N_20276);
nor U22329 (N_22329,N_19614,N_20336);
or U22330 (N_22330,N_21154,N_21245);
nor U22331 (N_22331,N_18819,N_20134);
xnor U22332 (N_22332,N_19512,N_21844);
nand U22333 (N_22333,N_19278,N_21397);
or U22334 (N_22334,N_20737,N_19601);
nor U22335 (N_22335,N_20078,N_20588);
nor U22336 (N_22336,N_21042,N_21139);
and U22337 (N_22337,N_19911,N_19867);
or U22338 (N_22338,N_20230,N_19188);
xor U22339 (N_22339,N_21088,N_19201);
or U22340 (N_22340,N_20342,N_20511);
and U22341 (N_22341,N_19158,N_21073);
xnor U22342 (N_22342,N_19126,N_20513);
and U22343 (N_22343,N_20945,N_20086);
or U22344 (N_22344,N_20618,N_21539);
nand U22345 (N_22345,N_19156,N_19341);
and U22346 (N_22346,N_20040,N_20073);
and U22347 (N_22347,N_20215,N_19468);
nor U22348 (N_22348,N_19289,N_20778);
nand U22349 (N_22349,N_21187,N_20344);
nor U22350 (N_22350,N_19104,N_20821);
or U22351 (N_22351,N_20757,N_19304);
xor U22352 (N_22352,N_20577,N_18971);
or U22353 (N_22353,N_20615,N_18925);
nor U22354 (N_22354,N_19701,N_21734);
nand U22355 (N_22355,N_21587,N_21360);
and U22356 (N_22356,N_18921,N_19472);
nand U22357 (N_22357,N_19699,N_20563);
xor U22358 (N_22358,N_20954,N_19269);
and U22359 (N_22359,N_20497,N_20605);
xor U22360 (N_22360,N_19439,N_18871);
or U22361 (N_22361,N_21331,N_20295);
nor U22362 (N_22362,N_18870,N_19249);
xor U22363 (N_22363,N_21036,N_18797);
or U22364 (N_22364,N_20550,N_20875);
nand U22365 (N_22365,N_19018,N_20675);
xor U22366 (N_22366,N_18977,N_19091);
and U22367 (N_22367,N_18840,N_20929);
nand U22368 (N_22368,N_21221,N_19901);
xnor U22369 (N_22369,N_21425,N_20826);
or U22370 (N_22370,N_21341,N_21599);
nand U22371 (N_22371,N_21500,N_21145);
nand U22372 (N_22372,N_20203,N_20673);
nand U22373 (N_22373,N_20789,N_21807);
nand U22374 (N_22374,N_20357,N_21507);
and U22375 (N_22375,N_21453,N_20256);
nand U22376 (N_22376,N_19307,N_20355);
xor U22377 (N_22377,N_20682,N_20185);
and U22378 (N_22378,N_20927,N_19050);
xnor U22379 (N_22379,N_19691,N_19176);
or U22380 (N_22380,N_21340,N_18901);
xnor U22381 (N_22381,N_20987,N_20551);
and U22382 (N_22382,N_21098,N_21445);
or U22383 (N_22383,N_21259,N_19088);
nand U22384 (N_22384,N_19784,N_21548);
xnor U22385 (N_22385,N_21578,N_20989);
xor U22386 (N_22386,N_19579,N_21402);
nand U22387 (N_22387,N_21419,N_20235);
or U22388 (N_22388,N_18919,N_21281);
and U22389 (N_22389,N_20106,N_19810);
nand U22390 (N_22390,N_21530,N_19719);
or U22391 (N_22391,N_20823,N_18927);
or U22392 (N_22392,N_20543,N_19769);
nand U22393 (N_22393,N_19221,N_21727);
xnor U22394 (N_22394,N_19507,N_19019);
or U22395 (N_22395,N_21405,N_19934);
nor U22396 (N_22396,N_20581,N_20573);
and U22397 (N_22397,N_21077,N_20888);
or U22398 (N_22398,N_21680,N_19939);
nand U22399 (N_22399,N_20808,N_20940);
nor U22400 (N_22400,N_19816,N_19037);
or U22401 (N_22401,N_19746,N_20735);
or U22402 (N_22402,N_20095,N_21029);
and U22403 (N_22403,N_19421,N_19162);
or U22404 (N_22404,N_21591,N_19725);
nand U22405 (N_22405,N_19009,N_18905);
nand U22406 (N_22406,N_20538,N_19590);
or U22407 (N_22407,N_21244,N_21642);
and U22408 (N_22408,N_21330,N_20741);
and U22409 (N_22409,N_19146,N_21228);
or U22410 (N_22410,N_20651,N_21580);
nor U22411 (N_22411,N_18782,N_21742);
xnor U22412 (N_22412,N_20270,N_21320);
and U22413 (N_22413,N_21485,N_21103);
or U22414 (N_22414,N_20653,N_21560);
or U22415 (N_22415,N_21596,N_20627);
nor U22416 (N_22416,N_19498,N_18761);
nand U22417 (N_22417,N_19150,N_20706);
xnor U22418 (N_22418,N_21167,N_21533);
nor U22419 (N_22419,N_20836,N_19892);
or U22420 (N_22420,N_21771,N_19499);
nor U22421 (N_22421,N_19479,N_19671);
and U22422 (N_22422,N_20397,N_19917);
xnor U22423 (N_22423,N_18850,N_19033);
and U22424 (N_22424,N_19982,N_21694);
and U22425 (N_22425,N_20152,N_21292);
xnor U22426 (N_22426,N_21449,N_20440);
nor U22427 (N_22427,N_19948,N_21054);
nand U22428 (N_22428,N_20131,N_19286);
nor U22429 (N_22429,N_19677,N_21329);
or U22430 (N_22430,N_20036,N_19329);
nor U22431 (N_22431,N_21373,N_20503);
nand U22432 (N_22432,N_19971,N_20466);
or U22433 (N_22433,N_21528,N_20609);
xnor U22434 (N_22434,N_21495,N_18980);
or U22435 (N_22435,N_18994,N_19041);
and U22436 (N_22436,N_20198,N_20450);
or U22437 (N_22437,N_20885,N_19697);
and U22438 (N_22438,N_19722,N_21431);
nand U22439 (N_22439,N_20980,N_21754);
xor U22440 (N_22440,N_20514,N_19808);
and U22441 (N_22441,N_20393,N_18924);
and U22442 (N_22442,N_19656,N_21607);
or U22443 (N_22443,N_21857,N_21553);
xor U22444 (N_22444,N_19625,N_19487);
or U22445 (N_22445,N_20908,N_20061);
nand U22446 (N_22446,N_20963,N_19449);
nor U22447 (N_22447,N_19315,N_18769);
nor U22448 (N_22448,N_20598,N_20273);
nor U22449 (N_22449,N_21124,N_19983);
xor U22450 (N_22450,N_18983,N_21514);
and U22451 (N_22451,N_20774,N_20359);
or U22452 (N_22452,N_20055,N_19829);
xnor U22453 (N_22453,N_19968,N_21400);
nand U22454 (N_22454,N_19381,N_20637);
nor U22455 (N_22455,N_21775,N_21123);
or U22456 (N_22456,N_18855,N_19535);
nand U22457 (N_22457,N_21597,N_19039);
xor U22458 (N_22458,N_20485,N_19559);
nor U22459 (N_22459,N_18918,N_18829);
nor U22460 (N_22460,N_20396,N_19125);
nor U22461 (N_22461,N_19277,N_20924);
nand U22462 (N_22462,N_21700,N_19568);
nand U22463 (N_22463,N_20859,N_21630);
nand U22464 (N_22464,N_20264,N_19229);
nor U22465 (N_22465,N_20593,N_18987);
xnor U22466 (N_22466,N_20481,N_20779);
xor U22467 (N_22467,N_20096,N_19930);
xnor U22468 (N_22468,N_19577,N_19856);
nor U22469 (N_22469,N_19492,N_20479);
nor U22470 (N_22470,N_21800,N_18831);
and U22471 (N_22471,N_20388,N_19185);
and U22472 (N_22472,N_18903,N_20248);
nor U22473 (N_22473,N_18822,N_21666);
and U22474 (N_22474,N_19413,N_20046);
and U22475 (N_22475,N_20730,N_20760);
and U22476 (N_22476,N_21127,N_20473);
or U22477 (N_22477,N_20953,N_21211);
xnor U22478 (N_22478,N_20345,N_19531);
nand U22479 (N_22479,N_19241,N_19175);
xor U22480 (N_22480,N_20250,N_19795);
and U22481 (N_22481,N_19955,N_19366);
nor U22482 (N_22482,N_19768,N_20935);
nor U22483 (N_22483,N_20476,N_19620);
nor U22484 (N_22484,N_20458,N_19303);
nor U22485 (N_22485,N_21398,N_18865);
xor U22486 (N_22486,N_19848,N_19169);
or U22487 (N_22487,N_20327,N_20726);
xor U22488 (N_22488,N_20995,N_21109);
nand U22489 (N_22489,N_19043,N_19951);
xor U22490 (N_22490,N_19225,N_19013);
and U22491 (N_22491,N_20415,N_21343);
and U22492 (N_22492,N_18912,N_19828);
and U22493 (N_22493,N_21708,N_21705);
nor U22494 (N_22494,N_19445,N_19754);
and U22495 (N_22495,N_21237,N_21041);
nand U22496 (N_22496,N_20045,N_20080);
or U22497 (N_22497,N_19872,N_21258);
xnor U22498 (N_22498,N_21126,N_19384);
nor U22499 (N_22499,N_21802,N_19533);
nor U22500 (N_22500,N_19944,N_21417);
nand U22501 (N_22501,N_20208,N_19981);
and U22502 (N_22502,N_20756,N_19131);
and U22503 (N_22503,N_21462,N_19463);
and U22504 (N_22504,N_20914,N_18934);
nor U22505 (N_22505,N_20714,N_20874);
xnor U22506 (N_22506,N_21833,N_21631);
and U22507 (N_22507,N_21414,N_19728);
xor U22508 (N_22508,N_19912,N_19317);
nand U22509 (N_22509,N_18848,N_20287);
and U22510 (N_22510,N_21284,N_21380);
xnor U22511 (N_22511,N_18888,N_19142);
nand U22512 (N_22512,N_21859,N_20689);
nor U22513 (N_22513,N_20411,N_20200);
nor U22514 (N_22514,N_20213,N_18805);
and U22515 (N_22515,N_19014,N_21484);
xnor U22516 (N_22516,N_20085,N_21224);
and U22517 (N_22517,N_19253,N_20312);
nand U22518 (N_22518,N_20445,N_19086);
or U22519 (N_22519,N_19584,N_19861);
and U22520 (N_22520,N_21759,N_21458);
or U22521 (N_22521,N_19800,N_19101);
nand U22522 (N_22522,N_18893,N_21428);
nand U22523 (N_22523,N_18770,N_19079);
nand U22524 (N_22524,N_19270,N_19884);
or U22525 (N_22525,N_20723,N_21219);
or U22526 (N_22526,N_21791,N_20661);
nor U22527 (N_22527,N_21829,N_20825);
nand U22528 (N_22528,N_20144,N_21238);
xnor U22529 (N_22529,N_20610,N_19866);
and U22530 (N_22530,N_21659,N_19514);
nor U22531 (N_22531,N_18938,N_18799);
xnor U22532 (N_22532,N_19257,N_20959);
and U22533 (N_22533,N_19330,N_21089);
and U22534 (N_22534,N_19476,N_19119);
nor U22535 (N_22535,N_19962,N_19256);
xnor U22536 (N_22536,N_21749,N_19462);
or U22537 (N_22537,N_21682,N_19794);
nand U22538 (N_22538,N_18810,N_19616);
xnor U22539 (N_22539,N_21741,N_19566);
xor U22540 (N_22540,N_20919,N_19987);
or U22541 (N_22541,N_20212,N_21522);
xor U22542 (N_22542,N_19574,N_19230);
nor U22543 (N_22543,N_19997,N_21724);
or U22544 (N_22544,N_19831,N_21020);
xor U22545 (N_22545,N_18779,N_20455);
xnor U22546 (N_22546,N_19252,N_19558);
nand U22547 (N_22547,N_21034,N_20285);
xor U22548 (N_22548,N_20978,N_19064);
nand U22549 (N_22549,N_20161,N_20110);
nor U22550 (N_22550,N_19224,N_20386);
nor U22551 (N_22551,N_18961,N_21023);
or U22552 (N_22552,N_21483,N_21810);
nor U22553 (N_22553,N_19681,N_20758);
or U22554 (N_22554,N_19694,N_19128);
xor U22555 (N_22555,N_20436,N_20221);
xor U22556 (N_22556,N_21672,N_19670);
or U22557 (N_22557,N_21226,N_20302);
nor U22558 (N_22558,N_20921,N_21623);
nand U22559 (N_22559,N_20156,N_20710);
and U22560 (N_22560,N_20260,N_20596);
or U22561 (N_22561,N_18818,N_18801);
nor U22562 (N_22562,N_20680,N_19084);
or U22563 (N_22563,N_21558,N_21674);
and U22564 (N_22564,N_19319,N_19555);
xnor U22565 (N_22565,N_21480,N_18766);
nand U22566 (N_22566,N_20979,N_21830);
nand U22567 (N_22567,N_20991,N_20169);
xnor U22568 (N_22568,N_18787,N_21722);
or U22569 (N_22569,N_20644,N_21277);
and U22570 (N_22570,N_20330,N_19628);
nor U22571 (N_22571,N_19525,N_19882);
or U22572 (N_22572,N_18853,N_21415);
nand U22573 (N_22573,N_18858,N_20722);
nor U22574 (N_22574,N_21335,N_19602);
and U22575 (N_22575,N_19323,N_21362);
xnor U22576 (N_22576,N_19308,N_19165);
xor U22577 (N_22577,N_20136,N_19600);
or U22578 (N_22578,N_21491,N_21834);
nand U22579 (N_22579,N_20404,N_19268);
nor U22580 (N_22580,N_19766,N_20717);
xnor U22581 (N_22581,N_20236,N_19921);
and U22582 (N_22582,N_21639,N_18869);
nor U22583 (N_22583,N_21782,N_19817);
nand U22584 (N_22584,N_21562,N_20590);
or U22585 (N_22585,N_19783,N_20183);
xnor U22586 (N_22586,N_20646,N_21868);
and U22587 (N_22587,N_20738,N_20383);
or U22588 (N_22588,N_19380,N_20243);
xor U22589 (N_22589,N_21332,N_21812);
and U22590 (N_22590,N_19973,N_19877);
nor U22591 (N_22591,N_20417,N_19368);
and U22592 (N_22592,N_21364,N_19918);
nand U22593 (N_22593,N_20352,N_21191);
nor U22594 (N_22594,N_21152,N_20904);
nand U22595 (N_22595,N_20361,N_21448);
xor U22596 (N_22596,N_19027,N_21786);
or U22597 (N_22597,N_21157,N_20528);
nor U22598 (N_22598,N_21605,N_21469);
and U22599 (N_22599,N_18765,N_19827);
nand U22600 (N_22600,N_20289,N_20034);
and U22601 (N_22601,N_18806,N_18836);
or U22602 (N_22602,N_21242,N_21856);
xor U22603 (N_22603,N_21387,N_21060);
xnor U22604 (N_22604,N_19772,N_19993);
or U22605 (N_22605,N_19849,N_20491);
or U22606 (N_22606,N_21604,N_21874);
nand U22607 (N_22607,N_19737,N_21196);
xnor U22608 (N_22608,N_21422,N_20010);
or U22609 (N_22609,N_18862,N_19940);
nor U22610 (N_22610,N_19928,N_19791);
xor U22611 (N_22611,N_20891,N_20209);
nand U22612 (N_22612,N_20234,N_18798);
or U22613 (N_22613,N_20246,N_20029);
or U22614 (N_22614,N_19733,N_19083);
nand U22615 (N_22615,N_20552,N_19597);
nand U22616 (N_22616,N_21633,N_19771);
nor U22617 (N_22617,N_19115,N_21208);
nor U22618 (N_22618,N_20426,N_21761);
nand U22619 (N_22619,N_19068,N_19035);
nor U22620 (N_22620,N_19464,N_19030);
xnor U22621 (N_22621,N_21602,N_20446);
nor U22622 (N_22622,N_19465,N_20048);
and U22623 (N_22623,N_20024,N_21410);
xor U22624 (N_22624,N_20606,N_20683);
and U22625 (N_22625,N_21540,N_21176);
or U22626 (N_22626,N_20930,N_21393);
and U22627 (N_22627,N_21033,N_19106);
nor U22628 (N_22628,N_19357,N_19686);
or U22629 (N_22629,N_21600,N_19143);
nor U22630 (N_22630,N_21647,N_18958);
or U22631 (N_22631,N_19474,N_21496);
nor U22632 (N_22632,N_19721,N_19715);
nand U22633 (N_22633,N_21432,N_20912);
xor U22634 (N_22634,N_19351,N_19496);
nor U22635 (N_22635,N_18899,N_20854);
and U22636 (N_22636,N_19193,N_21523);
nand U22637 (N_22637,N_19242,N_19328);
and U22638 (N_22638,N_21752,N_20665);
or U22639 (N_22639,N_20297,N_18981);
nor U22640 (N_22640,N_21186,N_21789);
or U22641 (N_22641,N_18941,N_18966);
nor U22642 (N_22642,N_19748,N_18931);
nor U22643 (N_22643,N_21873,N_20547);
nand U22644 (N_22644,N_18965,N_19870);
xor U22645 (N_22645,N_21476,N_18964);
nor U22646 (N_22646,N_19935,N_19284);
nand U22647 (N_22647,N_20998,N_20292);
nor U22648 (N_22648,N_21025,N_19399);
nand U22649 (N_22649,N_21404,N_20452);
nor U22650 (N_22650,N_20849,N_19387);
nor U22651 (N_22651,N_20138,N_21858);
nand U22652 (N_22652,N_21056,N_19151);
and U22653 (N_22653,N_20313,N_19556);
or U22654 (N_22654,N_20379,N_21262);
and U22655 (N_22655,N_21308,N_21764);
nor U22656 (N_22656,N_21336,N_21222);
nor U22657 (N_22657,N_20216,N_19891);
xor U22658 (N_22658,N_20591,N_20833);
xor U22659 (N_22659,N_21182,N_20822);
xnor U22660 (N_22660,N_21366,N_21204);
or U22661 (N_22661,N_21563,N_19897);
nor U22662 (N_22662,N_21223,N_21457);
nand U22663 (N_22663,N_19306,N_20354);
nand U22664 (N_22664,N_20102,N_19432);
or U22665 (N_22665,N_20962,N_20684);
nor U22666 (N_22666,N_20318,N_19941);
xnor U22667 (N_22667,N_19223,N_19377);
xor U22668 (N_22668,N_19520,N_21149);
or U22669 (N_22669,N_19910,N_19793);
nor U22670 (N_22670,N_20056,N_21418);
or U22671 (N_22671,N_19051,N_19818);
and U22672 (N_22672,N_21703,N_20329);
and U22673 (N_22673,N_21575,N_21654);
nand U22674 (N_22674,N_20013,N_19889);
nand U22675 (N_22675,N_21685,N_21493);
and U22676 (N_22676,N_19683,N_20107);
and U22677 (N_22677,N_21158,N_20444);
nand U22678 (N_22678,N_19426,N_20299);
nor U22679 (N_22679,N_19513,N_21451);
and U22680 (N_22680,N_19139,N_21467);
and U22681 (N_22681,N_21032,N_20193);
or U22682 (N_22682,N_19619,N_20678);
or U22683 (N_22683,N_21197,N_19552);
or U22684 (N_22684,N_20951,N_21836);
xnor U22685 (N_22685,N_18808,N_19360);
nand U22686 (N_22686,N_21319,N_21489);
nor U22687 (N_22687,N_21372,N_20494);
xnor U22688 (N_22688,N_19585,N_19425);
and U22689 (N_22689,N_20254,N_19154);
nor U22690 (N_22690,N_21128,N_18895);
nor U22691 (N_22691,N_20856,N_20788);
nor U22692 (N_22692,N_21200,N_20290);
nor U22693 (N_22693,N_20641,N_20835);
xor U22694 (N_22694,N_20845,N_21641);
nand U22695 (N_22695,N_18952,N_21823);
nand U22696 (N_22696,N_19203,N_18917);
nor U22697 (N_22697,N_21846,N_20448);
or U22698 (N_22698,N_21021,N_20994);
nand U22699 (N_22699,N_21012,N_20432);
and U22700 (N_22700,N_19386,N_19565);
xor U22701 (N_22701,N_21488,N_18884);
nor U22702 (N_22702,N_21267,N_21143);
or U22703 (N_22703,N_20842,N_18904);
nand U22704 (N_22704,N_21841,N_20047);
xor U22705 (N_22705,N_19979,N_19875);
xnor U22706 (N_22706,N_21711,N_18768);
nand U22707 (N_22707,N_19922,N_20755);
nand U22708 (N_22708,N_18849,N_20277);
nand U22709 (N_22709,N_21111,N_20694);
xor U22710 (N_22710,N_20873,N_21091);
nand U22711 (N_22711,N_18763,N_18760);
xnor U22712 (N_22712,N_20407,N_18817);
xor U22713 (N_22713,N_20526,N_20807);
or U22714 (N_22714,N_20483,N_19087);
xor U22715 (N_22715,N_18990,N_19433);
nor U22716 (N_22716,N_19454,N_20846);
or U22717 (N_22717,N_20634,N_21511);
or U22718 (N_22718,N_20791,N_20939);
xor U22719 (N_22719,N_21121,N_19501);
and U22720 (N_22720,N_20674,N_20252);
and U22721 (N_22721,N_21464,N_20687);
xnor U22722 (N_22722,N_21720,N_19883);
and U22723 (N_22723,N_20698,N_19526);
xnor U22724 (N_22724,N_19904,N_21537);
and U22725 (N_22725,N_21297,N_19473);
nand U22726 (N_22726,N_21210,N_19163);
nor U22727 (N_22727,N_19682,N_20378);
and U22728 (N_22728,N_21847,N_18997);
and U22729 (N_22729,N_19594,N_20633);
or U22730 (N_22730,N_20677,N_19248);
nor U22731 (N_22731,N_19516,N_20824);
nor U22732 (N_22732,N_19363,N_19076);
nand U22733 (N_22733,N_18953,N_20984);
and U22734 (N_22734,N_21804,N_19545);
nor U22735 (N_22735,N_20746,N_21295);
and U22736 (N_22736,N_21048,N_20434);
and U22737 (N_22737,N_19685,N_19226);
or U22738 (N_22738,N_20576,N_21850);
or U22739 (N_22739,N_19976,N_19031);
nor U22740 (N_22740,N_21768,N_19369);
or U22741 (N_22741,N_20291,N_19885);
or U22742 (N_22742,N_18940,N_21848);
xor U22743 (N_22743,N_20643,N_20799);
and U22744 (N_22744,N_20828,N_20907);
nor U22745 (N_22745,N_19611,N_19644);
or U22746 (N_22746,N_21456,N_21198);
nor U22747 (N_22747,N_18933,N_21443);
nor U22748 (N_22748,N_19335,N_20162);
xnor U22749 (N_22749,N_21028,N_20507);
and U22750 (N_22750,N_19239,N_19826);
nor U22751 (N_22751,N_19544,N_19097);
or U22752 (N_22752,N_19196,N_21826);
or U22753 (N_22753,N_19765,N_20098);
nor U22754 (N_22754,N_21407,N_19629);
nor U22755 (N_22755,N_21122,N_18866);
and U22756 (N_22756,N_20539,N_21095);
and U22757 (N_22757,N_19436,N_20520);
nand U22758 (N_22758,N_19605,N_19669);
or U22759 (N_22759,N_19734,N_21133);
and U22760 (N_22760,N_20559,N_20294);
or U22761 (N_22761,N_21777,N_21618);
nor U22762 (N_22762,N_20469,N_18991);
or U22763 (N_22763,N_19553,N_19481);
nor U22764 (N_22764,N_20320,N_20611);
nand U22765 (N_22765,N_20190,N_20505);
nand U22766 (N_22766,N_21367,N_21233);
nand U22767 (N_22767,N_21444,N_21675);
and U22768 (N_22768,N_18860,N_20020);
nand U22769 (N_22769,N_20541,N_19679);
xor U22770 (N_22770,N_20635,N_20420);
nor U22771 (N_22771,N_21160,N_20724);
xnor U22772 (N_22772,N_20189,N_20410);
or U22773 (N_22773,N_20304,N_18883);
and U22774 (N_22774,N_19325,N_21290);
xor U22775 (N_22775,N_21394,N_19343);
or U22776 (N_22776,N_21766,N_20113);
or U22777 (N_22777,N_19822,N_19727);
nand U22778 (N_22778,N_21635,N_19680);
and U22779 (N_22779,N_21490,N_19662);
nand U22780 (N_22780,N_19524,N_20993);
or U22781 (N_22781,N_19932,N_21112);
nor U22782 (N_22782,N_21792,N_21465);
nand U22783 (N_22783,N_19650,N_21130);
nand U22784 (N_22784,N_19926,N_21717);
or U22785 (N_22785,N_20504,N_18876);
or U22786 (N_22786,N_21676,N_20918);
nor U22787 (N_22787,N_18784,N_19312);
xnor U22788 (N_22788,N_20154,N_20589);
nor U22789 (N_22789,N_19530,N_20428);
nand U22790 (N_22790,N_21181,N_20628);
xnor U22791 (N_22791,N_20305,N_21498);
xnor U22792 (N_22792,N_21055,N_21699);
nand U22793 (N_22793,N_19843,N_20567);
nand U22794 (N_22794,N_21293,N_19880);
xor U22795 (N_22795,N_20412,N_21256);
nor U22796 (N_22796,N_19839,N_21532);
and U22797 (N_22797,N_20715,N_21615);
nand U22798 (N_22798,N_21207,N_19563);
and U22799 (N_22799,N_21344,N_20128);
nor U22800 (N_22800,N_19134,N_19989);
xor U22801 (N_22801,N_20140,N_19522);
and U22802 (N_22802,N_19711,N_20852);
xor U22803 (N_22803,N_19255,N_19275);
or U22804 (N_22804,N_19202,N_19495);
or U22805 (N_22805,N_19547,N_19356);
nor U22806 (N_22806,N_19812,N_19710);
or U22807 (N_22807,N_21559,N_21169);
and U22808 (N_22808,N_21565,N_20838);
and U22809 (N_22809,N_19923,N_19434);
xnor U22810 (N_22810,N_19785,N_21556);
nor U22811 (N_22811,N_21570,N_20402);
xnor U22812 (N_22812,N_20433,N_19896);
or U22813 (N_22813,N_21747,N_19132);
nor U22814 (N_22814,N_20053,N_20360);
or U22815 (N_22815,N_21304,N_20019);
nand U22816 (N_22816,N_20910,N_19942);
or U22817 (N_22817,N_19913,N_19376);
and U22818 (N_22818,N_21542,N_20229);
nor U22819 (N_22819,N_21071,N_21525);
xnor U22820 (N_22820,N_19285,N_20957);
xor U22821 (N_22821,N_20207,N_21194);
xor U22822 (N_22822,N_18890,N_21796);
nand U22823 (N_22823,N_20767,N_19178);
nand U22824 (N_22824,N_19034,N_21866);
and U22825 (N_22825,N_20347,N_20805);
and U22826 (N_22826,N_20184,N_20882);
nand U22827 (N_22827,N_21730,N_21094);
xor U22828 (N_22828,N_20575,N_21839);
or U22829 (N_22829,N_20535,N_21815);
nand U22830 (N_22830,N_20812,N_20851);
xnor U22831 (N_22831,N_21828,N_19578);
and U22832 (N_22832,N_20322,N_19238);
nand U22833 (N_22833,N_20204,N_20599);
and U22834 (N_22834,N_21821,N_18803);
or U22835 (N_22835,N_18794,N_18792);
xnor U22836 (N_22836,N_20558,N_19112);
xnor U22837 (N_22837,N_20122,N_20798);
nand U22838 (N_22838,N_21264,N_18894);
nor U22839 (N_22839,N_21018,N_20759);
or U22840 (N_22840,N_18857,N_19233);
and U22841 (N_22841,N_19214,N_19635);
xnor U22842 (N_22842,N_19314,N_20983);
nand U22843 (N_22843,N_19042,N_20197);
nand U22844 (N_22844,N_21662,N_19021);
nor U22845 (N_22845,N_21140,N_20255);
xor U22846 (N_22846,N_19025,N_20224);
and U22847 (N_22847,N_21546,N_21151);
nor U22848 (N_22848,N_20620,N_21626);
and U22849 (N_22849,N_19024,N_19408);
or U22850 (N_22850,N_20818,N_20083);
or U22851 (N_22851,N_19693,N_20191);
or U22852 (N_22852,N_20880,N_20317);
nand U22853 (N_22853,N_20565,N_20429);
nor U22854 (N_22854,N_19888,N_20732);
nand U22855 (N_22855,N_21632,N_20727);
and U22856 (N_22856,N_18955,N_21778);
xnor U22857 (N_22857,N_20960,N_20853);
xor U22858 (N_22858,N_21019,N_20695);
xor U22859 (N_22859,N_19854,N_18878);
xnor U22860 (N_22860,N_18791,N_19667);
or U22861 (N_22861,N_20941,N_20974);
xnor U22862 (N_22862,N_19991,N_21494);
xnor U22863 (N_22863,N_20314,N_19587);
nand U22864 (N_22864,N_21153,N_20516);
xnor U22865 (N_22865,N_20630,N_21644);
or U22866 (N_22866,N_19844,N_20014);
nor U22867 (N_22867,N_20961,N_21579);
nand U22868 (N_22868,N_19649,N_20971);
nand U22869 (N_22869,N_19004,N_19687);
nor U22870 (N_22870,N_18790,N_18832);
and U22871 (N_22871,N_20227,N_19945);
and U22872 (N_22872,N_20387,N_20409);
and U22873 (N_22873,N_20489,N_19346);
nand U22874 (N_22874,N_20827,N_20101);
nand U22875 (N_22875,N_19251,N_18812);
nor U22876 (N_22876,N_19581,N_20601);
or U22877 (N_22877,N_19527,N_18767);
nand U22878 (N_22878,N_19280,N_21566);
nor U22879 (N_22879,N_20087,N_19726);
nand U22880 (N_22880,N_20922,N_19992);
nor U22881 (N_22881,N_19168,N_20240);
nand U22882 (N_22882,N_20021,N_19490);
xnor U22883 (N_22883,N_19177,N_19259);
nor U22884 (N_22884,N_18837,N_20975);
nand U22885 (N_22885,N_20871,N_19972);
and U22886 (N_22886,N_19738,N_21235);
and U22887 (N_22887,N_21285,N_21342);
nand U22888 (N_22888,N_21861,N_21762);
xor U22889 (N_22889,N_18892,N_21100);
nand U22890 (N_22890,N_19540,N_19792);
and U22891 (N_22891,N_19198,N_19261);
nor U22892 (N_22892,N_21592,N_21683);
nand U22893 (N_22893,N_21477,N_21134);
and U22894 (N_22894,N_20150,N_20139);
or U22895 (N_22895,N_19640,N_21283);
and U22896 (N_22896,N_19696,N_21616);
or U22897 (N_22897,N_21388,N_21586);
nand U22898 (N_22898,N_21333,N_19393);
xnor U22899 (N_22899,N_18967,N_20218);
nor U22900 (N_22900,N_20192,N_19572);
nor U22901 (N_22901,N_21593,N_19874);
and U22902 (N_22902,N_20091,N_19503);
nand U22903 (N_22903,N_20662,N_19313);
nand U22904 (N_22904,N_18982,N_19536);
nor U22905 (N_22905,N_19778,N_19207);
or U22906 (N_22906,N_20005,N_19266);
or U22907 (N_22907,N_19789,N_19423);
nor U22908 (N_22908,N_19905,N_20422);
and U22909 (N_22909,N_21381,N_21084);
and U22910 (N_22910,N_20718,N_19372);
nand U22911 (N_22911,N_19077,N_21624);
nor U22912 (N_22912,N_19706,N_21481);
xor U22913 (N_22913,N_21291,N_20508);
and U22914 (N_22914,N_21479,N_20670);
or U22915 (N_22915,N_20697,N_19309);
nand U22916 (N_22916,N_20263,N_20237);
xnor U22917 (N_22917,N_20517,N_21252);
or U22918 (N_22918,N_19554,N_20331);
or U22919 (N_22919,N_18998,N_19927);
nor U22920 (N_22920,N_18882,N_19430);
nor U22921 (N_22921,N_19672,N_19576);
or U22922 (N_22922,N_19852,N_21691);
or U22923 (N_22923,N_20349,N_20819);
nand U22924 (N_22924,N_20222,N_19489);
nor U22925 (N_22925,N_21086,N_19502);
xor U22926 (N_22926,N_21052,N_20728);
or U22927 (N_22927,N_20750,N_21773);
or U22928 (N_22928,N_20199,N_21713);
or U22929 (N_22929,N_19819,N_19504);
nand U22930 (N_22930,N_19354,N_21738);
nand U22931 (N_22931,N_20749,N_20956);
and U22932 (N_22932,N_19428,N_19510);
xnor U22933 (N_22933,N_19618,N_19416);
nand U22934 (N_22934,N_20171,N_19595);
xnor U22935 (N_22935,N_19279,N_19103);
nand U22936 (N_22936,N_20594,N_20506);
or U22937 (N_22937,N_20002,N_21230);
xnor U22938 (N_22938,N_21743,N_18906);
and U22939 (N_22939,N_19823,N_20241);
or U22940 (N_22940,N_21707,N_20050);
and U22941 (N_22941,N_21038,N_19191);
nand U22942 (N_22942,N_21309,N_20527);
and U22943 (N_22943,N_20579,N_20206);
nor U22944 (N_22944,N_21022,N_20301);
or U22945 (N_22945,N_20059,N_20702);
xor U22946 (N_22946,N_21058,N_19641);
xor U22947 (N_22947,N_19352,N_19801);
nand U22948 (N_22948,N_21137,N_21737);
nand U22949 (N_22949,N_21087,N_21612);
nand U22950 (N_22950,N_19846,N_20947);
xor U22951 (N_22951,N_21102,N_21473);
nand U22952 (N_22952,N_21298,N_21656);
xor U22953 (N_22953,N_20583,N_19316);
nor U22954 (N_22954,N_19424,N_21770);
xnor U22955 (N_22955,N_21116,N_18780);
nand U22956 (N_22956,N_21403,N_19798);
and U22957 (N_22957,N_19294,N_19731);
and U22958 (N_22958,N_19075,N_18996);
nand U22959 (N_22959,N_20281,N_19089);
nor U22960 (N_22960,N_20081,N_19919);
xor U22961 (N_22961,N_20044,N_21232);
nand U22962 (N_22962,N_19751,N_19953);
or U22963 (N_22963,N_21218,N_21606);
nor U22964 (N_22964,N_20524,N_19184);
nand U22965 (N_22965,N_19405,N_18752);
or U22966 (N_22966,N_19073,N_20051);
nor U22967 (N_22967,N_21314,N_20307);
and U22968 (N_22968,N_21011,N_19603);
nand U22969 (N_22969,N_21050,N_21390);
xnor U22970 (N_22970,N_19943,N_18830);
nand U22971 (N_22971,N_21552,N_20736);
xor U22972 (N_22972,N_18978,N_20796);
and U22973 (N_22973,N_19160,N_20545);
or U22974 (N_22974,N_21543,N_18785);
nand U22975 (N_22975,N_20519,N_18947);
or U22976 (N_22976,N_21188,N_21669);
nor U22977 (N_22977,N_21640,N_19392);
or U22978 (N_22978,N_21125,N_20179);
nand U22979 (N_22979,N_20751,N_21044);
nand U22980 (N_22980,N_21227,N_19646);
xor U22981 (N_22981,N_18942,N_19634);
or U22982 (N_22982,N_20049,N_21053);
and U22983 (N_22983,N_20663,N_21628);
nor U22984 (N_22984,N_20372,N_19367);
xnor U22985 (N_22985,N_19781,N_21613);
or U22986 (N_22986,N_21827,N_21148);
and U22987 (N_22987,N_19648,N_19790);
and U22988 (N_22988,N_20600,N_20088);
nor U22989 (N_22989,N_20900,N_20174);
nor U22990 (N_22990,N_19643,N_21322);
xnor U22991 (N_22991,N_19950,N_21413);
xor U22992 (N_22992,N_20848,N_18750);
nand U22993 (N_22993,N_19045,N_21455);
nor U22994 (N_22994,N_21651,N_20509);
nor U22995 (N_22995,N_19333,N_21070);
nand U22996 (N_22996,N_19404,N_20421);
or U22997 (N_22997,N_21082,N_19549);
nor U22998 (N_22998,N_19517,N_20499);
xor U22999 (N_22999,N_20380,N_20972);
xnor U23000 (N_23000,N_18900,N_19244);
or U23001 (N_23001,N_19732,N_20878);
or U23002 (N_23002,N_18943,N_21648);
and U23003 (N_23003,N_21808,N_19906);
nand U23004 (N_23004,N_21108,N_19937);
nand U23005 (N_23005,N_19864,N_18920);
xnor U23006 (N_23006,N_21512,N_19802);
xor U23007 (N_23007,N_19924,N_19127);
and U23008 (N_23008,N_20546,N_21250);
nand U23009 (N_23009,N_19020,N_20990);
or U23010 (N_23010,N_19388,N_20895);
or U23011 (N_23011,N_21634,N_20077);
nor U23012 (N_23012,N_19638,N_20770);
xor U23013 (N_23013,N_19739,N_19336);
nor U23014 (N_23014,N_19340,N_19060);
and U23015 (N_23015,N_20242,N_21797);
and U23016 (N_23016,N_21101,N_18861);
nand U23017 (N_23017,N_20300,N_18762);
and U23018 (N_23018,N_20795,N_19952);
and U23019 (N_23019,N_19383,N_19596);
and U23020 (N_23020,N_20165,N_20743);
or U23021 (N_23021,N_19385,N_19032);
and U23022 (N_23022,N_20074,N_20655);
nor U23023 (N_23023,N_20707,N_21265);
or U23024 (N_23024,N_18816,N_18815);
or U23025 (N_23025,N_18851,N_21783);
xor U23026 (N_23026,N_20792,N_21468);
nor U23027 (N_23027,N_20465,N_19246);
nor U23028 (N_23028,N_21206,N_19859);
and U23029 (N_23029,N_19167,N_18838);
and U23030 (N_23030,N_19887,N_20093);
nand U23031 (N_23031,N_21526,N_21013);
or U23032 (N_23032,N_18847,N_21240);
xor U23033 (N_23033,N_19250,N_20510);
and U23034 (N_23034,N_21710,N_19541);
nand U23035 (N_23035,N_20339,N_19070);
and U23036 (N_23036,N_21165,N_21147);
or U23037 (N_23037,N_19511,N_19799);
nor U23038 (N_23038,N_21704,N_21780);
or U23039 (N_23039,N_20916,N_21779);
nand U23040 (N_23040,N_19344,N_18929);
or U23041 (N_23041,N_21581,N_21002);
nor U23042 (N_23042,N_20787,N_19028);
and U23043 (N_23043,N_19470,N_20137);
and U23044 (N_23044,N_19195,N_20001);
xnor U23045 (N_23045,N_21065,N_19379);
or U23046 (N_23046,N_20562,N_20768);
nand U23047 (N_23047,N_19966,N_21159);
nand U23048 (N_23048,N_21356,N_19857);
and U23049 (N_23049,N_21870,N_21809);
nor U23050 (N_23050,N_21492,N_20806);
and U23051 (N_23051,N_19716,N_21574);
xor U23052 (N_23052,N_19639,N_21475);
and U23053 (N_23053,N_18783,N_19519);
and U23054 (N_23054,N_21554,N_18896);
nand U23055 (N_23055,N_19651,N_19061);
nor U23056 (N_23056,N_19933,N_21795);
and U23057 (N_23057,N_19053,N_20748);
or U23058 (N_23058,N_19457,N_19663);
or U23059 (N_23059,N_18932,N_21421);
nand U23060 (N_23060,N_19109,N_20332);
or U23061 (N_23061,N_20041,N_18913);
nor U23062 (N_23062,N_19153,N_21300);
nor U23063 (N_23063,N_19074,N_20708);
nand U23064 (N_23064,N_21739,N_19443);
nand U23065 (N_23065,N_18802,N_19583);
nand U23066 (N_23066,N_19210,N_20027);
nand U23067 (N_23067,N_20389,N_20453);
and U23068 (N_23068,N_21254,N_18804);
nor U23069 (N_23069,N_20623,N_19114);
or U23070 (N_23070,N_20621,N_20720);
nand U23071 (N_23071,N_21547,N_19841);
nand U23072 (N_23072,N_20030,N_18826);
nor U23073 (N_23073,N_19569,N_19301);
or U23074 (N_23074,N_20253,N_19322);
nor U23075 (N_23075,N_19157,N_21557);
nand U23076 (N_23076,N_20333,N_21756);
nor U23077 (N_23077,N_18993,N_19124);
and U23078 (N_23078,N_21280,N_21767);
or U23079 (N_23079,N_21353,N_21712);
nor U23080 (N_23080,N_21572,N_20009);
nand U23081 (N_23081,N_20375,N_20195);
and U23082 (N_23082,N_21209,N_18842);
xnor U23083 (N_23083,N_21083,N_19108);
nor U23084 (N_23084,N_20769,N_19274);
xnor U23085 (N_23085,N_20973,N_20194);
or U23086 (N_23086,N_20747,N_20597);
or U23087 (N_23087,N_20158,N_19550);
xnor U23088 (N_23088,N_20864,N_19895);
or U23089 (N_23089,N_18937,N_19830);
and U23090 (N_23090,N_19349,N_19561);
nor U23091 (N_23091,N_21203,N_21118);
and U23092 (N_23092,N_20671,N_20456);
or U23093 (N_23093,N_21871,N_21031);
nand U23094 (N_23094,N_21466,N_19491);
and U23095 (N_23095,N_21007,N_19295);
nand U23096 (N_23096,N_21076,N_19776);
and U23097 (N_23097,N_21583,N_19532);
and U23098 (N_23098,N_20897,N_20926);
and U23099 (N_23099,N_19586,N_21437);
or U23100 (N_23100,N_19805,N_19881);
nor U23101 (N_23101,N_20804,N_20210);
nand U23102 (N_23102,N_21609,N_20071);
and U23103 (N_23103,N_20385,N_19359);
xor U23104 (N_23104,N_19389,N_20406);
nand U23105 (N_23105,N_20532,N_20876);
nor U23106 (N_23106,N_20894,N_21339);
and U23107 (N_23107,N_21003,N_20705);
xor U23108 (N_23108,N_21819,N_21851);
and U23109 (N_23109,N_20459,N_19929);
or U23110 (N_23110,N_21726,N_21867);
or U23111 (N_23111,N_21357,N_19467);
and U23112 (N_23112,N_20069,N_20887);
and U23113 (N_23113,N_21696,N_21793);
or U23114 (N_23114,N_20266,N_21040);
xor U23115 (N_23115,N_21506,N_21345);
xor U23116 (N_23116,N_21113,N_20977);
nor U23117 (N_23117,N_19626,N_21396);
xnor U23118 (N_23118,N_18776,N_19908);
and U23119 (N_23119,N_19370,N_19102);
nand U23120 (N_23120,N_21328,N_19219);
nor U23121 (N_23121,N_19661,N_18908);
nor U23122 (N_23122,N_19809,N_19938);
and U23123 (N_23123,N_20126,N_20201);
nor U23124 (N_23124,N_20232,N_21037);
or U23125 (N_23125,N_19607,N_21386);
nand U23126 (N_23126,N_21164,N_21241);
or U23127 (N_23127,N_20265,N_20667);
nand U23128 (N_23128,N_20739,N_21849);
and U23129 (N_23129,N_19551,N_18969);
xnor U23130 (N_23130,N_21129,N_20063);
nor U23131 (N_23131,N_21315,N_19419);
nor U23132 (N_23132,N_21085,N_20468);
xor U23133 (N_23133,N_19409,N_19960);
nor U23134 (N_23134,N_20692,N_21395);
nand U23135 (N_23135,N_19069,N_19774);
and U23136 (N_23136,N_18755,N_20414);
and U23137 (N_23137,N_19111,N_18859);
or U23138 (N_23138,N_20062,N_21236);
or U23139 (N_23139,N_20548,N_20462);
or U23140 (N_23140,N_21346,N_21535);
or U23141 (N_23141,N_21837,N_20120);
or U23142 (N_23142,N_19263,N_20148);
or U23143 (N_23143,N_21595,N_20928);
xnor U23144 (N_23144,N_18788,N_19164);
or U23145 (N_23145,N_19010,N_19023);
nor U23146 (N_23146,N_18777,N_20595);
or U23147 (N_23147,N_19373,N_20701);
nand U23148 (N_23148,N_20335,N_18992);
or U23149 (N_23149,N_21234,N_20275);
nor U23150 (N_23150,N_19842,N_21173);
and U23151 (N_23151,N_20525,N_19736);
and U23152 (N_23152,N_21736,N_20438);
nand U23153 (N_23153,N_19735,N_21671);
xnor U23154 (N_23154,N_21732,N_20570);
xor U23155 (N_23155,N_21097,N_19980);
and U23156 (N_23156,N_20693,N_21536);
nand U23157 (N_23157,N_21438,N_18939);
or U23158 (N_23158,N_21625,N_20172);
nand U23159 (N_23159,N_19886,N_19105);
nand U23160 (N_23160,N_20324,N_20181);
and U23161 (N_23161,N_19506,N_20986);
and U23162 (N_23162,N_20337,N_21286);
or U23163 (N_23163,N_21289,N_19500);
and U23164 (N_23164,N_19361,N_20401);
nor U23165 (N_23165,N_19515,N_21745);
nand U23166 (N_23166,N_20188,N_20267);
nand U23167 (N_23167,N_19521,N_20817);
nor U23168 (N_23168,N_19414,N_20319);
nand U23169 (N_23169,N_20112,N_21661);
xnor U23170 (N_23170,N_20374,N_19047);
and U23171 (N_23171,N_20368,N_21482);
or U23172 (N_23172,N_21504,N_20906);
nor U23173 (N_23173,N_21104,N_19570);
and U23174 (N_23174,N_21688,N_19907);
nor U23175 (N_23175,N_20556,N_20416);
or U23176 (N_23176,N_20966,N_19879);
xor U23177 (N_23177,N_20917,N_19334);
nor U23178 (N_23178,N_20070,N_20762);
nor U23179 (N_23179,N_19890,N_20245);
or U23180 (N_23180,N_19420,N_21527);
xnor U23181 (N_23181,N_19588,N_21435);
xor U23182 (N_23182,N_19078,N_21177);
nor U23183 (N_23183,N_19407,N_21843);
nor U23184 (N_23184,N_21161,N_20869);
or U23185 (N_23185,N_20109,N_20901);
or U23186 (N_23186,N_19750,N_21278);
nand U23187 (N_23187,N_20801,N_21585);
nand U23188 (N_23188,N_19362,N_21427);
nand U23189 (N_23189,N_20530,N_18820);
xor U23190 (N_23190,N_21305,N_21788);
and U23191 (N_23191,N_20776,N_18881);
nand U23192 (N_23192,N_20889,N_21627);
and U23193 (N_23193,N_19811,N_19478);
and U23194 (N_23194,N_21772,N_21629);
nor U23195 (N_23195,N_20523,N_20487);
nand U23196 (N_23196,N_19708,N_19450);
nand U23197 (N_23197,N_19755,N_21567);
or U23198 (N_23198,N_20381,N_18959);
xor U23199 (N_23199,N_19138,N_21610);
nand U23200 (N_23200,N_19477,N_21555);
nor U23201 (N_23201,N_19429,N_19749);
or U23202 (N_23202,N_21075,N_21275);
nand U23203 (N_23203,N_20052,N_21529);
nand U23204 (N_23204,N_20371,N_18854);
nor U23205 (N_23205,N_19240,N_21225);
nor U23206 (N_23206,N_19833,N_19339);
xnor U23207 (N_23207,N_19947,N_21541);
nand U23208 (N_23208,N_19456,N_21650);
xnor U23209 (N_23209,N_21119,N_21030);
and U23210 (N_23210,N_20439,N_20079);
or U23211 (N_23211,N_19137,N_20149);
nor U23212 (N_23212,N_18753,N_20461);
and U23213 (N_23213,N_19302,N_20413);
nor U23214 (N_23214,N_18951,N_21213);
and U23215 (N_23215,N_20068,N_19631);
nor U23216 (N_23216,N_19065,N_20813);
and U23217 (N_23217,N_20587,N_19094);
nor U23218 (N_23218,N_21860,N_21068);
nor U23219 (N_23219,N_19324,N_19832);
xnor U23220 (N_23220,N_20785,N_20490);
and U23221 (N_23221,N_19310,N_21313);
nand U23222 (N_23222,N_20855,N_20310);
or U23223 (N_23223,N_20777,N_18926);
or U23224 (N_23224,N_19080,N_18756);
nor U23225 (N_23225,N_20054,N_20364);
xor U23226 (N_23226,N_19402,N_19959);
xor U23227 (N_23227,N_20484,N_20340);
nand U23228 (N_23228,N_19534,N_19199);
xnor U23229 (N_23229,N_19123,N_19624);
nand U23230 (N_23230,N_19213,N_21069);
nand U23231 (N_23231,N_19136,N_21384);
and U23232 (N_23232,N_21374,N_20025);
and U23233 (N_23233,N_19753,N_20334);
nand U23234 (N_23234,N_19300,N_20170);
and U23235 (N_23235,N_19237,N_21008);
or U23236 (N_23236,N_19958,N_19647);
or U23237 (N_23237,N_20753,N_19946);
or U23238 (N_23238,N_19375,N_19371);
nor U23239 (N_23239,N_21478,N_19837);
nand U23240 (N_23240,N_19582,N_20157);
nor U23241 (N_23241,N_19863,N_19838);
nor U23242 (N_23242,N_19345,N_20740);
nor U23243 (N_23243,N_20249,N_20358);
nand U23244 (N_23244,N_20167,N_19898);
and U23245 (N_23245,N_21079,N_20716);
nand U23246 (N_23246,N_20669,N_21107);
nand U23247 (N_23247,N_19847,N_19627);
or U23248 (N_23248,N_20553,N_18828);
xnor U23249 (N_23249,N_21261,N_19775);
nand U23250 (N_23250,N_21832,N_20135);
xnor U23251 (N_23251,N_19655,N_20679);
nor U23252 (N_23252,N_19181,N_21436);
nand U23253 (N_23253,N_18825,N_20017);
or U23254 (N_23254,N_21389,N_19066);
or U23255 (N_23255,N_20554,N_19807);
nor U23256 (N_23256,N_20023,N_19235);
and U23257 (N_23257,N_20058,N_20841);
and U23258 (N_23258,N_20857,N_21774);
or U23259 (N_23259,N_20398,N_19318);
nand U23260 (N_23260,N_20968,N_20862);
nand U23261 (N_23261,N_20612,N_19017);
xor U23262 (N_23262,N_20443,N_19560);
and U23263 (N_23263,N_20729,N_20163);
nor U23264 (N_23264,N_20626,N_19147);
or U23265 (N_23265,N_20844,N_20863);
nand U23266 (N_23266,N_19005,N_18891);
xnor U23267 (N_23267,N_18793,N_20159);
xor U23268 (N_23268,N_21375,N_19190);
xor U23269 (N_23269,N_20457,N_18985);
and U23270 (N_23270,N_20472,N_20279);
nand U23271 (N_23271,N_18757,N_19954);
nor U23272 (N_23272,N_21725,N_19007);
or U23273 (N_23273,N_20540,N_19172);
and U23274 (N_23274,N_20771,N_18786);
or U23275 (N_23275,N_21637,N_20648);
and U23276 (N_23276,N_20153,N_20405);
and U23277 (N_23277,N_21487,N_19949);
and U23278 (N_23278,N_20831,N_20274);
nor U23279 (N_23279,N_20057,N_19260);
and U23280 (N_23280,N_21046,N_18758);
and U23281 (N_23281,N_21146,N_20584);
nor U23282 (N_23282,N_20315,N_20970);
nand U23283 (N_23283,N_21067,N_18821);
nand U23284 (N_23284,N_21695,N_19194);
and U23285 (N_23285,N_18910,N_20006);
xnor U23286 (N_23286,N_20117,N_21282);
nand U23287 (N_23287,N_21550,N_20704);
xnor U23288 (N_23288,N_20075,N_19209);
xor U23289 (N_23289,N_20182,N_21312);
xnor U23290 (N_23290,N_21447,N_20486);
nor U23291 (N_23291,N_20943,N_18979);
and U23292 (N_23292,N_20592,N_19804);
nor U23293 (N_23293,N_19505,N_19834);
nor U23294 (N_23294,N_20026,N_20008);
xnor U23295 (N_23295,N_19806,N_19397);
nand U23296 (N_23296,N_21163,N_21189);
or U23297 (N_23297,N_21684,N_20861);
nand U23298 (N_23298,N_20231,N_20377);
nor U23299 (N_23299,N_20323,N_21463);
nor U23300 (N_23300,N_20111,N_21461);
xor U23301 (N_23301,N_21825,N_20877);
xnor U23302 (N_23302,N_20477,N_19262);
nand U23303 (N_23303,N_19752,N_19777);
or U23304 (N_23304,N_19689,N_19871);
and U23305 (N_23305,N_20574,N_20176);
or U23306 (N_23306,N_19780,N_20082);
or U23307 (N_23307,N_20996,N_20555);
nand U23308 (N_23308,N_21709,N_20278);
nand U23309 (N_23309,N_21698,N_18841);
nor U23310 (N_23310,N_19598,N_20531);
nand U23311 (N_23311,N_19557,N_18864);
xor U23312 (N_23312,N_19970,N_19709);
xnor U23313 (N_23313,N_21074,N_20619);
or U23314 (N_23314,N_20390,N_21452);
and U23315 (N_23315,N_19063,N_19718);
nand U23316 (N_23316,N_19299,N_19347);
and U23317 (N_23317,N_18846,N_20328);
and U23318 (N_23318,N_20811,N_19853);
xnor U23319 (N_23319,N_18909,N_21302);
xor U23320 (N_23320,N_19714,N_21664);
nor U23321 (N_23321,N_19400,N_20155);
nor U23322 (N_23322,N_21516,N_20431);
nand U23323 (N_23323,N_19742,N_19012);
nor U23324 (N_23324,N_19093,N_21092);
nor U23325 (N_23325,N_21351,N_19730);
or U23326 (N_23326,N_21047,N_20765);
nand U23327 (N_23327,N_20933,N_19212);
xnor U23328 (N_23328,N_18873,N_20793);
nand U23329 (N_23329,N_20214,N_21296);
nor U23330 (N_23330,N_20173,N_20257);
or U23331 (N_23331,N_20964,N_19961);
xor U23332 (N_23332,N_21513,N_21399);
nor U23333 (N_23333,N_21266,N_21412);
xnor U23334 (N_23334,N_19113,N_21379);
xnor U23335 (N_23335,N_19058,N_21645);
xnor U23336 (N_23336,N_21692,N_21551);
nand U23337 (N_23337,N_18759,N_19902);
and U23338 (N_23338,N_21746,N_21170);
or U23339 (N_23339,N_21359,N_19440);
and U23340 (N_23340,N_21142,N_20108);
nand U23341 (N_23341,N_19821,N_18922);
and U23342 (N_23342,N_20321,N_21179);
or U23343 (N_23343,N_21582,N_20125);
and U23344 (N_23344,N_20427,N_20632);
and U23345 (N_23345,N_21385,N_19129);
and U23346 (N_23346,N_21649,N_21014);
nor U23347 (N_23347,N_18911,N_21670);
nand U23348 (N_23348,N_19287,N_20657);
or U23349 (N_23349,N_19258,N_19920);
nor U23350 (N_23350,N_20699,N_20442);
nor U23351 (N_23351,N_19401,N_20586);
and U23352 (N_23352,N_20952,N_20084);
xor U23353 (N_23353,N_20936,N_21757);
xor U23354 (N_23354,N_20622,N_20146);
and U23355 (N_23355,N_19461,N_21072);
nand U23356 (N_23356,N_19342,N_21735);
nor U23357 (N_23357,N_18962,N_21247);
and U23358 (N_23358,N_21818,N_21571);
and U23359 (N_23359,N_19770,N_21323);
xnor U23360 (N_23360,N_18916,N_21190);
nand U23361 (N_23361,N_21377,N_19161);
xor U23362 (N_23362,N_21004,N_20843);
nand U23363 (N_23363,N_20810,N_19539);
and U23364 (N_23364,N_20899,N_21081);
xnor U23365 (N_23365,N_20116,N_20650);
xor U23366 (N_23366,N_19116,N_19049);
nand U23367 (N_23367,N_18946,N_19015);
or U23368 (N_23368,N_19152,N_20614);
xor U23369 (N_23369,N_21534,N_19796);
nand U23370 (N_23370,N_19189,N_20326);
nand U23371 (N_23371,N_19729,N_21806);
nor U23372 (N_23372,N_20536,N_19621);
or U23373 (N_23373,N_18928,N_20376);
xor U23374 (N_23374,N_18845,N_21678);
nand U23375 (N_23375,N_20460,N_19447);
nand U23376 (N_23376,N_20934,N_21324);
or U23377 (N_23377,N_19803,N_21715);
nor U23378 (N_23378,N_20719,N_20658);
and U23379 (N_23379,N_19743,N_20636);
xnor U23380 (N_23380,N_20269,N_20482);
or U23381 (N_23381,N_20703,N_18814);
xor U23382 (N_23382,N_20309,N_20097);
and U23383 (N_23383,N_21156,N_19665);
nand U23384 (N_23384,N_21184,N_21051);
xnor U23385 (N_23385,N_18976,N_21199);
and U23386 (N_23386,N_19056,N_19779);
nand U23387 (N_23387,N_19218,N_19546);
nand U23388 (N_23388,N_21751,N_21269);
nand U23389 (N_23389,N_20119,N_20902);
and U23390 (N_23390,N_19637,N_20166);
nor U23391 (N_23391,N_21816,N_21321);
nor U23392 (N_23392,N_19110,N_21078);
nor U23393 (N_23393,N_20988,N_21472);
xor U23394 (N_23394,N_20981,N_21059);
nor U23395 (N_23395,N_20454,N_20830);
nor U23396 (N_23396,N_21263,N_19451);
xnor U23397 (N_23397,N_18751,N_21306);
nor U23398 (N_23398,N_18843,N_19403);
xor U23399 (N_23399,N_19528,N_19741);
nor U23400 (N_23400,N_19488,N_19096);
nand U23401 (N_23401,N_20733,N_20104);
nor U23402 (N_23402,N_19632,N_19296);
or U23403 (N_23403,N_19092,N_20284);
or U23404 (N_23404,N_19394,N_20028);
nand U23405 (N_23405,N_21420,N_21509);
or U23406 (N_23406,N_18889,N_20625);
nor U23407 (N_23407,N_21061,N_21677);
or U23408 (N_23408,N_21162,N_20501);
and U23409 (N_23409,N_20639,N_19293);
or U23410 (N_23410,N_19707,N_21503);
nor U23411 (N_23411,N_20868,N_21120);
or U23412 (N_23412,N_19186,N_21248);
nand U23413 (N_23413,N_18999,N_20879);
and U23414 (N_23414,N_20847,N_20463);
nor U23415 (N_23415,N_21117,N_18868);
nor U23416 (N_23416,N_21279,N_19893);
nor U23417 (N_23417,N_19391,N_20038);
and U23418 (N_23418,N_20418,N_19767);
nor U23419 (N_23419,N_21365,N_20296);
and U23420 (N_23420,N_21576,N_19187);
and U23421 (N_23421,N_21824,N_19417);
nor U23422 (N_23422,N_19247,N_19764);
and U23423 (N_23423,N_19850,N_19704);
or U23424 (N_23424,N_19493,N_21201);
nand U23425 (N_23425,N_20985,N_19700);
or U23426 (N_23426,N_20775,N_20435);
or U23427 (N_23427,N_21180,N_20430);
nor U23428 (N_23428,N_20259,N_20561);
xor U23429 (N_23429,N_19122,N_18963);
and U23430 (N_23430,N_20475,N_20280);
and U23431 (N_23431,N_19836,N_19455);
and U23432 (N_23432,N_21406,N_21141);
xor U23433 (N_23433,N_19654,N_21409);
or U23434 (N_23434,N_21748,N_20566);
or U23435 (N_23435,N_19996,N_19442);
or U23436 (N_23436,N_20258,N_21434);
xnor U23437 (N_23437,N_20186,N_20313);
nor U23438 (N_23438,N_21130,N_19369);
or U23439 (N_23439,N_19945,N_19417);
and U23440 (N_23440,N_20259,N_21628);
nor U23441 (N_23441,N_18751,N_21809);
nor U23442 (N_23442,N_20519,N_19237);
nand U23443 (N_23443,N_19517,N_19580);
or U23444 (N_23444,N_19478,N_19788);
and U23445 (N_23445,N_19547,N_21438);
nor U23446 (N_23446,N_19290,N_20750);
and U23447 (N_23447,N_21847,N_21033);
and U23448 (N_23448,N_21207,N_21409);
and U23449 (N_23449,N_18759,N_20621);
nor U23450 (N_23450,N_21788,N_20586);
and U23451 (N_23451,N_19177,N_20698);
nand U23452 (N_23452,N_20004,N_19076);
xnor U23453 (N_23453,N_19812,N_21416);
xor U23454 (N_23454,N_20559,N_19546);
or U23455 (N_23455,N_21147,N_20116);
or U23456 (N_23456,N_20713,N_19286);
nor U23457 (N_23457,N_18989,N_21702);
nor U23458 (N_23458,N_20391,N_21610);
nor U23459 (N_23459,N_21028,N_18883);
and U23460 (N_23460,N_20926,N_21385);
and U23461 (N_23461,N_19707,N_20897);
xor U23462 (N_23462,N_21199,N_21699);
nand U23463 (N_23463,N_18818,N_19722);
xor U23464 (N_23464,N_21682,N_21085);
or U23465 (N_23465,N_20865,N_20378);
or U23466 (N_23466,N_19478,N_19938);
or U23467 (N_23467,N_21310,N_18786);
and U23468 (N_23468,N_21672,N_20918);
or U23469 (N_23469,N_20399,N_20619);
nor U23470 (N_23470,N_19252,N_21858);
nor U23471 (N_23471,N_20424,N_21728);
and U23472 (N_23472,N_20522,N_20681);
xnor U23473 (N_23473,N_18916,N_19284);
xnor U23474 (N_23474,N_21640,N_20287);
xnor U23475 (N_23475,N_21324,N_20605);
or U23476 (N_23476,N_19150,N_20477);
xnor U23477 (N_23477,N_20480,N_19910);
or U23478 (N_23478,N_19573,N_20581);
and U23479 (N_23479,N_21415,N_18849);
and U23480 (N_23480,N_21095,N_20735);
or U23481 (N_23481,N_19562,N_18843);
nor U23482 (N_23482,N_21007,N_21195);
or U23483 (N_23483,N_18929,N_19720);
or U23484 (N_23484,N_19473,N_19911);
nand U23485 (N_23485,N_20992,N_19388);
xnor U23486 (N_23486,N_21246,N_21627);
nand U23487 (N_23487,N_20903,N_21284);
nand U23488 (N_23488,N_20057,N_21013);
and U23489 (N_23489,N_20234,N_19441);
xor U23490 (N_23490,N_20223,N_21171);
nor U23491 (N_23491,N_19989,N_21034);
xnor U23492 (N_23492,N_21368,N_19646);
xnor U23493 (N_23493,N_21228,N_19234);
and U23494 (N_23494,N_20503,N_19702);
nor U23495 (N_23495,N_21517,N_18965);
xor U23496 (N_23496,N_20273,N_21647);
nor U23497 (N_23497,N_18787,N_20501);
and U23498 (N_23498,N_19699,N_21622);
xor U23499 (N_23499,N_19852,N_21740);
and U23500 (N_23500,N_19087,N_21523);
nor U23501 (N_23501,N_20528,N_19360);
nand U23502 (N_23502,N_20759,N_21411);
or U23503 (N_23503,N_19663,N_18876);
nand U23504 (N_23504,N_21320,N_20231);
nor U23505 (N_23505,N_21833,N_20531);
and U23506 (N_23506,N_21034,N_20089);
xnor U23507 (N_23507,N_20528,N_21553);
and U23508 (N_23508,N_20626,N_20122);
xnor U23509 (N_23509,N_20329,N_19829);
nor U23510 (N_23510,N_21439,N_20370);
and U23511 (N_23511,N_19962,N_18965);
xor U23512 (N_23512,N_21353,N_18801);
or U23513 (N_23513,N_19285,N_21476);
or U23514 (N_23514,N_18983,N_20325);
or U23515 (N_23515,N_21001,N_21633);
nor U23516 (N_23516,N_21131,N_19783);
nand U23517 (N_23517,N_21639,N_21164);
and U23518 (N_23518,N_21583,N_20833);
nor U23519 (N_23519,N_18945,N_20837);
nand U23520 (N_23520,N_19921,N_21081);
and U23521 (N_23521,N_21464,N_19421);
and U23522 (N_23522,N_20311,N_18905);
xnor U23523 (N_23523,N_20004,N_19764);
and U23524 (N_23524,N_20019,N_21601);
nand U23525 (N_23525,N_21680,N_18901);
xor U23526 (N_23526,N_20777,N_19907);
and U23527 (N_23527,N_20806,N_20948);
xnor U23528 (N_23528,N_18774,N_20439);
nand U23529 (N_23529,N_20338,N_19495);
xor U23530 (N_23530,N_21158,N_21211);
and U23531 (N_23531,N_19386,N_20298);
nand U23532 (N_23532,N_19099,N_20821);
nand U23533 (N_23533,N_20157,N_21443);
xnor U23534 (N_23534,N_19170,N_18881);
or U23535 (N_23535,N_20406,N_20464);
and U23536 (N_23536,N_20040,N_21205);
or U23537 (N_23537,N_20818,N_19126);
xnor U23538 (N_23538,N_19586,N_20757);
xor U23539 (N_23539,N_18963,N_20182);
nand U23540 (N_23540,N_20017,N_20870);
and U23541 (N_23541,N_20759,N_21714);
xnor U23542 (N_23542,N_20065,N_20523);
xor U23543 (N_23543,N_20916,N_21355);
and U23544 (N_23544,N_20041,N_18922);
or U23545 (N_23545,N_19205,N_21161);
nor U23546 (N_23546,N_19440,N_21300);
or U23547 (N_23547,N_21738,N_19428);
or U23548 (N_23548,N_19406,N_19328);
and U23549 (N_23549,N_20970,N_21426);
and U23550 (N_23550,N_21628,N_21341);
or U23551 (N_23551,N_21075,N_21304);
xnor U23552 (N_23552,N_20628,N_21356);
nor U23553 (N_23553,N_18912,N_20438);
and U23554 (N_23554,N_21674,N_21779);
nor U23555 (N_23555,N_21150,N_20490);
xnor U23556 (N_23556,N_19798,N_21378);
nand U23557 (N_23557,N_20067,N_21311);
or U23558 (N_23558,N_19973,N_21108);
and U23559 (N_23559,N_19477,N_19807);
and U23560 (N_23560,N_20121,N_20558);
and U23561 (N_23561,N_19701,N_21270);
xnor U23562 (N_23562,N_18952,N_19439);
nor U23563 (N_23563,N_20770,N_19603);
nor U23564 (N_23564,N_18776,N_19811);
nand U23565 (N_23565,N_19382,N_21488);
nand U23566 (N_23566,N_21096,N_19842);
and U23567 (N_23567,N_18764,N_21515);
or U23568 (N_23568,N_19487,N_19205);
xor U23569 (N_23569,N_19690,N_19816);
and U23570 (N_23570,N_19644,N_19060);
and U23571 (N_23571,N_19744,N_20295);
xor U23572 (N_23572,N_20742,N_18783);
and U23573 (N_23573,N_20052,N_21138);
nand U23574 (N_23574,N_20833,N_20637);
nand U23575 (N_23575,N_21687,N_19142);
nor U23576 (N_23576,N_21871,N_20319);
or U23577 (N_23577,N_21165,N_20371);
and U23578 (N_23578,N_19445,N_20251);
nand U23579 (N_23579,N_18830,N_19247);
nand U23580 (N_23580,N_19170,N_19485);
nand U23581 (N_23581,N_19332,N_20626);
nor U23582 (N_23582,N_19491,N_20277);
xor U23583 (N_23583,N_20599,N_21355);
and U23584 (N_23584,N_19094,N_21160);
nor U23585 (N_23585,N_20160,N_20272);
and U23586 (N_23586,N_20293,N_21439);
nor U23587 (N_23587,N_20364,N_19508);
xnor U23588 (N_23588,N_20877,N_21374);
and U23589 (N_23589,N_21642,N_18889);
xor U23590 (N_23590,N_20685,N_20190);
nand U23591 (N_23591,N_19362,N_19634);
or U23592 (N_23592,N_21076,N_21332);
nand U23593 (N_23593,N_18924,N_19595);
and U23594 (N_23594,N_21483,N_18958);
and U23595 (N_23595,N_20439,N_19770);
and U23596 (N_23596,N_19447,N_21847);
nor U23597 (N_23597,N_21085,N_19717);
xor U23598 (N_23598,N_19604,N_21447);
or U23599 (N_23599,N_19398,N_20924);
nand U23600 (N_23600,N_19418,N_19487);
nor U23601 (N_23601,N_21574,N_21018);
xnor U23602 (N_23602,N_21019,N_21434);
xor U23603 (N_23603,N_20936,N_20202);
nor U23604 (N_23604,N_18931,N_18962);
or U23605 (N_23605,N_19138,N_19549);
nand U23606 (N_23606,N_19470,N_19237);
and U23607 (N_23607,N_19367,N_20453);
or U23608 (N_23608,N_19789,N_21291);
nand U23609 (N_23609,N_21838,N_21204);
and U23610 (N_23610,N_21237,N_18982);
xor U23611 (N_23611,N_21649,N_19050);
nand U23612 (N_23612,N_21164,N_19381);
nor U23613 (N_23613,N_19588,N_20330);
and U23614 (N_23614,N_20894,N_19439);
and U23615 (N_23615,N_19991,N_19439);
nand U23616 (N_23616,N_21849,N_20815);
nor U23617 (N_23617,N_18940,N_21746);
nor U23618 (N_23618,N_19843,N_21343);
nor U23619 (N_23619,N_18983,N_21023);
nor U23620 (N_23620,N_20628,N_19719);
and U23621 (N_23621,N_20003,N_18837);
or U23622 (N_23622,N_18849,N_21661);
or U23623 (N_23623,N_20380,N_19666);
and U23624 (N_23624,N_19230,N_20216);
or U23625 (N_23625,N_19548,N_21104);
nor U23626 (N_23626,N_18881,N_21569);
and U23627 (N_23627,N_18902,N_19984);
or U23628 (N_23628,N_18976,N_19971);
and U23629 (N_23629,N_19755,N_20923);
and U23630 (N_23630,N_18820,N_19374);
nand U23631 (N_23631,N_19588,N_21489);
xor U23632 (N_23632,N_19209,N_21753);
nor U23633 (N_23633,N_20836,N_19176);
nand U23634 (N_23634,N_19221,N_20755);
and U23635 (N_23635,N_18787,N_21445);
nand U23636 (N_23636,N_21469,N_21768);
xnor U23637 (N_23637,N_21615,N_19523);
nand U23638 (N_23638,N_19277,N_20891);
or U23639 (N_23639,N_19493,N_19166);
and U23640 (N_23640,N_21246,N_20395);
or U23641 (N_23641,N_20536,N_21498);
nor U23642 (N_23642,N_21707,N_20725);
and U23643 (N_23643,N_19657,N_21138);
nand U23644 (N_23644,N_19610,N_20695);
and U23645 (N_23645,N_21632,N_19898);
and U23646 (N_23646,N_20214,N_21390);
nor U23647 (N_23647,N_19774,N_20658);
and U23648 (N_23648,N_20191,N_20757);
and U23649 (N_23649,N_21014,N_21741);
xnor U23650 (N_23650,N_20792,N_19467);
nor U23651 (N_23651,N_18828,N_19663);
or U23652 (N_23652,N_19178,N_19413);
and U23653 (N_23653,N_20736,N_19148);
xnor U23654 (N_23654,N_19752,N_19849);
or U23655 (N_23655,N_21351,N_19561);
and U23656 (N_23656,N_20473,N_20332);
nand U23657 (N_23657,N_21545,N_20242);
or U23658 (N_23658,N_20824,N_21061);
or U23659 (N_23659,N_21799,N_21413);
and U23660 (N_23660,N_21729,N_20680);
and U23661 (N_23661,N_21698,N_21273);
nor U23662 (N_23662,N_20844,N_20442);
and U23663 (N_23663,N_20070,N_19918);
nand U23664 (N_23664,N_20336,N_21862);
nor U23665 (N_23665,N_19157,N_20087);
or U23666 (N_23666,N_19403,N_20487);
xor U23667 (N_23667,N_19706,N_20662);
nor U23668 (N_23668,N_20155,N_20731);
and U23669 (N_23669,N_21316,N_19959);
and U23670 (N_23670,N_20473,N_19416);
or U23671 (N_23671,N_20156,N_19399);
or U23672 (N_23672,N_21271,N_19162);
xnor U23673 (N_23673,N_20787,N_21069);
xor U23674 (N_23674,N_20855,N_18895);
or U23675 (N_23675,N_18838,N_21369);
nor U23676 (N_23676,N_20703,N_19640);
nor U23677 (N_23677,N_20408,N_20057);
nand U23678 (N_23678,N_18958,N_20897);
and U23679 (N_23679,N_20402,N_21631);
xor U23680 (N_23680,N_20117,N_20182);
nor U23681 (N_23681,N_21032,N_19873);
nor U23682 (N_23682,N_18889,N_20976);
and U23683 (N_23683,N_21655,N_19384);
nand U23684 (N_23684,N_20168,N_19367);
xor U23685 (N_23685,N_19732,N_21151);
nor U23686 (N_23686,N_19890,N_20750);
nor U23687 (N_23687,N_20453,N_19679);
or U23688 (N_23688,N_18946,N_19014);
or U23689 (N_23689,N_19588,N_19766);
nand U23690 (N_23690,N_19933,N_21279);
nand U23691 (N_23691,N_21308,N_19308);
xnor U23692 (N_23692,N_18829,N_19286);
and U23693 (N_23693,N_20273,N_21321);
nand U23694 (N_23694,N_20986,N_19948);
nor U23695 (N_23695,N_20555,N_20121);
and U23696 (N_23696,N_20888,N_20622);
nor U23697 (N_23697,N_18818,N_19330);
and U23698 (N_23698,N_21045,N_20223);
and U23699 (N_23699,N_21139,N_21076);
and U23700 (N_23700,N_20172,N_18869);
and U23701 (N_23701,N_18803,N_19446);
and U23702 (N_23702,N_20553,N_19690);
and U23703 (N_23703,N_19357,N_20631);
nand U23704 (N_23704,N_20289,N_20018);
or U23705 (N_23705,N_19360,N_20923);
and U23706 (N_23706,N_20529,N_20611);
or U23707 (N_23707,N_18774,N_21771);
or U23708 (N_23708,N_20204,N_20023);
nand U23709 (N_23709,N_20160,N_20221);
nand U23710 (N_23710,N_20406,N_20593);
nor U23711 (N_23711,N_20367,N_21291);
or U23712 (N_23712,N_19201,N_20807);
nand U23713 (N_23713,N_18975,N_19218);
xnor U23714 (N_23714,N_21133,N_20368);
or U23715 (N_23715,N_20247,N_19888);
xor U23716 (N_23716,N_19615,N_20392);
or U23717 (N_23717,N_21085,N_21425);
and U23718 (N_23718,N_19016,N_18965);
nand U23719 (N_23719,N_20088,N_21088);
nand U23720 (N_23720,N_19751,N_21765);
nor U23721 (N_23721,N_20946,N_18824);
xnor U23722 (N_23722,N_19483,N_19498);
or U23723 (N_23723,N_19794,N_18848);
nand U23724 (N_23724,N_20107,N_21390);
or U23725 (N_23725,N_20573,N_19342);
xnor U23726 (N_23726,N_20131,N_21412);
xor U23727 (N_23727,N_21829,N_19761);
nor U23728 (N_23728,N_19434,N_19328);
xor U23729 (N_23729,N_20881,N_19093);
nor U23730 (N_23730,N_19114,N_20964);
and U23731 (N_23731,N_20157,N_19291);
nand U23732 (N_23732,N_20176,N_21728);
nand U23733 (N_23733,N_20212,N_20606);
nor U23734 (N_23734,N_19243,N_21546);
nand U23735 (N_23735,N_20967,N_21413);
nor U23736 (N_23736,N_18990,N_19400);
and U23737 (N_23737,N_19505,N_20574);
nor U23738 (N_23738,N_20797,N_19847);
nor U23739 (N_23739,N_21379,N_21243);
nand U23740 (N_23740,N_20840,N_21683);
or U23741 (N_23741,N_18750,N_19652);
nand U23742 (N_23742,N_21219,N_20230);
xor U23743 (N_23743,N_20374,N_19406);
or U23744 (N_23744,N_20903,N_19021);
or U23745 (N_23745,N_20199,N_19578);
xnor U23746 (N_23746,N_21167,N_21851);
xor U23747 (N_23747,N_18845,N_20443);
xnor U23748 (N_23748,N_20042,N_18918);
nand U23749 (N_23749,N_19078,N_19237);
nand U23750 (N_23750,N_20119,N_21618);
nand U23751 (N_23751,N_18940,N_21450);
nand U23752 (N_23752,N_20288,N_20425);
or U23753 (N_23753,N_20822,N_21084);
and U23754 (N_23754,N_19723,N_19928);
or U23755 (N_23755,N_19529,N_20798);
and U23756 (N_23756,N_19966,N_20470);
or U23757 (N_23757,N_20252,N_20826);
xnor U23758 (N_23758,N_19232,N_21195);
nand U23759 (N_23759,N_20408,N_19506);
nor U23760 (N_23760,N_21156,N_20746);
and U23761 (N_23761,N_20091,N_19439);
and U23762 (N_23762,N_20113,N_20872);
nor U23763 (N_23763,N_20164,N_21546);
xnor U23764 (N_23764,N_18952,N_19095);
xor U23765 (N_23765,N_20223,N_19610);
and U23766 (N_23766,N_20768,N_18786);
and U23767 (N_23767,N_21678,N_19634);
nor U23768 (N_23768,N_20072,N_20542);
nand U23769 (N_23769,N_21525,N_19759);
or U23770 (N_23770,N_21676,N_19569);
xor U23771 (N_23771,N_19146,N_21112);
nand U23772 (N_23772,N_20825,N_19918);
or U23773 (N_23773,N_20652,N_19233);
xor U23774 (N_23774,N_19000,N_21733);
and U23775 (N_23775,N_20455,N_20535);
nand U23776 (N_23776,N_21436,N_18985);
xnor U23777 (N_23777,N_18948,N_19627);
or U23778 (N_23778,N_19627,N_21861);
nand U23779 (N_23779,N_21823,N_19286);
nor U23780 (N_23780,N_19202,N_20682);
and U23781 (N_23781,N_21581,N_21597);
nand U23782 (N_23782,N_19152,N_20330);
nand U23783 (N_23783,N_19689,N_19171);
nand U23784 (N_23784,N_18863,N_21688);
nand U23785 (N_23785,N_20792,N_20409);
nand U23786 (N_23786,N_18790,N_18767);
or U23787 (N_23787,N_18953,N_18980);
xor U23788 (N_23788,N_21258,N_20634);
nand U23789 (N_23789,N_19973,N_21645);
or U23790 (N_23790,N_21211,N_20850);
nor U23791 (N_23791,N_20351,N_19355);
and U23792 (N_23792,N_21148,N_21085);
nand U23793 (N_23793,N_19249,N_19028);
and U23794 (N_23794,N_19397,N_20526);
nand U23795 (N_23795,N_20753,N_19750);
nand U23796 (N_23796,N_21231,N_20843);
nand U23797 (N_23797,N_19463,N_20468);
and U23798 (N_23798,N_21767,N_19537);
nand U23799 (N_23799,N_19220,N_19842);
or U23800 (N_23800,N_19622,N_19261);
nand U23801 (N_23801,N_20530,N_20025);
or U23802 (N_23802,N_21090,N_20909);
nand U23803 (N_23803,N_19592,N_21052);
xnor U23804 (N_23804,N_19008,N_20660);
xor U23805 (N_23805,N_18869,N_19590);
xor U23806 (N_23806,N_18834,N_19385);
xor U23807 (N_23807,N_19248,N_19340);
and U23808 (N_23808,N_21477,N_21668);
or U23809 (N_23809,N_21220,N_18915);
or U23810 (N_23810,N_19197,N_20188);
nor U23811 (N_23811,N_18970,N_19544);
and U23812 (N_23812,N_20311,N_19572);
nand U23813 (N_23813,N_21576,N_20762);
or U23814 (N_23814,N_20429,N_21613);
nand U23815 (N_23815,N_21513,N_19060);
nand U23816 (N_23816,N_21682,N_21440);
and U23817 (N_23817,N_20983,N_19901);
or U23818 (N_23818,N_20169,N_19637);
or U23819 (N_23819,N_18793,N_19842);
nand U23820 (N_23820,N_21049,N_19333);
nor U23821 (N_23821,N_21696,N_20617);
nand U23822 (N_23822,N_20589,N_21794);
xor U23823 (N_23823,N_20021,N_21272);
xnor U23824 (N_23824,N_20561,N_21089);
nor U23825 (N_23825,N_21128,N_20998);
xnor U23826 (N_23826,N_19432,N_19838);
nor U23827 (N_23827,N_20803,N_20584);
xor U23828 (N_23828,N_20383,N_20068);
xnor U23829 (N_23829,N_19024,N_21686);
xnor U23830 (N_23830,N_19148,N_21316);
nor U23831 (N_23831,N_19507,N_19627);
nor U23832 (N_23832,N_21711,N_21288);
or U23833 (N_23833,N_21695,N_18787);
or U23834 (N_23834,N_20224,N_19745);
and U23835 (N_23835,N_19429,N_18848);
nand U23836 (N_23836,N_20054,N_21362);
nand U23837 (N_23837,N_21460,N_20042);
xor U23838 (N_23838,N_21090,N_18832);
nand U23839 (N_23839,N_21705,N_20701);
xor U23840 (N_23840,N_19660,N_19330);
and U23841 (N_23841,N_19981,N_20092);
or U23842 (N_23842,N_20867,N_20647);
or U23843 (N_23843,N_20233,N_19396);
or U23844 (N_23844,N_19007,N_19136);
and U23845 (N_23845,N_19401,N_19306);
and U23846 (N_23846,N_20662,N_21697);
nand U23847 (N_23847,N_19254,N_18866);
xnor U23848 (N_23848,N_18928,N_20474);
and U23849 (N_23849,N_20782,N_19459);
and U23850 (N_23850,N_21404,N_19966);
nor U23851 (N_23851,N_21446,N_20395);
and U23852 (N_23852,N_20804,N_19123);
nor U23853 (N_23853,N_21322,N_21750);
nor U23854 (N_23854,N_19329,N_19182);
nand U23855 (N_23855,N_20316,N_20909);
xor U23856 (N_23856,N_19398,N_21156);
xnor U23857 (N_23857,N_18907,N_19243);
or U23858 (N_23858,N_20972,N_18859);
nand U23859 (N_23859,N_19636,N_20559);
or U23860 (N_23860,N_21187,N_20054);
nor U23861 (N_23861,N_20016,N_21714);
and U23862 (N_23862,N_20323,N_18765);
and U23863 (N_23863,N_20866,N_21687);
or U23864 (N_23864,N_20254,N_19842);
xor U23865 (N_23865,N_20760,N_20280);
nor U23866 (N_23866,N_21263,N_19637);
nand U23867 (N_23867,N_20354,N_21332);
or U23868 (N_23868,N_20672,N_19335);
and U23869 (N_23869,N_20814,N_19562);
xnor U23870 (N_23870,N_20169,N_19002);
xnor U23871 (N_23871,N_20478,N_21031);
nor U23872 (N_23872,N_20641,N_19474);
or U23873 (N_23873,N_20978,N_18775);
or U23874 (N_23874,N_20266,N_21572);
nor U23875 (N_23875,N_21254,N_18884);
or U23876 (N_23876,N_20722,N_19579);
xnor U23877 (N_23877,N_19402,N_21629);
nand U23878 (N_23878,N_20748,N_21707);
xor U23879 (N_23879,N_21687,N_19560);
or U23880 (N_23880,N_21718,N_19185);
nor U23881 (N_23881,N_20412,N_21428);
or U23882 (N_23882,N_19202,N_19103);
or U23883 (N_23883,N_20859,N_18758);
xor U23884 (N_23884,N_21704,N_21519);
nand U23885 (N_23885,N_20732,N_21379);
nand U23886 (N_23886,N_21368,N_20036);
xor U23887 (N_23887,N_19980,N_20831);
and U23888 (N_23888,N_20250,N_20845);
xnor U23889 (N_23889,N_18963,N_20862);
xnor U23890 (N_23890,N_21519,N_18973);
nand U23891 (N_23891,N_19410,N_19772);
nor U23892 (N_23892,N_19236,N_19066);
xnor U23893 (N_23893,N_20900,N_20533);
and U23894 (N_23894,N_19892,N_21726);
nand U23895 (N_23895,N_21826,N_21547);
xnor U23896 (N_23896,N_21790,N_19859);
or U23897 (N_23897,N_20421,N_18883);
xor U23898 (N_23898,N_20677,N_19034);
and U23899 (N_23899,N_20950,N_19606);
nand U23900 (N_23900,N_19987,N_20774);
and U23901 (N_23901,N_20672,N_21859);
xor U23902 (N_23902,N_19740,N_20512);
xnor U23903 (N_23903,N_20814,N_20682);
or U23904 (N_23904,N_19118,N_19919);
nand U23905 (N_23905,N_18830,N_20720);
xor U23906 (N_23906,N_20846,N_20250);
nand U23907 (N_23907,N_21131,N_20287);
or U23908 (N_23908,N_21095,N_18923);
or U23909 (N_23909,N_19653,N_19357);
or U23910 (N_23910,N_21135,N_21171);
nand U23911 (N_23911,N_20489,N_21055);
xnor U23912 (N_23912,N_18883,N_20589);
xor U23913 (N_23913,N_21859,N_19209);
or U23914 (N_23914,N_20225,N_20099);
nand U23915 (N_23915,N_20450,N_19709);
and U23916 (N_23916,N_20707,N_20638);
or U23917 (N_23917,N_19783,N_20621);
and U23918 (N_23918,N_19828,N_18995);
and U23919 (N_23919,N_19097,N_20392);
or U23920 (N_23920,N_21825,N_20971);
xnor U23921 (N_23921,N_20667,N_20882);
nor U23922 (N_23922,N_20165,N_21359);
xor U23923 (N_23923,N_20817,N_21088);
xnor U23924 (N_23924,N_21829,N_20610);
nor U23925 (N_23925,N_19597,N_18941);
or U23926 (N_23926,N_20855,N_20957);
nor U23927 (N_23927,N_20563,N_20108);
xnor U23928 (N_23928,N_19289,N_19034);
nand U23929 (N_23929,N_21405,N_18845);
or U23930 (N_23930,N_20937,N_19019);
and U23931 (N_23931,N_19321,N_21733);
xor U23932 (N_23932,N_21661,N_21114);
nand U23933 (N_23933,N_21518,N_19878);
and U23934 (N_23934,N_19429,N_20202);
xnor U23935 (N_23935,N_21335,N_21792);
nand U23936 (N_23936,N_21841,N_21126);
nand U23937 (N_23937,N_19808,N_20659);
nand U23938 (N_23938,N_19354,N_20531);
nand U23939 (N_23939,N_19877,N_21120);
or U23940 (N_23940,N_20924,N_20629);
nor U23941 (N_23941,N_19060,N_20390);
nor U23942 (N_23942,N_20606,N_21438);
nand U23943 (N_23943,N_19618,N_20982);
nand U23944 (N_23944,N_20142,N_19352);
or U23945 (N_23945,N_18959,N_20143);
or U23946 (N_23946,N_20750,N_20498);
nor U23947 (N_23947,N_21266,N_19705);
and U23948 (N_23948,N_19391,N_18885);
nand U23949 (N_23949,N_21694,N_19470);
or U23950 (N_23950,N_18817,N_21421);
or U23951 (N_23951,N_20815,N_18997);
nor U23952 (N_23952,N_21270,N_21166);
nand U23953 (N_23953,N_20554,N_21775);
xor U23954 (N_23954,N_20643,N_19968);
and U23955 (N_23955,N_21771,N_20390);
xnor U23956 (N_23956,N_18853,N_20844);
xnor U23957 (N_23957,N_21163,N_20942);
nor U23958 (N_23958,N_19139,N_20118);
or U23959 (N_23959,N_21161,N_19340);
and U23960 (N_23960,N_21055,N_19332);
nand U23961 (N_23961,N_19829,N_21645);
or U23962 (N_23962,N_20663,N_20579);
nor U23963 (N_23963,N_19761,N_20901);
and U23964 (N_23964,N_20579,N_21757);
xnor U23965 (N_23965,N_20751,N_20676);
nor U23966 (N_23966,N_21556,N_19725);
nor U23967 (N_23967,N_19335,N_20456);
nand U23968 (N_23968,N_20056,N_20821);
nand U23969 (N_23969,N_20770,N_19957);
xor U23970 (N_23970,N_19104,N_20059);
nor U23971 (N_23971,N_21809,N_20670);
or U23972 (N_23972,N_20290,N_20408);
or U23973 (N_23973,N_20437,N_19820);
nor U23974 (N_23974,N_21820,N_21732);
or U23975 (N_23975,N_20957,N_21342);
nor U23976 (N_23976,N_18899,N_21424);
and U23977 (N_23977,N_21317,N_19837);
nand U23978 (N_23978,N_20210,N_19438);
and U23979 (N_23979,N_21790,N_19728);
or U23980 (N_23980,N_19822,N_19993);
and U23981 (N_23981,N_21655,N_20900);
nor U23982 (N_23982,N_21812,N_19609);
xnor U23983 (N_23983,N_19210,N_20205);
or U23984 (N_23984,N_19011,N_20641);
nand U23985 (N_23985,N_20803,N_21594);
and U23986 (N_23986,N_21391,N_21823);
nor U23987 (N_23987,N_20589,N_19967);
and U23988 (N_23988,N_20346,N_21679);
nand U23989 (N_23989,N_21667,N_20666);
and U23990 (N_23990,N_21842,N_21608);
xor U23991 (N_23991,N_19094,N_21529);
xor U23992 (N_23992,N_21116,N_20462);
nor U23993 (N_23993,N_21836,N_18856);
or U23994 (N_23994,N_19466,N_19973);
nor U23995 (N_23995,N_20091,N_19158);
and U23996 (N_23996,N_19367,N_20750);
or U23997 (N_23997,N_20869,N_21071);
nor U23998 (N_23998,N_20616,N_21201);
xor U23999 (N_23999,N_20513,N_18850);
or U24000 (N_24000,N_18975,N_21062);
nand U24001 (N_24001,N_20165,N_19388);
or U24002 (N_24002,N_19925,N_19880);
and U24003 (N_24003,N_21656,N_19540);
and U24004 (N_24004,N_21558,N_21790);
and U24005 (N_24005,N_19206,N_21634);
nand U24006 (N_24006,N_19026,N_19231);
nor U24007 (N_24007,N_20963,N_20066);
nand U24008 (N_24008,N_20513,N_18977);
nand U24009 (N_24009,N_21221,N_21743);
nand U24010 (N_24010,N_20983,N_21592);
and U24011 (N_24011,N_21468,N_20539);
and U24012 (N_24012,N_20288,N_19114);
nor U24013 (N_24013,N_21566,N_20823);
or U24014 (N_24014,N_20190,N_19598);
nand U24015 (N_24015,N_19795,N_20299);
and U24016 (N_24016,N_20649,N_21517);
and U24017 (N_24017,N_21133,N_19288);
xor U24018 (N_24018,N_19839,N_20931);
xnor U24019 (N_24019,N_21235,N_21060);
nand U24020 (N_24020,N_20955,N_20860);
and U24021 (N_24021,N_19100,N_19134);
xnor U24022 (N_24022,N_20414,N_20387);
xnor U24023 (N_24023,N_20259,N_20337);
nand U24024 (N_24024,N_20319,N_19671);
nand U24025 (N_24025,N_19528,N_19126);
xnor U24026 (N_24026,N_18784,N_20484);
nor U24027 (N_24027,N_19206,N_19689);
and U24028 (N_24028,N_20821,N_19269);
nor U24029 (N_24029,N_18904,N_20963);
nand U24030 (N_24030,N_20092,N_18994);
or U24031 (N_24031,N_20952,N_19648);
xnor U24032 (N_24032,N_21430,N_20208);
or U24033 (N_24033,N_19879,N_19168);
and U24034 (N_24034,N_19853,N_21185);
nor U24035 (N_24035,N_21369,N_20797);
and U24036 (N_24036,N_19243,N_18888);
and U24037 (N_24037,N_21731,N_21142);
nand U24038 (N_24038,N_19508,N_20462);
nand U24039 (N_24039,N_19984,N_21672);
and U24040 (N_24040,N_19450,N_19525);
xnor U24041 (N_24041,N_21764,N_20835);
xnor U24042 (N_24042,N_21650,N_19695);
or U24043 (N_24043,N_20072,N_20320);
or U24044 (N_24044,N_19775,N_20162);
xor U24045 (N_24045,N_21023,N_21191);
nand U24046 (N_24046,N_20067,N_19277);
xnor U24047 (N_24047,N_21099,N_18783);
nor U24048 (N_24048,N_21214,N_19457);
nand U24049 (N_24049,N_18847,N_21386);
nor U24050 (N_24050,N_19819,N_19370);
xor U24051 (N_24051,N_20539,N_20973);
nand U24052 (N_24052,N_21822,N_21719);
nand U24053 (N_24053,N_18869,N_20780);
nor U24054 (N_24054,N_20884,N_21064);
nor U24055 (N_24055,N_20220,N_18766);
nor U24056 (N_24056,N_19511,N_21834);
xnor U24057 (N_24057,N_21204,N_20480);
nand U24058 (N_24058,N_19235,N_20636);
nand U24059 (N_24059,N_19501,N_19784);
and U24060 (N_24060,N_20088,N_18796);
nand U24061 (N_24061,N_18800,N_21760);
nand U24062 (N_24062,N_20671,N_19409);
and U24063 (N_24063,N_18820,N_21777);
and U24064 (N_24064,N_19998,N_19426);
nand U24065 (N_24065,N_21046,N_18945);
or U24066 (N_24066,N_21874,N_20373);
nor U24067 (N_24067,N_20797,N_21348);
and U24068 (N_24068,N_21647,N_20691);
or U24069 (N_24069,N_19320,N_20598);
nand U24070 (N_24070,N_19107,N_19234);
nand U24071 (N_24071,N_20104,N_19334);
or U24072 (N_24072,N_18759,N_21691);
nand U24073 (N_24073,N_20234,N_18972);
and U24074 (N_24074,N_20545,N_19360);
nand U24075 (N_24075,N_20341,N_20355);
nand U24076 (N_24076,N_20141,N_19871);
and U24077 (N_24077,N_20636,N_21594);
nor U24078 (N_24078,N_20963,N_19470);
xor U24079 (N_24079,N_20515,N_21154);
nand U24080 (N_24080,N_19677,N_20352);
or U24081 (N_24081,N_20899,N_19321);
xnor U24082 (N_24082,N_20861,N_21029);
nand U24083 (N_24083,N_19206,N_20692);
or U24084 (N_24084,N_19881,N_19076);
nand U24085 (N_24085,N_19995,N_20392);
xnor U24086 (N_24086,N_18784,N_20277);
or U24087 (N_24087,N_21528,N_20910);
and U24088 (N_24088,N_20258,N_19631);
and U24089 (N_24089,N_21614,N_19387);
nor U24090 (N_24090,N_20126,N_19422);
and U24091 (N_24091,N_19540,N_20859);
or U24092 (N_24092,N_21376,N_20272);
and U24093 (N_24093,N_19489,N_21845);
xor U24094 (N_24094,N_19433,N_20223);
or U24095 (N_24095,N_19926,N_21172);
and U24096 (N_24096,N_21437,N_19911);
nand U24097 (N_24097,N_18848,N_21797);
xor U24098 (N_24098,N_20106,N_19435);
xor U24099 (N_24099,N_19438,N_20257);
nor U24100 (N_24100,N_20890,N_19254);
nand U24101 (N_24101,N_21187,N_18758);
nand U24102 (N_24102,N_19735,N_21261);
and U24103 (N_24103,N_20946,N_20730);
or U24104 (N_24104,N_21285,N_18832);
or U24105 (N_24105,N_20518,N_19759);
and U24106 (N_24106,N_20626,N_18755);
nand U24107 (N_24107,N_19227,N_19521);
xor U24108 (N_24108,N_21272,N_21467);
nand U24109 (N_24109,N_19953,N_20290);
nand U24110 (N_24110,N_20628,N_21828);
and U24111 (N_24111,N_20228,N_20295);
xor U24112 (N_24112,N_20092,N_20885);
nand U24113 (N_24113,N_19418,N_20800);
or U24114 (N_24114,N_21088,N_19919);
or U24115 (N_24115,N_21773,N_21527);
and U24116 (N_24116,N_21155,N_20737);
nor U24117 (N_24117,N_20712,N_21638);
and U24118 (N_24118,N_20594,N_20992);
nor U24119 (N_24119,N_21284,N_20280);
xnor U24120 (N_24120,N_20417,N_19286);
and U24121 (N_24121,N_20449,N_21644);
nor U24122 (N_24122,N_19924,N_20674);
nand U24123 (N_24123,N_19841,N_20770);
and U24124 (N_24124,N_21835,N_20156);
and U24125 (N_24125,N_18831,N_19323);
xor U24126 (N_24126,N_18926,N_20104);
nand U24127 (N_24127,N_20360,N_20704);
or U24128 (N_24128,N_19482,N_20231);
and U24129 (N_24129,N_20845,N_21008);
nand U24130 (N_24130,N_21628,N_20632);
nor U24131 (N_24131,N_21586,N_21499);
nand U24132 (N_24132,N_19422,N_19649);
xor U24133 (N_24133,N_19723,N_20925);
nand U24134 (N_24134,N_19216,N_19337);
nand U24135 (N_24135,N_21001,N_19540);
nand U24136 (N_24136,N_21240,N_20120);
nor U24137 (N_24137,N_20272,N_20284);
or U24138 (N_24138,N_19075,N_20045);
nand U24139 (N_24139,N_19707,N_19699);
nor U24140 (N_24140,N_20443,N_18907);
and U24141 (N_24141,N_21362,N_20728);
nand U24142 (N_24142,N_20115,N_19957);
and U24143 (N_24143,N_20973,N_20892);
nor U24144 (N_24144,N_19741,N_20870);
nor U24145 (N_24145,N_21682,N_18955);
xnor U24146 (N_24146,N_19464,N_19525);
nor U24147 (N_24147,N_21848,N_20994);
or U24148 (N_24148,N_19376,N_21721);
or U24149 (N_24149,N_21675,N_20787);
or U24150 (N_24150,N_21796,N_19772);
and U24151 (N_24151,N_20686,N_19120);
nor U24152 (N_24152,N_21130,N_20212);
xor U24153 (N_24153,N_20610,N_21015);
and U24154 (N_24154,N_19462,N_20763);
nor U24155 (N_24155,N_21180,N_20128);
nand U24156 (N_24156,N_18822,N_20601);
nor U24157 (N_24157,N_20842,N_20276);
nor U24158 (N_24158,N_20947,N_20477);
nand U24159 (N_24159,N_19895,N_21256);
nor U24160 (N_24160,N_19784,N_21716);
and U24161 (N_24161,N_21246,N_20402);
nor U24162 (N_24162,N_19508,N_20139);
nor U24163 (N_24163,N_19373,N_20946);
and U24164 (N_24164,N_19694,N_19072);
xor U24165 (N_24165,N_20849,N_19506);
xnor U24166 (N_24166,N_20694,N_20864);
xnor U24167 (N_24167,N_18846,N_19432);
and U24168 (N_24168,N_21531,N_19507);
xnor U24169 (N_24169,N_19458,N_20499);
and U24170 (N_24170,N_19184,N_19135);
and U24171 (N_24171,N_20762,N_19850);
xor U24172 (N_24172,N_20761,N_18960);
and U24173 (N_24173,N_20212,N_21707);
and U24174 (N_24174,N_21095,N_20869);
xor U24175 (N_24175,N_21299,N_20909);
or U24176 (N_24176,N_20883,N_21548);
or U24177 (N_24177,N_21381,N_19961);
nand U24178 (N_24178,N_21208,N_20542);
or U24179 (N_24179,N_20758,N_21785);
and U24180 (N_24180,N_18903,N_19014);
xor U24181 (N_24181,N_20200,N_19607);
xor U24182 (N_24182,N_20166,N_18999);
or U24183 (N_24183,N_21171,N_18876);
nor U24184 (N_24184,N_19021,N_18804);
and U24185 (N_24185,N_19715,N_20104);
or U24186 (N_24186,N_19469,N_19961);
nand U24187 (N_24187,N_19555,N_20079);
or U24188 (N_24188,N_20494,N_20215);
nor U24189 (N_24189,N_21008,N_21486);
xnor U24190 (N_24190,N_21161,N_21562);
nand U24191 (N_24191,N_20289,N_20109);
nand U24192 (N_24192,N_20856,N_20843);
and U24193 (N_24193,N_21364,N_19130);
and U24194 (N_24194,N_20412,N_21448);
xor U24195 (N_24195,N_18999,N_18880);
xor U24196 (N_24196,N_20476,N_20327);
and U24197 (N_24197,N_20680,N_20174);
or U24198 (N_24198,N_21091,N_20556);
and U24199 (N_24199,N_20042,N_21750);
and U24200 (N_24200,N_21424,N_18889);
nand U24201 (N_24201,N_21489,N_19360);
or U24202 (N_24202,N_20800,N_19134);
nand U24203 (N_24203,N_20553,N_21747);
nand U24204 (N_24204,N_20057,N_20692);
or U24205 (N_24205,N_19467,N_21503);
nand U24206 (N_24206,N_20394,N_20545);
xor U24207 (N_24207,N_18974,N_19002);
nor U24208 (N_24208,N_20053,N_18886);
nor U24209 (N_24209,N_20515,N_21691);
xnor U24210 (N_24210,N_18750,N_20219);
xnor U24211 (N_24211,N_19493,N_20280);
xnor U24212 (N_24212,N_20998,N_21248);
and U24213 (N_24213,N_20399,N_18885);
nand U24214 (N_24214,N_20477,N_21130);
and U24215 (N_24215,N_19154,N_21649);
and U24216 (N_24216,N_21501,N_21700);
nand U24217 (N_24217,N_20329,N_21168);
or U24218 (N_24218,N_18833,N_21701);
or U24219 (N_24219,N_20822,N_21605);
xnor U24220 (N_24220,N_21157,N_19558);
or U24221 (N_24221,N_19305,N_19791);
xnor U24222 (N_24222,N_19507,N_21821);
xor U24223 (N_24223,N_20063,N_21409);
and U24224 (N_24224,N_20709,N_19580);
or U24225 (N_24225,N_19499,N_20831);
xor U24226 (N_24226,N_18873,N_20754);
and U24227 (N_24227,N_20105,N_20822);
nor U24228 (N_24228,N_19648,N_21157);
nor U24229 (N_24229,N_20673,N_18842);
nor U24230 (N_24230,N_21397,N_21276);
nand U24231 (N_24231,N_20633,N_19311);
and U24232 (N_24232,N_21056,N_18892);
or U24233 (N_24233,N_18912,N_21693);
nand U24234 (N_24234,N_19814,N_21136);
nand U24235 (N_24235,N_20720,N_19315);
nand U24236 (N_24236,N_18867,N_21073);
nand U24237 (N_24237,N_18895,N_20654);
or U24238 (N_24238,N_21719,N_19864);
or U24239 (N_24239,N_20803,N_20511);
and U24240 (N_24240,N_21834,N_18795);
or U24241 (N_24241,N_21729,N_19983);
nand U24242 (N_24242,N_21512,N_20895);
nor U24243 (N_24243,N_21865,N_20790);
xnor U24244 (N_24244,N_21331,N_19566);
and U24245 (N_24245,N_19060,N_19611);
xor U24246 (N_24246,N_21628,N_21742);
nand U24247 (N_24247,N_21562,N_21780);
and U24248 (N_24248,N_19368,N_19221);
or U24249 (N_24249,N_21836,N_20641);
or U24250 (N_24250,N_18853,N_21322);
and U24251 (N_24251,N_20068,N_20062);
and U24252 (N_24252,N_20547,N_21255);
xor U24253 (N_24253,N_20014,N_20588);
and U24254 (N_24254,N_20735,N_21328);
nand U24255 (N_24255,N_21710,N_20124);
and U24256 (N_24256,N_19432,N_20603);
nand U24257 (N_24257,N_20554,N_20137);
nand U24258 (N_24258,N_19179,N_21716);
nor U24259 (N_24259,N_18845,N_19541);
or U24260 (N_24260,N_20535,N_21421);
xnor U24261 (N_24261,N_21151,N_21790);
nand U24262 (N_24262,N_18922,N_21494);
or U24263 (N_24263,N_21831,N_21279);
nor U24264 (N_24264,N_19312,N_21466);
xnor U24265 (N_24265,N_18770,N_21389);
nand U24266 (N_24266,N_20067,N_19507);
xnor U24267 (N_24267,N_21578,N_19927);
nand U24268 (N_24268,N_20399,N_19134);
nor U24269 (N_24269,N_21272,N_21578);
nand U24270 (N_24270,N_20456,N_21387);
and U24271 (N_24271,N_21377,N_18803);
nor U24272 (N_24272,N_20596,N_20811);
or U24273 (N_24273,N_19821,N_20564);
or U24274 (N_24274,N_20475,N_21272);
and U24275 (N_24275,N_20979,N_21551);
or U24276 (N_24276,N_20598,N_21165);
xor U24277 (N_24277,N_18809,N_20571);
and U24278 (N_24278,N_19717,N_19203);
nand U24279 (N_24279,N_21556,N_20848);
nand U24280 (N_24280,N_21232,N_21662);
nand U24281 (N_24281,N_19208,N_19020);
or U24282 (N_24282,N_18976,N_20958);
or U24283 (N_24283,N_21277,N_21391);
nand U24284 (N_24284,N_18856,N_21656);
or U24285 (N_24285,N_18859,N_21139);
or U24286 (N_24286,N_19693,N_19013);
and U24287 (N_24287,N_19102,N_21564);
or U24288 (N_24288,N_19950,N_20829);
xor U24289 (N_24289,N_18827,N_18869);
and U24290 (N_24290,N_21258,N_19690);
xnor U24291 (N_24291,N_20219,N_21692);
nor U24292 (N_24292,N_19589,N_20675);
and U24293 (N_24293,N_19688,N_20060);
nor U24294 (N_24294,N_20869,N_21041);
xnor U24295 (N_24295,N_20145,N_20010);
nor U24296 (N_24296,N_19050,N_20101);
and U24297 (N_24297,N_19096,N_19980);
and U24298 (N_24298,N_20777,N_20253);
xor U24299 (N_24299,N_21163,N_21450);
and U24300 (N_24300,N_18876,N_20087);
and U24301 (N_24301,N_19903,N_20313);
or U24302 (N_24302,N_20072,N_20701);
and U24303 (N_24303,N_19940,N_19672);
nor U24304 (N_24304,N_20310,N_20363);
or U24305 (N_24305,N_19645,N_21645);
nand U24306 (N_24306,N_20311,N_21477);
xnor U24307 (N_24307,N_21291,N_21277);
and U24308 (N_24308,N_19135,N_21273);
nand U24309 (N_24309,N_21194,N_21278);
nand U24310 (N_24310,N_20287,N_20347);
or U24311 (N_24311,N_20709,N_20120);
nor U24312 (N_24312,N_18974,N_20912);
nor U24313 (N_24313,N_21173,N_20296);
nor U24314 (N_24314,N_21000,N_19227);
or U24315 (N_24315,N_19683,N_19053);
or U24316 (N_24316,N_19705,N_19317);
or U24317 (N_24317,N_19388,N_20769);
and U24318 (N_24318,N_18806,N_19511);
nand U24319 (N_24319,N_21250,N_20569);
xor U24320 (N_24320,N_21551,N_20137);
and U24321 (N_24321,N_20157,N_21188);
xor U24322 (N_24322,N_21722,N_19951);
nor U24323 (N_24323,N_18768,N_19060);
xnor U24324 (N_24324,N_21694,N_20939);
xor U24325 (N_24325,N_19485,N_21386);
and U24326 (N_24326,N_18944,N_19265);
nand U24327 (N_24327,N_21469,N_21012);
and U24328 (N_24328,N_21681,N_19089);
xnor U24329 (N_24329,N_20453,N_19470);
and U24330 (N_24330,N_19709,N_18911);
or U24331 (N_24331,N_18996,N_21245);
nor U24332 (N_24332,N_19630,N_19933);
and U24333 (N_24333,N_20748,N_20740);
xnor U24334 (N_24334,N_19667,N_20494);
xor U24335 (N_24335,N_21545,N_20471);
xnor U24336 (N_24336,N_19682,N_21503);
and U24337 (N_24337,N_21397,N_20123);
xnor U24338 (N_24338,N_20246,N_20883);
nand U24339 (N_24339,N_19879,N_21515);
nand U24340 (N_24340,N_21248,N_21241);
or U24341 (N_24341,N_20569,N_21802);
and U24342 (N_24342,N_19956,N_20399);
nand U24343 (N_24343,N_18765,N_20744);
or U24344 (N_24344,N_21029,N_21100);
nand U24345 (N_24345,N_20870,N_20644);
nand U24346 (N_24346,N_18931,N_20537);
and U24347 (N_24347,N_18914,N_19185);
nand U24348 (N_24348,N_20438,N_19810);
or U24349 (N_24349,N_20033,N_18798);
xnor U24350 (N_24350,N_18790,N_20226);
or U24351 (N_24351,N_21412,N_21789);
xor U24352 (N_24352,N_19869,N_21186);
nand U24353 (N_24353,N_19200,N_19418);
and U24354 (N_24354,N_20231,N_19187);
nor U24355 (N_24355,N_19623,N_20230);
or U24356 (N_24356,N_20513,N_20626);
nor U24357 (N_24357,N_21344,N_20303);
nand U24358 (N_24358,N_18939,N_19527);
nor U24359 (N_24359,N_19461,N_20694);
nand U24360 (N_24360,N_20218,N_20391);
nand U24361 (N_24361,N_20455,N_19647);
or U24362 (N_24362,N_21570,N_20393);
and U24363 (N_24363,N_21142,N_21828);
or U24364 (N_24364,N_18965,N_20011);
nor U24365 (N_24365,N_20071,N_21530);
or U24366 (N_24366,N_19511,N_19474);
xor U24367 (N_24367,N_19518,N_20446);
xnor U24368 (N_24368,N_20779,N_20503);
or U24369 (N_24369,N_21370,N_20871);
nor U24370 (N_24370,N_20925,N_19892);
nand U24371 (N_24371,N_19224,N_19573);
xnor U24372 (N_24372,N_21134,N_19658);
nor U24373 (N_24373,N_18854,N_20713);
nand U24374 (N_24374,N_20444,N_18866);
nand U24375 (N_24375,N_19134,N_18773);
xnor U24376 (N_24376,N_19219,N_20849);
xnor U24377 (N_24377,N_20329,N_19416);
and U24378 (N_24378,N_19199,N_19548);
or U24379 (N_24379,N_19198,N_21521);
or U24380 (N_24380,N_19301,N_19163);
nand U24381 (N_24381,N_21061,N_20905);
nand U24382 (N_24382,N_20771,N_21509);
and U24383 (N_24383,N_21811,N_20983);
or U24384 (N_24384,N_20490,N_21386);
nand U24385 (N_24385,N_21669,N_19749);
and U24386 (N_24386,N_19903,N_20231);
nor U24387 (N_24387,N_21793,N_21711);
xor U24388 (N_24388,N_19598,N_21312);
nand U24389 (N_24389,N_21469,N_19455);
xor U24390 (N_24390,N_20153,N_21189);
xor U24391 (N_24391,N_21608,N_21122);
and U24392 (N_24392,N_21230,N_19521);
and U24393 (N_24393,N_21303,N_20343);
or U24394 (N_24394,N_20205,N_20284);
nand U24395 (N_24395,N_19692,N_19404);
and U24396 (N_24396,N_20128,N_21013);
or U24397 (N_24397,N_20871,N_20099);
nor U24398 (N_24398,N_20154,N_21560);
or U24399 (N_24399,N_18828,N_20188);
or U24400 (N_24400,N_21320,N_20111);
or U24401 (N_24401,N_21654,N_19814);
nand U24402 (N_24402,N_21169,N_18769);
xor U24403 (N_24403,N_20996,N_21114);
or U24404 (N_24404,N_19998,N_20818);
nor U24405 (N_24405,N_19914,N_21353);
or U24406 (N_24406,N_19691,N_21776);
xor U24407 (N_24407,N_19935,N_18930);
and U24408 (N_24408,N_21365,N_21137);
nor U24409 (N_24409,N_21467,N_21487);
or U24410 (N_24410,N_21757,N_20786);
nand U24411 (N_24411,N_21495,N_20663);
and U24412 (N_24412,N_18804,N_21831);
or U24413 (N_24413,N_20387,N_20203);
and U24414 (N_24414,N_20624,N_19805);
or U24415 (N_24415,N_19867,N_19649);
xnor U24416 (N_24416,N_20303,N_20630);
nor U24417 (N_24417,N_20309,N_21730);
xor U24418 (N_24418,N_21677,N_19661);
xor U24419 (N_24419,N_21461,N_20106);
and U24420 (N_24420,N_21316,N_21334);
xor U24421 (N_24421,N_18902,N_20333);
nor U24422 (N_24422,N_20572,N_21635);
nor U24423 (N_24423,N_19148,N_20094);
nand U24424 (N_24424,N_19706,N_21433);
or U24425 (N_24425,N_21457,N_21377);
nand U24426 (N_24426,N_19800,N_20695);
nor U24427 (N_24427,N_20564,N_21700);
or U24428 (N_24428,N_19887,N_20853);
or U24429 (N_24429,N_18759,N_19673);
and U24430 (N_24430,N_21129,N_21021);
and U24431 (N_24431,N_19954,N_19748);
nor U24432 (N_24432,N_20140,N_21326);
and U24433 (N_24433,N_20457,N_21582);
or U24434 (N_24434,N_19509,N_18776);
nor U24435 (N_24435,N_20570,N_20142);
and U24436 (N_24436,N_19021,N_21325);
nor U24437 (N_24437,N_19946,N_21536);
nand U24438 (N_24438,N_18966,N_21601);
and U24439 (N_24439,N_21559,N_21432);
and U24440 (N_24440,N_20671,N_20158);
or U24441 (N_24441,N_19751,N_20492);
nor U24442 (N_24442,N_21233,N_19798);
nor U24443 (N_24443,N_21584,N_21308);
xnor U24444 (N_24444,N_20131,N_20586);
nand U24445 (N_24445,N_20216,N_21574);
and U24446 (N_24446,N_20417,N_19751);
nor U24447 (N_24447,N_19673,N_21764);
nand U24448 (N_24448,N_19117,N_20624);
and U24449 (N_24449,N_21644,N_20600);
nand U24450 (N_24450,N_21361,N_21856);
nand U24451 (N_24451,N_19903,N_21550);
or U24452 (N_24452,N_20729,N_20439);
nand U24453 (N_24453,N_19383,N_19660);
and U24454 (N_24454,N_21729,N_20596);
xor U24455 (N_24455,N_21716,N_20956);
nor U24456 (N_24456,N_21308,N_18797);
nand U24457 (N_24457,N_21769,N_21379);
nor U24458 (N_24458,N_20952,N_21081);
and U24459 (N_24459,N_20298,N_21493);
and U24460 (N_24460,N_21812,N_20224);
nand U24461 (N_24461,N_21218,N_20606);
and U24462 (N_24462,N_19760,N_19458);
and U24463 (N_24463,N_19714,N_18755);
xor U24464 (N_24464,N_21205,N_21527);
nand U24465 (N_24465,N_19021,N_19948);
and U24466 (N_24466,N_19925,N_21564);
or U24467 (N_24467,N_19321,N_21817);
nor U24468 (N_24468,N_19247,N_21413);
nor U24469 (N_24469,N_21121,N_19663);
nand U24470 (N_24470,N_20677,N_20917);
nor U24471 (N_24471,N_21867,N_20617);
or U24472 (N_24472,N_19061,N_21840);
or U24473 (N_24473,N_20936,N_19556);
or U24474 (N_24474,N_20192,N_21498);
or U24475 (N_24475,N_20685,N_20881);
nand U24476 (N_24476,N_19921,N_20068);
nand U24477 (N_24477,N_18805,N_19145);
or U24478 (N_24478,N_20421,N_20988);
xnor U24479 (N_24479,N_21171,N_20871);
nand U24480 (N_24480,N_21673,N_20105);
xor U24481 (N_24481,N_21669,N_19198);
or U24482 (N_24482,N_21851,N_21185);
xor U24483 (N_24483,N_21482,N_20145);
nand U24484 (N_24484,N_21591,N_21505);
xnor U24485 (N_24485,N_19277,N_20297);
nor U24486 (N_24486,N_21732,N_19593);
nor U24487 (N_24487,N_21113,N_20566);
nand U24488 (N_24488,N_18994,N_21223);
nand U24489 (N_24489,N_19281,N_21321);
nand U24490 (N_24490,N_19647,N_20769);
nor U24491 (N_24491,N_19154,N_19563);
nor U24492 (N_24492,N_20123,N_21159);
xnor U24493 (N_24493,N_20411,N_21241);
and U24494 (N_24494,N_20969,N_20429);
xor U24495 (N_24495,N_21836,N_21175);
and U24496 (N_24496,N_20680,N_20898);
nor U24497 (N_24497,N_20969,N_19074);
or U24498 (N_24498,N_19916,N_20279);
xor U24499 (N_24499,N_20027,N_20195);
nand U24500 (N_24500,N_19579,N_20082);
and U24501 (N_24501,N_21264,N_20390);
nand U24502 (N_24502,N_20747,N_20103);
xnor U24503 (N_24503,N_20959,N_19045);
xnor U24504 (N_24504,N_19818,N_21628);
nand U24505 (N_24505,N_19984,N_20400);
nor U24506 (N_24506,N_19210,N_20350);
nand U24507 (N_24507,N_21063,N_21306);
and U24508 (N_24508,N_19032,N_19229);
nor U24509 (N_24509,N_21222,N_21350);
xnor U24510 (N_24510,N_21593,N_20429);
or U24511 (N_24511,N_20540,N_21269);
nand U24512 (N_24512,N_21346,N_19593);
nor U24513 (N_24513,N_18992,N_21013);
and U24514 (N_24514,N_20869,N_18774);
or U24515 (N_24515,N_20250,N_19073);
nand U24516 (N_24516,N_21031,N_20774);
xnor U24517 (N_24517,N_21160,N_19285);
nand U24518 (N_24518,N_20031,N_21199);
xor U24519 (N_24519,N_19460,N_20855);
or U24520 (N_24520,N_18922,N_19632);
or U24521 (N_24521,N_19951,N_21760);
nor U24522 (N_24522,N_19680,N_19547);
or U24523 (N_24523,N_18896,N_21578);
xnor U24524 (N_24524,N_20831,N_19083);
and U24525 (N_24525,N_20746,N_19419);
and U24526 (N_24526,N_20862,N_21257);
or U24527 (N_24527,N_18976,N_21455);
nand U24528 (N_24528,N_21816,N_20381);
or U24529 (N_24529,N_20640,N_20864);
nor U24530 (N_24530,N_19525,N_20958);
nand U24531 (N_24531,N_19725,N_19350);
xnor U24532 (N_24532,N_21742,N_19880);
and U24533 (N_24533,N_21569,N_20542);
nor U24534 (N_24534,N_20465,N_20156);
xnor U24535 (N_24535,N_20823,N_19721);
xor U24536 (N_24536,N_19562,N_21368);
or U24537 (N_24537,N_20650,N_18999);
xor U24538 (N_24538,N_19979,N_19585);
and U24539 (N_24539,N_19857,N_20449);
or U24540 (N_24540,N_20049,N_21576);
and U24541 (N_24541,N_19597,N_20730);
xnor U24542 (N_24542,N_20860,N_21351);
xor U24543 (N_24543,N_19397,N_21838);
and U24544 (N_24544,N_19760,N_21512);
or U24545 (N_24545,N_20677,N_21367);
xnor U24546 (N_24546,N_20093,N_19810);
nor U24547 (N_24547,N_20160,N_20124);
nand U24548 (N_24548,N_21332,N_21121);
nor U24549 (N_24549,N_19555,N_21781);
nor U24550 (N_24550,N_21195,N_19599);
xor U24551 (N_24551,N_21727,N_21668);
nor U24552 (N_24552,N_21797,N_20733);
and U24553 (N_24553,N_21491,N_19229);
and U24554 (N_24554,N_20000,N_18956);
nand U24555 (N_24555,N_18835,N_20587);
nand U24556 (N_24556,N_21749,N_20181);
xor U24557 (N_24557,N_21618,N_20370);
and U24558 (N_24558,N_19687,N_20119);
xnor U24559 (N_24559,N_19354,N_19536);
and U24560 (N_24560,N_20419,N_19792);
or U24561 (N_24561,N_19449,N_21238);
xnor U24562 (N_24562,N_21130,N_21280);
xnor U24563 (N_24563,N_21541,N_18915);
and U24564 (N_24564,N_19399,N_20823);
nor U24565 (N_24565,N_21392,N_19194);
nor U24566 (N_24566,N_21749,N_20125);
or U24567 (N_24567,N_19244,N_20275);
xor U24568 (N_24568,N_18756,N_20314);
or U24569 (N_24569,N_21424,N_21632);
xnor U24570 (N_24570,N_21289,N_19675);
nor U24571 (N_24571,N_19708,N_20676);
nor U24572 (N_24572,N_20662,N_19415);
nor U24573 (N_24573,N_19395,N_19677);
and U24574 (N_24574,N_21016,N_20161);
and U24575 (N_24575,N_19498,N_21145);
xnor U24576 (N_24576,N_19535,N_21784);
or U24577 (N_24577,N_19148,N_20900);
or U24578 (N_24578,N_20969,N_19295);
nand U24579 (N_24579,N_20587,N_20304);
or U24580 (N_24580,N_21785,N_19091);
and U24581 (N_24581,N_19106,N_21703);
and U24582 (N_24582,N_20904,N_18751);
xor U24583 (N_24583,N_19298,N_21608);
or U24584 (N_24584,N_21507,N_20828);
or U24585 (N_24585,N_18931,N_18870);
and U24586 (N_24586,N_20603,N_20845);
nor U24587 (N_24587,N_19991,N_20112);
and U24588 (N_24588,N_21194,N_21125);
xor U24589 (N_24589,N_19307,N_20307);
xor U24590 (N_24590,N_19212,N_18876);
xor U24591 (N_24591,N_21653,N_20860);
and U24592 (N_24592,N_21829,N_20737);
or U24593 (N_24593,N_19527,N_20925);
nor U24594 (N_24594,N_19870,N_18909);
nand U24595 (N_24595,N_19979,N_19277);
nand U24596 (N_24596,N_19543,N_20740);
or U24597 (N_24597,N_21261,N_21198);
and U24598 (N_24598,N_20329,N_19150);
nor U24599 (N_24599,N_20853,N_19776);
nor U24600 (N_24600,N_21792,N_19390);
xnor U24601 (N_24601,N_19620,N_20422);
and U24602 (N_24602,N_19292,N_21175);
nand U24603 (N_24603,N_18774,N_21597);
or U24604 (N_24604,N_21244,N_19436);
nand U24605 (N_24605,N_20569,N_19713);
xor U24606 (N_24606,N_21177,N_19340);
and U24607 (N_24607,N_21587,N_20700);
or U24608 (N_24608,N_19275,N_21285);
or U24609 (N_24609,N_19649,N_20369);
and U24610 (N_24610,N_19033,N_19101);
nor U24611 (N_24611,N_21219,N_18756);
nor U24612 (N_24612,N_20909,N_21666);
nand U24613 (N_24613,N_20627,N_19278);
nand U24614 (N_24614,N_20115,N_19744);
nand U24615 (N_24615,N_19724,N_20661);
and U24616 (N_24616,N_18849,N_21393);
nand U24617 (N_24617,N_21146,N_20275);
xnor U24618 (N_24618,N_19541,N_19116);
nor U24619 (N_24619,N_19666,N_20843);
and U24620 (N_24620,N_20926,N_19828);
or U24621 (N_24621,N_21577,N_19519);
and U24622 (N_24622,N_18829,N_21331);
nor U24623 (N_24623,N_21622,N_19229);
or U24624 (N_24624,N_21037,N_21177);
xnor U24625 (N_24625,N_19537,N_20107);
nand U24626 (N_24626,N_19025,N_19491);
nor U24627 (N_24627,N_18802,N_19593);
and U24628 (N_24628,N_20074,N_20647);
xnor U24629 (N_24629,N_20049,N_19728);
nand U24630 (N_24630,N_21429,N_21336);
nand U24631 (N_24631,N_21504,N_19725);
and U24632 (N_24632,N_19367,N_19714);
nand U24633 (N_24633,N_21300,N_21057);
nand U24634 (N_24634,N_21582,N_20572);
or U24635 (N_24635,N_21374,N_20042);
or U24636 (N_24636,N_20375,N_18754);
or U24637 (N_24637,N_19526,N_18751);
nor U24638 (N_24638,N_19856,N_20292);
nand U24639 (N_24639,N_21482,N_19079);
nand U24640 (N_24640,N_20132,N_21441);
nand U24641 (N_24641,N_19890,N_20711);
nor U24642 (N_24642,N_19424,N_19169);
xor U24643 (N_24643,N_18958,N_21599);
or U24644 (N_24644,N_21555,N_20266);
or U24645 (N_24645,N_21857,N_20259);
xnor U24646 (N_24646,N_19307,N_19306);
xor U24647 (N_24647,N_19460,N_21109);
xnor U24648 (N_24648,N_19543,N_21387);
xnor U24649 (N_24649,N_18955,N_19630);
nor U24650 (N_24650,N_20294,N_21312);
or U24651 (N_24651,N_19707,N_19827);
xnor U24652 (N_24652,N_19320,N_18805);
xor U24653 (N_24653,N_20565,N_20973);
xnor U24654 (N_24654,N_21636,N_19789);
nand U24655 (N_24655,N_19037,N_19554);
and U24656 (N_24656,N_21678,N_19328);
or U24657 (N_24657,N_21019,N_18994);
nand U24658 (N_24658,N_19714,N_20097);
nor U24659 (N_24659,N_19798,N_19289);
nor U24660 (N_24660,N_21284,N_18915);
xnor U24661 (N_24661,N_21601,N_19600);
nor U24662 (N_24662,N_20666,N_21019);
nand U24663 (N_24663,N_21046,N_20136);
xor U24664 (N_24664,N_19968,N_19930);
nand U24665 (N_24665,N_19285,N_20252);
nor U24666 (N_24666,N_19815,N_18769);
nand U24667 (N_24667,N_19264,N_18767);
and U24668 (N_24668,N_21070,N_20253);
nor U24669 (N_24669,N_21566,N_19333);
xor U24670 (N_24670,N_21095,N_21744);
or U24671 (N_24671,N_20191,N_20980);
nand U24672 (N_24672,N_19844,N_19876);
nor U24673 (N_24673,N_20112,N_19911);
xnor U24674 (N_24674,N_19029,N_20834);
and U24675 (N_24675,N_20280,N_20338);
nand U24676 (N_24676,N_19495,N_21181);
nand U24677 (N_24677,N_20294,N_19762);
and U24678 (N_24678,N_21344,N_19522);
nand U24679 (N_24679,N_21843,N_21050);
xor U24680 (N_24680,N_20934,N_19664);
xor U24681 (N_24681,N_21473,N_20241);
or U24682 (N_24682,N_19442,N_18937);
nand U24683 (N_24683,N_21399,N_19134);
nor U24684 (N_24684,N_19056,N_20767);
xor U24685 (N_24685,N_19868,N_19375);
nand U24686 (N_24686,N_21608,N_21801);
nand U24687 (N_24687,N_19890,N_19051);
xnor U24688 (N_24688,N_21654,N_19289);
nor U24689 (N_24689,N_20695,N_19580);
nand U24690 (N_24690,N_21461,N_20373);
and U24691 (N_24691,N_20805,N_21609);
nand U24692 (N_24692,N_19941,N_20630);
or U24693 (N_24693,N_21586,N_20122);
and U24694 (N_24694,N_20554,N_18755);
and U24695 (N_24695,N_20468,N_21222);
and U24696 (N_24696,N_21418,N_21829);
or U24697 (N_24697,N_19653,N_20758);
and U24698 (N_24698,N_19669,N_19311);
xnor U24699 (N_24699,N_20478,N_21872);
xnor U24700 (N_24700,N_20745,N_20532);
xor U24701 (N_24701,N_21751,N_20096);
xor U24702 (N_24702,N_20398,N_19590);
or U24703 (N_24703,N_19609,N_19604);
nand U24704 (N_24704,N_19051,N_20647);
nand U24705 (N_24705,N_21446,N_20769);
nor U24706 (N_24706,N_19861,N_21136);
or U24707 (N_24707,N_21679,N_20802);
nor U24708 (N_24708,N_20189,N_19068);
nand U24709 (N_24709,N_20496,N_19615);
and U24710 (N_24710,N_20007,N_21103);
or U24711 (N_24711,N_20062,N_20495);
or U24712 (N_24712,N_19823,N_18803);
and U24713 (N_24713,N_21225,N_21656);
xnor U24714 (N_24714,N_20672,N_20586);
nor U24715 (N_24715,N_19065,N_18951);
and U24716 (N_24716,N_19293,N_18998);
and U24717 (N_24717,N_19558,N_21320);
nand U24718 (N_24718,N_19738,N_20638);
and U24719 (N_24719,N_20386,N_21236);
xor U24720 (N_24720,N_21773,N_19863);
or U24721 (N_24721,N_21233,N_18864);
xor U24722 (N_24722,N_21036,N_19500);
xor U24723 (N_24723,N_20449,N_21610);
and U24724 (N_24724,N_19339,N_18758);
nor U24725 (N_24725,N_21699,N_20404);
or U24726 (N_24726,N_20766,N_21724);
and U24727 (N_24727,N_19931,N_20344);
and U24728 (N_24728,N_19028,N_20006);
nor U24729 (N_24729,N_19089,N_20413);
and U24730 (N_24730,N_21718,N_20525);
nor U24731 (N_24731,N_20722,N_18798);
nor U24732 (N_24732,N_19407,N_21011);
or U24733 (N_24733,N_19368,N_20691);
and U24734 (N_24734,N_21588,N_19305);
nor U24735 (N_24735,N_20411,N_19497);
nand U24736 (N_24736,N_18798,N_19189);
nand U24737 (N_24737,N_19616,N_21343);
xor U24738 (N_24738,N_21290,N_21812);
nor U24739 (N_24739,N_20534,N_21754);
nand U24740 (N_24740,N_18946,N_21826);
xor U24741 (N_24741,N_19492,N_21124);
or U24742 (N_24742,N_19348,N_18911);
or U24743 (N_24743,N_20082,N_20072);
nor U24744 (N_24744,N_20005,N_21127);
nor U24745 (N_24745,N_20576,N_20739);
nand U24746 (N_24746,N_20754,N_20587);
and U24747 (N_24747,N_20412,N_20267);
nor U24748 (N_24748,N_21376,N_19132);
nand U24749 (N_24749,N_21639,N_20403);
or U24750 (N_24750,N_19443,N_21106);
xor U24751 (N_24751,N_20175,N_18936);
nor U24752 (N_24752,N_20040,N_20581);
or U24753 (N_24753,N_19515,N_19137);
nor U24754 (N_24754,N_21051,N_20660);
and U24755 (N_24755,N_19178,N_19715);
or U24756 (N_24756,N_21726,N_21418);
xor U24757 (N_24757,N_20123,N_19672);
or U24758 (N_24758,N_20007,N_19016);
and U24759 (N_24759,N_21139,N_21827);
and U24760 (N_24760,N_18895,N_21198);
nor U24761 (N_24761,N_19863,N_20951);
nor U24762 (N_24762,N_18893,N_21738);
or U24763 (N_24763,N_20328,N_19258);
nand U24764 (N_24764,N_19447,N_21659);
nor U24765 (N_24765,N_21190,N_21637);
nand U24766 (N_24766,N_20310,N_21737);
and U24767 (N_24767,N_19121,N_19726);
xnor U24768 (N_24768,N_21198,N_20397);
xnor U24769 (N_24769,N_19066,N_20623);
nor U24770 (N_24770,N_21607,N_19068);
nand U24771 (N_24771,N_20501,N_21464);
nor U24772 (N_24772,N_21814,N_20366);
and U24773 (N_24773,N_21064,N_21342);
and U24774 (N_24774,N_21425,N_20277);
nand U24775 (N_24775,N_21724,N_21758);
or U24776 (N_24776,N_18862,N_21461);
or U24777 (N_24777,N_20906,N_19529);
and U24778 (N_24778,N_18932,N_19002);
xnor U24779 (N_24779,N_21258,N_20062);
and U24780 (N_24780,N_20145,N_21443);
and U24781 (N_24781,N_21575,N_19726);
nand U24782 (N_24782,N_19045,N_19165);
or U24783 (N_24783,N_19570,N_21464);
xnor U24784 (N_24784,N_19244,N_19517);
and U24785 (N_24785,N_19957,N_19693);
nand U24786 (N_24786,N_20886,N_20819);
and U24787 (N_24787,N_18876,N_20557);
nor U24788 (N_24788,N_21203,N_18973);
nor U24789 (N_24789,N_20661,N_18999);
and U24790 (N_24790,N_18979,N_20386);
and U24791 (N_24791,N_20941,N_20057);
xnor U24792 (N_24792,N_18765,N_19871);
nor U24793 (N_24793,N_21870,N_21754);
and U24794 (N_24794,N_21388,N_21741);
or U24795 (N_24795,N_20977,N_19399);
or U24796 (N_24796,N_20942,N_19971);
and U24797 (N_24797,N_20941,N_21702);
nor U24798 (N_24798,N_21833,N_20203);
xnor U24799 (N_24799,N_21027,N_19893);
nor U24800 (N_24800,N_21467,N_20710);
or U24801 (N_24801,N_19155,N_21754);
nor U24802 (N_24802,N_21280,N_20610);
and U24803 (N_24803,N_18945,N_20738);
nor U24804 (N_24804,N_20863,N_20357);
or U24805 (N_24805,N_19066,N_20649);
or U24806 (N_24806,N_20851,N_21120);
nand U24807 (N_24807,N_20988,N_21143);
nand U24808 (N_24808,N_20952,N_19660);
nor U24809 (N_24809,N_20780,N_20640);
xnor U24810 (N_24810,N_21768,N_20704);
xnor U24811 (N_24811,N_19994,N_20181);
xor U24812 (N_24812,N_21625,N_21859);
xor U24813 (N_24813,N_18773,N_20079);
nand U24814 (N_24814,N_19554,N_21291);
nor U24815 (N_24815,N_18801,N_18849);
and U24816 (N_24816,N_20028,N_19184);
nor U24817 (N_24817,N_19790,N_20488);
or U24818 (N_24818,N_19246,N_19243);
xor U24819 (N_24819,N_20779,N_20397);
nand U24820 (N_24820,N_19427,N_20899);
xnor U24821 (N_24821,N_21245,N_18847);
and U24822 (N_24822,N_21009,N_19428);
xor U24823 (N_24823,N_19972,N_20354);
xnor U24824 (N_24824,N_20527,N_21059);
and U24825 (N_24825,N_18973,N_19889);
nor U24826 (N_24826,N_20996,N_20040);
xnor U24827 (N_24827,N_20573,N_20007);
nand U24828 (N_24828,N_19828,N_20051);
nor U24829 (N_24829,N_20754,N_20696);
or U24830 (N_24830,N_18949,N_19321);
xor U24831 (N_24831,N_20804,N_21490);
and U24832 (N_24832,N_19944,N_20505);
or U24833 (N_24833,N_19481,N_21667);
nor U24834 (N_24834,N_19834,N_20601);
nor U24835 (N_24835,N_19676,N_21484);
or U24836 (N_24836,N_21732,N_19705);
and U24837 (N_24837,N_19975,N_21693);
nand U24838 (N_24838,N_19993,N_19959);
nor U24839 (N_24839,N_19195,N_21693);
xor U24840 (N_24840,N_18929,N_21782);
nand U24841 (N_24841,N_19739,N_20818);
nand U24842 (N_24842,N_20481,N_20114);
or U24843 (N_24843,N_20694,N_20836);
nor U24844 (N_24844,N_19334,N_19530);
xnor U24845 (N_24845,N_19619,N_21814);
or U24846 (N_24846,N_20924,N_21007);
xnor U24847 (N_24847,N_18895,N_21402);
and U24848 (N_24848,N_19559,N_19984);
or U24849 (N_24849,N_19904,N_21297);
nand U24850 (N_24850,N_18802,N_19591);
nand U24851 (N_24851,N_20537,N_18799);
or U24852 (N_24852,N_21678,N_21260);
or U24853 (N_24853,N_20946,N_21401);
or U24854 (N_24854,N_21787,N_19394);
nor U24855 (N_24855,N_18750,N_20535);
xor U24856 (N_24856,N_20440,N_20574);
nor U24857 (N_24857,N_21093,N_21740);
and U24858 (N_24858,N_20118,N_19052);
nand U24859 (N_24859,N_19077,N_20958);
or U24860 (N_24860,N_19024,N_19794);
nor U24861 (N_24861,N_18950,N_18903);
nand U24862 (N_24862,N_19728,N_21419);
xnor U24863 (N_24863,N_20665,N_20582);
xnor U24864 (N_24864,N_19603,N_20556);
nand U24865 (N_24865,N_20941,N_21687);
xor U24866 (N_24866,N_19436,N_21565);
or U24867 (N_24867,N_18936,N_20086);
and U24868 (N_24868,N_19362,N_19779);
nand U24869 (N_24869,N_19246,N_19841);
nor U24870 (N_24870,N_18927,N_21310);
or U24871 (N_24871,N_20840,N_19065);
nand U24872 (N_24872,N_19747,N_21573);
xnor U24873 (N_24873,N_19760,N_19143);
and U24874 (N_24874,N_19615,N_18940);
nand U24875 (N_24875,N_18779,N_19128);
or U24876 (N_24876,N_19183,N_20366);
nand U24877 (N_24877,N_19025,N_19887);
and U24878 (N_24878,N_20241,N_21415);
nand U24879 (N_24879,N_18937,N_18905);
nor U24880 (N_24880,N_21686,N_20818);
or U24881 (N_24881,N_20897,N_19386);
xnor U24882 (N_24882,N_20064,N_19617);
or U24883 (N_24883,N_20850,N_19262);
nand U24884 (N_24884,N_20631,N_19931);
nand U24885 (N_24885,N_21150,N_19755);
and U24886 (N_24886,N_19754,N_20672);
nor U24887 (N_24887,N_19001,N_21205);
xor U24888 (N_24888,N_20855,N_19334);
nand U24889 (N_24889,N_21259,N_21086);
or U24890 (N_24890,N_20701,N_20204);
xor U24891 (N_24891,N_20486,N_21037);
or U24892 (N_24892,N_19374,N_20987);
and U24893 (N_24893,N_19633,N_19156);
nand U24894 (N_24894,N_21618,N_19821);
nor U24895 (N_24895,N_18825,N_18997);
and U24896 (N_24896,N_19861,N_19893);
and U24897 (N_24897,N_21271,N_21874);
nor U24898 (N_24898,N_19979,N_20420);
nand U24899 (N_24899,N_19529,N_19440);
nand U24900 (N_24900,N_20844,N_19913);
or U24901 (N_24901,N_21320,N_20675);
nor U24902 (N_24902,N_20917,N_20838);
or U24903 (N_24903,N_18967,N_19584);
and U24904 (N_24904,N_18957,N_20743);
xnor U24905 (N_24905,N_19950,N_19801);
or U24906 (N_24906,N_19949,N_20378);
or U24907 (N_24907,N_19343,N_19278);
and U24908 (N_24908,N_20380,N_21106);
nor U24909 (N_24909,N_19252,N_21237);
or U24910 (N_24910,N_18970,N_18920);
nand U24911 (N_24911,N_21124,N_19747);
and U24912 (N_24912,N_20993,N_20865);
xor U24913 (N_24913,N_19868,N_19570);
or U24914 (N_24914,N_18856,N_20190);
or U24915 (N_24915,N_21751,N_19052);
or U24916 (N_24916,N_18893,N_19400);
nand U24917 (N_24917,N_21749,N_18992);
or U24918 (N_24918,N_21426,N_19119);
nor U24919 (N_24919,N_18862,N_21250);
xnor U24920 (N_24920,N_19404,N_21154);
xor U24921 (N_24921,N_21857,N_18922);
and U24922 (N_24922,N_21561,N_19885);
nand U24923 (N_24923,N_21702,N_19813);
xor U24924 (N_24924,N_19968,N_18755);
xnor U24925 (N_24925,N_20274,N_20576);
and U24926 (N_24926,N_21716,N_20760);
or U24927 (N_24927,N_20556,N_20001);
or U24928 (N_24928,N_19252,N_18789);
nand U24929 (N_24929,N_19194,N_18810);
nand U24930 (N_24930,N_18934,N_20724);
nor U24931 (N_24931,N_20037,N_19768);
or U24932 (N_24932,N_19464,N_21169);
xor U24933 (N_24933,N_21374,N_19798);
nand U24934 (N_24934,N_19821,N_19893);
and U24935 (N_24935,N_19640,N_20551);
or U24936 (N_24936,N_18858,N_20919);
and U24937 (N_24937,N_19195,N_21091);
and U24938 (N_24938,N_19142,N_21153);
xor U24939 (N_24939,N_21544,N_19763);
or U24940 (N_24940,N_20840,N_20180);
nand U24941 (N_24941,N_21625,N_19795);
nand U24942 (N_24942,N_19243,N_19075);
nand U24943 (N_24943,N_19345,N_20601);
xor U24944 (N_24944,N_19972,N_20013);
xor U24945 (N_24945,N_20590,N_18808);
nand U24946 (N_24946,N_19405,N_20570);
and U24947 (N_24947,N_20117,N_20465);
or U24948 (N_24948,N_20472,N_21208);
xnor U24949 (N_24949,N_19050,N_21231);
xnor U24950 (N_24950,N_19041,N_20131);
xor U24951 (N_24951,N_19397,N_21584);
xor U24952 (N_24952,N_20436,N_21526);
nand U24953 (N_24953,N_21823,N_18838);
and U24954 (N_24954,N_19264,N_18758);
nor U24955 (N_24955,N_21485,N_19719);
nand U24956 (N_24956,N_20117,N_18936);
nor U24957 (N_24957,N_20579,N_20426);
and U24958 (N_24958,N_19538,N_20849);
or U24959 (N_24959,N_21036,N_20875);
nand U24960 (N_24960,N_21103,N_20828);
or U24961 (N_24961,N_20795,N_20790);
or U24962 (N_24962,N_21531,N_19073);
nand U24963 (N_24963,N_19191,N_20431);
or U24964 (N_24964,N_19738,N_20200);
nor U24965 (N_24965,N_20562,N_20269);
nor U24966 (N_24966,N_19956,N_19708);
and U24967 (N_24967,N_21387,N_20581);
and U24968 (N_24968,N_21763,N_19071);
and U24969 (N_24969,N_19978,N_21683);
nor U24970 (N_24970,N_21840,N_19300);
xor U24971 (N_24971,N_21122,N_21813);
nand U24972 (N_24972,N_19470,N_19122);
nor U24973 (N_24973,N_20868,N_20309);
and U24974 (N_24974,N_19711,N_20108);
or U24975 (N_24975,N_21652,N_19727);
nand U24976 (N_24976,N_20836,N_20469);
xor U24977 (N_24977,N_20797,N_18883);
or U24978 (N_24978,N_20978,N_19802);
and U24979 (N_24979,N_18960,N_21380);
and U24980 (N_24980,N_21138,N_21401);
and U24981 (N_24981,N_21198,N_19191);
and U24982 (N_24982,N_18759,N_19008);
nand U24983 (N_24983,N_21755,N_21873);
and U24984 (N_24984,N_20488,N_19837);
nand U24985 (N_24985,N_19462,N_20754);
nand U24986 (N_24986,N_20061,N_20917);
xor U24987 (N_24987,N_21418,N_20752);
nor U24988 (N_24988,N_20358,N_18872);
xor U24989 (N_24989,N_21324,N_20026);
nor U24990 (N_24990,N_19925,N_19554);
or U24991 (N_24991,N_20149,N_21792);
nand U24992 (N_24992,N_19681,N_21085);
nor U24993 (N_24993,N_20607,N_18921);
nand U24994 (N_24994,N_21640,N_21063);
nand U24995 (N_24995,N_20502,N_20962);
and U24996 (N_24996,N_20030,N_19681);
xnor U24997 (N_24997,N_20350,N_20502);
nand U24998 (N_24998,N_21868,N_18830);
nand U24999 (N_24999,N_19733,N_21361);
and UO_0 (O_0,N_23758,N_24420);
nor UO_1 (O_1,N_22642,N_23330);
xor UO_2 (O_2,N_22495,N_23986);
and UO_3 (O_3,N_23731,N_21915);
nand UO_4 (O_4,N_24166,N_23005);
or UO_5 (O_5,N_23034,N_24544);
nand UO_6 (O_6,N_23571,N_24954);
nor UO_7 (O_7,N_22652,N_23805);
and UO_8 (O_8,N_22364,N_23182);
nand UO_9 (O_9,N_24724,N_22812);
and UO_10 (O_10,N_23595,N_24072);
and UO_11 (O_11,N_24964,N_23056);
or UO_12 (O_12,N_23911,N_23853);
xor UO_13 (O_13,N_22456,N_22749);
nand UO_14 (O_14,N_21913,N_24806);
xor UO_15 (O_15,N_22391,N_23055);
xor UO_16 (O_16,N_24585,N_24674);
or UO_17 (O_17,N_22727,N_24981);
and UO_18 (O_18,N_23541,N_23059);
nor UO_19 (O_19,N_23052,N_23438);
xor UO_20 (O_20,N_22855,N_22143);
and UO_21 (O_21,N_23638,N_22207);
nand UO_22 (O_22,N_23550,N_23905);
or UO_23 (O_23,N_22880,N_24345);
nand UO_24 (O_24,N_23944,N_24989);
and UO_25 (O_25,N_23299,N_23914);
or UO_26 (O_26,N_23185,N_23174);
and UO_27 (O_27,N_23763,N_22296);
and UO_28 (O_28,N_21950,N_22966);
nor UO_29 (O_29,N_24628,N_24975);
xnor UO_30 (O_30,N_23564,N_21953);
nor UO_31 (O_31,N_22424,N_24137);
nand UO_32 (O_32,N_24060,N_22845);
nand UO_33 (O_33,N_23077,N_24566);
xnor UO_34 (O_34,N_23753,N_23628);
xor UO_35 (O_35,N_22586,N_23768);
nand UO_36 (O_36,N_23012,N_22649);
nand UO_37 (O_37,N_23384,N_24050);
or UO_38 (O_38,N_23793,N_23149);
or UO_39 (O_39,N_24064,N_23388);
and UO_40 (O_40,N_22940,N_23367);
nand UO_41 (O_41,N_23007,N_22598);
and UO_42 (O_42,N_22362,N_23560);
xor UO_43 (O_43,N_24646,N_24071);
or UO_44 (O_44,N_22538,N_24282);
xnor UO_45 (O_45,N_24667,N_23206);
nor UO_46 (O_46,N_23436,N_22129);
xnor UO_47 (O_47,N_23127,N_23457);
and UO_48 (O_48,N_22286,N_23410);
xor UO_49 (O_49,N_23476,N_23485);
xor UO_50 (O_50,N_22071,N_24961);
and UO_51 (O_51,N_22146,N_24540);
nor UO_52 (O_52,N_21992,N_23265);
nand UO_53 (O_53,N_24762,N_22228);
nand UO_54 (O_54,N_24985,N_24398);
nand UO_55 (O_55,N_23930,N_22587);
nand UO_56 (O_56,N_22779,N_22202);
and UO_57 (O_57,N_24407,N_22405);
xnor UO_58 (O_58,N_22144,N_24347);
xnor UO_59 (O_59,N_23281,N_23808);
nand UO_60 (O_60,N_24133,N_22870);
xor UO_61 (O_61,N_21885,N_24506);
xor UO_62 (O_62,N_21927,N_22445);
and UO_63 (O_63,N_23501,N_23420);
nor UO_64 (O_64,N_24098,N_23656);
xnor UO_65 (O_65,N_24717,N_24059);
nand UO_66 (O_66,N_22250,N_22795);
and UO_67 (O_67,N_23667,N_23834);
nand UO_68 (O_68,N_23841,N_21975);
or UO_69 (O_69,N_24002,N_24163);
xor UO_70 (O_70,N_24690,N_23067);
or UO_71 (O_71,N_22962,N_22523);
xor UO_72 (O_72,N_22656,N_21881);
nor UO_73 (O_73,N_22086,N_22367);
nand UO_74 (O_74,N_24586,N_22638);
or UO_75 (O_75,N_23633,N_22684);
nand UO_76 (O_76,N_24545,N_24533);
or UO_77 (O_77,N_24156,N_24221);
xnor UO_78 (O_78,N_23934,N_23035);
nor UO_79 (O_79,N_22515,N_22145);
and UO_80 (O_80,N_23402,N_21890);
nand UO_81 (O_81,N_24031,N_21978);
nand UO_82 (O_82,N_24634,N_24534);
or UO_83 (O_83,N_21967,N_22050);
or UO_84 (O_84,N_24754,N_22725);
xnor UO_85 (O_85,N_23215,N_23585);
xor UO_86 (O_86,N_24310,N_24388);
nor UO_87 (O_87,N_22470,N_22458);
xor UO_88 (O_88,N_24291,N_24704);
nand UO_89 (O_89,N_22002,N_22699);
nand UO_90 (O_90,N_24154,N_22119);
xnor UO_91 (O_91,N_21990,N_23849);
xnor UO_92 (O_92,N_22361,N_24307);
nand UO_93 (O_93,N_22011,N_24945);
or UO_94 (O_94,N_23458,N_23788);
nand UO_95 (O_95,N_24439,N_22890);
and UO_96 (O_96,N_22745,N_22629);
or UO_97 (O_97,N_24449,N_24063);
nand UO_98 (O_98,N_23648,N_22401);
or UO_99 (O_99,N_23961,N_24573);
nand UO_100 (O_100,N_22720,N_23704);
xor UO_101 (O_101,N_24035,N_24253);
xnor UO_102 (O_102,N_22072,N_23061);
and UO_103 (O_103,N_22078,N_23023);
nor UO_104 (O_104,N_23379,N_23529);
xor UO_105 (O_105,N_23838,N_24250);
nand UO_106 (O_106,N_22517,N_24913);
nand UO_107 (O_107,N_23223,N_23686);
nor UO_108 (O_108,N_23707,N_24097);
xor UO_109 (O_109,N_23785,N_23176);
or UO_110 (O_110,N_23576,N_24316);
xor UO_111 (O_111,N_22904,N_24238);
and UO_112 (O_112,N_23732,N_24707);
xnor UO_113 (O_113,N_23448,N_24065);
xnor UO_114 (O_114,N_22199,N_24530);
nand UO_115 (O_115,N_24782,N_23407);
and UO_116 (O_116,N_24180,N_23578);
xor UO_117 (O_117,N_22167,N_24504);
nand UO_118 (O_118,N_24361,N_24962);
xor UO_119 (O_119,N_23714,N_24411);
or UO_120 (O_120,N_24046,N_24124);
or UO_121 (O_121,N_22178,N_23664);
and UO_122 (O_122,N_24592,N_23486);
nor UO_123 (O_123,N_24054,N_24703);
or UO_124 (O_124,N_22349,N_23635);
nor UO_125 (O_125,N_21970,N_22866);
xnor UO_126 (O_126,N_22980,N_24798);
nor UO_127 (O_127,N_22925,N_24326);
nand UO_128 (O_128,N_23974,N_22780);
nor UO_129 (O_129,N_22848,N_23075);
xor UO_130 (O_130,N_23693,N_22007);
and UO_131 (O_131,N_23722,N_23397);
or UO_132 (O_132,N_22793,N_23926);
nand UO_133 (O_133,N_24429,N_22112);
nor UO_134 (O_134,N_23818,N_23324);
nand UO_135 (O_135,N_22266,N_23734);
xor UO_136 (O_136,N_22110,N_23290);
nor UO_137 (O_137,N_24229,N_24480);
and UO_138 (O_138,N_22216,N_22645);
nand UO_139 (O_139,N_22746,N_22448);
and UO_140 (O_140,N_21875,N_24344);
and UO_141 (O_141,N_22528,N_23196);
and UO_142 (O_142,N_24753,N_23041);
xnor UO_143 (O_143,N_22956,N_22481);
xnor UO_144 (O_144,N_22691,N_24632);
nor UO_145 (O_145,N_22951,N_24218);
or UO_146 (O_146,N_23165,N_22695);
or UO_147 (O_147,N_23230,N_24893);
and UO_148 (O_148,N_23499,N_22839);
nand UO_149 (O_149,N_23243,N_22103);
xor UO_150 (O_150,N_21930,N_22338);
or UO_151 (O_151,N_23001,N_24817);
nand UO_152 (O_152,N_24616,N_24720);
nor UO_153 (O_153,N_23902,N_24744);
or UO_154 (O_154,N_22700,N_24998);
nor UO_155 (O_155,N_22898,N_22952);
xnor UO_156 (O_156,N_24702,N_22541);
or UO_157 (O_157,N_22460,N_22196);
xnor UO_158 (O_158,N_22504,N_24286);
xnor UO_159 (O_159,N_22408,N_24321);
xor UO_160 (O_160,N_24612,N_22045);
nand UO_161 (O_161,N_23432,N_24080);
and UO_162 (O_162,N_23952,N_24094);
nand UO_163 (O_163,N_22234,N_24805);
nand UO_164 (O_164,N_23452,N_22217);
or UO_165 (O_165,N_24808,N_24313);
or UO_166 (O_166,N_23478,N_24131);
or UO_167 (O_167,N_23446,N_24416);
or UO_168 (O_168,N_22844,N_22084);
and UO_169 (O_169,N_23355,N_22578);
nor UO_170 (O_170,N_22814,N_24173);
xor UO_171 (O_171,N_22469,N_24390);
nor UO_172 (O_172,N_24866,N_23396);
nor UO_173 (O_173,N_24652,N_24430);
and UO_174 (O_174,N_22923,N_22859);
xor UO_175 (O_175,N_22612,N_22766);
nor UO_176 (O_176,N_23235,N_23237);
nor UO_177 (O_177,N_22059,N_22789);
and UO_178 (O_178,N_24539,N_24887);
nand UO_179 (O_179,N_21986,N_23385);
or UO_180 (O_180,N_24497,N_22000);
xor UO_181 (O_181,N_24719,N_23147);
nor UO_182 (O_182,N_21982,N_22183);
and UO_183 (O_183,N_23445,N_24742);
xor UO_184 (O_184,N_24120,N_23749);
xnor UO_185 (O_185,N_24109,N_22139);
nor UO_186 (O_186,N_22534,N_24148);
nor UO_187 (O_187,N_22556,N_21880);
xnor UO_188 (O_188,N_24264,N_22466);
xor UO_189 (O_189,N_22340,N_23296);
xor UO_190 (O_190,N_22348,N_23601);
xor UO_191 (O_191,N_23117,N_24348);
xor UO_192 (O_192,N_22697,N_23003);
xnor UO_193 (O_193,N_22834,N_22751);
nor UO_194 (O_194,N_22376,N_22450);
nand UO_195 (O_195,N_23587,N_24809);
nor UO_196 (O_196,N_23241,N_23892);
and UO_197 (O_197,N_23573,N_23702);
nor UO_198 (O_198,N_24292,N_24931);
and UO_199 (O_199,N_21949,N_23931);
or UO_200 (O_200,N_23815,N_24821);
and UO_201 (O_201,N_22743,N_21893);
and UO_202 (O_202,N_23009,N_24765);
nor UO_203 (O_203,N_23256,N_23800);
xor UO_204 (O_204,N_24470,N_21946);
or UO_205 (O_205,N_22636,N_22594);
nor UO_206 (O_206,N_23234,N_24852);
xnor UO_207 (O_207,N_22579,N_23738);
xor UO_208 (O_208,N_22088,N_24763);
nand UO_209 (O_209,N_22963,N_24671);
xor UO_210 (O_210,N_22713,N_22404);
and UO_211 (O_211,N_23344,N_22117);
xor UO_212 (O_212,N_24297,N_23461);
xnor UO_213 (O_213,N_23205,N_23092);
or UO_214 (O_214,N_24233,N_24351);
or UO_215 (O_215,N_24062,N_24921);
or UO_216 (O_216,N_23246,N_22680);
or UO_217 (O_217,N_22809,N_23018);
or UO_218 (O_218,N_24587,N_22406);
and UO_219 (O_219,N_23646,N_23935);
nand UO_220 (O_220,N_24830,N_24368);
and UO_221 (O_221,N_24425,N_22849);
xnor UO_222 (O_222,N_22377,N_24761);
nand UO_223 (O_223,N_24142,N_23993);
or UO_224 (O_224,N_24898,N_22712);
and UO_225 (O_225,N_24146,N_24452);
nor UO_226 (O_226,N_23100,N_23300);
or UO_227 (O_227,N_24219,N_23840);
and UO_228 (O_228,N_23454,N_24028);
nand UO_229 (O_229,N_22551,N_22903);
and UO_230 (O_230,N_23473,N_22918);
and UO_231 (O_231,N_21891,N_24904);
or UO_232 (O_232,N_22794,N_23111);
or UO_233 (O_233,N_24729,N_22157);
nor UO_234 (O_234,N_22227,N_24341);
or UO_235 (O_235,N_24914,N_22182);
and UO_236 (O_236,N_22018,N_22505);
nor UO_237 (O_237,N_23058,N_22969);
xor UO_238 (O_238,N_23554,N_23705);
nand UO_239 (O_239,N_24865,N_23925);
xnor UO_240 (O_240,N_22156,N_22335);
nor UO_241 (O_241,N_22588,N_24546);
nor UO_242 (O_242,N_24900,N_23472);
nand UO_243 (O_243,N_23224,N_22514);
nand UO_244 (O_244,N_22488,N_23804);
nor UO_245 (O_245,N_22259,N_22563);
or UO_246 (O_246,N_23433,N_22576);
nor UO_247 (O_247,N_24726,N_22803);
xor UO_248 (O_248,N_23411,N_23988);
nand UO_249 (O_249,N_23570,N_24694);
or UO_250 (O_250,N_23668,N_22764);
nand UO_251 (O_251,N_21910,N_24069);
nor UO_252 (O_252,N_23426,N_21883);
or UO_253 (O_253,N_24289,N_23661);
and UO_254 (O_254,N_22105,N_24356);
xnor UO_255 (O_255,N_23311,N_23917);
or UO_256 (O_256,N_22577,N_24944);
nor UO_257 (O_257,N_22317,N_23002);
nor UO_258 (O_258,N_23483,N_21929);
nand UO_259 (O_259,N_21906,N_23033);
and UO_260 (O_260,N_24327,N_22027);
nand UO_261 (O_261,N_24928,N_24531);
nor UO_262 (O_262,N_23675,N_22717);
xnor UO_263 (O_263,N_23427,N_22566);
xor UO_264 (O_264,N_21976,N_23810);
nor UO_265 (O_265,N_22532,N_23423);
xnor UO_266 (O_266,N_24479,N_23885);
and UO_267 (O_267,N_24232,N_23137);
xor UO_268 (O_268,N_22961,N_24766);
nand UO_269 (O_269,N_24971,N_23096);
nand UO_270 (O_270,N_24227,N_23284);
or UO_271 (O_271,N_24192,N_24645);
nand UO_272 (O_272,N_24990,N_22388);
xor UO_273 (O_273,N_24771,N_24929);
nand UO_274 (O_274,N_23546,N_24487);
nand UO_275 (O_275,N_23364,N_24579);
nor UO_276 (O_276,N_22536,N_23293);
nand UO_277 (O_277,N_23776,N_22967);
and UO_278 (O_278,N_22454,N_24110);
nand UO_279 (O_279,N_22792,N_22476);
nand UO_280 (O_280,N_24240,N_22997);
xnor UO_281 (O_281,N_22729,N_24693);
nand UO_282 (O_282,N_22483,N_22097);
nor UO_283 (O_283,N_23042,N_23470);
or UO_284 (O_284,N_24455,N_23778);
and UO_285 (O_285,N_23950,N_23091);
nor UO_286 (O_286,N_22080,N_23263);
xor UO_287 (O_287,N_22651,N_22785);
xor UO_288 (O_288,N_24956,N_22336);
and UO_289 (O_289,N_23989,N_23698);
and UO_290 (O_290,N_22653,N_22273);
xor UO_291 (O_291,N_24024,N_22263);
and UO_292 (O_292,N_23360,N_22325);
nand UO_293 (O_293,N_22643,N_23118);
or UO_294 (O_294,N_23779,N_22521);
nand UO_295 (O_295,N_22245,N_24442);
or UO_296 (O_296,N_23053,N_23323);
or UO_297 (O_297,N_24359,N_23307);
or UO_298 (O_298,N_23534,N_22617);
or UO_299 (O_299,N_24635,N_22826);
nor UO_300 (O_300,N_24925,N_24270);
and UO_301 (O_301,N_23847,N_21954);
and UO_302 (O_302,N_24325,N_22831);
nand UO_303 (O_303,N_23106,N_23171);
nor UO_304 (O_304,N_24491,N_22718);
nand UO_305 (O_305,N_23369,N_23697);
nor UO_306 (O_306,N_22323,N_23424);
xnor UO_307 (O_307,N_22224,N_22920);
or UO_308 (O_308,N_24993,N_23188);
nand UO_309 (O_309,N_22300,N_23006);
nor UO_310 (O_310,N_24471,N_24603);
and UO_311 (O_311,N_23134,N_22229);
nor UO_312 (O_312,N_23492,N_24550);
or UO_313 (O_313,N_24433,N_22996);
and UO_314 (O_314,N_23659,N_22719);
or UO_315 (O_315,N_23039,N_24617);
and UO_316 (O_316,N_23863,N_22895);
and UO_317 (O_317,N_23875,N_22832);
or UO_318 (O_318,N_24795,N_23932);
xor UO_319 (O_319,N_24572,N_22331);
xor UO_320 (O_320,N_22285,N_24996);
nor UO_321 (O_321,N_23295,N_22808);
or UO_322 (O_322,N_22069,N_23679);
nor UO_323 (O_323,N_24885,N_24209);
xnor UO_324 (O_324,N_23801,N_21996);
and UO_325 (O_325,N_21916,N_22813);
nand UO_326 (O_326,N_22599,N_22398);
or UO_327 (O_327,N_23605,N_22128);
xnor UO_328 (O_328,N_24476,N_22138);
xor UO_329 (O_329,N_24537,N_24393);
nand UO_330 (O_330,N_23786,N_23947);
xor UO_331 (O_331,N_24543,N_21904);
nand UO_332 (O_332,N_23980,N_22955);
and UO_333 (O_333,N_23743,N_24023);
nand UO_334 (O_334,N_24651,N_24627);
nand UO_335 (O_335,N_24245,N_22004);
xor UO_336 (O_336,N_24385,N_24595);
and UO_337 (O_337,N_24330,N_23494);
xnor UO_338 (O_338,N_23399,N_24244);
nand UO_339 (O_339,N_24656,N_24338);
or UO_340 (O_340,N_22137,N_23191);
or UO_341 (O_341,N_22796,N_22647);
or UO_342 (O_342,N_23381,N_24105);
nor UO_343 (O_343,N_24854,N_22399);
xnor UO_344 (O_344,N_23378,N_23966);
xor UO_345 (O_345,N_22750,N_24926);
nand UO_346 (O_346,N_22822,N_24084);
and UO_347 (O_347,N_23238,N_22385);
nor UO_348 (O_348,N_22142,N_23062);
xnor UO_349 (O_349,N_22434,N_22624);
xnor UO_350 (O_350,N_23325,N_23609);
and UO_351 (O_351,N_22040,N_24932);
nand UO_352 (O_352,N_22574,N_23233);
nand UO_353 (O_353,N_24118,N_22530);
nor UO_354 (O_354,N_23321,N_23539);
and UO_355 (O_355,N_22274,N_23913);
or UO_356 (O_356,N_24556,N_23229);
or UO_357 (O_357,N_21924,N_22247);
xnor UO_358 (O_358,N_22929,N_23069);
xnor UO_359 (O_359,N_23011,N_23357);
or UO_360 (O_360,N_24623,N_24165);
and UO_361 (O_361,N_24189,N_24879);
or UO_362 (O_362,N_22676,N_23481);
and UO_363 (O_363,N_24483,N_22631);
nor UO_364 (O_364,N_23218,N_22922);
nand UO_365 (O_365,N_22108,N_24836);
xor UO_366 (O_366,N_22294,N_24561);
nor UO_367 (O_367,N_22508,N_22421);
or UO_368 (O_368,N_24644,N_22527);
and UO_369 (O_369,N_23363,N_24745);
or UO_370 (O_370,N_23694,N_24802);
nor UO_371 (O_371,N_22757,N_23563);
nand UO_372 (O_372,N_23507,N_22159);
and UO_373 (O_373,N_22744,N_21926);
xor UO_374 (O_374,N_24498,N_24965);
xnor UO_375 (O_375,N_24747,N_22650);
nor UO_376 (O_376,N_24026,N_23036);
nand UO_377 (O_377,N_22806,N_23395);
xor UO_378 (O_378,N_24367,N_23045);
or UO_379 (O_379,N_22035,N_21966);
and UO_380 (O_380,N_24977,N_24302);
xnor UO_381 (O_381,N_21944,N_21969);
and UO_382 (O_382,N_24811,N_24615);
or UO_383 (O_383,N_23741,N_24248);
xor UO_384 (O_384,N_23065,N_22797);
xor UO_385 (O_385,N_24349,N_22082);
nor UO_386 (O_386,N_22824,N_22584);
nor UO_387 (O_387,N_21933,N_22913);
nand UO_388 (O_388,N_22547,N_22120);
or UO_389 (O_389,N_23645,N_21898);
and UO_390 (O_390,N_24353,N_24285);
or UO_391 (O_391,N_23789,N_22706);
or UO_392 (O_392,N_24225,N_23998);
or UO_393 (O_393,N_24991,N_24224);
nand UO_394 (O_394,N_23145,N_22908);
and UO_395 (O_395,N_24369,N_22269);
or UO_396 (O_396,N_24169,N_22258);
nor UO_397 (O_397,N_21942,N_23456);
or UO_398 (O_398,N_23316,N_23287);
or UO_399 (O_399,N_21920,N_23639);
and UO_400 (O_400,N_22887,N_22569);
or UO_401 (O_401,N_22572,N_23594);
or UO_402 (O_402,N_23872,N_22012);
and UO_403 (O_403,N_22498,N_24360);
or UO_404 (O_404,N_22802,N_24841);
nor UO_405 (O_405,N_22418,N_23105);
and UO_406 (O_406,N_24636,N_24862);
or UO_407 (O_407,N_22909,N_24642);
or UO_408 (O_408,N_24672,N_24049);
xnor UO_409 (O_409,N_24737,N_24613);
nand UO_410 (O_410,N_23542,N_23963);
nand UO_411 (O_411,N_22185,N_24299);
xnor UO_412 (O_412,N_23496,N_23374);
and UO_413 (O_413,N_22260,N_22184);
xnor UO_414 (O_414,N_22827,N_24464);
or UO_415 (O_415,N_24933,N_22066);
xnor UO_416 (O_416,N_22308,N_24583);
xor UO_417 (O_417,N_23612,N_22395);
and UO_418 (O_418,N_21999,N_22380);
and UO_419 (O_419,N_23150,N_23959);
nand UO_420 (O_420,N_24610,N_24220);
or UO_421 (O_421,N_22627,N_23141);
or UO_422 (O_422,N_22519,N_23527);
and UO_423 (O_423,N_22902,N_22290);
and UO_424 (O_424,N_23831,N_24275);
nand UO_425 (O_425,N_24007,N_24317);
nor UO_426 (O_426,N_22169,N_24295);
nor UO_427 (O_427,N_22973,N_21963);
nand UO_428 (O_428,N_22622,N_22293);
or UO_429 (O_429,N_23401,N_22402);
nor UO_430 (O_430,N_22853,N_24228);
nand UO_431 (O_431,N_24378,N_23928);
nand UO_432 (O_432,N_23028,N_23102);
or UO_433 (O_433,N_22019,N_24401);
and UO_434 (O_434,N_24387,N_23482);
nor UO_435 (O_435,N_22816,N_24725);
xor UO_436 (O_436,N_22358,N_24590);
and UO_437 (O_437,N_23257,N_23070);
or UO_438 (O_438,N_21964,N_22060);
xnor UO_439 (O_439,N_24685,N_23469);
xnor UO_440 (O_440,N_22366,N_24828);
or UO_441 (O_441,N_22964,N_22937);
nand UO_442 (O_442,N_22878,N_22884);
xnor UO_443 (O_443,N_23538,N_21998);
or UO_444 (O_444,N_22787,N_22585);
xnor UO_445 (O_445,N_23121,N_23918);
and UO_446 (O_446,N_24731,N_24127);
nor UO_447 (O_447,N_23116,N_24058);
nor UO_448 (O_448,N_22447,N_22333);
xnor UO_449 (O_449,N_22026,N_23502);
nand UO_450 (O_450,N_22052,N_22784);
nor UO_451 (O_451,N_23739,N_24048);
or UO_452 (O_452,N_22277,N_22736);
or UO_453 (O_453,N_22249,N_22912);
xor UO_454 (O_454,N_23559,N_24789);
xor UO_455 (O_455,N_23212,N_24536);
xnor UO_456 (O_456,N_22513,N_24089);
or UO_457 (O_457,N_24373,N_24746);
and UO_458 (O_458,N_24328,N_22172);
nand UO_459 (O_459,N_22021,N_24655);
and UO_460 (O_460,N_24708,N_24437);
nor UO_461 (O_461,N_22092,N_23960);
nand UO_462 (O_462,N_23435,N_23579);
xnor UO_463 (O_463,N_23419,N_24174);
nand UO_464 (O_464,N_22425,N_22892);
xnor UO_465 (O_465,N_24008,N_24560);
and UO_466 (O_466,N_22024,N_22817);
or UO_467 (O_467,N_24357,N_23735);
or UO_468 (O_468,N_22819,N_23291);
nor UO_469 (O_469,N_23462,N_24750);
and UO_470 (O_470,N_24139,N_23726);
and UO_471 (O_471,N_22711,N_22379);
and UO_472 (O_472,N_24886,N_23881);
nand UO_473 (O_473,N_22982,N_24625);
nand UO_474 (O_474,N_24384,N_23415);
xor UO_475 (O_475,N_22089,N_23487);
nor UO_476 (O_476,N_23864,N_23761);
or UO_477 (O_477,N_22747,N_23509);
and UO_478 (O_478,N_23590,N_23288);
nor UO_479 (O_479,N_24421,N_22941);
and UO_480 (O_480,N_22393,N_24947);
or UO_481 (O_481,N_24010,N_24919);
nor UO_482 (O_482,N_22804,N_23510);
nor UO_483 (O_483,N_22067,N_23744);
or UO_484 (O_484,N_24051,N_21882);
and UO_485 (O_485,N_24950,N_21981);
nand UO_486 (O_486,N_24850,N_22359);
nand UO_487 (O_487,N_23076,N_23901);
xnor UO_488 (O_488,N_23562,N_22381);
and UO_489 (O_489,N_22791,N_24332);
nor UO_490 (O_490,N_22419,N_23136);
nand UO_491 (O_491,N_24278,N_24974);
xnor UO_492 (O_492,N_22368,N_24216);
or UO_493 (O_493,N_22321,N_23727);
xor UO_494 (O_494,N_24870,N_22554);
or UO_495 (O_495,N_24692,N_24596);
and UO_496 (O_496,N_23666,N_24864);
or UO_497 (O_497,N_22484,N_22432);
nand UO_498 (O_498,N_23418,N_22332);
nor UO_499 (O_499,N_21911,N_23687);
nand UO_500 (O_500,N_24888,N_23690);
and UO_501 (O_501,N_22921,N_24790);
xor UO_502 (O_502,N_23567,N_22989);
xnor UO_503 (O_503,N_22879,N_22270);
xor UO_504 (O_504,N_22439,N_23376);
or UO_505 (O_505,N_24303,N_23508);
and UO_506 (O_506,N_24440,N_24029);
or UO_507 (O_507,N_24591,N_22251);
and UO_508 (O_508,N_23214,N_23762);
xnor UO_509 (O_509,N_24884,N_24516);
nor UO_510 (O_510,N_22106,N_24057);
and UO_511 (O_511,N_22687,N_23782);
or UO_512 (O_512,N_22175,N_23268);
or UO_513 (O_513,N_23654,N_24812);
xnor UO_514 (O_514,N_23783,N_23370);
or UO_515 (O_515,N_23093,N_24858);
nor UO_516 (O_516,N_22934,N_22936);
or UO_517 (O_517,N_23000,N_24099);
and UO_518 (O_518,N_24078,N_23696);
and UO_519 (O_519,N_22218,N_22861);
xnor UO_520 (O_520,N_24276,N_23647);
or UO_521 (O_521,N_23549,N_23271);
xnor UO_522 (O_522,N_22383,N_22568);
and UO_523 (O_523,N_23561,N_23334);
nand UO_524 (O_524,N_24231,N_22254);
or UO_525 (O_525,N_23175,N_22134);
nor UO_526 (O_526,N_22047,N_21971);
and UO_527 (O_527,N_24214,N_22777);
nand UO_528 (O_528,N_24876,N_22553);
nand UO_529 (O_529,N_23195,N_24005);
nand UO_530 (O_530,N_22862,N_24714);
xor UO_531 (O_531,N_24151,N_23650);
nand UO_532 (O_532,N_22465,N_22346);
or UO_533 (O_533,N_24846,N_23375);
or UO_534 (O_534,N_22748,N_24386);
nor UO_535 (O_535,N_23392,N_22314);
nand UO_536 (O_536,N_24999,N_23489);
xor UO_537 (O_537,N_23900,N_22070);
nor UO_538 (O_538,N_22292,N_24458);
nor UO_539 (O_539,N_23692,N_22979);
and UO_540 (O_540,N_22557,N_22761);
or UO_541 (O_541,N_24940,N_23701);
and UO_542 (O_542,N_22707,N_22852);
or UO_543 (O_543,N_23429,N_23757);
nor UO_544 (O_544,N_23580,N_24459);
nor UO_545 (O_545,N_23671,N_24108);
nor UO_546 (O_546,N_23883,N_22931);
nor UO_547 (O_547,N_23685,N_22312);
nor UO_548 (O_548,N_24004,N_22153);
nor UO_549 (O_549,N_23975,N_23148);
or UO_550 (O_550,N_24706,N_22371);
nand UO_551 (O_551,N_24513,N_22363);
or UO_552 (O_552,N_22440,N_24404);
nor UO_553 (O_553,N_22926,N_23910);
and UO_554 (O_554,N_23021,N_23750);
xor UO_555 (O_555,N_22850,N_24682);
and UO_556 (O_556,N_23260,N_24336);
nor UO_557 (O_557,N_24447,N_24252);
xor UO_558 (O_558,N_23084,N_23751);
xnor UO_559 (O_559,N_22025,N_22949);
xor UO_560 (O_560,N_23715,N_24723);
nor UO_561 (O_561,N_23999,N_23660);
xor UO_562 (O_562,N_24265,N_24565);
or UO_563 (O_563,N_21945,N_24564);
and UO_564 (O_564,N_23674,N_24626);
and UO_565 (O_565,N_24037,N_22863);
or UO_566 (O_566,N_22665,N_24905);
and UO_567 (O_567,N_24605,N_23047);
or UO_568 (O_568,N_22467,N_24825);
xor UO_569 (O_569,N_22675,N_23575);
nand UO_570 (O_570,N_24294,N_24422);
and UO_571 (O_571,N_24223,N_24012);
nor UO_572 (O_572,N_22662,N_23090);
nor UO_573 (O_573,N_23830,N_24329);
and UO_574 (O_574,N_22613,N_24849);
or UO_575 (O_575,N_24178,N_23712);
or UO_576 (O_576,N_23547,N_24283);
xor UO_577 (O_577,N_22123,N_23078);
nor UO_578 (O_578,N_23143,N_22565);
xnor UO_579 (O_579,N_24482,N_23416);
xnor UO_580 (O_580,N_23941,N_23657);
xor UO_581 (O_581,N_24874,N_22561);
and UO_582 (O_582,N_23643,N_24117);
nand UO_583 (O_583,N_22013,N_22630);
or UO_584 (O_584,N_22552,N_23040);
and UO_585 (O_585,N_24017,N_23682);
or UO_586 (O_586,N_24512,N_23610);
or UO_587 (O_587,N_23520,N_22322);
or UO_588 (O_588,N_24473,N_24908);
nand UO_589 (O_589,N_22877,N_23389);
nand UO_590 (O_590,N_22571,N_24727);
nand UO_591 (O_591,N_23094,N_23604);
nand UO_592 (O_592,N_22102,N_24164);
and UO_593 (O_593,N_22226,N_22502);
nand UO_594 (O_594,N_24015,N_21947);
nor UO_595 (O_595,N_24686,N_24116);
nor UO_596 (O_596,N_22407,N_23368);
nand UO_597 (O_597,N_23072,N_23314);
or UO_598 (O_598,N_22267,N_22206);
or UO_599 (O_599,N_24150,N_23126);
xor UO_600 (O_600,N_23050,N_23120);
and UO_601 (O_601,N_23156,N_23994);
and UO_602 (O_602,N_23791,N_23479);
and UO_603 (O_603,N_24315,N_24391);
nor UO_604 (O_604,N_22345,N_24354);
and UO_605 (O_605,N_22140,N_23536);
nand UO_606 (O_606,N_23159,N_24515);
or UO_607 (O_607,N_22914,N_23219);
xnor UO_608 (O_608,N_22378,N_22131);
nor UO_609 (O_609,N_22104,N_22164);
xor UO_610 (O_610,N_24207,N_22705);
or UO_611 (O_611,N_24969,N_24705);
nand UO_612 (O_612,N_24868,N_22473);
or UO_613 (O_613,N_23336,N_23759);
nor UO_614 (O_614,N_24320,N_23755);
and UO_615 (O_615,N_22384,N_23642);
and UO_616 (O_616,N_22474,N_24792);
nor UO_617 (O_617,N_22664,N_23231);
xor UO_618 (O_618,N_23742,N_21958);
nor UO_619 (O_619,N_23909,N_22919);
xnor UO_620 (O_620,N_24241,N_24379);
nand UO_621 (O_621,N_24517,N_22305);
or UO_622 (O_622,N_22686,N_22628);
xor UO_623 (O_623,N_23203,N_22875);
and UO_624 (O_624,N_22355,N_24415);
and UO_625 (O_625,N_24432,N_24673);
xor UO_626 (O_626,N_22058,N_21940);
and UO_627 (O_627,N_22735,N_23278);
or UO_628 (O_628,N_24837,N_23254);
nand UO_629 (O_629,N_23101,N_23308);
or UO_630 (O_630,N_24436,N_23167);
nor UO_631 (O_631,N_24638,N_23097);
or UO_632 (O_632,N_22222,N_23807);
nor UO_633 (O_633,N_21955,N_22132);
nor UO_634 (O_634,N_23979,N_23443);
nor UO_635 (O_635,N_23286,N_23393);
nor UO_636 (O_636,N_24680,N_24794);
nor UO_637 (O_637,N_24713,N_22281);
and UO_638 (O_638,N_24260,N_23591);
nor UO_639 (O_639,N_21912,N_24243);
or UO_640 (O_640,N_23920,N_24259);
xor UO_641 (O_641,N_22546,N_22985);
nand UO_642 (O_642,N_23340,N_23382);
or UO_643 (O_643,N_24804,N_24370);
nor UO_644 (O_644,N_24405,N_24322);
nand UO_645 (O_645,N_24469,N_24472);
and UO_646 (O_646,N_24068,N_24532);
and UO_647 (O_647,N_23259,N_22243);
nand UO_648 (O_648,N_24637,N_23708);
xnor UO_649 (O_649,N_22529,N_23819);
nand UO_650 (O_650,N_22500,N_22490);
and UO_651 (O_651,N_24409,N_23850);
and UO_652 (O_652,N_24382,N_23839);
nor UO_653 (O_653,N_22633,N_24691);
nand UO_654 (O_654,N_23080,N_24606);
nand UO_655 (O_655,N_23627,N_22370);
nor UO_656 (O_656,N_23194,N_24462);
xnor UO_657 (O_657,N_23827,N_24783);
xor UO_658 (O_658,N_22022,N_23717);
or UO_659 (O_659,N_21943,N_22077);
nand UO_660 (O_660,N_22210,N_23390);
or UO_661 (O_661,N_22238,N_22600);
nand UO_662 (O_662,N_24978,N_23207);
or UO_663 (O_663,N_22968,N_22452);
nor UO_664 (O_664,N_24751,N_23204);
and UO_665 (O_665,N_24333,N_23616);
nor UO_666 (O_666,N_24123,N_24272);
and UO_667 (O_667,N_24288,N_24833);
nand UO_668 (O_668,N_23406,N_23162);
xor UO_669 (O_669,N_22315,N_22187);
xnor UO_670 (O_670,N_23946,N_22494);
xor UO_671 (O_671,N_22655,N_24624);
xor UO_672 (O_672,N_23361,N_24399);
nor UO_673 (O_673,N_22738,N_24033);
or UO_674 (O_674,N_23157,N_22728);
nor UO_675 (O_675,N_22620,N_23455);
or UO_676 (O_676,N_24593,N_22181);
xor UO_677 (O_677,N_22441,N_24427);
xor UO_678 (O_678,N_24235,N_24738);
or UO_679 (O_679,N_22436,N_24716);
xor UO_680 (O_680,N_22965,N_22595);
nand UO_681 (O_681,N_23377,N_22279);
xor UO_682 (O_682,N_22422,N_24641);
and UO_683 (O_683,N_22559,N_22625);
nor UO_684 (O_684,N_23964,N_23555);
xor UO_685 (O_685,N_24488,N_23967);
or UO_686 (O_686,N_23995,N_24114);
nor UO_687 (O_687,N_24363,N_22846);
xor UO_688 (O_688,N_23858,N_23027);
and UO_689 (O_689,N_23306,N_23498);
and UO_690 (O_690,N_23422,N_24249);
nand UO_691 (O_691,N_23480,N_24082);
and UO_692 (O_692,N_24683,N_22413);
nand UO_693 (O_693,N_22350,N_24824);
and UO_694 (O_694,N_23051,N_23641);
nand UO_695 (O_695,N_22756,N_22209);
nand UO_696 (O_696,N_22788,N_23026);
nand UO_697 (O_697,N_24045,N_24444);
nand UO_698 (O_698,N_24364,N_24001);
nor UO_699 (O_699,N_22076,N_24211);
and UO_700 (O_700,N_24183,N_23228);
or UO_701 (O_701,N_22428,N_23851);
nand UO_702 (O_702,N_23387,N_24549);
nand UO_703 (O_703,N_22606,N_24087);
nand UO_704 (O_704,N_22354,N_24261);
and UO_705 (O_705,N_23607,N_23372);
and UO_706 (O_706,N_23348,N_22255);
and UO_707 (O_707,N_23669,N_22589);
xnor UO_708 (O_708,N_23172,N_23471);
nand UO_709 (O_709,N_22329,N_23957);
xor UO_710 (O_710,N_22948,N_24269);
or UO_711 (O_711,N_23718,N_24927);
nand UO_712 (O_712,N_24514,N_23347);
nor UO_713 (O_713,N_23582,N_23916);
nor UO_714 (O_714,N_23373,N_22512);
nor UO_715 (O_715,N_22762,N_22090);
or UO_716 (O_716,N_24563,N_24149);
nand UO_717 (O_717,N_24733,N_23283);
or UO_718 (O_718,N_24016,N_22692);
and UO_719 (O_719,N_24077,N_22882);
nor UO_720 (O_720,N_24305,N_23301);
nand UO_721 (O_721,N_23730,N_22287);
or UO_722 (O_722,N_22171,N_24428);
xnor UO_723 (O_723,N_22865,N_22416);
xor UO_724 (O_724,N_24412,N_22324);
nor UO_725 (O_725,N_23859,N_22582);
xor UO_726 (O_726,N_24203,N_22382);
nand UO_727 (O_727,N_23584,N_23170);
and UO_728 (O_728,N_24780,N_22740);
and UO_729 (O_729,N_23891,N_24756);
xnor UO_730 (O_730,N_23922,N_21959);
nor UO_731 (O_731,N_22083,N_21968);
nand UO_732 (O_732,N_24659,N_23064);
and UO_733 (O_733,N_22999,N_22001);
xnor UO_734 (O_734,N_23927,N_24902);
nand UO_735 (O_735,N_22029,N_22661);
and UO_736 (O_736,N_23780,N_22959);
nor UO_737 (O_737,N_23201,N_24773);
xnor UO_738 (O_738,N_23569,N_23168);
and UO_739 (O_739,N_24757,N_24262);
xor UO_740 (O_740,N_23689,N_24167);
nor UO_741 (O_741,N_24206,N_23981);
or UO_742 (O_742,N_22390,N_23449);
nand UO_743 (O_743,N_23644,N_24665);
nor UO_744 (O_744,N_22213,N_22220);
xor UO_745 (O_745,N_22148,N_23114);
nor UO_746 (O_746,N_23518,N_22357);
nor UO_747 (O_747,N_24055,N_24907);
nor UO_748 (O_748,N_23294,N_23651);
nand UO_749 (O_749,N_22889,N_23285);
nor UO_750 (O_750,N_23318,N_24237);
and UO_751 (O_751,N_22858,N_23242);
or UO_752 (O_752,N_23317,N_23264);
nor UO_753 (O_753,N_22225,N_24222);
nand UO_754 (O_754,N_22201,N_24578);
nor UO_755 (O_755,N_24815,N_23319);
nor UO_756 (O_756,N_22596,N_22933);
nor UO_757 (O_757,N_22442,N_24621);
nor UO_758 (O_758,N_22896,N_24882);
nor UO_759 (O_759,N_24980,N_24842);
xor UO_760 (O_760,N_23574,N_24496);
or UO_761 (O_761,N_23703,N_22935);
xor UO_762 (O_762,N_22897,N_22240);
or UO_763 (O_763,N_24102,N_23197);
and UO_764 (O_764,N_23919,N_24461);
and UO_765 (O_765,N_24255,N_22907);
xnor UO_766 (O_766,N_22462,N_23414);
xor UO_767 (O_767,N_24758,N_23996);
or UO_768 (O_768,N_23088,N_23798);
and UO_769 (O_769,N_21889,N_22708);
nor UO_770 (O_770,N_23820,N_23765);
nand UO_771 (O_771,N_22970,N_23085);
xnor UO_772 (O_772,N_24869,N_24366);
xnor UO_773 (O_773,N_24197,N_23108);
xor UO_774 (O_774,N_24362,N_24381);
xor UO_775 (O_775,N_22978,N_22339);
and UO_776 (O_776,N_22981,N_23107);
nor UO_777 (O_777,N_24495,N_22790);
nor UO_778 (O_778,N_24614,N_23081);
and UO_779 (O_779,N_24711,N_24153);
and UO_780 (O_780,N_24735,N_23983);
or UO_781 (O_781,N_22174,N_23338);
and UO_782 (O_782,N_23086,N_22009);
nand UO_783 (O_783,N_24523,N_22041);
nor UO_784 (O_784,N_24318,N_24040);
nor UO_785 (O_785,N_24785,N_21941);
and UO_786 (O_786,N_21909,N_22755);
xnor UO_787 (O_787,N_23184,N_23544);
or UO_788 (O_788,N_22365,N_24414);
nand UO_789 (O_789,N_22330,N_22539);
or UO_790 (O_790,N_24200,N_22133);
nor UO_791 (O_791,N_24337,N_23971);
xnor UO_792 (O_792,N_23533,N_22189);
nand UO_793 (O_793,N_24855,N_22776);
or UO_794 (O_794,N_22396,N_23383);
xor UO_795 (O_795,N_23044,N_23262);
xnor UO_796 (O_796,N_23956,N_22626);
and UO_797 (O_797,N_22327,N_24340);
and UO_798 (O_798,N_22463,N_23342);
nor UO_799 (O_799,N_23279,N_23655);
xor UO_800 (O_800,N_23403,N_24650);
xor UO_801 (O_801,N_22723,N_22111);
or UO_802 (O_802,N_24557,N_23451);
and UO_803 (O_803,N_24856,N_24396);
and UO_804 (O_804,N_22983,N_24848);
and UO_805 (O_805,N_22198,N_24020);
nor UO_806 (O_806,N_22954,N_22304);
and UO_807 (O_807,N_23794,N_22417);
xor UO_808 (O_808,N_22810,N_24111);
nand UO_809 (O_809,N_23152,N_22990);
xor UO_810 (O_810,N_24562,N_23142);
or UO_811 (O_811,N_22734,N_24324);
or UO_812 (O_812,N_23977,N_23521);
nand UO_813 (O_813,N_24917,N_22200);
nor UO_814 (O_814,N_22352,N_24377);
nand UO_815 (O_815,N_23973,N_23110);
and UO_816 (O_816,N_23844,N_24113);
nor UO_817 (O_817,N_24630,N_23756);
or UO_818 (O_818,N_23766,N_24279);
nor UO_819 (O_819,N_23535,N_24748);
or UO_820 (O_820,N_22590,N_23954);
or UO_821 (O_821,N_23437,N_24520);
xor UO_822 (O_822,N_22550,N_23876);
and UO_823 (O_823,N_22044,N_24877);
and UO_824 (O_824,N_22095,N_23924);
and UO_825 (O_825,N_24826,N_24066);
and UO_826 (O_826,N_22028,N_23709);
nand UO_827 (O_827,N_24688,N_23202);
or UO_828 (O_828,N_24136,N_22497);
xnor UO_829 (O_829,N_23992,N_22489);
xor UO_830 (O_830,N_24027,N_24522);
nor UO_831 (O_831,N_24797,N_23421);
nor UO_832 (O_832,N_24389,N_24205);
nor UO_833 (O_833,N_23843,N_22732);
nand UO_834 (O_834,N_24553,N_24700);
or UO_835 (O_835,N_24267,N_24287);
xor UO_836 (O_836,N_23965,N_22854);
nand UO_837 (O_837,N_22101,N_24143);
nand UO_838 (O_838,N_21879,N_22306);
xnor UO_839 (O_839,N_24934,N_22397);
nand UO_840 (O_840,N_22288,N_23929);
xnor UO_841 (O_841,N_24937,N_22446);
xor UO_842 (O_842,N_22180,N_22107);
xor UO_843 (O_843,N_23272,N_23266);
and UO_844 (O_844,N_23057,N_24774);
or UO_845 (O_845,N_22668,N_22851);
xnor UO_846 (O_846,N_23493,N_22020);
or UO_847 (O_847,N_24274,N_24810);
xor UO_848 (O_848,N_23329,N_22016);
nand UO_849 (O_849,N_24582,N_22917);
xor UO_850 (O_850,N_24709,N_22065);
xor UO_851 (O_851,N_23198,N_23978);
nand UO_852 (O_852,N_24899,N_23888);
or UO_853 (O_853,N_24468,N_23322);
or UO_854 (O_854,N_22010,N_22696);
or UO_855 (O_855,N_24973,N_23104);
or UO_856 (O_856,N_21938,N_23836);
nand UO_857 (O_857,N_21965,N_24122);
xor UO_858 (O_858,N_24609,N_23129);
nor UO_859 (O_859,N_23211,N_23912);
nand UO_860 (O_860,N_23972,N_22160);
nand UO_861 (O_861,N_23320,N_23740);
and UO_862 (O_862,N_22122,N_24669);
nand UO_863 (O_863,N_24577,N_23602);
nand UO_864 (O_864,N_22389,N_24920);
and UO_865 (O_865,N_22055,N_22485);
nor UO_866 (O_866,N_22930,N_24196);
and UO_867 (O_867,N_23796,N_22236);
or UO_868 (O_868,N_22660,N_23135);
nand UO_869 (O_869,N_24176,N_22644);
nand UO_870 (O_870,N_24441,N_23054);
nand UO_871 (O_871,N_23189,N_24246);
xor UO_872 (O_872,N_22886,N_24507);
and UO_873 (O_873,N_22257,N_23861);
xor UO_874 (O_874,N_22972,N_24552);
xnor UO_875 (O_875,N_24843,N_24450);
or UO_876 (O_876,N_22953,N_21876);
xnor UO_877 (O_877,N_24633,N_23354);
or UO_878 (O_878,N_24551,N_24293);
or UO_879 (O_879,N_24352,N_23577);
and UO_880 (O_880,N_23439,N_24518);
or UO_881 (O_881,N_22161,N_22888);
nor UO_882 (O_882,N_24505,N_22562);
nand UO_883 (O_883,N_23404,N_22062);
nand UO_884 (O_884,N_22205,N_22038);
or UO_885 (O_885,N_23109,N_23553);
and UO_886 (O_886,N_24600,N_22242);
nand UO_887 (O_887,N_23173,N_22995);
xor UO_888 (O_888,N_24660,N_23904);
or UO_889 (O_889,N_23468,N_23710);
xor UO_890 (O_890,N_24647,N_22420);
nand UO_891 (O_891,N_22592,N_21903);
and UO_892 (O_892,N_21939,N_23275);
nand UO_893 (O_893,N_24380,N_24073);
nor UO_894 (O_894,N_23984,N_23315);
xnor UO_895 (O_895,N_21900,N_23032);
xnor UO_896 (O_896,N_23227,N_24791);
nor UO_897 (O_897,N_21905,N_23122);
nor UO_898 (O_898,N_23155,N_24649);
xor UO_899 (O_899,N_23049,N_22373);
xnor UO_900 (O_900,N_21894,N_22894);
or UO_901 (O_901,N_23251,N_24280);
or UO_902 (O_902,N_22960,N_23985);
or UO_903 (O_903,N_22152,N_24161);
xor UO_904 (O_904,N_24916,N_22455);
nand UO_905 (O_905,N_24053,N_24086);
nor UO_906 (O_906,N_24715,N_22526);
and UO_907 (O_907,N_23860,N_23592);
or UO_908 (O_908,N_22522,N_22194);
nand UO_909 (O_909,N_22615,N_24760);
nand UO_910 (O_910,N_24984,N_21884);
or UO_911 (O_911,N_22942,N_24273);
nor UO_912 (O_912,N_23622,N_24668);
or UO_913 (O_913,N_22558,N_24254);
nand UO_914 (O_914,N_24435,N_23345);
nor UO_915 (O_915,N_24034,N_24580);
xnor UO_916 (O_916,N_24859,N_22946);
nor UO_917 (O_917,N_22975,N_23297);
xor UO_918 (O_918,N_22482,N_23095);
and UO_919 (O_919,N_24011,N_21914);
and UO_920 (O_920,N_22278,N_23723);
and UO_921 (O_921,N_22211,N_24312);
or UO_922 (O_922,N_23332,N_22042);
and UO_923 (O_923,N_21962,N_24159);
nor UO_924 (O_924,N_24734,N_24924);
nor UO_925 (O_925,N_23177,N_22109);
nor UO_926 (O_926,N_23048,N_22639);
nor UO_927 (O_927,N_24201,N_23871);
and UO_928 (O_928,N_24730,N_23277);
nor UO_929 (O_929,N_23444,N_22690);
and UO_930 (O_930,N_24485,N_23936);
xor UO_931 (O_931,N_24951,N_23823);
nor UO_932 (O_932,N_24039,N_24499);
and UO_933 (O_933,N_24074,N_24448);
or UO_934 (O_934,N_22524,N_23326);
or UO_935 (O_935,N_24867,N_23772);
nand UO_936 (O_936,N_24199,N_22872);
or UO_937 (O_937,N_22444,N_23884);
xor UO_938 (O_938,N_23600,N_23046);
nor UO_939 (O_939,N_23232,N_22864);
nand UO_940 (O_940,N_22015,N_24987);
and UO_941 (O_941,N_24047,N_22737);
and UO_942 (O_942,N_22033,N_23169);
xnor UO_943 (O_943,N_23082,N_23835);
or UO_944 (O_944,N_23144,N_24881);
nand UO_945 (O_945,N_23013,N_24787);
nand UO_946 (O_946,N_22341,N_23852);
nor UO_947 (O_947,N_24170,N_22769);
nand UO_948 (O_948,N_21917,N_22127);
and UO_949 (O_949,N_22261,N_24814);
nor UO_950 (O_950,N_22621,N_22369);
and UO_951 (O_951,N_21897,N_24141);
nand UO_952 (O_952,N_24144,N_24698);
nand UO_953 (O_953,N_23737,N_22219);
and UO_954 (O_954,N_24208,N_24777);
and UO_955 (O_955,N_24752,N_21887);
and UO_956 (O_956,N_23706,N_23495);
xor UO_957 (O_957,N_23313,N_24967);
nand UO_958 (O_958,N_24217,N_23349);
nor UO_959 (O_959,N_24589,N_24851);
or UO_960 (O_960,N_23298,N_23970);
and UO_961 (O_961,N_22471,N_23138);
xnor UO_962 (O_962,N_23637,N_23532);
or UO_963 (O_963,N_21973,N_23769);
xnor UO_964 (O_964,N_24298,N_24508);
nand UO_965 (O_965,N_24104,N_23289);
xnor UO_966 (O_966,N_24853,N_24400);
xor UO_967 (O_967,N_24739,N_22503);
nor UO_968 (O_968,N_24466,N_23551);
or UO_969 (O_969,N_24355,N_22567);
xor UO_970 (O_970,N_24157,N_23514);
and UO_971 (O_971,N_24309,N_22535);
or UO_972 (O_972,N_23413,N_24819);
nand UO_973 (O_973,N_22938,N_23192);
nor UO_974 (O_974,N_22560,N_22130);
nor UO_975 (O_975,N_22114,N_24014);
or UO_976 (O_976,N_23589,N_22415);
nand UO_977 (O_977,N_24554,N_24239);
xor UO_978 (O_978,N_24607,N_23352);
nor UO_979 (O_979,N_23099,N_23991);
nand UO_980 (O_980,N_24038,N_22392);
and UO_981 (O_981,N_22073,N_22017);
xnor UO_982 (O_982,N_24284,N_22555);
xnor UO_983 (O_983,N_24134,N_24845);
nor UO_984 (O_984,N_23140,N_23799);
and UO_985 (O_985,N_24397,N_23405);
xor UO_986 (O_986,N_21878,N_24675);
nand UO_987 (O_987,N_22427,N_24643);
and UO_988 (O_988,N_22318,N_23711);
xor UO_989 (O_989,N_23133,N_23269);
or UO_990 (O_990,N_24190,N_24912);
nand UO_991 (O_991,N_24574,N_24188);
nand UO_992 (O_992,N_24608,N_22163);
nand UO_993 (O_993,N_21928,N_23811);
xnor UO_994 (O_994,N_24681,N_22611);
nand UO_995 (O_995,N_23530,N_24743);
xor UO_996 (O_996,N_24070,N_22272);
nor UO_997 (O_997,N_24187,N_24446);
xnor UO_998 (O_998,N_22932,N_21935);
nand UO_999 (O_999,N_22099,N_22403);
nand UO_1000 (O_1000,N_23621,N_23548);
nand UO_1001 (O_1001,N_22320,N_24569);
nand UO_1002 (O_1002,N_22874,N_24677);
nor UO_1003 (O_1003,N_22950,N_21988);
or UO_1004 (O_1004,N_23619,N_24394);
xor UO_1005 (O_1005,N_21951,N_24477);
nand UO_1006 (O_1006,N_24710,N_24339);
nor UO_1007 (O_1007,N_22602,N_23200);
and UO_1008 (O_1008,N_23990,N_23700);
nor UO_1009 (O_1009,N_22468,N_22230);
nand UO_1010 (O_1010,N_24323,N_23833);
xnor UO_1011 (O_1011,N_24465,N_24604);
or UO_1012 (O_1012,N_23771,N_24524);
or UO_1013 (O_1013,N_24194,N_24521);
nor UO_1014 (O_1014,N_23166,N_22709);
xnor UO_1015 (O_1015,N_23098,N_23653);
or UO_1016 (O_1016,N_22670,N_23625);
and UO_1017 (O_1017,N_22893,N_22694);
nand UO_1018 (O_1018,N_22741,N_24258);
xor UO_1019 (O_1019,N_24277,N_24903);
or UO_1020 (O_1020,N_22716,N_23817);
nand UO_1021 (O_1021,N_23328,N_22842);
or UO_1022 (O_1022,N_24873,N_22433);
xnor UO_1023 (O_1023,N_23131,N_24036);
nor UO_1024 (O_1024,N_22063,N_24403);
or UO_1025 (O_1025,N_22815,N_22299);
and UO_1026 (O_1026,N_22464,N_23879);
nor UO_1027 (O_1027,N_22608,N_23537);
or UO_1028 (O_1028,N_24775,N_22682);
xnor UO_1029 (O_1029,N_23292,N_22733);
nand UO_1030 (O_1030,N_22360,N_23652);
nor UO_1031 (O_1031,N_23124,N_24793);
and UO_1032 (O_1032,N_24096,N_22186);
xnor UO_1033 (O_1033,N_23583,N_24901);
xor UO_1034 (O_1034,N_24115,N_24500);
and UO_1035 (O_1035,N_24226,N_21888);
xor UO_1036 (O_1036,N_22770,N_22492);
nand UO_1037 (O_1037,N_24032,N_24191);
nand UO_1038 (O_1038,N_24083,N_22679);
and UO_1039 (O_1039,N_23878,N_22141);
or UO_1040 (O_1040,N_22195,N_23945);
nor UO_1041 (O_1041,N_22542,N_23430);
nand UO_1042 (O_1042,N_24107,N_22006);
or UO_1043 (O_1043,N_24992,N_24949);
xnor UO_1044 (O_1044,N_22353,N_22531);
xnor UO_1045 (O_1045,N_24475,N_22121);
or UO_1046 (O_1046,N_24542,N_23898);
xnor UO_1047 (O_1047,N_22564,N_23681);
or UO_1048 (O_1048,N_24119,N_23014);
nand UO_1049 (O_1049,N_22900,N_22268);
or UO_1050 (O_1050,N_22619,N_24210);
and UO_1051 (O_1051,N_24679,N_23475);
and UO_1052 (O_1052,N_23193,N_22724);
xor UO_1053 (O_1053,N_24079,N_23512);
xor UO_1054 (O_1054,N_23631,N_24213);
xor UO_1055 (O_1055,N_23103,N_24424);
nor UO_1056 (O_1056,N_24701,N_24781);
xor UO_1057 (O_1057,N_23558,N_23380);
nand UO_1058 (O_1058,N_23987,N_24687);
nor UO_1059 (O_1059,N_23225,N_23620);
xor UO_1060 (O_1060,N_22867,N_22507);
nor UO_1061 (O_1061,N_24997,N_24654);
or UO_1062 (O_1062,N_22944,N_22614);
and UO_1063 (O_1063,N_23236,N_23597);
nand UO_1064 (O_1064,N_23611,N_23431);
or UO_1065 (O_1065,N_21892,N_24081);
and UO_1066 (O_1066,N_23365,N_23691);
and UO_1067 (O_1067,N_23958,N_24678);
nor UO_1068 (O_1068,N_24529,N_22265);
nor UO_1069 (O_1069,N_23854,N_22873);
xnor UO_1070 (O_1070,N_22911,N_24100);
nand UO_1071 (O_1071,N_24718,N_23672);
xnor UO_1072 (O_1072,N_22739,N_22698);
nor UO_1073 (O_1073,N_24588,N_24883);
nor UO_1074 (O_1074,N_24813,N_23465);
xor UO_1075 (O_1075,N_24803,N_23398);
and UO_1076 (O_1076,N_22666,N_22451);
nor UO_1077 (O_1077,N_22688,N_22658);
nand UO_1078 (O_1078,N_24594,N_22673);
nor UO_1079 (O_1079,N_23459,N_21956);
nand UO_1080 (O_1080,N_23953,N_24417);
xnor UO_1081 (O_1081,N_23802,N_23907);
nor UO_1082 (O_1082,N_24160,N_21931);
nand UO_1083 (O_1083,N_24172,N_24639);
nor UO_1084 (O_1084,N_23822,N_23181);
and UO_1085 (O_1085,N_23425,N_22158);
xnor UO_1086 (O_1086,N_24818,N_22486);
xor UO_1087 (O_1087,N_24314,N_24611);
or UO_1088 (O_1088,N_24132,N_24052);
and UO_1089 (O_1089,N_23037,N_22678);
xnor UO_1090 (O_1090,N_23736,N_24983);
and UO_1091 (O_1091,N_24319,N_22943);
xnor UO_1092 (O_1092,N_23440,N_22876);
nor UO_1093 (O_1093,N_22828,N_24042);
xor UO_1094 (O_1094,N_24571,N_22607);
nor UO_1095 (O_1095,N_23358,N_24184);
or UO_1096 (O_1096,N_23729,N_23677);
xor UO_1097 (O_1097,N_24101,N_23240);
nor UO_1098 (O_1098,N_22275,N_22253);
or UO_1099 (O_1099,N_22191,N_23792);
and UO_1100 (O_1100,N_24493,N_23221);
xnor UO_1101 (O_1101,N_23806,N_23506);
and UO_1102 (O_1102,N_24779,N_23845);
or UO_1103 (O_1103,N_22998,N_24445);
or UO_1104 (O_1104,N_23341,N_24130);
nand UO_1105 (O_1105,N_21923,N_21991);
nand UO_1106 (O_1106,N_24152,N_23066);
and UO_1107 (O_1107,N_23676,N_22125);
or UO_1108 (O_1108,N_21979,N_24025);
or UO_1109 (O_1109,N_24930,N_22193);
nor UO_1110 (O_1110,N_24171,N_23442);
xnor UO_1111 (O_1111,N_24006,N_24304);
or UO_1112 (O_1112,N_24942,N_23767);
nand UO_1113 (O_1113,N_23216,N_24618);
xnor UO_1114 (O_1114,N_23030,N_21957);
xnor UO_1115 (O_1115,N_23255,N_23773);
nand UO_1116 (O_1116,N_23728,N_23614);
nand UO_1117 (O_1117,N_22641,N_23745);
and UO_1118 (O_1118,N_24832,N_21983);
and UO_1119 (O_1119,N_23312,N_24648);
and UO_1120 (O_1120,N_23812,N_21932);
xnor UO_1121 (O_1121,N_24619,N_22298);
xor UO_1122 (O_1122,N_22496,N_22927);
nor UO_1123 (O_1123,N_24202,N_24056);
xor UO_1124 (O_1124,N_22414,N_22048);
or UO_1125 (O_1125,N_23083,N_22722);
xnor UO_1126 (O_1126,N_24622,N_23524);
or UO_1127 (O_1127,N_23764,N_24918);
nand UO_1128 (O_1128,N_23089,N_23982);
or UO_1129 (O_1129,N_23217,N_24541);
or UO_1130 (O_1130,N_21952,N_21961);
or UO_1131 (O_1131,N_24696,N_22593);
or UO_1132 (O_1132,N_24281,N_24375);
or UO_1133 (O_1133,N_23366,N_23491);
and UO_1134 (O_1134,N_24875,N_22068);
or UO_1135 (O_1135,N_22623,N_22545);
or UO_1136 (O_1136,N_23797,N_24509);
and UO_1137 (O_1137,N_22905,N_22235);
nand UO_1138 (O_1138,N_23408,N_23213);
xnor UO_1139 (O_1139,N_24129,N_22232);
and UO_1140 (O_1140,N_23350,N_23873);
xnor UO_1141 (O_1141,N_22031,N_22984);
xnor UO_1142 (O_1142,N_24438,N_24568);
nor UO_1143 (O_1143,N_23874,N_23477);
nand UO_1144 (O_1144,N_22343,N_24095);
nand UO_1145 (O_1145,N_24021,N_24776);
nand UO_1146 (O_1146,N_23581,N_23832);
or UO_1147 (O_1147,N_23603,N_23933);
nor UO_1148 (O_1148,N_22303,N_22573);
nor UO_1149 (O_1149,N_22449,N_24019);
xnor UO_1150 (O_1150,N_23938,N_22977);
xnor UO_1151 (O_1151,N_22347,N_24910);
nand UO_1152 (O_1152,N_23304,N_22715);
or UO_1153 (O_1153,N_22291,N_24451);
nand UO_1154 (O_1154,N_24527,N_22190);
xnor UO_1155 (O_1155,N_21907,N_23760);
and UO_1156 (O_1156,N_24195,N_22276);
and UO_1157 (O_1157,N_23453,N_22663);
or UO_1158 (O_1158,N_24492,N_22192);
nand UO_1159 (O_1159,N_23400,N_22674);
xnor UO_1160 (O_1160,N_23346,N_22081);
xnor UO_1161 (O_1161,N_22493,N_22916);
nor UO_1162 (O_1162,N_24878,N_22801);
nand UO_1163 (O_1163,N_24268,N_23123);
and UO_1164 (O_1164,N_22847,N_23825);
nand UO_1165 (O_1165,N_24179,N_24778);
xor UO_1166 (O_1166,N_22049,N_24519);
nor UO_1167 (O_1167,N_24266,N_23566);
nor UO_1168 (O_1168,N_24061,N_22043);
xor UO_1169 (O_1169,N_23889,N_24423);
xnor UO_1170 (O_1170,N_22098,N_22667);
nor UO_1171 (O_1171,N_24022,N_22409);
or UO_1172 (O_1172,N_24955,N_22034);
xnor UO_1173 (O_1173,N_23226,N_24695);
nor UO_1174 (O_1174,N_24767,N_24860);
xor UO_1175 (O_1175,N_23754,N_22212);
or UO_1176 (O_1176,N_22509,N_22993);
or UO_1177 (O_1177,N_24454,N_24257);
nand UO_1178 (O_1178,N_22056,N_23695);
nand UO_1179 (O_1179,N_23258,N_23210);
and UO_1180 (O_1180,N_23640,N_22244);
or UO_1181 (O_1181,N_24484,N_23187);
nor UO_1182 (O_1182,N_24510,N_24177);
xnor UO_1183 (O_1183,N_24308,N_23178);
or UO_1184 (O_1184,N_24181,N_23282);
and UO_1185 (O_1185,N_23273,N_23523);
xor UO_1186 (O_1186,N_22772,N_21995);
xor UO_1187 (O_1187,N_22411,N_22683);
nor UO_1188 (O_1188,N_24467,N_22540);
and UO_1189 (O_1189,N_22992,N_23158);
and UO_1190 (O_1190,N_24212,N_24670);
nand UO_1191 (O_1191,N_22657,N_24663);
or UO_1192 (O_1192,N_22188,N_22150);
and UO_1193 (O_1193,N_23606,N_24525);
and UO_1194 (O_1194,N_24911,N_24372);
nor UO_1195 (O_1195,N_24799,N_24909);
xor UO_1196 (O_1196,N_24000,N_22681);
nand UO_1197 (O_1197,N_24121,N_23163);
and UO_1198 (O_1198,N_21886,N_23450);
nor UO_1199 (O_1199,N_24343,N_24871);
or UO_1200 (O_1200,N_22689,N_22326);
xnor UO_1201 (O_1201,N_22609,N_23848);
nand UO_1202 (O_1202,N_24494,N_22113);
nand UO_1203 (O_1203,N_24555,N_22309);
nor UO_1204 (O_1204,N_24894,N_24041);
xnor UO_1205 (O_1205,N_24759,N_24511);
nor UO_1206 (O_1206,N_23896,N_23526);
and UO_1207 (O_1207,N_23008,N_24247);
xnor UO_1208 (O_1208,N_24970,N_22241);
nor UO_1209 (O_1209,N_24979,N_22742);
nand UO_1210 (O_1210,N_22438,N_23781);
xor UO_1211 (O_1211,N_21994,N_24915);
xor UO_1212 (O_1212,N_23531,N_24722);
nand UO_1213 (O_1213,N_22208,N_24959);
nor UO_1214 (O_1214,N_24145,N_23747);
nor UO_1215 (O_1215,N_22064,N_23010);
nor UO_1216 (O_1216,N_22976,N_24570);
or UO_1217 (O_1217,N_22533,N_23869);
xnor UO_1218 (O_1218,N_23183,N_22374);
or UO_1219 (O_1219,N_22730,N_24982);
nor UO_1220 (O_1220,N_22800,N_24755);
nor UO_1221 (O_1221,N_23497,N_24090);
nor UO_1222 (O_1222,N_24088,N_22430);
nand UO_1223 (O_1223,N_23516,N_22475);
or UO_1224 (O_1224,N_23327,N_22386);
or UO_1225 (O_1225,N_22057,N_23842);
or UO_1226 (O_1226,N_23132,N_23252);
nor UO_1227 (O_1227,N_23125,N_22833);
or UO_1228 (O_1228,N_23305,N_24960);
and UO_1229 (O_1229,N_24584,N_22256);
xnor UO_1230 (O_1230,N_23545,N_21899);
xor UO_1231 (O_1231,N_24838,N_23017);
nand UO_1232 (O_1232,N_24816,N_23593);
xor UO_1233 (O_1233,N_24044,N_22710);
nor UO_1234 (O_1234,N_23467,N_22491);
xor UO_1235 (O_1235,N_22085,N_23940);
nor UO_1236 (O_1236,N_23434,N_22214);
nand UO_1237 (O_1237,N_22731,N_24193);
and UO_1238 (O_1238,N_22094,N_21934);
xnor UO_1239 (O_1239,N_24800,N_23886);
nand UO_1240 (O_1240,N_22974,N_23190);
or UO_1241 (O_1241,N_24406,N_22246);
or UO_1242 (O_1242,N_23019,N_22351);
and UO_1243 (O_1243,N_24296,N_22231);
xnor UO_1244 (O_1244,N_22003,N_24457);
and UO_1245 (O_1245,N_22991,N_24558);
xnor UO_1246 (O_1246,N_24182,N_23598);
and UO_1247 (O_1247,N_24075,N_24943);
xor UO_1248 (O_1248,N_22753,N_23244);
xnor UO_1249 (O_1249,N_24147,N_23572);
nor UO_1250 (O_1250,N_22173,N_23813);
or UO_1251 (O_1251,N_22506,N_23955);
and UO_1252 (O_1252,N_24185,N_24526);
xor UO_1253 (O_1253,N_23031,N_22701);
and UO_1254 (O_1254,N_23809,N_22752);
or UO_1255 (O_1255,N_24952,N_23474);
nand UO_1256 (O_1256,N_22400,N_23894);
xor UO_1257 (O_1257,N_24827,N_22075);
and UO_1258 (O_1258,N_22221,N_23087);
nand UO_1259 (O_1259,N_23680,N_22197);
or UO_1260 (O_1260,N_22841,N_23826);
nor UO_1261 (O_1261,N_23517,N_24697);
or UO_1262 (O_1262,N_23733,N_22605);
or UO_1263 (O_1263,N_23253,N_21985);
or UO_1264 (O_1264,N_23828,N_24576);
and UO_1265 (O_1265,N_23725,N_22051);
xor UO_1266 (O_1266,N_23447,N_24271);
or UO_1267 (O_1267,N_23856,N_23557);
nor UO_1268 (O_1268,N_23463,N_23139);
and UO_1269 (O_1269,N_23915,N_22036);
xor UO_1270 (O_1270,N_22525,N_22939);
nor UO_1271 (O_1271,N_22165,N_23528);
xor UO_1272 (O_1272,N_22435,N_24946);
xnor UO_1273 (O_1273,N_21901,N_24863);
and UO_1274 (O_1274,N_23303,N_24300);
xnor UO_1275 (O_1275,N_23568,N_23937);
xor UO_1276 (O_1276,N_22581,N_24236);
xnor UO_1277 (O_1277,N_24112,N_23113);
xnor UO_1278 (O_1278,N_24402,N_22501);
or UO_1279 (O_1279,N_23942,N_22124);
xor UO_1280 (O_1280,N_22659,N_24741);
and UO_1281 (O_1281,N_24128,N_22387);
xor UO_1282 (O_1282,N_23337,N_24620);
nand UO_1283 (O_1283,N_22426,N_22477);
nor UO_1284 (O_1284,N_22168,N_23351);
xnor UO_1285 (O_1285,N_23897,N_23519);
nor UO_1286 (O_1286,N_24092,N_24085);
xor UO_1287 (O_1287,N_24358,N_22829);
or UO_1288 (O_1288,N_22924,N_23949);
nand UO_1289 (O_1289,N_23038,N_23079);
nand UO_1290 (O_1290,N_24043,N_24418);
and UO_1291 (O_1291,N_24431,N_24953);
nand UO_1292 (O_1292,N_22037,N_24204);
and UO_1293 (O_1293,N_22100,N_22215);
and UO_1294 (O_1294,N_22994,N_24676);
nor UO_1295 (O_1295,N_24426,N_22248);
and UO_1296 (O_1296,N_21937,N_24030);
xnor UO_1297 (O_1297,N_23588,N_22881);
nand UO_1298 (O_1298,N_24958,N_22721);
nor UO_1299 (O_1299,N_23777,N_23029);
and UO_1300 (O_1300,N_24003,N_22838);
xnor UO_1301 (O_1301,N_22289,N_22014);
and UO_1302 (O_1302,N_23890,N_23513);
or UO_1303 (O_1303,N_24801,N_24602);
nor UO_1304 (O_1304,N_22778,N_22499);
nand UO_1305 (O_1305,N_22549,N_24168);
nor UO_1306 (O_1306,N_22118,N_24311);
xnor UO_1307 (O_1307,N_24658,N_22835);
xnor UO_1308 (O_1308,N_24597,N_22091);
nand UO_1309 (O_1309,N_24453,N_22429);
xor UO_1310 (O_1310,N_22799,N_22431);
or UO_1311 (O_1311,N_24664,N_22836);
nand UO_1312 (O_1312,N_24976,N_24481);
nand UO_1313 (O_1313,N_23043,N_21989);
or UO_1314 (O_1314,N_22344,N_23683);
or UO_1315 (O_1315,N_22704,N_24897);
or UO_1316 (O_1316,N_24895,N_22334);
nand UO_1317 (O_1317,N_22899,N_24242);
xor UO_1318 (O_1318,N_24067,N_24290);
or UO_1319 (O_1319,N_22821,N_23220);
or UO_1320 (O_1320,N_24770,N_24721);
and UO_1321 (O_1321,N_22767,N_22774);
and UO_1322 (O_1322,N_23015,N_22986);
and UO_1323 (O_1323,N_23868,N_22126);
or UO_1324 (O_1324,N_22591,N_24601);
xor UO_1325 (O_1325,N_22883,N_24889);
and UO_1326 (O_1326,N_22947,N_22008);
and UO_1327 (O_1327,N_22179,N_22583);
and UO_1328 (O_1328,N_22646,N_23276);
or UO_1329 (O_1329,N_24598,N_22280);
and UO_1330 (O_1330,N_22837,N_24749);
and UO_1331 (O_1331,N_22685,N_23164);
nand UO_1332 (O_1332,N_23309,N_24820);
xnor UO_1333 (O_1333,N_22754,N_22807);
or UO_1334 (O_1334,N_22915,N_22149);
nand UO_1335 (O_1335,N_24125,N_23948);
or UO_1336 (O_1336,N_23837,N_22310);
and UO_1337 (O_1337,N_22356,N_24478);
nor UO_1338 (O_1338,N_23068,N_23270);
or UO_1339 (O_1339,N_23417,N_22957);
nand UO_1340 (O_1340,N_23119,N_23333);
nand UO_1341 (O_1341,N_22597,N_22264);
nor UO_1342 (O_1342,N_24575,N_22610);
nand UO_1343 (O_1343,N_23356,N_23071);
and UO_1344 (O_1344,N_24419,N_22823);
nor UO_1345 (O_1345,N_22510,N_24740);
nand UO_1346 (O_1346,N_21877,N_22518);
or UO_1347 (O_1347,N_21936,N_22702);
or UO_1348 (O_1348,N_23908,N_23608);
and UO_1349 (O_1349,N_24922,N_24547);
nand UO_1350 (O_1350,N_22311,N_22885);
xnor UO_1351 (O_1351,N_22910,N_22781);
xnor UO_1352 (O_1352,N_23673,N_24839);
and UO_1353 (O_1353,N_24840,N_23719);
nor UO_1354 (O_1354,N_24736,N_24186);
nand UO_1355 (O_1355,N_23716,N_22805);
and UO_1356 (O_1356,N_22763,N_23074);
xor UO_1357 (O_1357,N_24861,N_23613);
or UO_1358 (O_1358,N_22511,N_22637);
and UO_1359 (O_1359,N_22857,N_23540);
nand UO_1360 (O_1360,N_24788,N_23857);
xor UO_1361 (O_1361,N_22891,N_23359);
xnor UO_1362 (O_1362,N_23623,N_22548);
and UO_1363 (O_1363,N_23814,N_22634);
xnor UO_1364 (O_1364,N_23490,N_24374);
nor UO_1365 (O_1365,N_24661,N_21895);
nand UO_1366 (O_1366,N_23208,N_23261);
nand UO_1367 (O_1367,N_22830,N_22958);
and UO_1368 (O_1368,N_23335,N_23245);
and UO_1369 (O_1369,N_24823,N_23247);
and UO_1370 (O_1370,N_24175,N_22782);
nor UO_1371 (O_1371,N_24599,N_22632);
xnor UO_1372 (O_1372,N_24138,N_22760);
and UO_1373 (O_1373,N_23522,N_24126);
nor UO_1374 (O_1374,N_22603,N_24198);
xor UO_1375 (O_1375,N_24684,N_23025);
xor UO_1376 (O_1376,N_23249,N_22319);
and UO_1377 (O_1377,N_24891,N_22901);
or UO_1378 (O_1378,N_23128,N_23409);
nor UO_1379 (O_1379,N_23816,N_24251);
or UO_1380 (O_1380,N_23877,N_22453);
nand UO_1381 (O_1381,N_23969,N_23209);
nor UO_1382 (O_1382,N_22825,N_23649);
nor UO_1383 (O_1383,N_22771,N_23146);
and UO_1384 (O_1384,N_24772,N_22677);
nor UO_1385 (O_1385,N_23887,N_24640);
nand UO_1386 (O_1386,N_23391,N_22170);
xor UO_1387 (O_1387,N_23153,N_24559);
and UO_1388 (O_1388,N_22616,N_24013);
xnor UO_1389 (O_1389,N_23618,N_24786);
or UO_1390 (O_1390,N_22671,N_24784);
xor UO_1391 (O_1391,N_23867,N_23824);
nand UO_1392 (O_1392,N_24548,N_22039);
nor UO_1393 (O_1393,N_24972,N_22703);
and UO_1394 (O_1394,N_24653,N_24968);
xor UO_1395 (O_1395,N_22176,N_22798);
and UO_1396 (O_1396,N_22412,N_22177);
xor UO_1397 (O_1397,N_23790,N_22461);
nand UO_1398 (O_1398,N_23505,N_22478);
or UO_1399 (O_1399,N_23115,N_23511);
xor UO_1400 (O_1400,N_24103,N_22437);
and UO_1401 (O_1401,N_23670,N_22459);
nand UO_1402 (O_1402,N_24460,N_24158);
xnor UO_1403 (O_1403,N_22096,N_24383);
and UO_1404 (O_1404,N_23248,N_24890);
or UO_1405 (O_1405,N_23962,N_23921);
nand UO_1406 (O_1406,N_24831,N_24896);
and UO_1407 (O_1407,N_24135,N_23882);
nand UO_1408 (O_1408,N_23684,N_23016);
nor UO_1409 (O_1409,N_22223,N_23624);
xor UO_1410 (O_1410,N_23923,N_23310);
xor UO_1411 (O_1411,N_23302,N_22284);
nor UO_1412 (O_1412,N_23724,N_22147);
nand UO_1413 (O_1413,N_22295,N_23239);
nor UO_1414 (O_1414,N_22443,N_24662);
nor UO_1415 (O_1415,N_24941,N_23484);
or UO_1416 (O_1416,N_21908,N_24834);
or UO_1417 (O_1417,N_22239,N_23596);
or UO_1418 (O_1418,N_24935,N_22987);
and UO_1419 (O_1419,N_23699,N_22151);
and UO_1420 (O_1420,N_23060,N_23073);
nand UO_1421 (O_1421,N_22635,N_24857);
nand UO_1422 (O_1422,N_23130,N_22906);
and UO_1423 (O_1423,N_22116,N_23865);
xnor UO_1424 (O_1424,N_24501,N_22759);
nand UO_1425 (O_1425,N_23866,N_22297);
and UO_1426 (O_1426,N_23746,N_24769);
nand UO_1427 (O_1427,N_24844,N_24413);
nand UO_1428 (O_1428,N_23748,N_24689);
nor UO_1429 (O_1429,N_23274,N_23862);
nand UO_1430 (O_1430,N_23552,N_23880);
and UO_1431 (O_1431,N_23280,N_22237);
nand UO_1432 (O_1432,N_24306,N_22030);
nor UO_1433 (O_1433,N_22971,N_22543);
nor UO_1434 (O_1434,N_23179,N_23460);
or UO_1435 (O_1435,N_22868,N_23331);
and UO_1436 (O_1436,N_22410,N_24994);
nand UO_1437 (O_1437,N_23503,N_24796);
nand UO_1438 (O_1438,N_22479,N_23466);
or UO_1439 (O_1439,N_21919,N_22307);
and UO_1440 (O_1440,N_22135,N_22115);
xor UO_1441 (O_1441,N_22457,N_22537);
or UO_1442 (O_1442,N_22328,N_22375);
nand UO_1443 (O_1443,N_23488,N_24581);
nor UO_1444 (O_1444,N_23855,N_22945);
xor UO_1445 (O_1445,N_22860,N_23004);
and UO_1446 (O_1446,N_24301,N_24966);
nand UO_1447 (O_1447,N_22693,N_22046);
and UO_1448 (O_1448,N_23997,N_22726);
or UO_1449 (O_1449,N_22301,N_23024);
xor UO_1450 (O_1450,N_23720,N_22765);
or UO_1451 (O_1451,N_21918,N_23186);
xor UO_1452 (O_1452,N_23976,N_23795);
and UO_1453 (O_1453,N_22162,N_23556);
or UO_1454 (O_1454,N_22840,N_24091);
or UO_1455 (O_1455,N_24822,N_22775);
xnor UO_1456 (O_1456,N_23713,N_22337);
xnor UO_1457 (O_1457,N_23678,N_22604);
xor UO_1458 (O_1458,N_23525,N_22871);
and UO_1459 (O_1459,N_23630,N_22053);
nand UO_1460 (O_1460,N_21977,N_23752);
xor UO_1461 (O_1461,N_22580,N_22768);
nand UO_1462 (O_1462,N_24371,N_24699);
nor UO_1463 (O_1463,N_23500,N_23770);
nor UO_1464 (O_1464,N_23543,N_24076);
nor UO_1465 (O_1465,N_24936,N_24106);
and UO_1466 (O_1466,N_24456,N_24892);
nand UO_1467 (O_1467,N_22079,N_22342);
xnor UO_1468 (O_1468,N_24807,N_22640);
nand UO_1469 (O_1469,N_24331,N_24923);
or UO_1470 (O_1470,N_22654,N_22316);
xor UO_1471 (O_1471,N_24350,N_23063);
nand UO_1472 (O_1472,N_21922,N_23662);
xor UO_1473 (O_1473,N_22093,N_22783);
or UO_1474 (O_1474,N_23629,N_24986);
or UO_1475 (O_1475,N_22005,N_23663);
xnor UO_1476 (O_1476,N_22988,N_23504);
nor UO_1477 (O_1477,N_22061,N_23803);
nand UO_1478 (O_1478,N_21896,N_24535);
and UO_1479 (O_1479,N_22023,N_24215);
and UO_1480 (O_1480,N_22820,N_22648);
xnor UO_1481 (O_1481,N_24009,N_23565);
nor UO_1482 (O_1482,N_22154,N_22869);
nor UO_1483 (O_1483,N_23222,N_23441);
and UO_1484 (O_1484,N_24939,N_22204);
nor UO_1485 (O_1485,N_22233,N_22669);
xnor UO_1486 (O_1486,N_22283,N_22618);
nor UO_1487 (O_1487,N_24835,N_24629);
or UO_1488 (O_1488,N_22520,N_24732);
and UO_1489 (O_1489,N_23160,N_23362);
nor UO_1490 (O_1490,N_24093,N_22282);
xnor UO_1491 (O_1491,N_21980,N_24346);
and UO_1492 (O_1492,N_23343,N_23951);
or UO_1493 (O_1493,N_23784,N_24995);
or UO_1494 (O_1494,N_23394,N_21993);
nor UO_1495 (O_1495,N_22672,N_24567);
and UO_1496 (O_1496,N_23626,N_22758);
nand UO_1497 (O_1497,N_24963,N_24256);
xnor UO_1498 (O_1498,N_22575,N_22087);
or UO_1499 (O_1499,N_21921,N_24906);
or UO_1500 (O_1500,N_24335,N_22074);
nand UO_1501 (O_1501,N_24502,N_23586);
xnor UO_1502 (O_1502,N_23688,N_22472);
nand UO_1503 (O_1503,N_24728,N_24410);
and UO_1504 (O_1504,N_24486,N_24829);
nor UO_1505 (O_1505,N_23893,N_23154);
nor UO_1506 (O_1506,N_22155,N_23829);
nor UO_1507 (O_1507,N_23615,N_24263);
and UO_1508 (O_1508,N_24938,N_23412);
or UO_1509 (O_1509,N_23199,N_22843);
and UO_1510 (O_1510,N_24392,N_22313);
nor UO_1511 (O_1511,N_22544,N_23180);
nor UO_1512 (O_1512,N_23846,N_24365);
xor UO_1513 (O_1513,N_23151,N_21960);
nand UO_1514 (O_1514,N_23774,N_22714);
nand UO_1515 (O_1515,N_23632,N_24489);
and UO_1516 (O_1516,N_24988,N_23895);
and UO_1517 (O_1517,N_23371,N_22601);
nand UO_1518 (O_1518,N_24443,N_22818);
nand UO_1519 (O_1519,N_24230,N_23464);
xnor UO_1520 (O_1520,N_23428,N_23353);
nor UO_1521 (O_1521,N_24474,N_24155);
xor UO_1522 (O_1522,N_22252,N_21974);
nand UO_1523 (O_1523,N_23939,N_22856);
or UO_1524 (O_1524,N_21997,N_22032);
or UO_1525 (O_1525,N_21902,N_24376);
and UO_1526 (O_1526,N_24342,N_23636);
or UO_1527 (O_1527,N_24768,N_24395);
xnor UO_1528 (O_1528,N_22203,N_23787);
nand UO_1529 (O_1529,N_23899,N_22773);
nand UO_1530 (O_1530,N_23821,N_24657);
nor UO_1531 (O_1531,N_23903,N_22054);
nor UO_1532 (O_1532,N_23665,N_22136);
xor UO_1533 (O_1533,N_23112,N_22271);
nor UO_1534 (O_1534,N_23161,N_24764);
xor UO_1535 (O_1535,N_24666,N_22480);
nand UO_1536 (O_1536,N_24140,N_21925);
or UO_1537 (O_1537,N_23386,N_24872);
nand UO_1538 (O_1538,N_24528,N_23617);
or UO_1539 (O_1539,N_23515,N_21984);
xnor UO_1540 (O_1540,N_23020,N_22811);
and UO_1541 (O_1541,N_22786,N_22262);
nor UO_1542 (O_1542,N_24018,N_24948);
or UO_1543 (O_1543,N_23721,N_21972);
nand UO_1544 (O_1544,N_23968,N_23775);
or UO_1545 (O_1545,N_23943,N_24408);
nor UO_1546 (O_1546,N_24631,N_23634);
or UO_1547 (O_1547,N_24538,N_24434);
and UO_1548 (O_1548,N_23658,N_23599);
or UO_1549 (O_1549,N_22372,N_23267);
and UO_1550 (O_1550,N_24847,N_24463);
and UO_1551 (O_1551,N_23906,N_24712);
nor UO_1552 (O_1552,N_22423,N_24490);
nor UO_1553 (O_1553,N_22928,N_21987);
xor UO_1554 (O_1554,N_24334,N_23339);
nand UO_1555 (O_1555,N_22394,N_23870);
xor UO_1556 (O_1556,N_23022,N_24162);
or UO_1557 (O_1557,N_24503,N_22166);
or UO_1558 (O_1558,N_21948,N_22487);
or UO_1559 (O_1559,N_22302,N_24880);
or UO_1560 (O_1560,N_22570,N_23250);
nor UO_1561 (O_1561,N_22516,N_24234);
nor UO_1562 (O_1562,N_24957,N_24181);
xnor UO_1563 (O_1563,N_24110,N_22178);
xor UO_1564 (O_1564,N_21893,N_23757);
nor UO_1565 (O_1565,N_21897,N_24467);
xnor UO_1566 (O_1566,N_23298,N_23629);
nor UO_1567 (O_1567,N_24108,N_22245);
or UO_1568 (O_1568,N_23751,N_23870);
or UO_1569 (O_1569,N_24714,N_23358);
nand UO_1570 (O_1570,N_24620,N_24534);
nor UO_1571 (O_1571,N_24142,N_22156);
and UO_1572 (O_1572,N_23518,N_24172);
nor UO_1573 (O_1573,N_24432,N_23546);
xnor UO_1574 (O_1574,N_22416,N_23311);
xor UO_1575 (O_1575,N_22819,N_22946);
xor UO_1576 (O_1576,N_22377,N_24600);
nand UO_1577 (O_1577,N_22360,N_23591);
nand UO_1578 (O_1578,N_24174,N_23313);
or UO_1579 (O_1579,N_22434,N_22264);
or UO_1580 (O_1580,N_22303,N_23497);
or UO_1581 (O_1581,N_24394,N_24903);
xor UO_1582 (O_1582,N_23796,N_22002);
nor UO_1583 (O_1583,N_23710,N_23473);
nand UO_1584 (O_1584,N_24084,N_22087);
xnor UO_1585 (O_1585,N_22154,N_24137);
and UO_1586 (O_1586,N_24471,N_24092);
nor UO_1587 (O_1587,N_22784,N_24939);
xor UO_1588 (O_1588,N_23747,N_23610);
or UO_1589 (O_1589,N_24381,N_24999);
nor UO_1590 (O_1590,N_22565,N_22169);
and UO_1591 (O_1591,N_22486,N_24796);
nor UO_1592 (O_1592,N_23214,N_22370);
nor UO_1593 (O_1593,N_22565,N_23818);
nor UO_1594 (O_1594,N_24446,N_23456);
nand UO_1595 (O_1595,N_23809,N_24077);
and UO_1596 (O_1596,N_22421,N_24420);
nor UO_1597 (O_1597,N_21988,N_22419);
nand UO_1598 (O_1598,N_24487,N_23332);
and UO_1599 (O_1599,N_22380,N_24079);
or UO_1600 (O_1600,N_23485,N_23597);
and UO_1601 (O_1601,N_22539,N_23790);
and UO_1602 (O_1602,N_22994,N_22315);
nand UO_1603 (O_1603,N_23757,N_23981);
nor UO_1604 (O_1604,N_24234,N_23632);
nand UO_1605 (O_1605,N_23429,N_22961);
nor UO_1606 (O_1606,N_24837,N_23620);
or UO_1607 (O_1607,N_23645,N_23593);
nor UO_1608 (O_1608,N_22864,N_24795);
xor UO_1609 (O_1609,N_22458,N_22308);
and UO_1610 (O_1610,N_24344,N_24221);
nand UO_1611 (O_1611,N_24860,N_23073);
nand UO_1612 (O_1612,N_24604,N_22117);
nor UO_1613 (O_1613,N_22705,N_22917);
nor UO_1614 (O_1614,N_24416,N_24812);
nor UO_1615 (O_1615,N_24024,N_24035);
nor UO_1616 (O_1616,N_22633,N_24346);
xnor UO_1617 (O_1617,N_22305,N_23234);
xor UO_1618 (O_1618,N_24089,N_23870);
xor UO_1619 (O_1619,N_24830,N_22466);
xnor UO_1620 (O_1620,N_24595,N_23399);
or UO_1621 (O_1621,N_24240,N_24150);
nor UO_1622 (O_1622,N_24704,N_22016);
nor UO_1623 (O_1623,N_21955,N_23898);
and UO_1624 (O_1624,N_22777,N_23792);
nand UO_1625 (O_1625,N_23464,N_22038);
xnor UO_1626 (O_1626,N_24570,N_23029);
nor UO_1627 (O_1627,N_24424,N_22018);
and UO_1628 (O_1628,N_23974,N_22037);
nand UO_1629 (O_1629,N_23662,N_22656);
nor UO_1630 (O_1630,N_23065,N_23759);
and UO_1631 (O_1631,N_23404,N_22106);
and UO_1632 (O_1632,N_23300,N_24530);
or UO_1633 (O_1633,N_24031,N_22023);
nand UO_1634 (O_1634,N_22293,N_22374);
nor UO_1635 (O_1635,N_22152,N_23617);
and UO_1636 (O_1636,N_21925,N_22053);
or UO_1637 (O_1637,N_22226,N_22759);
xnor UO_1638 (O_1638,N_22670,N_23675);
or UO_1639 (O_1639,N_24289,N_24970);
and UO_1640 (O_1640,N_23612,N_23022);
and UO_1641 (O_1641,N_23492,N_22933);
or UO_1642 (O_1642,N_23588,N_24084);
and UO_1643 (O_1643,N_24015,N_22252);
nor UO_1644 (O_1644,N_23121,N_22063);
or UO_1645 (O_1645,N_22658,N_23946);
xnor UO_1646 (O_1646,N_23864,N_24592);
or UO_1647 (O_1647,N_24693,N_22934);
nand UO_1648 (O_1648,N_22407,N_23388);
or UO_1649 (O_1649,N_23327,N_23174);
xnor UO_1650 (O_1650,N_23874,N_23725);
nand UO_1651 (O_1651,N_24444,N_22386);
nor UO_1652 (O_1652,N_21887,N_24090);
and UO_1653 (O_1653,N_22460,N_23831);
nor UO_1654 (O_1654,N_24920,N_22021);
nor UO_1655 (O_1655,N_22628,N_24037);
xnor UO_1656 (O_1656,N_22931,N_24170);
or UO_1657 (O_1657,N_22356,N_24356);
or UO_1658 (O_1658,N_21890,N_24990);
and UO_1659 (O_1659,N_21912,N_21936);
and UO_1660 (O_1660,N_23354,N_22849);
nor UO_1661 (O_1661,N_21957,N_22943);
nor UO_1662 (O_1662,N_22410,N_24916);
or UO_1663 (O_1663,N_22082,N_24168);
or UO_1664 (O_1664,N_24169,N_22938);
and UO_1665 (O_1665,N_23800,N_24840);
nand UO_1666 (O_1666,N_23728,N_22578);
and UO_1667 (O_1667,N_21938,N_22973);
nand UO_1668 (O_1668,N_23199,N_22760);
nand UO_1669 (O_1669,N_22917,N_24967);
and UO_1670 (O_1670,N_22561,N_22017);
or UO_1671 (O_1671,N_24184,N_22503);
xnor UO_1672 (O_1672,N_23636,N_22476);
and UO_1673 (O_1673,N_23846,N_22302);
nand UO_1674 (O_1674,N_22506,N_24259);
nor UO_1675 (O_1675,N_22199,N_24571);
nand UO_1676 (O_1676,N_23296,N_23247);
or UO_1677 (O_1677,N_22581,N_23294);
nand UO_1678 (O_1678,N_24549,N_22845);
nor UO_1679 (O_1679,N_23309,N_22021);
nor UO_1680 (O_1680,N_22696,N_23977);
xnor UO_1681 (O_1681,N_24093,N_24574);
or UO_1682 (O_1682,N_22590,N_23560);
nand UO_1683 (O_1683,N_23710,N_21973);
or UO_1684 (O_1684,N_22064,N_23922);
and UO_1685 (O_1685,N_22816,N_24644);
and UO_1686 (O_1686,N_22221,N_22610);
nand UO_1687 (O_1687,N_23645,N_23058);
nor UO_1688 (O_1688,N_24702,N_24458);
or UO_1689 (O_1689,N_23853,N_22479);
nand UO_1690 (O_1690,N_24832,N_23267);
nor UO_1691 (O_1691,N_23214,N_23442);
nor UO_1692 (O_1692,N_24661,N_24159);
and UO_1693 (O_1693,N_23700,N_23437);
nor UO_1694 (O_1694,N_22439,N_24585);
nand UO_1695 (O_1695,N_21920,N_24440);
and UO_1696 (O_1696,N_23828,N_23145);
xnor UO_1697 (O_1697,N_21953,N_24175);
or UO_1698 (O_1698,N_22867,N_24202);
xor UO_1699 (O_1699,N_23947,N_22619);
and UO_1700 (O_1700,N_24658,N_22293);
nand UO_1701 (O_1701,N_24582,N_23632);
nand UO_1702 (O_1702,N_22165,N_22390);
xor UO_1703 (O_1703,N_23219,N_23169);
nor UO_1704 (O_1704,N_22898,N_24912);
nor UO_1705 (O_1705,N_23194,N_24687);
nand UO_1706 (O_1706,N_22882,N_23062);
or UO_1707 (O_1707,N_22892,N_24943);
xnor UO_1708 (O_1708,N_23327,N_24977);
xnor UO_1709 (O_1709,N_24200,N_23392);
or UO_1710 (O_1710,N_23049,N_22732);
nand UO_1711 (O_1711,N_22922,N_23790);
xor UO_1712 (O_1712,N_24257,N_23897);
nand UO_1713 (O_1713,N_22299,N_24264);
xnor UO_1714 (O_1714,N_22626,N_23848);
nand UO_1715 (O_1715,N_21888,N_22245);
xnor UO_1716 (O_1716,N_22674,N_22142);
xnor UO_1717 (O_1717,N_24086,N_24326);
or UO_1718 (O_1718,N_24245,N_24853);
nand UO_1719 (O_1719,N_22723,N_23403);
nor UO_1720 (O_1720,N_22840,N_23171);
or UO_1721 (O_1721,N_24709,N_22860);
nand UO_1722 (O_1722,N_23530,N_23162);
nand UO_1723 (O_1723,N_24831,N_22249);
or UO_1724 (O_1724,N_24099,N_22367);
or UO_1725 (O_1725,N_23261,N_24973);
and UO_1726 (O_1726,N_23099,N_22798);
nor UO_1727 (O_1727,N_24074,N_21969);
nand UO_1728 (O_1728,N_22729,N_24358);
or UO_1729 (O_1729,N_22024,N_23763);
or UO_1730 (O_1730,N_22497,N_22492);
xor UO_1731 (O_1731,N_24820,N_23507);
and UO_1732 (O_1732,N_21958,N_22517);
or UO_1733 (O_1733,N_22834,N_22338);
or UO_1734 (O_1734,N_24876,N_22511);
nand UO_1735 (O_1735,N_23069,N_24938);
xor UO_1736 (O_1736,N_22247,N_23771);
nor UO_1737 (O_1737,N_22697,N_24013);
xor UO_1738 (O_1738,N_22257,N_22813);
and UO_1739 (O_1739,N_24102,N_23674);
and UO_1740 (O_1740,N_23310,N_24252);
nor UO_1741 (O_1741,N_22619,N_24015);
or UO_1742 (O_1742,N_22760,N_23061);
or UO_1743 (O_1743,N_24144,N_22066);
nand UO_1744 (O_1744,N_24649,N_24320);
or UO_1745 (O_1745,N_23540,N_22582);
and UO_1746 (O_1746,N_22821,N_21998);
or UO_1747 (O_1747,N_24184,N_23132);
nor UO_1748 (O_1748,N_22419,N_22494);
nand UO_1749 (O_1749,N_23513,N_24753);
or UO_1750 (O_1750,N_23431,N_23724);
nand UO_1751 (O_1751,N_23527,N_22129);
xnor UO_1752 (O_1752,N_24371,N_22129);
xor UO_1753 (O_1753,N_24509,N_22612);
and UO_1754 (O_1754,N_24069,N_24135);
xor UO_1755 (O_1755,N_24737,N_22402);
xnor UO_1756 (O_1756,N_24910,N_24195);
or UO_1757 (O_1757,N_23794,N_24095);
or UO_1758 (O_1758,N_22110,N_22045);
nor UO_1759 (O_1759,N_23391,N_24727);
nand UO_1760 (O_1760,N_22278,N_23950);
nand UO_1761 (O_1761,N_22416,N_21975);
and UO_1762 (O_1762,N_22661,N_22283);
nand UO_1763 (O_1763,N_22733,N_22495);
nor UO_1764 (O_1764,N_23509,N_24299);
xnor UO_1765 (O_1765,N_23526,N_22666);
or UO_1766 (O_1766,N_23239,N_24461);
nand UO_1767 (O_1767,N_23577,N_24430);
nor UO_1768 (O_1768,N_22942,N_24663);
or UO_1769 (O_1769,N_22712,N_24677);
and UO_1770 (O_1770,N_22720,N_22683);
xor UO_1771 (O_1771,N_21901,N_23316);
nand UO_1772 (O_1772,N_22295,N_22711);
nand UO_1773 (O_1773,N_22046,N_22836);
nor UO_1774 (O_1774,N_22480,N_23487);
nand UO_1775 (O_1775,N_22446,N_21882);
xnor UO_1776 (O_1776,N_24801,N_24489);
nand UO_1777 (O_1777,N_23148,N_22318);
xor UO_1778 (O_1778,N_23285,N_22609);
and UO_1779 (O_1779,N_22463,N_24488);
or UO_1780 (O_1780,N_23153,N_24552);
xor UO_1781 (O_1781,N_24255,N_24571);
or UO_1782 (O_1782,N_22267,N_24743);
or UO_1783 (O_1783,N_24487,N_24998);
nand UO_1784 (O_1784,N_22461,N_22524);
or UO_1785 (O_1785,N_24801,N_24352);
or UO_1786 (O_1786,N_24895,N_24006);
and UO_1787 (O_1787,N_24045,N_24796);
and UO_1788 (O_1788,N_22370,N_24566);
xnor UO_1789 (O_1789,N_23451,N_23525);
nand UO_1790 (O_1790,N_22521,N_24933);
xor UO_1791 (O_1791,N_24204,N_23866);
and UO_1792 (O_1792,N_24074,N_24757);
nor UO_1793 (O_1793,N_22820,N_22617);
nor UO_1794 (O_1794,N_23720,N_23482);
or UO_1795 (O_1795,N_24419,N_24087);
or UO_1796 (O_1796,N_23323,N_24989);
and UO_1797 (O_1797,N_22834,N_22660);
and UO_1798 (O_1798,N_23125,N_23515);
nor UO_1799 (O_1799,N_24543,N_24142);
or UO_1800 (O_1800,N_24127,N_22814);
nor UO_1801 (O_1801,N_22482,N_23772);
nand UO_1802 (O_1802,N_24386,N_23328);
xor UO_1803 (O_1803,N_21881,N_23535);
or UO_1804 (O_1804,N_22494,N_24818);
xnor UO_1805 (O_1805,N_22982,N_23603);
nand UO_1806 (O_1806,N_24743,N_24281);
xnor UO_1807 (O_1807,N_22704,N_24409);
and UO_1808 (O_1808,N_22162,N_22857);
and UO_1809 (O_1809,N_23925,N_22078);
xor UO_1810 (O_1810,N_22617,N_21964);
and UO_1811 (O_1811,N_24907,N_22449);
and UO_1812 (O_1812,N_23681,N_23263);
nand UO_1813 (O_1813,N_24090,N_23770);
xor UO_1814 (O_1814,N_24946,N_24957);
nor UO_1815 (O_1815,N_22726,N_23747);
nand UO_1816 (O_1816,N_24282,N_21996);
nor UO_1817 (O_1817,N_22615,N_22398);
nand UO_1818 (O_1818,N_23299,N_23808);
or UO_1819 (O_1819,N_23791,N_24383);
nor UO_1820 (O_1820,N_21896,N_22523);
and UO_1821 (O_1821,N_23304,N_22863);
and UO_1822 (O_1822,N_22435,N_24569);
or UO_1823 (O_1823,N_24908,N_22798);
xnor UO_1824 (O_1824,N_24471,N_23446);
xnor UO_1825 (O_1825,N_22459,N_22133);
xnor UO_1826 (O_1826,N_23925,N_24663);
and UO_1827 (O_1827,N_24248,N_22249);
or UO_1828 (O_1828,N_22021,N_24939);
or UO_1829 (O_1829,N_22966,N_23254);
and UO_1830 (O_1830,N_24792,N_23249);
xor UO_1831 (O_1831,N_24738,N_24961);
and UO_1832 (O_1832,N_22968,N_23359);
nand UO_1833 (O_1833,N_23319,N_23303);
nor UO_1834 (O_1834,N_22145,N_24023);
and UO_1835 (O_1835,N_22980,N_22227);
nor UO_1836 (O_1836,N_23706,N_21877);
nor UO_1837 (O_1837,N_21988,N_22059);
nor UO_1838 (O_1838,N_24574,N_24571);
xnor UO_1839 (O_1839,N_22123,N_24491);
or UO_1840 (O_1840,N_23823,N_21934);
and UO_1841 (O_1841,N_24060,N_22088);
nand UO_1842 (O_1842,N_22361,N_22656);
nor UO_1843 (O_1843,N_24087,N_22395);
nand UO_1844 (O_1844,N_24645,N_23211);
xnor UO_1845 (O_1845,N_23446,N_24175);
nand UO_1846 (O_1846,N_23296,N_22321);
xnor UO_1847 (O_1847,N_22227,N_22759);
and UO_1848 (O_1848,N_24119,N_23687);
or UO_1849 (O_1849,N_24025,N_22296);
and UO_1850 (O_1850,N_23744,N_24037);
nor UO_1851 (O_1851,N_23871,N_24881);
nor UO_1852 (O_1852,N_24748,N_21968);
and UO_1853 (O_1853,N_24074,N_23569);
nor UO_1854 (O_1854,N_23285,N_21907);
and UO_1855 (O_1855,N_23220,N_23559);
xor UO_1856 (O_1856,N_22472,N_22227);
or UO_1857 (O_1857,N_22621,N_24861);
nand UO_1858 (O_1858,N_22364,N_24985);
nor UO_1859 (O_1859,N_22403,N_23748);
nand UO_1860 (O_1860,N_22466,N_24679);
and UO_1861 (O_1861,N_24034,N_24790);
xor UO_1862 (O_1862,N_23332,N_23268);
or UO_1863 (O_1863,N_22445,N_24013);
xor UO_1864 (O_1864,N_24208,N_23306);
xnor UO_1865 (O_1865,N_22022,N_22468);
nor UO_1866 (O_1866,N_22751,N_23432);
or UO_1867 (O_1867,N_23972,N_22270);
or UO_1868 (O_1868,N_24721,N_23853);
nand UO_1869 (O_1869,N_23911,N_22242);
or UO_1870 (O_1870,N_24544,N_21876);
or UO_1871 (O_1871,N_24157,N_22906);
and UO_1872 (O_1872,N_22797,N_23824);
nand UO_1873 (O_1873,N_24110,N_22111);
or UO_1874 (O_1874,N_22994,N_22235);
nand UO_1875 (O_1875,N_23192,N_24155);
or UO_1876 (O_1876,N_24721,N_24715);
and UO_1877 (O_1877,N_24292,N_22131);
nand UO_1878 (O_1878,N_22678,N_23697);
or UO_1879 (O_1879,N_22607,N_24223);
xor UO_1880 (O_1880,N_24530,N_24053);
nand UO_1881 (O_1881,N_23962,N_22600);
xor UO_1882 (O_1882,N_22408,N_24460);
xor UO_1883 (O_1883,N_22448,N_23350);
and UO_1884 (O_1884,N_23000,N_22193);
xor UO_1885 (O_1885,N_24577,N_23961);
nor UO_1886 (O_1886,N_24977,N_23482);
nand UO_1887 (O_1887,N_22730,N_23972);
nand UO_1888 (O_1888,N_23930,N_24655);
and UO_1889 (O_1889,N_22775,N_23958);
xnor UO_1890 (O_1890,N_22318,N_22605);
nand UO_1891 (O_1891,N_24465,N_23183);
nand UO_1892 (O_1892,N_24755,N_24650);
and UO_1893 (O_1893,N_22317,N_24614);
nand UO_1894 (O_1894,N_22677,N_23246);
and UO_1895 (O_1895,N_22313,N_24780);
nand UO_1896 (O_1896,N_23405,N_24010);
and UO_1897 (O_1897,N_22565,N_24018);
nor UO_1898 (O_1898,N_24074,N_22175);
nand UO_1899 (O_1899,N_22940,N_22457);
or UO_1900 (O_1900,N_22027,N_22654);
nand UO_1901 (O_1901,N_23750,N_24743);
and UO_1902 (O_1902,N_24850,N_22686);
or UO_1903 (O_1903,N_23712,N_22466);
and UO_1904 (O_1904,N_24713,N_24737);
or UO_1905 (O_1905,N_23881,N_23649);
or UO_1906 (O_1906,N_23983,N_22895);
nor UO_1907 (O_1907,N_22556,N_22203);
nand UO_1908 (O_1908,N_22448,N_24925);
or UO_1909 (O_1909,N_23255,N_23737);
nor UO_1910 (O_1910,N_23557,N_23258);
xnor UO_1911 (O_1911,N_22714,N_24483);
nor UO_1912 (O_1912,N_23774,N_22877);
nand UO_1913 (O_1913,N_23119,N_24588);
nor UO_1914 (O_1914,N_24132,N_22670);
and UO_1915 (O_1915,N_24794,N_22771);
or UO_1916 (O_1916,N_22466,N_23650);
or UO_1917 (O_1917,N_22326,N_24315);
nor UO_1918 (O_1918,N_22921,N_24026);
nor UO_1919 (O_1919,N_22436,N_23624);
xor UO_1920 (O_1920,N_22706,N_23842);
nor UO_1921 (O_1921,N_22420,N_23497);
nand UO_1922 (O_1922,N_21905,N_24678);
or UO_1923 (O_1923,N_24413,N_24892);
or UO_1924 (O_1924,N_22517,N_22219);
or UO_1925 (O_1925,N_24458,N_22550);
nand UO_1926 (O_1926,N_22496,N_23984);
nor UO_1927 (O_1927,N_22005,N_22778);
and UO_1928 (O_1928,N_22258,N_22561);
nand UO_1929 (O_1929,N_23130,N_23275);
and UO_1930 (O_1930,N_23209,N_24319);
xnor UO_1931 (O_1931,N_24964,N_24572);
or UO_1932 (O_1932,N_22855,N_24725);
nand UO_1933 (O_1933,N_24477,N_24721);
or UO_1934 (O_1934,N_24177,N_22118);
nor UO_1935 (O_1935,N_23397,N_23632);
nor UO_1936 (O_1936,N_24878,N_22846);
xnor UO_1937 (O_1937,N_23611,N_24723);
xnor UO_1938 (O_1938,N_22140,N_22462);
nand UO_1939 (O_1939,N_22403,N_24220);
xnor UO_1940 (O_1940,N_23392,N_23551);
or UO_1941 (O_1941,N_22607,N_24997);
and UO_1942 (O_1942,N_23511,N_22381);
xnor UO_1943 (O_1943,N_22776,N_23634);
xnor UO_1944 (O_1944,N_22786,N_23291);
and UO_1945 (O_1945,N_22686,N_24274);
nor UO_1946 (O_1946,N_24635,N_23032);
or UO_1947 (O_1947,N_24783,N_22153);
xor UO_1948 (O_1948,N_24538,N_23744);
nor UO_1949 (O_1949,N_21984,N_24957);
and UO_1950 (O_1950,N_21974,N_24534);
nand UO_1951 (O_1951,N_24510,N_22769);
nand UO_1952 (O_1952,N_22764,N_23692);
and UO_1953 (O_1953,N_21984,N_22694);
xnor UO_1954 (O_1954,N_22051,N_23171);
nand UO_1955 (O_1955,N_22487,N_21979);
or UO_1956 (O_1956,N_23988,N_22267);
nor UO_1957 (O_1957,N_23718,N_23916);
nor UO_1958 (O_1958,N_23636,N_23174);
xor UO_1959 (O_1959,N_23721,N_23801);
xnor UO_1960 (O_1960,N_23849,N_23495);
or UO_1961 (O_1961,N_24189,N_23893);
nor UO_1962 (O_1962,N_22833,N_22465);
and UO_1963 (O_1963,N_22280,N_22803);
nor UO_1964 (O_1964,N_23150,N_23285);
nand UO_1965 (O_1965,N_24085,N_23825);
nor UO_1966 (O_1966,N_22231,N_24264);
xor UO_1967 (O_1967,N_23038,N_24190);
nand UO_1968 (O_1968,N_24379,N_24483);
nor UO_1969 (O_1969,N_22793,N_24668);
nor UO_1970 (O_1970,N_22387,N_24285);
xor UO_1971 (O_1971,N_22797,N_23668);
nand UO_1972 (O_1972,N_22126,N_22680);
nand UO_1973 (O_1973,N_22415,N_22119);
nor UO_1974 (O_1974,N_24184,N_24307);
and UO_1975 (O_1975,N_23195,N_23900);
xnor UO_1976 (O_1976,N_24589,N_21915);
or UO_1977 (O_1977,N_23407,N_22290);
and UO_1978 (O_1978,N_23283,N_22141);
nor UO_1979 (O_1979,N_24465,N_23007);
nor UO_1980 (O_1980,N_23076,N_24984);
nand UO_1981 (O_1981,N_24221,N_24529);
nand UO_1982 (O_1982,N_23642,N_23292);
xnor UO_1983 (O_1983,N_24079,N_24460);
or UO_1984 (O_1984,N_22052,N_23029);
or UO_1985 (O_1985,N_23971,N_23462);
or UO_1986 (O_1986,N_22351,N_22456);
or UO_1987 (O_1987,N_23704,N_24238);
nand UO_1988 (O_1988,N_22356,N_23469);
xor UO_1989 (O_1989,N_23927,N_24203);
xnor UO_1990 (O_1990,N_22684,N_22822);
nand UO_1991 (O_1991,N_24341,N_22842);
or UO_1992 (O_1992,N_24908,N_23475);
xnor UO_1993 (O_1993,N_23477,N_22832);
nand UO_1994 (O_1994,N_23067,N_22647);
or UO_1995 (O_1995,N_24127,N_22418);
xnor UO_1996 (O_1996,N_21968,N_22454);
or UO_1997 (O_1997,N_24128,N_23195);
or UO_1998 (O_1998,N_22852,N_23191);
nand UO_1999 (O_1999,N_24070,N_21981);
or UO_2000 (O_2000,N_23817,N_23282);
nor UO_2001 (O_2001,N_23756,N_22123);
xnor UO_2002 (O_2002,N_24899,N_24330);
and UO_2003 (O_2003,N_24137,N_21991);
and UO_2004 (O_2004,N_23521,N_23956);
xnor UO_2005 (O_2005,N_23891,N_24426);
nor UO_2006 (O_2006,N_22509,N_24660);
or UO_2007 (O_2007,N_24220,N_24717);
nand UO_2008 (O_2008,N_22606,N_22441);
nor UO_2009 (O_2009,N_23720,N_24920);
and UO_2010 (O_2010,N_21955,N_22539);
xnor UO_2011 (O_2011,N_22167,N_24843);
xnor UO_2012 (O_2012,N_22257,N_22586);
and UO_2013 (O_2013,N_23275,N_24135);
and UO_2014 (O_2014,N_23324,N_22462);
or UO_2015 (O_2015,N_23677,N_24833);
or UO_2016 (O_2016,N_24785,N_24537);
or UO_2017 (O_2017,N_23810,N_24533);
or UO_2018 (O_2018,N_24656,N_24247);
nand UO_2019 (O_2019,N_24381,N_24499);
nor UO_2020 (O_2020,N_23771,N_22605);
nand UO_2021 (O_2021,N_22128,N_24626);
or UO_2022 (O_2022,N_23982,N_23850);
xnor UO_2023 (O_2023,N_24318,N_24133);
or UO_2024 (O_2024,N_22379,N_23578);
or UO_2025 (O_2025,N_24882,N_22658);
nand UO_2026 (O_2026,N_24126,N_22484);
xnor UO_2027 (O_2027,N_24769,N_24165);
xor UO_2028 (O_2028,N_24866,N_22033);
nand UO_2029 (O_2029,N_23492,N_24494);
nand UO_2030 (O_2030,N_22861,N_23798);
nor UO_2031 (O_2031,N_23136,N_23339);
or UO_2032 (O_2032,N_23955,N_22174);
nand UO_2033 (O_2033,N_22261,N_23124);
xor UO_2034 (O_2034,N_23059,N_24162);
nor UO_2035 (O_2035,N_23660,N_21940);
xor UO_2036 (O_2036,N_23776,N_23650);
nand UO_2037 (O_2037,N_23383,N_24586);
nand UO_2038 (O_2038,N_24506,N_22337);
or UO_2039 (O_2039,N_23299,N_23863);
or UO_2040 (O_2040,N_24055,N_22688);
and UO_2041 (O_2041,N_22171,N_22709);
and UO_2042 (O_2042,N_24425,N_22458);
nor UO_2043 (O_2043,N_24419,N_22183);
and UO_2044 (O_2044,N_23737,N_23246);
or UO_2045 (O_2045,N_24877,N_23459);
and UO_2046 (O_2046,N_24603,N_22003);
and UO_2047 (O_2047,N_22826,N_24570);
xor UO_2048 (O_2048,N_22587,N_24861);
or UO_2049 (O_2049,N_24977,N_22102);
xor UO_2050 (O_2050,N_22147,N_23933);
or UO_2051 (O_2051,N_24729,N_24920);
xnor UO_2052 (O_2052,N_22239,N_24356);
xnor UO_2053 (O_2053,N_22697,N_22705);
nand UO_2054 (O_2054,N_23158,N_22480);
nor UO_2055 (O_2055,N_22383,N_21981);
xor UO_2056 (O_2056,N_23085,N_23162);
nand UO_2057 (O_2057,N_23597,N_23867);
nor UO_2058 (O_2058,N_21905,N_24075);
xnor UO_2059 (O_2059,N_22790,N_24087);
nand UO_2060 (O_2060,N_24064,N_23414);
nor UO_2061 (O_2061,N_22815,N_23914);
and UO_2062 (O_2062,N_22748,N_23038);
xor UO_2063 (O_2063,N_23590,N_23057);
nor UO_2064 (O_2064,N_24101,N_24376);
nor UO_2065 (O_2065,N_23920,N_24914);
and UO_2066 (O_2066,N_21988,N_24378);
nand UO_2067 (O_2067,N_24790,N_22491);
or UO_2068 (O_2068,N_23362,N_23977);
nand UO_2069 (O_2069,N_24668,N_23211);
xnor UO_2070 (O_2070,N_24380,N_23565);
and UO_2071 (O_2071,N_23412,N_22853);
or UO_2072 (O_2072,N_23497,N_22774);
and UO_2073 (O_2073,N_22411,N_24724);
and UO_2074 (O_2074,N_24799,N_24008);
or UO_2075 (O_2075,N_24607,N_22522);
and UO_2076 (O_2076,N_24705,N_24434);
nand UO_2077 (O_2077,N_24322,N_23011);
or UO_2078 (O_2078,N_24166,N_22957);
or UO_2079 (O_2079,N_22133,N_24561);
or UO_2080 (O_2080,N_22789,N_24223);
and UO_2081 (O_2081,N_22629,N_22018);
and UO_2082 (O_2082,N_23456,N_21926);
nor UO_2083 (O_2083,N_23842,N_24322);
nor UO_2084 (O_2084,N_24134,N_23956);
and UO_2085 (O_2085,N_23468,N_22570);
nand UO_2086 (O_2086,N_24839,N_22332);
and UO_2087 (O_2087,N_23492,N_23194);
nor UO_2088 (O_2088,N_22752,N_23189);
and UO_2089 (O_2089,N_23266,N_24799);
or UO_2090 (O_2090,N_23703,N_24393);
nand UO_2091 (O_2091,N_23061,N_22126);
or UO_2092 (O_2092,N_21921,N_22051);
or UO_2093 (O_2093,N_24858,N_22308);
or UO_2094 (O_2094,N_23346,N_24136);
xnor UO_2095 (O_2095,N_22568,N_23123);
nand UO_2096 (O_2096,N_22640,N_23660);
and UO_2097 (O_2097,N_22877,N_21964);
or UO_2098 (O_2098,N_23856,N_22845);
or UO_2099 (O_2099,N_24265,N_22544);
xnor UO_2100 (O_2100,N_24634,N_23530);
xor UO_2101 (O_2101,N_23778,N_23131);
xnor UO_2102 (O_2102,N_23581,N_22261);
xnor UO_2103 (O_2103,N_23084,N_23116);
nand UO_2104 (O_2104,N_22906,N_22160);
xor UO_2105 (O_2105,N_22738,N_23675);
xor UO_2106 (O_2106,N_23513,N_24564);
xor UO_2107 (O_2107,N_22792,N_24534);
nor UO_2108 (O_2108,N_22439,N_24188);
or UO_2109 (O_2109,N_22343,N_23336);
nand UO_2110 (O_2110,N_24956,N_24499);
or UO_2111 (O_2111,N_23517,N_23103);
and UO_2112 (O_2112,N_23216,N_23662);
nor UO_2113 (O_2113,N_22368,N_24544);
nand UO_2114 (O_2114,N_22924,N_24789);
and UO_2115 (O_2115,N_24996,N_22790);
nand UO_2116 (O_2116,N_22151,N_23294);
and UO_2117 (O_2117,N_24880,N_22923);
nor UO_2118 (O_2118,N_24075,N_22588);
or UO_2119 (O_2119,N_24699,N_24516);
or UO_2120 (O_2120,N_22627,N_22750);
nor UO_2121 (O_2121,N_24590,N_24979);
and UO_2122 (O_2122,N_24053,N_23399);
nand UO_2123 (O_2123,N_22504,N_21970);
xor UO_2124 (O_2124,N_23549,N_23495);
or UO_2125 (O_2125,N_23847,N_23295);
nand UO_2126 (O_2126,N_24633,N_23209);
xor UO_2127 (O_2127,N_23627,N_24456);
and UO_2128 (O_2128,N_22724,N_24351);
nor UO_2129 (O_2129,N_22664,N_24374);
nand UO_2130 (O_2130,N_24385,N_23568);
or UO_2131 (O_2131,N_22151,N_22883);
nand UO_2132 (O_2132,N_22619,N_22055);
xnor UO_2133 (O_2133,N_23256,N_22362);
nor UO_2134 (O_2134,N_22195,N_23127);
nor UO_2135 (O_2135,N_22816,N_22511);
xnor UO_2136 (O_2136,N_21966,N_23872);
nor UO_2137 (O_2137,N_22462,N_23272);
nand UO_2138 (O_2138,N_22073,N_22480);
nand UO_2139 (O_2139,N_21964,N_22979);
nand UO_2140 (O_2140,N_23022,N_24281);
xor UO_2141 (O_2141,N_22007,N_24297);
and UO_2142 (O_2142,N_24610,N_23195);
or UO_2143 (O_2143,N_24793,N_22216);
nor UO_2144 (O_2144,N_24180,N_24037);
xor UO_2145 (O_2145,N_24946,N_23505);
and UO_2146 (O_2146,N_24466,N_24119);
nor UO_2147 (O_2147,N_22836,N_22396);
nor UO_2148 (O_2148,N_23892,N_22237);
nor UO_2149 (O_2149,N_23234,N_22597);
xor UO_2150 (O_2150,N_22075,N_22216);
and UO_2151 (O_2151,N_24079,N_23005);
and UO_2152 (O_2152,N_22763,N_22933);
nor UO_2153 (O_2153,N_23518,N_22719);
and UO_2154 (O_2154,N_24569,N_24323);
xnor UO_2155 (O_2155,N_24602,N_22100);
nor UO_2156 (O_2156,N_23826,N_22525);
nor UO_2157 (O_2157,N_22997,N_24750);
and UO_2158 (O_2158,N_24528,N_24169);
nor UO_2159 (O_2159,N_23302,N_23062);
nand UO_2160 (O_2160,N_23199,N_24197);
nand UO_2161 (O_2161,N_24668,N_22329);
nand UO_2162 (O_2162,N_22144,N_23063);
nor UO_2163 (O_2163,N_24894,N_24116);
nor UO_2164 (O_2164,N_22595,N_22235);
nor UO_2165 (O_2165,N_22632,N_22115);
xor UO_2166 (O_2166,N_24468,N_22423);
nor UO_2167 (O_2167,N_24692,N_23674);
or UO_2168 (O_2168,N_22833,N_22800);
xor UO_2169 (O_2169,N_24117,N_24426);
xnor UO_2170 (O_2170,N_24385,N_23171);
nand UO_2171 (O_2171,N_24630,N_24175);
or UO_2172 (O_2172,N_24863,N_23472);
or UO_2173 (O_2173,N_23734,N_23687);
or UO_2174 (O_2174,N_23676,N_23831);
nand UO_2175 (O_2175,N_24929,N_24479);
and UO_2176 (O_2176,N_24669,N_22051);
nand UO_2177 (O_2177,N_23570,N_23328);
xnor UO_2178 (O_2178,N_22895,N_23558);
nor UO_2179 (O_2179,N_22882,N_22342);
xor UO_2180 (O_2180,N_22515,N_23687);
nand UO_2181 (O_2181,N_23646,N_23432);
xor UO_2182 (O_2182,N_22031,N_23226);
xor UO_2183 (O_2183,N_21887,N_23093);
or UO_2184 (O_2184,N_24678,N_23203);
xnor UO_2185 (O_2185,N_24068,N_24740);
nor UO_2186 (O_2186,N_22418,N_23868);
and UO_2187 (O_2187,N_22353,N_24885);
or UO_2188 (O_2188,N_22837,N_24058);
nor UO_2189 (O_2189,N_24829,N_24704);
xnor UO_2190 (O_2190,N_22963,N_24836);
xnor UO_2191 (O_2191,N_23565,N_22508);
and UO_2192 (O_2192,N_23582,N_22793);
or UO_2193 (O_2193,N_24432,N_23093);
nor UO_2194 (O_2194,N_22408,N_24943);
or UO_2195 (O_2195,N_23426,N_23158);
or UO_2196 (O_2196,N_22459,N_24933);
nor UO_2197 (O_2197,N_24463,N_22430);
and UO_2198 (O_2198,N_22956,N_24074);
nand UO_2199 (O_2199,N_22975,N_24037);
nand UO_2200 (O_2200,N_24404,N_21898);
or UO_2201 (O_2201,N_24107,N_24488);
and UO_2202 (O_2202,N_23609,N_24561);
and UO_2203 (O_2203,N_24692,N_24629);
nand UO_2204 (O_2204,N_24707,N_23978);
nand UO_2205 (O_2205,N_22718,N_24713);
and UO_2206 (O_2206,N_22527,N_24777);
and UO_2207 (O_2207,N_23426,N_23477);
and UO_2208 (O_2208,N_23251,N_22493);
xor UO_2209 (O_2209,N_21921,N_22641);
or UO_2210 (O_2210,N_22040,N_22664);
nand UO_2211 (O_2211,N_22708,N_22365);
or UO_2212 (O_2212,N_24690,N_23285);
nor UO_2213 (O_2213,N_24613,N_24348);
xnor UO_2214 (O_2214,N_23552,N_24748);
or UO_2215 (O_2215,N_23353,N_23990);
xor UO_2216 (O_2216,N_24726,N_24254);
nand UO_2217 (O_2217,N_24694,N_23268);
xnor UO_2218 (O_2218,N_23010,N_22447);
xor UO_2219 (O_2219,N_23535,N_24726);
or UO_2220 (O_2220,N_22132,N_22081);
xnor UO_2221 (O_2221,N_24608,N_22629);
nand UO_2222 (O_2222,N_23200,N_24636);
or UO_2223 (O_2223,N_24363,N_24997);
and UO_2224 (O_2224,N_23917,N_23097);
and UO_2225 (O_2225,N_22453,N_23545);
or UO_2226 (O_2226,N_24598,N_22841);
or UO_2227 (O_2227,N_22638,N_23017);
nor UO_2228 (O_2228,N_23145,N_23704);
xor UO_2229 (O_2229,N_22138,N_22946);
xnor UO_2230 (O_2230,N_23254,N_22106);
and UO_2231 (O_2231,N_24587,N_24394);
xor UO_2232 (O_2232,N_23790,N_24184);
or UO_2233 (O_2233,N_23358,N_21890);
or UO_2234 (O_2234,N_24643,N_22837);
nand UO_2235 (O_2235,N_23898,N_22923);
or UO_2236 (O_2236,N_24276,N_23376);
and UO_2237 (O_2237,N_22759,N_23043);
or UO_2238 (O_2238,N_23853,N_23803);
and UO_2239 (O_2239,N_24936,N_23540);
xnor UO_2240 (O_2240,N_24370,N_24488);
nor UO_2241 (O_2241,N_23833,N_21895);
nor UO_2242 (O_2242,N_22632,N_23062);
or UO_2243 (O_2243,N_23862,N_22603);
nand UO_2244 (O_2244,N_23772,N_22312);
xor UO_2245 (O_2245,N_23320,N_23595);
and UO_2246 (O_2246,N_22989,N_22781);
nand UO_2247 (O_2247,N_23306,N_23996);
nor UO_2248 (O_2248,N_23416,N_23902);
xor UO_2249 (O_2249,N_23382,N_22671);
xnor UO_2250 (O_2250,N_22622,N_22174);
nor UO_2251 (O_2251,N_22076,N_24309);
nor UO_2252 (O_2252,N_22524,N_22212);
nor UO_2253 (O_2253,N_23426,N_24582);
xnor UO_2254 (O_2254,N_24420,N_24884);
nor UO_2255 (O_2255,N_23966,N_23839);
or UO_2256 (O_2256,N_24496,N_23568);
nand UO_2257 (O_2257,N_24725,N_24271);
or UO_2258 (O_2258,N_23910,N_23576);
nand UO_2259 (O_2259,N_23246,N_24646);
nor UO_2260 (O_2260,N_23652,N_21958);
nor UO_2261 (O_2261,N_22490,N_23113);
nor UO_2262 (O_2262,N_22152,N_23391);
nor UO_2263 (O_2263,N_24561,N_21897);
nand UO_2264 (O_2264,N_21903,N_23418);
and UO_2265 (O_2265,N_23446,N_24916);
nor UO_2266 (O_2266,N_24000,N_23614);
or UO_2267 (O_2267,N_23965,N_24316);
nand UO_2268 (O_2268,N_24356,N_24851);
nand UO_2269 (O_2269,N_23220,N_22947);
and UO_2270 (O_2270,N_23622,N_22116);
and UO_2271 (O_2271,N_22641,N_23948);
nor UO_2272 (O_2272,N_22323,N_23289);
nand UO_2273 (O_2273,N_22924,N_22079);
and UO_2274 (O_2274,N_24232,N_24455);
nand UO_2275 (O_2275,N_23944,N_23060);
xor UO_2276 (O_2276,N_24436,N_24802);
xor UO_2277 (O_2277,N_22220,N_24581);
nand UO_2278 (O_2278,N_22281,N_24460);
and UO_2279 (O_2279,N_22351,N_22158);
nand UO_2280 (O_2280,N_24947,N_22602);
nor UO_2281 (O_2281,N_24874,N_23395);
nor UO_2282 (O_2282,N_24151,N_22474);
xnor UO_2283 (O_2283,N_23641,N_23413);
nand UO_2284 (O_2284,N_24882,N_22693);
nand UO_2285 (O_2285,N_22419,N_23205);
xnor UO_2286 (O_2286,N_24164,N_22231);
nand UO_2287 (O_2287,N_24859,N_22342);
and UO_2288 (O_2288,N_22410,N_24716);
nand UO_2289 (O_2289,N_23186,N_24137);
nor UO_2290 (O_2290,N_22989,N_22758);
nor UO_2291 (O_2291,N_23947,N_22130);
nor UO_2292 (O_2292,N_22668,N_23168);
xor UO_2293 (O_2293,N_22516,N_22658);
xnor UO_2294 (O_2294,N_23017,N_24277);
nand UO_2295 (O_2295,N_22520,N_23456);
or UO_2296 (O_2296,N_22625,N_22173);
xnor UO_2297 (O_2297,N_24035,N_22876);
nor UO_2298 (O_2298,N_23560,N_22875);
or UO_2299 (O_2299,N_23791,N_24368);
and UO_2300 (O_2300,N_22493,N_23306);
nor UO_2301 (O_2301,N_24865,N_23209);
nor UO_2302 (O_2302,N_24233,N_24814);
xnor UO_2303 (O_2303,N_24497,N_23783);
and UO_2304 (O_2304,N_23702,N_24466);
and UO_2305 (O_2305,N_24821,N_22349);
nor UO_2306 (O_2306,N_23467,N_24423);
nand UO_2307 (O_2307,N_23024,N_24570);
nor UO_2308 (O_2308,N_22068,N_23266);
nor UO_2309 (O_2309,N_23639,N_24180);
and UO_2310 (O_2310,N_21887,N_23746);
xor UO_2311 (O_2311,N_22331,N_24938);
xor UO_2312 (O_2312,N_24022,N_22499);
nand UO_2313 (O_2313,N_23178,N_23982);
xnor UO_2314 (O_2314,N_22741,N_22299);
and UO_2315 (O_2315,N_22808,N_24442);
or UO_2316 (O_2316,N_23084,N_24828);
and UO_2317 (O_2317,N_23518,N_24554);
xor UO_2318 (O_2318,N_22371,N_23682);
nor UO_2319 (O_2319,N_22403,N_24124);
and UO_2320 (O_2320,N_22905,N_22325);
nand UO_2321 (O_2321,N_22321,N_24272);
or UO_2322 (O_2322,N_24173,N_22723);
nor UO_2323 (O_2323,N_24850,N_22085);
xnor UO_2324 (O_2324,N_24717,N_22294);
or UO_2325 (O_2325,N_23895,N_24133);
and UO_2326 (O_2326,N_23138,N_23885);
nand UO_2327 (O_2327,N_22654,N_24340);
nor UO_2328 (O_2328,N_23991,N_22237);
or UO_2329 (O_2329,N_23346,N_24256);
nor UO_2330 (O_2330,N_22130,N_24161);
nor UO_2331 (O_2331,N_24019,N_22525);
and UO_2332 (O_2332,N_22484,N_24619);
nand UO_2333 (O_2333,N_23734,N_24484);
or UO_2334 (O_2334,N_23804,N_22378);
and UO_2335 (O_2335,N_24770,N_23632);
or UO_2336 (O_2336,N_23822,N_24879);
nor UO_2337 (O_2337,N_23903,N_22271);
nand UO_2338 (O_2338,N_22747,N_23911);
nor UO_2339 (O_2339,N_24153,N_23568);
nor UO_2340 (O_2340,N_23100,N_22288);
and UO_2341 (O_2341,N_23221,N_23819);
or UO_2342 (O_2342,N_22584,N_21901);
and UO_2343 (O_2343,N_22775,N_24112);
and UO_2344 (O_2344,N_24270,N_24658);
or UO_2345 (O_2345,N_23090,N_22958);
nor UO_2346 (O_2346,N_22517,N_23199);
or UO_2347 (O_2347,N_22122,N_23575);
nor UO_2348 (O_2348,N_23080,N_24807);
nor UO_2349 (O_2349,N_23183,N_23127);
or UO_2350 (O_2350,N_24631,N_24099);
or UO_2351 (O_2351,N_24581,N_22485);
nand UO_2352 (O_2352,N_22254,N_23823);
nor UO_2353 (O_2353,N_23205,N_23034);
and UO_2354 (O_2354,N_24933,N_22131);
xor UO_2355 (O_2355,N_22256,N_23436);
nor UO_2356 (O_2356,N_23127,N_22759);
nor UO_2357 (O_2357,N_22232,N_23087);
nor UO_2358 (O_2358,N_24079,N_22517);
or UO_2359 (O_2359,N_22127,N_24107);
nand UO_2360 (O_2360,N_23458,N_24755);
xnor UO_2361 (O_2361,N_23328,N_24583);
or UO_2362 (O_2362,N_23749,N_23760);
and UO_2363 (O_2363,N_24151,N_22253);
or UO_2364 (O_2364,N_24485,N_23623);
and UO_2365 (O_2365,N_23036,N_24588);
xor UO_2366 (O_2366,N_23769,N_24679);
or UO_2367 (O_2367,N_24328,N_24090);
xnor UO_2368 (O_2368,N_24316,N_23612);
xor UO_2369 (O_2369,N_23209,N_22419);
and UO_2370 (O_2370,N_24241,N_23427);
nor UO_2371 (O_2371,N_23398,N_24737);
or UO_2372 (O_2372,N_23024,N_23953);
and UO_2373 (O_2373,N_23328,N_22032);
nor UO_2374 (O_2374,N_24011,N_23492);
xnor UO_2375 (O_2375,N_24313,N_22409);
and UO_2376 (O_2376,N_24848,N_22157);
or UO_2377 (O_2377,N_23868,N_23478);
xor UO_2378 (O_2378,N_23451,N_23845);
or UO_2379 (O_2379,N_23783,N_24960);
nand UO_2380 (O_2380,N_22404,N_22726);
xor UO_2381 (O_2381,N_22289,N_23891);
nand UO_2382 (O_2382,N_24924,N_22609);
nand UO_2383 (O_2383,N_22176,N_23522);
nor UO_2384 (O_2384,N_22378,N_23222);
or UO_2385 (O_2385,N_23836,N_22484);
nand UO_2386 (O_2386,N_23748,N_24628);
or UO_2387 (O_2387,N_22432,N_23708);
nand UO_2388 (O_2388,N_24282,N_24257);
nand UO_2389 (O_2389,N_22945,N_22425);
nand UO_2390 (O_2390,N_22635,N_22397);
xnor UO_2391 (O_2391,N_22276,N_23934);
and UO_2392 (O_2392,N_23012,N_23346);
nand UO_2393 (O_2393,N_23216,N_23724);
and UO_2394 (O_2394,N_24004,N_23266);
or UO_2395 (O_2395,N_22926,N_23237);
xor UO_2396 (O_2396,N_21953,N_24287);
and UO_2397 (O_2397,N_22379,N_24785);
or UO_2398 (O_2398,N_24011,N_23856);
xnor UO_2399 (O_2399,N_22324,N_24100);
and UO_2400 (O_2400,N_21985,N_23502);
xnor UO_2401 (O_2401,N_23745,N_24505);
nand UO_2402 (O_2402,N_24073,N_24876);
nand UO_2403 (O_2403,N_22388,N_24233);
or UO_2404 (O_2404,N_22411,N_23585);
and UO_2405 (O_2405,N_23907,N_22689);
nor UO_2406 (O_2406,N_24448,N_21900);
or UO_2407 (O_2407,N_24312,N_23942);
xnor UO_2408 (O_2408,N_24820,N_22028);
nand UO_2409 (O_2409,N_23802,N_22802);
and UO_2410 (O_2410,N_24515,N_24347);
or UO_2411 (O_2411,N_22535,N_24895);
and UO_2412 (O_2412,N_24569,N_24020);
or UO_2413 (O_2413,N_23881,N_24466);
and UO_2414 (O_2414,N_23584,N_22324);
nor UO_2415 (O_2415,N_22395,N_23552);
nand UO_2416 (O_2416,N_22184,N_22675);
xor UO_2417 (O_2417,N_24921,N_23500);
xor UO_2418 (O_2418,N_21944,N_23335);
xor UO_2419 (O_2419,N_23310,N_24201);
nand UO_2420 (O_2420,N_22338,N_24483);
and UO_2421 (O_2421,N_23296,N_23931);
nor UO_2422 (O_2422,N_24852,N_23088);
xnor UO_2423 (O_2423,N_24554,N_23994);
or UO_2424 (O_2424,N_23903,N_22750);
nand UO_2425 (O_2425,N_24697,N_23388);
nor UO_2426 (O_2426,N_23734,N_24958);
xor UO_2427 (O_2427,N_24433,N_22926);
nor UO_2428 (O_2428,N_22015,N_21905);
xnor UO_2429 (O_2429,N_24133,N_22416);
nand UO_2430 (O_2430,N_24992,N_23991);
or UO_2431 (O_2431,N_24566,N_22170);
or UO_2432 (O_2432,N_22840,N_22048);
nor UO_2433 (O_2433,N_22008,N_24467);
nand UO_2434 (O_2434,N_23021,N_23250);
and UO_2435 (O_2435,N_24553,N_23618);
nor UO_2436 (O_2436,N_22634,N_24479);
nand UO_2437 (O_2437,N_23000,N_24260);
nand UO_2438 (O_2438,N_24289,N_21901);
or UO_2439 (O_2439,N_24076,N_23383);
nor UO_2440 (O_2440,N_24186,N_23073);
nor UO_2441 (O_2441,N_23071,N_22633);
or UO_2442 (O_2442,N_24366,N_22762);
xnor UO_2443 (O_2443,N_24369,N_24011);
nor UO_2444 (O_2444,N_21980,N_22508);
xnor UO_2445 (O_2445,N_23938,N_24186);
and UO_2446 (O_2446,N_24998,N_22020);
and UO_2447 (O_2447,N_23752,N_23564);
nor UO_2448 (O_2448,N_22138,N_22473);
nand UO_2449 (O_2449,N_24259,N_23699);
xnor UO_2450 (O_2450,N_23748,N_24826);
nor UO_2451 (O_2451,N_22189,N_24102);
nor UO_2452 (O_2452,N_23382,N_21961);
or UO_2453 (O_2453,N_22361,N_24911);
nand UO_2454 (O_2454,N_24789,N_22686);
nor UO_2455 (O_2455,N_23846,N_22685);
xnor UO_2456 (O_2456,N_24671,N_22989);
or UO_2457 (O_2457,N_22035,N_23029);
nand UO_2458 (O_2458,N_24657,N_22709);
nand UO_2459 (O_2459,N_24594,N_22504);
nand UO_2460 (O_2460,N_22864,N_24951);
nand UO_2461 (O_2461,N_21903,N_22047);
nor UO_2462 (O_2462,N_21892,N_21925);
nand UO_2463 (O_2463,N_23422,N_22369);
xor UO_2464 (O_2464,N_22227,N_24879);
or UO_2465 (O_2465,N_22218,N_22610);
nor UO_2466 (O_2466,N_24196,N_22991);
and UO_2467 (O_2467,N_21969,N_22848);
nor UO_2468 (O_2468,N_24653,N_24476);
nand UO_2469 (O_2469,N_23299,N_22706);
nor UO_2470 (O_2470,N_23674,N_24424);
nand UO_2471 (O_2471,N_23044,N_24940);
or UO_2472 (O_2472,N_23935,N_23283);
xor UO_2473 (O_2473,N_22315,N_22071);
or UO_2474 (O_2474,N_21988,N_24078);
or UO_2475 (O_2475,N_21960,N_23222);
nor UO_2476 (O_2476,N_22775,N_22043);
nand UO_2477 (O_2477,N_23497,N_22792);
nand UO_2478 (O_2478,N_22477,N_24013);
nand UO_2479 (O_2479,N_23942,N_24713);
nor UO_2480 (O_2480,N_24864,N_24865);
and UO_2481 (O_2481,N_23317,N_23176);
xnor UO_2482 (O_2482,N_22582,N_22581);
or UO_2483 (O_2483,N_22795,N_24584);
xor UO_2484 (O_2484,N_22089,N_22685);
nor UO_2485 (O_2485,N_22195,N_24603);
nand UO_2486 (O_2486,N_23830,N_24838);
and UO_2487 (O_2487,N_24291,N_24591);
and UO_2488 (O_2488,N_23774,N_22598);
or UO_2489 (O_2489,N_22479,N_24581);
nand UO_2490 (O_2490,N_22446,N_24695);
and UO_2491 (O_2491,N_24625,N_21924);
xnor UO_2492 (O_2492,N_24964,N_22175);
nand UO_2493 (O_2493,N_22766,N_24626);
or UO_2494 (O_2494,N_23608,N_22448);
and UO_2495 (O_2495,N_22440,N_23683);
nor UO_2496 (O_2496,N_22345,N_22029);
xnor UO_2497 (O_2497,N_23320,N_21974);
nand UO_2498 (O_2498,N_22360,N_23295);
xnor UO_2499 (O_2499,N_22403,N_23638);
nor UO_2500 (O_2500,N_23851,N_23388);
or UO_2501 (O_2501,N_24348,N_21916);
xnor UO_2502 (O_2502,N_24461,N_23263);
xnor UO_2503 (O_2503,N_22391,N_23603);
nor UO_2504 (O_2504,N_23230,N_22678);
xor UO_2505 (O_2505,N_22320,N_22845);
xor UO_2506 (O_2506,N_22462,N_23714);
or UO_2507 (O_2507,N_22960,N_23956);
nor UO_2508 (O_2508,N_22271,N_24168);
nor UO_2509 (O_2509,N_23992,N_22455);
nand UO_2510 (O_2510,N_22576,N_23189);
or UO_2511 (O_2511,N_22032,N_22898);
nand UO_2512 (O_2512,N_23500,N_22347);
or UO_2513 (O_2513,N_22512,N_22356);
or UO_2514 (O_2514,N_23758,N_22316);
or UO_2515 (O_2515,N_24533,N_24653);
nor UO_2516 (O_2516,N_22027,N_24971);
and UO_2517 (O_2517,N_22721,N_24316);
or UO_2518 (O_2518,N_22721,N_24889);
and UO_2519 (O_2519,N_23488,N_22838);
and UO_2520 (O_2520,N_24208,N_23968);
xnor UO_2521 (O_2521,N_24118,N_24389);
nor UO_2522 (O_2522,N_22585,N_23955);
nand UO_2523 (O_2523,N_22034,N_23428);
nor UO_2524 (O_2524,N_22320,N_21916);
nand UO_2525 (O_2525,N_23507,N_22231);
and UO_2526 (O_2526,N_24308,N_24663);
and UO_2527 (O_2527,N_23831,N_23103);
xor UO_2528 (O_2528,N_24559,N_23753);
nor UO_2529 (O_2529,N_22505,N_22283);
nand UO_2530 (O_2530,N_22412,N_24970);
nor UO_2531 (O_2531,N_23114,N_24793);
nand UO_2532 (O_2532,N_22743,N_22184);
or UO_2533 (O_2533,N_24897,N_23939);
or UO_2534 (O_2534,N_21951,N_23072);
nor UO_2535 (O_2535,N_23825,N_24237);
and UO_2536 (O_2536,N_22711,N_23687);
xnor UO_2537 (O_2537,N_22962,N_23027);
nand UO_2538 (O_2538,N_22519,N_22392);
and UO_2539 (O_2539,N_22318,N_22388);
or UO_2540 (O_2540,N_24094,N_23587);
or UO_2541 (O_2541,N_24737,N_23991);
and UO_2542 (O_2542,N_24728,N_22016);
and UO_2543 (O_2543,N_21942,N_22803);
nand UO_2544 (O_2544,N_24436,N_23259);
nor UO_2545 (O_2545,N_23862,N_23194);
or UO_2546 (O_2546,N_22844,N_24631);
or UO_2547 (O_2547,N_23673,N_24963);
xnor UO_2548 (O_2548,N_22352,N_22039);
xor UO_2549 (O_2549,N_24382,N_24896);
nand UO_2550 (O_2550,N_23045,N_24655);
or UO_2551 (O_2551,N_24128,N_22993);
nor UO_2552 (O_2552,N_23669,N_22908);
and UO_2553 (O_2553,N_24137,N_23911);
nand UO_2554 (O_2554,N_22253,N_24103);
or UO_2555 (O_2555,N_21973,N_24824);
xor UO_2556 (O_2556,N_24661,N_24098);
nand UO_2557 (O_2557,N_23205,N_24159);
nand UO_2558 (O_2558,N_22588,N_23632);
xnor UO_2559 (O_2559,N_24556,N_23410);
xnor UO_2560 (O_2560,N_24529,N_22731);
and UO_2561 (O_2561,N_23423,N_22897);
nand UO_2562 (O_2562,N_23884,N_22241);
or UO_2563 (O_2563,N_23103,N_22228);
xor UO_2564 (O_2564,N_23108,N_24598);
or UO_2565 (O_2565,N_23090,N_22960);
xnor UO_2566 (O_2566,N_22517,N_23636);
nor UO_2567 (O_2567,N_23233,N_22102);
and UO_2568 (O_2568,N_22893,N_22126);
nor UO_2569 (O_2569,N_21881,N_24315);
nand UO_2570 (O_2570,N_22908,N_24277);
nand UO_2571 (O_2571,N_23304,N_22245);
nand UO_2572 (O_2572,N_22362,N_24683);
and UO_2573 (O_2573,N_23135,N_22441);
and UO_2574 (O_2574,N_23730,N_22186);
xor UO_2575 (O_2575,N_22459,N_24298);
nor UO_2576 (O_2576,N_22642,N_23387);
nand UO_2577 (O_2577,N_23107,N_24042);
nor UO_2578 (O_2578,N_22903,N_22124);
xor UO_2579 (O_2579,N_22070,N_22188);
and UO_2580 (O_2580,N_24199,N_22139);
xnor UO_2581 (O_2581,N_23103,N_22679);
xnor UO_2582 (O_2582,N_22981,N_22360);
nand UO_2583 (O_2583,N_22028,N_23160);
nor UO_2584 (O_2584,N_22129,N_23026);
nor UO_2585 (O_2585,N_22181,N_22275);
or UO_2586 (O_2586,N_23040,N_21927);
xor UO_2587 (O_2587,N_22883,N_23132);
xor UO_2588 (O_2588,N_23249,N_23515);
or UO_2589 (O_2589,N_22069,N_24598);
nand UO_2590 (O_2590,N_23261,N_23245);
nand UO_2591 (O_2591,N_22155,N_22177);
nand UO_2592 (O_2592,N_23436,N_22173);
xor UO_2593 (O_2593,N_22348,N_24087);
or UO_2594 (O_2594,N_24704,N_23147);
and UO_2595 (O_2595,N_24480,N_21883);
and UO_2596 (O_2596,N_24615,N_24317);
xor UO_2597 (O_2597,N_23488,N_22668);
and UO_2598 (O_2598,N_22676,N_22269);
or UO_2599 (O_2599,N_24097,N_24520);
or UO_2600 (O_2600,N_22338,N_23856);
or UO_2601 (O_2601,N_23199,N_24726);
nor UO_2602 (O_2602,N_23726,N_24147);
or UO_2603 (O_2603,N_23480,N_24443);
and UO_2604 (O_2604,N_23824,N_22080);
nor UO_2605 (O_2605,N_23782,N_22385);
and UO_2606 (O_2606,N_23455,N_23138);
or UO_2607 (O_2607,N_22734,N_24983);
nand UO_2608 (O_2608,N_24760,N_23945);
nor UO_2609 (O_2609,N_21945,N_22247);
and UO_2610 (O_2610,N_22661,N_23668);
or UO_2611 (O_2611,N_23774,N_23893);
nand UO_2612 (O_2612,N_23347,N_22625);
nand UO_2613 (O_2613,N_23377,N_23524);
xnor UO_2614 (O_2614,N_24641,N_22021);
and UO_2615 (O_2615,N_23804,N_24767);
nand UO_2616 (O_2616,N_23968,N_22896);
xor UO_2617 (O_2617,N_21930,N_22085);
or UO_2618 (O_2618,N_22051,N_23507);
nor UO_2619 (O_2619,N_22923,N_24901);
nor UO_2620 (O_2620,N_22773,N_22101);
and UO_2621 (O_2621,N_22882,N_22753);
and UO_2622 (O_2622,N_24965,N_24610);
nand UO_2623 (O_2623,N_23019,N_24742);
nor UO_2624 (O_2624,N_24842,N_22164);
nor UO_2625 (O_2625,N_22325,N_22552);
and UO_2626 (O_2626,N_24222,N_23707);
xor UO_2627 (O_2627,N_24285,N_22983);
nand UO_2628 (O_2628,N_24135,N_21955);
nor UO_2629 (O_2629,N_23883,N_22595);
nand UO_2630 (O_2630,N_24209,N_23975);
and UO_2631 (O_2631,N_23022,N_24145);
or UO_2632 (O_2632,N_24591,N_23235);
xor UO_2633 (O_2633,N_24594,N_24390);
nor UO_2634 (O_2634,N_22683,N_22359);
nand UO_2635 (O_2635,N_23894,N_22668);
and UO_2636 (O_2636,N_24181,N_24124);
xor UO_2637 (O_2637,N_21962,N_22423);
or UO_2638 (O_2638,N_23032,N_21904);
nand UO_2639 (O_2639,N_24535,N_24184);
and UO_2640 (O_2640,N_23570,N_24386);
or UO_2641 (O_2641,N_22860,N_24870);
or UO_2642 (O_2642,N_23796,N_22592);
and UO_2643 (O_2643,N_22935,N_22156);
nand UO_2644 (O_2644,N_24780,N_24669);
or UO_2645 (O_2645,N_24729,N_21997);
or UO_2646 (O_2646,N_23548,N_21875);
or UO_2647 (O_2647,N_24507,N_22844);
and UO_2648 (O_2648,N_24863,N_24938);
nor UO_2649 (O_2649,N_24118,N_22211);
xnor UO_2650 (O_2650,N_23356,N_23701);
and UO_2651 (O_2651,N_24093,N_24647);
or UO_2652 (O_2652,N_22866,N_24233);
nor UO_2653 (O_2653,N_24941,N_22526);
nor UO_2654 (O_2654,N_22280,N_22628);
nand UO_2655 (O_2655,N_24682,N_23306);
and UO_2656 (O_2656,N_22321,N_22804);
nand UO_2657 (O_2657,N_24372,N_24064);
or UO_2658 (O_2658,N_22664,N_24301);
nor UO_2659 (O_2659,N_22574,N_23558);
nor UO_2660 (O_2660,N_23240,N_22136);
and UO_2661 (O_2661,N_22610,N_22106);
and UO_2662 (O_2662,N_23175,N_23923);
nor UO_2663 (O_2663,N_23985,N_22577);
or UO_2664 (O_2664,N_24338,N_23653);
nor UO_2665 (O_2665,N_22367,N_23199);
nor UO_2666 (O_2666,N_23170,N_23368);
or UO_2667 (O_2667,N_23902,N_22976);
and UO_2668 (O_2668,N_22266,N_23005);
nor UO_2669 (O_2669,N_22960,N_24740);
xnor UO_2670 (O_2670,N_24770,N_24408);
nand UO_2671 (O_2671,N_22863,N_21992);
and UO_2672 (O_2672,N_23498,N_22650);
nand UO_2673 (O_2673,N_24217,N_24772);
nor UO_2674 (O_2674,N_23274,N_22901);
or UO_2675 (O_2675,N_24510,N_24750);
nor UO_2676 (O_2676,N_23490,N_23502);
xnor UO_2677 (O_2677,N_22052,N_23264);
and UO_2678 (O_2678,N_22969,N_22330);
xnor UO_2679 (O_2679,N_24940,N_22559);
nand UO_2680 (O_2680,N_24847,N_22862);
or UO_2681 (O_2681,N_24396,N_22355);
nand UO_2682 (O_2682,N_23981,N_22757);
nor UO_2683 (O_2683,N_23404,N_24212);
or UO_2684 (O_2684,N_23152,N_22234);
or UO_2685 (O_2685,N_24568,N_23882);
and UO_2686 (O_2686,N_22988,N_21913);
or UO_2687 (O_2687,N_24795,N_24021);
and UO_2688 (O_2688,N_22834,N_24389);
or UO_2689 (O_2689,N_23850,N_24607);
or UO_2690 (O_2690,N_22316,N_22784);
xor UO_2691 (O_2691,N_23862,N_23386);
or UO_2692 (O_2692,N_23163,N_23533);
or UO_2693 (O_2693,N_24744,N_22190);
xnor UO_2694 (O_2694,N_24390,N_24386);
or UO_2695 (O_2695,N_24002,N_24958);
or UO_2696 (O_2696,N_21888,N_24680);
and UO_2697 (O_2697,N_21891,N_23376);
or UO_2698 (O_2698,N_23591,N_23319);
nand UO_2699 (O_2699,N_24628,N_23355);
or UO_2700 (O_2700,N_24885,N_22198);
nand UO_2701 (O_2701,N_24831,N_24031);
or UO_2702 (O_2702,N_21997,N_23067);
nand UO_2703 (O_2703,N_22278,N_23107);
or UO_2704 (O_2704,N_22596,N_22463);
and UO_2705 (O_2705,N_24946,N_22902);
nand UO_2706 (O_2706,N_22648,N_24553);
and UO_2707 (O_2707,N_24358,N_22169);
and UO_2708 (O_2708,N_24462,N_24289);
nor UO_2709 (O_2709,N_22553,N_23521);
or UO_2710 (O_2710,N_22760,N_23906);
or UO_2711 (O_2711,N_24189,N_22939);
or UO_2712 (O_2712,N_24688,N_24551);
nor UO_2713 (O_2713,N_23535,N_23393);
or UO_2714 (O_2714,N_24426,N_22170);
or UO_2715 (O_2715,N_22321,N_24748);
nor UO_2716 (O_2716,N_24219,N_22477);
and UO_2717 (O_2717,N_23400,N_24472);
xor UO_2718 (O_2718,N_23628,N_24431);
nor UO_2719 (O_2719,N_23010,N_24862);
nand UO_2720 (O_2720,N_24241,N_22428);
xor UO_2721 (O_2721,N_23674,N_24987);
or UO_2722 (O_2722,N_23522,N_22887);
and UO_2723 (O_2723,N_23161,N_23393);
nand UO_2724 (O_2724,N_24623,N_24027);
and UO_2725 (O_2725,N_24833,N_24715);
nand UO_2726 (O_2726,N_22784,N_22524);
and UO_2727 (O_2727,N_23539,N_24938);
nor UO_2728 (O_2728,N_23914,N_23483);
xnor UO_2729 (O_2729,N_24124,N_24449);
or UO_2730 (O_2730,N_21897,N_23110);
and UO_2731 (O_2731,N_22060,N_23763);
and UO_2732 (O_2732,N_22139,N_21875);
nand UO_2733 (O_2733,N_22509,N_22187);
nor UO_2734 (O_2734,N_21940,N_24767);
or UO_2735 (O_2735,N_24158,N_24314);
nor UO_2736 (O_2736,N_22609,N_24485);
or UO_2737 (O_2737,N_22879,N_24697);
nand UO_2738 (O_2738,N_23686,N_23568);
or UO_2739 (O_2739,N_24252,N_22986);
nand UO_2740 (O_2740,N_21983,N_23453);
xor UO_2741 (O_2741,N_22468,N_23850);
and UO_2742 (O_2742,N_22405,N_24066);
nand UO_2743 (O_2743,N_24790,N_23472);
xor UO_2744 (O_2744,N_22580,N_23302);
and UO_2745 (O_2745,N_22099,N_22629);
nor UO_2746 (O_2746,N_22810,N_22616);
nand UO_2747 (O_2747,N_24490,N_23260);
and UO_2748 (O_2748,N_24223,N_22894);
and UO_2749 (O_2749,N_24357,N_22234);
or UO_2750 (O_2750,N_22300,N_22414);
nand UO_2751 (O_2751,N_23407,N_23746);
xnor UO_2752 (O_2752,N_23784,N_22420);
nand UO_2753 (O_2753,N_21880,N_22857);
or UO_2754 (O_2754,N_24615,N_21913);
and UO_2755 (O_2755,N_22284,N_22841);
nor UO_2756 (O_2756,N_23852,N_24441);
or UO_2757 (O_2757,N_23964,N_22483);
xor UO_2758 (O_2758,N_21913,N_23409);
xor UO_2759 (O_2759,N_23723,N_24642);
or UO_2760 (O_2760,N_24456,N_23302);
nand UO_2761 (O_2761,N_22286,N_23745);
or UO_2762 (O_2762,N_23690,N_24247);
or UO_2763 (O_2763,N_24605,N_22871);
nand UO_2764 (O_2764,N_22486,N_22685);
xnor UO_2765 (O_2765,N_24149,N_23065);
and UO_2766 (O_2766,N_24688,N_23837);
or UO_2767 (O_2767,N_23018,N_23338);
nand UO_2768 (O_2768,N_22962,N_24911);
nand UO_2769 (O_2769,N_22576,N_23726);
xor UO_2770 (O_2770,N_24332,N_22693);
nand UO_2771 (O_2771,N_24082,N_23554);
xnor UO_2772 (O_2772,N_24843,N_24730);
or UO_2773 (O_2773,N_23815,N_23954);
nand UO_2774 (O_2774,N_22018,N_22246);
xnor UO_2775 (O_2775,N_22756,N_22463);
xor UO_2776 (O_2776,N_24019,N_23076);
or UO_2777 (O_2777,N_22463,N_23167);
and UO_2778 (O_2778,N_23906,N_22162);
xnor UO_2779 (O_2779,N_23329,N_24385);
nand UO_2780 (O_2780,N_24563,N_23444);
or UO_2781 (O_2781,N_23774,N_24497);
nor UO_2782 (O_2782,N_22135,N_23839);
or UO_2783 (O_2783,N_24002,N_24328);
nand UO_2784 (O_2784,N_22173,N_24159);
and UO_2785 (O_2785,N_22450,N_24277);
nand UO_2786 (O_2786,N_24465,N_23367);
xnor UO_2787 (O_2787,N_22486,N_22956);
or UO_2788 (O_2788,N_22241,N_24921);
or UO_2789 (O_2789,N_23420,N_22427);
or UO_2790 (O_2790,N_22929,N_23612);
xnor UO_2791 (O_2791,N_21880,N_24377);
xnor UO_2792 (O_2792,N_23582,N_24549);
and UO_2793 (O_2793,N_22627,N_22784);
nor UO_2794 (O_2794,N_22072,N_22612);
nand UO_2795 (O_2795,N_24842,N_24927);
xnor UO_2796 (O_2796,N_22613,N_23779);
xor UO_2797 (O_2797,N_22291,N_23092);
nand UO_2798 (O_2798,N_24641,N_23272);
or UO_2799 (O_2799,N_22247,N_24591);
nand UO_2800 (O_2800,N_24010,N_22217);
nand UO_2801 (O_2801,N_22296,N_24987);
xor UO_2802 (O_2802,N_22628,N_24675);
nand UO_2803 (O_2803,N_24229,N_24473);
and UO_2804 (O_2804,N_22124,N_24084);
or UO_2805 (O_2805,N_23670,N_24750);
or UO_2806 (O_2806,N_24402,N_24370);
and UO_2807 (O_2807,N_22983,N_24245);
nand UO_2808 (O_2808,N_24633,N_22395);
nand UO_2809 (O_2809,N_23782,N_23289);
and UO_2810 (O_2810,N_23837,N_24764);
and UO_2811 (O_2811,N_23344,N_22474);
and UO_2812 (O_2812,N_23459,N_23867);
and UO_2813 (O_2813,N_24937,N_23235);
and UO_2814 (O_2814,N_24916,N_22356);
and UO_2815 (O_2815,N_24703,N_23572);
and UO_2816 (O_2816,N_24830,N_22694);
and UO_2817 (O_2817,N_23693,N_22597);
and UO_2818 (O_2818,N_22545,N_22828);
nand UO_2819 (O_2819,N_24639,N_24457);
or UO_2820 (O_2820,N_24050,N_24129);
nand UO_2821 (O_2821,N_24196,N_22334);
nand UO_2822 (O_2822,N_24514,N_21907);
or UO_2823 (O_2823,N_24004,N_23117);
nand UO_2824 (O_2824,N_22483,N_24587);
or UO_2825 (O_2825,N_24699,N_23560);
and UO_2826 (O_2826,N_23123,N_23274);
or UO_2827 (O_2827,N_22067,N_24855);
nand UO_2828 (O_2828,N_24452,N_23574);
and UO_2829 (O_2829,N_24172,N_22548);
xnor UO_2830 (O_2830,N_24427,N_23551);
xor UO_2831 (O_2831,N_22078,N_23011);
and UO_2832 (O_2832,N_23908,N_22254);
and UO_2833 (O_2833,N_23413,N_22325);
or UO_2834 (O_2834,N_23184,N_24875);
nand UO_2835 (O_2835,N_23344,N_24629);
xnor UO_2836 (O_2836,N_24892,N_23376);
nand UO_2837 (O_2837,N_24147,N_22140);
xnor UO_2838 (O_2838,N_24726,N_24979);
or UO_2839 (O_2839,N_23651,N_24025);
or UO_2840 (O_2840,N_23367,N_24785);
or UO_2841 (O_2841,N_23762,N_22921);
xnor UO_2842 (O_2842,N_24447,N_23330);
and UO_2843 (O_2843,N_22027,N_23431);
xor UO_2844 (O_2844,N_24496,N_24744);
or UO_2845 (O_2845,N_23941,N_23431);
nand UO_2846 (O_2846,N_24773,N_24013);
nand UO_2847 (O_2847,N_23929,N_24275);
or UO_2848 (O_2848,N_22484,N_23577);
nor UO_2849 (O_2849,N_22368,N_22707);
nor UO_2850 (O_2850,N_24238,N_22919);
nor UO_2851 (O_2851,N_24274,N_22349);
nand UO_2852 (O_2852,N_22095,N_24417);
and UO_2853 (O_2853,N_23380,N_24514);
or UO_2854 (O_2854,N_22864,N_22031);
or UO_2855 (O_2855,N_22795,N_22263);
xnor UO_2856 (O_2856,N_24196,N_23455);
and UO_2857 (O_2857,N_22325,N_23514);
or UO_2858 (O_2858,N_23701,N_22441);
and UO_2859 (O_2859,N_24008,N_23651);
nor UO_2860 (O_2860,N_23813,N_22898);
nor UO_2861 (O_2861,N_24248,N_22433);
and UO_2862 (O_2862,N_22877,N_23862);
nor UO_2863 (O_2863,N_24703,N_23264);
xor UO_2864 (O_2864,N_22643,N_24171);
or UO_2865 (O_2865,N_24591,N_24951);
nor UO_2866 (O_2866,N_23817,N_24669);
nand UO_2867 (O_2867,N_23178,N_24674);
nand UO_2868 (O_2868,N_23489,N_23255);
nor UO_2869 (O_2869,N_23417,N_23558);
and UO_2870 (O_2870,N_22113,N_23607);
xnor UO_2871 (O_2871,N_23786,N_23129);
and UO_2872 (O_2872,N_23389,N_22727);
xnor UO_2873 (O_2873,N_23350,N_23335);
or UO_2874 (O_2874,N_22278,N_23681);
nor UO_2875 (O_2875,N_24991,N_23092);
nor UO_2876 (O_2876,N_22210,N_22096);
or UO_2877 (O_2877,N_22241,N_23232);
nand UO_2878 (O_2878,N_23176,N_22218);
or UO_2879 (O_2879,N_22867,N_22330);
nand UO_2880 (O_2880,N_22337,N_24357);
and UO_2881 (O_2881,N_23073,N_24895);
nand UO_2882 (O_2882,N_23549,N_22866);
xnor UO_2883 (O_2883,N_22673,N_23548);
nor UO_2884 (O_2884,N_24293,N_23563);
xnor UO_2885 (O_2885,N_23405,N_23370);
and UO_2886 (O_2886,N_22046,N_22585);
nor UO_2887 (O_2887,N_24899,N_22390);
nor UO_2888 (O_2888,N_24863,N_22499);
and UO_2889 (O_2889,N_22381,N_24332);
or UO_2890 (O_2890,N_23240,N_22890);
and UO_2891 (O_2891,N_23594,N_22430);
or UO_2892 (O_2892,N_23501,N_24036);
xor UO_2893 (O_2893,N_24956,N_22849);
nor UO_2894 (O_2894,N_24543,N_24937);
or UO_2895 (O_2895,N_24743,N_24037);
and UO_2896 (O_2896,N_24001,N_24293);
nand UO_2897 (O_2897,N_22781,N_22275);
nand UO_2898 (O_2898,N_23835,N_22365);
xor UO_2899 (O_2899,N_23235,N_21973);
nand UO_2900 (O_2900,N_22516,N_21985);
or UO_2901 (O_2901,N_22488,N_22167);
nor UO_2902 (O_2902,N_22621,N_23079);
nand UO_2903 (O_2903,N_22585,N_23103);
and UO_2904 (O_2904,N_24932,N_22045);
and UO_2905 (O_2905,N_22755,N_24888);
nand UO_2906 (O_2906,N_23531,N_23305);
nor UO_2907 (O_2907,N_24437,N_22911);
nand UO_2908 (O_2908,N_22930,N_23782);
nand UO_2909 (O_2909,N_22325,N_23567);
or UO_2910 (O_2910,N_22967,N_24055);
and UO_2911 (O_2911,N_23207,N_23231);
nor UO_2912 (O_2912,N_22569,N_23412);
xnor UO_2913 (O_2913,N_23475,N_24248);
nand UO_2914 (O_2914,N_22974,N_24590);
xnor UO_2915 (O_2915,N_23359,N_22093);
and UO_2916 (O_2916,N_22440,N_23751);
nand UO_2917 (O_2917,N_23194,N_23097);
nand UO_2918 (O_2918,N_22683,N_23925);
nor UO_2919 (O_2919,N_24334,N_23557);
and UO_2920 (O_2920,N_23924,N_24892);
or UO_2921 (O_2921,N_23674,N_22919);
xor UO_2922 (O_2922,N_22333,N_24896);
or UO_2923 (O_2923,N_24558,N_22825);
nor UO_2924 (O_2924,N_23836,N_22142);
xor UO_2925 (O_2925,N_23795,N_21898);
or UO_2926 (O_2926,N_24659,N_24655);
xnor UO_2927 (O_2927,N_23884,N_22598);
nor UO_2928 (O_2928,N_22901,N_22137);
nor UO_2929 (O_2929,N_22360,N_23043);
and UO_2930 (O_2930,N_23503,N_24078);
and UO_2931 (O_2931,N_23008,N_22108);
nand UO_2932 (O_2932,N_23061,N_24488);
nand UO_2933 (O_2933,N_23555,N_22892);
and UO_2934 (O_2934,N_24134,N_24613);
nor UO_2935 (O_2935,N_22592,N_24534);
nand UO_2936 (O_2936,N_23994,N_23999);
xor UO_2937 (O_2937,N_24824,N_24746);
xor UO_2938 (O_2938,N_23564,N_24665);
and UO_2939 (O_2939,N_23927,N_23201);
and UO_2940 (O_2940,N_23619,N_23302);
or UO_2941 (O_2941,N_24518,N_22913);
nand UO_2942 (O_2942,N_24088,N_23496);
or UO_2943 (O_2943,N_22446,N_22967);
nor UO_2944 (O_2944,N_23880,N_23441);
nor UO_2945 (O_2945,N_24928,N_22307);
or UO_2946 (O_2946,N_23990,N_22593);
nor UO_2947 (O_2947,N_24533,N_23413);
or UO_2948 (O_2948,N_22315,N_23075);
or UO_2949 (O_2949,N_23825,N_22498);
and UO_2950 (O_2950,N_22181,N_22866);
and UO_2951 (O_2951,N_23574,N_23114);
nor UO_2952 (O_2952,N_22582,N_23896);
nand UO_2953 (O_2953,N_24055,N_24330);
or UO_2954 (O_2954,N_22650,N_23381);
nand UO_2955 (O_2955,N_21965,N_22330);
nand UO_2956 (O_2956,N_23063,N_23623);
nand UO_2957 (O_2957,N_22655,N_23158);
nand UO_2958 (O_2958,N_23878,N_24958);
nand UO_2959 (O_2959,N_23317,N_24498);
and UO_2960 (O_2960,N_24065,N_22963);
or UO_2961 (O_2961,N_23385,N_22108);
or UO_2962 (O_2962,N_24379,N_24762);
and UO_2963 (O_2963,N_23157,N_24000);
xnor UO_2964 (O_2964,N_24599,N_23784);
nor UO_2965 (O_2965,N_22412,N_24562);
and UO_2966 (O_2966,N_23254,N_22188);
nand UO_2967 (O_2967,N_22913,N_24042);
nor UO_2968 (O_2968,N_23301,N_22951);
nor UO_2969 (O_2969,N_22543,N_23827);
and UO_2970 (O_2970,N_24058,N_24881);
and UO_2971 (O_2971,N_23531,N_22717);
and UO_2972 (O_2972,N_23311,N_24347);
nand UO_2973 (O_2973,N_22675,N_24082);
nor UO_2974 (O_2974,N_23602,N_22992);
xnor UO_2975 (O_2975,N_24495,N_24702);
nand UO_2976 (O_2976,N_22504,N_21974);
or UO_2977 (O_2977,N_24471,N_22627);
xor UO_2978 (O_2978,N_23661,N_22302);
or UO_2979 (O_2979,N_24222,N_24132);
nand UO_2980 (O_2980,N_22934,N_22543);
or UO_2981 (O_2981,N_24497,N_23546);
nor UO_2982 (O_2982,N_22190,N_23300);
xnor UO_2983 (O_2983,N_24615,N_23858);
nor UO_2984 (O_2984,N_21998,N_24918);
or UO_2985 (O_2985,N_22878,N_24012);
and UO_2986 (O_2986,N_23396,N_23783);
or UO_2987 (O_2987,N_23847,N_24228);
nor UO_2988 (O_2988,N_23439,N_23733);
or UO_2989 (O_2989,N_23078,N_22315);
xnor UO_2990 (O_2990,N_24679,N_24531);
nand UO_2991 (O_2991,N_23147,N_23278);
nor UO_2992 (O_2992,N_24790,N_23499);
nor UO_2993 (O_2993,N_24768,N_21944);
or UO_2994 (O_2994,N_22960,N_24694);
or UO_2995 (O_2995,N_24250,N_22444);
and UO_2996 (O_2996,N_23688,N_21928);
and UO_2997 (O_2997,N_24233,N_24102);
and UO_2998 (O_2998,N_24666,N_23770);
nor UO_2999 (O_2999,N_22983,N_23738);
endmodule