module basic_3000_30000_3500_3_levels_1xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20003,N_20004,N_20005,N_20006,N_20009,N_20011,N_20013,N_20014,N_20015,N_20016,N_20017,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20027,N_20028,N_20030,N_20034,N_20035,N_20037,N_20039,N_20040,N_20041,N_20043,N_20045,N_20046,N_20047,N_20048,N_20050,N_20051,N_20052,N_20054,N_20056,N_20057,N_20059,N_20060,N_20062,N_20063,N_20065,N_20066,N_20067,N_20070,N_20071,N_20072,N_20074,N_20075,N_20076,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20091,N_20092,N_20093,N_20095,N_20098,N_20099,N_20100,N_20101,N_20102,N_20104,N_20105,N_20106,N_20107,N_20108,N_20110,N_20111,N_20113,N_20114,N_20115,N_20116,N_20118,N_20119,N_20120,N_20121,N_20123,N_20124,N_20125,N_20127,N_20129,N_20130,N_20131,N_20133,N_20134,N_20136,N_20137,N_20138,N_20140,N_20141,N_20143,N_20144,N_20146,N_20147,N_20148,N_20149,N_20150,N_20152,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20166,N_20167,N_20168,N_20171,N_20172,N_20175,N_20176,N_20177,N_20178,N_20180,N_20181,N_20182,N_20184,N_20185,N_20189,N_20190,N_20191,N_20193,N_20194,N_20197,N_20202,N_20204,N_20205,N_20206,N_20208,N_20210,N_20211,N_20212,N_20214,N_20215,N_20216,N_20218,N_20220,N_20222,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20233,N_20234,N_20235,N_20237,N_20239,N_20242,N_20244,N_20246,N_20248,N_20249,N_20252,N_20253,N_20255,N_20256,N_20259,N_20260,N_20261,N_20263,N_20265,N_20266,N_20267,N_20268,N_20269,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20298,N_20299,N_20300,N_20303,N_20304,N_20305,N_20306,N_20307,N_20310,N_20311,N_20312,N_20313,N_20314,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20323,N_20324,N_20329,N_20330,N_20333,N_20336,N_20337,N_20339,N_20340,N_20342,N_20345,N_20346,N_20348,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20363,N_20364,N_20365,N_20366,N_20367,N_20369,N_20370,N_20371,N_20375,N_20377,N_20378,N_20379,N_20382,N_20383,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20392,N_20393,N_20395,N_20396,N_20397,N_20399,N_20400,N_20401,N_20402,N_20403,N_20405,N_20406,N_20407,N_20408,N_20409,N_20412,N_20413,N_20415,N_20416,N_20419,N_20420,N_20421,N_20422,N_20423,N_20425,N_20427,N_20430,N_20431,N_20432,N_20433,N_20435,N_20437,N_20438,N_20440,N_20441,N_20442,N_20443,N_20444,N_20446,N_20447,N_20448,N_20449,N_20453,N_20454,N_20455,N_20456,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20469,N_20470,N_20472,N_20473,N_20474,N_20476,N_20477,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20492,N_20493,N_20494,N_20497,N_20498,N_20499,N_20500,N_20502,N_20503,N_20505,N_20506,N_20507,N_20510,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20531,N_20532,N_20533,N_20534,N_20538,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20548,N_20549,N_20550,N_20552,N_20553,N_20554,N_20555,N_20557,N_20558,N_20559,N_20560,N_20562,N_20563,N_20565,N_20566,N_20568,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20577,N_20579,N_20585,N_20586,N_20587,N_20588,N_20591,N_20593,N_20594,N_20595,N_20596,N_20597,N_20599,N_20600,N_20602,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20611,N_20613,N_20614,N_20615,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20627,N_20628,N_20629,N_20631,N_20632,N_20633,N_20635,N_20636,N_20637,N_20638,N_20640,N_20641,N_20642,N_20643,N_20646,N_20648,N_20649,N_20650,N_20651,N_20652,N_20654,N_20655,N_20657,N_20659,N_20660,N_20661,N_20663,N_20666,N_20667,N_20668,N_20669,N_20670,N_20672,N_20673,N_20676,N_20679,N_20682,N_20683,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20701,N_20702,N_20703,N_20704,N_20706,N_20707,N_20709,N_20711,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20730,N_20731,N_20732,N_20733,N_20737,N_20738,N_20741,N_20744,N_20745,N_20746,N_20747,N_20752,N_20753,N_20754,N_20757,N_20758,N_20759,N_20761,N_20763,N_20764,N_20765,N_20766,N_20767,N_20769,N_20770,N_20771,N_20772,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20781,N_20782,N_20783,N_20784,N_20785,N_20788,N_20789,N_20792,N_20793,N_20794,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20803,N_20804,N_20805,N_20807,N_20809,N_20810,N_20811,N_20812,N_20813,N_20816,N_20817,N_20818,N_20819,N_20821,N_20823,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20842,N_20843,N_20844,N_20846,N_20847,N_20848,N_20849,N_20852,N_20854,N_20855,N_20856,N_20858,N_20859,N_20860,N_20863,N_20864,N_20866,N_20867,N_20868,N_20869,N_20871,N_20872,N_20873,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20886,N_20888,N_20889,N_20891,N_20893,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20905,N_20907,N_20908,N_20909,N_20912,N_20914,N_20915,N_20917,N_20918,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20940,N_20941,N_20942,N_20944,N_20947,N_20949,N_20950,N_20951,N_20952,N_20954,N_20957,N_20958,N_20959,N_20960,N_20963,N_20964,N_20965,N_20967,N_20968,N_20969,N_20975,N_20976,N_20977,N_20979,N_20981,N_20982,N_20983,N_20984,N_20985,N_20987,N_20989,N_20991,N_20992,N_20994,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21015,N_21017,N_21018,N_21021,N_21023,N_21025,N_21026,N_21027,N_21028,N_21029,N_21031,N_21032,N_21034,N_21035,N_21036,N_21037,N_21039,N_21040,N_21042,N_21043,N_21044,N_21045,N_21046,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21057,N_21060,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21086,N_21087,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21098,N_21100,N_21101,N_21103,N_21105,N_21107,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21126,N_21127,N_21128,N_21129,N_21130,N_21132,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21142,N_21144,N_21145,N_21147,N_21148,N_21151,N_21152,N_21153,N_21154,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21173,N_21174,N_21175,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21193,N_21194,N_21195,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21207,N_21209,N_21213,N_21214,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21226,N_21227,N_21229,N_21230,N_21232,N_21234,N_21235,N_21236,N_21240,N_21241,N_21242,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21251,N_21252,N_21253,N_21254,N_21255,N_21257,N_21258,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21269,N_21270,N_21271,N_21272,N_21274,N_21276,N_21277,N_21278,N_21281,N_21283,N_21284,N_21285,N_21286,N_21287,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21302,N_21303,N_21304,N_21305,N_21307,N_21311,N_21313,N_21315,N_21316,N_21317,N_21318,N_21320,N_21321,N_21322,N_21324,N_21326,N_21327,N_21328,N_21329,N_21330,N_21332,N_21333,N_21334,N_21337,N_21338,N_21341,N_21342,N_21344,N_21345,N_21346,N_21348,N_21349,N_21350,N_21351,N_21353,N_21354,N_21355,N_21356,N_21358,N_21359,N_21360,N_21361,N_21363,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21380,N_21381,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21391,N_21392,N_21393,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21403,N_21405,N_21406,N_21407,N_21410,N_21412,N_21413,N_21415,N_21416,N_21417,N_21418,N_21421,N_21422,N_21423,N_21424,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21480,N_21481,N_21483,N_21485,N_21486,N_21487,N_21488,N_21490,N_21495,N_21496,N_21497,N_21498,N_21501,N_21504,N_21505,N_21506,N_21507,N_21508,N_21510,N_21511,N_21513,N_21515,N_21516,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21526,N_21528,N_21530,N_21533,N_21538,N_21541,N_21543,N_21546,N_21547,N_21548,N_21549,N_21551,N_21552,N_21553,N_21555,N_21559,N_21560,N_21562,N_21563,N_21564,N_21565,N_21566,N_21568,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21591,N_21592,N_21594,N_21595,N_21596,N_21597,N_21599,N_21600,N_21601,N_21602,N_21603,N_21605,N_21606,N_21607,N_21610,N_21611,N_21612,N_21614,N_21615,N_21618,N_21620,N_21622,N_21624,N_21626,N_21628,N_21630,N_21631,N_21633,N_21634,N_21636,N_21638,N_21639,N_21641,N_21642,N_21644,N_21645,N_21647,N_21649,N_21652,N_21654,N_21656,N_21657,N_21660,N_21664,N_21665,N_21666,N_21667,N_21668,N_21670,N_21671,N_21674,N_21675,N_21676,N_21678,N_21679,N_21680,N_21681,N_21683,N_21684,N_21685,N_21687,N_21688,N_21690,N_21692,N_21694,N_21695,N_21696,N_21697,N_21699,N_21701,N_21702,N_21703,N_21711,N_21712,N_21713,N_21714,N_21717,N_21719,N_21720,N_21721,N_21722,N_21725,N_21726,N_21728,N_21729,N_21732,N_21733,N_21734,N_21735,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21758,N_21759,N_21761,N_21762,N_21763,N_21764,N_21765,N_21767,N_21770,N_21771,N_21773,N_21775,N_21776,N_21782,N_21783,N_21784,N_21785,N_21786,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21801,N_21802,N_21803,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21819,N_21820,N_21822,N_21824,N_21827,N_21831,N_21832,N_21835,N_21836,N_21838,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21848,N_21849,N_21851,N_21852,N_21853,N_21854,N_21856,N_21857,N_21858,N_21859,N_21861,N_21864,N_21865,N_21866,N_21867,N_21868,N_21871,N_21873,N_21874,N_21876,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21888,N_21889,N_21890,N_21891,N_21894,N_21897,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21908,N_21909,N_21910,N_21911,N_21912,N_21914,N_21915,N_21916,N_21919,N_21920,N_21921,N_21923,N_21924,N_21926,N_21929,N_21933,N_21934,N_21936,N_21938,N_21941,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21976,N_21977,N_21978,N_21979,N_21980,N_21983,N_21986,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22007,N_22009,N_22010,N_22011,N_22013,N_22014,N_22016,N_22018,N_22020,N_22021,N_22024,N_22026,N_22027,N_22028,N_22029,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22042,N_22044,N_22046,N_22047,N_22049,N_22051,N_22052,N_22053,N_22054,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22065,N_22067,N_22068,N_22069,N_22070,N_22072,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22106,N_22107,N_22110,N_22112,N_22114,N_22119,N_22120,N_22121,N_22123,N_22124,N_22125,N_22126,N_22128,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22140,N_22141,N_22142,N_22143,N_22145,N_22146,N_22147,N_22148,N_22150,N_22152,N_22153,N_22155,N_22157,N_22158,N_22159,N_22160,N_22161,N_22163,N_22164,N_22165,N_22166,N_22169,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22183,N_22185,N_22186,N_22188,N_22189,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22203,N_22205,N_22206,N_22207,N_22209,N_22211,N_22212,N_22213,N_22215,N_22216,N_22217,N_22219,N_22220,N_22221,N_22222,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22235,N_22236,N_22239,N_22242,N_22243,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22254,N_22255,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22268,N_22269,N_22271,N_22272,N_22273,N_22274,N_22275,N_22278,N_22280,N_22281,N_22282,N_22283,N_22285,N_22286,N_22288,N_22290,N_22292,N_22294,N_22295,N_22296,N_22298,N_22299,N_22300,N_22301,N_22303,N_22305,N_22306,N_22307,N_22308,N_22309,N_22311,N_22312,N_22315,N_22319,N_22320,N_22321,N_22323,N_22324,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22336,N_22341,N_22342,N_22343,N_22345,N_22346,N_22347,N_22348,N_22350,N_22351,N_22352,N_22353,N_22354,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22366,N_22367,N_22370,N_22371,N_22373,N_22374,N_22375,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22408,N_22409,N_22411,N_22415,N_22417,N_22418,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22428,N_22430,N_22431,N_22432,N_22435,N_22436,N_22437,N_22438,N_22440,N_22443,N_22444,N_22445,N_22446,N_22449,N_22450,N_22451,N_22453,N_22455,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22473,N_22474,N_22475,N_22477,N_22478,N_22479,N_22480,N_22482,N_22483,N_22485,N_22487,N_22489,N_22490,N_22491,N_22492,N_22493,N_22495,N_22496,N_22498,N_22499,N_22500,N_22501,N_22503,N_22505,N_22507,N_22508,N_22509,N_22511,N_22512,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22523,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22534,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22544,N_22545,N_22546,N_22547,N_22549,N_22550,N_22551,N_22553,N_22555,N_22556,N_22558,N_22559,N_22562,N_22563,N_22564,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22576,N_22577,N_22578,N_22579,N_22580,N_22582,N_22584,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22594,N_22595,N_22596,N_22598,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22609,N_22610,N_22611,N_22614,N_22615,N_22616,N_22619,N_22621,N_22623,N_22624,N_22625,N_22628,N_22630,N_22631,N_22634,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22644,N_22645,N_22646,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22655,N_22656,N_22657,N_22659,N_22660,N_22661,N_22663,N_22664,N_22665,N_22667,N_22670,N_22671,N_22672,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22684,N_22685,N_22686,N_22687,N_22688,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22705,N_22708,N_22709,N_22710,N_22712,N_22714,N_22715,N_22716,N_22717,N_22719,N_22721,N_22722,N_22723,N_22724,N_22726,N_22727,N_22728,N_22730,N_22733,N_22735,N_22736,N_22737,N_22738,N_22739,N_22741,N_22742,N_22743,N_22744,N_22746,N_22747,N_22748,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22759,N_22761,N_22763,N_22764,N_22766,N_22767,N_22768,N_22769,N_22770,N_22773,N_22774,N_22775,N_22776,N_22779,N_22780,N_22781,N_22782,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22793,N_22795,N_22796,N_22797,N_22798,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22816,N_22817,N_22818,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22832,N_22836,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22849,N_22850,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22880,N_22883,N_22884,N_22885,N_22886,N_22887,N_22890,N_22891,N_22893,N_22894,N_22895,N_22896,N_22898,N_22901,N_22902,N_22903,N_22904,N_22906,N_22907,N_22908,N_22910,N_22911,N_22912,N_22913,N_22914,N_22916,N_22917,N_22918,N_22919,N_22922,N_22923,N_22925,N_22926,N_22927,N_22928,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22938,N_22940,N_22941,N_22943,N_22944,N_22945,N_22947,N_22948,N_22949,N_22950,N_22951,N_22953,N_22954,N_22955,N_22957,N_22958,N_22959,N_22960,N_22962,N_22963,N_22965,N_22966,N_22968,N_22970,N_22975,N_22976,N_22979,N_22980,N_22981,N_22982,N_22983,N_22985,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22997,N_22998,N_23000,N_23001,N_23003,N_23006,N_23007,N_23008,N_23010,N_23011,N_23012,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23021,N_23022,N_23023,N_23025,N_23027,N_23028,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23038,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23055,N_23056,N_23057,N_23058,N_23059,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23068,N_23069,N_23071,N_23072,N_23074,N_23075,N_23076,N_23077,N_23078,N_23082,N_23083,N_23085,N_23087,N_23088,N_23090,N_23091,N_23096,N_23099,N_23100,N_23101,N_23103,N_23104,N_23107,N_23108,N_23109,N_23111,N_23112,N_23113,N_23115,N_23117,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23126,N_23128,N_23129,N_23130,N_23131,N_23134,N_23136,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23160,N_23161,N_23164,N_23165,N_23167,N_23168,N_23172,N_23174,N_23176,N_23178,N_23179,N_23180,N_23181,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23192,N_23193,N_23195,N_23196,N_23198,N_23199,N_23201,N_23202,N_23204,N_23205,N_23207,N_23208,N_23210,N_23212,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23223,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23236,N_23237,N_23238,N_23239,N_23242,N_23243,N_23247,N_23249,N_23250,N_23251,N_23252,N_23254,N_23255,N_23256,N_23257,N_23260,N_23261,N_23262,N_23264,N_23265,N_23266,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23280,N_23281,N_23282,N_23284,N_23285,N_23286,N_23288,N_23289,N_23291,N_23292,N_23294,N_23296,N_23297,N_23300,N_23301,N_23303,N_23304,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23319,N_23320,N_23321,N_23323,N_23324,N_23325,N_23326,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23359,N_23361,N_23362,N_23363,N_23364,N_23365,N_23367,N_23370,N_23371,N_23372,N_23373,N_23378,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23389,N_23390,N_23391,N_23392,N_23393,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23404,N_23405,N_23407,N_23408,N_23409,N_23410,N_23412,N_23413,N_23415,N_23416,N_23417,N_23418,N_23419,N_23421,N_23423,N_23424,N_23426,N_23427,N_23428,N_23429,N_23431,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23443,N_23445,N_23446,N_23448,N_23451,N_23454,N_23456,N_23457,N_23459,N_23460,N_23461,N_23462,N_23463,N_23465,N_23466,N_23467,N_23469,N_23470,N_23471,N_23473,N_23475,N_23477,N_23478,N_23480,N_23481,N_23482,N_23483,N_23488,N_23490,N_23491,N_23492,N_23493,N_23495,N_23496,N_23497,N_23499,N_23501,N_23504,N_23505,N_23506,N_23508,N_23509,N_23511,N_23512,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23538,N_23539,N_23540,N_23541,N_23542,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23553,N_23554,N_23557,N_23558,N_23559,N_23561,N_23562,N_23563,N_23564,N_23566,N_23567,N_23571,N_23572,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23592,N_23594,N_23595,N_23596,N_23598,N_23599,N_23600,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23626,N_23627,N_23628,N_23629,N_23630,N_23632,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23642,N_23645,N_23646,N_23648,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23670,N_23671,N_23672,N_23673,N_23674,N_23676,N_23678,N_23680,N_23682,N_23684,N_23685,N_23688,N_23689,N_23691,N_23694,N_23695,N_23696,N_23697,N_23699,N_23700,N_23701,N_23702,N_23706,N_23707,N_23708,N_23710,N_23711,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23720,N_23721,N_23722,N_23724,N_23725,N_23728,N_23736,N_23738,N_23740,N_23741,N_23742,N_23744,N_23746,N_23747,N_23748,N_23750,N_23751,N_23754,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23764,N_23765,N_23766,N_23768,N_23769,N_23770,N_23774,N_23776,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23787,N_23788,N_23790,N_23792,N_23793,N_23794,N_23795,N_23798,N_23799,N_23800,N_23801,N_23803,N_23805,N_23806,N_23807,N_23808,N_23810,N_23811,N_23814,N_23815,N_23818,N_23819,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23829,N_23830,N_23831,N_23833,N_23834,N_23835,N_23836,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23846,N_23847,N_23848,N_23849,N_23850,N_23852,N_23856,N_23857,N_23859,N_23861,N_23864,N_23865,N_23866,N_23867,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23877,N_23878,N_23879,N_23880,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23898,N_23899,N_23900,N_23903,N_23905,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23927,N_23935,N_23936,N_23938,N_23940,N_23941,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23953,N_23954,N_23955,N_23956,N_23958,N_23959,N_23960,N_23962,N_23965,N_23967,N_23970,N_23971,N_23972,N_23973,N_23974,N_23976,N_23977,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23990,N_23992,N_23994,N_23995,N_23996,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24008,N_24009,N_24010,N_24011,N_24013,N_24014,N_24015,N_24016,N_24017,N_24020,N_24022,N_24023,N_24025,N_24028,N_24029,N_24032,N_24034,N_24036,N_24037,N_24039,N_24040,N_24042,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24052,N_24053,N_24054,N_24055,N_24057,N_24060,N_24061,N_24062,N_24063,N_24065,N_24068,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24082,N_24083,N_24084,N_24085,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24098,N_24102,N_24105,N_24107,N_24109,N_24110,N_24112,N_24115,N_24116,N_24117,N_24121,N_24122,N_24125,N_24126,N_24129,N_24130,N_24131,N_24135,N_24136,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24148,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24167,N_24169,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24178,N_24179,N_24182,N_24183,N_24186,N_24188,N_24189,N_24190,N_24191,N_24192,N_24194,N_24201,N_24202,N_24203,N_24205,N_24206,N_24209,N_24212,N_24214,N_24215,N_24219,N_24221,N_24224,N_24225,N_24226,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24240,N_24241,N_24243,N_24244,N_24247,N_24248,N_24249,N_24250,N_24253,N_24254,N_24256,N_24257,N_24258,N_24260,N_24261,N_24263,N_24264,N_24265,N_24267,N_24268,N_24269,N_24270,N_24272,N_24273,N_24275,N_24276,N_24278,N_24279,N_24281,N_24282,N_24283,N_24284,N_24286,N_24288,N_24289,N_24290,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24301,N_24305,N_24307,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24320,N_24321,N_24322,N_24325,N_24327,N_24328,N_24329,N_24330,N_24331,N_24333,N_24334,N_24338,N_24340,N_24341,N_24342,N_24343,N_24344,N_24347,N_24348,N_24349,N_24350,N_24352,N_24354,N_24355,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24364,N_24365,N_24366,N_24367,N_24370,N_24372,N_24373,N_24374,N_24375,N_24377,N_24378,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24393,N_24394,N_24395,N_24397,N_24399,N_24402,N_24403,N_24404,N_24405,N_24408,N_24410,N_24411,N_24412,N_24413,N_24415,N_24416,N_24417,N_24423,N_24425,N_24426,N_24428,N_24429,N_24430,N_24431,N_24433,N_24434,N_24437,N_24439,N_24440,N_24441,N_24442,N_24443,N_24445,N_24446,N_24447,N_24448,N_24450,N_24451,N_24452,N_24454,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24473,N_24474,N_24475,N_24476,N_24478,N_24479,N_24480,N_24481,N_24482,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24496,N_24497,N_24498,N_24499,N_24502,N_24504,N_24505,N_24506,N_24508,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24519,N_24521,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24547,N_24550,N_24551,N_24554,N_24555,N_24556,N_24557,N_24559,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24571,N_24573,N_24574,N_24575,N_24577,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24588,N_24589,N_24591,N_24593,N_24594,N_24596,N_24599,N_24601,N_24602,N_24603,N_24605,N_24608,N_24609,N_24610,N_24612,N_24613,N_24617,N_24618,N_24619,N_24621,N_24622,N_24623,N_24624,N_24626,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24637,N_24638,N_24640,N_24641,N_24642,N_24645,N_24646,N_24647,N_24650,N_24651,N_24652,N_24653,N_24654,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24668,N_24669,N_24670,N_24672,N_24673,N_24674,N_24675,N_24678,N_24680,N_24681,N_24683,N_24684,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24706,N_24707,N_24710,N_24711,N_24712,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24721,N_24722,N_24723,N_24725,N_24727,N_24728,N_24731,N_24732,N_24733,N_24734,N_24735,N_24737,N_24738,N_24740,N_24741,N_24743,N_24744,N_24745,N_24746,N_24747,N_24749,N_24750,N_24753,N_24754,N_24756,N_24757,N_24758,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24767,N_24771,N_24774,N_24775,N_24776,N_24777,N_24779,N_24782,N_24784,N_24785,N_24786,N_24788,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24800,N_24801,N_24802,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24811,N_24812,N_24813,N_24814,N_24815,N_24818,N_24819,N_24824,N_24825,N_24826,N_24828,N_24830,N_24832,N_24833,N_24834,N_24836,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24849,N_24853,N_24854,N_24855,N_24857,N_24858,N_24859,N_24863,N_24865,N_24867,N_24870,N_24871,N_24872,N_24873,N_24875,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24887,N_24888,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24910,N_24915,N_24917,N_24919,N_24921,N_24922,N_24923,N_24925,N_24926,N_24927,N_24929,N_24931,N_24932,N_24933,N_24934,N_24936,N_24937,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24950,N_24951,N_24952,N_24953,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24963,N_24964,N_24965,N_24967,N_24968,N_24969,N_24971,N_24972,N_24973,N_24974,N_24975,N_24977,N_24982,N_24983,N_24984,N_24987,N_24988,N_24989,N_24990,N_24994,N_24995,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25006,N_25007,N_25009,N_25010,N_25012,N_25014,N_25017,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25035,N_25037,N_25039,N_25041,N_25043,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25054,N_25055,N_25056,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25076,N_25077,N_25078,N_25081,N_25082,N_25083,N_25089,N_25090,N_25091,N_25092,N_25094,N_25095,N_25096,N_25099,N_25100,N_25102,N_25103,N_25104,N_25105,N_25106,N_25109,N_25110,N_25111,N_25116,N_25118,N_25119,N_25120,N_25124,N_25125,N_25126,N_25127,N_25128,N_25130,N_25133,N_25134,N_25135,N_25138,N_25141,N_25142,N_25144,N_25147,N_25149,N_25150,N_25151,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25160,N_25162,N_25164,N_25165,N_25170,N_25171,N_25172,N_25174,N_25176,N_25177,N_25178,N_25179,N_25180,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25192,N_25194,N_25196,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25209,N_25210,N_25211,N_25213,N_25215,N_25216,N_25217,N_25218,N_25219,N_25221,N_25222,N_25224,N_25225,N_25226,N_25227,N_25229,N_25231,N_25232,N_25233,N_25236,N_25237,N_25238,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25250,N_25251,N_25252,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25263,N_25264,N_25265,N_25266,N_25267,N_25269,N_25271,N_25272,N_25275,N_25276,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25287,N_25288,N_25290,N_25291,N_25293,N_25294,N_25296,N_25297,N_25298,N_25299,N_25300,N_25302,N_25303,N_25304,N_25305,N_25307,N_25309,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25320,N_25321,N_25323,N_25324,N_25325,N_25327,N_25328,N_25330,N_25331,N_25333,N_25334,N_25335,N_25337,N_25338,N_25340,N_25341,N_25342,N_25344,N_25345,N_25346,N_25347,N_25348,N_25350,N_25351,N_25352,N_25353,N_25354,N_25356,N_25357,N_25359,N_25360,N_25361,N_25363,N_25364,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25374,N_25375,N_25377,N_25379,N_25380,N_25381,N_25382,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25396,N_25397,N_25398,N_25399,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25411,N_25412,N_25413,N_25414,N_25416,N_25417,N_25420,N_25424,N_25425,N_25426,N_25427,N_25429,N_25430,N_25431,N_25432,N_25433,N_25436,N_25438,N_25439,N_25440,N_25441,N_25444,N_25446,N_25447,N_25449,N_25450,N_25451,N_25452,N_25454,N_25455,N_25456,N_25457,N_25458,N_25461,N_25462,N_25463,N_25464,N_25465,N_25467,N_25469,N_25470,N_25471,N_25472,N_25474,N_25475,N_25476,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25489,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25500,N_25501,N_25502,N_25503,N_25505,N_25506,N_25509,N_25512,N_25513,N_25514,N_25515,N_25517,N_25518,N_25520,N_25522,N_25523,N_25525,N_25526,N_25527,N_25529,N_25530,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25539,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25549,N_25550,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25561,N_25562,N_25566,N_25567,N_25568,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25579,N_25580,N_25581,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25591,N_25592,N_25593,N_25594,N_25596,N_25597,N_25599,N_25600,N_25601,N_25602,N_25603,N_25606,N_25608,N_25609,N_25610,N_25611,N_25612,N_25614,N_25615,N_25616,N_25619,N_25620,N_25621,N_25622,N_25625,N_25626,N_25627,N_25629,N_25630,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25639,N_25640,N_25642,N_25644,N_25645,N_25646,N_25647,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25661,N_25662,N_25663,N_25664,N_25665,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25677,N_25679,N_25681,N_25682,N_25684,N_25685,N_25687,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25700,N_25702,N_25707,N_25708,N_25709,N_25710,N_25711,N_25715,N_25716,N_25718,N_25720,N_25721,N_25722,N_25724,N_25731,N_25732,N_25733,N_25734,N_25736,N_25738,N_25739,N_25741,N_25743,N_25744,N_25745,N_25747,N_25748,N_25749,N_25751,N_25753,N_25754,N_25756,N_25758,N_25759,N_25761,N_25762,N_25763,N_25766,N_25767,N_25768,N_25769,N_25770,N_25772,N_25776,N_25777,N_25778,N_25779,N_25781,N_25783,N_25785,N_25786,N_25787,N_25788,N_25789,N_25791,N_25792,N_25793,N_25794,N_25796,N_25798,N_25799,N_25800,N_25801,N_25804,N_25805,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25815,N_25816,N_25818,N_25821,N_25823,N_25824,N_25825,N_25828,N_25829,N_25830,N_25831,N_25833,N_25834,N_25835,N_25836,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25848,N_25850,N_25851,N_25853,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25867,N_25868,N_25870,N_25871,N_25872,N_25873,N_25875,N_25878,N_25879,N_25880,N_25881,N_25882,N_25885,N_25886,N_25888,N_25890,N_25892,N_25893,N_25895,N_25896,N_25900,N_25903,N_25904,N_25905,N_25906,N_25907,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25919,N_25922,N_25925,N_25927,N_25928,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25951,N_25952,N_25954,N_25955,N_25956,N_25957,N_25958,N_25960,N_25961,N_25963,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25973,N_25974,N_25976,N_25977,N_25978,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25989,N_25990,N_25991,N_25992,N_25994,N_25995,N_25997,N_25998,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26007,N_26008,N_26009,N_26011,N_26012,N_26013,N_26017,N_26018,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26039,N_26040,N_26041,N_26042,N_26044,N_26046,N_26049,N_26051,N_26052,N_26054,N_26055,N_26057,N_26059,N_26060,N_26062,N_26063,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26073,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26086,N_26088,N_26089,N_26090,N_26091,N_26092,N_26094,N_26095,N_26097,N_26098,N_26099,N_26100,N_26101,N_26103,N_26104,N_26105,N_26106,N_26108,N_26109,N_26112,N_26115,N_26117,N_26118,N_26119,N_26120,N_26122,N_26123,N_26124,N_26127,N_26128,N_26129,N_26131,N_26132,N_26133,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26143,N_26145,N_26147,N_26148,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26159,N_26161,N_26163,N_26164,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26173,N_26175,N_26178,N_26179,N_26180,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26192,N_26194,N_26195,N_26197,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26209,N_26210,N_26213,N_26215,N_26219,N_26220,N_26221,N_26222,N_26225,N_26226,N_26227,N_26228,N_26229,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26238,N_26240,N_26243,N_26244,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26257,N_26258,N_26261,N_26262,N_26263,N_26265,N_26266,N_26267,N_26269,N_26270,N_26271,N_26272,N_26274,N_26278,N_26280,N_26281,N_26283,N_26284,N_26285,N_26286,N_26288,N_26289,N_26291,N_26292,N_26294,N_26295,N_26296,N_26298,N_26299,N_26300,N_26303,N_26304,N_26305,N_26306,N_26307,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26316,N_26317,N_26319,N_26320,N_26322,N_26323,N_26324,N_26325,N_26326,N_26328,N_26329,N_26330,N_26331,N_26333,N_26334,N_26335,N_26336,N_26338,N_26340,N_26341,N_26342,N_26343,N_26344,N_26347,N_26349,N_26352,N_26353,N_26355,N_26356,N_26357,N_26360,N_26361,N_26362,N_26364,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26389,N_26390,N_26393,N_26396,N_26398,N_26399,N_26400,N_26401,N_26402,N_26404,N_26405,N_26406,N_26408,N_26409,N_26410,N_26411,N_26413,N_26415,N_26417,N_26418,N_26420,N_26421,N_26422,N_26423,N_26424,N_26426,N_26427,N_26428,N_26429,N_26431,N_26432,N_26433,N_26437,N_26438,N_26439,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26449,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26460,N_26461,N_26462,N_26463,N_26465,N_26466,N_26467,N_26468,N_26470,N_26471,N_26472,N_26474,N_26475,N_26476,N_26478,N_26479,N_26480,N_26482,N_26484,N_26487,N_26490,N_26491,N_26492,N_26493,N_26494,N_26496,N_26497,N_26498,N_26499,N_26501,N_26502,N_26504,N_26509,N_26510,N_26512,N_26513,N_26516,N_26517,N_26518,N_26520,N_26521,N_26522,N_26523,N_26525,N_26527,N_26529,N_26531,N_26533,N_26535,N_26536,N_26537,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26549,N_26551,N_26552,N_26554,N_26555,N_26556,N_26557,N_26558,N_26560,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26569,N_26571,N_26572,N_26574,N_26575,N_26576,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26588,N_26589,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26606,N_26607,N_26609,N_26610,N_26611,N_26613,N_26614,N_26615,N_26616,N_26618,N_26619,N_26620,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26634,N_26635,N_26636,N_26637,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26660,N_26661,N_26662,N_26663,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26686,N_26687,N_26688,N_26689,N_26690,N_26692,N_26694,N_26695,N_26697,N_26700,N_26701,N_26703,N_26705,N_26707,N_26709,N_26710,N_26712,N_26714,N_26715,N_26716,N_26717,N_26719,N_26722,N_26723,N_26724,N_26726,N_26727,N_26728,N_26730,N_26731,N_26732,N_26734,N_26735,N_26737,N_26738,N_26742,N_26743,N_26745,N_26746,N_26747,N_26749,N_26753,N_26754,N_26755,N_26757,N_26758,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26773,N_26775,N_26776,N_26779,N_26780,N_26781,N_26783,N_26784,N_26785,N_26787,N_26788,N_26789,N_26790,N_26792,N_26793,N_26794,N_26796,N_26798,N_26799,N_26800,N_26801,N_26804,N_26806,N_26809,N_26810,N_26812,N_26815,N_26816,N_26819,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26843,N_26846,N_26847,N_26849,N_26850,N_26851,N_26852,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26862,N_26863,N_26864,N_26866,N_26867,N_26868,N_26869,N_26871,N_26872,N_26874,N_26875,N_26878,N_26880,N_26881,N_26883,N_26885,N_26886,N_26890,N_26891,N_26894,N_26895,N_26897,N_26898,N_26900,N_26901,N_26902,N_26904,N_26905,N_26906,N_26909,N_26910,N_26912,N_26913,N_26914,N_26915,N_26918,N_26920,N_26921,N_26922,N_26923,N_26924,N_26927,N_26928,N_26931,N_26932,N_26933,N_26935,N_26938,N_26939,N_26940,N_26943,N_26944,N_26947,N_26948,N_26949,N_26951,N_26952,N_26953,N_26955,N_26956,N_26957,N_26958,N_26959,N_26962,N_26964,N_26965,N_26966,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26989,N_26992,N_26993,N_26995,N_26996,N_26997,N_26999,N_27003,N_27004,N_27007,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27020,N_27021,N_27024,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27040,N_27041,N_27044,N_27045,N_27046,N_27047,N_27050,N_27051,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27060,N_27061,N_27062,N_27063,N_27065,N_27066,N_27067,N_27068,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27081,N_27082,N_27084,N_27086,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27097,N_27098,N_27099,N_27100,N_27101,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27111,N_27112,N_27113,N_27115,N_27116,N_27117,N_27119,N_27121,N_27122,N_27123,N_27124,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27133,N_27134,N_27135,N_27136,N_27138,N_27140,N_27141,N_27142,N_27144,N_27146,N_27148,N_27150,N_27151,N_27154,N_27155,N_27156,N_27157,N_27158,N_27160,N_27161,N_27162,N_27163,N_27166,N_27167,N_27168,N_27170,N_27171,N_27172,N_27173,N_27176,N_27178,N_27179,N_27180,N_27183,N_27185,N_27186,N_27187,N_27188,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27200,N_27201,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27217,N_27218,N_27219,N_27220,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27231,N_27233,N_27234,N_27235,N_27237,N_27238,N_27241,N_27242,N_27243,N_27247,N_27248,N_27249,N_27253,N_27254,N_27255,N_27257,N_27258,N_27259,N_27260,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27274,N_27275,N_27278,N_27280,N_27281,N_27282,N_27285,N_27287,N_27288,N_27289,N_27291,N_27292,N_27294,N_27295,N_27296,N_27297,N_27298,N_27300,N_27301,N_27302,N_27304,N_27306,N_27307,N_27308,N_27310,N_27311,N_27312,N_27313,N_27315,N_27316,N_27317,N_27318,N_27319,N_27321,N_27322,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27333,N_27334,N_27335,N_27336,N_27337,N_27339,N_27342,N_27343,N_27344,N_27346,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27357,N_27359,N_27360,N_27361,N_27363,N_27364,N_27365,N_27366,N_27367,N_27369,N_27371,N_27372,N_27373,N_27375,N_27376,N_27378,N_27379,N_27380,N_27381,N_27383,N_27384,N_27386,N_27387,N_27390,N_27391,N_27393,N_27394,N_27395,N_27396,N_27397,N_27399,N_27401,N_27402,N_27403,N_27404,N_27405,N_27407,N_27409,N_27410,N_27411,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27421,N_27424,N_27425,N_27426,N_27427,N_27429,N_27430,N_27432,N_27434,N_27435,N_27436,N_27438,N_27439,N_27441,N_27442,N_27443,N_27445,N_27446,N_27449,N_27450,N_27451,N_27455,N_27462,N_27463,N_27465,N_27467,N_27468,N_27469,N_27470,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27482,N_27483,N_27484,N_27487,N_27488,N_27491,N_27492,N_27493,N_27494,N_27495,N_27497,N_27498,N_27500,N_27501,N_27502,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27512,N_27513,N_27517,N_27518,N_27520,N_27522,N_27523,N_27525,N_27528,N_27529,N_27530,N_27531,N_27532,N_27535,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27544,N_27545,N_27548,N_27551,N_27555,N_27556,N_27557,N_27558,N_27559,N_27562,N_27563,N_27564,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27573,N_27574,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27595,N_27596,N_27598,N_27603,N_27604,N_27605,N_27607,N_27608,N_27609,N_27611,N_27612,N_27614,N_27616,N_27617,N_27618,N_27620,N_27623,N_27624,N_27625,N_27626,N_27628,N_27629,N_27630,N_27631,N_27632,N_27634,N_27635,N_27636,N_27637,N_27639,N_27640,N_27641,N_27644,N_27645,N_27646,N_27647,N_27648,N_27650,N_27651,N_27653,N_27654,N_27656,N_27658,N_27659,N_27660,N_27663,N_27664,N_27665,N_27666,N_27667,N_27669,N_27670,N_27673,N_27674,N_27675,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27687,N_27689,N_27690,N_27691,N_27692,N_27695,N_27697,N_27700,N_27701,N_27702,N_27703,N_27706,N_27707,N_27709,N_27712,N_27714,N_27716,N_27719,N_27720,N_27721,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27737,N_27738,N_27739,N_27741,N_27742,N_27743,N_27746,N_27748,N_27749,N_27751,N_27753,N_27754,N_27755,N_27756,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27777,N_27778,N_27780,N_27781,N_27782,N_27783,N_27785,N_27786,N_27787,N_27789,N_27790,N_27791,N_27793,N_27794,N_27797,N_27800,N_27802,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27816,N_27817,N_27818,N_27821,N_27823,N_27824,N_27826,N_27827,N_27829,N_27833,N_27834,N_27836,N_27838,N_27840,N_27841,N_27842,N_27845,N_27846,N_27847,N_27849,N_27851,N_27852,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27867,N_27869,N_27870,N_27871,N_27872,N_27873,N_27875,N_27876,N_27877,N_27879,N_27880,N_27881,N_27882,N_27883,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27896,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27923,N_27925,N_27926,N_27927,N_27930,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27946,N_27947,N_27948,N_27951,N_27952,N_27953,N_27954,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27965,N_27966,N_27968,N_27969,N_27972,N_27973,N_27974,N_27975,N_27979,N_27981,N_27982,N_27983,N_27984,N_27985,N_27987,N_27988,N_27989,N_27990,N_27991,N_27993,N_27995,N_27997,N_27998,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28010,N_28012,N_28013,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28024,N_28025,N_28026,N_28028,N_28029,N_28032,N_28033,N_28035,N_28036,N_28038,N_28039,N_28041,N_28045,N_28047,N_28048,N_28049,N_28050,N_28054,N_28055,N_28056,N_28057,N_28058,N_28060,N_28061,N_28062,N_28066,N_28067,N_28068,N_28069,N_28071,N_28072,N_28073,N_28075,N_28076,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28101,N_28104,N_28106,N_28108,N_28111,N_28112,N_28114,N_28117,N_28118,N_28119,N_28122,N_28125,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28135,N_28137,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28146,N_28147,N_28148,N_28149,N_28150,N_28152,N_28153,N_28154,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28183,N_28184,N_28185,N_28187,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28201,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28210,N_28211,N_28212,N_28213,N_28214,N_28217,N_28218,N_28219,N_28223,N_28224,N_28225,N_28226,N_28229,N_28230,N_28231,N_28234,N_28235,N_28236,N_28237,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28249,N_28251,N_28252,N_28253,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28265,N_28267,N_28268,N_28270,N_28271,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28308,N_28309,N_28310,N_28312,N_28313,N_28315,N_28316,N_28317,N_28322,N_28324,N_28326,N_28327,N_28328,N_28330,N_28331,N_28332,N_28333,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28344,N_28345,N_28347,N_28349,N_28350,N_28352,N_28353,N_28355,N_28356,N_28358,N_28359,N_28363,N_28364,N_28365,N_28367,N_28368,N_28369,N_28370,N_28371,N_28373,N_28375,N_28376,N_28378,N_28380,N_28381,N_28383,N_28389,N_28390,N_28391,N_28392,N_28393,N_28398,N_28399,N_28400,N_28403,N_28404,N_28405,N_28406,N_28409,N_28410,N_28411,N_28412,N_28413,N_28415,N_28416,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28428,N_28431,N_28433,N_28434,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28461,N_28462,N_28463,N_28465,N_28466,N_28467,N_28469,N_28470,N_28471,N_28472,N_28473,N_28475,N_28476,N_28478,N_28479,N_28481,N_28483,N_28484,N_28485,N_28486,N_28488,N_28490,N_28492,N_28493,N_28494,N_28496,N_28497,N_28498,N_28499,N_28500,N_28503,N_28504,N_28505,N_28506,N_28507,N_28509,N_28510,N_28516,N_28519,N_28520,N_28521,N_28523,N_28528,N_28529,N_28530,N_28531,N_28532,N_28534,N_28535,N_28540,N_28541,N_28542,N_28543,N_28544,N_28548,N_28550,N_28552,N_28553,N_28554,N_28555,N_28556,N_28559,N_28561,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28573,N_28574,N_28577,N_28579,N_28580,N_28581,N_28583,N_28584,N_28585,N_28586,N_28588,N_28589,N_28592,N_28593,N_28594,N_28596,N_28597,N_28598,N_28600,N_28602,N_28604,N_28605,N_28606,N_28608,N_28610,N_28611,N_28613,N_28614,N_28616,N_28618,N_28620,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28629,N_28632,N_28633,N_28634,N_28636,N_28637,N_28638,N_28640,N_28641,N_28642,N_28644,N_28646,N_28647,N_28650,N_28651,N_28654,N_28655,N_28657,N_28658,N_28660,N_28661,N_28662,N_28663,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28677,N_28678,N_28679,N_28680,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28693,N_28694,N_28695,N_28696,N_28698,N_28699,N_28703,N_28704,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28721,N_28724,N_28725,N_28726,N_28727,N_28728,N_28730,N_28731,N_28733,N_28734,N_28736,N_28737,N_28738,N_28740,N_28742,N_28743,N_28744,N_28746,N_28747,N_28748,N_28749,N_28750,N_28752,N_28753,N_28754,N_28756,N_28759,N_28760,N_28762,N_28763,N_28765,N_28766,N_28768,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28783,N_28784,N_28785,N_28787,N_28788,N_28789,N_28791,N_28792,N_28794,N_28796,N_28798,N_28799,N_28800,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28810,N_28811,N_28812,N_28813,N_28814,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28830,N_28832,N_28833,N_28835,N_28837,N_28839,N_28840,N_28841,N_28843,N_28844,N_28846,N_28847,N_28850,N_28851,N_28852,N_28856,N_28857,N_28858,N_28859,N_28861,N_28862,N_28864,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28874,N_28876,N_28878,N_28880,N_28881,N_28882,N_28883,N_28884,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28893,N_28895,N_28897,N_28898,N_28899,N_28900,N_28901,N_28903,N_28904,N_28905,N_28906,N_28907,N_28910,N_28911,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28920,N_28922,N_28923,N_28924,N_28925,N_28926,N_28928,N_28929,N_28930,N_28931,N_28933,N_28934,N_28937,N_28938,N_28941,N_28943,N_28945,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28956,N_28957,N_28959,N_28961,N_28964,N_28965,N_28966,N_28968,N_28970,N_28971,N_28975,N_28977,N_28979,N_28980,N_28981,N_28983,N_28984,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28998,N_28999,N_29000,N_29001,N_29003,N_29004,N_29005,N_29006,N_29009,N_29012,N_29013,N_29015,N_29016,N_29017,N_29021,N_29022,N_29024,N_29025,N_29028,N_29029,N_29030,N_29031,N_29032,N_29034,N_29037,N_29038,N_29040,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29050,N_29051,N_29052,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29064,N_29065,N_29066,N_29067,N_29068,N_29070,N_29072,N_29073,N_29074,N_29075,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29085,N_29086,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29101,N_29103,N_29104,N_29106,N_29107,N_29113,N_29115,N_29116,N_29117,N_29118,N_29119,N_29121,N_29122,N_29123,N_29124,N_29125,N_29127,N_29129,N_29135,N_29136,N_29140,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29149,N_29150,N_29151,N_29153,N_29155,N_29156,N_29157,N_29158,N_29159,N_29161,N_29162,N_29165,N_29166,N_29168,N_29169,N_29172,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29185,N_29186,N_29187,N_29188,N_29189,N_29192,N_29193,N_29195,N_29197,N_29198,N_29201,N_29203,N_29205,N_29207,N_29208,N_29209,N_29211,N_29212,N_29214,N_29215,N_29216,N_29217,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29231,N_29232,N_29234,N_29235,N_29238,N_29239,N_29241,N_29242,N_29244,N_29245,N_29246,N_29247,N_29250,N_29251,N_29253,N_29255,N_29256,N_29257,N_29258,N_29261,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29281,N_29282,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29298,N_29299,N_29300,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29310,N_29311,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29323,N_29325,N_29326,N_29328,N_29329,N_29330,N_29331,N_29332,N_29334,N_29335,N_29337,N_29338,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29351,N_29353,N_29354,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29369,N_29370,N_29373,N_29374,N_29375,N_29376,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29387,N_29389,N_29391,N_29392,N_29393,N_29394,N_29396,N_29397,N_29398,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29407,N_29409,N_29410,N_29413,N_29415,N_29416,N_29417,N_29418,N_29419,N_29421,N_29423,N_29424,N_29425,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29437,N_29438,N_29439,N_29441,N_29443,N_29444,N_29445,N_29446,N_29447,N_29450,N_29451,N_29452,N_29455,N_29458,N_29459,N_29462,N_29463,N_29465,N_29467,N_29468,N_29470,N_29473,N_29474,N_29475,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29491,N_29494,N_29495,N_29496,N_29499,N_29501,N_29502,N_29504,N_29507,N_29509,N_29510,N_29511,N_29514,N_29515,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29539,N_29541,N_29542,N_29544,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29578,N_29580,N_29582,N_29583,N_29584,N_29586,N_29588,N_29589,N_29590,N_29591,N_29592,N_29594,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29603,N_29604,N_29606,N_29607,N_29608,N_29609,N_29610,N_29612,N_29613,N_29617,N_29619,N_29620,N_29621,N_29622,N_29624,N_29625,N_29626,N_29628,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29642,N_29643,N_29644,N_29646,N_29647,N_29648,N_29649,N_29650,N_29652,N_29653,N_29655,N_29658,N_29660,N_29661,N_29663,N_29664,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29683,N_29685,N_29688,N_29689,N_29690,N_29692,N_29693,N_29694,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29705,N_29706,N_29707,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29717,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29744,N_29746,N_29747,N_29749,N_29750,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29767,N_29771,N_29772,N_29773,N_29774,N_29775,N_29777,N_29778,N_29779,N_29780,N_29781,N_29784,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29796,N_29797,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29813,N_29816,N_29817,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29826,N_29827,N_29828,N_29830,N_29831,N_29832,N_29837,N_29838,N_29839,N_29841,N_29842,N_29843,N_29844,N_29848,N_29849,N_29850,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29860,N_29863,N_29864,N_29865,N_29866,N_29867,N_29869,N_29870,N_29871,N_29872,N_29875,N_29876,N_29877,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29886,N_29887,N_29891,N_29893,N_29895,N_29896,N_29897,N_29898,N_29899,N_29901,N_29902,N_29905,N_29906,N_29907,N_29908,N_29911,N_29912,N_29913,N_29914,N_29915,N_29918,N_29919,N_29923,N_29925,N_29926,N_29927,N_29929,N_29932,N_29933,N_29934,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29957,N_29958,N_29959,N_29960,N_29961,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29974,N_29975,N_29976,N_29978,N_29980,N_29981,N_29983,N_29984,N_29986,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29995,N_29996,N_29998;
and U0 (N_0,In_2283,In_952);
nand U1 (N_1,In_2221,In_2170);
and U2 (N_2,In_161,In_1798);
or U3 (N_3,In_939,In_2709);
or U4 (N_4,In_2760,In_396);
and U5 (N_5,In_961,In_2713);
nand U6 (N_6,In_2467,In_1594);
nor U7 (N_7,In_1925,In_1879);
or U8 (N_8,In_351,In_2062);
or U9 (N_9,In_76,In_1801);
nor U10 (N_10,In_889,In_359);
or U11 (N_11,In_1061,In_1201);
and U12 (N_12,In_428,In_1101);
and U13 (N_13,In_2448,In_2483);
and U14 (N_14,In_2823,In_67);
and U15 (N_15,In_444,In_2535);
and U16 (N_16,In_339,In_392);
nor U17 (N_17,In_18,In_1397);
nand U18 (N_18,In_943,In_1804);
nand U19 (N_19,In_2345,In_1107);
and U20 (N_20,In_1122,In_703);
or U21 (N_21,In_1985,In_518);
and U22 (N_22,In_2039,In_464);
and U23 (N_23,In_852,In_661);
and U24 (N_24,In_2788,In_2601);
or U25 (N_25,In_915,In_1001);
or U26 (N_26,In_1547,In_822);
nand U27 (N_27,In_818,In_2817);
nor U28 (N_28,In_483,In_1639);
or U29 (N_29,In_2209,In_2860);
and U30 (N_30,In_1981,In_1811);
and U31 (N_31,In_1419,In_1288);
nor U32 (N_32,In_2060,In_1095);
or U33 (N_33,In_167,In_1004);
and U34 (N_34,In_1672,In_2637);
nor U35 (N_35,In_305,In_1293);
nand U36 (N_36,In_264,In_272);
and U37 (N_37,In_2832,In_2123);
or U38 (N_38,In_1844,In_1545);
nor U39 (N_39,In_311,In_755);
or U40 (N_40,In_240,In_1439);
or U41 (N_41,In_448,In_2865);
nor U42 (N_42,In_761,In_37);
or U43 (N_43,In_698,In_813);
or U44 (N_44,In_2482,In_2631);
and U45 (N_45,In_1418,In_1366);
or U46 (N_46,In_1992,In_206);
or U47 (N_47,In_2936,In_1889);
nand U48 (N_48,In_1258,In_2449);
or U49 (N_49,In_2479,In_217);
nor U50 (N_50,In_1239,In_2340);
nor U51 (N_51,In_1161,In_2789);
nor U52 (N_52,In_1148,In_2462);
or U53 (N_53,In_417,In_2566);
and U54 (N_54,In_2643,In_82);
nor U55 (N_55,In_2526,In_2412);
nand U56 (N_56,In_2762,In_225);
nand U57 (N_57,In_2879,In_54);
or U58 (N_58,In_1822,In_110);
nor U59 (N_59,In_2026,In_2066);
or U60 (N_60,In_2228,In_1349);
nor U61 (N_61,In_2584,In_960);
nand U62 (N_62,In_1245,In_1338);
or U63 (N_63,In_834,In_1323);
nand U64 (N_64,In_2282,In_2811);
and U65 (N_65,In_2249,In_1238);
or U66 (N_66,In_2125,In_2935);
nand U67 (N_67,In_974,In_2986);
nor U68 (N_68,In_1795,In_1387);
or U69 (N_69,In_1880,In_2528);
or U70 (N_70,In_101,In_2881);
or U71 (N_71,In_1799,In_2357);
and U72 (N_72,In_2710,In_17);
xnor U73 (N_73,In_2518,In_474);
and U74 (N_74,In_602,In_222);
nand U75 (N_75,In_154,In_919);
or U76 (N_76,In_2645,In_651);
or U77 (N_77,In_2147,In_2625);
or U78 (N_78,In_466,In_1946);
or U79 (N_79,In_2044,In_2155);
or U80 (N_80,In_1021,In_1763);
and U81 (N_81,In_789,In_425);
xnor U82 (N_82,In_1993,In_1678);
or U83 (N_83,In_182,In_1566);
nor U84 (N_84,In_528,In_1028);
or U85 (N_85,In_512,In_729);
nor U86 (N_86,In_1104,In_713);
nor U87 (N_87,In_2609,In_2399);
nor U88 (N_88,In_2852,In_2627);
and U89 (N_89,In_197,In_310);
nor U90 (N_90,In_1688,In_918);
nand U91 (N_91,In_2456,In_1048);
nor U92 (N_92,In_2966,In_1908);
nand U93 (N_93,In_1573,In_220);
nand U94 (N_94,In_2910,In_2900);
nor U95 (N_95,In_493,In_1731);
nor U96 (N_96,In_1394,In_1863);
or U97 (N_97,In_1308,In_2501);
and U98 (N_98,In_656,In_2670);
and U99 (N_99,In_733,In_437);
or U100 (N_100,In_838,In_2604);
and U101 (N_101,In_2455,In_1666);
nand U102 (N_102,In_979,In_1110);
nor U103 (N_103,In_242,In_285);
nand U104 (N_104,In_779,In_883);
nand U105 (N_105,In_1559,In_1489);
xor U106 (N_106,In_2049,In_2752);
and U107 (N_107,In_843,In_1528);
nand U108 (N_108,In_2263,In_117);
nor U109 (N_109,In_2262,In_1959);
nand U110 (N_110,In_1907,In_633);
nand U111 (N_111,In_1139,In_587);
nand U112 (N_112,In_2746,In_160);
nand U113 (N_113,In_2094,In_219);
nand U114 (N_114,In_1120,In_1793);
nor U115 (N_115,In_2682,In_2949);
or U116 (N_116,In_1674,In_1128);
or U117 (N_117,In_758,In_519);
nor U118 (N_118,In_2215,In_1124);
nor U119 (N_119,In_1249,In_840);
nor U120 (N_120,In_1466,In_2838);
and U121 (N_121,In_1125,In_2715);
nand U122 (N_122,In_77,In_1170);
nor U123 (N_123,In_1949,In_957);
nor U124 (N_124,In_844,In_1442);
nor U125 (N_125,In_2397,In_2106);
nor U126 (N_126,In_368,In_2976);
and U127 (N_127,In_20,In_583);
nor U128 (N_128,In_566,In_1003);
nor U129 (N_129,In_2320,In_1924);
nand U130 (N_130,In_1613,In_454);
nor U131 (N_131,In_1138,In_1108);
and U132 (N_132,In_1824,In_2260);
or U133 (N_133,In_97,In_1734);
and U134 (N_134,In_2922,In_1851);
and U135 (N_135,In_649,In_1092);
nand U136 (N_136,In_1585,In_1284);
nand U137 (N_137,In_1029,In_2488);
nand U138 (N_138,In_2258,In_520);
or U139 (N_139,In_2723,In_1752);
and U140 (N_140,In_1742,In_395);
and U141 (N_141,In_2565,In_1060);
and U142 (N_142,In_1381,In_643);
or U143 (N_143,In_2463,In_1750);
and U144 (N_144,In_2697,In_684);
or U145 (N_145,In_2222,In_880);
and U146 (N_146,In_2248,In_2395);
nand U147 (N_147,In_215,In_694);
or U148 (N_148,In_1624,In_2621);
nor U149 (N_149,In_2906,In_1701);
nand U150 (N_150,In_1237,In_2265);
or U151 (N_151,In_2524,In_741);
nor U152 (N_152,In_2800,In_1205);
nand U153 (N_153,In_2694,In_207);
or U154 (N_154,In_878,In_2751);
nor U155 (N_155,In_760,In_301);
and U156 (N_156,In_2580,In_2116);
nand U157 (N_157,In_704,In_2748);
and U158 (N_158,In_1438,In_923);
nand U159 (N_159,In_1414,In_2154);
nand U160 (N_160,In_1667,In_2770);
nand U161 (N_161,In_699,In_2538);
nor U162 (N_162,In_1350,In_2591);
and U163 (N_163,In_679,In_531);
or U164 (N_164,In_588,In_2046);
nor U165 (N_165,In_2515,In_398);
and U166 (N_166,In_2257,In_1073);
nor U167 (N_167,In_1789,In_2998);
or U168 (N_168,In_1459,In_1272);
or U169 (N_169,In_2310,In_440);
or U170 (N_170,In_1332,In_2909);
and U171 (N_171,In_500,In_12);
and U172 (N_172,In_1541,In_2244);
or U173 (N_173,In_1670,In_2065);
nand U174 (N_174,In_2912,In_1204);
or U175 (N_175,In_1448,In_1151);
and U176 (N_176,In_1597,In_1754);
and U177 (N_177,In_36,In_2562);
and U178 (N_178,In_1746,In_2045);
and U179 (N_179,In_155,In_1227);
nand U180 (N_180,In_2992,In_1867);
nor U181 (N_181,In_969,In_2204);
nand U182 (N_182,In_599,In_1885);
and U183 (N_183,In_763,In_744);
nand U184 (N_184,In_2465,In_1369);
and U185 (N_185,In_1821,In_935);
or U186 (N_186,In_1966,In_2989);
nand U187 (N_187,In_1089,In_2272);
nand U188 (N_188,In_1728,In_2613);
and U189 (N_189,In_1479,In_781);
or U190 (N_190,In_1725,In_2680);
nand U191 (N_191,In_1391,In_2899);
nand U192 (N_192,In_127,In_2761);
and U193 (N_193,In_1546,In_2707);
xnor U194 (N_194,In_435,In_176);
and U195 (N_195,In_2203,In_542);
or U196 (N_196,In_1719,In_1625);
and U197 (N_197,In_1134,In_1978);
or U198 (N_198,In_1434,In_1552);
nor U199 (N_199,In_1888,In_992);
nand U200 (N_200,In_1032,In_2575);
or U201 (N_201,In_324,In_2348);
and U202 (N_202,In_2121,In_1916);
nor U203 (N_203,In_701,In_2740);
or U204 (N_204,In_857,In_2181);
and U205 (N_205,In_737,In_1972);
or U206 (N_206,In_625,In_2361);
nand U207 (N_207,In_2520,In_876);
or U208 (N_208,In_2275,In_1346);
nand U209 (N_209,In_1214,In_1361);
nor U210 (N_210,In_459,In_546);
and U211 (N_211,In_1891,In_2019);
nor U212 (N_212,In_35,In_1254);
or U213 (N_213,In_2496,In_1511);
nor U214 (N_214,In_244,In_491);
and U215 (N_215,In_58,In_1301);
and U216 (N_216,In_2122,In_2952);
and U217 (N_217,In_2166,In_2884);
nor U218 (N_218,In_2,In_2419);
or U219 (N_219,In_1650,In_1524);
nand U220 (N_220,In_1159,In_819);
nor U221 (N_221,In_1102,In_1392);
or U222 (N_222,In_2768,In_2880);
nand U223 (N_223,In_1020,In_1886);
nand U224 (N_224,In_2730,In_1975);
and U225 (N_225,In_1316,In_329);
or U226 (N_226,In_1222,In_2539);
nand U227 (N_227,In_463,In_263);
or U228 (N_228,In_1747,In_1026);
and U229 (N_229,In_190,In_564);
nand U230 (N_230,In_746,In_2117);
and U231 (N_231,In_1510,In_1112);
or U232 (N_232,In_2274,In_2938);
nor U233 (N_233,In_2163,In_2895);
and U234 (N_234,In_1808,In_1197);
nor U235 (N_235,In_2886,In_2537);
and U236 (N_236,In_1839,In_2440);
or U237 (N_237,In_125,In_1570);
and U238 (N_238,In_1034,In_2557);
nand U239 (N_239,In_2072,In_2527);
and U240 (N_240,In_2431,In_2224);
nor U241 (N_241,In_2634,In_600);
or U242 (N_242,In_2738,In_2574);
and U243 (N_243,In_2192,In_2338);
nor U244 (N_244,In_2716,In_1292);
or U245 (N_245,In_2600,In_2319);
and U246 (N_246,In_1266,In_268);
and U247 (N_247,In_2944,In_1996);
or U248 (N_248,In_949,In_2316);
and U249 (N_249,In_2299,In_2023);
nor U250 (N_250,In_971,In_279);
or U251 (N_251,In_1962,In_2371);
and U252 (N_252,In_2896,In_670);
or U253 (N_253,In_1603,In_348);
and U254 (N_254,In_628,In_836);
or U255 (N_255,In_1388,In_2514);
nor U256 (N_256,In_1873,In_2400);
and U257 (N_257,In_2599,In_296);
nor U258 (N_258,In_214,In_2835);
nor U259 (N_259,In_941,In_2350);
nor U260 (N_260,In_41,In_1958);
or U261 (N_261,In_2693,In_1923);
nor U262 (N_262,In_964,In_1109);
nand U263 (N_263,In_1567,In_2306);
nand U264 (N_264,In_2069,In_1760);
and U265 (N_265,In_1351,In_2383);
and U266 (N_266,In_1311,In_2516);
nor U267 (N_267,In_2688,In_2389);
or U268 (N_268,In_1454,In_189);
or U269 (N_269,In_2855,In_1321);
or U270 (N_270,In_2194,In_895);
and U271 (N_271,In_1607,In_2184);
and U272 (N_272,In_1035,In_2200);
and U273 (N_273,In_1711,In_2882);
nand U274 (N_274,In_1263,In_2165);
and U275 (N_275,In_2784,In_132);
nand U276 (N_276,In_2547,In_1800);
and U277 (N_277,In_1848,In_2644);
nor U278 (N_278,In_422,In_808);
or U279 (N_279,In_350,In_2076);
nand U280 (N_280,In_2152,In_886);
nand U281 (N_281,In_2169,In_480);
or U282 (N_282,In_1869,In_1582);
nand U283 (N_283,In_1297,In_2285);
nor U284 (N_284,In_1519,In_1598);
or U285 (N_285,In_371,In_2925);
and U286 (N_286,In_2372,In_2161);
nand U287 (N_287,In_707,In_1070);
and U288 (N_288,In_854,In_2632);
nand U289 (N_289,In_1832,In_2665);
nand U290 (N_290,In_292,In_201);
or U291 (N_291,In_1036,In_697);
nand U292 (N_292,In_2552,In_2726);
nand U293 (N_293,In_1997,In_1649);
nor U294 (N_294,In_2782,In_1553);
or U295 (N_295,In_859,In_2646);
or U296 (N_296,In_1841,In_275);
or U297 (N_297,In_2120,In_1481);
nand U298 (N_298,In_2425,In_254);
or U299 (N_299,In_2010,In_1192);
or U300 (N_300,In_318,In_708);
nor U301 (N_301,In_2003,In_1467);
nor U302 (N_302,In_2294,In_2111);
and U303 (N_303,In_1512,In_2517);
nor U304 (N_304,In_357,In_2377);
nor U305 (N_305,In_811,In_1770);
and U306 (N_306,In_2336,In_1665);
or U307 (N_307,In_1915,In_191);
and U308 (N_308,In_2022,In_1304);
or U309 (N_309,In_1372,In_962);
nor U310 (N_310,In_2783,In_38);
and U311 (N_311,In_950,In_109);
nor U312 (N_312,In_2616,In_340);
nand U313 (N_313,In_105,In_1508);
nand U314 (N_314,In_159,In_1240);
nand U315 (N_315,In_1939,In_907);
and U316 (N_316,In_175,In_1368);
nand U317 (N_317,In_1733,In_2522);
nand U318 (N_318,In_1160,In_629);
nor U319 (N_319,In_1934,In_1591);
and U320 (N_320,In_2541,In_2975);
or U321 (N_321,In_1098,In_615);
or U322 (N_322,In_2858,In_2423);
or U323 (N_323,In_2819,In_1922);
and U324 (N_324,In_650,In_1840);
or U325 (N_325,In_2287,In_1698);
nor U326 (N_326,In_800,In_934);
nor U327 (N_327,In_2284,In_1773);
and U328 (N_328,In_1951,In_1359);
or U329 (N_329,In_2027,In_618);
nor U330 (N_330,In_1890,In_1187);
and U331 (N_331,In_1378,In_342);
or U332 (N_332,In_685,In_56);
and U333 (N_333,In_484,In_997);
nor U334 (N_334,In_2826,In_163);
nand U335 (N_335,In_1684,In_15);
nand U336 (N_336,In_1445,In_11);
or U337 (N_337,In_710,In_2914);
nand U338 (N_338,In_784,In_180);
nor U339 (N_339,In_2772,In_2205);
nand U340 (N_340,In_1636,In_2491);
nand U341 (N_341,In_864,In_617);
nand U342 (N_342,In_556,In_2135);
and U343 (N_343,In_576,In_796);
nand U344 (N_344,In_2384,In_1347);
or U345 (N_345,In_2733,In_2341);
or U346 (N_346,In_471,In_1080);
nand U347 (N_347,In_794,In_2174);
nand U348 (N_348,In_198,In_2534);
nor U349 (N_349,In_2363,In_2421);
nor U350 (N_350,In_2302,In_1153);
nand U351 (N_351,In_229,In_1791);
or U352 (N_352,In_22,In_407);
nor U353 (N_353,In_1579,In_28);
or U354 (N_354,In_313,In_1450);
or U355 (N_355,In_2326,In_936);
nor U356 (N_356,In_1574,In_309);
and U357 (N_357,In_2785,In_2136);
nor U358 (N_358,In_1433,In_902);
and U359 (N_359,In_1903,In_1250);
or U360 (N_360,In_829,In_1283);
or U361 (N_361,In_2842,In_1371);
or U362 (N_362,In_2530,In_2824);
and U363 (N_363,In_91,In_1940);
or U364 (N_364,In_1947,In_1490);
nand U365 (N_365,In_2402,In_468);
nand U366 (N_366,In_2280,In_1919);
or U367 (N_367,In_258,In_524);
nor U368 (N_368,In_605,In_2335);
or U369 (N_369,In_2267,In_1954);
nor U370 (N_370,In_434,In_2671);
and U371 (N_371,In_94,In_1623);
or U372 (N_372,In_2484,In_2655);
and U373 (N_373,In_646,In_498);
nand U374 (N_374,In_560,In_1937);
nand U375 (N_375,In_2963,In_208);
or U376 (N_376,In_2814,In_2349);
or U377 (N_377,In_2756,In_1342);
nor U378 (N_378,In_1252,In_2521);
or U379 (N_379,In_2696,In_170);
nor U380 (N_380,In_2273,In_388);
and U381 (N_381,In_648,In_80);
nand U382 (N_382,In_443,In_1044);
nor U383 (N_383,In_2705,In_81);
and U384 (N_384,In_509,In_71);
nand U385 (N_385,In_644,In_1334);
nor U386 (N_386,In_2159,In_416);
nor U387 (N_387,In_2208,In_2322);
nor U388 (N_388,In_1162,In_1953);
nand U389 (N_389,In_975,In_2358);
nand U390 (N_390,In_2701,In_660);
nor U391 (N_391,In_1988,In_1364);
nor U392 (N_392,In_2666,In_355);
and U393 (N_393,In_1006,In_2633);
nand U394 (N_394,In_966,In_2853);
nand U395 (N_395,In_1052,In_2663);
and U396 (N_396,In_2226,In_447);
and U397 (N_397,In_1462,In_2093);
nand U398 (N_398,In_616,In_2764);
and U399 (N_399,In_2904,In_2129);
or U400 (N_400,In_1893,In_2352);
nor U401 (N_401,In_2151,In_1717);
xnor U402 (N_402,In_1732,In_597);
or U403 (N_403,In_319,In_1005);
nand U404 (N_404,In_284,In_2277);
nand U405 (N_405,In_2695,In_1175);
or U406 (N_406,In_104,In_1611);
and U407 (N_407,In_2930,In_575);
nand U408 (N_408,In_1782,In_1569);
nand U409 (N_409,In_2157,In_1259);
and U410 (N_410,In_1682,In_2825);
and U411 (N_411,In_1335,In_640);
or U412 (N_412,In_57,In_2640);
nor U413 (N_413,In_619,In_2105);
and U414 (N_414,In_2190,In_2589);
and U415 (N_415,In_1707,In_2243);
nor U416 (N_416,In_2686,In_1792);
or U417 (N_417,In_231,In_1493);
nor U418 (N_418,In_1726,In_1831);
nand U419 (N_419,In_16,In_1430);
and U420 (N_420,In_230,In_1526);
nand U421 (N_421,In_2237,In_1212);
or U422 (N_422,In_2991,In_73);
and U423 (N_423,In_1735,In_100);
and U424 (N_424,In_715,In_2183);
nand U425 (N_425,In_551,In_2816);
and U426 (N_426,In_128,In_1865);
or U427 (N_427,In_1154,In_659);
or U428 (N_428,In_2508,In_1514);
and U429 (N_429,In_2923,In_79);
and U430 (N_430,In_2493,In_139);
or U431 (N_431,In_976,In_436);
and U432 (N_432,In_1143,In_2704);
and U433 (N_433,In_89,In_2393);
nor U434 (N_434,In_2873,In_2685);
and U435 (N_435,In_990,In_2658);
and U436 (N_436,In_1592,In_705);
nor U437 (N_437,In_933,In_1322);
and U438 (N_438,In_2863,In_978);
or U439 (N_439,In_1189,In_2791);
nand U440 (N_440,In_2362,In_606);
nor U441 (N_441,In_1870,In_1722);
or U442 (N_442,In_2074,In_2314);
nor U443 (N_443,In_2652,In_774);
nand U444 (N_444,In_2498,In_1492);
nand U445 (N_445,In_2550,In_1543);
nor U446 (N_446,In_1976,In_2286);
nor U447 (N_447,In_1324,In_192);
nor U448 (N_448,In_1797,In_2605);
nand U449 (N_449,In_1012,In_320);
nand U450 (N_450,In_2269,In_1568);
and U451 (N_451,In_508,In_1944);
or U452 (N_452,In_1638,In_1426);
or U453 (N_453,In_1681,In_365);
and U454 (N_454,In_2919,In_1765);
and U455 (N_455,In_184,In_188);
nor U456 (N_456,In_664,In_652);
or U457 (N_457,In_2820,In_2617);
or U458 (N_458,In_449,In_1827);
and U459 (N_459,In_678,In_2387);
nand U460 (N_460,In_845,In_2486);
nand U461 (N_461,In_2119,In_378);
and U462 (N_462,In_552,In_1609);
and U463 (N_463,In_1991,In_247);
nor U464 (N_464,In_86,In_40);
nor U465 (N_465,In_1630,In_1131);
nand U466 (N_466,In_1,In_1050);
nor U467 (N_467,In_363,In_882);
nor U468 (N_468,In_1756,In_559);
or U469 (N_469,In_148,In_470);
nor U470 (N_470,In_164,In_1406);
or U471 (N_471,In_2885,In_2353);
nand U472 (N_472,In_2712,In_1040);
nor U473 (N_473,In_367,In_544);
or U474 (N_474,In_820,In_2141);
and U475 (N_475,In_1617,In_384);
or U476 (N_476,In_987,In_2869);
and U477 (N_477,In_194,In_1601);
or U478 (N_478,In_347,In_70);
and U479 (N_479,In_2172,In_693);
nor U480 (N_480,In_686,In_914);
nor U481 (N_481,In_45,In_2030);
nand U482 (N_482,In_1019,In_877);
and U483 (N_483,In_1241,In_146);
or U484 (N_484,In_2623,In_1142);
nand U485 (N_485,In_1480,In_1499);
nand U486 (N_486,In_775,In_2968);
and U487 (N_487,In_2289,In_66);
and U488 (N_488,In_2586,In_867);
or U489 (N_489,In_2965,In_1296);
nand U490 (N_490,In_1470,In_1926);
or U491 (N_491,In_1208,In_2365);
and U492 (N_492,In_1920,In_2669);
or U493 (N_493,In_2101,In_1825);
nor U494 (N_494,In_2216,In_277);
nor U495 (N_495,In_1794,In_2597);
or U496 (N_496,In_304,In_1041);
nand U497 (N_497,In_2137,In_1500);
nand U498 (N_498,In_2579,In_375);
or U499 (N_499,In_1251,In_2581);
xnor U500 (N_500,In_291,In_802);
nor U501 (N_501,In_604,In_754);
nor U502 (N_502,In_223,In_797);
or U503 (N_503,In_896,In_2446);
or U504 (N_504,In_2787,In_233);
and U505 (N_505,In_680,In_529);
or U506 (N_506,In_2202,In_2898);
nor U507 (N_507,In_533,In_591);
and U508 (N_508,In_1921,In_727);
nand U509 (N_509,In_2773,In_1668);
nor U510 (N_510,In_2276,In_1039);
or U511 (N_511,In_503,In_1646);
nor U512 (N_512,In_486,In_1096);
nor U513 (N_513,In_562,In_1713);
and U514 (N_514,In_2354,In_2638);
and U515 (N_515,In_2176,In_1723);
nand U516 (N_516,In_1810,In_1084);
nand U517 (N_517,In_994,In_2197);
nor U518 (N_518,In_460,In_2847);
and U519 (N_519,In_1228,In_2815);
or U520 (N_520,In_1843,In_738);
nand U521 (N_521,In_2794,In_145);
nor U522 (N_522,In_134,In_2343);
nor U523 (N_523,In_2021,In_2126);
or U524 (N_524,In_373,In_671);
nand U525 (N_525,In_2210,In_1659);
or U526 (N_526,In_766,In_585);
nor U527 (N_527,In_1219,In_1847);
or U528 (N_528,In_322,In_803);
nor U529 (N_529,In_1928,In_2901);
nor U530 (N_530,In_536,In_1357);
nor U531 (N_531,In_2502,In_956);
nor U532 (N_532,In_634,In_2171);
nor U533 (N_533,In_234,In_673);
nor U534 (N_534,In_432,In_2821);
or U535 (N_535,In_2386,In_1912);
or U536 (N_536,In_1375,In_1812);
nor U537 (N_537,In_415,In_2648);
or U538 (N_538,In_502,In_136);
nor U539 (N_539,In_2635,In_1116);
nand U540 (N_540,In_441,In_1712);
nor U541 (N_541,In_2214,In_2769);
xnor U542 (N_542,In_114,In_74);
nor U543 (N_543,In_2972,In_2596);
or U544 (N_544,In_582,In_52);
and U545 (N_545,In_1188,In_2594);
nand U546 (N_546,In_561,In_955);
or U547 (N_547,In_824,In_2291);
or U548 (N_548,In_2953,In_1158);
nand U549 (N_549,In_2982,In_237);
nand U550 (N_550,In_2934,In_288);
nor U551 (N_551,In_1932,In_1059);
nand U552 (N_552,In_152,In_1820);
nand U553 (N_553,In_403,In_2813);
xnor U554 (N_554,In_2720,In_1772);
nor U555 (N_555,In_1780,In_112);
and U556 (N_556,In_972,In_1018);
nand U557 (N_557,In_2029,In_2559);
and U558 (N_558,In_2413,In_144);
nand U559 (N_559,In_2839,In_102);
and U560 (N_560,In_2042,In_25);
and U561 (N_561,In_269,In_782);
nand U562 (N_562,In_1353,In_1505);
nand U563 (N_563,In_2339,In_1087);
and U564 (N_564,In_2388,In_149);
nor U565 (N_565,In_1498,In_2943);
or U566 (N_566,In_1523,In_2999);
and U567 (N_567,In_938,In_516);
or U568 (N_568,In_620,In_2391);
nand U569 (N_569,In_1340,In_1169);
and U570 (N_570,In_866,In_1640);
nor U571 (N_571,In_2679,In_2690);
and U572 (N_572,In_1745,In_2841);
or U573 (N_573,In_1078,In_912);
and U574 (N_574,In_1491,In_2114);
nand U575 (N_575,In_894,In_236);
and U576 (N_576,In_2139,In_1117);
or U577 (N_577,In_2469,In_1876);
and U578 (N_578,In_2312,In_1805);
nor U579 (N_579,In_124,In_801);
or U580 (N_580,In_259,In_1358);
and U581 (N_581,In_2344,In_2702);
or U582 (N_582,In_2037,In_1231);
and U583 (N_583,In_2959,In_2311);
and U584 (N_584,In_361,In_2755);
xnor U585 (N_585,In_1590,In_1743);
nor U586 (N_586,In_2628,In_1413);
and U587 (N_587,In_2464,In_814);
and U588 (N_588,In_2718,In_522);
nor U589 (N_589,In_885,In_1699);
nor U590 (N_590,In_1017,In_742);
or U591 (N_591,In_925,In_1412);
and U592 (N_592,In_2681,In_1677);
and U593 (N_593,In_870,In_1533);
and U594 (N_594,In_2073,In_455);
and U595 (N_595,In_658,In_1088);
and U596 (N_596,In_1520,In_289);
nor U597 (N_597,In_286,In_623);
or U598 (N_598,In_2892,In_2055);
nand U599 (N_599,In_2757,In_2540);
nor U600 (N_600,In_1693,In_1702);
and U601 (N_601,In_2854,In_706);
and U602 (N_602,In_2743,In_1390);
or U603 (N_603,In_2005,In_2068);
nor U604 (N_604,In_60,In_2911);
nor U605 (N_605,In_143,In_406);
or U606 (N_606,In_453,In_487);
nor U607 (N_607,In_2929,In_2545);
nand U608 (N_608,In_1269,In_2315);
or U609 (N_609,In_1815,In_609);
or U610 (N_610,In_1216,In_3);
nand U611 (N_611,In_1589,In_266);
and U612 (N_612,In_2744,In_849);
and U613 (N_613,In_2560,In_2133);
and U614 (N_614,In_2654,In_2115);
nor U615 (N_615,In_709,In_356);
nand U616 (N_616,In_926,In_1642);
or U617 (N_617,In_1739,In_1785);
nand U618 (N_618,In_722,In_1179);
nand U619 (N_619,In_816,In_1310);
and U620 (N_620,In_1982,In_2618);
and U621 (N_621,In_2085,In_475);
nor U622 (N_622,In_177,In_1984);
nand U623 (N_623,In_2677,In_1176);
xnor U624 (N_624,In_2667,In_2924);
nor U625 (N_625,In_892,In_1037);
nand U626 (N_626,In_2647,In_2888);
nor U627 (N_627,In_2043,In_2849);
nand U628 (N_628,In_1248,In_1538);
or U629 (N_629,In_1509,In_1558);
or U630 (N_630,In_213,In_2711);
nand U631 (N_631,In_967,In_391);
and U632 (N_632,In_1186,In_624);
nor U633 (N_633,In_1486,In_221);
or U634 (N_634,In_1955,In_307);
or U635 (N_635,In_32,In_1431);
nand U636 (N_636,In_581,In_1280);
nand U637 (N_637,In_1729,In_2956);
nor U638 (N_638,In_1900,In_1302);
and U639 (N_639,In_1146,In_2369);
and U640 (N_640,In_5,In_362);
or U641 (N_641,In_1286,In_1622);
nand U642 (N_642,In_1849,In_2432);
or U643 (N_643,In_1016,In_563);
or U644 (N_644,In_83,In_404);
nor U645 (N_645,In_202,In_1516);
and U646 (N_646,In_1660,In_2337);
nor U647 (N_647,In_832,In_541);
nand U648 (N_648,In_2317,In_1274);
nor U649 (N_649,In_2661,In_2422);
nor U650 (N_650,In_2439,In_1305);
or U651 (N_651,In_1163,In_2461);
and U652 (N_652,In_655,In_1884);
and U653 (N_653,In_764,In_2025);
or U654 (N_654,In_2032,In_344);
and U655 (N_655,In_2983,In_2827);
or U656 (N_656,In_439,In_9);
nor U657 (N_657,In_1326,In_2630);
and U658 (N_658,In_1894,In_1809);
or U659 (N_659,In_750,In_712);
nor U660 (N_660,In_2890,In_2664);
and U661 (N_661,In_239,In_412);
nor U662 (N_662,In_1676,In_989);
nor U663 (N_663,In_543,In_1898);
nand U664 (N_664,In_1437,In_2735);
nand U665 (N_665,In_590,In_2563);
nand U666 (N_666,In_887,In_720);
nor U667 (N_667,In_1199,In_631);
or U668 (N_668,In_2444,In_2608);
and U669 (N_669,In_2495,In_2031);
nor U670 (N_670,In_1654,In_2146);
nand U671 (N_671,In_1577,In_1690);
nor U672 (N_672,In_1398,In_442);
nor U673 (N_673,In_1330,In_62);
nor U674 (N_674,In_2342,In_1917);
or U675 (N_675,In_1950,In_1918);
nor U676 (N_676,In_90,In_2356);
nor U677 (N_677,In_2295,In_2851);
nor U678 (N_678,In_88,In_2009);
nand U679 (N_679,In_49,In_1675);
or U680 (N_680,In_1458,In_2551);
or U681 (N_681,In_1030,In_2590);
and U682 (N_682,In_2771,In_2240);
and U683 (N_683,In_1265,In_2799);
and U684 (N_684,In_2845,In_2107);
nor U685 (N_685,In_2201,In_821);
nand U686 (N_686,In_1385,In_179);
or U687 (N_687,In_2971,In_1056);
nand U688 (N_688,In_1618,In_2962);
or U689 (N_689,In_2098,In_2434);
or U690 (N_690,In_1679,In_2109);
and U691 (N_691,In_478,In_831);
and U692 (N_692,In_2305,In_2795);
nor U693 (N_693,In_2438,In_1776);
or U694 (N_694,In_358,In_511);
nor U695 (N_695,In_1471,In_1850);
nand U696 (N_696,In_399,In_1755);
nor U697 (N_697,In_2908,In_2411);
nor U698 (N_698,In_2719,In_848);
nand U699 (N_699,In_1071,In_1653);
or U700 (N_700,In_1877,In_168);
and U701 (N_701,In_2102,In_1525);
nand U702 (N_702,In_2687,In_335);
or U703 (N_703,In_232,In_642);
nor U704 (N_704,In_2261,In_46);
nor U705 (N_705,In_349,In_1121);
or U706 (N_706,In_2058,In_1560);
xnor U707 (N_707,In_1402,In_1790);
or U708 (N_708,In_1474,In_2700);
or U709 (N_709,In_2668,In_69);
xor U710 (N_710,In_2987,In_1111);
nor U711 (N_711,In_1861,In_662);
xor U712 (N_712,In_1536,In_2187);
nand U713 (N_713,In_2233,In_2721);
nor U714 (N_714,In_1282,In_1696);
nand U715 (N_715,In_731,In_723);
nand U716 (N_716,In_667,In_1695);
nand U717 (N_717,In_2951,In_795);
and U718 (N_718,In_873,In_2092);
nand U719 (N_719,In_2497,In_2195);
nor U720 (N_720,In_481,In_2213);
or U721 (N_721,In_2149,In_1572);
nor U722 (N_722,In_2973,In_1025);
nor U723 (N_723,In_218,In_1718);
nand U724 (N_724,In_1881,In_1806);
nand U725 (N_725,In_1902,In_1551);
nand U726 (N_726,In_711,In_2619);
and U727 (N_727,In_565,In_1673);
xor U728 (N_728,In_2255,In_0);
nor U729 (N_729,In_1692,In_2406);
and U730 (N_730,In_1429,In_751);
nor U731 (N_731,In_924,In_1683);
nand U732 (N_732,In_545,In_1064);
and U733 (N_733,In_1610,In_2856);
or U734 (N_734,In_1529,In_2734);
or U735 (N_735,In_2251,In_1503);
nor U736 (N_736,In_2876,In_1930);
or U737 (N_737,In_1631,In_645);
and U738 (N_738,In_2028,In_2064);
nor U739 (N_739,In_540,In_1076);
and U740 (N_740,In_900,In_2503);
or U741 (N_741,In_861,In_2454);
or U742 (N_742,In_98,In_669);
nor U743 (N_743,In_382,In_2212);
nand U744 (N_744,In_730,In_1370);
nor U745 (N_745,In_59,In_1010);
nor U746 (N_746,In_903,In_2512);
nand U747 (N_747,In_690,In_1771);
nand U748 (N_748,In_842,In_959);
nand U749 (N_749,In_1452,In_982);
nor U750 (N_750,In_1453,In_517);
or U751 (N_751,In_2610,In_2303);
or U752 (N_752,In_1669,In_1226);
or U753 (N_753,In_2466,In_419);
and U754 (N_754,In_2034,In_807);
and U755 (N_755,In_2252,In_2728);
xnor U756 (N_756,In_1113,In_121);
and U757 (N_757,In_1336,In_1393);
or U758 (N_758,In_2451,In_1270);
nand U759 (N_759,In_890,In_1172);
or U760 (N_760,In_653,In_2916);
nor U761 (N_761,In_2708,In_1952);
and U762 (N_762,In_2370,In_2404);
xor U763 (N_763,In_734,In_346);
nor U764 (N_764,In_1232,In_1367);
nor U765 (N_765,In_75,In_2850);
nor U766 (N_766,In_1027,In_2447);
or U767 (N_767,In_1178,In_2227);
and U768 (N_768,In_1475,In_397);
nor U769 (N_769,In_2090,In_1000);
and U770 (N_770,In_2472,In_1933);
nand U771 (N_771,In_1964,In_92);
or U772 (N_772,In_668,In_2766);
or U773 (N_773,In_881,In_2714);
and U774 (N_774,In_1317,In_1449);
or U775 (N_775,In_2653,In_806);
or U776 (N_776,In_1436,In_2225);
or U777 (N_777,In_336,In_2985);
nor U778 (N_778,In_2883,In_851);
nand U779 (N_779,In_869,In_334);
nand U780 (N_780,In_507,In_1339);
or U781 (N_781,In_2238,In_991);
or U782 (N_782,In_1544,In_1769);
or U783 (N_783,In_980,In_2487);
and U784 (N_784,In_2620,In_1857);
nor U785 (N_785,In_2767,In_1909);
nor U786 (N_786,In_1319,In_584);
nand U787 (N_787,In_501,In_856);
nor U788 (N_788,In_2615,In_1031);
or U789 (N_789,In_2128,In_769);
and U790 (N_790,In_2253,In_1714);
nor U791 (N_791,In_1986,In_2629);
nor U792 (N_792,In_1215,In_1709);
and U793 (N_793,In_1294,In_195);
nor U794 (N_794,In_596,In_535);
and U795 (N_795,In_1218,In_1753);
nor U796 (N_796,In_2796,In_2780);
xor U797 (N_797,In_527,In_2778);
nand U798 (N_798,In_1356,In_2724);
or U799 (N_799,In_1816,In_1401);
nand U800 (N_800,In_1147,In_745);
nand U801 (N_801,In_1002,In_394);
and U802 (N_802,In_2920,In_2583);
nor U803 (N_803,In_1126,In_2300);
nand U804 (N_804,In_386,In_308);
and U805 (N_805,In_212,In_612);
or U806 (N_806,In_462,In_899);
nor U807 (N_807,In_345,In_1077);
nand U808 (N_808,In_930,In_1775);
or U809 (N_809,In_1561,In_666);
and U810 (N_810,In_1312,In_492);
or U811 (N_811,In_2351,In_2684);
nor U812 (N_812,In_2864,In_1164);
nand U813 (N_813,In_917,In_2519);
nor U814 (N_814,In_2941,In_2232);
or U815 (N_815,In_241,In_1328);
nor U816 (N_816,In_2321,In_2651);
nor U817 (N_817,In_1046,In_2793);
nor U818 (N_818,In_96,In_2378);
nand U819 (N_819,In_6,In_376);
nor U820 (N_820,In_2774,In_1648);
nor U821 (N_821,In_1069,In_2553);
and U822 (N_822,In_672,In_736);
nand U823 (N_823,In_1663,In_1097);
nand U824 (N_824,In_916,In_557);
nand U825 (N_825,In_1817,In_771);
nand U826 (N_826,In_1862,In_988);
nor U827 (N_827,In_1846,In_2394);
nand U828 (N_828,In_2250,In_1853);
or U829 (N_829,In_2418,In_1522);
and U830 (N_830,In_1365,In_2083);
nor U831 (N_831,In_216,In_1913);
or U832 (N_832,In_2499,In_2080);
or U833 (N_833,In_753,In_1969);
or U834 (N_834,In_579,In_2011);
or U835 (N_835,In_408,In_872);
or U836 (N_836,In_2359,In_2598);
nand U837 (N_837,In_1929,In_898);
nand U838 (N_838,In_162,In_2164);
or U839 (N_839,In_2776,In_875);
or U840 (N_840,In_947,In_433);
nor U841 (N_841,In_1224,In_2416);
and U842 (N_842,In_1396,In_421);
nor U843 (N_843,In_374,In_526);
nor U844 (N_844,In_1960,In_2872);
or U845 (N_845,In_595,In_2436);
and U846 (N_846,In_830,In_1834);
nor U847 (N_847,In_1457,In_2144);
and U848 (N_848,In_1315,In_1229);
nor U849 (N_849,In_2650,In_2132);
or U850 (N_850,In_1606,In_732);
nand U851 (N_851,In_1276,In_1090);
nor U852 (N_852,In_968,In_405);
and U853 (N_853,In_1914,In_1091);
or U854 (N_854,In_985,In_513);
nor U855 (N_855,In_1127,In_1168);
nor U856 (N_856,In_610,In_1830);
nand U857 (N_857,In_402,In_2576);
or U858 (N_858,In_1194,In_1540);
and U859 (N_859,In_1852,In_1945);
nor U860 (N_860,In_1584,In_1537);
nand U861 (N_861,In_1337,In_2875);
or U862 (N_862,In_226,In_1444);
and U863 (N_863,In_1141,In_2186);
nor U864 (N_864,In_2614,In_2955);
nor U865 (N_865,In_1008,In_825);
xnor U866 (N_866,In_2100,In_2199);
and U867 (N_867,In_1751,In_2367);
nand U868 (N_868,In_203,In_1477);
or U869 (N_869,In_1386,In_2995);
and U870 (N_870,In_2996,In_2427);
nor U871 (N_871,In_1463,In_2582);
nor U872 (N_872,In_2001,In_1703);
or U873 (N_873,In_2296,In_951);
or U874 (N_874,In_2798,In_2636);
nor U875 (N_875,In_641,In_2364);
nand U876 (N_876,In_749,In_2937);
and U877 (N_877,In_986,In_325);
and U878 (N_878,In_725,In_137);
nor U879 (N_879,In_1106,In_321);
nor U880 (N_880,In_2450,In_2443);
and U881 (N_881,In_717,In_2298);
nor U882 (N_882,In_1983,In_1565);
and U883 (N_883,In_341,In_2167);
nand U884 (N_884,In_2529,In_2329);
and U885 (N_885,In_451,In_2002);
or U886 (N_886,In_2473,In_1363);
and U887 (N_887,In_756,In_2572);
and U888 (N_888,In_1748,In_438);
nand U889 (N_889,In_1271,In_490);
nor U890 (N_890,In_696,In_2368);
nand U891 (N_891,In_1757,In_2471);
nand U892 (N_892,In_1706,In_1185);
nand U893 (N_893,In_2834,In_2790);
and U894 (N_894,In_2327,In_172);
nand U895 (N_895,In_85,In_1562);
nand U896 (N_896,In_884,In_657);
or U897 (N_897,In_390,In_1911);
nand U898 (N_898,In_1156,In_780);
and U899 (N_899,In_2020,In_1114);
nor U900 (N_900,In_1464,In_2889);
and U901 (N_901,In_2392,In_1022);
nor U902 (N_902,In_2585,In_2797);
and U903 (N_903,In_793,In_1644);
nand U904 (N_904,In_1472,In_337);
nand U905 (N_905,In_714,In_2806);
and U906 (N_906,In_2417,In_874);
nor U907 (N_907,In_762,In_115);
nand U908 (N_908,In_333,In_457);
nand U909 (N_909,In_1478,In_2818);
or U910 (N_910,In_2981,In_523);
or U911 (N_911,In_721,In_768);
nand U912 (N_912,In_2893,In_1990);
or U913 (N_913,In_2108,In_2504);
or U914 (N_914,In_2247,In_2477);
nor U915 (N_915,In_1604,In_2836);
nor U916 (N_916,In_853,In_283);
or U917 (N_917,In_2830,In_1556);
nor U918 (N_918,In_965,In_835);
nor U919 (N_919,In_2753,In_1587);
nand U920 (N_920,In_2006,In_1626);
and U921 (N_921,In_1038,In_2558);
nor U922 (N_922,In_2867,In_1766);
or U923 (N_923,In_2866,In_2672);
and U924 (N_924,In_532,In_2082);
nor U925 (N_925,In_1740,In_1155);
or U926 (N_926,In_2245,In_1994);
nand U927 (N_927,In_2587,In_2729);
nand U928 (N_928,In_893,In_4);
and U929 (N_929,In_2103,In_210);
and U930 (N_930,In_614,In_2331);
and U931 (N_931,In_228,In_1072);
nand U932 (N_932,In_1506,In_1497);
or U933 (N_933,In_68,In_2606);
nand U934 (N_934,In_1233,In_573);
and U935 (N_935,In_1935,In_2536);
or U936 (N_936,In_1583,In_1736);
nand U937 (N_937,In_2829,In_1860);
and U938 (N_938,In_2235,In_65);
nor U939 (N_939,In_1094,In_2242);
nor U940 (N_940,In_2731,In_2086);
or U941 (N_941,In_1015,In_1469);
or U942 (N_942,In_1354,In_1255);
nand U943 (N_943,In_315,In_280);
nand U944 (N_944,In_1262,In_120);
xor U945 (N_945,In_785,In_2414);
nor U946 (N_946,In_150,In_1023);
nor U947 (N_947,In_2091,In_2196);
nor U948 (N_948,In_1079,In_2008);
nand U949 (N_949,In_586,In_2859);
and U950 (N_950,In_171,In_7);
and U951 (N_951,In_2877,In_977);
nor U952 (N_952,In_2642,In_2293);
and U953 (N_953,In_2831,In_1967);
nor U954 (N_954,In_2138,In_1416);
and U955 (N_955,In_456,In_2290);
nor U956 (N_956,In_1425,In_998);
or U957 (N_957,In_303,In_1287);
or U958 (N_958,In_2570,In_2948);
nand U959 (N_959,In_626,In_1267);
and U960 (N_960,In_1878,In_2150);
nor U961 (N_961,In_637,In_2510);
nand U962 (N_962,In_2506,In_2857);
and U963 (N_963,In_2173,In_1260);
nand U964 (N_964,In_23,In_476);
nor U965 (N_965,In_929,In_1842);
and U966 (N_966,In_450,In_2969);
or U967 (N_967,In_1099,In_156);
nand U968 (N_968,In_783,In_1530);
and U969 (N_969,In_2588,In_2067);
nand U970 (N_970,In_1586,In_2124);
and U971 (N_971,In_2355,In_908);
nor U972 (N_972,In_1685,In_1422);
and U973 (N_973,In_506,In_1671);
or U974 (N_974,In_1761,In_1235);
and U975 (N_975,In_1133,In_515);
and U976 (N_976,In_24,In_2382);
nand U977 (N_977,In_2759,In_1400);
nand U978 (N_978,In_2994,In_2441);
or U979 (N_979,In_2140,In_1517);
or U980 (N_980,In_2492,In_2390);
and U981 (N_981,In_2057,In_1836);
nand U982 (N_982,In_906,In_1803);
nor U983 (N_983,In_2268,In_1230);
nand U984 (N_984,In_1768,In_33);
nor U985 (N_985,In_791,In_2410);
nand U986 (N_986,In_1063,In_158);
nor U987 (N_987,In_812,In_1833);
and U988 (N_988,In_1054,In_809);
nand U989 (N_989,In_954,In_871);
xnor U990 (N_990,In_477,In_2546);
nor U991 (N_991,In_1303,In_187);
nand U992 (N_992,In_426,In_1534);
and U993 (N_993,In_2409,In_2346);
nand U994 (N_994,In_2266,In_2309);
nor U995 (N_995,In_630,In_1783);
nor U996 (N_996,In_31,In_1115);
and U997 (N_997,In_973,In_1362);
or U998 (N_998,In_636,In_2958);
nand U999 (N_999,In_2480,In_411);
nor U1000 (N_1000,In_2660,In_2014);
nor U1001 (N_1001,In_1826,In_1970);
and U1002 (N_1002,In_1838,In_2870);
nor U1003 (N_1003,In_1882,In_360);
or U1004 (N_1004,In_2500,In_1864);
and U1005 (N_1005,In_1987,In_1074);
nor U1006 (N_1006,In_249,In_1465);
and U1007 (N_1007,In_1432,In_2175);
and U1008 (N_1008,In_2833,In_1807);
or U1009 (N_1009,In_123,In_2297);
nand U1010 (N_1010,In_865,In_2077);
and U1011 (N_1011,In_1554,In_1829);
nor U1012 (N_1012,In_2739,In_1417);
and U1013 (N_1013,In_1710,In_2040);
nor U1014 (N_1014,In_2578,In_2523);
nand U1015 (N_1015,In_2907,In_1956);
nand U1016 (N_1016,In_2013,In_550);
nor U1017 (N_1017,In_116,In_1580);
nor U1018 (N_1018,In_1166,In_2481);
nor U1019 (N_1019,In_1614,In_1376);
nand U1020 (N_1020,In_1440,In_2977);
nand U1021 (N_1021,In_424,In_996);
or U1022 (N_1022,In_2786,In_2641);
and U1023 (N_1023,In_1243,In_51);
nor U1024 (N_1024,In_1223,In_2603);
or U1025 (N_1025,In_2112,In_1645);
or U1026 (N_1026,In_1202,In_1314);
and U1027 (N_1027,In_2288,In_905);
and U1028 (N_1028,In_2980,In_135);
or U1029 (N_1029,In_1936,In_485);
or U1030 (N_1030,In_141,In_879);
or U1031 (N_1031,In_2960,In_13);
or U1032 (N_1032,In_1132,In_1150);
and U1033 (N_1033,In_1504,In_2548);
nand U1034 (N_1034,In_580,In_1557);
and U1035 (N_1035,In_1331,In_525);
and U1036 (N_1036,In_2095,In_2577);
nor U1037 (N_1037,In_186,In_2230);
and U1038 (N_1038,In_521,In_253);
or U1039 (N_1039,In_211,In_257);
or U1040 (N_1040,In_2542,In_1275);
or U1041 (N_1041,In_1167,In_1268);
nand U1042 (N_1042,In_1129,In_293);
or U1043 (N_1043,In_2624,In_1007);
nor U1044 (N_1044,In_862,In_1144);
or U1045 (N_1045,In_2142,In_2511);
nor U1046 (N_1046,In_183,In_2189);
nor U1047 (N_1047,In_504,In_904);
and U1048 (N_1048,In_910,In_2532);
nand U1049 (N_1049,In_1043,In_1715);
or U1050 (N_1050,In_2328,In_1473);
or U1051 (N_1051,In_2239,In_1483);
or U1052 (N_1052,In_2217,In_2915);
nor U1053 (N_1053,In_246,In_2012);
and U1054 (N_1054,In_1307,In_255);
nor U1055 (N_1055,In_1191,In_1066);
or U1056 (N_1056,In_2513,In_261);
or U1057 (N_1057,In_151,In_294);
or U1058 (N_1058,In_499,In_2234);
and U1059 (N_1059,In_2803,In_282);
nor U1060 (N_1060,In_1858,In_743);
nor U1061 (N_1061,In_2279,In_251);
and U1062 (N_1062,In_1995,In_497);
nor U1063 (N_1063,In_281,In_2219);
and U1064 (N_1064,In_1818,In_2078);
or U1065 (N_1065,In_2038,In_1256);
nand U1066 (N_1066,In_1875,In_1395);
nand U1067 (N_1067,In_330,In_1716);
nand U1068 (N_1068,In_627,In_752);
nor U1069 (N_1069,In_1868,In_2458);
nor U1070 (N_1070,In_2612,In_1837);
nand U1071 (N_1071,In_2840,In_2318);
nand U1072 (N_1072,In_43,In_2741);
or U1073 (N_1073,In_1596,In_1866);
nor U1074 (N_1074,In_2323,In_539);
nor U1075 (N_1075,In_427,In_55);
or U1076 (N_1076,In_1502,In_2079);
nor U1077 (N_1077,In_804,In_2437);
nand U1078 (N_1078,In_767,In_1343);
nor U1079 (N_1079,In_270,In_2940);
or U1080 (N_1080,In_103,In_34);
or U1081 (N_1081,In_1643,In_944);
nand U1082 (N_1082,In_2292,In_2063);
nand U1083 (N_1083,In_2193,In_2942);
and U1084 (N_1084,In_1182,In_2932);
nor U1085 (N_1085,In_2802,In_2894);
and U1086 (N_1086,In_2229,In_739);
nand U1087 (N_1087,In_1494,In_1062);
or U1088 (N_1088,In_2271,In_2571);
nor U1089 (N_1089,In_1211,In_765);
or U1090 (N_1090,In_142,In_2903);
and U1091 (N_1091,In_2779,In_1535);
or U1092 (N_1092,In_676,In_773);
and U1093 (N_1093,In_84,In_306);
and U1094 (N_1094,In_1652,In_2084);
nand U1095 (N_1095,In_593,In_577);
or U1096 (N_1096,In_1571,In_2385);
and U1097 (N_1097,In_928,In_87);
or U1098 (N_1098,In_1119,In_787);
or U1099 (N_1099,In_252,In_2004);
and U1100 (N_1100,In_2015,In_328);
or U1101 (N_1101,In_1399,In_2745);
nand U1102 (N_1102,In_2374,In_287);
xor U1103 (N_1103,In_1989,In_140);
nand U1104 (N_1104,In_1819,In_1217);
nor U1105 (N_1105,In_2017,In_93);
nor U1106 (N_1106,In_2460,In_47);
nor U1107 (N_1107,In_2075,In_314);
nor U1108 (N_1108,In_1291,In_370);
and U1109 (N_1109,In_1575,In_1384);
nand U1110 (N_1110,In_2148,In_778);
nand U1111 (N_1111,In_2198,In_1427);
nor U1112 (N_1112,In_1355,In_2891);
and U1113 (N_1113,In_1379,In_1333);
or U1114 (N_1114,In_2007,In_353);
nor U1115 (N_1115,In_2333,In_846);
and U1116 (N_1116,In_29,In_1203);
nand U1117 (N_1117,In_1068,In_2478);
nand U1118 (N_1118,In_2946,In_209);
or U1119 (N_1119,In_482,In_2179);
nand U1120 (N_1120,In_1081,In_2659);
or U1121 (N_1121,In_1374,In_578);
and U1122 (N_1122,In_675,In_1198);
or U1123 (N_1123,In_2104,In_2961);
nand U1124 (N_1124,In_2675,In_1521);
and U1125 (N_1125,In_1196,In_1758);
and U1126 (N_1126,In_735,In_817);
nand U1127 (N_1127,In_2231,In_2424);
or U1128 (N_1128,In_1157,In_1383);
nand U1129 (N_1129,In_1588,In_2134);
or U1130 (N_1130,In_298,In_2270);
nand U1131 (N_1131,In_2453,In_410);
or U1132 (N_1132,In_2380,In_1737);
and U1133 (N_1133,In_2505,In_1802);
and U1134 (N_1134,In_2678,In_1943);
nor U1135 (N_1135,In_1661,In_1428);
nand U1136 (N_1136,In_1941,In_665);
nand U1137 (N_1137,In_431,In_423);
or U1138 (N_1138,In_2089,In_635);
and U1139 (N_1139,In_1484,In_1777);
nor U1140 (N_1140,In_174,In_1152);
and U1141 (N_1141,In_2979,In_868);
and U1142 (N_1142,In_467,In_828);
nor U1143 (N_1143,In_2544,In_235);
or U1144 (N_1144,In_2763,In_1550);
nand U1145 (N_1145,In_494,In_1700);
and U1146 (N_1146,In_327,In_10);
nand U1147 (N_1147,In_1424,In_181);
nor U1148 (N_1148,In_1633,In_21);
nor U1149 (N_1149,In_2947,In_2689);
and U1150 (N_1150,In_1651,In_2048);
or U1151 (N_1151,In_724,In_1961);
nor U1152 (N_1152,In_1593,In_50);
or U1153 (N_1153,In_1137,In_1468);
nor U1154 (N_1154,In_385,In_64);
or U1155 (N_1155,In_446,In_1341);
and U1156 (N_1156,In_227,In_2970);
or U1157 (N_1157,In_2902,In_1764);
nor U1158 (N_1158,In_747,In_570);
or U1159 (N_1159,In_1998,In_1828);
or U1160 (N_1160,In_2430,In_2822);
or U1161 (N_1161,In_2593,In_2649);
nor U1162 (N_1162,In_2555,In_927);
nand U1163 (N_1163,In_2113,In_553);
and U1164 (N_1164,In_413,In_469);
or U1165 (N_1165,In_2933,In_1637);
nor U1166 (N_1166,In_27,In_2278);
and U1167 (N_1167,In_1136,In_2396);
nand U1168 (N_1168,In_354,In_639);
nor U1169 (N_1169,In_1045,In_479);
or U1170 (N_1170,In_1931,In_2990);
or U1171 (N_1171,In_1047,In_1277);
or U1172 (N_1172,In_776,In_2254);
nor U1173 (N_1173,In_1542,In_243);
and U1174 (N_1174,In_2087,In_1871);
nor U1175 (N_1175,In_173,In_133);
or U1176 (N_1176,In_389,In_248);
and U1177 (N_1177,In_2792,In_1662);
nor U1178 (N_1178,In_2507,In_1246);
nor U1179 (N_1179,In_290,In_414);
or U1180 (N_1180,In_1352,In_2602);
nand U1181 (N_1181,In_1380,In_2639);
or U1182 (N_1182,In_1555,In_2156);
and U1183 (N_1183,In_2622,In_1065);
or U1184 (N_1184,In_1446,In_1415);
nor U1185 (N_1185,In_1796,In_920);
nor U1186 (N_1186,In_204,In_2099);
and U1187 (N_1187,In_1778,In_726);
and U1188 (N_1188,In_547,In_1093);
and U1189 (N_1189,In_505,In_1441);
and U1190 (N_1190,In_2754,In_1173);
nand U1191 (N_1191,In_728,In_1657);
nor U1192 (N_1192,In_1595,In_1100);
nor U1193 (N_1193,In_2052,In_1184);
nor U1194 (N_1194,In_14,In_1895);
nand U1195 (N_1195,In_1904,In_592);
nor U1196 (N_1196,In_1014,In_2801);
and U1197 (N_1197,In_2913,In_1299);
and U1198 (N_1198,In_2673,In_1906);
nand U1199 (N_1199,In_909,In_1403);
and U1200 (N_1200,In_2474,In_274);
and U1201 (N_1201,In_530,In_473);
nor U1202 (N_1202,In_1456,In_2993);
or U1203 (N_1203,In_1694,In_823);
and U1204 (N_1204,In_1942,In_1377);
or U1205 (N_1205,In_1075,In_937);
or U1206 (N_1206,In_1974,In_855);
or U1207 (N_1207,In_1612,In_2717);
xor U1208 (N_1208,In_2804,In_2828);
or U1209 (N_1209,In_1686,In_827);
nor U1210 (N_1210,In_429,In_1289);
nand U1211 (N_1211,In_1253,In_995);
nand U1212 (N_1212,In_1704,In_1620);
and U1213 (N_1213,In_1655,In_571);
and U1214 (N_1214,In_647,In_601);
nor U1215 (N_1215,In_953,In_2657);
or U1216 (N_1216,In_2177,In_2927);
or U1217 (N_1217,In_1180,In_2207);
or U1218 (N_1218,In_2878,In_465);
or U1219 (N_1219,In_2662,In_1859);
and U1220 (N_1220,In_1874,In_1207);
or U1221 (N_1221,In_1634,In_555);
nor U1222 (N_1222,In_331,In_1306);
nand U1223 (N_1223,In_2307,In_393);
and U1224 (N_1224,In_383,In_496);
or U1225 (N_1225,In_1689,In_1856);
and U1226 (N_1226,In_2917,In_169);
and U1227 (N_1227,In_1300,In_1236);
or U1228 (N_1228,In_2118,In_1787);
nand U1229 (N_1229,In_1409,In_238);
and U1230 (N_1230,In_2452,In_2626);
nor U1231 (N_1231,In_113,In_2347);
xor U1232 (N_1232,In_2088,In_1264);
nand U1233 (N_1233,In_2153,In_1602);
nor U1234 (N_1234,In_2567,In_1447);
nor U1235 (N_1235,In_1730,In_554);
nor U1236 (N_1236,In_922,In_1327);
or U1237 (N_1237,In_757,In_2725);
or U1238 (N_1238,In_2168,In_1149);
or U1239 (N_1239,In_1927,In_837);
nand U1240 (N_1240,In_2143,In_111);
nor U1241 (N_1241,In_833,In_1697);
and U1242 (N_1242,In_983,In_2554);
or U1243 (N_1243,In_2490,In_2223);
nand U1244 (N_1244,In_2056,In_245);
and U1245 (N_1245,In_78,In_338);
and U1246 (N_1246,In_138,In_1774);
and U1247 (N_1247,In_948,In_2281);
nor U1248 (N_1248,In_1767,In_364);
and U1249 (N_1249,In_1724,In_1647);
nor U1250 (N_1250,In_1527,In_993);
and U1251 (N_1251,In_654,In_2018);
and U1252 (N_1252,In_1957,In_42);
and U1253 (N_1253,In_1123,In_1348);
nor U1254 (N_1254,In_568,In_1210);
or U1255 (N_1255,In_677,In_2158);
and U1256 (N_1256,In_1420,In_2691);
nor U1257 (N_1257,In_1329,In_810);
and U1258 (N_1258,In_537,In_2050);
nand U1259 (N_1259,In_1938,In_788);
or U1260 (N_1260,In_2703,In_2313);
or U1261 (N_1261,In_420,In_1118);
or U1262 (N_1262,In_1507,In_1563);
or U1263 (N_1263,In_1281,In_1318);
nor U1264 (N_1264,In_2758,In_118);
nor U1265 (N_1265,In_224,In_1680);
nor U1266 (N_1266,In_1641,In_1999);
or U1267 (N_1267,In_2061,In_1910);
and U1268 (N_1268,In_1313,In_1247);
or U1269 (N_1269,In_1405,In_2592);
xnor U1270 (N_1270,In_607,In_2241);
or U1271 (N_1271,In_472,In_1576);
and U1272 (N_1272,In_1174,In_1067);
or U1273 (N_1273,In_2897,In_2926);
nand U1274 (N_1274,In_2407,In_683);
and U1275 (N_1275,In_2964,In_1404);
or U1276 (N_1276,In_2211,In_2096);
and U1277 (N_1277,In_2054,In_2843);
nor U1278 (N_1278,In_2549,In_2070);
nor U1279 (N_1279,In_534,In_2024);
and U1280 (N_1280,In_2749,In_931);
and U1281 (N_1281,In_2160,In_418);
and U1282 (N_1282,In_1181,In_847);
and U1283 (N_1283,In_2304,In_1225);
and U1284 (N_1284,In_2561,In_2805);
or U1285 (N_1285,In_1741,In_1053);
and U1286 (N_1286,In_2033,In_2420);
nor U1287 (N_1287,In_2984,In_1658);
or U1288 (N_1288,In_2706,In_2401);
and U1289 (N_1289,In_1049,In_981);
or U1290 (N_1290,In_2442,In_2110);
and U1291 (N_1291,In_891,In_1779);
and U1292 (N_1292,In_44,In_2595);
or U1293 (N_1293,In_2954,In_2978);
and U1294 (N_1294,In_1345,In_2494);
and U1295 (N_1295,In_2556,In_1977);
nor U1296 (N_1296,In_2398,In_2742);
nand U1297 (N_1297,In_2945,In_2459);
nor U1298 (N_1298,In_1382,In_2191);
nand U1299 (N_1299,In_1410,In_2564);
or U1300 (N_1300,In_1140,In_858);
or U1301 (N_1301,In_963,In_295);
nand U1302 (N_1302,In_256,In_126);
nand U1303 (N_1303,In_681,In_2868);
nor U1304 (N_1304,In_689,In_2435);
and U1305 (N_1305,In_199,In_1177);
and U1306 (N_1306,In_790,In_2525);
or U1307 (N_1307,In_2874,In_1261);
nor U1308 (N_1308,In_2967,In_2777);
or U1309 (N_1309,In_1896,In_2533);
nor U1310 (N_1310,In_2569,In_2206);
nand U1311 (N_1311,In_2844,In_692);
nand U1312 (N_1312,In_262,In_1024);
and U1313 (N_1313,In_2264,In_1082);
nor U1314 (N_1314,In_300,In_2429);
nand U1315 (N_1315,In_2000,In_1285);
and U1316 (N_1316,In_1781,In_488);
nand U1317 (N_1317,In_72,In_1600);
nor U1318 (N_1318,In_1033,In_317);
and U1319 (N_1319,In_719,In_663);
or U1320 (N_1320,In_608,In_30);
and U1321 (N_1321,In_379,In_1721);
and U1322 (N_1322,In_19,In_622);
nand U1323 (N_1323,In_2747,In_1629);
and U1324 (N_1324,In_1855,In_53);
nor U1325 (N_1325,In_594,In_2325);
or U1326 (N_1326,In_2861,In_1055);
nor U1327 (N_1327,In_2812,In_2918);
nor U1328 (N_1328,In_2445,In_2433);
and U1329 (N_1329,In_2543,In_1421);
or U1330 (N_1330,In_2053,In_196);
nand U1331 (N_1331,In_2810,In_2426);
and U1332 (N_1332,In_2676,In_999);
or U1333 (N_1333,In_1183,In_1605);
nand U1334 (N_1334,In_178,In_409);
and U1335 (N_1335,In_911,In_2887);
and U1336 (N_1336,In_2848,In_1165);
nor U1337 (N_1337,In_1145,In_1814);
nand U1338 (N_1338,In_1621,In_2846);
nor U1339 (N_1339,In_1244,In_1518);
and U1340 (N_1340,In_1892,In_1476);
nor U1341 (N_1341,In_2457,In_1897);
and U1342 (N_1342,In_1619,In_1501);
nor U1343 (N_1343,In_1451,In_1057);
nor U1344 (N_1344,In_1549,In_1320);
or U1345 (N_1345,In_538,In_1171);
nor U1346 (N_1346,In_278,In_2381);
or U1347 (N_1347,In_759,In_1979);
or U1348 (N_1348,In_205,In_387);
nand U1349 (N_1349,In_185,In_1581);
or U1350 (N_1350,In_567,In_2047);
nor U1351 (N_1351,In_271,In_166);
and U1352 (N_1352,In_548,In_1786);
nand U1353 (N_1353,In_273,In_549);
nor U1354 (N_1354,In_2674,In_1963);
nor U1355 (N_1355,In_1548,In_265);
nand U1356 (N_1356,In_2489,In_119);
or U1357 (N_1357,In_2862,In_1762);
nand U1358 (N_1358,In_332,In_1083);
and U1359 (N_1359,In_1213,In_1487);
nor U1360 (N_1360,In_401,In_718);
nor U1361 (N_1361,In_1411,In_1373);
nor U1362 (N_1362,In_613,In_2750);
nand U1363 (N_1363,In_2509,In_2324);
or U1364 (N_1364,In_250,In_2531);
nand U1365 (N_1365,In_1234,In_2950);
nor U1366 (N_1366,In_621,In_326);
nor U1367 (N_1367,In_946,In_569);
and U1368 (N_1368,In_2016,In_792);
or U1369 (N_1369,In_1749,In_1759);
and U1370 (N_1370,In_2957,In_1130);
or U1371 (N_1371,In_942,In_2373);
or U1372 (N_1372,In_1632,In_716);
nor U1373 (N_1373,In_2568,In_1845);
nand U1374 (N_1374,In_1013,In_297);
nor U1375 (N_1375,In_99,In_863);
nand U1376 (N_1376,In_1257,In_2727);
nand U1377 (N_1377,In_2807,In_1708);
or U1378 (N_1378,In_1691,In_1389);
and U1379 (N_1379,In_1105,In_2683);
nor U1380 (N_1380,In_1905,In_1058);
nor U1381 (N_1381,In_2611,In_2334);
and U1382 (N_1382,In_1539,In_1495);
nor U1383 (N_1383,In_2041,In_302);
and U1384 (N_1384,In_2182,In_2131);
nor U1385 (N_1385,In_740,In_2360);
or U1386 (N_1386,In_312,In_702);
nand U1387 (N_1387,In_1532,In_153);
or U1388 (N_1388,In_2781,In_2468);
and U1389 (N_1389,In_1279,In_1513);
or U1390 (N_1390,In_2931,In_2366);
and U1391 (N_1391,In_2485,In_1485);
or U1392 (N_1392,In_1784,In_2997);
nor U1393 (N_1393,In_129,In_1309);
nand U1394 (N_1394,In_2036,In_1488);
and U1395 (N_1395,In_770,In_1460);
and U1396 (N_1396,In_1738,In_1973);
or U1397 (N_1397,In_299,In_514);
nor U1398 (N_1398,In_2939,In_921);
nor U1399 (N_1399,In_815,In_901);
nor U1400 (N_1400,In_772,In_1206);
and U1401 (N_1401,In_1823,In_1242);
nor U1402 (N_1402,In_380,In_897);
nand U1403 (N_1403,In_2974,In_1195);
and U1404 (N_1404,In_26,In_2405);
nor U1405 (N_1405,In_1407,In_430);
nor U1406 (N_1406,In_826,In_777);
nor U1407 (N_1407,In_1628,In_8);
or U1408 (N_1408,In_1360,In_2145);
nor U1409 (N_1409,In_799,In_638);
nand U1410 (N_1410,In_984,In_323);
and U1411 (N_1411,In_2988,In_1564);
nand U1412 (N_1412,In_2809,In_107);
and U1413 (N_1413,In_932,In_1608);
or U1414 (N_1414,In_1705,In_2736);
and U1415 (N_1415,In_1011,In_1664);
and U1416 (N_1416,In_63,In_352);
and U1417 (N_1417,In_860,In_2415);
or U1418 (N_1418,In_674,In_2607);
nor U1419 (N_1419,In_558,In_839);
and U1420 (N_1420,In_276,In_1899);
nand U1421 (N_1421,In_458,In_1656);
nand U1422 (N_1422,In_2162,In_2428);
nor U1423 (N_1423,In_1635,In_1744);
nand U1424 (N_1424,In_805,In_970);
nor U1425 (N_1425,In_1221,In_1971);
nand U1426 (N_1426,In_2332,In_1887);
or U1427 (N_1427,In_2330,In_2808);
and U1428 (N_1428,In_1578,In_572);
nor U1429 (N_1429,In_589,In_603);
and U1430 (N_1430,In_1298,In_366);
nand U1431 (N_1431,In_369,In_2178);
nor U1432 (N_1432,In_2236,In_574);
and U1433 (N_1433,In_343,In_798);
xnor U1434 (N_1434,In_2403,In_1968);
or U1435 (N_1435,In_611,In_1443);
nor U1436 (N_1436,In_381,In_2699);
nand U1437 (N_1437,In_1455,In_1435);
nand U1438 (N_1438,In_61,In_2722);
nand U1439 (N_1439,In_2573,In_2185);
nor U1440 (N_1440,In_1616,In_2475);
and U1441 (N_1441,In_1325,In_2218);
nor U1442 (N_1442,In_1687,In_748);
nand U1443 (N_1443,In_1220,In_2180);
nor U1444 (N_1444,In_1813,In_1531);
nand U1445 (N_1445,In_695,In_1948);
nor U1446 (N_1446,In_2379,In_377);
or U1447 (N_1447,In_1788,In_495);
nor U1448 (N_1448,In_1720,In_95);
nand U1449 (N_1449,In_1599,In_2656);
nor U1450 (N_1450,In_1965,In_147);
nor U1451 (N_1451,In_1190,In_691);
nand U1452 (N_1452,In_1461,In_700);
or U1453 (N_1453,In_682,In_786);
nand U1454 (N_1454,In_1883,In_193);
nor U1455 (N_1455,In_2765,In_1344);
or U1456 (N_1456,In_200,In_2059);
nor U1457 (N_1457,In_510,In_108);
and U1458 (N_1458,In_2408,In_452);
or U1459 (N_1459,In_157,In_2698);
nor U1460 (N_1460,In_2188,In_850);
nand U1461 (N_1461,In_2928,In_2308);
nand U1462 (N_1462,In_122,In_1980);
or U1463 (N_1463,In_48,In_1209);
and U1464 (N_1464,In_2376,In_131);
or U1465 (N_1465,In_688,In_267);
or U1466 (N_1466,In_945,In_260);
nand U1467 (N_1467,In_165,In_2081);
nor U1468 (N_1468,In_958,In_1835);
nor U1469 (N_1469,In_2732,In_106);
and U1470 (N_1470,In_489,In_1200);
nand U1471 (N_1471,In_2097,In_2301);
nor U1472 (N_1472,In_2692,In_39);
xnor U1473 (N_1473,In_2905,In_2470);
and U1474 (N_1474,In_1872,In_2035);
and U1475 (N_1475,In_687,In_1627);
or U1476 (N_1476,In_1135,In_1086);
and U1477 (N_1477,In_2071,In_1295);
and U1478 (N_1478,In_1273,In_1515);
nor U1479 (N_1479,In_316,In_1009);
xnor U1480 (N_1480,In_1901,In_2775);
nand U1481 (N_1481,In_632,In_1278);
or U1482 (N_1482,In_1408,In_2375);
and U1483 (N_1483,In_1042,In_940);
and U1484 (N_1484,In_130,In_2051);
and U1485 (N_1485,In_1615,In_400);
nor U1486 (N_1486,In_2737,In_2130);
or U1487 (N_1487,In_372,In_2127);
nor U1488 (N_1488,In_1085,In_1193);
nand U1489 (N_1489,In_2921,In_841);
and U1490 (N_1490,In_2259,In_913);
and U1491 (N_1491,In_888,In_1482);
nand U1492 (N_1492,In_598,In_2476);
nand U1493 (N_1493,In_1423,In_1496);
or U1494 (N_1494,In_1051,In_2246);
nand U1495 (N_1495,In_1854,In_2837);
and U1496 (N_1496,In_2871,In_2220);
xor U1497 (N_1497,In_445,In_2256);
nand U1498 (N_1498,In_1290,In_1103);
and U1499 (N_1499,In_461,In_1727);
or U1500 (N_1500,In_532,In_603);
nor U1501 (N_1501,In_1168,In_189);
nand U1502 (N_1502,In_662,In_54);
and U1503 (N_1503,In_425,In_2302);
or U1504 (N_1504,In_786,In_2040);
nor U1505 (N_1505,In_980,In_2630);
nand U1506 (N_1506,In_1100,In_2248);
and U1507 (N_1507,In_2921,In_2874);
or U1508 (N_1508,In_230,In_2470);
or U1509 (N_1509,In_2166,In_738);
xor U1510 (N_1510,In_2913,In_839);
and U1511 (N_1511,In_1297,In_1685);
nor U1512 (N_1512,In_1724,In_1422);
nand U1513 (N_1513,In_2843,In_998);
nand U1514 (N_1514,In_2855,In_1655);
nand U1515 (N_1515,In_58,In_397);
or U1516 (N_1516,In_755,In_1137);
nand U1517 (N_1517,In_997,In_1650);
xor U1518 (N_1518,In_1115,In_1918);
nand U1519 (N_1519,In_1420,In_2968);
and U1520 (N_1520,In_2145,In_1794);
nor U1521 (N_1521,In_1888,In_1986);
and U1522 (N_1522,In_1328,In_2186);
nand U1523 (N_1523,In_1082,In_662);
and U1524 (N_1524,In_2056,In_1595);
nand U1525 (N_1525,In_702,In_223);
or U1526 (N_1526,In_2224,In_567);
nand U1527 (N_1527,In_2127,In_2536);
nor U1528 (N_1528,In_371,In_716);
nand U1529 (N_1529,In_1155,In_1455);
and U1530 (N_1530,In_984,In_1300);
nor U1531 (N_1531,In_2271,In_2821);
nand U1532 (N_1532,In_2523,In_45);
nor U1533 (N_1533,In_2534,In_211);
nand U1534 (N_1534,In_2784,In_1993);
nand U1535 (N_1535,In_2277,In_825);
nor U1536 (N_1536,In_1012,In_61);
or U1537 (N_1537,In_30,In_1496);
nand U1538 (N_1538,In_2445,In_2262);
nor U1539 (N_1539,In_999,In_2277);
nand U1540 (N_1540,In_613,In_1957);
nand U1541 (N_1541,In_629,In_1689);
and U1542 (N_1542,In_2513,In_2027);
and U1543 (N_1543,In_1049,In_747);
nor U1544 (N_1544,In_2195,In_1301);
nor U1545 (N_1545,In_2004,In_1743);
nand U1546 (N_1546,In_2299,In_1137);
nor U1547 (N_1547,In_2271,In_766);
nor U1548 (N_1548,In_16,In_2856);
or U1549 (N_1549,In_1692,In_2156);
or U1550 (N_1550,In_2302,In_898);
nand U1551 (N_1551,In_1742,In_1463);
or U1552 (N_1552,In_619,In_2049);
and U1553 (N_1553,In_2282,In_1266);
or U1554 (N_1554,In_608,In_496);
and U1555 (N_1555,In_2911,In_289);
and U1556 (N_1556,In_2921,In_1842);
nor U1557 (N_1557,In_477,In_1746);
nand U1558 (N_1558,In_2636,In_139);
or U1559 (N_1559,In_2287,In_618);
nor U1560 (N_1560,In_2880,In_2811);
nor U1561 (N_1561,In_832,In_422);
nand U1562 (N_1562,In_411,In_2306);
nor U1563 (N_1563,In_332,In_2386);
nor U1564 (N_1564,In_37,In_1569);
nor U1565 (N_1565,In_997,In_2199);
nor U1566 (N_1566,In_624,In_2591);
nand U1567 (N_1567,In_89,In_1181);
or U1568 (N_1568,In_2467,In_2100);
nand U1569 (N_1569,In_1332,In_1751);
nand U1570 (N_1570,In_2159,In_459);
nand U1571 (N_1571,In_2608,In_1249);
and U1572 (N_1572,In_732,In_150);
and U1573 (N_1573,In_1678,In_2513);
and U1574 (N_1574,In_2079,In_2737);
nand U1575 (N_1575,In_561,In_216);
or U1576 (N_1576,In_847,In_2312);
and U1577 (N_1577,In_2279,In_157);
nor U1578 (N_1578,In_647,In_162);
nand U1579 (N_1579,In_121,In_1094);
or U1580 (N_1580,In_2423,In_101);
nor U1581 (N_1581,In_984,In_2566);
or U1582 (N_1582,In_2823,In_1441);
nor U1583 (N_1583,In_1252,In_1545);
nor U1584 (N_1584,In_1837,In_1842);
nor U1585 (N_1585,In_157,In_1774);
and U1586 (N_1586,In_92,In_2496);
nor U1587 (N_1587,In_2346,In_347);
or U1588 (N_1588,In_1273,In_2787);
nand U1589 (N_1589,In_2831,In_740);
and U1590 (N_1590,In_2159,In_408);
or U1591 (N_1591,In_2601,In_1549);
nand U1592 (N_1592,In_2420,In_2310);
nor U1593 (N_1593,In_1141,In_1717);
or U1594 (N_1594,In_258,In_2928);
and U1595 (N_1595,In_1407,In_2793);
or U1596 (N_1596,In_2894,In_517);
or U1597 (N_1597,In_1145,In_2280);
nor U1598 (N_1598,In_658,In_2082);
and U1599 (N_1599,In_1164,In_1664);
nor U1600 (N_1600,In_2518,In_1600);
or U1601 (N_1601,In_1591,In_359);
and U1602 (N_1602,In_1017,In_2254);
nor U1603 (N_1603,In_1130,In_1371);
and U1604 (N_1604,In_826,In_1498);
or U1605 (N_1605,In_1727,In_870);
nor U1606 (N_1606,In_2957,In_1580);
nor U1607 (N_1607,In_1364,In_517);
nand U1608 (N_1608,In_1784,In_2261);
and U1609 (N_1609,In_2836,In_1928);
nor U1610 (N_1610,In_2844,In_5);
or U1611 (N_1611,In_2828,In_1715);
nand U1612 (N_1612,In_2910,In_2542);
nand U1613 (N_1613,In_1702,In_837);
and U1614 (N_1614,In_526,In_1606);
nor U1615 (N_1615,In_1740,In_2617);
or U1616 (N_1616,In_1665,In_2604);
nor U1617 (N_1617,In_1245,In_2412);
or U1618 (N_1618,In_460,In_852);
or U1619 (N_1619,In_1311,In_373);
or U1620 (N_1620,In_2922,In_2605);
nor U1621 (N_1621,In_1704,In_1150);
or U1622 (N_1622,In_2765,In_3);
nand U1623 (N_1623,In_1446,In_728);
or U1624 (N_1624,In_2109,In_495);
or U1625 (N_1625,In_475,In_223);
or U1626 (N_1626,In_1160,In_2820);
nand U1627 (N_1627,In_1061,In_745);
nor U1628 (N_1628,In_920,In_2612);
nor U1629 (N_1629,In_1995,In_2271);
nor U1630 (N_1630,In_966,In_1816);
and U1631 (N_1631,In_1743,In_721);
nor U1632 (N_1632,In_1712,In_26);
nor U1633 (N_1633,In_2149,In_1354);
nand U1634 (N_1634,In_2538,In_1029);
nor U1635 (N_1635,In_2457,In_2315);
and U1636 (N_1636,In_1133,In_600);
nor U1637 (N_1637,In_1728,In_2270);
and U1638 (N_1638,In_1779,In_65);
and U1639 (N_1639,In_1285,In_1249);
xor U1640 (N_1640,In_2828,In_1677);
and U1641 (N_1641,In_1666,In_2846);
and U1642 (N_1642,In_2297,In_2112);
xor U1643 (N_1643,In_2290,In_551);
nand U1644 (N_1644,In_748,In_2535);
and U1645 (N_1645,In_1928,In_2706);
nor U1646 (N_1646,In_435,In_2873);
and U1647 (N_1647,In_1172,In_1340);
nor U1648 (N_1648,In_440,In_2628);
and U1649 (N_1649,In_1281,In_2966);
nand U1650 (N_1650,In_2935,In_1513);
and U1651 (N_1651,In_1442,In_2052);
nor U1652 (N_1652,In_45,In_1478);
and U1653 (N_1653,In_1259,In_1860);
or U1654 (N_1654,In_2878,In_1006);
nand U1655 (N_1655,In_896,In_2024);
and U1656 (N_1656,In_1308,In_2473);
nor U1657 (N_1657,In_1358,In_1673);
nand U1658 (N_1658,In_432,In_2810);
or U1659 (N_1659,In_219,In_551);
or U1660 (N_1660,In_923,In_742);
or U1661 (N_1661,In_2965,In_2621);
nor U1662 (N_1662,In_913,In_2679);
and U1663 (N_1663,In_2999,In_2466);
nor U1664 (N_1664,In_2351,In_2663);
nand U1665 (N_1665,In_882,In_2010);
nor U1666 (N_1666,In_1644,In_1983);
xnor U1667 (N_1667,In_165,In_182);
and U1668 (N_1668,In_1614,In_427);
or U1669 (N_1669,In_2492,In_2163);
nor U1670 (N_1670,In_1000,In_1338);
nor U1671 (N_1671,In_2331,In_1443);
nand U1672 (N_1672,In_1941,In_1208);
nor U1673 (N_1673,In_1174,In_398);
or U1674 (N_1674,In_572,In_719);
nand U1675 (N_1675,In_247,In_960);
and U1676 (N_1676,In_2934,In_915);
and U1677 (N_1677,In_376,In_1911);
nand U1678 (N_1678,In_1780,In_1572);
nand U1679 (N_1679,In_2460,In_2865);
nor U1680 (N_1680,In_25,In_880);
nor U1681 (N_1681,In_542,In_2061);
nor U1682 (N_1682,In_1090,In_381);
nand U1683 (N_1683,In_2546,In_2542);
nor U1684 (N_1684,In_2036,In_97);
and U1685 (N_1685,In_1906,In_2985);
nand U1686 (N_1686,In_1894,In_2082);
and U1687 (N_1687,In_1677,In_2050);
and U1688 (N_1688,In_1808,In_2226);
nor U1689 (N_1689,In_1885,In_744);
nor U1690 (N_1690,In_426,In_1756);
or U1691 (N_1691,In_1668,In_404);
or U1692 (N_1692,In_913,In_1373);
or U1693 (N_1693,In_2667,In_1225);
nand U1694 (N_1694,In_893,In_2671);
or U1695 (N_1695,In_883,In_974);
nor U1696 (N_1696,In_0,In_490);
or U1697 (N_1697,In_289,In_1284);
and U1698 (N_1698,In_2222,In_50);
and U1699 (N_1699,In_2306,In_2581);
and U1700 (N_1700,In_1044,In_649);
nand U1701 (N_1701,In_441,In_2672);
nand U1702 (N_1702,In_2404,In_2530);
or U1703 (N_1703,In_1305,In_2055);
and U1704 (N_1704,In_647,In_504);
or U1705 (N_1705,In_324,In_1776);
and U1706 (N_1706,In_2563,In_1746);
and U1707 (N_1707,In_932,In_11);
nor U1708 (N_1708,In_677,In_2585);
and U1709 (N_1709,In_1966,In_1634);
nor U1710 (N_1710,In_2133,In_715);
or U1711 (N_1711,In_1044,In_1789);
and U1712 (N_1712,In_177,In_1159);
nor U1713 (N_1713,In_2179,In_1988);
nand U1714 (N_1714,In_1449,In_643);
nand U1715 (N_1715,In_1089,In_1421);
or U1716 (N_1716,In_2542,In_1352);
nand U1717 (N_1717,In_867,In_557);
nor U1718 (N_1718,In_1344,In_1865);
nor U1719 (N_1719,In_2059,In_2376);
nand U1720 (N_1720,In_1028,In_2534);
nand U1721 (N_1721,In_495,In_2727);
nor U1722 (N_1722,In_1305,In_1712);
or U1723 (N_1723,In_1555,In_2572);
and U1724 (N_1724,In_1112,In_2780);
nor U1725 (N_1725,In_1875,In_2073);
and U1726 (N_1726,In_614,In_2821);
and U1727 (N_1727,In_2992,In_1122);
nand U1728 (N_1728,In_911,In_509);
or U1729 (N_1729,In_1058,In_512);
nor U1730 (N_1730,In_1446,In_1726);
and U1731 (N_1731,In_2685,In_2515);
nand U1732 (N_1732,In_1030,In_146);
and U1733 (N_1733,In_2394,In_2431);
or U1734 (N_1734,In_2795,In_651);
nor U1735 (N_1735,In_2715,In_1495);
nor U1736 (N_1736,In_656,In_2688);
or U1737 (N_1737,In_2890,In_1279);
or U1738 (N_1738,In_860,In_2932);
nand U1739 (N_1739,In_1832,In_623);
or U1740 (N_1740,In_2429,In_2215);
and U1741 (N_1741,In_434,In_372);
and U1742 (N_1742,In_609,In_2410);
nor U1743 (N_1743,In_983,In_995);
nand U1744 (N_1744,In_2569,In_46);
nor U1745 (N_1745,In_1089,In_308);
and U1746 (N_1746,In_1198,In_1875);
nand U1747 (N_1747,In_1217,In_1835);
or U1748 (N_1748,In_2002,In_0);
nand U1749 (N_1749,In_1993,In_2872);
or U1750 (N_1750,In_2544,In_2364);
and U1751 (N_1751,In_1044,In_1488);
nor U1752 (N_1752,In_2546,In_1632);
or U1753 (N_1753,In_2575,In_492);
nand U1754 (N_1754,In_1965,In_685);
or U1755 (N_1755,In_1384,In_972);
nor U1756 (N_1756,In_269,In_1373);
or U1757 (N_1757,In_2385,In_2587);
nand U1758 (N_1758,In_1659,In_1363);
nand U1759 (N_1759,In_1628,In_343);
or U1760 (N_1760,In_1037,In_1667);
or U1761 (N_1761,In_948,In_1196);
or U1762 (N_1762,In_157,In_2275);
nor U1763 (N_1763,In_974,In_1205);
and U1764 (N_1764,In_515,In_2498);
or U1765 (N_1765,In_122,In_1003);
and U1766 (N_1766,In_2763,In_1338);
xor U1767 (N_1767,In_1643,In_205);
nand U1768 (N_1768,In_987,In_1226);
or U1769 (N_1769,In_1331,In_450);
or U1770 (N_1770,In_943,In_659);
nor U1771 (N_1771,In_811,In_1938);
and U1772 (N_1772,In_2168,In_580);
or U1773 (N_1773,In_1718,In_1241);
nand U1774 (N_1774,In_2658,In_2786);
or U1775 (N_1775,In_2015,In_306);
nor U1776 (N_1776,In_661,In_2782);
and U1777 (N_1777,In_2161,In_2402);
nand U1778 (N_1778,In_37,In_2539);
nand U1779 (N_1779,In_2348,In_2215);
and U1780 (N_1780,In_2648,In_765);
or U1781 (N_1781,In_198,In_1118);
nor U1782 (N_1782,In_967,In_763);
and U1783 (N_1783,In_2009,In_1914);
and U1784 (N_1784,In_1593,In_2230);
nor U1785 (N_1785,In_1288,In_2517);
nand U1786 (N_1786,In_1612,In_2095);
or U1787 (N_1787,In_1623,In_2072);
nand U1788 (N_1788,In_2907,In_1140);
nor U1789 (N_1789,In_2394,In_633);
nand U1790 (N_1790,In_1889,In_1578);
nor U1791 (N_1791,In_1072,In_512);
and U1792 (N_1792,In_625,In_2830);
and U1793 (N_1793,In_201,In_1625);
and U1794 (N_1794,In_590,In_406);
nor U1795 (N_1795,In_1534,In_229);
and U1796 (N_1796,In_1951,In_864);
nand U1797 (N_1797,In_1255,In_82);
and U1798 (N_1798,In_1375,In_2981);
nand U1799 (N_1799,In_374,In_2288);
nand U1800 (N_1800,In_270,In_674);
and U1801 (N_1801,In_2004,In_1129);
or U1802 (N_1802,In_1269,In_2786);
nor U1803 (N_1803,In_1635,In_2161);
nor U1804 (N_1804,In_585,In_440);
nor U1805 (N_1805,In_96,In_1298);
or U1806 (N_1806,In_131,In_2395);
nand U1807 (N_1807,In_202,In_1610);
and U1808 (N_1808,In_331,In_1663);
and U1809 (N_1809,In_2330,In_1725);
nand U1810 (N_1810,In_2831,In_2832);
nor U1811 (N_1811,In_704,In_467);
nor U1812 (N_1812,In_257,In_1735);
nand U1813 (N_1813,In_859,In_271);
and U1814 (N_1814,In_1893,In_1751);
nand U1815 (N_1815,In_1628,In_75);
or U1816 (N_1816,In_1059,In_1241);
nor U1817 (N_1817,In_799,In_1199);
or U1818 (N_1818,In_1110,In_1464);
nor U1819 (N_1819,In_1018,In_2140);
and U1820 (N_1820,In_175,In_1298);
nor U1821 (N_1821,In_103,In_633);
or U1822 (N_1822,In_1543,In_1985);
and U1823 (N_1823,In_2943,In_1817);
and U1824 (N_1824,In_105,In_620);
nor U1825 (N_1825,In_2965,In_1322);
nor U1826 (N_1826,In_1327,In_1573);
xnor U1827 (N_1827,In_12,In_838);
nand U1828 (N_1828,In_0,In_639);
or U1829 (N_1829,In_419,In_1413);
nand U1830 (N_1830,In_543,In_1723);
or U1831 (N_1831,In_2674,In_615);
nor U1832 (N_1832,In_1803,In_1875);
nand U1833 (N_1833,In_840,In_1386);
nand U1834 (N_1834,In_318,In_1501);
nand U1835 (N_1835,In_1536,In_2183);
or U1836 (N_1836,In_1206,In_1791);
nand U1837 (N_1837,In_2066,In_2388);
and U1838 (N_1838,In_2227,In_681);
nand U1839 (N_1839,In_1549,In_698);
nand U1840 (N_1840,In_387,In_26);
and U1841 (N_1841,In_2822,In_2020);
nand U1842 (N_1842,In_2133,In_928);
nand U1843 (N_1843,In_759,In_1431);
nor U1844 (N_1844,In_1553,In_853);
and U1845 (N_1845,In_2106,In_2974);
or U1846 (N_1846,In_41,In_1672);
and U1847 (N_1847,In_1179,In_329);
nand U1848 (N_1848,In_864,In_321);
or U1849 (N_1849,In_2133,In_917);
nand U1850 (N_1850,In_2037,In_1963);
nor U1851 (N_1851,In_2725,In_785);
and U1852 (N_1852,In_2478,In_160);
nand U1853 (N_1853,In_2306,In_493);
or U1854 (N_1854,In_890,In_87);
nor U1855 (N_1855,In_1274,In_1198);
and U1856 (N_1856,In_2596,In_1787);
or U1857 (N_1857,In_1903,In_1197);
nor U1858 (N_1858,In_2577,In_38);
or U1859 (N_1859,In_1861,In_2534);
nand U1860 (N_1860,In_1903,In_1117);
nand U1861 (N_1861,In_1210,In_1738);
or U1862 (N_1862,In_1747,In_142);
nor U1863 (N_1863,In_1350,In_1936);
nand U1864 (N_1864,In_229,In_794);
nand U1865 (N_1865,In_2583,In_958);
nand U1866 (N_1866,In_2392,In_2365);
nand U1867 (N_1867,In_1011,In_838);
and U1868 (N_1868,In_840,In_457);
or U1869 (N_1869,In_1482,In_1349);
or U1870 (N_1870,In_2478,In_2548);
nand U1871 (N_1871,In_2827,In_2213);
nor U1872 (N_1872,In_2265,In_152);
and U1873 (N_1873,In_250,In_638);
or U1874 (N_1874,In_1704,In_952);
and U1875 (N_1875,In_1652,In_2615);
or U1876 (N_1876,In_2865,In_303);
or U1877 (N_1877,In_1076,In_2762);
nor U1878 (N_1878,In_2713,In_2777);
nor U1879 (N_1879,In_425,In_1671);
and U1880 (N_1880,In_307,In_1305);
and U1881 (N_1881,In_520,In_680);
nor U1882 (N_1882,In_2505,In_2858);
or U1883 (N_1883,In_1933,In_992);
nand U1884 (N_1884,In_2047,In_2840);
nand U1885 (N_1885,In_683,In_2297);
and U1886 (N_1886,In_2765,In_7);
and U1887 (N_1887,In_732,In_2528);
or U1888 (N_1888,In_1212,In_2529);
or U1889 (N_1889,In_1540,In_1465);
nor U1890 (N_1890,In_497,In_1920);
and U1891 (N_1891,In_2453,In_2281);
and U1892 (N_1892,In_2638,In_1485);
and U1893 (N_1893,In_2407,In_75);
nand U1894 (N_1894,In_2755,In_2053);
and U1895 (N_1895,In_349,In_1063);
or U1896 (N_1896,In_1561,In_2258);
nor U1897 (N_1897,In_1522,In_337);
and U1898 (N_1898,In_183,In_206);
or U1899 (N_1899,In_1757,In_2370);
nor U1900 (N_1900,In_594,In_2003);
and U1901 (N_1901,In_2787,In_1953);
nand U1902 (N_1902,In_388,In_1768);
nor U1903 (N_1903,In_638,In_830);
or U1904 (N_1904,In_643,In_413);
or U1905 (N_1905,In_1826,In_236);
or U1906 (N_1906,In_2637,In_1278);
nand U1907 (N_1907,In_1205,In_643);
or U1908 (N_1908,In_1210,In_434);
nor U1909 (N_1909,In_2060,In_1205);
and U1910 (N_1910,In_1839,In_2520);
and U1911 (N_1911,In_2107,In_2852);
or U1912 (N_1912,In_104,In_2303);
nor U1913 (N_1913,In_2811,In_698);
or U1914 (N_1914,In_1506,In_124);
nand U1915 (N_1915,In_2539,In_2);
and U1916 (N_1916,In_2769,In_607);
nand U1917 (N_1917,In_137,In_600);
nor U1918 (N_1918,In_741,In_1594);
or U1919 (N_1919,In_1656,In_228);
and U1920 (N_1920,In_1061,In_1343);
or U1921 (N_1921,In_2440,In_2174);
or U1922 (N_1922,In_1624,In_153);
nand U1923 (N_1923,In_683,In_1011);
nor U1924 (N_1924,In_316,In_2541);
nand U1925 (N_1925,In_2354,In_525);
or U1926 (N_1926,In_2929,In_1055);
nor U1927 (N_1927,In_1479,In_2390);
and U1928 (N_1928,In_2764,In_749);
xor U1929 (N_1929,In_2702,In_750);
nand U1930 (N_1930,In_2705,In_1081);
nor U1931 (N_1931,In_2229,In_2640);
nor U1932 (N_1932,In_384,In_2680);
and U1933 (N_1933,In_2089,In_2809);
or U1934 (N_1934,In_2366,In_821);
and U1935 (N_1935,In_1806,In_910);
nor U1936 (N_1936,In_1256,In_531);
nand U1937 (N_1937,In_1084,In_959);
nand U1938 (N_1938,In_1808,In_817);
and U1939 (N_1939,In_68,In_506);
nor U1940 (N_1940,In_1306,In_2862);
nor U1941 (N_1941,In_2965,In_1530);
and U1942 (N_1942,In_2471,In_942);
and U1943 (N_1943,In_2524,In_1427);
nor U1944 (N_1944,In_2399,In_1354);
nand U1945 (N_1945,In_706,In_1379);
or U1946 (N_1946,In_2059,In_1837);
and U1947 (N_1947,In_1206,In_1587);
nor U1948 (N_1948,In_2936,In_1085);
and U1949 (N_1949,In_575,In_6);
nor U1950 (N_1950,In_787,In_1971);
or U1951 (N_1951,In_2358,In_1911);
nor U1952 (N_1952,In_1923,In_570);
and U1953 (N_1953,In_1168,In_926);
nor U1954 (N_1954,In_1395,In_1865);
or U1955 (N_1955,In_1612,In_2561);
nor U1956 (N_1956,In_1956,In_2808);
nor U1957 (N_1957,In_2917,In_471);
and U1958 (N_1958,In_545,In_394);
nor U1959 (N_1959,In_1814,In_2952);
nand U1960 (N_1960,In_1577,In_1902);
nor U1961 (N_1961,In_1342,In_965);
or U1962 (N_1962,In_2166,In_1433);
and U1963 (N_1963,In_880,In_1046);
and U1964 (N_1964,In_819,In_1052);
nand U1965 (N_1965,In_1067,In_816);
nor U1966 (N_1966,In_621,In_1892);
nor U1967 (N_1967,In_2958,In_148);
nor U1968 (N_1968,In_1405,In_2429);
and U1969 (N_1969,In_1868,In_1303);
and U1970 (N_1970,In_289,In_1994);
or U1971 (N_1971,In_1349,In_662);
and U1972 (N_1972,In_1806,In_389);
nand U1973 (N_1973,In_356,In_2358);
nor U1974 (N_1974,In_598,In_267);
nor U1975 (N_1975,In_538,In_1752);
nand U1976 (N_1976,In_1399,In_470);
xnor U1977 (N_1977,In_2101,In_28);
nor U1978 (N_1978,In_117,In_1486);
nand U1979 (N_1979,In_2762,In_2779);
xnor U1980 (N_1980,In_416,In_2016);
and U1981 (N_1981,In_1892,In_1284);
and U1982 (N_1982,In_2669,In_1319);
and U1983 (N_1983,In_1829,In_2350);
nand U1984 (N_1984,In_2467,In_2704);
nor U1985 (N_1985,In_124,In_278);
or U1986 (N_1986,In_257,In_182);
or U1987 (N_1987,In_2432,In_2224);
and U1988 (N_1988,In_720,In_2272);
nor U1989 (N_1989,In_841,In_67);
or U1990 (N_1990,In_844,In_2404);
nor U1991 (N_1991,In_2467,In_629);
nand U1992 (N_1992,In_2360,In_370);
or U1993 (N_1993,In_29,In_1358);
or U1994 (N_1994,In_1309,In_2159);
nor U1995 (N_1995,In_2203,In_830);
nor U1996 (N_1996,In_2955,In_536);
nor U1997 (N_1997,In_158,In_962);
or U1998 (N_1998,In_2642,In_2641);
or U1999 (N_1999,In_606,In_867);
and U2000 (N_2000,In_2055,In_820);
and U2001 (N_2001,In_359,In_2626);
nand U2002 (N_2002,In_1632,In_2286);
or U2003 (N_2003,In_1292,In_1681);
nor U2004 (N_2004,In_1716,In_2126);
or U2005 (N_2005,In_144,In_243);
or U2006 (N_2006,In_1860,In_1591);
and U2007 (N_2007,In_46,In_1196);
and U2008 (N_2008,In_2692,In_465);
and U2009 (N_2009,In_2968,In_1644);
or U2010 (N_2010,In_644,In_1282);
and U2011 (N_2011,In_550,In_773);
or U2012 (N_2012,In_2304,In_2062);
or U2013 (N_2013,In_1246,In_1382);
and U2014 (N_2014,In_1320,In_389);
and U2015 (N_2015,In_2951,In_694);
and U2016 (N_2016,In_2969,In_1827);
nand U2017 (N_2017,In_618,In_410);
or U2018 (N_2018,In_798,In_805);
or U2019 (N_2019,In_2849,In_2660);
nor U2020 (N_2020,In_1788,In_2190);
nor U2021 (N_2021,In_1010,In_1438);
nand U2022 (N_2022,In_1048,In_2230);
and U2023 (N_2023,In_512,In_1594);
nor U2024 (N_2024,In_574,In_1191);
or U2025 (N_2025,In_2501,In_2193);
nor U2026 (N_2026,In_1880,In_2040);
nor U2027 (N_2027,In_17,In_124);
and U2028 (N_2028,In_835,In_971);
and U2029 (N_2029,In_1262,In_1329);
or U2030 (N_2030,In_2007,In_1711);
nand U2031 (N_2031,In_2774,In_382);
nor U2032 (N_2032,In_385,In_2553);
nand U2033 (N_2033,In_819,In_2210);
nor U2034 (N_2034,In_2046,In_1033);
nor U2035 (N_2035,In_807,In_2817);
nand U2036 (N_2036,In_918,In_624);
and U2037 (N_2037,In_2903,In_307);
nand U2038 (N_2038,In_396,In_732);
and U2039 (N_2039,In_771,In_2823);
nand U2040 (N_2040,In_405,In_125);
and U2041 (N_2041,In_494,In_2721);
nor U2042 (N_2042,In_390,In_2976);
or U2043 (N_2043,In_2248,In_1952);
and U2044 (N_2044,In_2568,In_2497);
nor U2045 (N_2045,In_1336,In_1208);
nand U2046 (N_2046,In_1196,In_2640);
and U2047 (N_2047,In_1188,In_2253);
or U2048 (N_2048,In_2973,In_553);
nand U2049 (N_2049,In_1455,In_668);
nand U2050 (N_2050,In_2243,In_2161);
nand U2051 (N_2051,In_1321,In_180);
nor U2052 (N_2052,In_638,In_452);
and U2053 (N_2053,In_2202,In_2355);
nand U2054 (N_2054,In_1323,In_1960);
nand U2055 (N_2055,In_1645,In_812);
or U2056 (N_2056,In_2457,In_1462);
nor U2057 (N_2057,In_180,In_1189);
or U2058 (N_2058,In_72,In_2567);
nand U2059 (N_2059,In_2492,In_1542);
and U2060 (N_2060,In_478,In_922);
and U2061 (N_2061,In_339,In_1691);
or U2062 (N_2062,In_61,In_2753);
nand U2063 (N_2063,In_1076,In_2822);
and U2064 (N_2064,In_682,In_1862);
nand U2065 (N_2065,In_2233,In_2182);
or U2066 (N_2066,In_1459,In_178);
or U2067 (N_2067,In_1921,In_2045);
or U2068 (N_2068,In_915,In_964);
nand U2069 (N_2069,In_333,In_1717);
nand U2070 (N_2070,In_1942,In_1455);
or U2071 (N_2071,In_602,In_2602);
or U2072 (N_2072,In_326,In_2233);
nor U2073 (N_2073,In_1688,In_2289);
nand U2074 (N_2074,In_566,In_1016);
nand U2075 (N_2075,In_548,In_294);
nand U2076 (N_2076,In_2831,In_2021);
nor U2077 (N_2077,In_1474,In_2266);
or U2078 (N_2078,In_2533,In_2422);
nor U2079 (N_2079,In_2122,In_1712);
nor U2080 (N_2080,In_632,In_2382);
or U2081 (N_2081,In_1004,In_1342);
nand U2082 (N_2082,In_1627,In_1238);
nand U2083 (N_2083,In_1495,In_118);
or U2084 (N_2084,In_1180,In_2817);
nand U2085 (N_2085,In_750,In_313);
nor U2086 (N_2086,In_2245,In_2105);
nor U2087 (N_2087,In_2941,In_336);
nand U2088 (N_2088,In_2614,In_781);
nor U2089 (N_2089,In_1974,In_2866);
nor U2090 (N_2090,In_894,In_508);
or U2091 (N_2091,In_1575,In_2685);
nand U2092 (N_2092,In_2084,In_480);
and U2093 (N_2093,In_730,In_492);
or U2094 (N_2094,In_1276,In_176);
or U2095 (N_2095,In_2962,In_727);
or U2096 (N_2096,In_1785,In_295);
and U2097 (N_2097,In_147,In_92);
nand U2098 (N_2098,In_2192,In_2070);
nand U2099 (N_2099,In_710,In_1647);
or U2100 (N_2100,In_928,In_2303);
or U2101 (N_2101,In_334,In_2685);
nand U2102 (N_2102,In_1282,In_990);
nor U2103 (N_2103,In_1020,In_1001);
and U2104 (N_2104,In_2019,In_2044);
and U2105 (N_2105,In_1389,In_2345);
nand U2106 (N_2106,In_194,In_898);
nand U2107 (N_2107,In_565,In_222);
nor U2108 (N_2108,In_37,In_2978);
nand U2109 (N_2109,In_1714,In_1261);
or U2110 (N_2110,In_762,In_866);
and U2111 (N_2111,In_270,In_2088);
and U2112 (N_2112,In_290,In_2803);
nor U2113 (N_2113,In_2018,In_2327);
nor U2114 (N_2114,In_1646,In_1045);
nor U2115 (N_2115,In_2501,In_2109);
nand U2116 (N_2116,In_680,In_2830);
nand U2117 (N_2117,In_2630,In_183);
or U2118 (N_2118,In_2247,In_2437);
nand U2119 (N_2119,In_1746,In_208);
and U2120 (N_2120,In_440,In_234);
nor U2121 (N_2121,In_2194,In_1659);
or U2122 (N_2122,In_2564,In_2050);
or U2123 (N_2123,In_1220,In_2402);
or U2124 (N_2124,In_1874,In_1682);
or U2125 (N_2125,In_433,In_1319);
and U2126 (N_2126,In_522,In_1312);
or U2127 (N_2127,In_2857,In_2887);
or U2128 (N_2128,In_1414,In_1122);
nand U2129 (N_2129,In_583,In_1803);
nor U2130 (N_2130,In_588,In_716);
or U2131 (N_2131,In_2065,In_2107);
and U2132 (N_2132,In_2744,In_2480);
and U2133 (N_2133,In_1003,In_2254);
nand U2134 (N_2134,In_1405,In_2605);
nor U2135 (N_2135,In_1239,In_1333);
nand U2136 (N_2136,In_790,In_2432);
and U2137 (N_2137,In_1928,In_2893);
or U2138 (N_2138,In_1127,In_294);
or U2139 (N_2139,In_908,In_60);
and U2140 (N_2140,In_333,In_2660);
and U2141 (N_2141,In_1512,In_2290);
nand U2142 (N_2142,In_829,In_176);
nand U2143 (N_2143,In_431,In_277);
and U2144 (N_2144,In_923,In_2388);
and U2145 (N_2145,In_2814,In_2853);
nand U2146 (N_2146,In_1384,In_1943);
and U2147 (N_2147,In_2304,In_1833);
nor U2148 (N_2148,In_298,In_806);
nor U2149 (N_2149,In_791,In_2551);
or U2150 (N_2150,In_2736,In_452);
nand U2151 (N_2151,In_1826,In_1954);
nand U2152 (N_2152,In_278,In_2002);
and U2153 (N_2153,In_1823,In_516);
nor U2154 (N_2154,In_725,In_2087);
nor U2155 (N_2155,In_306,In_646);
or U2156 (N_2156,In_2794,In_2410);
nor U2157 (N_2157,In_1509,In_67);
nor U2158 (N_2158,In_2560,In_409);
nand U2159 (N_2159,In_2255,In_2570);
and U2160 (N_2160,In_1466,In_2250);
nor U2161 (N_2161,In_2079,In_1795);
nand U2162 (N_2162,In_107,In_1533);
nor U2163 (N_2163,In_1952,In_2236);
nand U2164 (N_2164,In_910,In_2144);
and U2165 (N_2165,In_1968,In_622);
and U2166 (N_2166,In_1864,In_410);
and U2167 (N_2167,In_1483,In_2780);
and U2168 (N_2168,In_344,In_2480);
nor U2169 (N_2169,In_1218,In_2373);
and U2170 (N_2170,In_636,In_1232);
nor U2171 (N_2171,In_1628,In_2407);
nor U2172 (N_2172,In_1829,In_964);
or U2173 (N_2173,In_2072,In_631);
nor U2174 (N_2174,In_2437,In_287);
and U2175 (N_2175,In_2622,In_413);
and U2176 (N_2176,In_1607,In_850);
or U2177 (N_2177,In_879,In_1511);
and U2178 (N_2178,In_1574,In_720);
and U2179 (N_2179,In_35,In_1253);
or U2180 (N_2180,In_1435,In_1507);
xnor U2181 (N_2181,In_575,In_2341);
nand U2182 (N_2182,In_1260,In_806);
and U2183 (N_2183,In_1039,In_2286);
or U2184 (N_2184,In_2719,In_884);
or U2185 (N_2185,In_1875,In_2032);
and U2186 (N_2186,In_2579,In_1785);
nor U2187 (N_2187,In_2795,In_230);
nor U2188 (N_2188,In_1740,In_518);
or U2189 (N_2189,In_1049,In_1457);
nor U2190 (N_2190,In_820,In_2912);
nand U2191 (N_2191,In_2050,In_2352);
nor U2192 (N_2192,In_725,In_2150);
nor U2193 (N_2193,In_224,In_1223);
nor U2194 (N_2194,In_1628,In_314);
and U2195 (N_2195,In_1532,In_1834);
nand U2196 (N_2196,In_985,In_603);
and U2197 (N_2197,In_2041,In_2310);
or U2198 (N_2198,In_881,In_713);
nor U2199 (N_2199,In_2564,In_578);
nand U2200 (N_2200,In_554,In_2592);
nand U2201 (N_2201,In_1776,In_2318);
nand U2202 (N_2202,In_1651,In_1428);
nor U2203 (N_2203,In_1557,In_876);
or U2204 (N_2204,In_1739,In_2011);
nor U2205 (N_2205,In_414,In_107);
and U2206 (N_2206,In_1742,In_804);
nor U2207 (N_2207,In_2401,In_2274);
nand U2208 (N_2208,In_2955,In_312);
nand U2209 (N_2209,In_1914,In_667);
nand U2210 (N_2210,In_1238,In_301);
or U2211 (N_2211,In_2860,In_1989);
nor U2212 (N_2212,In_1412,In_2516);
nor U2213 (N_2213,In_2038,In_177);
and U2214 (N_2214,In_1800,In_1221);
and U2215 (N_2215,In_1751,In_2534);
nor U2216 (N_2216,In_766,In_2567);
nor U2217 (N_2217,In_529,In_1209);
nor U2218 (N_2218,In_555,In_101);
and U2219 (N_2219,In_2160,In_701);
nor U2220 (N_2220,In_1953,In_1156);
and U2221 (N_2221,In_2743,In_1020);
and U2222 (N_2222,In_979,In_1815);
or U2223 (N_2223,In_1712,In_714);
nor U2224 (N_2224,In_178,In_1040);
nand U2225 (N_2225,In_2707,In_2276);
nor U2226 (N_2226,In_2339,In_1705);
nand U2227 (N_2227,In_1573,In_2854);
xor U2228 (N_2228,In_190,In_1828);
nor U2229 (N_2229,In_145,In_442);
and U2230 (N_2230,In_2301,In_309);
or U2231 (N_2231,In_2093,In_2014);
or U2232 (N_2232,In_753,In_2812);
and U2233 (N_2233,In_2826,In_1853);
nor U2234 (N_2234,In_1513,In_101);
or U2235 (N_2235,In_1930,In_62);
nand U2236 (N_2236,In_84,In_2345);
or U2237 (N_2237,In_1468,In_1875);
and U2238 (N_2238,In_352,In_537);
nor U2239 (N_2239,In_2541,In_1652);
or U2240 (N_2240,In_641,In_1284);
or U2241 (N_2241,In_1504,In_1347);
nor U2242 (N_2242,In_2225,In_2792);
nand U2243 (N_2243,In_2021,In_41);
nand U2244 (N_2244,In_820,In_1099);
and U2245 (N_2245,In_1047,In_2109);
and U2246 (N_2246,In_922,In_1238);
nor U2247 (N_2247,In_388,In_2303);
nand U2248 (N_2248,In_2165,In_2630);
and U2249 (N_2249,In_528,In_2203);
and U2250 (N_2250,In_613,In_2027);
nand U2251 (N_2251,In_764,In_2944);
nand U2252 (N_2252,In_2206,In_1772);
or U2253 (N_2253,In_583,In_992);
xnor U2254 (N_2254,In_2987,In_1225);
nand U2255 (N_2255,In_265,In_2951);
and U2256 (N_2256,In_2540,In_894);
or U2257 (N_2257,In_983,In_283);
nand U2258 (N_2258,In_2845,In_2727);
nor U2259 (N_2259,In_192,In_1159);
and U2260 (N_2260,In_2058,In_197);
nand U2261 (N_2261,In_1779,In_2074);
or U2262 (N_2262,In_635,In_2157);
or U2263 (N_2263,In_2864,In_1504);
and U2264 (N_2264,In_153,In_2859);
and U2265 (N_2265,In_2494,In_2883);
xor U2266 (N_2266,In_94,In_832);
or U2267 (N_2267,In_666,In_142);
nand U2268 (N_2268,In_2654,In_1103);
and U2269 (N_2269,In_2569,In_1747);
xor U2270 (N_2270,In_2060,In_112);
nor U2271 (N_2271,In_1489,In_1741);
or U2272 (N_2272,In_1803,In_1005);
nor U2273 (N_2273,In_563,In_1736);
nand U2274 (N_2274,In_389,In_212);
and U2275 (N_2275,In_2607,In_725);
nor U2276 (N_2276,In_1405,In_1526);
nor U2277 (N_2277,In_2135,In_1712);
nand U2278 (N_2278,In_2395,In_2700);
or U2279 (N_2279,In_2797,In_2215);
nor U2280 (N_2280,In_21,In_1504);
nor U2281 (N_2281,In_1672,In_2547);
nor U2282 (N_2282,In_950,In_1548);
nand U2283 (N_2283,In_2028,In_1511);
nand U2284 (N_2284,In_2375,In_2737);
nand U2285 (N_2285,In_2246,In_1321);
and U2286 (N_2286,In_896,In_620);
or U2287 (N_2287,In_1770,In_1072);
and U2288 (N_2288,In_2054,In_1174);
nor U2289 (N_2289,In_1472,In_2964);
or U2290 (N_2290,In_1915,In_1713);
nor U2291 (N_2291,In_2883,In_284);
and U2292 (N_2292,In_2715,In_726);
nand U2293 (N_2293,In_749,In_35);
nor U2294 (N_2294,In_2739,In_2130);
nor U2295 (N_2295,In_1059,In_716);
nor U2296 (N_2296,In_1214,In_2972);
or U2297 (N_2297,In_2929,In_455);
and U2298 (N_2298,In_2140,In_2080);
nand U2299 (N_2299,In_1425,In_2584);
and U2300 (N_2300,In_2861,In_2138);
or U2301 (N_2301,In_304,In_372);
nand U2302 (N_2302,In_2890,In_2969);
or U2303 (N_2303,In_2013,In_1087);
nor U2304 (N_2304,In_1873,In_509);
or U2305 (N_2305,In_380,In_603);
nor U2306 (N_2306,In_871,In_2064);
nand U2307 (N_2307,In_485,In_622);
and U2308 (N_2308,In_2521,In_141);
or U2309 (N_2309,In_1841,In_1694);
or U2310 (N_2310,In_533,In_1057);
and U2311 (N_2311,In_1222,In_2773);
and U2312 (N_2312,In_2258,In_1994);
and U2313 (N_2313,In_986,In_2868);
or U2314 (N_2314,In_1448,In_1019);
and U2315 (N_2315,In_2690,In_1126);
nand U2316 (N_2316,In_1764,In_2922);
and U2317 (N_2317,In_1158,In_2944);
or U2318 (N_2318,In_2270,In_2201);
or U2319 (N_2319,In_682,In_1210);
nor U2320 (N_2320,In_1430,In_864);
nand U2321 (N_2321,In_246,In_886);
or U2322 (N_2322,In_649,In_152);
and U2323 (N_2323,In_2797,In_371);
and U2324 (N_2324,In_1473,In_2250);
nand U2325 (N_2325,In_2184,In_940);
nor U2326 (N_2326,In_244,In_134);
or U2327 (N_2327,In_1320,In_1270);
nand U2328 (N_2328,In_2040,In_374);
or U2329 (N_2329,In_1987,In_1557);
nor U2330 (N_2330,In_2004,In_1185);
and U2331 (N_2331,In_1567,In_226);
nor U2332 (N_2332,In_1595,In_1768);
nand U2333 (N_2333,In_2088,In_666);
and U2334 (N_2334,In_2790,In_1226);
nor U2335 (N_2335,In_848,In_408);
nand U2336 (N_2336,In_1632,In_1287);
xnor U2337 (N_2337,In_2972,In_1206);
and U2338 (N_2338,In_2938,In_1698);
nand U2339 (N_2339,In_1334,In_2452);
nor U2340 (N_2340,In_464,In_489);
nor U2341 (N_2341,In_72,In_587);
nor U2342 (N_2342,In_1760,In_2668);
nor U2343 (N_2343,In_1759,In_930);
nor U2344 (N_2344,In_2180,In_1100);
and U2345 (N_2345,In_2569,In_1477);
or U2346 (N_2346,In_2599,In_2249);
nand U2347 (N_2347,In_1134,In_98);
or U2348 (N_2348,In_1608,In_1205);
nor U2349 (N_2349,In_1677,In_611);
or U2350 (N_2350,In_2204,In_456);
and U2351 (N_2351,In_84,In_277);
and U2352 (N_2352,In_2766,In_2769);
and U2353 (N_2353,In_1504,In_2019);
nor U2354 (N_2354,In_33,In_2014);
and U2355 (N_2355,In_2694,In_2166);
and U2356 (N_2356,In_2656,In_662);
and U2357 (N_2357,In_2457,In_2092);
nor U2358 (N_2358,In_982,In_2681);
and U2359 (N_2359,In_1535,In_2464);
nor U2360 (N_2360,In_2428,In_2918);
nand U2361 (N_2361,In_1699,In_2242);
or U2362 (N_2362,In_1967,In_1998);
nor U2363 (N_2363,In_1252,In_1193);
and U2364 (N_2364,In_125,In_1861);
and U2365 (N_2365,In_2717,In_2154);
or U2366 (N_2366,In_319,In_1242);
nand U2367 (N_2367,In_1334,In_2732);
and U2368 (N_2368,In_2733,In_1300);
or U2369 (N_2369,In_2091,In_1760);
and U2370 (N_2370,In_1972,In_717);
nand U2371 (N_2371,In_2864,In_1425);
or U2372 (N_2372,In_1977,In_2659);
nor U2373 (N_2373,In_994,In_476);
nand U2374 (N_2374,In_689,In_226);
or U2375 (N_2375,In_1527,In_2814);
nand U2376 (N_2376,In_1207,In_224);
nand U2377 (N_2377,In_1434,In_1498);
or U2378 (N_2378,In_2580,In_583);
or U2379 (N_2379,In_2060,In_2983);
and U2380 (N_2380,In_244,In_1411);
and U2381 (N_2381,In_2879,In_705);
nor U2382 (N_2382,In_186,In_1721);
and U2383 (N_2383,In_1920,In_2295);
nor U2384 (N_2384,In_2305,In_2209);
and U2385 (N_2385,In_279,In_1272);
or U2386 (N_2386,In_78,In_2116);
or U2387 (N_2387,In_776,In_1561);
nand U2388 (N_2388,In_1633,In_99);
or U2389 (N_2389,In_503,In_1316);
nand U2390 (N_2390,In_1339,In_1179);
nand U2391 (N_2391,In_790,In_1921);
and U2392 (N_2392,In_207,In_2182);
nand U2393 (N_2393,In_499,In_380);
nor U2394 (N_2394,In_1991,In_153);
nor U2395 (N_2395,In_1359,In_2916);
nor U2396 (N_2396,In_221,In_2412);
or U2397 (N_2397,In_257,In_288);
or U2398 (N_2398,In_895,In_2470);
and U2399 (N_2399,In_1264,In_974);
nand U2400 (N_2400,In_371,In_2613);
nand U2401 (N_2401,In_1409,In_121);
and U2402 (N_2402,In_805,In_359);
nand U2403 (N_2403,In_2207,In_2728);
and U2404 (N_2404,In_1728,In_1558);
or U2405 (N_2405,In_1729,In_2836);
nand U2406 (N_2406,In_2750,In_668);
nor U2407 (N_2407,In_659,In_2654);
nand U2408 (N_2408,In_1656,In_1337);
nor U2409 (N_2409,In_925,In_1839);
and U2410 (N_2410,In_304,In_1339);
nand U2411 (N_2411,In_1723,In_2967);
nand U2412 (N_2412,In_2464,In_2905);
nand U2413 (N_2413,In_1355,In_1352);
and U2414 (N_2414,In_1416,In_2306);
or U2415 (N_2415,In_2448,In_983);
and U2416 (N_2416,In_1914,In_1198);
nor U2417 (N_2417,In_576,In_2353);
nand U2418 (N_2418,In_2387,In_1570);
nor U2419 (N_2419,In_2961,In_1523);
nand U2420 (N_2420,In_1777,In_779);
or U2421 (N_2421,In_2205,In_2778);
nor U2422 (N_2422,In_502,In_668);
nor U2423 (N_2423,In_810,In_2544);
nor U2424 (N_2424,In_1602,In_303);
nor U2425 (N_2425,In_1368,In_1335);
nand U2426 (N_2426,In_1393,In_74);
or U2427 (N_2427,In_1452,In_2133);
and U2428 (N_2428,In_681,In_955);
and U2429 (N_2429,In_44,In_2278);
nand U2430 (N_2430,In_381,In_1671);
or U2431 (N_2431,In_275,In_1881);
or U2432 (N_2432,In_801,In_2621);
nor U2433 (N_2433,In_744,In_2758);
nor U2434 (N_2434,In_983,In_2356);
nand U2435 (N_2435,In_2352,In_2695);
nand U2436 (N_2436,In_901,In_2674);
nor U2437 (N_2437,In_2213,In_1017);
nor U2438 (N_2438,In_2699,In_1382);
nand U2439 (N_2439,In_356,In_2337);
or U2440 (N_2440,In_2772,In_950);
or U2441 (N_2441,In_1795,In_124);
and U2442 (N_2442,In_1682,In_1580);
and U2443 (N_2443,In_1278,In_2660);
and U2444 (N_2444,In_584,In_13);
nand U2445 (N_2445,In_1448,In_2444);
xor U2446 (N_2446,In_2674,In_708);
nor U2447 (N_2447,In_890,In_1650);
nor U2448 (N_2448,In_2048,In_448);
nand U2449 (N_2449,In_226,In_645);
nand U2450 (N_2450,In_1081,In_2074);
nor U2451 (N_2451,In_27,In_1910);
nand U2452 (N_2452,In_2264,In_123);
nor U2453 (N_2453,In_1607,In_772);
or U2454 (N_2454,In_174,In_122);
or U2455 (N_2455,In_2375,In_2642);
and U2456 (N_2456,In_2826,In_1477);
nor U2457 (N_2457,In_1852,In_718);
nand U2458 (N_2458,In_1932,In_2133);
and U2459 (N_2459,In_1317,In_2842);
or U2460 (N_2460,In_2979,In_1649);
nand U2461 (N_2461,In_2051,In_899);
or U2462 (N_2462,In_2423,In_374);
and U2463 (N_2463,In_2593,In_0);
nand U2464 (N_2464,In_1932,In_1529);
nand U2465 (N_2465,In_2118,In_399);
nand U2466 (N_2466,In_426,In_2063);
nor U2467 (N_2467,In_1089,In_1298);
and U2468 (N_2468,In_1908,In_1778);
nand U2469 (N_2469,In_2894,In_1103);
nor U2470 (N_2470,In_773,In_1748);
and U2471 (N_2471,In_489,In_217);
and U2472 (N_2472,In_1373,In_1803);
or U2473 (N_2473,In_892,In_2961);
nand U2474 (N_2474,In_901,In_2592);
nor U2475 (N_2475,In_2675,In_2568);
nor U2476 (N_2476,In_1622,In_227);
or U2477 (N_2477,In_1927,In_1429);
or U2478 (N_2478,In_1032,In_2769);
or U2479 (N_2479,In_1069,In_431);
and U2480 (N_2480,In_1450,In_2178);
or U2481 (N_2481,In_445,In_2975);
nor U2482 (N_2482,In_2901,In_1193);
or U2483 (N_2483,In_2838,In_2533);
and U2484 (N_2484,In_356,In_314);
nor U2485 (N_2485,In_2462,In_1993);
and U2486 (N_2486,In_35,In_954);
or U2487 (N_2487,In_356,In_1544);
nand U2488 (N_2488,In_2421,In_1626);
and U2489 (N_2489,In_2010,In_861);
nor U2490 (N_2490,In_497,In_2774);
or U2491 (N_2491,In_572,In_2252);
or U2492 (N_2492,In_954,In_274);
nor U2493 (N_2493,In_1574,In_386);
nor U2494 (N_2494,In_1638,In_443);
nand U2495 (N_2495,In_868,In_2263);
nand U2496 (N_2496,In_2482,In_1170);
or U2497 (N_2497,In_1165,In_232);
or U2498 (N_2498,In_1365,In_2164);
nand U2499 (N_2499,In_807,In_2189);
or U2500 (N_2500,In_2341,In_1633);
or U2501 (N_2501,In_1985,In_1462);
or U2502 (N_2502,In_651,In_2821);
or U2503 (N_2503,In_2447,In_992);
nand U2504 (N_2504,In_1361,In_1395);
nand U2505 (N_2505,In_1100,In_495);
and U2506 (N_2506,In_1783,In_1080);
nor U2507 (N_2507,In_2336,In_2231);
or U2508 (N_2508,In_1733,In_801);
nand U2509 (N_2509,In_1120,In_923);
and U2510 (N_2510,In_1883,In_184);
nand U2511 (N_2511,In_519,In_58);
or U2512 (N_2512,In_2984,In_302);
or U2513 (N_2513,In_1355,In_496);
nand U2514 (N_2514,In_2814,In_1436);
or U2515 (N_2515,In_748,In_2321);
or U2516 (N_2516,In_615,In_385);
and U2517 (N_2517,In_899,In_2202);
nand U2518 (N_2518,In_1606,In_1254);
or U2519 (N_2519,In_1625,In_2305);
or U2520 (N_2520,In_2560,In_1743);
or U2521 (N_2521,In_163,In_1243);
and U2522 (N_2522,In_2532,In_602);
nor U2523 (N_2523,In_2758,In_2393);
nand U2524 (N_2524,In_2359,In_2277);
nor U2525 (N_2525,In_1217,In_1399);
or U2526 (N_2526,In_2209,In_366);
nand U2527 (N_2527,In_2783,In_1257);
and U2528 (N_2528,In_2179,In_1879);
nand U2529 (N_2529,In_1745,In_1091);
nand U2530 (N_2530,In_594,In_45);
nand U2531 (N_2531,In_1578,In_2767);
and U2532 (N_2532,In_2673,In_446);
or U2533 (N_2533,In_2874,In_1803);
nand U2534 (N_2534,In_2275,In_531);
or U2535 (N_2535,In_1385,In_1496);
nor U2536 (N_2536,In_854,In_1994);
or U2537 (N_2537,In_2722,In_1376);
nor U2538 (N_2538,In_399,In_746);
or U2539 (N_2539,In_2687,In_1798);
or U2540 (N_2540,In_1604,In_787);
and U2541 (N_2541,In_2159,In_77);
xnor U2542 (N_2542,In_981,In_723);
nand U2543 (N_2543,In_404,In_2358);
or U2544 (N_2544,In_2940,In_1094);
and U2545 (N_2545,In_2346,In_2626);
nor U2546 (N_2546,In_1255,In_1889);
nor U2547 (N_2547,In_509,In_1563);
nand U2548 (N_2548,In_2516,In_1381);
nand U2549 (N_2549,In_394,In_2332);
nand U2550 (N_2550,In_1823,In_350);
and U2551 (N_2551,In_766,In_596);
or U2552 (N_2552,In_2369,In_723);
and U2553 (N_2553,In_2810,In_2068);
or U2554 (N_2554,In_361,In_2764);
nor U2555 (N_2555,In_2091,In_1271);
nand U2556 (N_2556,In_797,In_2657);
or U2557 (N_2557,In_692,In_2416);
nor U2558 (N_2558,In_2530,In_1657);
or U2559 (N_2559,In_1589,In_1026);
nor U2560 (N_2560,In_787,In_151);
and U2561 (N_2561,In_2666,In_2516);
nor U2562 (N_2562,In_1872,In_525);
nor U2563 (N_2563,In_1380,In_1806);
nand U2564 (N_2564,In_2243,In_1845);
or U2565 (N_2565,In_2065,In_1148);
nor U2566 (N_2566,In_2609,In_2368);
nor U2567 (N_2567,In_2521,In_41);
or U2568 (N_2568,In_2758,In_166);
and U2569 (N_2569,In_3,In_1137);
nand U2570 (N_2570,In_1246,In_2097);
nor U2571 (N_2571,In_790,In_2331);
or U2572 (N_2572,In_170,In_1190);
or U2573 (N_2573,In_156,In_2956);
or U2574 (N_2574,In_2301,In_1210);
xor U2575 (N_2575,In_2218,In_206);
and U2576 (N_2576,In_2815,In_423);
nor U2577 (N_2577,In_386,In_118);
nor U2578 (N_2578,In_441,In_740);
and U2579 (N_2579,In_2430,In_182);
nand U2580 (N_2580,In_403,In_2420);
nor U2581 (N_2581,In_435,In_2223);
nor U2582 (N_2582,In_1624,In_292);
nand U2583 (N_2583,In_1607,In_2521);
or U2584 (N_2584,In_1335,In_594);
nor U2585 (N_2585,In_602,In_1989);
or U2586 (N_2586,In_1245,In_1147);
or U2587 (N_2587,In_665,In_626);
nand U2588 (N_2588,In_123,In_2134);
nand U2589 (N_2589,In_1707,In_2005);
nand U2590 (N_2590,In_2220,In_448);
or U2591 (N_2591,In_2443,In_2828);
or U2592 (N_2592,In_1259,In_225);
nand U2593 (N_2593,In_2270,In_1739);
nor U2594 (N_2594,In_2873,In_2986);
and U2595 (N_2595,In_2852,In_2148);
and U2596 (N_2596,In_444,In_2948);
or U2597 (N_2597,In_2937,In_697);
or U2598 (N_2598,In_2782,In_1403);
nor U2599 (N_2599,In_1765,In_1007);
nand U2600 (N_2600,In_2045,In_530);
nor U2601 (N_2601,In_176,In_1333);
nand U2602 (N_2602,In_2596,In_650);
and U2603 (N_2603,In_2849,In_587);
or U2604 (N_2604,In_127,In_2695);
or U2605 (N_2605,In_2073,In_54);
nand U2606 (N_2606,In_2926,In_1171);
nor U2607 (N_2607,In_2181,In_1472);
or U2608 (N_2608,In_971,In_107);
or U2609 (N_2609,In_2498,In_1838);
or U2610 (N_2610,In_963,In_83);
nor U2611 (N_2611,In_926,In_100);
nand U2612 (N_2612,In_916,In_1182);
or U2613 (N_2613,In_2436,In_2853);
xnor U2614 (N_2614,In_1103,In_209);
and U2615 (N_2615,In_249,In_614);
nor U2616 (N_2616,In_2682,In_2331);
and U2617 (N_2617,In_2427,In_1050);
nand U2618 (N_2618,In_458,In_241);
or U2619 (N_2619,In_1796,In_839);
nand U2620 (N_2620,In_538,In_1107);
nor U2621 (N_2621,In_2961,In_2423);
nor U2622 (N_2622,In_2322,In_2844);
and U2623 (N_2623,In_2401,In_2120);
nor U2624 (N_2624,In_1457,In_2877);
and U2625 (N_2625,In_1892,In_768);
and U2626 (N_2626,In_908,In_2693);
and U2627 (N_2627,In_2125,In_2210);
nand U2628 (N_2628,In_1881,In_1667);
nor U2629 (N_2629,In_2992,In_781);
nor U2630 (N_2630,In_2420,In_2138);
and U2631 (N_2631,In_264,In_2833);
or U2632 (N_2632,In_2673,In_2880);
and U2633 (N_2633,In_2437,In_1116);
nand U2634 (N_2634,In_835,In_2452);
or U2635 (N_2635,In_1958,In_2277);
nor U2636 (N_2636,In_1539,In_1549);
or U2637 (N_2637,In_1845,In_1161);
nand U2638 (N_2638,In_630,In_741);
nand U2639 (N_2639,In_2261,In_1528);
and U2640 (N_2640,In_563,In_704);
xnor U2641 (N_2641,In_941,In_663);
or U2642 (N_2642,In_560,In_2684);
or U2643 (N_2643,In_444,In_2854);
nor U2644 (N_2644,In_1258,In_2921);
nor U2645 (N_2645,In_742,In_2953);
nor U2646 (N_2646,In_589,In_677);
and U2647 (N_2647,In_1052,In_2079);
nand U2648 (N_2648,In_1699,In_922);
nand U2649 (N_2649,In_2763,In_1255);
nand U2650 (N_2650,In_2657,In_882);
nand U2651 (N_2651,In_2579,In_1799);
and U2652 (N_2652,In_2426,In_509);
nand U2653 (N_2653,In_895,In_1478);
or U2654 (N_2654,In_2874,In_1949);
xor U2655 (N_2655,In_783,In_915);
and U2656 (N_2656,In_720,In_611);
or U2657 (N_2657,In_520,In_1277);
nor U2658 (N_2658,In_1688,In_163);
nor U2659 (N_2659,In_1508,In_1693);
nand U2660 (N_2660,In_2021,In_276);
nand U2661 (N_2661,In_1879,In_1837);
and U2662 (N_2662,In_2700,In_1983);
nor U2663 (N_2663,In_2081,In_530);
or U2664 (N_2664,In_711,In_1823);
nor U2665 (N_2665,In_1553,In_2647);
and U2666 (N_2666,In_1287,In_892);
xnor U2667 (N_2667,In_847,In_125);
and U2668 (N_2668,In_1244,In_1617);
nor U2669 (N_2669,In_834,In_225);
and U2670 (N_2670,In_606,In_495);
nand U2671 (N_2671,In_2000,In_2653);
or U2672 (N_2672,In_1344,In_420);
nand U2673 (N_2673,In_1984,In_644);
nor U2674 (N_2674,In_2294,In_1650);
and U2675 (N_2675,In_22,In_223);
and U2676 (N_2676,In_523,In_2690);
nor U2677 (N_2677,In_893,In_2280);
nand U2678 (N_2678,In_2495,In_2796);
or U2679 (N_2679,In_1770,In_199);
or U2680 (N_2680,In_915,In_1390);
nand U2681 (N_2681,In_1735,In_2711);
nor U2682 (N_2682,In_901,In_1121);
or U2683 (N_2683,In_816,In_493);
or U2684 (N_2684,In_449,In_1793);
or U2685 (N_2685,In_1124,In_2511);
or U2686 (N_2686,In_2919,In_1623);
or U2687 (N_2687,In_998,In_1770);
nand U2688 (N_2688,In_368,In_555);
nor U2689 (N_2689,In_1113,In_1351);
or U2690 (N_2690,In_465,In_720);
nor U2691 (N_2691,In_884,In_2736);
and U2692 (N_2692,In_1772,In_335);
and U2693 (N_2693,In_71,In_2914);
nand U2694 (N_2694,In_258,In_841);
and U2695 (N_2695,In_2125,In_2042);
and U2696 (N_2696,In_2674,In_1041);
nand U2697 (N_2697,In_1154,In_2169);
or U2698 (N_2698,In_1847,In_2574);
nand U2699 (N_2699,In_2411,In_381);
and U2700 (N_2700,In_2605,In_1652);
nand U2701 (N_2701,In_1456,In_2236);
nor U2702 (N_2702,In_917,In_2106);
or U2703 (N_2703,In_2344,In_1098);
or U2704 (N_2704,In_505,In_1006);
nand U2705 (N_2705,In_1992,In_1401);
nor U2706 (N_2706,In_2913,In_115);
or U2707 (N_2707,In_810,In_449);
and U2708 (N_2708,In_331,In_857);
nand U2709 (N_2709,In_2139,In_1495);
nor U2710 (N_2710,In_92,In_386);
and U2711 (N_2711,In_1166,In_57);
and U2712 (N_2712,In_2076,In_2025);
or U2713 (N_2713,In_2675,In_2545);
and U2714 (N_2714,In_2899,In_1439);
nand U2715 (N_2715,In_1748,In_180);
nand U2716 (N_2716,In_2999,In_215);
nor U2717 (N_2717,In_2501,In_2617);
or U2718 (N_2718,In_1949,In_463);
and U2719 (N_2719,In_1482,In_1435);
nand U2720 (N_2720,In_852,In_1327);
nor U2721 (N_2721,In_1557,In_945);
and U2722 (N_2722,In_2795,In_782);
and U2723 (N_2723,In_564,In_1058);
and U2724 (N_2724,In_2875,In_259);
and U2725 (N_2725,In_1091,In_519);
or U2726 (N_2726,In_892,In_19);
and U2727 (N_2727,In_2627,In_70);
or U2728 (N_2728,In_2978,In_470);
or U2729 (N_2729,In_2605,In_1988);
nand U2730 (N_2730,In_2644,In_1863);
or U2731 (N_2731,In_1254,In_1172);
or U2732 (N_2732,In_1501,In_2934);
nand U2733 (N_2733,In_2995,In_784);
xor U2734 (N_2734,In_2731,In_1726);
nor U2735 (N_2735,In_2210,In_1767);
nand U2736 (N_2736,In_381,In_1014);
nand U2737 (N_2737,In_1591,In_75);
nand U2738 (N_2738,In_1362,In_1674);
nor U2739 (N_2739,In_63,In_1735);
and U2740 (N_2740,In_1356,In_1480);
nor U2741 (N_2741,In_191,In_2661);
nor U2742 (N_2742,In_2891,In_2185);
and U2743 (N_2743,In_1908,In_979);
and U2744 (N_2744,In_584,In_835);
and U2745 (N_2745,In_1128,In_2652);
and U2746 (N_2746,In_1114,In_2157);
and U2747 (N_2747,In_482,In_1207);
or U2748 (N_2748,In_2748,In_1013);
or U2749 (N_2749,In_2102,In_1128);
nand U2750 (N_2750,In_1278,In_93);
nand U2751 (N_2751,In_490,In_923);
and U2752 (N_2752,In_964,In_1922);
nor U2753 (N_2753,In_2410,In_2984);
nand U2754 (N_2754,In_1622,In_367);
and U2755 (N_2755,In_300,In_2168);
nor U2756 (N_2756,In_546,In_2955);
or U2757 (N_2757,In_2828,In_1349);
and U2758 (N_2758,In_2335,In_2865);
nor U2759 (N_2759,In_2141,In_1682);
nand U2760 (N_2760,In_1707,In_901);
nand U2761 (N_2761,In_2083,In_708);
and U2762 (N_2762,In_437,In_2303);
nor U2763 (N_2763,In_2638,In_2131);
nand U2764 (N_2764,In_631,In_1481);
or U2765 (N_2765,In_338,In_2900);
nor U2766 (N_2766,In_2554,In_824);
and U2767 (N_2767,In_860,In_2151);
nor U2768 (N_2768,In_1842,In_944);
nand U2769 (N_2769,In_228,In_1061);
nor U2770 (N_2770,In_1645,In_314);
nand U2771 (N_2771,In_2089,In_1520);
nor U2772 (N_2772,In_2221,In_1902);
and U2773 (N_2773,In_762,In_2545);
nand U2774 (N_2774,In_1434,In_2084);
and U2775 (N_2775,In_8,In_2697);
or U2776 (N_2776,In_2684,In_1746);
and U2777 (N_2777,In_525,In_1536);
nand U2778 (N_2778,In_1565,In_543);
nor U2779 (N_2779,In_155,In_2014);
and U2780 (N_2780,In_258,In_1966);
or U2781 (N_2781,In_1480,In_412);
and U2782 (N_2782,In_1268,In_272);
nand U2783 (N_2783,In_1438,In_1617);
and U2784 (N_2784,In_954,In_675);
nor U2785 (N_2785,In_28,In_127);
or U2786 (N_2786,In_1462,In_2706);
nor U2787 (N_2787,In_1263,In_711);
nor U2788 (N_2788,In_2993,In_2520);
nand U2789 (N_2789,In_1030,In_2408);
nand U2790 (N_2790,In_2381,In_2310);
nand U2791 (N_2791,In_648,In_69);
nor U2792 (N_2792,In_922,In_2530);
nor U2793 (N_2793,In_2980,In_2135);
nor U2794 (N_2794,In_1787,In_1801);
nor U2795 (N_2795,In_1082,In_2379);
or U2796 (N_2796,In_1240,In_2073);
nand U2797 (N_2797,In_278,In_1719);
and U2798 (N_2798,In_1844,In_1924);
nand U2799 (N_2799,In_706,In_1474);
or U2800 (N_2800,In_743,In_1276);
or U2801 (N_2801,In_1838,In_1126);
nand U2802 (N_2802,In_807,In_2180);
nor U2803 (N_2803,In_1401,In_270);
and U2804 (N_2804,In_282,In_2609);
nand U2805 (N_2805,In_91,In_2751);
nand U2806 (N_2806,In_1735,In_807);
nand U2807 (N_2807,In_1371,In_1743);
nand U2808 (N_2808,In_2256,In_1468);
nor U2809 (N_2809,In_1871,In_686);
nor U2810 (N_2810,In_1837,In_1851);
or U2811 (N_2811,In_132,In_2327);
and U2812 (N_2812,In_438,In_553);
nor U2813 (N_2813,In_1368,In_649);
nand U2814 (N_2814,In_822,In_2918);
nand U2815 (N_2815,In_1070,In_450);
nor U2816 (N_2816,In_216,In_2635);
and U2817 (N_2817,In_1339,In_1437);
nor U2818 (N_2818,In_1414,In_675);
nand U2819 (N_2819,In_2159,In_252);
or U2820 (N_2820,In_2287,In_407);
nor U2821 (N_2821,In_1741,In_607);
nor U2822 (N_2822,In_1530,In_198);
nor U2823 (N_2823,In_2294,In_2078);
or U2824 (N_2824,In_345,In_2237);
and U2825 (N_2825,In_2859,In_443);
and U2826 (N_2826,In_1719,In_1841);
nor U2827 (N_2827,In_958,In_1887);
nor U2828 (N_2828,In_828,In_935);
nand U2829 (N_2829,In_2724,In_76);
nor U2830 (N_2830,In_2733,In_955);
and U2831 (N_2831,In_2298,In_2178);
and U2832 (N_2832,In_1640,In_2638);
nand U2833 (N_2833,In_2499,In_220);
nor U2834 (N_2834,In_1438,In_797);
and U2835 (N_2835,In_571,In_538);
nor U2836 (N_2836,In_1515,In_1074);
or U2837 (N_2837,In_1487,In_1342);
and U2838 (N_2838,In_1947,In_2565);
nand U2839 (N_2839,In_2651,In_2756);
nor U2840 (N_2840,In_2613,In_2787);
and U2841 (N_2841,In_2124,In_307);
or U2842 (N_2842,In_1350,In_1299);
or U2843 (N_2843,In_447,In_1313);
and U2844 (N_2844,In_802,In_1813);
nand U2845 (N_2845,In_2918,In_1274);
nand U2846 (N_2846,In_2997,In_1306);
nand U2847 (N_2847,In_2353,In_1663);
or U2848 (N_2848,In_1608,In_265);
nor U2849 (N_2849,In_2452,In_528);
or U2850 (N_2850,In_2117,In_1242);
nor U2851 (N_2851,In_1405,In_2032);
and U2852 (N_2852,In_1428,In_2262);
or U2853 (N_2853,In_518,In_653);
nand U2854 (N_2854,In_2337,In_1763);
nor U2855 (N_2855,In_928,In_1964);
nor U2856 (N_2856,In_1006,In_1814);
or U2857 (N_2857,In_325,In_2313);
or U2858 (N_2858,In_2538,In_1220);
nor U2859 (N_2859,In_75,In_1963);
nand U2860 (N_2860,In_2754,In_758);
or U2861 (N_2861,In_133,In_1581);
xor U2862 (N_2862,In_1966,In_1841);
or U2863 (N_2863,In_1604,In_1612);
nor U2864 (N_2864,In_1147,In_2167);
nand U2865 (N_2865,In_1801,In_1044);
or U2866 (N_2866,In_896,In_1032);
nand U2867 (N_2867,In_630,In_1444);
xor U2868 (N_2868,In_1304,In_1114);
or U2869 (N_2869,In_1007,In_721);
and U2870 (N_2870,In_635,In_963);
nor U2871 (N_2871,In_1382,In_1133);
and U2872 (N_2872,In_476,In_694);
and U2873 (N_2873,In_313,In_492);
nand U2874 (N_2874,In_2876,In_1360);
nand U2875 (N_2875,In_204,In_2151);
and U2876 (N_2876,In_556,In_786);
nand U2877 (N_2877,In_1193,In_2924);
and U2878 (N_2878,In_2222,In_1440);
nor U2879 (N_2879,In_2761,In_267);
nand U2880 (N_2880,In_2908,In_2455);
nand U2881 (N_2881,In_547,In_2413);
or U2882 (N_2882,In_2545,In_118);
nand U2883 (N_2883,In_895,In_1983);
or U2884 (N_2884,In_173,In_2419);
or U2885 (N_2885,In_2818,In_2419);
nand U2886 (N_2886,In_208,In_2252);
nor U2887 (N_2887,In_2725,In_1830);
and U2888 (N_2888,In_35,In_756);
nand U2889 (N_2889,In_1191,In_1054);
nor U2890 (N_2890,In_960,In_1823);
nor U2891 (N_2891,In_2814,In_2128);
nor U2892 (N_2892,In_768,In_302);
and U2893 (N_2893,In_675,In_2764);
and U2894 (N_2894,In_1324,In_2026);
nor U2895 (N_2895,In_1152,In_1998);
nand U2896 (N_2896,In_1325,In_2072);
and U2897 (N_2897,In_1129,In_2743);
and U2898 (N_2898,In_1053,In_1590);
nand U2899 (N_2899,In_2264,In_1929);
and U2900 (N_2900,In_463,In_611);
nand U2901 (N_2901,In_1348,In_244);
nor U2902 (N_2902,In_2532,In_553);
nand U2903 (N_2903,In_116,In_1254);
nand U2904 (N_2904,In_296,In_361);
and U2905 (N_2905,In_492,In_1113);
nand U2906 (N_2906,In_2190,In_353);
nor U2907 (N_2907,In_150,In_308);
and U2908 (N_2908,In_2346,In_2830);
or U2909 (N_2909,In_2222,In_2450);
or U2910 (N_2910,In_243,In_2908);
nand U2911 (N_2911,In_2566,In_2370);
nand U2912 (N_2912,In_2771,In_1762);
and U2913 (N_2913,In_1209,In_2329);
and U2914 (N_2914,In_1835,In_641);
and U2915 (N_2915,In_863,In_1669);
nand U2916 (N_2916,In_769,In_1728);
nand U2917 (N_2917,In_1074,In_892);
nor U2918 (N_2918,In_435,In_2046);
nand U2919 (N_2919,In_124,In_1843);
and U2920 (N_2920,In_1845,In_1727);
nor U2921 (N_2921,In_2603,In_561);
nand U2922 (N_2922,In_1052,In_2650);
and U2923 (N_2923,In_2337,In_2084);
and U2924 (N_2924,In_229,In_1831);
xor U2925 (N_2925,In_2381,In_1009);
nand U2926 (N_2926,In_1638,In_935);
or U2927 (N_2927,In_2067,In_994);
and U2928 (N_2928,In_1534,In_2862);
and U2929 (N_2929,In_2204,In_2810);
nor U2930 (N_2930,In_472,In_1064);
nand U2931 (N_2931,In_95,In_611);
and U2932 (N_2932,In_2245,In_871);
and U2933 (N_2933,In_2272,In_478);
nor U2934 (N_2934,In_775,In_2189);
and U2935 (N_2935,In_210,In_2716);
nand U2936 (N_2936,In_200,In_2808);
nand U2937 (N_2937,In_2433,In_727);
nand U2938 (N_2938,In_441,In_1764);
nor U2939 (N_2939,In_784,In_2454);
and U2940 (N_2940,In_1174,In_201);
nand U2941 (N_2941,In_299,In_1207);
and U2942 (N_2942,In_2942,In_2716);
nor U2943 (N_2943,In_805,In_1932);
or U2944 (N_2944,In_598,In_2417);
nor U2945 (N_2945,In_2964,In_807);
nand U2946 (N_2946,In_1513,In_2461);
nor U2947 (N_2947,In_2672,In_1559);
or U2948 (N_2948,In_72,In_2406);
nor U2949 (N_2949,In_1763,In_1353);
nor U2950 (N_2950,In_1651,In_2026);
nor U2951 (N_2951,In_2300,In_1703);
nand U2952 (N_2952,In_1678,In_1473);
or U2953 (N_2953,In_1391,In_786);
or U2954 (N_2954,In_1747,In_333);
nor U2955 (N_2955,In_773,In_406);
or U2956 (N_2956,In_1855,In_2174);
and U2957 (N_2957,In_59,In_2997);
and U2958 (N_2958,In_505,In_1068);
xnor U2959 (N_2959,In_2122,In_2994);
or U2960 (N_2960,In_238,In_1177);
or U2961 (N_2961,In_2638,In_2056);
and U2962 (N_2962,In_956,In_965);
or U2963 (N_2963,In_1353,In_2079);
nand U2964 (N_2964,In_966,In_1655);
nor U2965 (N_2965,In_561,In_918);
nand U2966 (N_2966,In_813,In_454);
and U2967 (N_2967,In_667,In_1145);
or U2968 (N_2968,In_818,In_545);
xnor U2969 (N_2969,In_1181,In_177);
nor U2970 (N_2970,In_310,In_1925);
or U2971 (N_2971,In_1817,In_315);
nor U2972 (N_2972,In_789,In_1249);
nand U2973 (N_2973,In_1557,In_2702);
or U2974 (N_2974,In_1682,In_843);
nand U2975 (N_2975,In_1185,In_806);
nor U2976 (N_2976,In_1208,In_277);
or U2977 (N_2977,In_340,In_347);
or U2978 (N_2978,In_1015,In_2911);
and U2979 (N_2979,In_1582,In_107);
nand U2980 (N_2980,In_1255,In_2056);
or U2981 (N_2981,In_1503,In_2090);
nor U2982 (N_2982,In_1702,In_962);
or U2983 (N_2983,In_2329,In_2743);
and U2984 (N_2984,In_2362,In_272);
or U2985 (N_2985,In_490,In_507);
nand U2986 (N_2986,In_2181,In_2530);
nand U2987 (N_2987,In_174,In_252);
nor U2988 (N_2988,In_920,In_2738);
and U2989 (N_2989,In_2754,In_469);
and U2990 (N_2990,In_1289,In_1557);
or U2991 (N_2991,In_576,In_707);
and U2992 (N_2992,In_2429,In_2060);
nand U2993 (N_2993,In_2522,In_1171);
and U2994 (N_2994,In_2319,In_2271);
or U2995 (N_2995,In_2999,In_2327);
and U2996 (N_2996,In_2857,In_2962);
nor U2997 (N_2997,In_2509,In_1835);
nor U2998 (N_2998,In_2026,In_1433);
nor U2999 (N_2999,In_2212,In_804);
nor U3000 (N_3000,In_659,In_804);
or U3001 (N_3001,In_622,In_2555);
and U3002 (N_3002,In_1874,In_2623);
or U3003 (N_3003,In_2686,In_2767);
and U3004 (N_3004,In_2731,In_1677);
nor U3005 (N_3005,In_71,In_1726);
and U3006 (N_3006,In_420,In_285);
nor U3007 (N_3007,In_1610,In_2833);
nor U3008 (N_3008,In_1891,In_2524);
or U3009 (N_3009,In_539,In_2734);
and U3010 (N_3010,In_1675,In_2965);
nor U3011 (N_3011,In_1441,In_852);
nor U3012 (N_3012,In_514,In_1351);
xnor U3013 (N_3013,In_2921,In_1355);
and U3014 (N_3014,In_659,In_2089);
or U3015 (N_3015,In_235,In_846);
and U3016 (N_3016,In_2585,In_2027);
nor U3017 (N_3017,In_16,In_408);
and U3018 (N_3018,In_1222,In_1820);
and U3019 (N_3019,In_211,In_1212);
or U3020 (N_3020,In_2498,In_2275);
nor U3021 (N_3021,In_393,In_2971);
nor U3022 (N_3022,In_2900,In_1471);
or U3023 (N_3023,In_1805,In_184);
nor U3024 (N_3024,In_2086,In_2123);
nand U3025 (N_3025,In_2689,In_412);
nor U3026 (N_3026,In_2839,In_799);
and U3027 (N_3027,In_286,In_2724);
nor U3028 (N_3028,In_673,In_1139);
or U3029 (N_3029,In_1246,In_1061);
and U3030 (N_3030,In_2159,In_1665);
nor U3031 (N_3031,In_2404,In_1702);
nand U3032 (N_3032,In_835,In_2398);
nand U3033 (N_3033,In_744,In_777);
or U3034 (N_3034,In_2797,In_1551);
or U3035 (N_3035,In_392,In_2085);
and U3036 (N_3036,In_2602,In_512);
and U3037 (N_3037,In_2042,In_2111);
nor U3038 (N_3038,In_1767,In_449);
or U3039 (N_3039,In_2678,In_1435);
nand U3040 (N_3040,In_1777,In_1319);
nand U3041 (N_3041,In_1472,In_203);
nand U3042 (N_3042,In_789,In_2761);
nand U3043 (N_3043,In_1248,In_1890);
nor U3044 (N_3044,In_231,In_2247);
or U3045 (N_3045,In_2200,In_1520);
or U3046 (N_3046,In_1030,In_1969);
and U3047 (N_3047,In_977,In_2464);
or U3048 (N_3048,In_491,In_781);
nor U3049 (N_3049,In_1338,In_1137);
or U3050 (N_3050,In_560,In_2274);
or U3051 (N_3051,In_60,In_2594);
and U3052 (N_3052,In_1650,In_2623);
nor U3053 (N_3053,In_2494,In_2392);
nor U3054 (N_3054,In_1368,In_170);
nand U3055 (N_3055,In_2006,In_2719);
nand U3056 (N_3056,In_1965,In_2787);
or U3057 (N_3057,In_2667,In_2539);
nand U3058 (N_3058,In_2109,In_1701);
nand U3059 (N_3059,In_2011,In_2000);
nand U3060 (N_3060,In_2728,In_1395);
or U3061 (N_3061,In_657,In_2431);
nand U3062 (N_3062,In_589,In_974);
nor U3063 (N_3063,In_1111,In_1855);
nand U3064 (N_3064,In_1455,In_124);
and U3065 (N_3065,In_2330,In_1362);
or U3066 (N_3066,In_65,In_2089);
or U3067 (N_3067,In_933,In_1174);
and U3068 (N_3068,In_2243,In_1084);
nand U3069 (N_3069,In_1332,In_2201);
or U3070 (N_3070,In_2149,In_2459);
or U3071 (N_3071,In_276,In_148);
or U3072 (N_3072,In_852,In_1099);
and U3073 (N_3073,In_2892,In_103);
or U3074 (N_3074,In_351,In_1546);
nand U3075 (N_3075,In_1197,In_2026);
or U3076 (N_3076,In_1452,In_957);
xor U3077 (N_3077,In_887,In_913);
and U3078 (N_3078,In_1122,In_1417);
nor U3079 (N_3079,In_2985,In_89);
nand U3080 (N_3080,In_322,In_2793);
and U3081 (N_3081,In_765,In_1938);
xnor U3082 (N_3082,In_1226,In_2167);
nand U3083 (N_3083,In_1204,In_2319);
nand U3084 (N_3084,In_2969,In_25);
nor U3085 (N_3085,In_230,In_2734);
or U3086 (N_3086,In_845,In_2394);
nor U3087 (N_3087,In_440,In_380);
nand U3088 (N_3088,In_1482,In_2913);
and U3089 (N_3089,In_2289,In_1047);
and U3090 (N_3090,In_1140,In_2151);
nand U3091 (N_3091,In_412,In_138);
nor U3092 (N_3092,In_2195,In_1673);
or U3093 (N_3093,In_2077,In_753);
and U3094 (N_3094,In_1469,In_1470);
nor U3095 (N_3095,In_592,In_978);
nor U3096 (N_3096,In_2547,In_2890);
or U3097 (N_3097,In_564,In_2761);
and U3098 (N_3098,In_669,In_1396);
xor U3099 (N_3099,In_373,In_1191);
nand U3100 (N_3100,In_1004,In_2986);
or U3101 (N_3101,In_285,In_2676);
and U3102 (N_3102,In_1392,In_2866);
nand U3103 (N_3103,In_5,In_1137);
or U3104 (N_3104,In_414,In_2704);
nand U3105 (N_3105,In_2486,In_1376);
or U3106 (N_3106,In_882,In_1483);
nand U3107 (N_3107,In_988,In_396);
nor U3108 (N_3108,In_2243,In_1659);
or U3109 (N_3109,In_2287,In_2902);
nand U3110 (N_3110,In_2644,In_2729);
and U3111 (N_3111,In_2771,In_1139);
nand U3112 (N_3112,In_909,In_549);
or U3113 (N_3113,In_2599,In_1674);
nor U3114 (N_3114,In_2043,In_2984);
or U3115 (N_3115,In_1258,In_201);
and U3116 (N_3116,In_1942,In_2407);
nand U3117 (N_3117,In_1620,In_2077);
nand U3118 (N_3118,In_2844,In_2189);
or U3119 (N_3119,In_1009,In_2756);
and U3120 (N_3120,In_1736,In_2282);
or U3121 (N_3121,In_470,In_911);
or U3122 (N_3122,In_1867,In_2745);
xnor U3123 (N_3123,In_2585,In_2002);
or U3124 (N_3124,In_713,In_500);
nor U3125 (N_3125,In_1993,In_2438);
nand U3126 (N_3126,In_2263,In_2180);
or U3127 (N_3127,In_2591,In_1366);
and U3128 (N_3128,In_860,In_289);
nand U3129 (N_3129,In_318,In_468);
or U3130 (N_3130,In_1507,In_1499);
and U3131 (N_3131,In_728,In_827);
or U3132 (N_3132,In_790,In_2996);
and U3133 (N_3133,In_417,In_2367);
or U3134 (N_3134,In_793,In_690);
and U3135 (N_3135,In_987,In_1676);
nand U3136 (N_3136,In_98,In_2561);
nand U3137 (N_3137,In_1191,In_588);
nand U3138 (N_3138,In_1025,In_2385);
or U3139 (N_3139,In_2919,In_35);
or U3140 (N_3140,In_2116,In_804);
and U3141 (N_3141,In_106,In_486);
nor U3142 (N_3142,In_711,In_2034);
or U3143 (N_3143,In_335,In_228);
nand U3144 (N_3144,In_1441,In_881);
nor U3145 (N_3145,In_388,In_2682);
nand U3146 (N_3146,In_2389,In_389);
nand U3147 (N_3147,In_2729,In_751);
nor U3148 (N_3148,In_518,In_779);
nor U3149 (N_3149,In_1415,In_929);
and U3150 (N_3150,In_1465,In_1238);
and U3151 (N_3151,In_2160,In_367);
nand U3152 (N_3152,In_1462,In_2870);
nand U3153 (N_3153,In_1611,In_1725);
nand U3154 (N_3154,In_1165,In_2849);
nand U3155 (N_3155,In_1134,In_1282);
or U3156 (N_3156,In_1920,In_1580);
nor U3157 (N_3157,In_2837,In_275);
nand U3158 (N_3158,In_2740,In_2315);
nand U3159 (N_3159,In_659,In_928);
nor U3160 (N_3160,In_43,In_311);
nand U3161 (N_3161,In_110,In_1105);
or U3162 (N_3162,In_961,In_2407);
nor U3163 (N_3163,In_2151,In_2563);
and U3164 (N_3164,In_257,In_2556);
nand U3165 (N_3165,In_1513,In_1347);
nand U3166 (N_3166,In_453,In_2832);
xnor U3167 (N_3167,In_2323,In_2317);
nor U3168 (N_3168,In_368,In_492);
nand U3169 (N_3169,In_2429,In_1195);
and U3170 (N_3170,In_851,In_1919);
and U3171 (N_3171,In_1896,In_1861);
nor U3172 (N_3172,In_86,In_1187);
nor U3173 (N_3173,In_402,In_415);
nand U3174 (N_3174,In_217,In_2216);
or U3175 (N_3175,In_918,In_197);
or U3176 (N_3176,In_2895,In_664);
or U3177 (N_3177,In_1693,In_2993);
nand U3178 (N_3178,In_138,In_297);
or U3179 (N_3179,In_1102,In_2289);
nand U3180 (N_3180,In_1798,In_447);
and U3181 (N_3181,In_1367,In_1534);
nand U3182 (N_3182,In_534,In_2378);
nor U3183 (N_3183,In_303,In_1671);
nand U3184 (N_3184,In_1111,In_97);
or U3185 (N_3185,In_716,In_1405);
and U3186 (N_3186,In_1121,In_1005);
nand U3187 (N_3187,In_1596,In_956);
nor U3188 (N_3188,In_1867,In_609);
or U3189 (N_3189,In_2013,In_2149);
or U3190 (N_3190,In_1381,In_1970);
and U3191 (N_3191,In_236,In_81);
nor U3192 (N_3192,In_445,In_610);
or U3193 (N_3193,In_29,In_587);
nand U3194 (N_3194,In_768,In_1343);
nand U3195 (N_3195,In_2125,In_1641);
and U3196 (N_3196,In_434,In_1095);
and U3197 (N_3197,In_2727,In_1712);
or U3198 (N_3198,In_647,In_1681);
nor U3199 (N_3199,In_1018,In_1360);
or U3200 (N_3200,In_2016,In_810);
or U3201 (N_3201,In_1076,In_939);
and U3202 (N_3202,In_2087,In_897);
and U3203 (N_3203,In_801,In_2755);
nand U3204 (N_3204,In_2354,In_340);
and U3205 (N_3205,In_2887,In_928);
or U3206 (N_3206,In_1404,In_2181);
and U3207 (N_3207,In_992,In_2472);
nand U3208 (N_3208,In_1759,In_2155);
nor U3209 (N_3209,In_18,In_456);
and U3210 (N_3210,In_1563,In_479);
nand U3211 (N_3211,In_1114,In_1574);
and U3212 (N_3212,In_687,In_2043);
nor U3213 (N_3213,In_977,In_406);
or U3214 (N_3214,In_81,In_2350);
nor U3215 (N_3215,In_2531,In_2427);
or U3216 (N_3216,In_2257,In_2278);
nor U3217 (N_3217,In_1840,In_365);
nor U3218 (N_3218,In_1704,In_946);
or U3219 (N_3219,In_228,In_146);
nand U3220 (N_3220,In_1718,In_1141);
and U3221 (N_3221,In_1258,In_148);
and U3222 (N_3222,In_717,In_1474);
or U3223 (N_3223,In_895,In_95);
and U3224 (N_3224,In_483,In_405);
or U3225 (N_3225,In_897,In_2349);
nor U3226 (N_3226,In_2284,In_179);
and U3227 (N_3227,In_2383,In_2231);
nor U3228 (N_3228,In_211,In_1376);
or U3229 (N_3229,In_96,In_2716);
nand U3230 (N_3230,In_541,In_1340);
nand U3231 (N_3231,In_1334,In_875);
or U3232 (N_3232,In_1484,In_254);
or U3233 (N_3233,In_2811,In_2346);
or U3234 (N_3234,In_2693,In_489);
and U3235 (N_3235,In_2435,In_1981);
or U3236 (N_3236,In_1024,In_1955);
nand U3237 (N_3237,In_2464,In_1387);
and U3238 (N_3238,In_1173,In_2954);
nor U3239 (N_3239,In_1851,In_1768);
nand U3240 (N_3240,In_1747,In_667);
and U3241 (N_3241,In_1403,In_242);
nand U3242 (N_3242,In_680,In_831);
nand U3243 (N_3243,In_1440,In_678);
nor U3244 (N_3244,In_2940,In_1012);
nor U3245 (N_3245,In_2687,In_1935);
nand U3246 (N_3246,In_2021,In_1148);
or U3247 (N_3247,In_2870,In_2574);
nand U3248 (N_3248,In_137,In_732);
nand U3249 (N_3249,In_298,In_2670);
nand U3250 (N_3250,In_1167,In_2592);
nand U3251 (N_3251,In_204,In_2978);
nor U3252 (N_3252,In_2403,In_1164);
nor U3253 (N_3253,In_527,In_2644);
nor U3254 (N_3254,In_2052,In_1829);
or U3255 (N_3255,In_2071,In_1559);
nand U3256 (N_3256,In_1926,In_2344);
nand U3257 (N_3257,In_1464,In_2547);
nand U3258 (N_3258,In_921,In_959);
and U3259 (N_3259,In_2967,In_1912);
nand U3260 (N_3260,In_1499,In_971);
nor U3261 (N_3261,In_1900,In_2746);
nor U3262 (N_3262,In_2776,In_21);
and U3263 (N_3263,In_315,In_2074);
and U3264 (N_3264,In_2730,In_94);
or U3265 (N_3265,In_2859,In_1694);
or U3266 (N_3266,In_188,In_2289);
nor U3267 (N_3267,In_378,In_1517);
and U3268 (N_3268,In_2534,In_1576);
and U3269 (N_3269,In_211,In_1079);
nand U3270 (N_3270,In_630,In_427);
nand U3271 (N_3271,In_1145,In_1803);
or U3272 (N_3272,In_538,In_1052);
and U3273 (N_3273,In_979,In_1980);
and U3274 (N_3274,In_992,In_1350);
or U3275 (N_3275,In_2031,In_1074);
or U3276 (N_3276,In_106,In_2624);
nand U3277 (N_3277,In_2490,In_107);
and U3278 (N_3278,In_2003,In_1571);
nor U3279 (N_3279,In_2052,In_2932);
nand U3280 (N_3280,In_2592,In_1477);
or U3281 (N_3281,In_869,In_2186);
nor U3282 (N_3282,In_139,In_1425);
or U3283 (N_3283,In_2551,In_2122);
or U3284 (N_3284,In_2793,In_2866);
and U3285 (N_3285,In_1254,In_2517);
or U3286 (N_3286,In_2693,In_2690);
nor U3287 (N_3287,In_648,In_540);
and U3288 (N_3288,In_1783,In_1970);
nand U3289 (N_3289,In_1113,In_2130);
nand U3290 (N_3290,In_2952,In_949);
nand U3291 (N_3291,In_625,In_1313);
nor U3292 (N_3292,In_2837,In_2172);
nand U3293 (N_3293,In_1257,In_2429);
and U3294 (N_3294,In_800,In_363);
nand U3295 (N_3295,In_1831,In_17);
and U3296 (N_3296,In_1308,In_622);
and U3297 (N_3297,In_142,In_209);
and U3298 (N_3298,In_2953,In_1354);
nor U3299 (N_3299,In_2528,In_186);
and U3300 (N_3300,In_386,In_1611);
nand U3301 (N_3301,In_743,In_966);
or U3302 (N_3302,In_2331,In_2311);
and U3303 (N_3303,In_101,In_2099);
nor U3304 (N_3304,In_1613,In_486);
or U3305 (N_3305,In_1716,In_284);
nand U3306 (N_3306,In_534,In_1943);
or U3307 (N_3307,In_2805,In_1875);
or U3308 (N_3308,In_879,In_1633);
nor U3309 (N_3309,In_585,In_1909);
nand U3310 (N_3310,In_948,In_418);
or U3311 (N_3311,In_2951,In_873);
nand U3312 (N_3312,In_684,In_1337);
nor U3313 (N_3313,In_575,In_887);
nor U3314 (N_3314,In_1580,In_496);
and U3315 (N_3315,In_205,In_2629);
and U3316 (N_3316,In_775,In_891);
or U3317 (N_3317,In_2388,In_573);
and U3318 (N_3318,In_809,In_2076);
or U3319 (N_3319,In_2230,In_520);
nand U3320 (N_3320,In_59,In_427);
nor U3321 (N_3321,In_134,In_2698);
or U3322 (N_3322,In_1708,In_2196);
nand U3323 (N_3323,In_418,In_1332);
and U3324 (N_3324,In_1520,In_1142);
nand U3325 (N_3325,In_158,In_43);
nand U3326 (N_3326,In_1475,In_830);
and U3327 (N_3327,In_2600,In_2576);
and U3328 (N_3328,In_1107,In_267);
or U3329 (N_3329,In_1256,In_1204);
nor U3330 (N_3330,In_1449,In_455);
nand U3331 (N_3331,In_1772,In_1751);
and U3332 (N_3332,In_906,In_1824);
nand U3333 (N_3333,In_1124,In_711);
nor U3334 (N_3334,In_1806,In_2463);
or U3335 (N_3335,In_1292,In_2407);
or U3336 (N_3336,In_987,In_820);
and U3337 (N_3337,In_2886,In_1979);
and U3338 (N_3338,In_1141,In_594);
nor U3339 (N_3339,In_1671,In_2577);
nor U3340 (N_3340,In_1663,In_179);
and U3341 (N_3341,In_1888,In_1150);
nand U3342 (N_3342,In_2569,In_2279);
nand U3343 (N_3343,In_97,In_1172);
nor U3344 (N_3344,In_1020,In_581);
or U3345 (N_3345,In_2341,In_1483);
or U3346 (N_3346,In_371,In_82);
and U3347 (N_3347,In_722,In_2328);
and U3348 (N_3348,In_215,In_1374);
nor U3349 (N_3349,In_2840,In_2271);
or U3350 (N_3350,In_789,In_930);
xor U3351 (N_3351,In_749,In_1187);
nand U3352 (N_3352,In_1510,In_2932);
nand U3353 (N_3353,In_2246,In_2075);
and U3354 (N_3354,In_1427,In_1003);
or U3355 (N_3355,In_692,In_1481);
or U3356 (N_3356,In_2865,In_802);
nor U3357 (N_3357,In_834,In_731);
and U3358 (N_3358,In_1381,In_2806);
nor U3359 (N_3359,In_2747,In_1689);
nor U3360 (N_3360,In_2880,In_2158);
and U3361 (N_3361,In_2949,In_1905);
or U3362 (N_3362,In_2486,In_1299);
or U3363 (N_3363,In_1638,In_1716);
or U3364 (N_3364,In_443,In_0);
and U3365 (N_3365,In_2577,In_505);
nor U3366 (N_3366,In_2742,In_2772);
nand U3367 (N_3367,In_2520,In_602);
xor U3368 (N_3368,In_2802,In_2999);
nor U3369 (N_3369,In_369,In_212);
nor U3370 (N_3370,In_429,In_1399);
or U3371 (N_3371,In_583,In_2327);
nor U3372 (N_3372,In_2821,In_2466);
nand U3373 (N_3373,In_606,In_2193);
or U3374 (N_3374,In_170,In_2663);
and U3375 (N_3375,In_2990,In_24);
and U3376 (N_3376,In_2690,In_1049);
and U3377 (N_3377,In_1801,In_2158);
and U3378 (N_3378,In_1665,In_2176);
nor U3379 (N_3379,In_2674,In_2289);
and U3380 (N_3380,In_2445,In_1076);
and U3381 (N_3381,In_805,In_1551);
and U3382 (N_3382,In_1592,In_2826);
nor U3383 (N_3383,In_1308,In_2907);
or U3384 (N_3384,In_2069,In_1237);
nor U3385 (N_3385,In_2263,In_611);
and U3386 (N_3386,In_2434,In_2208);
and U3387 (N_3387,In_945,In_2966);
and U3388 (N_3388,In_784,In_340);
nor U3389 (N_3389,In_2202,In_39);
nand U3390 (N_3390,In_2655,In_260);
or U3391 (N_3391,In_2829,In_1653);
nor U3392 (N_3392,In_353,In_1998);
nor U3393 (N_3393,In_858,In_870);
or U3394 (N_3394,In_801,In_2729);
nor U3395 (N_3395,In_1025,In_1733);
nor U3396 (N_3396,In_1865,In_203);
nand U3397 (N_3397,In_2088,In_1207);
or U3398 (N_3398,In_1081,In_1413);
or U3399 (N_3399,In_280,In_462);
and U3400 (N_3400,In_623,In_1523);
and U3401 (N_3401,In_2867,In_2793);
and U3402 (N_3402,In_544,In_454);
nor U3403 (N_3403,In_579,In_974);
and U3404 (N_3404,In_1634,In_1218);
xnor U3405 (N_3405,In_2412,In_1908);
nor U3406 (N_3406,In_615,In_128);
nor U3407 (N_3407,In_991,In_1343);
nand U3408 (N_3408,In_1397,In_2263);
or U3409 (N_3409,In_1180,In_1727);
or U3410 (N_3410,In_152,In_965);
or U3411 (N_3411,In_2775,In_834);
and U3412 (N_3412,In_2483,In_866);
and U3413 (N_3413,In_2877,In_2189);
and U3414 (N_3414,In_1611,In_77);
and U3415 (N_3415,In_644,In_1829);
nor U3416 (N_3416,In_1161,In_2411);
nor U3417 (N_3417,In_118,In_2750);
and U3418 (N_3418,In_543,In_1464);
and U3419 (N_3419,In_2797,In_1016);
or U3420 (N_3420,In_1760,In_2003);
nor U3421 (N_3421,In_678,In_1234);
nand U3422 (N_3422,In_2405,In_1281);
and U3423 (N_3423,In_990,In_1992);
nor U3424 (N_3424,In_401,In_2691);
and U3425 (N_3425,In_1650,In_125);
and U3426 (N_3426,In_461,In_33);
or U3427 (N_3427,In_438,In_86);
or U3428 (N_3428,In_1270,In_2165);
nand U3429 (N_3429,In_327,In_950);
or U3430 (N_3430,In_2041,In_2639);
or U3431 (N_3431,In_1515,In_394);
and U3432 (N_3432,In_2597,In_2823);
or U3433 (N_3433,In_1568,In_781);
nor U3434 (N_3434,In_2729,In_2504);
nor U3435 (N_3435,In_1565,In_1571);
nor U3436 (N_3436,In_1338,In_333);
nand U3437 (N_3437,In_1087,In_1213);
nand U3438 (N_3438,In_590,In_1463);
or U3439 (N_3439,In_2531,In_254);
or U3440 (N_3440,In_1651,In_1435);
nor U3441 (N_3441,In_2889,In_2670);
or U3442 (N_3442,In_928,In_255);
or U3443 (N_3443,In_2965,In_2736);
nor U3444 (N_3444,In_2926,In_1256);
or U3445 (N_3445,In_1890,In_1027);
nor U3446 (N_3446,In_1208,In_2666);
nand U3447 (N_3447,In_553,In_2107);
nand U3448 (N_3448,In_223,In_534);
or U3449 (N_3449,In_318,In_2794);
nand U3450 (N_3450,In_2822,In_903);
nor U3451 (N_3451,In_234,In_2433);
nand U3452 (N_3452,In_693,In_2857);
nor U3453 (N_3453,In_2472,In_650);
nand U3454 (N_3454,In_1735,In_198);
or U3455 (N_3455,In_518,In_1834);
nor U3456 (N_3456,In_564,In_1002);
nor U3457 (N_3457,In_1399,In_2026);
or U3458 (N_3458,In_2288,In_2406);
nor U3459 (N_3459,In_343,In_850);
nand U3460 (N_3460,In_1393,In_550);
and U3461 (N_3461,In_473,In_1419);
and U3462 (N_3462,In_243,In_2712);
nand U3463 (N_3463,In_2019,In_1832);
nand U3464 (N_3464,In_1986,In_2574);
or U3465 (N_3465,In_743,In_1857);
or U3466 (N_3466,In_412,In_1392);
nor U3467 (N_3467,In_2525,In_81);
or U3468 (N_3468,In_2528,In_495);
and U3469 (N_3469,In_507,In_1437);
or U3470 (N_3470,In_1706,In_899);
nor U3471 (N_3471,In_1136,In_1990);
nand U3472 (N_3472,In_2550,In_2256);
nor U3473 (N_3473,In_2310,In_198);
nand U3474 (N_3474,In_1491,In_2261);
nor U3475 (N_3475,In_656,In_1873);
or U3476 (N_3476,In_1460,In_370);
and U3477 (N_3477,In_834,In_2880);
xnor U3478 (N_3478,In_2388,In_1305);
nor U3479 (N_3479,In_1046,In_312);
nand U3480 (N_3480,In_2610,In_1018);
nor U3481 (N_3481,In_396,In_30);
nand U3482 (N_3482,In_2672,In_2760);
nor U3483 (N_3483,In_1402,In_434);
and U3484 (N_3484,In_586,In_1776);
nand U3485 (N_3485,In_267,In_75);
and U3486 (N_3486,In_2670,In_457);
and U3487 (N_3487,In_40,In_308);
and U3488 (N_3488,In_618,In_2180);
nand U3489 (N_3489,In_2756,In_1947);
nor U3490 (N_3490,In_1227,In_1493);
nand U3491 (N_3491,In_636,In_1174);
and U3492 (N_3492,In_927,In_2936);
and U3493 (N_3493,In_507,In_2770);
and U3494 (N_3494,In_1170,In_183);
or U3495 (N_3495,In_1894,In_1856);
nor U3496 (N_3496,In_1847,In_556);
or U3497 (N_3497,In_2359,In_557);
or U3498 (N_3498,In_1805,In_850);
nand U3499 (N_3499,In_1832,In_2624);
nand U3500 (N_3500,In_2478,In_2606);
nor U3501 (N_3501,In_1422,In_1307);
nand U3502 (N_3502,In_1251,In_639);
nor U3503 (N_3503,In_2045,In_2456);
nand U3504 (N_3504,In_1497,In_2516);
and U3505 (N_3505,In_1821,In_1563);
and U3506 (N_3506,In_310,In_922);
or U3507 (N_3507,In_1795,In_1764);
nor U3508 (N_3508,In_1772,In_748);
or U3509 (N_3509,In_2793,In_1328);
or U3510 (N_3510,In_1018,In_1582);
or U3511 (N_3511,In_276,In_410);
nor U3512 (N_3512,In_2609,In_2834);
or U3513 (N_3513,In_909,In_1944);
nor U3514 (N_3514,In_2527,In_1027);
or U3515 (N_3515,In_1668,In_803);
and U3516 (N_3516,In_1003,In_2634);
nor U3517 (N_3517,In_1881,In_2997);
nand U3518 (N_3518,In_2979,In_2748);
or U3519 (N_3519,In_2710,In_962);
xor U3520 (N_3520,In_1816,In_2527);
nor U3521 (N_3521,In_1086,In_1649);
and U3522 (N_3522,In_1767,In_1321);
nand U3523 (N_3523,In_426,In_2861);
nand U3524 (N_3524,In_54,In_2256);
nor U3525 (N_3525,In_2707,In_2679);
or U3526 (N_3526,In_780,In_1748);
nor U3527 (N_3527,In_422,In_2123);
or U3528 (N_3528,In_2987,In_2524);
nor U3529 (N_3529,In_2349,In_2690);
or U3530 (N_3530,In_2097,In_2488);
nor U3531 (N_3531,In_563,In_774);
nand U3532 (N_3532,In_1182,In_2620);
nor U3533 (N_3533,In_682,In_92);
nand U3534 (N_3534,In_2005,In_2377);
or U3535 (N_3535,In_2348,In_1004);
or U3536 (N_3536,In_2699,In_1804);
xnor U3537 (N_3537,In_1976,In_673);
nor U3538 (N_3538,In_2844,In_2836);
nor U3539 (N_3539,In_2223,In_2893);
or U3540 (N_3540,In_2938,In_2912);
or U3541 (N_3541,In_2502,In_1008);
or U3542 (N_3542,In_1706,In_21);
nor U3543 (N_3543,In_839,In_2285);
and U3544 (N_3544,In_108,In_1513);
or U3545 (N_3545,In_807,In_727);
nor U3546 (N_3546,In_2307,In_2484);
nand U3547 (N_3547,In_1534,In_2389);
nor U3548 (N_3548,In_2017,In_1483);
and U3549 (N_3549,In_760,In_2598);
or U3550 (N_3550,In_84,In_2888);
nand U3551 (N_3551,In_1721,In_1204);
and U3552 (N_3552,In_704,In_156);
nor U3553 (N_3553,In_399,In_2355);
and U3554 (N_3554,In_861,In_573);
or U3555 (N_3555,In_1036,In_2159);
or U3556 (N_3556,In_2191,In_229);
nor U3557 (N_3557,In_2981,In_1566);
or U3558 (N_3558,In_902,In_1806);
nor U3559 (N_3559,In_501,In_544);
nand U3560 (N_3560,In_421,In_2559);
and U3561 (N_3561,In_970,In_2629);
and U3562 (N_3562,In_1194,In_1602);
and U3563 (N_3563,In_2965,In_2091);
nand U3564 (N_3564,In_844,In_2011);
or U3565 (N_3565,In_2342,In_2837);
nand U3566 (N_3566,In_782,In_621);
and U3567 (N_3567,In_488,In_2497);
nor U3568 (N_3568,In_723,In_453);
nand U3569 (N_3569,In_1737,In_1730);
and U3570 (N_3570,In_2930,In_2227);
or U3571 (N_3571,In_2407,In_2697);
nor U3572 (N_3572,In_627,In_2476);
nor U3573 (N_3573,In_2918,In_1300);
nand U3574 (N_3574,In_2452,In_1014);
and U3575 (N_3575,In_292,In_817);
and U3576 (N_3576,In_416,In_2143);
nand U3577 (N_3577,In_814,In_2752);
nand U3578 (N_3578,In_2423,In_2796);
and U3579 (N_3579,In_212,In_2288);
or U3580 (N_3580,In_340,In_654);
nand U3581 (N_3581,In_2610,In_924);
and U3582 (N_3582,In_775,In_2985);
or U3583 (N_3583,In_1297,In_2787);
nand U3584 (N_3584,In_568,In_678);
and U3585 (N_3585,In_1806,In_2533);
nand U3586 (N_3586,In_1996,In_2507);
nor U3587 (N_3587,In_749,In_299);
and U3588 (N_3588,In_1098,In_2628);
and U3589 (N_3589,In_358,In_2752);
nand U3590 (N_3590,In_1479,In_2437);
or U3591 (N_3591,In_402,In_1481);
nor U3592 (N_3592,In_1873,In_1044);
nand U3593 (N_3593,In_1891,In_71);
and U3594 (N_3594,In_1044,In_948);
nand U3595 (N_3595,In_1357,In_1597);
nor U3596 (N_3596,In_529,In_1596);
and U3597 (N_3597,In_422,In_2460);
nand U3598 (N_3598,In_2710,In_1708);
or U3599 (N_3599,In_2950,In_1648);
and U3600 (N_3600,In_207,In_2631);
or U3601 (N_3601,In_1646,In_2649);
and U3602 (N_3602,In_1307,In_1131);
nor U3603 (N_3603,In_1611,In_1346);
nand U3604 (N_3604,In_1991,In_2409);
or U3605 (N_3605,In_2020,In_1110);
or U3606 (N_3606,In_2068,In_1077);
and U3607 (N_3607,In_2260,In_134);
nor U3608 (N_3608,In_1447,In_1746);
nor U3609 (N_3609,In_1509,In_423);
and U3610 (N_3610,In_2393,In_1260);
or U3611 (N_3611,In_1104,In_1328);
nor U3612 (N_3612,In_1100,In_1716);
nand U3613 (N_3613,In_2583,In_2736);
nand U3614 (N_3614,In_2767,In_800);
nand U3615 (N_3615,In_838,In_650);
or U3616 (N_3616,In_1548,In_1389);
nand U3617 (N_3617,In_711,In_379);
or U3618 (N_3618,In_2446,In_2807);
and U3619 (N_3619,In_1062,In_1217);
nor U3620 (N_3620,In_259,In_2051);
and U3621 (N_3621,In_2351,In_2167);
and U3622 (N_3622,In_2377,In_813);
or U3623 (N_3623,In_1073,In_858);
or U3624 (N_3624,In_809,In_649);
nor U3625 (N_3625,In_2881,In_259);
or U3626 (N_3626,In_385,In_2141);
or U3627 (N_3627,In_2918,In_1866);
nor U3628 (N_3628,In_658,In_2496);
and U3629 (N_3629,In_1341,In_2220);
and U3630 (N_3630,In_365,In_2667);
and U3631 (N_3631,In_1718,In_2920);
nand U3632 (N_3632,In_2493,In_1081);
and U3633 (N_3633,In_2052,In_2252);
and U3634 (N_3634,In_2333,In_1300);
or U3635 (N_3635,In_1037,In_21);
or U3636 (N_3636,In_1936,In_2987);
and U3637 (N_3637,In_2788,In_822);
and U3638 (N_3638,In_1615,In_1961);
nor U3639 (N_3639,In_2144,In_320);
and U3640 (N_3640,In_141,In_1459);
nand U3641 (N_3641,In_1256,In_1459);
and U3642 (N_3642,In_687,In_1494);
or U3643 (N_3643,In_497,In_1177);
and U3644 (N_3644,In_826,In_52);
nand U3645 (N_3645,In_265,In_1007);
and U3646 (N_3646,In_2329,In_2885);
or U3647 (N_3647,In_375,In_1831);
nand U3648 (N_3648,In_30,In_1301);
xor U3649 (N_3649,In_2755,In_291);
nand U3650 (N_3650,In_2713,In_1652);
or U3651 (N_3651,In_739,In_2451);
xor U3652 (N_3652,In_2921,In_1930);
nand U3653 (N_3653,In_2042,In_410);
or U3654 (N_3654,In_2784,In_570);
nand U3655 (N_3655,In_1119,In_2813);
or U3656 (N_3656,In_2778,In_982);
or U3657 (N_3657,In_2426,In_2301);
and U3658 (N_3658,In_736,In_1591);
nor U3659 (N_3659,In_459,In_819);
nand U3660 (N_3660,In_2019,In_17);
and U3661 (N_3661,In_2396,In_2492);
and U3662 (N_3662,In_2745,In_1556);
nor U3663 (N_3663,In_2286,In_2089);
and U3664 (N_3664,In_1297,In_1354);
and U3665 (N_3665,In_725,In_8);
and U3666 (N_3666,In_726,In_2028);
or U3667 (N_3667,In_2018,In_968);
nand U3668 (N_3668,In_2211,In_1474);
nor U3669 (N_3669,In_1948,In_1490);
or U3670 (N_3670,In_1267,In_833);
or U3671 (N_3671,In_849,In_1495);
nand U3672 (N_3672,In_2764,In_23);
or U3673 (N_3673,In_1743,In_1782);
and U3674 (N_3674,In_476,In_2423);
and U3675 (N_3675,In_2334,In_1958);
nor U3676 (N_3676,In_2266,In_991);
nand U3677 (N_3677,In_1606,In_1179);
or U3678 (N_3678,In_2780,In_2167);
nand U3679 (N_3679,In_1045,In_1420);
and U3680 (N_3680,In_1169,In_2813);
nand U3681 (N_3681,In_109,In_942);
nand U3682 (N_3682,In_302,In_2547);
and U3683 (N_3683,In_2653,In_2811);
nand U3684 (N_3684,In_751,In_33);
nand U3685 (N_3685,In_511,In_2295);
nor U3686 (N_3686,In_223,In_309);
nand U3687 (N_3687,In_173,In_746);
and U3688 (N_3688,In_1139,In_2611);
nor U3689 (N_3689,In_2488,In_1788);
nor U3690 (N_3690,In_2410,In_2238);
nand U3691 (N_3691,In_2483,In_1791);
or U3692 (N_3692,In_1080,In_1850);
nand U3693 (N_3693,In_1372,In_694);
or U3694 (N_3694,In_2227,In_2222);
nand U3695 (N_3695,In_1240,In_1070);
and U3696 (N_3696,In_1723,In_1412);
and U3697 (N_3697,In_1667,In_922);
nand U3698 (N_3698,In_2542,In_161);
and U3699 (N_3699,In_2397,In_1378);
and U3700 (N_3700,In_2878,In_1014);
and U3701 (N_3701,In_1802,In_1352);
nand U3702 (N_3702,In_2233,In_518);
nor U3703 (N_3703,In_180,In_1598);
nand U3704 (N_3704,In_1790,In_285);
nand U3705 (N_3705,In_897,In_277);
nor U3706 (N_3706,In_531,In_2253);
nand U3707 (N_3707,In_956,In_1516);
and U3708 (N_3708,In_741,In_1555);
or U3709 (N_3709,In_2150,In_1714);
or U3710 (N_3710,In_2820,In_1394);
nand U3711 (N_3711,In_1959,In_2419);
nand U3712 (N_3712,In_1585,In_2176);
or U3713 (N_3713,In_2024,In_208);
xor U3714 (N_3714,In_1550,In_1928);
nand U3715 (N_3715,In_1947,In_2920);
or U3716 (N_3716,In_2145,In_1073);
or U3717 (N_3717,In_2813,In_402);
nand U3718 (N_3718,In_585,In_1262);
nand U3719 (N_3719,In_1381,In_115);
nand U3720 (N_3720,In_31,In_815);
nand U3721 (N_3721,In_1753,In_2863);
nor U3722 (N_3722,In_289,In_550);
and U3723 (N_3723,In_2487,In_2328);
and U3724 (N_3724,In_1661,In_2108);
and U3725 (N_3725,In_1901,In_2504);
or U3726 (N_3726,In_2779,In_253);
nand U3727 (N_3727,In_1085,In_1963);
nor U3728 (N_3728,In_556,In_2758);
or U3729 (N_3729,In_1584,In_92);
nand U3730 (N_3730,In_435,In_2667);
nand U3731 (N_3731,In_2497,In_2410);
and U3732 (N_3732,In_1998,In_1723);
nand U3733 (N_3733,In_1991,In_335);
and U3734 (N_3734,In_990,In_934);
nor U3735 (N_3735,In_2669,In_667);
nand U3736 (N_3736,In_567,In_1386);
or U3737 (N_3737,In_610,In_748);
nand U3738 (N_3738,In_547,In_2949);
or U3739 (N_3739,In_1784,In_2483);
nand U3740 (N_3740,In_2526,In_1324);
or U3741 (N_3741,In_2278,In_1761);
nor U3742 (N_3742,In_2962,In_2577);
and U3743 (N_3743,In_2290,In_1735);
nor U3744 (N_3744,In_1964,In_121);
and U3745 (N_3745,In_888,In_2309);
or U3746 (N_3746,In_1516,In_2092);
nand U3747 (N_3747,In_185,In_2558);
and U3748 (N_3748,In_1314,In_1600);
or U3749 (N_3749,In_937,In_2734);
nand U3750 (N_3750,In_1460,In_1983);
and U3751 (N_3751,In_746,In_2009);
or U3752 (N_3752,In_79,In_727);
nor U3753 (N_3753,In_679,In_708);
and U3754 (N_3754,In_845,In_2330);
nand U3755 (N_3755,In_516,In_887);
nand U3756 (N_3756,In_1190,In_212);
nor U3757 (N_3757,In_1417,In_380);
or U3758 (N_3758,In_1952,In_407);
nand U3759 (N_3759,In_2078,In_2408);
nor U3760 (N_3760,In_2233,In_568);
or U3761 (N_3761,In_215,In_2576);
nor U3762 (N_3762,In_14,In_76);
nand U3763 (N_3763,In_432,In_448);
nor U3764 (N_3764,In_450,In_1025);
nand U3765 (N_3765,In_2426,In_700);
nor U3766 (N_3766,In_495,In_2696);
or U3767 (N_3767,In_315,In_2411);
nor U3768 (N_3768,In_349,In_1129);
nor U3769 (N_3769,In_2162,In_1376);
or U3770 (N_3770,In_1918,In_1805);
xnor U3771 (N_3771,In_897,In_1569);
nor U3772 (N_3772,In_2232,In_337);
nand U3773 (N_3773,In_607,In_341);
or U3774 (N_3774,In_137,In_2947);
and U3775 (N_3775,In_442,In_1591);
and U3776 (N_3776,In_1644,In_336);
and U3777 (N_3777,In_2222,In_867);
nor U3778 (N_3778,In_1138,In_710);
and U3779 (N_3779,In_1453,In_2238);
and U3780 (N_3780,In_2957,In_1142);
nand U3781 (N_3781,In_861,In_1709);
or U3782 (N_3782,In_1132,In_283);
and U3783 (N_3783,In_1641,In_1666);
or U3784 (N_3784,In_242,In_635);
or U3785 (N_3785,In_1516,In_469);
or U3786 (N_3786,In_2498,In_706);
and U3787 (N_3787,In_2688,In_496);
or U3788 (N_3788,In_2852,In_1615);
and U3789 (N_3789,In_1227,In_2674);
and U3790 (N_3790,In_1845,In_1135);
nand U3791 (N_3791,In_2725,In_606);
nand U3792 (N_3792,In_1628,In_1144);
nand U3793 (N_3793,In_802,In_2280);
nand U3794 (N_3794,In_1974,In_2217);
and U3795 (N_3795,In_738,In_2429);
and U3796 (N_3796,In_2570,In_1083);
and U3797 (N_3797,In_1900,In_127);
nor U3798 (N_3798,In_1289,In_1827);
nand U3799 (N_3799,In_519,In_141);
and U3800 (N_3800,In_1711,In_965);
nor U3801 (N_3801,In_2305,In_2746);
nand U3802 (N_3802,In_691,In_1407);
nand U3803 (N_3803,In_727,In_196);
or U3804 (N_3804,In_1859,In_1386);
and U3805 (N_3805,In_1302,In_612);
nand U3806 (N_3806,In_2850,In_19);
nor U3807 (N_3807,In_625,In_2538);
and U3808 (N_3808,In_2515,In_1770);
and U3809 (N_3809,In_1404,In_1677);
nand U3810 (N_3810,In_2262,In_707);
and U3811 (N_3811,In_2631,In_177);
nor U3812 (N_3812,In_2579,In_1099);
and U3813 (N_3813,In_2112,In_2784);
nand U3814 (N_3814,In_1525,In_2506);
nor U3815 (N_3815,In_2196,In_2207);
or U3816 (N_3816,In_2061,In_148);
and U3817 (N_3817,In_2529,In_839);
or U3818 (N_3818,In_385,In_2337);
and U3819 (N_3819,In_561,In_1791);
nor U3820 (N_3820,In_1146,In_409);
or U3821 (N_3821,In_1620,In_2913);
nor U3822 (N_3822,In_806,In_1933);
or U3823 (N_3823,In_292,In_2634);
nor U3824 (N_3824,In_2897,In_1717);
nand U3825 (N_3825,In_1381,In_1078);
or U3826 (N_3826,In_2787,In_897);
or U3827 (N_3827,In_365,In_1588);
and U3828 (N_3828,In_2213,In_1584);
and U3829 (N_3829,In_2645,In_1147);
nand U3830 (N_3830,In_1797,In_407);
and U3831 (N_3831,In_1951,In_2378);
or U3832 (N_3832,In_231,In_2406);
nand U3833 (N_3833,In_1757,In_1503);
or U3834 (N_3834,In_2309,In_902);
nor U3835 (N_3835,In_108,In_2184);
and U3836 (N_3836,In_480,In_671);
nor U3837 (N_3837,In_1393,In_2587);
or U3838 (N_3838,In_1005,In_1807);
nand U3839 (N_3839,In_2563,In_1776);
nor U3840 (N_3840,In_1534,In_2924);
nand U3841 (N_3841,In_2338,In_544);
or U3842 (N_3842,In_649,In_688);
or U3843 (N_3843,In_2963,In_1742);
and U3844 (N_3844,In_2512,In_2756);
nor U3845 (N_3845,In_1138,In_930);
or U3846 (N_3846,In_2883,In_2189);
nor U3847 (N_3847,In_1449,In_1233);
nor U3848 (N_3848,In_1373,In_1141);
nor U3849 (N_3849,In_2832,In_241);
nor U3850 (N_3850,In_2190,In_14);
nand U3851 (N_3851,In_757,In_869);
nor U3852 (N_3852,In_2806,In_1894);
nand U3853 (N_3853,In_913,In_739);
and U3854 (N_3854,In_2501,In_334);
nor U3855 (N_3855,In_621,In_1230);
and U3856 (N_3856,In_1625,In_423);
xnor U3857 (N_3857,In_2538,In_1443);
and U3858 (N_3858,In_1017,In_2195);
nand U3859 (N_3859,In_951,In_240);
and U3860 (N_3860,In_808,In_1205);
nor U3861 (N_3861,In_1875,In_1538);
nand U3862 (N_3862,In_744,In_1744);
and U3863 (N_3863,In_2833,In_2327);
or U3864 (N_3864,In_2223,In_1415);
nand U3865 (N_3865,In_392,In_2597);
nor U3866 (N_3866,In_469,In_1216);
and U3867 (N_3867,In_108,In_1229);
nor U3868 (N_3868,In_721,In_956);
or U3869 (N_3869,In_997,In_2870);
nor U3870 (N_3870,In_184,In_1697);
nor U3871 (N_3871,In_777,In_573);
and U3872 (N_3872,In_1509,In_1748);
and U3873 (N_3873,In_1845,In_2148);
or U3874 (N_3874,In_2009,In_2111);
or U3875 (N_3875,In_998,In_9);
nand U3876 (N_3876,In_2562,In_1315);
or U3877 (N_3877,In_2788,In_2599);
xnor U3878 (N_3878,In_298,In_2342);
or U3879 (N_3879,In_1915,In_1859);
nor U3880 (N_3880,In_2119,In_338);
and U3881 (N_3881,In_2667,In_946);
or U3882 (N_3882,In_1730,In_2963);
and U3883 (N_3883,In_2243,In_1226);
nor U3884 (N_3884,In_424,In_1180);
and U3885 (N_3885,In_1963,In_2885);
or U3886 (N_3886,In_1113,In_1972);
nor U3887 (N_3887,In_1181,In_1257);
and U3888 (N_3888,In_1065,In_1837);
nand U3889 (N_3889,In_2932,In_1985);
and U3890 (N_3890,In_2154,In_2065);
nor U3891 (N_3891,In_1983,In_405);
or U3892 (N_3892,In_2318,In_2741);
nand U3893 (N_3893,In_234,In_2301);
and U3894 (N_3894,In_2354,In_883);
and U3895 (N_3895,In_878,In_50);
or U3896 (N_3896,In_940,In_266);
or U3897 (N_3897,In_821,In_1056);
or U3898 (N_3898,In_1700,In_1991);
nand U3899 (N_3899,In_2006,In_876);
nand U3900 (N_3900,In_1574,In_2361);
or U3901 (N_3901,In_2317,In_1037);
or U3902 (N_3902,In_253,In_2440);
or U3903 (N_3903,In_1417,In_1858);
and U3904 (N_3904,In_1098,In_1429);
and U3905 (N_3905,In_187,In_975);
nand U3906 (N_3906,In_2563,In_2559);
or U3907 (N_3907,In_1248,In_1513);
nand U3908 (N_3908,In_406,In_806);
nor U3909 (N_3909,In_1025,In_1057);
nor U3910 (N_3910,In_1768,In_2321);
nand U3911 (N_3911,In_2312,In_1166);
xor U3912 (N_3912,In_2159,In_2921);
and U3913 (N_3913,In_222,In_1326);
or U3914 (N_3914,In_2197,In_1853);
or U3915 (N_3915,In_2259,In_2090);
nor U3916 (N_3916,In_1786,In_1249);
nor U3917 (N_3917,In_447,In_2528);
or U3918 (N_3918,In_2316,In_553);
or U3919 (N_3919,In_1889,In_505);
nor U3920 (N_3920,In_680,In_1054);
nand U3921 (N_3921,In_2331,In_626);
nand U3922 (N_3922,In_1847,In_288);
nand U3923 (N_3923,In_2794,In_243);
and U3924 (N_3924,In_481,In_2682);
or U3925 (N_3925,In_1692,In_719);
xor U3926 (N_3926,In_415,In_481);
or U3927 (N_3927,In_591,In_1315);
and U3928 (N_3928,In_686,In_1357);
nor U3929 (N_3929,In_2883,In_264);
and U3930 (N_3930,In_1219,In_766);
nand U3931 (N_3931,In_1553,In_1825);
or U3932 (N_3932,In_2002,In_1604);
or U3933 (N_3933,In_2532,In_1695);
and U3934 (N_3934,In_1550,In_782);
nor U3935 (N_3935,In_774,In_443);
and U3936 (N_3936,In_1524,In_1987);
xor U3937 (N_3937,In_2871,In_2064);
nor U3938 (N_3938,In_1797,In_2731);
and U3939 (N_3939,In_2520,In_1767);
and U3940 (N_3940,In_1246,In_632);
or U3941 (N_3941,In_1626,In_1158);
or U3942 (N_3942,In_1847,In_11);
nor U3943 (N_3943,In_2108,In_2985);
nor U3944 (N_3944,In_442,In_594);
or U3945 (N_3945,In_191,In_2550);
and U3946 (N_3946,In_2251,In_2928);
and U3947 (N_3947,In_1128,In_2326);
nor U3948 (N_3948,In_652,In_2806);
nand U3949 (N_3949,In_66,In_528);
nand U3950 (N_3950,In_753,In_2894);
nor U3951 (N_3951,In_176,In_196);
nor U3952 (N_3952,In_1719,In_1226);
nor U3953 (N_3953,In_320,In_2146);
and U3954 (N_3954,In_2779,In_2128);
or U3955 (N_3955,In_695,In_1160);
and U3956 (N_3956,In_835,In_2166);
nor U3957 (N_3957,In_2373,In_901);
nand U3958 (N_3958,In_1676,In_2737);
nand U3959 (N_3959,In_2061,In_2334);
nand U3960 (N_3960,In_1768,In_2460);
nor U3961 (N_3961,In_1721,In_948);
and U3962 (N_3962,In_2245,In_2881);
nor U3963 (N_3963,In_1986,In_90);
nor U3964 (N_3964,In_1185,In_961);
nor U3965 (N_3965,In_543,In_1911);
or U3966 (N_3966,In_516,In_2357);
and U3967 (N_3967,In_2390,In_342);
or U3968 (N_3968,In_1373,In_883);
or U3969 (N_3969,In_925,In_2239);
or U3970 (N_3970,In_1775,In_1521);
nand U3971 (N_3971,In_258,In_981);
nand U3972 (N_3972,In_2110,In_2386);
and U3973 (N_3973,In_1522,In_22);
nor U3974 (N_3974,In_1833,In_1684);
or U3975 (N_3975,In_2575,In_1439);
and U3976 (N_3976,In_1147,In_2598);
nor U3977 (N_3977,In_1796,In_2383);
and U3978 (N_3978,In_2120,In_44);
nand U3979 (N_3979,In_1114,In_2346);
or U3980 (N_3980,In_2603,In_2564);
or U3981 (N_3981,In_1154,In_2967);
and U3982 (N_3982,In_929,In_327);
and U3983 (N_3983,In_1121,In_958);
and U3984 (N_3984,In_2312,In_2125);
nand U3985 (N_3985,In_612,In_1704);
nor U3986 (N_3986,In_1582,In_2096);
or U3987 (N_3987,In_2613,In_2309);
nor U3988 (N_3988,In_1437,In_521);
nor U3989 (N_3989,In_50,In_1646);
nand U3990 (N_3990,In_2341,In_674);
xnor U3991 (N_3991,In_1373,In_666);
and U3992 (N_3992,In_471,In_2396);
or U3993 (N_3993,In_1881,In_426);
and U3994 (N_3994,In_689,In_1612);
and U3995 (N_3995,In_813,In_62);
nor U3996 (N_3996,In_1418,In_1664);
nand U3997 (N_3997,In_598,In_308);
or U3998 (N_3998,In_2889,In_739);
nand U3999 (N_3999,In_2104,In_1517);
or U4000 (N_4000,In_1344,In_1801);
nor U4001 (N_4001,In_1441,In_2668);
and U4002 (N_4002,In_294,In_563);
or U4003 (N_4003,In_835,In_2106);
or U4004 (N_4004,In_920,In_2007);
nor U4005 (N_4005,In_1020,In_2063);
or U4006 (N_4006,In_219,In_2227);
and U4007 (N_4007,In_1887,In_2408);
or U4008 (N_4008,In_2783,In_1678);
nor U4009 (N_4009,In_2265,In_2555);
nand U4010 (N_4010,In_1688,In_465);
or U4011 (N_4011,In_1329,In_612);
and U4012 (N_4012,In_1058,In_1001);
nor U4013 (N_4013,In_2776,In_719);
nand U4014 (N_4014,In_924,In_124);
nand U4015 (N_4015,In_2566,In_2913);
nand U4016 (N_4016,In_2285,In_462);
or U4017 (N_4017,In_2776,In_367);
and U4018 (N_4018,In_474,In_991);
nor U4019 (N_4019,In_398,In_2493);
nor U4020 (N_4020,In_512,In_345);
nand U4021 (N_4021,In_1946,In_1388);
nor U4022 (N_4022,In_566,In_92);
nor U4023 (N_4023,In_1654,In_2142);
and U4024 (N_4024,In_1690,In_2605);
nand U4025 (N_4025,In_2556,In_1732);
nand U4026 (N_4026,In_1108,In_1266);
or U4027 (N_4027,In_2369,In_2211);
nand U4028 (N_4028,In_2912,In_769);
nor U4029 (N_4029,In_1086,In_624);
nor U4030 (N_4030,In_2645,In_2131);
xor U4031 (N_4031,In_2318,In_2443);
nor U4032 (N_4032,In_86,In_1787);
nand U4033 (N_4033,In_2714,In_2287);
or U4034 (N_4034,In_2634,In_2843);
and U4035 (N_4035,In_2368,In_354);
nor U4036 (N_4036,In_2466,In_964);
or U4037 (N_4037,In_1807,In_678);
and U4038 (N_4038,In_2080,In_1356);
nor U4039 (N_4039,In_1266,In_1406);
and U4040 (N_4040,In_2419,In_1755);
or U4041 (N_4041,In_1590,In_2816);
and U4042 (N_4042,In_2004,In_1933);
nor U4043 (N_4043,In_2097,In_1494);
and U4044 (N_4044,In_960,In_1067);
or U4045 (N_4045,In_1109,In_216);
nor U4046 (N_4046,In_2056,In_1384);
nand U4047 (N_4047,In_1897,In_1095);
nand U4048 (N_4048,In_1343,In_1282);
or U4049 (N_4049,In_2651,In_561);
nor U4050 (N_4050,In_194,In_1218);
xor U4051 (N_4051,In_2437,In_527);
nor U4052 (N_4052,In_2024,In_1834);
nand U4053 (N_4053,In_2507,In_1011);
nor U4054 (N_4054,In_1050,In_17);
or U4055 (N_4055,In_1829,In_422);
or U4056 (N_4056,In_147,In_787);
nand U4057 (N_4057,In_1958,In_626);
nor U4058 (N_4058,In_1855,In_2883);
and U4059 (N_4059,In_399,In_1270);
nand U4060 (N_4060,In_836,In_2851);
nand U4061 (N_4061,In_181,In_2757);
or U4062 (N_4062,In_1614,In_2382);
or U4063 (N_4063,In_2041,In_1304);
nor U4064 (N_4064,In_1075,In_444);
or U4065 (N_4065,In_770,In_2194);
or U4066 (N_4066,In_526,In_337);
or U4067 (N_4067,In_561,In_2848);
or U4068 (N_4068,In_21,In_972);
and U4069 (N_4069,In_588,In_435);
or U4070 (N_4070,In_858,In_222);
and U4071 (N_4071,In_1260,In_1453);
xor U4072 (N_4072,In_2323,In_111);
nor U4073 (N_4073,In_115,In_1614);
or U4074 (N_4074,In_2891,In_1528);
and U4075 (N_4075,In_1086,In_445);
and U4076 (N_4076,In_1232,In_1710);
or U4077 (N_4077,In_2531,In_661);
and U4078 (N_4078,In_209,In_728);
or U4079 (N_4079,In_1204,In_2925);
nand U4080 (N_4080,In_1125,In_2869);
nand U4081 (N_4081,In_703,In_1927);
or U4082 (N_4082,In_2772,In_2177);
or U4083 (N_4083,In_2671,In_213);
nor U4084 (N_4084,In_2987,In_1726);
nor U4085 (N_4085,In_2645,In_2343);
nand U4086 (N_4086,In_721,In_775);
nor U4087 (N_4087,In_2915,In_1523);
and U4088 (N_4088,In_2733,In_2521);
nor U4089 (N_4089,In_2386,In_2206);
or U4090 (N_4090,In_282,In_2690);
or U4091 (N_4091,In_1277,In_1856);
nor U4092 (N_4092,In_645,In_2643);
nand U4093 (N_4093,In_242,In_2735);
and U4094 (N_4094,In_2445,In_1679);
and U4095 (N_4095,In_1961,In_1788);
or U4096 (N_4096,In_5,In_379);
nor U4097 (N_4097,In_2279,In_1655);
nor U4098 (N_4098,In_2597,In_1812);
or U4099 (N_4099,In_1473,In_1258);
nor U4100 (N_4100,In_1375,In_2755);
or U4101 (N_4101,In_2675,In_413);
or U4102 (N_4102,In_370,In_1505);
nor U4103 (N_4103,In_1924,In_555);
and U4104 (N_4104,In_1063,In_213);
nand U4105 (N_4105,In_2349,In_2906);
nor U4106 (N_4106,In_203,In_2302);
nor U4107 (N_4107,In_1442,In_805);
nor U4108 (N_4108,In_1927,In_688);
nand U4109 (N_4109,In_679,In_1857);
nor U4110 (N_4110,In_1158,In_80);
nand U4111 (N_4111,In_1278,In_779);
nor U4112 (N_4112,In_1894,In_2271);
and U4113 (N_4113,In_1710,In_1977);
nand U4114 (N_4114,In_2064,In_2751);
or U4115 (N_4115,In_2480,In_2658);
or U4116 (N_4116,In_2929,In_2625);
or U4117 (N_4117,In_1926,In_2186);
or U4118 (N_4118,In_2403,In_2834);
and U4119 (N_4119,In_2080,In_1260);
and U4120 (N_4120,In_1682,In_2838);
nor U4121 (N_4121,In_558,In_341);
nor U4122 (N_4122,In_2616,In_1087);
or U4123 (N_4123,In_2248,In_2051);
or U4124 (N_4124,In_2039,In_570);
or U4125 (N_4125,In_2802,In_1207);
nor U4126 (N_4126,In_463,In_2623);
and U4127 (N_4127,In_2701,In_1054);
nand U4128 (N_4128,In_638,In_1462);
or U4129 (N_4129,In_1878,In_1422);
or U4130 (N_4130,In_1258,In_308);
or U4131 (N_4131,In_2887,In_131);
or U4132 (N_4132,In_2284,In_506);
nor U4133 (N_4133,In_592,In_684);
nand U4134 (N_4134,In_2622,In_1333);
and U4135 (N_4135,In_1868,In_1197);
nand U4136 (N_4136,In_838,In_2692);
xor U4137 (N_4137,In_2814,In_1159);
nor U4138 (N_4138,In_2461,In_2336);
or U4139 (N_4139,In_1830,In_2576);
nor U4140 (N_4140,In_1445,In_2931);
nand U4141 (N_4141,In_920,In_2563);
or U4142 (N_4142,In_2952,In_1144);
nor U4143 (N_4143,In_1637,In_1052);
nor U4144 (N_4144,In_600,In_36);
nor U4145 (N_4145,In_2628,In_1859);
and U4146 (N_4146,In_2571,In_1159);
or U4147 (N_4147,In_390,In_2863);
and U4148 (N_4148,In_239,In_1749);
nor U4149 (N_4149,In_318,In_2485);
nor U4150 (N_4150,In_1425,In_1059);
xor U4151 (N_4151,In_1040,In_2103);
or U4152 (N_4152,In_15,In_31);
or U4153 (N_4153,In_2012,In_1742);
nand U4154 (N_4154,In_1638,In_2188);
and U4155 (N_4155,In_2585,In_1113);
and U4156 (N_4156,In_1089,In_1194);
and U4157 (N_4157,In_740,In_1231);
nor U4158 (N_4158,In_887,In_2337);
or U4159 (N_4159,In_396,In_1706);
xnor U4160 (N_4160,In_2918,In_2401);
nand U4161 (N_4161,In_2515,In_1796);
nor U4162 (N_4162,In_916,In_2576);
or U4163 (N_4163,In_2203,In_532);
and U4164 (N_4164,In_1542,In_2595);
nor U4165 (N_4165,In_598,In_607);
or U4166 (N_4166,In_2891,In_885);
nor U4167 (N_4167,In_1836,In_868);
nor U4168 (N_4168,In_919,In_1406);
nand U4169 (N_4169,In_2444,In_896);
nand U4170 (N_4170,In_2838,In_1640);
or U4171 (N_4171,In_2251,In_775);
and U4172 (N_4172,In_1805,In_1128);
and U4173 (N_4173,In_2322,In_526);
nor U4174 (N_4174,In_2871,In_2207);
or U4175 (N_4175,In_2333,In_1494);
and U4176 (N_4176,In_2154,In_996);
nor U4177 (N_4177,In_2394,In_373);
nor U4178 (N_4178,In_1485,In_309);
and U4179 (N_4179,In_309,In_856);
or U4180 (N_4180,In_1989,In_1624);
and U4181 (N_4181,In_2729,In_2263);
nand U4182 (N_4182,In_1830,In_1617);
nand U4183 (N_4183,In_1589,In_2676);
nor U4184 (N_4184,In_2243,In_128);
nor U4185 (N_4185,In_1488,In_2762);
nand U4186 (N_4186,In_100,In_607);
nand U4187 (N_4187,In_2568,In_2448);
and U4188 (N_4188,In_2125,In_1513);
xnor U4189 (N_4189,In_947,In_363);
or U4190 (N_4190,In_1146,In_2611);
or U4191 (N_4191,In_2150,In_1141);
nand U4192 (N_4192,In_2633,In_2212);
and U4193 (N_4193,In_1640,In_1910);
nor U4194 (N_4194,In_2743,In_1057);
nor U4195 (N_4195,In_1154,In_1806);
nand U4196 (N_4196,In_1939,In_564);
or U4197 (N_4197,In_888,In_1264);
or U4198 (N_4198,In_2841,In_2109);
and U4199 (N_4199,In_2570,In_1487);
nor U4200 (N_4200,In_1934,In_1632);
or U4201 (N_4201,In_2929,In_1554);
nand U4202 (N_4202,In_2793,In_1916);
nor U4203 (N_4203,In_784,In_2672);
nor U4204 (N_4204,In_2974,In_2493);
nor U4205 (N_4205,In_441,In_144);
nand U4206 (N_4206,In_2188,In_1153);
and U4207 (N_4207,In_2436,In_787);
or U4208 (N_4208,In_1153,In_81);
nand U4209 (N_4209,In_192,In_2664);
nand U4210 (N_4210,In_1280,In_1178);
nand U4211 (N_4211,In_1300,In_891);
and U4212 (N_4212,In_819,In_1659);
or U4213 (N_4213,In_1276,In_74);
nor U4214 (N_4214,In_2235,In_1627);
or U4215 (N_4215,In_2480,In_1793);
nand U4216 (N_4216,In_1198,In_40);
nand U4217 (N_4217,In_1196,In_514);
and U4218 (N_4218,In_776,In_1742);
nand U4219 (N_4219,In_2175,In_2481);
and U4220 (N_4220,In_1447,In_1899);
or U4221 (N_4221,In_652,In_723);
nand U4222 (N_4222,In_1537,In_2279);
or U4223 (N_4223,In_1131,In_195);
and U4224 (N_4224,In_2626,In_2578);
and U4225 (N_4225,In_2217,In_1573);
nor U4226 (N_4226,In_2787,In_1945);
nand U4227 (N_4227,In_2231,In_1810);
nand U4228 (N_4228,In_848,In_913);
nand U4229 (N_4229,In_1220,In_1242);
nor U4230 (N_4230,In_2293,In_1795);
nor U4231 (N_4231,In_2373,In_2708);
nor U4232 (N_4232,In_765,In_981);
nand U4233 (N_4233,In_2031,In_1905);
and U4234 (N_4234,In_915,In_1315);
and U4235 (N_4235,In_1810,In_2406);
and U4236 (N_4236,In_1581,In_1746);
and U4237 (N_4237,In_1424,In_1118);
and U4238 (N_4238,In_2204,In_2220);
nand U4239 (N_4239,In_1037,In_2406);
and U4240 (N_4240,In_2944,In_2054);
nor U4241 (N_4241,In_138,In_1115);
or U4242 (N_4242,In_1828,In_1833);
and U4243 (N_4243,In_473,In_2188);
nor U4244 (N_4244,In_2562,In_1281);
and U4245 (N_4245,In_779,In_961);
nand U4246 (N_4246,In_643,In_2889);
nand U4247 (N_4247,In_2661,In_2033);
and U4248 (N_4248,In_1185,In_523);
and U4249 (N_4249,In_1572,In_2060);
nand U4250 (N_4250,In_1584,In_1948);
or U4251 (N_4251,In_1842,In_91);
xor U4252 (N_4252,In_165,In_2747);
and U4253 (N_4253,In_248,In_597);
or U4254 (N_4254,In_673,In_939);
nor U4255 (N_4255,In_1690,In_849);
nand U4256 (N_4256,In_2216,In_469);
and U4257 (N_4257,In_2204,In_687);
or U4258 (N_4258,In_2111,In_25);
nor U4259 (N_4259,In_2912,In_889);
and U4260 (N_4260,In_2591,In_2489);
or U4261 (N_4261,In_1438,In_1588);
or U4262 (N_4262,In_1542,In_224);
nor U4263 (N_4263,In_2237,In_2549);
nor U4264 (N_4264,In_931,In_530);
or U4265 (N_4265,In_2682,In_1875);
or U4266 (N_4266,In_2266,In_2571);
nand U4267 (N_4267,In_2560,In_1741);
and U4268 (N_4268,In_1541,In_659);
nand U4269 (N_4269,In_274,In_1967);
or U4270 (N_4270,In_2067,In_1496);
nor U4271 (N_4271,In_1592,In_1181);
nor U4272 (N_4272,In_709,In_2941);
nand U4273 (N_4273,In_40,In_1392);
or U4274 (N_4274,In_1358,In_254);
or U4275 (N_4275,In_2963,In_2918);
or U4276 (N_4276,In_1138,In_673);
nor U4277 (N_4277,In_1265,In_2952);
or U4278 (N_4278,In_243,In_2756);
or U4279 (N_4279,In_2020,In_57);
and U4280 (N_4280,In_2965,In_2227);
and U4281 (N_4281,In_1966,In_1815);
or U4282 (N_4282,In_2816,In_545);
nor U4283 (N_4283,In_2696,In_623);
nand U4284 (N_4284,In_1235,In_1906);
and U4285 (N_4285,In_1784,In_510);
and U4286 (N_4286,In_1424,In_1205);
nor U4287 (N_4287,In_89,In_1538);
and U4288 (N_4288,In_902,In_819);
nor U4289 (N_4289,In_1465,In_2742);
nand U4290 (N_4290,In_1851,In_164);
and U4291 (N_4291,In_1024,In_1470);
nor U4292 (N_4292,In_1340,In_900);
or U4293 (N_4293,In_1522,In_245);
nor U4294 (N_4294,In_333,In_2941);
nor U4295 (N_4295,In_710,In_2159);
nand U4296 (N_4296,In_1734,In_520);
nand U4297 (N_4297,In_572,In_2924);
nand U4298 (N_4298,In_1994,In_852);
nand U4299 (N_4299,In_440,In_1542);
and U4300 (N_4300,In_1853,In_1742);
nor U4301 (N_4301,In_978,In_2162);
nor U4302 (N_4302,In_2774,In_1886);
or U4303 (N_4303,In_268,In_574);
and U4304 (N_4304,In_1761,In_1949);
and U4305 (N_4305,In_610,In_1484);
or U4306 (N_4306,In_1956,In_1473);
or U4307 (N_4307,In_2102,In_1213);
and U4308 (N_4308,In_163,In_2680);
nor U4309 (N_4309,In_2784,In_1830);
or U4310 (N_4310,In_913,In_1810);
nand U4311 (N_4311,In_2748,In_2415);
and U4312 (N_4312,In_1309,In_77);
nor U4313 (N_4313,In_910,In_950);
and U4314 (N_4314,In_1477,In_2019);
and U4315 (N_4315,In_2740,In_136);
and U4316 (N_4316,In_431,In_1109);
or U4317 (N_4317,In_2784,In_2303);
nor U4318 (N_4318,In_2922,In_1365);
or U4319 (N_4319,In_2054,In_1696);
nor U4320 (N_4320,In_580,In_1366);
or U4321 (N_4321,In_2777,In_2015);
or U4322 (N_4322,In_547,In_2110);
nand U4323 (N_4323,In_1820,In_1809);
nor U4324 (N_4324,In_2740,In_2383);
and U4325 (N_4325,In_2682,In_275);
and U4326 (N_4326,In_646,In_1117);
nor U4327 (N_4327,In_1993,In_2027);
or U4328 (N_4328,In_2329,In_2644);
nor U4329 (N_4329,In_654,In_2401);
or U4330 (N_4330,In_2109,In_1804);
nor U4331 (N_4331,In_592,In_1432);
nor U4332 (N_4332,In_2093,In_1423);
or U4333 (N_4333,In_871,In_916);
and U4334 (N_4334,In_2548,In_2786);
or U4335 (N_4335,In_1231,In_1518);
or U4336 (N_4336,In_475,In_2526);
nand U4337 (N_4337,In_2923,In_1055);
or U4338 (N_4338,In_2602,In_2908);
nor U4339 (N_4339,In_2195,In_2776);
nor U4340 (N_4340,In_114,In_1883);
nor U4341 (N_4341,In_1576,In_2684);
and U4342 (N_4342,In_1032,In_1918);
nand U4343 (N_4343,In_2949,In_695);
and U4344 (N_4344,In_1055,In_2538);
or U4345 (N_4345,In_1795,In_116);
or U4346 (N_4346,In_1965,In_2681);
nor U4347 (N_4347,In_1359,In_2618);
and U4348 (N_4348,In_2900,In_409);
nand U4349 (N_4349,In_2294,In_1089);
and U4350 (N_4350,In_2546,In_2977);
and U4351 (N_4351,In_1339,In_2617);
nand U4352 (N_4352,In_1926,In_800);
or U4353 (N_4353,In_82,In_2106);
nand U4354 (N_4354,In_679,In_876);
nor U4355 (N_4355,In_576,In_595);
nand U4356 (N_4356,In_797,In_2448);
nor U4357 (N_4357,In_1411,In_771);
nand U4358 (N_4358,In_374,In_1840);
nand U4359 (N_4359,In_874,In_2902);
nor U4360 (N_4360,In_1619,In_631);
and U4361 (N_4361,In_872,In_1171);
nor U4362 (N_4362,In_1111,In_2774);
xnor U4363 (N_4363,In_1409,In_1917);
nor U4364 (N_4364,In_1622,In_2977);
nor U4365 (N_4365,In_1602,In_2099);
or U4366 (N_4366,In_463,In_2985);
nand U4367 (N_4367,In_223,In_2441);
nand U4368 (N_4368,In_2010,In_2209);
and U4369 (N_4369,In_1925,In_936);
nor U4370 (N_4370,In_957,In_2467);
nand U4371 (N_4371,In_1027,In_153);
nand U4372 (N_4372,In_2896,In_294);
and U4373 (N_4373,In_361,In_485);
and U4374 (N_4374,In_2028,In_260);
nor U4375 (N_4375,In_1423,In_2154);
or U4376 (N_4376,In_477,In_2704);
or U4377 (N_4377,In_2012,In_1644);
or U4378 (N_4378,In_594,In_2370);
and U4379 (N_4379,In_136,In_699);
nor U4380 (N_4380,In_1607,In_1036);
and U4381 (N_4381,In_1513,In_1470);
nand U4382 (N_4382,In_2369,In_119);
nor U4383 (N_4383,In_347,In_437);
nand U4384 (N_4384,In_134,In_1487);
xor U4385 (N_4385,In_1522,In_560);
nor U4386 (N_4386,In_330,In_1890);
nor U4387 (N_4387,In_708,In_17);
and U4388 (N_4388,In_967,In_2188);
or U4389 (N_4389,In_2214,In_1104);
nand U4390 (N_4390,In_2045,In_2398);
and U4391 (N_4391,In_2160,In_672);
xnor U4392 (N_4392,In_1382,In_2176);
and U4393 (N_4393,In_521,In_2909);
and U4394 (N_4394,In_314,In_2541);
nor U4395 (N_4395,In_94,In_2344);
or U4396 (N_4396,In_549,In_2989);
nand U4397 (N_4397,In_1441,In_2678);
nand U4398 (N_4398,In_1211,In_1888);
nand U4399 (N_4399,In_172,In_2751);
and U4400 (N_4400,In_2319,In_2858);
xor U4401 (N_4401,In_477,In_1083);
nand U4402 (N_4402,In_537,In_59);
and U4403 (N_4403,In_571,In_2479);
and U4404 (N_4404,In_2913,In_773);
nor U4405 (N_4405,In_1221,In_2786);
and U4406 (N_4406,In_1262,In_2700);
nand U4407 (N_4407,In_2916,In_1832);
and U4408 (N_4408,In_1980,In_913);
and U4409 (N_4409,In_761,In_925);
and U4410 (N_4410,In_155,In_1272);
nand U4411 (N_4411,In_2940,In_1417);
nor U4412 (N_4412,In_847,In_2153);
or U4413 (N_4413,In_2334,In_784);
nand U4414 (N_4414,In_1325,In_899);
or U4415 (N_4415,In_1372,In_1829);
nor U4416 (N_4416,In_1254,In_2310);
nand U4417 (N_4417,In_2499,In_244);
and U4418 (N_4418,In_244,In_1837);
nand U4419 (N_4419,In_2653,In_2257);
nand U4420 (N_4420,In_2885,In_1533);
nand U4421 (N_4421,In_1572,In_2550);
or U4422 (N_4422,In_2922,In_965);
or U4423 (N_4423,In_1682,In_262);
nand U4424 (N_4424,In_2581,In_1600);
nand U4425 (N_4425,In_2434,In_2992);
nand U4426 (N_4426,In_211,In_2537);
and U4427 (N_4427,In_2616,In_2330);
nand U4428 (N_4428,In_440,In_1610);
nand U4429 (N_4429,In_452,In_1251);
nor U4430 (N_4430,In_2220,In_212);
nor U4431 (N_4431,In_1536,In_2354);
nor U4432 (N_4432,In_1548,In_591);
nand U4433 (N_4433,In_1072,In_340);
and U4434 (N_4434,In_2584,In_1465);
nand U4435 (N_4435,In_2544,In_2157);
and U4436 (N_4436,In_187,In_2036);
xnor U4437 (N_4437,In_227,In_1104);
nor U4438 (N_4438,In_1502,In_2746);
or U4439 (N_4439,In_2810,In_2256);
nand U4440 (N_4440,In_2942,In_2619);
or U4441 (N_4441,In_1359,In_2954);
and U4442 (N_4442,In_284,In_1240);
nor U4443 (N_4443,In_1282,In_1541);
or U4444 (N_4444,In_2173,In_59);
nand U4445 (N_4445,In_1208,In_2785);
or U4446 (N_4446,In_1472,In_2698);
and U4447 (N_4447,In_2498,In_2545);
nor U4448 (N_4448,In_592,In_2308);
nand U4449 (N_4449,In_2115,In_891);
and U4450 (N_4450,In_502,In_266);
and U4451 (N_4451,In_1063,In_1299);
nor U4452 (N_4452,In_1803,In_1215);
and U4453 (N_4453,In_989,In_109);
nand U4454 (N_4454,In_1721,In_2659);
nand U4455 (N_4455,In_521,In_1812);
and U4456 (N_4456,In_726,In_50);
or U4457 (N_4457,In_2686,In_1265);
or U4458 (N_4458,In_557,In_960);
xor U4459 (N_4459,In_948,In_1612);
and U4460 (N_4460,In_733,In_2422);
nor U4461 (N_4461,In_2256,In_422);
and U4462 (N_4462,In_177,In_2948);
or U4463 (N_4463,In_536,In_860);
or U4464 (N_4464,In_1382,In_196);
and U4465 (N_4465,In_2418,In_287);
or U4466 (N_4466,In_984,In_497);
and U4467 (N_4467,In_198,In_2891);
or U4468 (N_4468,In_1391,In_341);
and U4469 (N_4469,In_1421,In_2304);
nor U4470 (N_4470,In_2393,In_1419);
and U4471 (N_4471,In_839,In_262);
nand U4472 (N_4472,In_1099,In_612);
or U4473 (N_4473,In_1192,In_1002);
nor U4474 (N_4474,In_2636,In_1350);
nand U4475 (N_4475,In_1015,In_977);
nor U4476 (N_4476,In_1626,In_2533);
or U4477 (N_4477,In_1853,In_1348);
or U4478 (N_4478,In_209,In_1572);
or U4479 (N_4479,In_291,In_2273);
nand U4480 (N_4480,In_2003,In_848);
and U4481 (N_4481,In_636,In_148);
and U4482 (N_4482,In_440,In_645);
or U4483 (N_4483,In_1031,In_1212);
nand U4484 (N_4484,In_2869,In_1732);
nor U4485 (N_4485,In_2571,In_1187);
or U4486 (N_4486,In_384,In_2784);
or U4487 (N_4487,In_2695,In_1866);
nor U4488 (N_4488,In_1931,In_1222);
nor U4489 (N_4489,In_411,In_1111);
and U4490 (N_4490,In_1453,In_580);
or U4491 (N_4491,In_255,In_2003);
nor U4492 (N_4492,In_2147,In_797);
and U4493 (N_4493,In_18,In_372);
nor U4494 (N_4494,In_913,In_1875);
or U4495 (N_4495,In_1440,In_2791);
or U4496 (N_4496,In_2130,In_1510);
nand U4497 (N_4497,In_2924,In_1619);
or U4498 (N_4498,In_2629,In_1364);
nor U4499 (N_4499,In_2815,In_2107);
and U4500 (N_4500,In_598,In_2279);
or U4501 (N_4501,In_1407,In_1377);
or U4502 (N_4502,In_2709,In_2555);
and U4503 (N_4503,In_1508,In_1641);
or U4504 (N_4504,In_766,In_1032);
and U4505 (N_4505,In_2936,In_522);
and U4506 (N_4506,In_431,In_1261);
and U4507 (N_4507,In_40,In_762);
or U4508 (N_4508,In_304,In_1806);
nor U4509 (N_4509,In_1765,In_1464);
nand U4510 (N_4510,In_1245,In_2357);
or U4511 (N_4511,In_20,In_2431);
nand U4512 (N_4512,In_825,In_1093);
and U4513 (N_4513,In_2035,In_2805);
or U4514 (N_4514,In_2411,In_996);
nor U4515 (N_4515,In_2413,In_1584);
or U4516 (N_4516,In_2251,In_1713);
and U4517 (N_4517,In_793,In_877);
or U4518 (N_4518,In_675,In_898);
nor U4519 (N_4519,In_2625,In_1614);
or U4520 (N_4520,In_1023,In_2241);
nand U4521 (N_4521,In_2720,In_1651);
nand U4522 (N_4522,In_2658,In_2828);
nand U4523 (N_4523,In_2245,In_1751);
or U4524 (N_4524,In_1067,In_1414);
xnor U4525 (N_4525,In_1301,In_368);
and U4526 (N_4526,In_2645,In_1462);
nor U4527 (N_4527,In_258,In_2793);
and U4528 (N_4528,In_1688,In_1408);
nand U4529 (N_4529,In_2011,In_1726);
nor U4530 (N_4530,In_1470,In_1115);
nand U4531 (N_4531,In_461,In_1464);
and U4532 (N_4532,In_2167,In_2873);
and U4533 (N_4533,In_1782,In_2029);
nand U4534 (N_4534,In_2293,In_2411);
or U4535 (N_4535,In_28,In_1536);
or U4536 (N_4536,In_608,In_341);
nor U4537 (N_4537,In_1801,In_611);
or U4538 (N_4538,In_2520,In_1846);
nand U4539 (N_4539,In_2519,In_682);
and U4540 (N_4540,In_2205,In_737);
xnor U4541 (N_4541,In_2248,In_2618);
nor U4542 (N_4542,In_2115,In_951);
or U4543 (N_4543,In_88,In_2976);
or U4544 (N_4544,In_2195,In_1080);
nor U4545 (N_4545,In_48,In_2856);
nand U4546 (N_4546,In_1110,In_1188);
and U4547 (N_4547,In_1728,In_1476);
nor U4548 (N_4548,In_2468,In_88);
nor U4549 (N_4549,In_2371,In_1891);
or U4550 (N_4550,In_2560,In_1573);
or U4551 (N_4551,In_1205,In_2110);
nand U4552 (N_4552,In_2210,In_376);
nand U4553 (N_4553,In_1706,In_644);
nor U4554 (N_4554,In_1008,In_111);
nand U4555 (N_4555,In_143,In_41);
and U4556 (N_4556,In_236,In_2882);
nor U4557 (N_4557,In_1348,In_151);
and U4558 (N_4558,In_575,In_252);
and U4559 (N_4559,In_1993,In_2535);
nand U4560 (N_4560,In_300,In_1515);
nand U4561 (N_4561,In_1371,In_1237);
or U4562 (N_4562,In_1515,In_2912);
nor U4563 (N_4563,In_174,In_330);
nor U4564 (N_4564,In_55,In_2015);
nand U4565 (N_4565,In_146,In_1127);
nor U4566 (N_4566,In_1406,In_2755);
and U4567 (N_4567,In_1915,In_1260);
xnor U4568 (N_4568,In_2505,In_2545);
and U4569 (N_4569,In_2322,In_826);
nor U4570 (N_4570,In_1758,In_2109);
nand U4571 (N_4571,In_1534,In_1122);
nand U4572 (N_4572,In_2423,In_1859);
xor U4573 (N_4573,In_1619,In_1429);
or U4574 (N_4574,In_1009,In_1843);
and U4575 (N_4575,In_150,In_2848);
or U4576 (N_4576,In_2305,In_1423);
nor U4577 (N_4577,In_2061,In_2982);
nor U4578 (N_4578,In_1100,In_2760);
or U4579 (N_4579,In_1079,In_1320);
nor U4580 (N_4580,In_1343,In_564);
or U4581 (N_4581,In_167,In_1583);
nor U4582 (N_4582,In_1563,In_1689);
nand U4583 (N_4583,In_2868,In_1372);
or U4584 (N_4584,In_2106,In_2864);
or U4585 (N_4585,In_1404,In_1800);
nand U4586 (N_4586,In_2617,In_2756);
nand U4587 (N_4587,In_1679,In_2232);
nand U4588 (N_4588,In_2722,In_1940);
nand U4589 (N_4589,In_1985,In_1280);
and U4590 (N_4590,In_927,In_2954);
nand U4591 (N_4591,In_1187,In_236);
nand U4592 (N_4592,In_2898,In_298);
nand U4593 (N_4593,In_2304,In_1834);
and U4594 (N_4594,In_847,In_2500);
nor U4595 (N_4595,In_401,In_427);
and U4596 (N_4596,In_153,In_1607);
nor U4597 (N_4597,In_2242,In_2743);
or U4598 (N_4598,In_1167,In_1934);
and U4599 (N_4599,In_422,In_2534);
or U4600 (N_4600,In_1474,In_2121);
and U4601 (N_4601,In_1276,In_2329);
and U4602 (N_4602,In_593,In_2060);
nor U4603 (N_4603,In_108,In_2852);
and U4604 (N_4604,In_113,In_2010);
nand U4605 (N_4605,In_505,In_113);
and U4606 (N_4606,In_918,In_2900);
nor U4607 (N_4607,In_1695,In_1162);
or U4608 (N_4608,In_1081,In_1819);
xor U4609 (N_4609,In_2775,In_1994);
xor U4610 (N_4610,In_1675,In_565);
nand U4611 (N_4611,In_1476,In_2632);
nor U4612 (N_4612,In_937,In_1067);
xor U4613 (N_4613,In_1637,In_779);
nor U4614 (N_4614,In_461,In_2061);
nor U4615 (N_4615,In_1313,In_480);
or U4616 (N_4616,In_2927,In_618);
or U4617 (N_4617,In_2148,In_2931);
nor U4618 (N_4618,In_1027,In_924);
nand U4619 (N_4619,In_2809,In_1622);
nand U4620 (N_4620,In_543,In_1579);
nor U4621 (N_4621,In_956,In_2128);
nor U4622 (N_4622,In_198,In_1286);
nand U4623 (N_4623,In_1936,In_2909);
or U4624 (N_4624,In_925,In_1661);
nand U4625 (N_4625,In_454,In_1475);
and U4626 (N_4626,In_2473,In_2237);
nor U4627 (N_4627,In_2415,In_88);
or U4628 (N_4628,In_1618,In_312);
nand U4629 (N_4629,In_2699,In_1423);
or U4630 (N_4630,In_897,In_1957);
and U4631 (N_4631,In_1315,In_1737);
or U4632 (N_4632,In_2380,In_2555);
or U4633 (N_4633,In_964,In_1649);
nand U4634 (N_4634,In_2582,In_2105);
nor U4635 (N_4635,In_812,In_2553);
or U4636 (N_4636,In_1609,In_362);
nand U4637 (N_4637,In_85,In_1677);
nor U4638 (N_4638,In_1330,In_2168);
and U4639 (N_4639,In_1335,In_1045);
and U4640 (N_4640,In_2568,In_2577);
nand U4641 (N_4641,In_1104,In_1126);
and U4642 (N_4642,In_466,In_715);
and U4643 (N_4643,In_888,In_861);
and U4644 (N_4644,In_1849,In_2766);
nor U4645 (N_4645,In_898,In_787);
nor U4646 (N_4646,In_539,In_208);
nor U4647 (N_4647,In_2556,In_2576);
or U4648 (N_4648,In_1839,In_670);
nand U4649 (N_4649,In_2713,In_2646);
and U4650 (N_4650,In_2657,In_432);
and U4651 (N_4651,In_2307,In_2020);
nand U4652 (N_4652,In_1655,In_1058);
or U4653 (N_4653,In_2782,In_1268);
nor U4654 (N_4654,In_2147,In_2531);
and U4655 (N_4655,In_1701,In_2862);
nor U4656 (N_4656,In_2772,In_2410);
and U4657 (N_4657,In_1839,In_1157);
nand U4658 (N_4658,In_2049,In_1428);
and U4659 (N_4659,In_59,In_84);
and U4660 (N_4660,In_510,In_1350);
nor U4661 (N_4661,In_1613,In_1912);
nand U4662 (N_4662,In_2561,In_1567);
and U4663 (N_4663,In_2658,In_2118);
nor U4664 (N_4664,In_1225,In_2546);
or U4665 (N_4665,In_1890,In_696);
nand U4666 (N_4666,In_878,In_1036);
and U4667 (N_4667,In_2258,In_1379);
nor U4668 (N_4668,In_2077,In_1205);
nor U4669 (N_4669,In_1031,In_2608);
and U4670 (N_4670,In_566,In_159);
xor U4671 (N_4671,In_1134,In_1875);
nand U4672 (N_4672,In_2061,In_1727);
or U4673 (N_4673,In_1869,In_856);
and U4674 (N_4674,In_2119,In_2951);
and U4675 (N_4675,In_2149,In_2451);
nor U4676 (N_4676,In_2039,In_191);
nand U4677 (N_4677,In_396,In_1333);
nand U4678 (N_4678,In_1520,In_2912);
and U4679 (N_4679,In_575,In_361);
nand U4680 (N_4680,In_57,In_2977);
nand U4681 (N_4681,In_2711,In_2982);
or U4682 (N_4682,In_512,In_1793);
nor U4683 (N_4683,In_1559,In_2240);
or U4684 (N_4684,In_467,In_1364);
nand U4685 (N_4685,In_243,In_361);
nand U4686 (N_4686,In_1520,In_2530);
and U4687 (N_4687,In_944,In_665);
and U4688 (N_4688,In_2955,In_2223);
and U4689 (N_4689,In_1229,In_2153);
or U4690 (N_4690,In_2781,In_897);
and U4691 (N_4691,In_122,In_501);
nor U4692 (N_4692,In_1954,In_902);
nor U4693 (N_4693,In_1098,In_2911);
or U4694 (N_4694,In_2130,In_1542);
nor U4695 (N_4695,In_1958,In_2652);
nand U4696 (N_4696,In_764,In_398);
nand U4697 (N_4697,In_730,In_2136);
nor U4698 (N_4698,In_2026,In_1474);
or U4699 (N_4699,In_889,In_1954);
and U4700 (N_4700,In_462,In_2342);
nor U4701 (N_4701,In_1063,In_1097);
and U4702 (N_4702,In_2610,In_1367);
nand U4703 (N_4703,In_1729,In_2941);
nand U4704 (N_4704,In_2815,In_1986);
and U4705 (N_4705,In_199,In_1528);
nand U4706 (N_4706,In_456,In_2428);
nor U4707 (N_4707,In_1282,In_628);
nand U4708 (N_4708,In_2981,In_1196);
or U4709 (N_4709,In_2930,In_2761);
or U4710 (N_4710,In_2450,In_901);
or U4711 (N_4711,In_2521,In_382);
or U4712 (N_4712,In_2030,In_2506);
and U4713 (N_4713,In_2401,In_882);
nand U4714 (N_4714,In_263,In_1611);
and U4715 (N_4715,In_2469,In_1154);
nand U4716 (N_4716,In_716,In_2820);
or U4717 (N_4717,In_2890,In_1943);
nor U4718 (N_4718,In_770,In_1722);
nor U4719 (N_4719,In_2821,In_2948);
nor U4720 (N_4720,In_2262,In_677);
and U4721 (N_4721,In_307,In_1675);
or U4722 (N_4722,In_701,In_1088);
nor U4723 (N_4723,In_1342,In_2423);
nor U4724 (N_4724,In_894,In_2868);
and U4725 (N_4725,In_994,In_1537);
and U4726 (N_4726,In_1213,In_1098);
or U4727 (N_4727,In_40,In_1305);
and U4728 (N_4728,In_1953,In_1233);
nand U4729 (N_4729,In_2440,In_32);
and U4730 (N_4730,In_850,In_695);
nand U4731 (N_4731,In_1991,In_1351);
nand U4732 (N_4732,In_2556,In_918);
and U4733 (N_4733,In_451,In_1161);
nand U4734 (N_4734,In_383,In_1313);
or U4735 (N_4735,In_2435,In_571);
and U4736 (N_4736,In_2702,In_890);
nand U4737 (N_4737,In_2764,In_465);
or U4738 (N_4738,In_2009,In_879);
and U4739 (N_4739,In_1039,In_563);
nor U4740 (N_4740,In_2305,In_241);
nand U4741 (N_4741,In_2906,In_1834);
nand U4742 (N_4742,In_2576,In_609);
nand U4743 (N_4743,In_2111,In_501);
nor U4744 (N_4744,In_2584,In_1011);
nor U4745 (N_4745,In_2748,In_386);
and U4746 (N_4746,In_101,In_249);
and U4747 (N_4747,In_1151,In_667);
or U4748 (N_4748,In_2264,In_2844);
nor U4749 (N_4749,In_2166,In_1106);
or U4750 (N_4750,In_2037,In_2004);
nor U4751 (N_4751,In_2641,In_552);
nand U4752 (N_4752,In_963,In_878);
or U4753 (N_4753,In_2086,In_2814);
nand U4754 (N_4754,In_1698,In_261);
and U4755 (N_4755,In_2242,In_843);
and U4756 (N_4756,In_2464,In_1445);
nand U4757 (N_4757,In_1552,In_1693);
nor U4758 (N_4758,In_2491,In_1787);
nor U4759 (N_4759,In_1680,In_673);
nor U4760 (N_4760,In_1404,In_63);
nand U4761 (N_4761,In_600,In_360);
and U4762 (N_4762,In_68,In_2834);
nand U4763 (N_4763,In_1553,In_2324);
nor U4764 (N_4764,In_973,In_2123);
or U4765 (N_4765,In_1209,In_266);
nor U4766 (N_4766,In_2478,In_2052);
or U4767 (N_4767,In_743,In_389);
nor U4768 (N_4768,In_2129,In_1448);
xnor U4769 (N_4769,In_634,In_2942);
or U4770 (N_4770,In_792,In_1230);
nor U4771 (N_4771,In_2516,In_964);
nand U4772 (N_4772,In_2781,In_1050);
nor U4773 (N_4773,In_789,In_163);
and U4774 (N_4774,In_617,In_2623);
nand U4775 (N_4775,In_2105,In_2622);
or U4776 (N_4776,In_1199,In_1018);
nor U4777 (N_4777,In_1195,In_1088);
or U4778 (N_4778,In_2676,In_1732);
and U4779 (N_4779,In_1254,In_2083);
nand U4780 (N_4780,In_2924,In_2363);
and U4781 (N_4781,In_471,In_1152);
nand U4782 (N_4782,In_11,In_1380);
nor U4783 (N_4783,In_1174,In_118);
nand U4784 (N_4784,In_1556,In_1967);
nand U4785 (N_4785,In_2376,In_2851);
and U4786 (N_4786,In_730,In_1314);
nor U4787 (N_4787,In_1226,In_149);
and U4788 (N_4788,In_2100,In_1698);
or U4789 (N_4789,In_1916,In_2787);
nand U4790 (N_4790,In_836,In_1439);
and U4791 (N_4791,In_2018,In_1439);
nand U4792 (N_4792,In_1393,In_1799);
nand U4793 (N_4793,In_1465,In_238);
and U4794 (N_4794,In_1432,In_1940);
nand U4795 (N_4795,In_1898,In_1888);
nand U4796 (N_4796,In_2060,In_538);
nor U4797 (N_4797,In_600,In_558);
or U4798 (N_4798,In_370,In_1289);
and U4799 (N_4799,In_2557,In_1599);
and U4800 (N_4800,In_35,In_1270);
nand U4801 (N_4801,In_2188,In_1770);
or U4802 (N_4802,In_1047,In_2746);
nand U4803 (N_4803,In_2753,In_2841);
nand U4804 (N_4804,In_9,In_152);
or U4805 (N_4805,In_1486,In_2911);
or U4806 (N_4806,In_1246,In_1406);
and U4807 (N_4807,In_1534,In_826);
nor U4808 (N_4808,In_2809,In_427);
or U4809 (N_4809,In_712,In_298);
or U4810 (N_4810,In_2825,In_877);
nor U4811 (N_4811,In_2716,In_1758);
and U4812 (N_4812,In_2575,In_2587);
nor U4813 (N_4813,In_1033,In_2013);
nand U4814 (N_4814,In_1677,In_2569);
nand U4815 (N_4815,In_990,In_1594);
or U4816 (N_4816,In_549,In_994);
or U4817 (N_4817,In_2780,In_2884);
nand U4818 (N_4818,In_1536,In_1980);
or U4819 (N_4819,In_1293,In_1218);
nor U4820 (N_4820,In_2152,In_621);
nor U4821 (N_4821,In_1672,In_972);
nor U4822 (N_4822,In_2924,In_1690);
or U4823 (N_4823,In_1312,In_1696);
nand U4824 (N_4824,In_2022,In_682);
or U4825 (N_4825,In_877,In_2349);
or U4826 (N_4826,In_334,In_651);
or U4827 (N_4827,In_655,In_2456);
or U4828 (N_4828,In_1140,In_64);
nand U4829 (N_4829,In_1859,In_2506);
and U4830 (N_4830,In_2619,In_2579);
xor U4831 (N_4831,In_193,In_2522);
nand U4832 (N_4832,In_1711,In_188);
nand U4833 (N_4833,In_916,In_1628);
nand U4834 (N_4834,In_1178,In_1726);
or U4835 (N_4835,In_1707,In_2840);
nor U4836 (N_4836,In_2499,In_2850);
nor U4837 (N_4837,In_2881,In_2959);
and U4838 (N_4838,In_1445,In_750);
nand U4839 (N_4839,In_1317,In_613);
or U4840 (N_4840,In_990,In_153);
nand U4841 (N_4841,In_690,In_648);
and U4842 (N_4842,In_2717,In_1338);
nand U4843 (N_4843,In_1763,In_536);
or U4844 (N_4844,In_291,In_2672);
or U4845 (N_4845,In_1881,In_670);
and U4846 (N_4846,In_2839,In_2011);
nand U4847 (N_4847,In_1947,In_965);
nor U4848 (N_4848,In_682,In_1729);
and U4849 (N_4849,In_437,In_1131);
nor U4850 (N_4850,In_357,In_2061);
and U4851 (N_4851,In_444,In_2248);
nand U4852 (N_4852,In_1219,In_2020);
nand U4853 (N_4853,In_1358,In_1017);
nor U4854 (N_4854,In_143,In_1064);
and U4855 (N_4855,In_297,In_126);
and U4856 (N_4856,In_2469,In_604);
nand U4857 (N_4857,In_606,In_557);
or U4858 (N_4858,In_2581,In_2649);
and U4859 (N_4859,In_916,In_2524);
nor U4860 (N_4860,In_1643,In_2029);
or U4861 (N_4861,In_203,In_1963);
nor U4862 (N_4862,In_53,In_2636);
nor U4863 (N_4863,In_2033,In_833);
nor U4864 (N_4864,In_141,In_632);
nand U4865 (N_4865,In_266,In_2988);
nor U4866 (N_4866,In_398,In_1820);
or U4867 (N_4867,In_56,In_421);
nor U4868 (N_4868,In_1628,In_424);
nor U4869 (N_4869,In_1004,In_2076);
and U4870 (N_4870,In_1545,In_1036);
nand U4871 (N_4871,In_2146,In_425);
or U4872 (N_4872,In_2529,In_841);
nand U4873 (N_4873,In_2976,In_2180);
and U4874 (N_4874,In_2037,In_2589);
and U4875 (N_4875,In_772,In_188);
and U4876 (N_4876,In_2789,In_714);
and U4877 (N_4877,In_935,In_2832);
or U4878 (N_4878,In_2124,In_904);
and U4879 (N_4879,In_513,In_2353);
nand U4880 (N_4880,In_2312,In_1821);
or U4881 (N_4881,In_181,In_2057);
nand U4882 (N_4882,In_542,In_1973);
or U4883 (N_4883,In_2462,In_1714);
nor U4884 (N_4884,In_1554,In_1501);
or U4885 (N_4885,In_1828,In_750);
nand U4886 (N_4886,In_503,In_470);
nor U4887 (N_4887,In_2936,In_302);
nor U4888 (N_4888,In_2447,In_2847);
or U4889 (N_4889,In_2270,In_2080);
nand U4890 (N_4890,In_591,In_688);
and U4891 (N_4891,In_357,In_869);
nor U4892 (N_4892,In_90,In_1093);
and U4893 (N_4893,In_2739,In_2158);
nor U4894 (N_4894,In_2185,In_2995);
or U4895 (N_4895,In_485,In_2992);
or U4896 (N_4896,In_1846,In_2533);
nor U4897 (N_4897,In_76,In_1903);
or U4898 (N_4898,In_278,In_2431);
or U4899 (N_4899,In_2685,In_1761);
and U4900 (N_4900,In_2919,In_2429);
nand U4901 (N_4901,In_1881,In_422);
nor U4902 (N_4902,In_395,In_2402);
or U4903 (N_4903,In_852,In_2093);
nand U4904 (N_4904,In_81,In_1437);
nor U4905 (N_4905,In_2771,In_817);
or U4906 (N_4906,In_1508,In_934);
and U4907 (N_4907,In_2997,In_1356);
and U4908 (N_4908,In_1605,In_2138);
or U4909 (N_4909,In_1677,In_2071);
nor U4910 (N_4910,In_1094,In_156);
nand U4911 (N_4911,In_1492,In_1127);
or U4912 (N_4912,In_893,In_1252);
nand U4913 (N_4913,In_2675,In_2919);
nor U4914 (N_4914,In_1105,In_2111);
nand U4915 (N_4915,In_83,In_2924);
and U4916 (N_4916,In_2754,In_246);
or U4917 (N_4917,In_1513,In_2751);
nand U4918 (N_4918,In_1190,In_1583);
or U4919 (N_4919,In_1913,In_1695);
and U4920 (N_4920,In_2552,In_1928);
nor U4921 (N_4921,In_1002,In_2238);
and U4922 (N_4922,In_1906,In_2688);
and U4923 (N_4923,In_32,In_2645);
nor U4924 (N_4924,In_1520,In_933);
nor U4925 (N_4925,In_341,In_1009);
and U4926 (N_4926,In_764,In_1133);
nand U4927 (N_4927,In_2826,In_2807);
nand U4928 (N_4928,In_2318,In_1114);
and U4929 (N_4929,In_2415,In_25);
or U4930 (N_4930,In_751,In_2596);
and U4931 (N_4931,In_1206,In_2094);
and U4932 (N_4932,In_4,In_2368);
and U4933 (N_4933,In_1702,In_2373);
or U4934 (N_4934,In_787,In_115);
or U4935 (N_4935,In_1468,In_2286);
and U4936 (N_4936,In_110,In_657);
nand U4937 (N_4937,In_2960,In_1239);
or U4938 (N_4938,In_1158,In_1442);
or U4939 (N_4939,In_2111,In_2153);
xnor U4940 (N_4940,In_379,In_2860);
nand U4941 (N_4941,In_1170,In_1364);
xnor U4942 (N_4942,In_1751,In_256);
nand U4943 (N_4943,In_2062,In_1333);
and U4944 (N_4944,In_280,In_1653);
nor U4945 (N_4945,In_1704,In_150);
nand U4946 (N_4946,In_2018,In_422);
or U4947 (N_4947,In_514,In_912);
nor U4948 (N_4948,In_287,In_690);
or U4949 (N_4949,In_887,In_904);
and U4950 (N_4950,In_1568,In_1297);
nor U4951 (N_4951,In_1577,In_1738);
or U4952 (N_4952,In_1372,In_1401);
nor U4953 (N_4953,In_1846,In_1563);
nor U4954 (N_4954,In_2795,In_715);
nor U4955 (N_4955,In_957,In_623);
nor U4956 (N_4956,In_771,In_912);
or U4957 (N_4957,In_2911,In_1899);
nor U4958 (N_4958,In_1306,In_313);
or U4959 (N_4959,In_2454,In_2304);
or U4960 (N_4960,In_760,In_2689);
nor U4961 (N_4961,In_2089,In_1805);
and U4962 (N_4962,In_1530,In_2702);
and U4963 (N_4963,In_281,In_1293);
or U4964 (N_4964,In_806,In_2433);
nand U4965 (N_4965,In_2338,In_1312);
or U4966 (N_4966,In_899,In_1739);
nor U4967 (N_4967,In_1866,In_1144);
and U4968 (N_4968,In_2700,In_1626);
or U4969 (N_4969,In_1986,In_2250);
nand U4970 (N_4970,In_2404,In_258);
nand U4971 (N_4971,In_1069,In_112);
nand U4972 (N_4972,In_278,In_1955);
nand U4973 (N_4973,In_1110,In_1898);
or U4974 (N_4974,In_2713,In_1274);
nor U4975 (N_4975,In_2391,In_1087);
nor U4976 (N_4976,In_1131,In_323);
nor U4977 (N_4977,In_813,In_2242);
nand U4978 (N_4978,In_1771,In_1875);
nand U4979 (N_4979,In_2948,In_370);
or U4980 (N_4980,In_608,In_833);
nand U4981 (N_4981,In_2333,In_1460);
nor U4982 (N_4982,In_73,In_1392);
nor U4983 (N_4983,In_2208,In_1923);
nor U4984 (N_4984,In_1316,In_2693);
nand U4985 (N_4985,In_761,In_1900);
nand U4986 (N_4986,In_2291,In_2727);
and U4987 (N_4987,In_1791,In_638);
or U4988 (N_4988,In_2451,In_1165);
or U4989 (N_4989,In_1089,In_11);
nor U4990 (N_4990,In_2444,In_1017);
nand U4991 (N_4991,In_1552,In_1471);
or U4992 (N_4992,In_2716,In_1699);
or U4993 (N_4993,In_2645,In_1293);
nand U4994 (N_4994,In_862,In_1168);
nand U4995 (N_4995,In_857,In_470);
or U4996 (N_4996,In_252,In_415);
or U4997 (N_4997,In_851,In_2575);
and U4998 (N_4998,In_2062,In_507);
and U4999 (N_4999,In_411,In_1268);
or U5000 (N_5000,In_2035,In_961);
or U5001 (N_5001,In_932,In_2119);
nor U5002 (N_5002,In_2072,In_390);
or U5003 (N_5003,In_1149,In_1290);
and U5004 (N_5004,In_336,In_428);
or U5005 (N_5005,In_1477,In_1035);
or U5006 (N_5006,In_1817,In_619);
and U5007 (N_5007,In_476,In_68);
nor U5008 (N_5008,In_1986,In_2339);
nand U5009 (N_5009,In_2329,In_752);
and U5010 (N_5010,In_2192,In_2879);
xor U5011 (N_5011,In_2700,In_1728);
and U5012 (N_5012,In_2301,In_47);
nand U5013 (N_5013,In_1678,In_1775);
and U5014 (N_5014,In_914,In_281);
nor U5015 (N_5015,In_72,In_1859);
and U5016 (N_5016,In_404,In_56);
nand U5017 (N_5017,In_842,In_197);
nor U5018 (N_5018,In_2391,In_323);
or U5019 (N_5019,In_1068,In_1842);
or U5020 (N_5020,In_2133,In_220);
xnor U5021 (N_5021,In_1552,In_2413);
or U5022 (N_5022,In_741,In_1206);
or U5023 (N_5023,In_1982,In_1579);
nor U5024 (N_5024,In_952,In_625);
and U5025 (N_5025,In_1184,In_620);
nand U5026 (N_5026,In_2158,In_933);
nand U5027 (N_5027,In_1061,In_2722);
or U5028 (N_5028,In_2924,In_2534);
nand U5029 (N_5029,In_2988,In_766);
or U5030 (N_5030,In_739,In_1381);
xor U5031 (N_5031,In_2932,In_627);
or U5032 (N_5032,In_2394,In_1496);
or U5033 (N_5033,In_2519,In_2876);
and U5034 (N_5034,In_2736,In_1773);
or U5035 (N_5035,In_1962,In_1821);
and U5036 (N_5036,In_1132,In_889);
or U5037 (N_5037,In_79,In_2816);
nand U5038 (N_5038,In_2815,In_469);
nor U5039 (N_5039,In_2239,In_156);
and U5040 (N_5040,In_1605,In_1591);
xor U5041 (N_5041,In_1846,In_440);
nand U5042 (N_5042,In_2661,In_1412);
or U5043 (N_5043,In_1826,In_29);
or U5044 (N_5044,In_919,In_2662);
and U5045 (N_5045,In_1519,In_1980);
nand U5046 (N_5046,In_1590,In_1520);
or U5047 (N_5047,In_1141,In_2381);
and U5048 (N_5048,In_2604,In_260);
nor U5049 (N_5049,In_366,In_878);
nor U5050 (N_5050,In_73,In_1374);
and U5051 (N_5051,In_2143,In_1078);
nand U5052 (N_5052,In_1253,In_1747);
nor U5053 (N_5053,In_672,In_1711);
or U5054 (N_5054,In_743,In_2662);
nor U5055 (N_5055,In_1165,In_2115);
nand U5056 (N_5056,In_1796,In_2036);
xor U5057 (N_5057,In_886,In_371);
or U5058 (N_5058,In_2530,In_1755);
nor U5059 (N_5059,In_2508,In_2802);
nor U5060 (N_5060,In_386,In_517);
and U5061 (N_5061,In_2813,In_865);
or U5062 (N_5062,In_616,In_1472);
or U5063 (N_5063,In_2067,In_1028);
or U5064 (N_5064,In_1101,In_2583);
nor U5065 (N_5065,In_267,In_728);
or U5066 (N_5066,In_348,In_2729);
and U5067 (N_5067,In_555,In_708);
and U5068 (N_5068,In_1114,In_1754);
or U5069 (N_5069,In_558,In_1469);
and U5070 (N_5070,In_1712,In_365);
nand U5071 (N_5071,In_1312,In_881);
or U5072 (N_5072,In_2398,In_1291);
and U5073 (N_5073,In_399,In_2338);
nand U5074 (N_5074,In_1405,In_1745);
nor U5075 (N_5075,In_2974,In_135);
nand U5076 (N_5076,In_2366,In_1643);
and U5077 (N_5077,In_1973,In_1933);
nor U5078 (N_5078,In_2538,In_1872);
and U5079 (N_5079,In_2900,In_560);
nand U5080 (N_5080,In_105,In_1604);
nor U5081 (N_5081,In_1395,In_1811);
nor U5082 (N_5082,In_2079,In_1600);
and U5083 (N_5083,In_2066,In_2228);
nand U5084 (N_5084,In_947,In_2621);
or U5085 (N_5085,In_2608,In_499);
or U5086 (N_5086,In_1621,In_2373);
and U5087 (N_5087,In_1214,In_2945);
or U5088 (N_5088,In_1395,In_838);
and U5089 (N_5089,In_308,In_2156);
nand U5090 (N_5090,In_2906,In_181);
or U5091 (N_5091,In_2606,In_622);
nor U5092 (N_5092,In_1768,In_1143);
or U5093 (N_5093,In_2105,In_2629);
nor U5094 (N_5094,In_1822,In_2075);
nor U5095 (N_5095,In_1090,In_2334);
nor U5096 (N_5096,In_2866,In_834);
nand U5097 (N_5097,In_2889,In_1817);
nor U5098 (N_5098,In_1017,In_2437);
nand U5099 (N_5099,In_2983,In_2672);
nor U5100 (N_5100,In_1223,In_554);
and U5101 (N_5101,In_2605,In_539);
nand U5102 (N_5102,In_941,In_2580);
nand U5103 (N_5103,In_2935,In_1071);
and U5104 (N_5104,In_1117,In_952);
and U5105 (N_5105,In_1421,In_11);
and U5106 (N_5106,In_2228,In_1635);
or U5107 (N_5107,In_253,In_1248);
nor U5108 (N_5108,In_930,In_2529);
nor U5109 (N_5109,In_1424,In_423);
or U5110 (N_5110,In_380,In_1956);
or U5111 (N_5111,In_1571,In_2504);
and U5112 (N_5112,In_291,In_1195);
and U5113 (N_5113,In_1886,In_2647);
or U5114 (N_5114,In_623,In_2547);
nand U5115 (N_5115,In_725,In_2368);
nand U5116 (N_5116,In_2215,In_1609);
nand U5117 (N_5117,In_1811,In_1794);
or U5118 (N_5118,In_1452,In_807);
or U5119 (N_5119,In_494,In_926);
and U5120 (N_5120,In_2590,In_2342);
and U5121 (N_5121,In_2876,In_303);
or U5122 (N_5122,In_1076,In_1552);
nor U5123 (N_5123,In_1834,In_2849);
or U5124 (N_5124,In_327,In_2412);
or U5125 (N_5125,In_2888,In_2925);
nand U5126 (N_5126,In_996,In_2479);
or U5127 (N_5127,In_2048,In_2291);
and U5128 (N_5128,In_96,In_2925);
nor U5129 (N_5129,In_1506,In_1823);
and U5130 (N_5130,In_2684,In_2144);
nand U5131 (N_5131,In_1337,In_591);
nor U5132 (N_5132,In_437,In_102);
or U5133 (N_5133,In_2593,In_2296);
nand U5134 (N_5134,In_2741,In_2930);
nand U5135 (N_5135,In_1254,In_1154);
or U5136 (N_5136,In_760,In_737);
or U5137 (N_5137,In_2648,In_2296);
and U5138 (N_5138,In_1219,In_505);
nand U5139 (N_5139,In_1018,In_2923);
nor U5140 (N_5140,In_1529,In_1352);
or U5141 (N_5141,In_2922,In_512);
and U5142 (N_5142,In_2712,In_2909);
or U5143 (N_5143,In_812,In_1268);
nand U5144 (N_5144,In_1526,In_490);
or U5145 (N_5145,In_1502,In_216);
or U5146 (N_5146,In_1018,In_1964);
and U5147 (N_5147,In_2118,In_2898);
nand U5148 (N_5148,In_906,In_1302);
nor U5149 (N_5149,In_456,In_857);
nor U5150 (N_5150,In_2163,In_2753);
and U5151 (N_5151,In_2219,In_375);
and U5152 (N_5152,In_547,In_2938);
nand U5153 (N_5153,In_2021,In_2069);
or U5154 (N_5154,In_1982,In_2140);
nand U5155 (N_5155,In_2929,In_1684);
nor U5156 (N_5156,In_1422,In_1178);
and U5157 (N_5157,In_794,In_1691);
nor U5158 (N_5158,In_1162,In_2850);
nor U5159 (N_5159,In_2037,In_666);
or U5160 (N_5160,In_1281,In_1376);
nor U5161 (N_5161,In_1406,In_1759);
and U5162 (N_5162,In_1279,In_565);
nor U5163 (N_5163,In_1841,In_764);
or U5164 (N_5164,In_813,In_465);
or U5165 (N_5165,In_454,In_1487);
nor U5166 (N_5166,In_1116,In_150);
nand U5167 (N_5167,In_38,In_2939);
and U5168 (N_5168,In_872,In_2372);
nand U5169 (N_5169,In_1739,In_2973);
and U5170 (N_5170,In_563,In_870);
nor U5171 (N_5171,In_2072,In_1666);
nand U5172 (N_5172,In_701,In_2586);
or U5173 (N_5173,In_2821,In_2097);
or U5174 (N_5174,In_2119,In_1349);
nor U5175 (N_5175,In_1547,In_512);
nor U5176 (N_5176,In_2725,In_577);
nand U5177 (N_5177,In_2771,In_1055);
and U5178 (N_5178,In_2012,In_1097);
and U5179 (N_5179,In_2429,In_2112);
nand U5180 (N_5180,In_1502,In_1374);
nand U5181 (N_5181,In_2438,In_2926);
or U5182 (N_5182,In_849,In_8);
or U5183 (N_5183,In_109,In_2514);
or U5184 (N_5184,In_2517,In_1935);
nand U5185 (N_5185,In_2128,In_2360);
nand U5186 (N_5186,In_2644,In_2667);
nand U5187 (N_5187,In_2588,In_1912);
nor U5188 (N_5188,In_1413,In_2967);
nand U5189 (N_5189,In_791,In_2858);
or U5190 (N_5190,In_2235,In_2323);
nor U5191 (N_5191,In_1841,In_624);
nor U5192 (N_5192,In_1696,In_2776);
nor U5193 (N_5193,In_2846,In_129);
nor U5194 (N_5194,In_504,In_681);
nor U5195 (N_5195,In_666,In_2827);
nand U5196 (N_5196,In_2020,In_601);
nand U5197 (N_5197,In_19,In_1078);
nor U5198 (N_5198,In_2323,In_2268);
or U5199 (N_5199,In_1162,In_2617);
or U5200 (N_5200,In_2188,In_1987);
nand U5201 (N_5201,In_2764,In_2570);
nor U5202 (N_5202,In_1141,In_1273);
or U5203 (N_5203,In_921,In_489);
xor U5204 (N_5204,In_1551,In_1538);
or U5205 (N_5205,In_132,In_1657);
or U5206 (N_5206,In_175,In_187);
xor U5207 (N_5207,In_2441,In_1805);
nand U5208 (N_5208,In_380,In_1349);
and U5209 (N_5209,In_653,In_2164);
nand U5210 (N_5210,In_1688,In_142);
and U5211 (N_5211,In_2755,In_870);
and U5212 (N_5212,In_1027,In_2962);
nand U5213 (N_5213,In_2190,In_2276);
or U5214 (N_5214,In_2828,In_1542);
nor U5215 (N_5215,In_1435,In_1427);
and U5216 (N_5216,In_1080,In_2381);
and U5217 (N_5217,In_1077,In_2110);
and U5218 (N_5218,In_77,In_469);
nand U5219 (N_5219,In_1847,In_1495);
and U5220 (N_5220,In_2149,In_2192);
nand U5221 (N_5221,In_1200,In_62);
and U5222 (N_5222,In_866,In_227);
nor U5223 (N_5223,In_1414,In_201);
nand U5224 (N_5224,In_2844,In_1206);
and U5225 (N_5225,In_1862,In_1488);
nand U5226 (N_5226,In_1134,In_850);
and U5227 (N_5227,In_819,In_0);
nor U5228 (N_5228,In_1802,In_2987);
nand U5229 (N_5229,In_175,In_762);
or U5230 (N_5230,In_2539,In_2534);
or U5231 (N_5231,In_640,In_1328);
nor U5232 (N_5232,In_1029,In_1608);
nand U5233 (N_5233,In_1058,In_2047);
nor U5234 (N_5234,In_1766,In_180);
and U5235 (N_5235,In_1420,In_282);
nor U5236 (N_5236,In_1028,In_106);
and U5237 (N_5237,In_1391,In_1141);
and U5238 (N_5238,In_2760,In_325);
or U5239 (N_5239,In_1119,In_2894);
nor U5240 (N_5240,In_544,In_2876);
nand U5241 (N_5241,In_2453,In_206);
nand U5242 (N_5242,In_2037,In_831);
or U5243 (N_5243,In_157,In_248);
or U5244 (N_5244,In_2974,In_1321);
nand U5245 (N_5245,In_1792,In_10);
nand U5246 (N_5246,In_2768,In_2719);
or U5247 (N_5247,In_1530,In_1231);
or U5248 (N_5248,In_2627,In_109);
nor U5249 (N_5249,In_2286,In_1682);
or U5250 (N_5250,In_320,In_58);
and U5251 (N_5251,In_1963,In_1696);
nor U5252 (N_5252,In_549,In_133);
nand U5253 (N_5253,In_974,In_1458);
or U5254 (N_5254,In_1745,In_2041);
xnor U5255 (N_5255,In_2066,In_2417);
nand U5256 (N_5256,In_2569,In_303);
and U5257 (N_5257,In_1854,In_2997);
nor U5258 (N_5258,In_615,In_2127);
and U5259 (N_5259,In_113,In_2698);
or U5260 (N_5260,In_2934,In_276);
and U5261 (N_5261,In_2946,In_2390);
and U5262 (N_5262,In_159,In_1987);
or U5263 (N_5263,In_2089,In_2383);
and U5264 (N_5264,In_2255,In_2449);
or U5265 (N_5265,In_2094,In_2564);
or U5266 (N_5266,In_2510,In_568);
nand U5267 (N_5267,In_1209,In_2996);
nand U5268 (N_5268,In_1507,In_1939);
nor U5269 (N_5269,In_301,In_2515);
nor U5270 (N_5270,In_1562,In_2888);
or U5271 (N_5271,In_2061,In_2395);
or U5272 (N_5272,In_392,In_1362);
or U5273 (N_5273,In_2178,In_462);
nand U5274 (N_5274,In_1271,In_2916);
nand U5275 (N_5275,In_1814,In_218);
and U5276 (N_5276,In_2768,In_1110);
nor U5277 (N_5277,In_1696,In_2672);
nand U5278 (N_5278,In_2803,In_1876);
nor U5279 (N_5279,In_1220,In_1121);
nor U5280 (N_5280,In_753,In_2840);
nor U5281 (N_5281,In_1420,In_1535);
nand U5282 (N_5282,In_1545,In_1038);
and U5283 (N_5283,In_618,In_2464);
nor U5284 (N_5284,In_988,In_1264);
nand U5285 (N_5285,In_731,In_1963);
and U5286 (N_5286,In_1508,In_2673);
nor U5287 (N_5287,In_1364,In_904);
nor U5288 (N_5288,In_184,In_2245);
and U5289 (N_5289,In_1737,In_168);
or U5290 (N_5290,In_2349,In_1943);
or U5291 (N_5291,In_2284,In_261);
or U5292 (N_5292,In_503,In_1050);
and U5293 (N_5293,In_128,In_2437);
nor U5294 (N_5294,In_1437,In_1195);
or U5295 (N_5295,In_2973,In_351);
or U5296 (N_5296,In_2018,In_2863);
or U5297 (N_5297,In_2439,In_879);
nand U5298 (N_5298,In_1755,In_670);
nand U5299 (N_5299,In_1430,In_166);
xor U5300 (N_5300,In_62,In_1276);
or U5301 (N_5301,In_1432,In_859);
and U5302 (N_5302,In_702,In_1721);
nand U5303 (N_5303,In_1658,In_1029);
nor U5304 (N_5304,In_370,In_1322);
nand U5305 (N_5305,In_927,In_953);
nor U5306 (N_5306,In_2771,In_849);
nand U5307 (N_5307,In_1750,In_2524);
nor U5308 (N_5308,In_358,In_328);
and U5309 (N_5309,In_1688,In_775);
nor U5310 (N_5310,In_2899,In_1854);
nor U5311 (N_5311,In_2077,In_2347);
nor U5312 (N_5312,In_1004,In_1349);
and U5313 (N_5313,In_2061,In_204);
or U5314 (N_5314,In_260,In_2230);
or U5315 (N_5315,In_2338,In_2337);
nand U5316 (N_5316,In_2098,In_1570);
and U5317 (N_5317,In_975,In_493);
nor U5318 (N_5318,In_806,In_744);
and U5319 (N_5319,In_1177,In_2092);
or U5320 (N_5320,In_2271,In_2752);
nand U5321 (N_5321,In_1798,In_2501);
and U5322 (N_5322,In_379,In_912);
nand U5323 (N_5323,In_716,In_1673);
nand U5324 (N_5324,In_2909,In_2025);
and U5325 (N_5325,In_2565,In_206);
or U5326 (N_5326,In_2787,In_2390);
nand U5327 (N_5327,In_2563,In_2344);
and U5328 (N_5328,In_1227,In_442);
or U5329 (N_5329,In_1088,In_2356);
nor U5330 (N_5330,In_291,In_1859);
and U5331 (N_5331,In_2221,In_2263);
nor U5332 (N_5332,In_2064,In_2230);
or U5333 (N_5333,In_2961,In_2046);
nor U5334 (N_5334,In_353,In_623);
nor U5335 (N_5335,In_1961,In_2882);
nand U5336 (N_5336,In_739,In_879);
and U5337 (N_5337,In_236,In_2450);
nor U5338 (N_5338,In_1340,In_1812);
and U5339 (N_5339,In_675,In_373);
and U5340 (N_5340,In_5,In_859);
nor U5341 (N_5341,In_1276,In_1789);
nand U5342 (N_5342,In_1465,In_1709);
or U5343 (N_5343,In_886,In_1737);
or U5344 (N_5344,In_1513,In_190);
nand U5345 (N_5345,In_1242,In_2076);
and U5346 (N_5346,In_1429,In_2818);
or U5347 (N_5347,In_56,In_2249);
nor U5348 (N_5348,In_566,In_1951);
xor U5349 (N_5349,In_1715,In_1836);
or U5350 (N_5350,In_2780,In_726);
and U5351 (N_5351,In_2253,In_1003);
and U5352 (N_5352,In_2420,In_472);
or U5353 (N_5353,In_1683,In_1892);
nand U5354 (N_5354,In_883,In_2285);
nor U5355 (N_5355,In_292,In_690);
and U5356 (N_5356,In_1469,In_44);
nand U5357 (N_5357,In_2763,In_1682);
nand U5358 (N_5358,In_20,In_1351);
or U5359 (N_5359,In_105,In_1767);
or U5360 (N_5360,In_2436,In_1429);
nand U5361 (N_5361,In_1435,In_2444);
nand U5362 (N_5362,In_969,In_493);
xnor U5363 (N_5363,In_1420,In_590);
nand U5364 (N_5364,In_2636,In_1613);
or U5365 (N_5365,In_2624,In_1210);
and U5366 (N_5366,In_1187,In_1721);
nor U5367 (N_5367,In_2935,In_1699);
nand U5368 (N_5368,In_656,In_477);
nand U5369 (N_5369,In_2752,In_2302);
nor U5370 (N_5370,In_49,In_1736);
nand U5371 (N_5371,In_2982,In_638);
and U5372 (N_5372,In_577,In_2186);
and U5373 (N_5373,In_1234,In_1531);
nand U5374 (N_5374,In_388,In_215);
and U5375 (N_5375,In_1242,In_1208);
nor U5376 (N_5376,In_252,In_1125);
or U5377 (N_5377,In_1387,In_755);
and U5378 (N_5378,In_1465,In_1588);
nor U5379 (N_5379,In_283,In_354);
nand U5380 (N_5380,In_461,In_440);
or U5381 (N_5381,In_370,In_458);
nand U5382 (N_5382,In_799,In_338);
and U5383 (N_5383,In_427,In_2614);
nand U5384 (N_5384,In_729,In_1330);
or U5385 (N_5385,In_2595,In_1370);
and U5386 (N_5386,In_2027,In_2909);
nor U5387 (N_5387,In_212,In_1347);
nor U5388 (N_5388,In_1046,In_2997);
or U5389 (N_5389,In_2881,In_1719);
and U5390 (N_5390,In_2091,In_2377);
nand U5391 (N_5391,In_1255,In_1493);
or U5392 (N_5392,In_179,In_1398);
and U5393 (N_5393,In_1972,In_1229);
and U5394 (N_5394,In_358,In_880);
nor U5395 (N_5395,In_1615,In_967);
or U5396 (N_5396,In_214,In_2349);
nor U5397 (N_5397,In_746,In_2755);
or U5398 (N_5398,In_2424,In_754);
and U5399 (N_5399,In_2574,In_1028);
nand U5400 (N_5400,In_1089,In_1020);
or U5401 (N_5401,In_480,In_566);
or U5402 (N_5402,In_1285,In_2089);
and U5403 (N_5403,In_397,In_2639);
nand U5404 (N_5404,In_1650,In_1651);
and U5405 (N_5405,In_2494,In_2697);
nand U5406 (N_5406,In_2883,In_1569);
nand U5407 (N_5407,In_983,In_1373);
or U5408 (N_5408,In_1129,In_1729);
nor U5409 (N_5409,In_1651,In_901);
nand U5410 (N_5410,In_2548,In_1025);
nand U5411 (N_5411,In_2753,In_2869);
and U5412 (N_5412,In_2348,In_1276);
nand U5413 (N_5413,In_2383,In_1048);
and U5414 (N_5414,In_2591,In_628);
and U5415 (N_5415,In_844,In_1461);
and U5416 (N_5416,In_2887,In_1119);
nand U5417 (N_5417,In_1488,In_1476);
nor U5418 (N_5418,In_1776,In_274);
nand U5419 (N_5419,In_660,In_2347);
nand U5420 (N_5420,In_921,In_979);
nand U5421 (N_5421,In_2015,In_975);
and U5422 (N_5422,In_2254,In_857);
nor U5423 (N_5423,In_1544,In_2065);
and U5424 (N_5424,In_2489,In_1421);
nand U5425 (N_5425,In_426,In_419);
or U5426 (N_5426,In_1594,In_184);
and U5427 (N_5427,In_2674,In_2164);
nand U5428 (N_5428,In_157,In_240);
nand U5429 (N_5429,In_1183,In_1340);
nor U5430 (N_5430,In_2852,In_53);
or U5431 (N_5431,In_137,In_1181);
and U5432 (N_5432,In_440,In_1188);
or U5433 (N_5433,In_2816,In_2858);
nor U5434 (N_5434,In_2819,In_2480);
and U5435 (N_5435,In_1752,In_1288);
and U5436 (N_5436,In_2633,In_2566);
or U5437 (N_5437,In_1214,In_2123);
and U5438 (N_5438,In_1390,In_798);
or U5439 (N_5439,In_2073,In_2499);
and U5440 (N_5440,In_2423,In_155);
nor U5441 (N_5441,In_131,In_581);
and U5442 (N_5442,In_2121,In_2745);
or U5443 (N_5443,In_2358,In_546);
or U5444 (N_5444,In_391,In_1413);
xnor U5445 (N_5445,In_2588,In_1971);
or U5446 (N_5446,In_1910,In_915);
and U5447 (N_5447,In_2430,In_1400);
nor U5448 (N_5448,In_2910,In_2417);
or U5449 (N_5449,In_1188,In_2348);
or U5450 (N_5450,In_451,In_2057);
nor U5451 (N_5451,In_1650,In_353);
or U5452 (N_5452,In_2670,In_91);
nor U5453 (N_5453,In_386,In_2081);
nand U5454 (N_5454,In_1419,In_661);
nand U5455 (N_5455,In_1853,In_1404);
or U5456 (N_5456,In_1465,In_1896);
nor U5457 (N_5457,In_1792,In_615);
and U5458 (N_5458,In_640,In_1672);
or U5459 (N_5459,In_2087,In_2984);
nor U5460 (N_5460,In_984,In_50);
and U5461 (N_5461,In_1131,In_943);
nor U5462 (N_5462,In_2306,In_840);
nor U5463 (N_5463,In_2494,In_1020);
or U5464 (N_5464,In_1991,In_1209);
nor U5465 (N_5465,In_1420,In_1808);
and U5466 (N_5466,In_804,In_642);
nand U5467 (N_5467,In_800,In_797);
nor U5468 (N_5468,In_725,In_1375);
or U5469 (N_5469,In_1026,In_755);
nand U5470 (N_5470,In_2670,In_2426);
and U5471 (N_5471,In_1473,In_608);
or U5472 (N_5472,In_1700,In_265);
xnor U5473 (N_5473,In_2367,In_765);
or U5474 (N_5474,In_283,In_760);
nor U5475 (N_5475,In_1730,In_2130);
and U5476 (N_5476,In_2480,In_548);
and U5477 (N_5477,In_2226,In_254);
or U5478 (N_5478,In_23,In_2254);
and U5479 (N_5479,In_620,In_2769);
nor U5480 (N_5480,In_1609,In_817);
and U5481 (N_5481,In_2852,In_884);
and U5482 (N_5482,In_470,In_2242);
and U5483 (N_5483,In_1920,In_342);
nor U5484 (N_5484,In_208,In_1091);
or U5485 (N_5485,In_2601,In_2998);
or U5486 (N_5486,In_493,In_2368);
nand U5487 (N_5487,In_1902,In_1990);
nand U5488 (N_5488,In_1610,In_1326);
nand U5489 (N_5489,In_880,In_1856);
and U5490 (N_5490,In_1101,In_1575);
nand U5491 (N_5491,In_2533,In_1022);
nor U5492 (N_5492,In_2077,In_89);
nor U5493 (N_5493,In_336,In_2912);
and U5494 (N_5494,In_2663,In_2855);
nand U5495 (N_5495,In_894,In_1873);
and U5496 (N_5496,In_1762,In_2953);
and U5497 (N_5497,In_1097,In_2079);
nor U5498 (N_5498,In_376,In_1121);
and U5499 (N_5499,In_2864,In_842);
nor U5500 (N_5500,In_2533,In_2471);
nor U5501 (N_5501,In_1729,In_117);
nand U5502 (N_5502,In_868,In_2171);
or U5503 (N_5503,In_1099,In_1333);
nand U5504 (N_5504,In_2818,In_726);
nor U5505 (N_5505,In_1146,In_614);
and U5506 (N_5506,In_1054,In_2858);
nand U5507 (N_5507,In_1689,In_498);
or U5508 (N_5508,In_1411,In_471);
or U5509 (N_5509,In_173,In_686);
or U5510 (N_5510,In_2568,In_1108);
nand U5511 (N_5511,In_1862,In_2565);
or U5512 (N_5512,In_2718,In_1603);
and U5513 (N_5513,In_287,In_359);
nor U5514 (N_5514,In_610,In_2815);
nand U5515 (N_5515,In_943,In_676);
xnor U5516 (N_5516,In_1351,In_1428);
or U5517 (N_5517,In_2898,In_1476);
nor U5518 (N_5518,In_2717,In_1470);
nand U5519 (N_5519,In_1148,In_1433);
nor U5520 (N_5520,In_2554,In_2199);
or U5521 (N_5521,In_1683,In_1393);
nand U5522 (N_5522,In_336,In_2450);
and U5523 (N_5523,In_2461,In_294);
nand U5524 (N_5524,In_1498,In_779);
or U5525 (N_5525,In_1887,In_1270);
and U5526 (N_5526,In_2333,In_1892);
and U5527 (N_5527,In_2391,In_2889);
nand U5528 (N_5528,In_2847,In_2189);
or U5529 (N_5529,In_2130,In_511);
nor U5530 (N_5530,In_2216,In_2927);
and U5531 (N_5531,In_1270,In_1039);
nand U5532 (N_5532,In_395,In_872);
xor U5533 (N_5533,In_2157,In_385);
or U5534 (N_5534,In_2815,In_2247);
or U5535 (N_5535,In_213,In_2911);
or U5536 (N_5536,In_1620,In_2172);
and U5537 (N_5537,In_948,In_1495);
nor U5538 (N_5538,In_1793,In_2962);
and U5539 (N_5539,In_448,In_2213);
or U5540 (N_5540,In_90,In_1350);
nand U5541 (N_5541,In_2127,In_2627);
or U5542 (N_5542,In_997,In_2705);
nor U5543 (N_5543,In_817,In_96);
or U5544 (N_5544,In_1219,In_654);
nor U5545 (N_5545,In_860,In_2258);
nor U5546 (N_5546,In_162,In_132);
nand U5547 (N_5547,In_2336,In_1901);
nor U5548 (N_5548,In_838,In_818);
nand U5549 (N_5549,In_2792,In_797);
or U5550 (N_5550,In_2557,In_224);
and U5551 (N_5551,In_2848,In_1303);
nand U5552 (N_5552,In_280,In_2996);
or U5553 (N_5553,In_1891,In_996);
and U5554 (N_5554,In_201,In_2341);
nor U5555 (N_5555,In_1637,In_2604);
or U5556 (N_5556,In_15,In_106);
or U5557 (N_5557,In_36,In_1938);
nor U5558 (N_5558,In_261,In_1052);
or U5559 (N_5559,In_2551,In_1236);
nor U5560 (N_5560,In_2748,In_1087);
and U5561 (N_5561,In_1913,In_1461);
nand U5562 (N_5562,In_508,In_1876);
or U5563 (N_5563,In_2249,In_582);
nand U5564 (N_5564,In_328,In_986);
nand U5565 (N_5565,In_1425,In_1108);
or U5566 (N_5566,In_1660,In_1667);
nand U5567 (N_5567,In_2071,In_2775);
nor U5568 (N_5568,In_324,In_245);
xor U5569 (N_5569,In_2487,In_1642);
nand U5570 (N_5570,In_2955,In_1679);
and U5571 (N_5571,In_1815,In_1209);
nor U5572 (N_5572,In_1814,In_336);
and U5573 (N_5573,In_873,In_1479);
nand U5574 (N_5574,In_2116,In_1849);
and U5575 (N_5575,In_338,In_2314);
or U5576 (N_5576,In_194,In_1471);
and U5577 (N_5577,In_2396,In_1848);
or U5578 (N_5578,In_1837,In_2662);
and U5579 (N_5579,In_177,In_1371);
or U5580 (N_5580,In_1251,In_40);
nor U5581 (N_5581,In_2238,In_1917);
nor U5582 (N_5582,In_683,In_2970);
xor U5583 (N_5583,In_150,In_2437);
and U5584 (N_5584,In_2242,In_2713);
xnor U5585 (N_5585,In_1366,In_1798);
nor U5586 (N_5586,In_2409,In_1683);
nand U5587 (N_5587,In_1183,In_255);
or U5588 (N_5588,In_2099,In_1328);
nand U5589 (N_5589,In_1386,In_2461);
or U5590 (N_5590,In_2475,In_1476);
nor U5591 (N_5591,In_2005,In_2079);
nand U5592 (N_5592,In_2585,In_754);
nand U5593 (N_5593,In_2902,In_2875);
nor U5594 (N_5594,In_544,In_2896);
nor U5595 (N_5595,In_1264,In_797);
and U5596 (N_5596,In_2519,In_1943);
nand U5597 (N_5597,In_1966,In_1328);
and U5598 (N_5598,In_112,In_67);
and U5599 (N_5599,In_2194,In_744);
nor U5600 (N_5600,In_2079,In_2885);
nor U5601 (N_5601,In_2620,In_2255);
nor U5602 (N_5602,In_145,In_1205);
nand U5603 (N_5603,In_1171,In_121);
nor U5604 (N_5604,In_399,In_730);
or U5605 (N_5605,In_2535,In_1272);
nor U5606 (N_5606,In_2901,In_2357);
or U5607 (N_5607,In_302,In_2360);
and U5608 (N_5608,In_2198,In_1186);
and U5609 (N_5609,In_1140,In_713);
or U5610 (N_5610,In_2572,In_180);
and U5611 (N_5611,In_944,In_98);
nor U5612 (N_5612,In_84,In_991);
or U5613 (N_5613,In_2417,In_2823);
or U5614 (N_5614,In_451,In_762);
and U5615 (N_5615,In_2047,In_1745);
nor U5616 (N_5616,In_2352,In_2696);
nand U5617 (N_5617,In_527,In_274);
nor U5618 (N_5618,In_912,In_2597);
nand U5619 (N_5619,In_2201,In_2458);
nand U5620 (N_5620,In_2467,In_2459);
nand U5621 (N_5621,In_2685,In_308);
and U5622 (N_5622,In_2872,In_780);
or U5623 (N_5623,In_833,In_2794);
or U5624 (N_5624,In_1238,In_2560);
nor U5625 (N_5625,In_2829,In_2049);
nand U5626 (N_5626,In_1217,In_1410);
and U5627 (N_5627,In_213,In_2967);
or U5628 (N_5628,In_1669,In_2425);
and U5629 (N_5629,In_1233,In_445);
or U5630 (N_5630,In_2291,In_891);
or U5631 (N_5631,In_1350,In_2040);
and U5632 (N_5632,In_896,In_2561);
and U5633 (N_5633,In_29,In_98);
or U5634 (N_5634,In_840,In_112);
and U5635 (N_5635,In_2650,In_658);
and U5636 (N_5636,In_2778,In_2142);
nand U5637 (N_5637,In_2974,In_1369);
nor U5638 (N_5638,In_2966,In_2702);
nor U5639 (N_5639,In_2530,In_124);
nor U5640 (N_5640,In_180,In_482);
or U5641 (N_5641,In_1172,In_1353);
nand U5642 (N_5642,In_2446,In_1147);
nand U5643 (N_5643,In_1248,In_1837);
and U5644 (N_5644,In_2490,In_1433);
nand U5645 (N_5645,In_2083,In_1783);
and U5646 (N_5646,In_1823,In_28);
and U5647 (N_5647,In_513,In_1673);
xor U5648 (N_5648,In_1456,In_654);
nand U5649 (N_5649,In_60,In_415);
nor U5650 (N_5650,In_1300,In_1888);
nor U5651 (N_5651,In_39,In_753);
or U5652 (N_5652,In_2267,In_1315);
and U5653 (N_5653,In_2713,In_1407);
or U5654 (N_5654,In_949,In_2323);
nor U5655 (N_5655,In_1826,In_841);
or U5656 (N_5656,In_670,In_10);
and U5657 (N_5657,In_801,In_1315);
or U5658 (N_5658,In_214,In_2459);
and U5659 (N_5659,In_243,In_346);
nor U5660 (N_5660,In_1792,In_2668);
and U5661 (N_5661,In_908,In_1136);
and U5662 (N_5662,In_1585,In_2046);
nor U5663 (N_5663,In_2839,In_703);
nand U5664 (N_5664,In_1677,In_1082);
nor U5665 (N_5665,In_2335,In_1817);
or U5666 (N_5666,In_1975,In_2943);
nor U5667 (N_5667,In_2850,In_603);
nor U5668 (N_5668,In_1016,In_667);
nor U5669 (N_5669,In_2979,In_369);
and U5670 (N_5670,In_2091,In_1803);
or U5671 (N_5671,In_1388,In_224);
nand U5672 (N_5672,In_160,In_386);
or U5673 (N_5673,In_2482,In_2426);
and U5674 (N_5674,In_872,In_2927);
nor U5675 (N_5675,In_1189,In_609);
nand U5676 (N_5676,In_1705,In_2686);
or U5677 (N_5677,In_2971,In_1603);
and U5678 (N_5678,In_1269,In_1222);
nor U5679 (N_5679,In_1554,In_2601);
nand U5680 (N_5680,In_2129,In_2165);
or U5681 (N_5681,In_2984,In_1130);
or U5682 (N_5682,In_2767,In_2103);
nor U5683 (N_5683,In_506,In_2163);
or U5684 (N_5684,In_2485,In_895);
nor U5685 (N_5685,In_1361,In_570);
or U5686 (N_5686,In_2660,In_1707);
nand U5687 (N_5687,In_2495,In_109);
or U5688 (N_5688,In_1580,In_601);
or U5689 (N_5689,In_1439,In_1554);
and U5690 (N_5690,In_861,In_234);
and U5691 (N_5691,In_2560,In_794);
nor U5692 (N_5692,In_248,In_1213);
nand U5693 (N_5693,In_338,In_1171);
or U5694 (N_5694,In_852,In_2143);
nand U5695 (N_5695,In_693,In_1252);
nand U5696 (N_5696,In_1158,In_1010);
nor U5697 (N_5697,In_516,In_1883);
or U5698 (N_5698,In_732,In_453);
or U5699 (N_5699,In_1320,In_626);
and U5700 (N_5700,In_256,In_1967);
nand U5701 (N_5701,In_337,In_2004);
or U5702 (N_5702,In_1245,In_312);
and U5703 (N_5703,In_1468,In_2129);
or U5704 (N_5704,In_2349,In_2578);
nor U5705 (N_5705,In_1440,In_456);
and U5706 (N_5706,In_683,In_830);
or U5707 (N_5707,In_1833,In_764);
or U5708 (N_5708,In_2967,In_1828);
and U5709 (N_5709,In_2090,In_553);
or U5710 (N_5710,In_861,In_2259);
nor U5711 (N_5711,In_1836,In_1496);
nand U5712 (N_5712,In_1897,In_2218);
or U5713 (N_5713,In_1870,In_221);
or U5714 (N_5714,In_1153,In_1388);
and U5715 (N_5715,In_1044,In_1621);
nand U5716 (N_5716,In_693,In_1177);
and U5717 (N_5717,In_162,In_645);
and U5718 (N_5718,In_729,In_2880);
or U5719 (N_5719,In_2814,In_2562);
nor U5720 (N_5720,In_830,In_1203);
nor U5721 (N_5721,In_2741,In_1297);
nor U5722 (N_5722,In_1067,In_1168);
nor U5723 (N_5723,In_82,In_836);
and U5724 (N_5724,In_329,In_1443);
and U5725 (N_5725,In_2030,In_138);
xor U5726 (N_5726,In_2734,In_1910);
nor U5727 (N_5727,In_2859,In_1401);
nand U5728 (N_5728,In_18,In_2275);
nor U5729 (N_5729,In_1000,In_755);
nand U5730 (N_5730,In_1639,In_974);
or U5731 (N_5731,In_2004,In_1051);
or U5732 (N_5732,In_2327,In_2579);
and U5733 (N_5733,In_1370,In_1392);
and U5734 (N_5734,In_411,In_1129);
nor U5735 (N_5735,In_1237,In_1957);
nand U5736 (N_5736,In_2319,In_2071);
and U5737 (N_5737,In_2503,In_2837);
nand U5738 (N_5738,In_1908,In_2078);
and U5739 (N_5739,In_2509,In_1385);
nand U5740 (N_5740,In_1979,In_2887);
nand U5741 (N_5741,In_2788,In_1201);
or U5742 (N_5742,In_2205,In_2492);
or U5743 (N_5743,In_2950,In_1471);
nand U5744 (N_5744,In_11,In_2516);
nor U5745 (N_5745,In_456,In_1712);
nor U5746 (N_5746,In_1223,In_282);
and U5747 (N_5747,In_2845,In_2931);
and U5748 (N_5748,In_1486,In_2819);
nor U5749 (N_5749,In_2243,In_1884);
nand U5750 (N_5750,In_1911,In_77);
or U5751 (N_5751,In_207,In_817);
nand U5752 (N_5752,In_1836,In_648);
nand U5753 (N_5753,In_1161,In_435);
nand U5754 (N_5754,In_2613,In_72);
and U5755 (N_5755,In_1813,In_1799);
nor U5756 (N_5756,In_2188,In_521);
nand U5757 (N_5757,In_857,In_1712);
or U5758 (N_5758,In_2153,In_637);
nor U5759 (N_5759,In_1059,In_323);
nor U5760 (N_5760,In_1481,In_871);
and U5761 (N_5761,In_275,In_1780);
nand U5762 (N_5762,In_491,In_2008);
nand U5763 (N_5763,In_781,In_877);
nand U5764 (N_5764,In_2210,In_2840);
nor U5765 (N_5765,In_1466,In_1276);
or U5766 (N_5766,In_997,In_554);
nor U5767 (N_5767,In_731,In_2225);
nor U5768 (N_5768,In_2799,In_2294);
nand U5769 (N_5769,In_906,In_1592);
nor U5770 (N_5770,In_416,In_1846);
nand U5771 (N_5771,In_1506,In_2245);
nor U5772 (N_5772,In_1402,In_2801);
nand U5773 (N_5773,In_1159,In_257);
nor U5774 (N_5774,In_1176,In_2504);
nand U5775 (N_5775,In_1315,In_2435);
nand U5776 (N_5776,In_1632,In_1202);
and U5777 (N_5777,In_2537,In_745);
and U5778 (N_5778,In_2749,In_1811);
nand U5779 (N_5779,In_2011,In_586);
or U5780 (N_5780,In_232,In_2803);
nor U5781 (N_5781,In_636,In_1218);
or U5782 (N_5782,In_2384,In_1162);
nor U5783 (N_5783,In_1450,In_673);
nor U5784 (N_5784,In_1236,In_815);
nand U5785 (N_5785,In_2850,In_507);
nor U5786 (N_5786,In_2165,In_584);
or U5787 (N_5787,In_1220,In_2500);
nor U5788 (N_5788,In_1014,In_2480);
nor U5789 (N_5789,In_1660,In_345);
nand U5790 (N_5790,In_2777,In_1221);
and U5791 (N_5791,In_746,In_2933);
nand U5792 (N_5792,In_1323,In_78);
nor U5793 (N_5793,In_43,In_2669);
nand U5794 (N_5794,In_2288,In_2400);
and U5795 (N_5795,In_129,In_2853);
and U5796 (N_5796,In_1860,In_610);
nor U5797 (N_5797,In_1909,In_286);
nor U5798 (N_5798,In_1340,In_2984);
nand U5799 (N_5799,In_2206,In_294);
or U5800 (N_5800,In_2250,In_1892);
and U5801 (N_5801,In_787,In_2464);
or U5802 (N_5802,In_19,In_1357);
nand U5803 (N_5803,In_72,In_2397);
nand U5804 (N_5804,In_2137,In_2072);
nand U5805 (N_5805,In_1704,In_2611);
or U5806 (N_5806,In_2169,In_1236);
nand U5807 (N_5807,In_2923,In_1488);
and U5808 (N_5808,In_2901,In_1039);
or U5809 (N_5809,In_2198,In_2236);
or U5810 (N_5810,In_1491,In_2747);
nand U5811 (N_5811,In_2126,In_907);
nor U5812 (N_5812,In_163,In_2278);
or U5813 (N_5813,In_1530,In_2225);
and U5814 (N_5814,In_1364,In_2850);
nand U5815 (N_5815,In_2942,In_1722);
and U5816 (N_5816,In_1480,In_1146);
nand U5817 (N_5817,In_661,In_1061);
nand U5818 (N_5818,In_759,In_93);
nand U5819 (N_5819,In_727,In_1707);
and U5820 (N_5820,In_2621,In_561);
and U5821 (N_5821,In_1156,In_2401);
nor U5822 (N_5822,In_1130,In_268);
nor U5823 (N_5823,In_2997,In_2047);
nor U5824 (N_5824,In_594,In_2545);
and U5825 (N_5825,In_2384,In_1583);
nand U5826 (N_5826,In_2660,In_1437);
or U5827 (N_5827,In_2130,In_1319);
nor U5828 (N_5828,In_1177,In_153);
nor U5829 (N_5829,In_1324,In_2185);
nand U5830 (N_5830,In_1270,In_720);
nor U5831 (N_5831,In_2224,In_2272);
or U5832 (N_5832,In_931,In_1562);
or U5833 (N_5833,In_1242,In_949);
or U5834 (N_5834,In_416,In_131);
nor U5835 (N_5835,In_1583,In_1211);
nor U5836 (N_5836,In_1640,In_407);
nor U5837 (N_5837,In_2455,In_1877);
or U5838 (N_5838,In_737,In_2557);
or U5839 (N_5839,In_497,In_1890);
nor U5840 (N_5840,In_1945,In_1672);
or U5841 (N_5841,In_271,In_2148);
nand U5842 (N_5842,In_1017,In_1702);
nor U5843 (N_5843,In_2067,In_191);
nor U5844 (N_5844,In_1970,In_388);
nand U5845 (N_5845,In_2169,In_1316);
or U5846 (N_5846,In_1973,In_1792);
nor U5847 (N_5847,In_1164,In_1566);
or U5848 (N_5848,In_1066,In_2310);
nor U5849 (N_5849,In_2419,In_1278);
nand U5850 (N_5850,In_2192,In_2838);
and U5851 (N_5851,In_2616,In_2293);
or U5852 (N_5852,In_1681,In_1404);
or U5853 (N_5853,In_811,In_1565);
and U5854 (N_5854,In_224,In_1123);
and U5855 (N_5855,In_2413,In_859);
nor U5856 (N_5856,In_2675,In_1421);
and U5857 (N_5857,In_586,In_628);
nand U5858 (N_5858,In_2962,In_2049);
and U5859 (N_5859,In_2377,In_2219);
nor U5860 (N_5860,In_340,In_374);
nand U5861 (N_5861,In_484,In_710);
nor U5862 (N_5862,In_2654,In_380);
and U5863 (N_5863,In_790,In_2718);
nand U5864 (N_5864,In_1633,In_594);
nand U5865 (N_5865,In_2487,In_1134);
and U5866 (N_5866,In_2596,In_597);
and U5867 (N_5867,In_1128,In_1797);
or U5868 (N_5868,In_1370,In_2511);
nor U5869 (N_5869,In_1230,In_129);
or U5870 (N_5870,In_1715,In_2301);
and U5871 (N_5871,In_2342,In_1538);
and U5872 (N_5872,In_997,In_1862);
and U5873 (N_5873,In_1783,In_2832);
nand U5874 (N_5874,In_349,In_2759);
nand U5875 (N_5875,In_688,In_1859);
nor U5876 (N_5876,In_2785,In_1503);
and U5877 (N_5877,In_1427,In_2693);
or U5878 (N_5878,In_313,In_1532);
or U5879 (N_5879,In_1908,In_1837);
or U5880 (N_5880,In_1663,In_2263);
or U5881 (N_5881,In_1845,In_2775);
or U5882 (N_5882,In_1270,In_1150);
and U5883 (N_5883,In_2563,In_1480);
nand U5884 (N_5884,In_2314,In_155);
nor U5885 (N_5885,In_2386,In_2203);
nor U5886 (N_5886,In_379,In_1144);
and U5887 (N_5887,In_1611,In_2841);
and U5888 (N_5888,In_2581,In_2964);
and U5889 (N_5889,In_1273,In_2724);
or U5890 (N_5890,In_2025,In_2849);
nor U5891 (N_5891,In_433,In_2522);
nor U5892 (N_5892,In_2019,In_2374);
and U5893 (N_5893,In_1172,In_802);
or U5894 (N_5894,In_718,In_1272);
or U5895 (N_5895,In_496,In_2970);
or U5896 (N_5896,In_650,In_1713);
nor U5897 (N_5897,In_1949,In_1109);
nor U5898 (N_5898,In_445,In_240);
or U5899 (N_5899,In_2050,In_981);
nor U5900 (N_5900,In_264,In_1764);
or U5901 (N_5901,In_1637,In_1901);
and U5902 (N_5902,In_1778,In_1922);
nand U5903 (N_5903,In_508,In_2887);
and U5904 (N_5904,In_834,In_2738);
or U5905 (N_5905,In_1988,In_2525);
nand U5906 (N_5906,In_2765,In_710);
or U5907 (N_5907,In_883,In_2985);
and U5908 (N_5908,In_1371,In_66);
or U5909 (N_5909,In_373,In_1472);
and U5910 (N_5910,In_654,In_1889);
nor U5911 (N_5911,In_2981,In_1322);
nor U5912 (N_5912,In_1341,In_718);
nand U5913 (N_5913,In_46,In_2783);
nand U5914 (N_5914,In_2785,In_593);
nor U5915 (N_5915,In_2614,In_2016);
and U5916 (N_5916,In_1600,In_295);
nor U5917 (N_5917,In_625,In_2807);
nand U5918 (N_5918,In_916,In_2890);
or U5919 (N_5919,In_1175,In_748);
nor U5920 (N_5920,In_1548,In_2645);
nand U5921 (N_5921,In_2724,In_187);
nor U5922 (N_5922,In_2964,In_106);
or U5923 (N_5923,In_556,In_2410);
nand U5924 (N_5924,In_2203,In_1023);
nor U5925 (N_5925,In_945,In_245);
nand U5926 (N_5926,In_2648,In_101);
or U5927 (N_5927,In_779,In_2533);
nor U5928 (N_5928,In_519,In_2685);
nor U5929 (N_5929,In_1405,In_2822);
and U5930 (N_5930,In_525,In_918);
nand U5931 (N_5931,In_270,In_2645);
nand U5932 (N_5932,In_362,In_1591);
nand U5933 (N_5933,In_1060,In_1726);
and U5934 (N_5934,In_2820,In_1342);
nand U5935 (N_5935,In_2498,In_658);
and U5936 (N_5936,In_880,In_1873);
and U5937 (N_5937,In_1248,In_2298);
nor U5938 (N_5938,In_1047,In_1838);
nor U5939 (N_5939,In_2575,In_2711);
and U5940 (N_5940,In_1834,In_2907);
and U5941 (N_5941,In_682,In_884);
or U5942 (N_5942,In_435,In_2341);
and U5943 (N_5943,In_1124,In_1099);
nor U5944 (N_5944,In_2725,In_2734);
or U5945 (N_5945,In_1781,In_41);
nand U5946 (N_5946,In_2428,In_983);
and U5947 (N_5947,In_833,In_2242);
nor U5948 (N_5948,In_1987,In_615);
nand U5949 (N_5949,In_2363,In_1716);
nor U5950 (N_5950,In_1338,In_341);
or U5951 (N_5951,In_894,In_412);
and U5952 (N_5952,In_1399,In_1198);
nand U5953 (N_5953,In_638,In_1289);
or U5954 (N_5954,In_1192,In_1312);
nand U5955 (N_5955,In_1376,In_2809);
nand U5956 (N_5956,In_175,In_1970);
or U5957 (N_5957,In_1361,In_261);
and U5958 (N_5958,In_2927,In_613);
or U5959 (N_5959,In_624,In_1964);
and U5960 (N_5960,In_2936,In_2428);
nor U5961 (N_5961,In_2202,In_2504);
nand U5962 (N_5962,In_469,In_1524);
nor U5963 (N_5963,In_942,In_2712);
and U5964 (N_5964,In_970,In_1220);
and U5965 (N_5965,In_953,In_72);
or U5966 (N_5966,In_2708,In_2603);
nand U5967 (N_5967,In_446,In_724);
and U5968 (N_5968,In_2524,In_2015);
and U5969 (N_5969,In_1746,In_2597);
nand U5970 (N_5970,In_1327,In_2695);
nand U5971 (N_5971,In_866,In_11);
nand U5972 (N_5972,In_1955,In_1240);
or U5973 (N_5973,In_2369,In_790);
or U5974 (N_5974,In_1087,In_1645);
or U5975 (N_5975,In_2739,In_1578);
or U5976 (N_5976,In_566,In_1890);
and U5977 (N_5977,In_1088,In_216);
nor U5978 (N_5978,In_2250,In_850);
nor U5979 (N_5979,In_125,In_2702);
nand U5980 (N_5980,In_1146,In_2944);
nor U5981 (N_5981,In_2693,In_678);
nor U5982 (N_5982,In_1007,In_1293);
and U5983 (N_5983,In_1332,In_1709);
nor U5984 (N_5984,In_1781,In_875);
or U5985 (N_5985,In_1691,In_2198);
and U5986 (N_5986,In_84,In_2802);
and U5987 (N_5987,In_2005,In_1102);
nand U5988 (N_5988,In_1293,In_1265);
or U5989 (N_5989,In_78,In_1956);
nand U5990 (N_5990,In_2826,In_1903);
nor U5991 (N_5991,In_795,In_2738);
or U5992 (N_5992,In_2530,In_1285);
nor U5993 (N_5993,In_2274,In_2599);
or U5994 (N_5994,In_397,In_1293);
and U5995 (N_5995,In_1400,In_2953);
and U5996 (N_5996,In_2921,In_159);
or U5997 (N_5997,In_2877,In_1304);
and U5998 (N_5998,In_1521,In_2408);
or U5999 (N_5999,In_2391,In_2339);
or U6000 (N_6000,In_2617,In_224);
nor U6001 (N_6001,In_929,In_2408);
and U6002 (N_6002,In_866,In_529);
and U6003 (N_6003,In_1627,In_1377);
and U6004 (N_6004,In_1992,In_699);
nand U6005 (N_6005,In_1953,In_1425);
nand U6006 (N_6006,In_803,In_1391);
nand U6007 (N_6007,In_970,In_1830);
nor U6008 (N_6008,In_1260,In_2054);
nand U6009 (N_6009,In_468,In_2395);
nor U6010 (N_6010,In_2731,In_158);
and U6011 (N_6011,In_2421,In_2996);
and U6012 (N_6012,In_75,In_1552);
nor U6013 (N_6013,In_662,In_1679);
nor U6014 (N_6014,In_2273,In_750);
nand U6015 (N_6015,In_2779,In_658);
nand U6016 (N_6016,In_2292,In_1241);
or U6017 (N_6017,In_301,In_173);
and U6018 (N_6018,In_1884,In_1779);
or U6019 (N_6019,In_564,In_2996);
and U6020 (N_6020,In_1161,In_938);
or U6021 (N_6021,In_2645,In_2282);
and U6022 (N_6022,In_1414,In_2537);
or U6023 (N_6023,In_2720,In_1046);
and U6024 (N_6024,In_904,In_1504);
nor U6025 (N_6025,In_1788,In_2434);
nand U6026 (N_6026,In_773,In_569);
and U6027 (N_6027,In_692,In_44);
or U6028 (N_6028,In_2078,In_774);
nand U6029 (N_6029,In_1875,In_2136);
or U6030 (N_6030,In_1913,In_2791);
and U6031 (N_6031,In_1815,In_1451);
nor U6032 (N_6032,In_1073,In_2791);
nand U6033 (N_6033,In_978,In_1471);
nor U6034 (N_6034,In_2284,In_2159);
or U6035 (N_6035,In_1366,In_485);
nor U6036 (N_6036,In_2414,In_2255);
or U6037 (N_6037,In_529,In_464);
or U6038 (N_6038,In_2413,In_409);
and U6039 (N_6039,In_10,In_999);
nor U6040 (N_6040,In_922,In_285);
and U6041 (N_6041,In_684,In_2200);
nand U6042 (N_6042,In_2864,In_1008);
nor U6043 (N_6043,In_1395,In_771);
or U6044 (N_6044,In_1473,In_1372);
nor U6045 (N_6045,In_2149,In_791);
nor U6046 (N_6046,In_2624,In_2768);
or U6047 (N_6047,In_2233,In_2795);
or U6048 (N_6048,In_911,In_754);
or U6049 (N_6049,In_1876,In_490);
nand U6050 (N_6050,In_2593,In_1605);
or U6051 (N_6051,In_71,In_1725);
nand U6052 (N_6052,In_2034,In_780);
and U6053 (N_6053,In_717,In_1271);
nand U6054 (N_6054,In_2823,In_1463);
and U6055 (N_6055,In_2843,In_664);
or U6056 (N_6056,In_1795,In_2694);
and U6057 (N_6057,In_2529,In_2278);
or U6058 (N_6058,In_1156,In_2030);
nor U6059 (N_6059,In_1021,In_1601);
and U6060 (N_6060,In_8,In_916);
and U6061 (N_6061,In_356,In_674);
nand U6062 (N_6062,In_924,In_1345);
nor U6063 (N_6063,In_2042,In_1735);
or U6064 (N_6064,In_818,In_788);
nand U6065 (N_6065,In_1800,In_1157);
nand U6066 (N_6066,In_1709,In_2314);
nand U6067 (N_6067,In_2725,In_2814);
or U6068 (N_6068,In_2384,In_2925);
and U6069 (N_6069,In_536,In_1132);
nand U6070 (N_6070,In_809,In_465);
nor U6071 (N_6071,In_2252,In_1195);
nor U6072 (N_6072,In_2356,In_2532);
nor U6073 (N_6073,In_415,In_18);
nand U6074 (N_6074,In_1904,In_2229);
nor U6075 (N_6075,In_1418,In_881);
or U6076 (N_6076,In_1343,In_883);
and U6077 (N_6077,In_2279,In_2142);
or U6078 (N_6078,In_546,In_395);
nor U6079 (N_6079,In_667,In_1786);
nand U6080 (N_6080,In_2452,In_111);
nand U6081 (N_6081,In_1087,In_2104);
or U6082 (N_6082,In_2027,In_448);
and U6083 (N_6083,In_1314,In_806);
or U6084 (N_6084,In_2091,In_1501);
nand U6085 (N_6085,In_248,In_2491);
nand U6086 (N_6086,In_1141,In_2269);
and U6087 (N_6087,In_2612,In_129);
or U6088 (N_6088,In_1995,In_1055);
nor U6089 (N_6089,In_2173,In_2566);
nor U6090 (N_6090,In_447,In_2468);
nor U6091 (N_6091,In_2077,In_561);
and U6092 (N_6092,In_590,In_1881);
nor U6093 (N_6093,In_25,In_163);
nand U6094 (N_6094,In_2010,In_227);
nor U6095 (N_6095,In_1384,In_779);
or U6096 (N_6096,In_2440,In_821);
nand U6097 (N_6097,In_588,In_2496);
and U6098 (N_6098,In_2938,In_2942);
nor U6099 (N_6099,In_1373,In_1746);
nor U6100 (N_6100,In_1565,In_2556);
nand U6101 (N_6101,In_2003,In_2627);
or U6102 (N_6102,In_1841,In_1737);
or U6103 (N_6103,In_1490,In_277);
nand U6104 (N_6104,In_859,In_1824);
and U6105 (N_6105,In_737,In_1913);
or U6106 (N_6106,In_1862,In_2920);
nor U6107 (N_6107,In_894,In_2739);
nor U6108 (N_6108,In_1423,In_1918);
nand U6109 (N_6109,In_606,In_2136);
or U6110 (N_6110,In_1767,In_2947);
and U6111 (N_6111,In_846,In_789);
and U6112 (N_6112,In_2067,In_891);
and U6113 (N_6113,In_258,In_1193);
or U6114 (N_6114,In_2242,In_327);
or U6115 (N_6115,In_1608,In_1646);
or U6116 (N_6116,In_1419,In_2781);
nor U6117 (N_6117,In_771,In_2331);
and U6118 (N_6118,In_2282,In_2775);
or U6119 (N_6119,In_2052,In_794);
nor U6120 (N_6120,In_1666,In_896);
nand U6121 (N_6121,In_2145,In_674);
nand U6122 (N_6122,In_2005,In_819);
and U6123 (N_6123,In_1174,In_558);
nand U6124 (N_6124,In_273,In_821);
nor U6125 (N_6125,In_1131,In_2653);
nand U6126 (N_6126,In_2856,In_1102);
nor U6127 (N_6127,In_1571,In_717);
and U6128 (N_6128,In_1144,In_2801);
or U6129 (N_6129,In_750,In_1013);
nor U6130 (N_6130,In_338,In_2762);
nor U6131 (N_6131,In_227,In_2380);
nor U6132 (N_6132,In_171,In_2788);
nand U6133 (N_6133,In_1936,In_193);
or U6134 (N_6134,In_2111,In_500);
or U6135 (N_6135,In_1394,In_1117);
nand U6136 (N_6136,In_1952,In_226);
nand U6137 (N_6137,In_2702,In_2698);
and U6138 (N_6138,In_2190,In_1862);
or U6139 (N_6139,In_2726,In_1699);
and U6140 (N_6140,In_1365,In_2600);
or U6141 (N_6141,In_570,In_860);
nand U6142 (N_6142,In_2188,In_2308);
nand U6143 (N_6143,In_856,In_224);
and U6144 (N_6144,In_2726,In_1121);
nand U6145 (N_6145,In_1659,In_1346);
nor U6146 (N_6146,In_2306,In_849);
or U6147 (N_6147,In_571,In_2358);
or U6148 (N_6148,In_1865,In_1741);
nor U6149 (N_6149,In_547,In_279);
and U6150 (N_6150,In_1389,In_668);
and U6151 (N_6151,In_2000,In_1601);
and U6152 (N_6152,In_595,In_893);
nor U6153 (N_6153,In_1901,In_2924);
or U6154 (N_6154,In_1499,In_2298);
and U6155 (N_6155,In_2186,In_1997);
nand U6156 (N_6156,In_1942,In_1644);
and U6157 (N_6157,In_2118,In_2575);
or U6158 (N_6158,In_1858,In_719);
nor U6159 (N_6159,In_1408,In_628);
nand U6160 (N_6160,In_1503,In_1460);
nand U6161 (N_6161,In_989,In_940);
or U6162 (N_6162,In_2604,In_2034);
nand U6163 (N_6163,In_2135,In_350);
and U6164 (N_6164,In_2135,In_1731);
nand U6165 (N_6165,In_1199,In_2977);
and U6166 (N_6166,In_1583,In_422);
nor U6167 (N_6167,In_2644,In_1951);
nand U6168 (N_6168,In_672,In_2900);
or U6169 (N_6169,In_1282,In_2204);
nor U6170 (N_6170,In_671,In_1297);
nand U6171 (N_6171,In_2980,In_2936);
and U6172 (N_6172,In_2016,In_2059);
and U6173 (N_6173,In_400,In_302);
and U6174 (N_6174,In_1706,In_229);
nor U6175 (N_6175,In_157,In_1194);
and U6176 (N_6176,In_146,In_1342);
nand U6177 (N_6177,In_2352,In_1852);
or U6178 (N_6178,In_2972,In_1615);
nand U6179 (N_6179,In_2665,In_1340);
nand U6180 (N_6180,In_2587,In_1292);
nor U6181 (N_6181,In_621,In_1371);
nor U6182 (N_6182,In_644,In_2262);
and U6183 (N_6183,In_2272,In_2770);
or U6184 (N_6184,In_1999,In_2145);
or U6185 (N_6185,In_1388,In_1750);
nor U6186 (N_6186,In_808,In_2922);
and U6187 (N_6187,In_1410,In_205);
or U6188 (N_6188,In_766,In_2166);
nor U6189 (N_6189,In_1449,In_1101);
or U6190 (N_6190,In_139,In_220);
nand U6191 (N_6191,In_267,In_2367);
or U6192 (N_6192,In_2651,In_1754);
nor U6193 (N_6193,In_378,In_1139);
nand U6194 (N_6194,In_1431,In_2849);
nor U6195 (N_6195,In_2346,In_1220);
or U6196 (N_6196,In_2596,In_2825);
nand U6197 (N_6197,In_421,In_2795);
and U6198 (N_6198,In_446,In_483);
or U6199 (N_6199,In_2945,In_368);
and U6200 (N_6200,In_933,In_152);
nor U6201 (N_6201,In_567,In_1183);
or U6202 (N_6202,In_2361,In_216);
nand U6203 (N_6203,In_2614,In_1067);
and U6204 (N_6204,In_1194,In_242);
and U6205 (N_6205,In_1596,In_1004);
nand U6206 (N_6206,In_492,In_979);
nand U6207 (N_6207,In_1148,In_1471);
or U6208 (N_6208,In_2983,In_1589);
nand U6209 (N_6209,In_577,In_1275);
nand U6210 (N_6210,In_2017,In_2273);
and U6211 (N_6211,In_2583,In_1872);
or U6212 (N_6212,In_463,In_1921);
and U6213 (N_6213,In_1238,In_1018);
nor U6214 (N_6214,In_1043,In_2818);
nor U6215 (N_6215,In_207,In_1015);
nand U6216 (N_6216,In_793,In_531);
and U6217 (N_6217,In_2685,In_1191);
or U6218 (N_6218,In_252,In_1382);
nor U6219 (N_6219,In_1370,In_579);
nor U6220 (N_6220,In_1142,In_329);
nand U6221 (N_6221,In_1781,In_1699);
or U6222 (N_6222,In_1589,In_194);
nor U6223 (N_6223,In_1504,In_2563);
or U6224 (N_6224,In_437,In_1905);
and U6225 (N_6225,In_1832,In_2111);
and U6226 (N_6226,In_2945,In_902);
nand U6227 (N_6227,In_2408,In_2087);
and U6228 (N_6228,In_1041,In_2224);
or U6229 (N_6229,In_1032,In_1478);
and U6230 (N_6230,In_1444,In_657);
nand U6231 (N_6231,In_362,In_1026);
nor U6232 (N_6232,In_771,In_524);
nand U6233 (N_6233,In_1245,In_1791);
nand U6234 (N_6234,In_86,In_894);
or U6235 (N_6235,In_1392,In_1403);
nor U6236 (N_6236,In_214,In_319);
xor U6237 (N_6237,In_2936,In_728);
or U6238 (N_6238,In_196,In_2207);
or U6239 (N_6239,In_2175,In_1158);
nor U6240 (N_6240,In_1044,In_1500);
or U6241 (N_6241,In_118,In_2140);
nand U6242 (N_6242,In_1584,In_1211);
nand U6243 (N_6243,In_740,In_90);
nand U6244 (N_6244,In_2639,In_2311);
nor U6245 (N_6245,In_8,In_2195);
and U6246 (N_6246,In_2149,In_2948);
nand U6247 (N_6247,In_2387,In_1018);
nor U6248 (N_6248,In_54,In_896);
nor U6249 (N_6249,In_574,In_956);
nor U6250 (N_6250,In_699,In_582);
nand U6251 (N_6251,In_564,In_2585);
or U6252 (N_6252,In_2921,In_2439);
and U6253 (N_6253,In_2811,In_1215);
nor U6254 (N_6254,In_840,In_1963);
and U6255 (N_6255,In_2990,In_1186);
or U6256 (N_6256,In_1776,In_321);
or U6257 (N_6257,In_1659,In_32);
and U6258 (N_6258,In_1826,In_1045);
nand U6259 (N_6259,In_246,In_1921);
nor U6260 (N_6260,In_288,In_2168);
and U6261 (N_6261,In_809,In_2622);
and U6262 (N_6262,In_194,In_2784);
or U6263 (N_6263,In_1047,In_545);
and U6264 (N_6264,In_1625,In_1847);
and U6265 (N_6265,In_2262,In_254);
nor U6266 (N_6266,In_235,In_1727);
or U6267 (N_6267,In_2853,In_2860);
and U6268 (N_6268,In_1902,In_1467);
or U6269 (N_6269,In_799,In_184);
or U6270 (N_6270,In_719,In_1970);
and U6271 (N_6271,In_550,In_635);
and U6272 (N_6272,In_1235,In_678);
and U6273 (N_6273,In_1589,In_2389);
and U6274 (N_6274,In_2275,In_171);
or U6275 (N_6275,In_2020,In_1618);
and U6276 (N_6276,In_1123,In_1731);
nor U6277 (N_6277,In_373,In_2623);
nand U6278 (N_6278,In_1116,In_2163);
or U6279 (N_6279,In_1754,In_2698);
or U6280 (N_6280,In_895,In_2075);
xor U6281 (N_6281,In_1799,In_1930);
or U6282 (N_6282,In_186,In_14);
nand U6283 (N_6283,In_1640,In_2995);
or U6284 (N_6284,In_377,In_932);
nand U6285 (N_6285,In_331,In_2194);
and U6286 (N_6286,In_2835,In_454);
nor U6287 (N_6287,In_1018,In_2929);
nor U6288 (N_6288,In_750,In_2048);
nor U6289 (N_6289,In_1542,In_2183);
or U6290 (N_6290,In_2825,In_2069);
and U6291 (N_6291,In_2757,In_813);
and U6292 (N_6292,In_2616,In_2280);
xor U6293 (N_6293,In_2062,In_1623);
or U6294 (N_6294,In_2310,In_2286);
and U6295 (N_6295,In_1079,In_2822);
nand U6296 (N_6296,In_1577,In_175);
or U6297 (N_6297,In_901,In_32);
nor U6298 (N_6298,In_2490,In_2625);
and U6299 (N_6299,In_88,In_1212);
and U6300 (N_6300,In_786,In_846);
or U6301 (N_6301,In_1668,In_2287);
nor U6302 (N_6302,In_1131,In_830);
nor U6303 (N_6303,In_1218,In_1846);
or U6304 (N_6304,In_2476,In_1273);
nor U6305 (N_6305,In_1279,In_1608);
nor U6306 (N_6306,In_904,In_3);
nand U6307 (N_6307,In_2320,In_2571);
or U6308 (N_6308,In_2729,In_2084);
and U6309 (N_6309,In_2014,In_2951);
or U6310 (N_6310,In_2862,In_1418);
nand U6311 (N_6311,In_2165,In_1626);
nand U6312 (N_6312,In_2126,In_1299);
nand U6313 (N_6313,In_1442,In_1754);
or U6314 (N_6314,In_1116,In_2024);
and U6315 (N_6315,In_1873,In_38);
nand U6316 (N_6316,In_2945,In_658);
and U6317 (N_6317,In_1554,In_1204);
or U6318 (N_6318,In_2881,In_703);
nand U6319 (N_6319,In_1544,In_2852);
and U6320 (N_6320,In_2313,In_2996);
nand U6321 (N_6321,In_470,In_677);
nor U6322 (N_6322,In_1351,In_1871);
nand U6323 (N_6323,In_2442,In_2104);
nand U6324 (N_6324,In_1744,In_2452);
nor U6325 (N_6325,In_1225,In_1345);
and U6326 (N_6326,In_2063,In_2934);
nor U6327 (N_6327,In_2962,In_2668);
and U6328 (N_6328,In_1530,In_1692);
or U6329 (N_6329,In_1530,In_234);
and U6330 (N_6330,In_702,In_1174);
and U6331 (N_6331,In_1119,In_1490);
nand U6332 (N_6332,In_1283,In_1500);
or U6333 (N_6333,In_1574,In_1329);
or U6334 (N_6334,In_1832,In_633);
nand U6335 (N_6335,In_1353,In_896);
nor U6336 (N_6336,In_1779,In_1806);
nand U6337 (N_6337,In_2153,In_138);
nor U6338 (N_6338,In_1890,In_2117);
or U6339 (N_6339,In_35,In_1428);
nand U6340 (N_6340,In_425,In_2375);
nor U6341 (N_6341,In_2392,In_201);
nor U6342 (N_6342,In_983,In_2348);
nand U6343 (N_6343,In_2815,In_1517);
nor U6344 (N_6344,In_2156,In_446);
or U6345 (N_6345,In_492,In_2463);
nand U6346 (N_6346,In_1774,In_1892);
nor U6347 (N_6347,In_482,In_1320);
nor U6348 (N_6348,In_1901,In_1921);
or U6349 (N_6349,In_311,In_828);
and U6350 (N_6350,In_1320,In_2770);
and U6351 (N_6351,In_1748,In_1182);
nand U6352 (N_6352,In_2676,In_1706);
or U6353 (N_6353,In_424,In_838);
nand U6354 (N_6354,In_720,In_2029);
nand U6355 (N_6355,In_2329,In_2917);
nand U6356 (N_6356,In_573,In_2777);
and U6357 (N_6357,In_468,In_301);
nor U6358 (N_6358,In_1846,In_2005);
or U6359 (N_6359,In_1127,In_369);
or U6360 (N_6360,In_2930,In_165);
or U6361 (N_6361,In_2394,In_2279);
and U6362 (N_6362,In_329,In_457);
or U6363 (N_6363,In_1475,In_639);
or U6364 (N_6364,In_2384,In_620);
or U6365 (N_6365,In_2770,In_556);
nand U6366 (N_6366,In_554,In_1638);
nor U6367 (N_6367,In_591,In_2626);
nand U6368 (N_6368,In_2489,In_775);
nand U6369 (N_6369,In_2287,In_258);
nor U6370 (N_6370,In_1328,In_1219);
and U6371 (N_6371,In_1095,In_1144);
and U6372 (N_6372,In_2831,In_195);
nor U6373 (N_6373,In_2479,In_1225);
xor U6374 (N_6374,In_2259,In_438);
and U6375 (N_6375,In_2353,In_2354);
nand U6376 (N_6376,In_1404,In_2317);
and U6377 (N_6377,In_2777,In_2351);
nand U6378 (N_6378,In_551,In_1277);
and U6379 (N_6379,In_345,In_2450);
nor U6380 (N_6380,In_2141,In_1066);
nor U6381 (N_6381,In_1918,In_2131);
nor U6382 (N_6382,In_1519,In_1762);
and U6383 (N_6383,In_2749,In_2720);
nand U6384 (N_6384,In_538,In_2529);
xor U6385 (N_6385,In_1527,In_766);
or U6386 (N_6386,In_1853,In_2153);
nor U6387 (N_6387,In_2008,In_852);
or U6388 (N_6388,In_664,In_2581);
and U6389 (N_6389,In_1570,In_2520);
and U6390 (N_6390,In_1906,In_2134);
nor U6391 (N_6391,In_2589,In_2460);
nor U6392 (N_6392,In_2893,In_2811);
and U6393 (N_6393,In_1159,In_2326);
nand U6394 (N_6394,In_2557,In_2432);
nor U6395 (N_6395,In_2161,In_2643);
nand U6396 (N_6396,In_645,In_1151);
or U6397 (N_6397,In_2104,In_1403);
or U6398 (N_6398,In_792,In_1474);
and U6399 (N_6399,In_2509,In_1227);
nor U6400 (N_6400,In_501,In_896);
nor U6401 (N_6401,In_1153,In_1054);
or U6402 (N_6402,In_764,In_2928);
and U6403 (N_6403,In_1391,In_2295);
nor U6404 (N_6404,In_503,In_378);
nand U6405 (N_6405,In_2157,In_2279);
nand U6406 (N_6406,In_736,In_250);
and U6407 (N_6407,In_183,In_2804);
or U6408 (N_6408,In_2879,In_328);
and U6409 (N_6409,In_383,In_184);
or U6410 (N_6410,In_1277,In_276);
nand U6411 (N_6411,In_417,In_325);
nand U6412 (N_6412,In_1111,In_603);
or U6413 (N_6413,In_1346,In_2264);
nand U6414 (N_6414,In_2342,In_2247);
and U6415 (N_6415,In_1224,In_617);
nand U6416 (N_6416,In_2045,In_2137);
and U6417 (N_6417,In_2970,In_1165);
and U6418 (N_6418,In_66,In_465);
and U6419 (N_6419,In_2911,In_932);
and U6420 (N_6420,In_2034,In_1846);
and U6421 (N_6421,In_569,In_1924);
nand U6422 (N_6422,In_1046,In_939);
or U6423 (N_6423,In_2106,In_1158);
and U6424 (N_6424,In_2978,In_80);
nand U6425 (N_6425,In_1860,In_1233);
or U6426 (N_6426,In_1334,In_544);
or U6427 (N_6427,In_2161,In_2955);
or U6428 (N_6428,In_1532,In_1768);
or U6429 (N_6429,In_2374,In_900);
nor U6430 (N_6430,In_522,In_1514);
nand U6431 (N_6431,In_2875,In_1647);
and U6432 (N_6432,In_998,In_2011);
or U6433 (N_6433,In_1074,In_1329);
nor U6434 (N_6434,In_2755,In_916);
or U6435 (N_6435,In_2461,In_1944);
nor U6436 (N_6436,In_1910,In_1548);
nand U6437 (N_6437,In_323,In_935);
nor U6438 (N_6438,In_2900,In_1055);
xnor U6439 (N_6439,In_1534,In_1054);
and U6440 (N_6440,In_144,In_811);
nor U6441 (N_6441,In_97,In_1966);
nand U6442 (N_6442,In_1789,In_266);
or U6443 (N_6443,In_1676,In_1608);
nand U6444 (N_6444,In_116,In_1658);
or U6445 (N_6445,In_1885,In_2009);
nor U6446 (N_6446,In_1287,In_383);
and U6447 (N_6447,In_508,In_1369);
nor U6448 (N_6448,In_1021,In_1101);
or U6449 (N_6449,In_1797,In_1004);
nand U6450 (N_6450,In_2261,In_322);
nor U6451 (N_6451,In_2668,In_576);
or U6452 (N_6452,In_2225,In_543);
and U6453 (N_6453,In_493,In_1945);
nand U6454 (N_6454,In_2134,In_809);
or U6455 (N_6455,In_2822,In_2705);
nor U6456 (N_6456,In_1129,In_1523);
nor U6457 (N_6457,In_2009,In_1152);
nor U6458 (N_6458,In_1857,In_2210);
or U6459 (N_6459,In_716,In_93);
or U6460 (N_6460,In_2646,In_2005);
nand U6461 (N_6461,In_2962,In_873);
or U6462 (N_6462,In_2451,In_2065);
or U6463 (N_6463,In_901,In_2694);
and U6464 (N_6464,In_2591,In_726);
and U6465 (N_6465,In_723,In_2253);
nor U6466 (N_6466,In_401,In_28);
and U6467 (N_6467,In_1502,In_2696);
nor U6468 (N_6468,In_767,In_2445);
nor U6469 (N_6469,In_342,In_1059);
nor U6470 (N_6470,In_220,In_217);
and U6471 (N_6471,In_1384,In_2907);
or U6472 (N_6472,In_1508,In_351);
nor U6473 (N_6473,In_794,In_1835);
and U6474 (N_6474,In_120,In_216);
and U6475 (N_6475,In_2914,In_128);
and U6476 (N_6476,In_1130,In_1301);
or U6477 (N_6477,In_2389,In_793);
and U6478 (N_6478,In_401,In_2309);
and U6479 (N_6479,In_2842,In_2519);
nand U6480 (N_6480,In_572,In_1274);
nand U6481 (N_6481,In_2958,In_921);
or U6482 (N_6482,In_2929,In_2149);
or U6483 (N_6483,In_342,In_79);
and U6484 (N_6484,In_1816,In_2863);
nand U6485 (N_6485,In_1252,In_538);
and U6486 (N_6486,In_123,In_1258);
nand U6487 (N_6487,In_715,In_491);
nor U6488 (N_6488,In_578,In_2368);
nand U6489 (N_6489,In_1,In_2);
or U6490 (N_6490,In_1519,In_2864);
nand U6491 (N_6491,In_521,In_608);
nand U6492 (N_6492,In_2911,In_2009);
nand U6493 (N_6493,In_155,In_352);
and U6494 (N_6494,In_1375,In_311);
nor U6495 (N_6495,In_2751,In_2813);
and U6496 (N_6496,In_289,In_39);
and U6497 (N_6497,In_1045,In_526);
or U6498 (N_6498,In_2839,In_2499);
nand U6499 (N_6499,In_2144,In_311);
nor U6500 (N_6500,In_1939,In_1853);
and U6501 (N_6501,In_2790,In_2737);
or U6502 (N_6502,In_2441,In_975);
and U6503 (N_6503,In_2663,In_1546);
or U6504 (N_6504,In_1275,In_90);
or U6505 (N_6505,In_2074,In_855);
or U6506 (N_6506,In_745,In_2223);
or U6507 (N_6507,In_458,In_2135);
nand U6508 (N_6508,In_1166,In_1898);
nand U6509 (N_6509,In_2112,In_1426);
nand U6510 (N_6510,In_3,In_217);
and U6511 (N_6511,In_1650,In_1824);
or U6512 (N_6512,In_463,In_45);
nor U6513 (N_6513,In_2192,In_2015);
nor U6514 (N_6514,In_337,In_659);
nor U6515 (N_6515,In_2312,In_948);
and U6516 (N_6516,In_940,In_2725);
and U6517 (N_6517,In_314,In_1710);
nand U6518 (N_6518,In_58,In_1209);
nor U6519 (N_6519,In_1020,In_1259);
nor U6520 (N_6520,In_1709,In_1204);
xnor U6521 (N_6521,In_1298,In_1943);
and U6522 (N_6522,In_2151,In_830);
or U6523 (N_6523,In_1038,In_169);
nand U6524 (N_6524,In_1142,In_1331);
and U6525 (N_6525,In_2723,In_2903);
nand U6526 (N_6526,In_1259,In_2026);
nand U6527 (N_6527,In_1389,In_404);
and U6528 (N_6528,In_1087,In_1910);
or U6529 (N_6529,In_608,In_536);
or U6530 (N_6530,In_1366,In_952);
xnor U6531 (N_6531,In_757,In_1853);
and U6532 (N_6532,In_761,In_1981);
and U6533 (N_6533,In_2487,In_243);
nand U6534 (N_6534,In_796,In_951);
nor U6535 (N_6535,In_2918,In_1879);
nand U6536 (N_6536,In_2519,In_888);
and U6537 (N_6537,In_2319,In_1403);
and U6538 (N_6538,In_2470,In_1635);
nand U6539 (N_6539,In_1458,In_2952);
nand U6540 (N_6540,In_2652,In_417);
nor U6541 (N_6541,In_583,In_833);
or U6542 (N_6542,In_2571,In_1594);
nand U6543 (N_6543,In_1476,In_34);
and U6544 (N_6544,In_1102,In_209);
nand U6545 (N_6545,In_1845,In_1512);
and U6546 (N_6546,In_2881,In_1578);
nor U6547 (N_6547,In_1554,In_2265);
or U6548 (N_6548,In_1066,In_2442);
nor U6549 (N_6549,In_1877,In_1480);
or U6550 (N_6550,In_251,In_943);
nor U6551 (N_6551,In_73,In_2755);
or U6552 (N_6552,In_1165,In_2872);
and U6553 (N_6553,In_1196,In_2387);
nand U6554 (N_6554,In_842,In_1982);
nand U6555 (N_6555,In_2766,In_2028);
and U6556 (N_6556,In_1479,In_1750);
nor U6557 (N_6557,In_699,In_333);
or U6558 (N_6558,In_1294,In_1057);
nand U6559 (N_6559,In_1220,In_2707);
or U6560 (N_6560,In_1936,In_1624);
or U6561 (N_6561,In_2967,In_1919);
and U6562 (N_6562,In_104,In_2070);
or U6563 (N_6563,In_1557,In_135);
or U6564 (N_6564,In_2875,In_2977);
and U6565 (N_6565,In_2282,In_1497);
nand U6566 (N_6566,In_757,In_1587);
nand U6567 (N_6567,In_2389,In_2081);
nand U6568 (N_6568,In_787,In_2936);
or U6569 (N_6569,In_2036,In_2972);
nor U6570 (N_6570,In_2697,In_245);
nand U6571 (N_6571,In_1340,In_2489);
and U6572 (N_6572,In_2635,In_1845);
or U6573 (N_6573,In_989,In_2552);
and U6574 (N_6574,In_2257,In_1633);
and U6575 (N_6575,In_467,In_2179);
xor U6576 (N_6576,In_2248,In_194);
nor U6577 (N_6577,In_171,In_882);
and U6578 (N_6578,In_846,In_670);
nand U6579 (N_6579,In_1201,In_967);
or U6580 (N_6580,In_1355,In_1366);
nor U6581 (N_6581,In_558,In_1929);
nand U6582 (N_6582,In_766,In_2990);
and U6583 (N_6583,In_1865,In_892);
and U6584 (N_6584,In_2017,In_1054);
nor U6585 (N_6585,In_33,In_2633);
nand U6586 (N_6586,In_2706,In_425);
nor U6587 (N_6587,In_24,In_793);
nor U6588 (N_6588,In_2607,In_2111);
nand U6589 (N_6589,In_2545,In_378);
or U6590 (N_6590,In_393,In_474);
nor U6591 (N_6591,In_1415,In_2315);
and U6592 (N_6592,In_1802,In_1973);
and U6593 (N_6593,In_2613,In_1944);
or U6594 (N_6594,In_2568,In_1060);
and U6595 (N_6595,In_2767,In_1949);
and U6596 (N_6596,In_2203,In_798);
nand U6597 (N_6597,In_2316,In_2377);
or U6598 (N_6598,In_74,In_1701);
or U6599 (N_6599,In_288,In_2142);
nor U6600 (N_6600,In_658,In_2442);
or U6601 (N_6601,In_2020,In_993);
nand U6602 (N_6602,In_662,In_2379);
or U6603 (N_6603,In_1304,In_1677);
nor U6604 (N_6604,In_118,In_1);
and U6605 (N_6605,In_1692,In_1846);
and U6606 (N_6606,In_2304,In_109);
nand U6607 (N_6607,In_678,In_2310);
or U6608 (N_6608,In_921,In_2467);
or U6609 (N_6609,In_2760,In_1458);
nand U6610 (N_6610,In_52,In_969);
and U6611 (N_6611,In_2451,In_2412);
nor U6612 (N_6612,In_305,In_739);
and U6613 (N_6613,In_2164,In_2927);
or U6614 (N_6614,In_2240,In_181);
nand U6615 (N_6615,In_103,In_587);
or U6616 (N_6616,In_430,In_1679);
nand U6617 (N_6617,In_1802,In_1681);
nand U6618 (N_6618,In_1373,In_83);
and U6619 (N_6619,In_2663,In_1595);
or U6620 (N_6620,In_2748,In_2464);
nand U6621 (N_6621,In_966,In_1667);
nor U6622 (N_6622,In_2671,In_1570);
and U6623 (N_6623,In_1944,In_1313);
and U6624 (N_6624,In_1238,In_962);
nand U6625 (N_6625,In_29,In_1501);
or U6626 (N_6626,In_1101,In_1942);
nor U6627 (N_6627,In_2809,In_2810);
or U6628 (N_6628,In_2865,In_2472);
or U6629 (N_6629,In_2504,In_619);
nor U6630 (N_6630,In_41,In_1862);
nand U6631 (N_6631,In_1471,In_1544);
and U6632 (N_6632,In_1300,In_1877);
and U6633 (N_6633,In_1593,In_2913);
nor U6634 (N_6634,In_2138,In_1293);
nand U6635 (N_6635,In_277,In_1245);
xnor U6636 (N_6636,In_1199,In_1807);
nor U6637 (N_6637,In_234,In_2869);
or U6638 (N_6638,In_2052,In_1065);
or U6639 (N_6639,In_2021,In_2041);
or U6640 (N_6640,In_2348,In_770);
and U6641 (N_6641,In_350,In_468);
nor U6642 (N_6642,In_761,In_1299);
nand U6643 (N_6643,In_2309,In_935);
and U6644 (N_6644,In_849,In_902);
and U6645 (N_6645,In_2656,In_2781);
nand U6646 (N_6646,In_1810,In_2677);
or U6647 (N_6647,In_2287,In_1316);
and U6648 (N_6648,In_1162,In_841);
nor U6649 (N_6649,In_2636,In_2378);
nand U6650 (N_6650,In_448,In_1599);
or U6651 (N_6651,In_2977,In_1484);
or U6652 (N_6652,In_721,In_1704);
nor U6653 (N_6653,In_859,In_1110);
nand U6654 (N_6654,In_1657,In_576);
and U6655 (N_6655,In_701,In_423);
nand U6656 (N_6656,In_2195,In_555);
or U6657 (N_6657,In_246,In_209);
xnor U6658 (N_6658,In_420,In_1129);
or U6659 (N_6659,In_774,In_1165);
nor U6660 (N_6660,In_2200,In_1493);
xor U6661 (N_6661,In_2035,In_501);
nor U6662 (N_6662,In_1379,In_2604);
and U6663 (N_6663,In_1168,In_2549);
nand U6664 (N_6664,In_2040,In_69);
and U6665 (N_6665,In_2892,In_2471);
nor U6666 (N_6666,In_2229,In_1085);
and U6667 (N_6667,In_37,In_2877);
nor U6668 (N_6668,In_1987,In_2663);
and U6669 (N_6669,In_2545,In_609);
nor U6670 (N_6670,In_146,In_1646);
nor U6671 (N_6671,In_936,In_132);
nand U6672 (N_6672,In_679,In_1093);
and U6673 (N_6673,In_1482,In_1829);
nand U6674 (N_6674,In_1809,In_152);
or U6675 (N_6675,In_1249,In_2966);
nand U6676 (N_6676,In_2255,In_2561);
nand U6677 (N_6677,In_1598,In_984);
or U6678 (N_6678,In_2218,In_1983);
nand U6679 (N_6679,In_893,In_939);
and U6680 (N_6680,In_310,In_2110);
or U6681 (N_6681,In_872,In_1253);
and U6682 (N_6682,In_2736,In_2014);
nor U6683 (N_6683,In_2471,In_787);
or U6684 (N_6684,In_623,In_2942);
and U6685 (N_6685,In_1104,In_2630);
nand U6686 (N_6686,In_2698,In_2879);
nor U6687 (N_6687,In_2315,In_2267);
nand U6688 (N_6688,In_757,In_2135);
nor U6689 (N_6689,In_478,In_2418);
nor U6690 (N_6690,In_1810,In_951);
nand U6691 (N_6691,In_1705,In_2178);
nor U6692 (N_6692,In_885,In_2140);
nor U6693 (N_6693,In_122,In_1339);
nand U6694 (N_6694,In_796,In_2595);
nor U6695 (N_6695,In_816,In_1034);
and U6696 (N_6696,In_798,In_534);
or U6697 (N_6697,In_590,In_1530);
and U6698 (N_6698,In_604,In_516);
nor U6699 (N_6699,In_2133,In_2034);
nor U6700 (N_6700,In_334,In_2974);
and U6701 (N_6701,In_2651,In_1943);
nor U6702 (N_6702,In_1620,In_79);
and U6703 (N_6703,In_2484,In_2868);
or U6704 (N_6704,In_2188,In_2399);
and U6705 (N_6705,In_2552,In_2504);
and U6706 (N_6706,In_2501,In_2877);
nand U6707 (N_6707,In_2139,In_1831);
nand U6708 (N_6708,In_1028,In_2459);
and U6709 (N_6709,In_889,In_2865);
nor U6710 (N_6710,In_1135,In_703);
nor U6711 (N_6711,In_539,In_61);
or U6712 (N_6712,In_1074,In_1749);
nand U6713 (N_6713,In_842,In_812);
nand U6714 (N_6714,In_255,In_270);
and U6715 (N_6715,In_2422,In_837);
or U6716 (N_6716,In_1446,In_709);
nand U6717 (N_6717,In_2773,In_149);
nand U6718 (N_6718,In_1081,In_1913);
or U6719 (N_6719,In_2402,In_2673);
nand U6720 (N_6720,In_1186,In_2822);
or U6721 (N_6721,In_2118,In_756);
and U6722 (N_6722,In_1464,In_2057);
nor U6723 (N_6723,In_1677,In_2485);
nand U6724 (N_6724,In_640,In_1636);
and U6725 (N_6725,In_2268,In_2525);
nand U6726 (N_6726,In_437,In_2495);
or U6727 (N_6727,In_1674,In_159);
nor U6728 (N_6728,In_1735,In_2764);
and U6729 (N_6729,In_2968,In_2853);
or U6730 (N_6730,In_68,In_2679);
and U6731 (N_6731,In_2471,In_1827);
and U6732 (N_6732,In_2831,In_780);
nor U6733 (N_6733,In_253,In_2321);
or U6734 (N_6734,In_1128,In_1576);
and U6735 (N_6735,In_144,In_1553);
and U6736 (N_6736,In_48,In_305);
and U6737 (N_6737,In_2759,In_62);
and U6738 (N_6738,In_909,In_1988);
nand U6739 (N_6739,In_1216,In_1564);
or U6740 (N_6740,In_1893,In_108);
or U6741 (N_6741,In_1718,In_1481);
and U6742 (N_6742,In_1965,In_850);
and U6743 (N_6743,In_1539,In_1867);
or U6744 (N_6744,In_15,In_1199);
and U6745 (N_6745,In_702,In_1230);
nor U6746 (N_6746,In_1030,In_229);
or U6747 (N_6747,In_2850,In_580);
nor U6748 (N_6748,In_2466,In_486);
nand U6749 (N_6749,In_2478,In_1505);
nor U6750 (N_6750,In_200,In_155);
and U6751 (N_6751,In_2211,In_2941);
and U6752 (N_6752,In_2356,In_1719);
nor U6753 (N_6753,In_2697,In_2886);
nand U6754 (N_6754,In_880,In_906);
nor U6755 (N_6755,In_1508,In_623);
and U6756 (N_6756,In_1234,In_1935);
or U6757 (N_6757,In_2048,In_192);
nand U6758 (N_6758,In_2024,In_68);
xor U6759 (N_6759,In_59,In_168);
or U6760 (N_6760,In_2534,In_1615);
or U6761 (N_6761,In_526,In_2423);
nor U6762 (N_6762,In_2332,In_2702);
or U6763 (N_6763,In_175,In_1675);
and U6764 (N_6764,In_854,In_2717);
nor U6765 (N_6765,In_2692,In_1189);
nor U6766 (N_6766,In_962,In_470);
or U6767 (N_6767,In_1948,In_1518);
or U6768 (N_6768,In_1742,In_1169);
nor U6769 (N_6769,In_124,In_2633);
or U6770 (N_6770,In_587,In_1010);
nor U6771 (N_6771,In_2143,In_210);
or U6772 (N_6772,In_566,In_1130);
or U6773 (N_6773,In_789,In_1831);
and U6774 (N_6774,In_29,In_2579);
and U6775 (N_6775,In_1070,In_1906);
and U6776 (N_6776,In_1472,In_255);
or U6777 (N_6777,In_32,In_2323);
or U6778 (N_6778,In_543,In_940);
nand U6779 (N_6779,In_142,In_219);
and U6780 (N_6780,In_78,In_377);
or U6781 (N_6781,In_242,In_756);
nand U6782 (N_6782,In_35,In_821);
nor U6783 (N_6783,In_413,In_1373);
or U6784 (N_6784,In_544,In_1694);
and U6785 (N_6785,In_955,In_887);
nor U6786 (N_6786,In_1848,In_2247);
nand U6787 (N_6787,In_743,In_1340);
or U6788 (N_6788,In_1224,In_1079);
and U6789 (N_6789,In_704,In_2788);
nor U6790 (N_6790,In_2479,In_1732);
or U6791 (N_6791,In_720,In_256);
nand U6792 (N_6792,In_181,In_570);
nand U6793 (N_6793,In_1230,In_194);
nand U6794 (N_6794,In_1155,In_597);
nor U6795 (N_6795,In_1423,In_330);
and U6796 (N_6796,In_2589,In_1985);
nand U6797 (N_6797,In_2169,In_146);
and U6798 (N_6798,In_1569,In_2278);
nor U6799 (N_6799,In_1244,In_298);
and U6800 (N_6800,In_1823,In_1787);
nor U6801 (N_6801,In_353,In_1032);
or U6802 (N_6802,In_2899,In_1792);
nor U6803 (N_6803,In_2121,In_437);
or U6804 (N_6804,In_466,In_1773);
nand U6805 (N_6805,In_1817,In_2494);
nor U6806 (N_6806,In_529,In_820);
and U6807 (N_6807,In_67,In_155);
or U6808 (N_6808,In_2195,In_1046);
nor U6809 (N_6809,In_928,In_2801);
xnor U6810 (N_6810,In_2012,In_1713);
nand U6811 (N_6811,In_1245,In_1618);
and U6812 (N_6812,In_1477,In_135);
nand U6813 (N_6813,In_2994,In_2026);
or U6814 (N_6814,In_2560,In_1434);
nand U6815 (N_6815,In_1489,In_160);
and U6816 (N_6816,In_2045,In_2054);
and U6817 (N_6817,In_1055,In_872);
or U6818 (N_6818,In_922,In_2951);
nand U6819 (N_6819,In_501,In_1086);
nand U6820 (N_6820,In_681,In_2072);
or U6821 (N_6821,In_2892,In_1902);
or U6822 (N_6822,In_2075,In_2481);
nand U6823 (N_6823,In_1528,In_1934);
and U6824 (N_6824,In_504,In_262);
and U6825 (N_6825,In_157,In_896);
nand U6826 (N_6826,In_2463,In_1032);
or U6827 (N_6827,In_908,In_440);
nand U6828 (N_6828,In_1338,In_1363);
xnor U6829 (N_6829,In_2165,In_284);
nor U6830 (N_6830,In_2035,In_2856);
nand U6831 (N_6831,In_2297,In_1976);
nand U6832 (N_6832,In_527,In_2818);
and U6833 (N_6833,In_940,In_2526);
and U6834 (N_6834,In_1183,In_1484);
and U6835 (N_6835,In_185,In_1880);
nand U6836 (N_6836,In_2659,In_309);
and U6837 (N_6837,In_1859,In_659);
and U6838 (N_6838,In_1379,In_1958);
nand U6839 (N_6839,In_53,In_1154);
nor U6840 (N_6840,In_2692,In_2863);
or U6841 (N_6841,In_2744,In_2222);
or U6842 (N_6842,In_2771,In_2152);
nor U6843 (N_6843,In_70,In_2722);
nor U6844 (N_6844,In_1358,In_2699);
nor U6845 (N_6845,In_2058,In_360);
xor U6846 (N_6846,In_83,In_110);
nand U6847 (N_6847,In_2859,In_733);
nand U6848 (N_6848,In_275,In_1099);
nor U6849 (N_6849,In_2494,In_1475);
and U6850 (N_6850,In_2140,In_1145);
nor U6851 (N_6851,In_2166,In_2329);
or U6852 (N_6852,In_1450,In_360);
nand U6853 (N_6853,In_1085,In_2120);
or U6854 (N_6854,In_851,In_2898);
and U6855 (N_6855,In_1032,In_40);
or U6856 (N_6856,In_1089,In_863);
or U6857 (N_6857,In_311,In_743);
nor U6858 (N_6858,In_2497,In_482);
or U6859 (N_6859,In_2387,In_191);
nand U6860 (N_6860,In_2446,In_2174);
nand U6861 (N_6861,In_1326,In_949);
and U6862 (N_6862,In_371,In_362);
or U6863 (N_6863,In_1841,In_2252);
or U6864 (N_6864,In_1225,In_2797);
or U6865 (N_6865,In_2757,In_2511);
nand U6866 (N_6866,In_2419,In_2834);
nand U6867 (N_6867,In_1921,In_2453);
or U6868 (N_6868,In_2153,In_1106);
nor U6869 (N_6869,In_1157,In_866);
nor U6870 (N_6870,In_1532,In_730);
nor U6871 (N_6871,In_2076,In_1311);
and U6872 (N_6872,In_1574,In_1825);
nor U6873 (N_6873,In_218,In_1587);
and U6874 (N_6874,In_1377,In_2613);
or U6875 (N_6875,In_2098,In_2393);
and U6876 (N_6876,In_2444,In_486);
nor U6877 (N_6877,In_770,In_1613);
or U6878 (N_6878,In_1151,In_767);
nand U6879 (N_6879,In_2801,In_2026);
or U6880 (N_6880,In_619,In_745);
or U6881 (N_6881,In_2036,In_1527);
and U6882 (N_6882,In_1853,In_1615);
or U6883 (N_6883,In_2590,In_1880);
nand U6884 (N_6884,In_1383,In_2235);
and U6885 (N_6885,In_1584,In_1279);
or U6886 (N_6886,In_2427,In_623);
and U6887 (N_6887,In_481,In_2445);
nor U6888 (N_6888,In_1294,In_2784);
or U6889 (N_6889,In_1427,In_2595);
or U6890 (N_6890,In_642,In_79);
nor U6891 (N_6891,In_2495,In_2402);
nor U6892 (N_6892,In_1830,In_1014);
or U6893 (N_6893,In_2505,In_2298);
or U6894 (N_6894,In_517,In_120);
or U6895 (N_6895,In_539,In_211);
nand U6896 (N_6896,In_1506,In_1088);
and U6897 (N_6897,In_1677,In_1410);
nand U6898 (N_6898,In_1592,In_273);
or U6899 (N_6899,In_1570,In_243);
or U6900 (N_6900,In_88,In_1320);
nor U6901 (N_6901,In_2024,In_148);
nor U6902 (N_6902,In_1118,In_2514);
or U6903 (N_6903,In_2928,In_2949);
nor U6904 (N_6904,In_1372,In_1733);
nor U6905 (N_6905,In_27,In_1914);
and U6906 (N_6906,In_1912,In_626);
nand U6907 (N_6907,In_823,In_2977);
nor U6908 (N_6908,In_2833,In_2521);
nor U6909 (N_6909,In_918,In_2242);
and U6910 (N_6910,In_735,In_221);
or U6911 (N_6911,In_2802,In_28);
and U6912 (N_6912,In_1010,In_1120);
or U6913 (N_6913,In_728,In_647);
and U6914 (N_6914,In_471,In_294);
nor U6915 (N_6915,In_1433,In_299);
nand U6916 (N_6916,In_1955,In_1247);
nor U6917 (N_6917,In_1932,In_109);
and U6918 (N_6918,In_2309,In_793);
xor U6919 (N_6919,In_1763,In_1070);
nor U6920 (N_6920,In_2314,In_150);
nand U6921 (N_6921,In_877,In_2418);
and U6922 (N_6922,In_2889,In_1563);
and U6923 (N_6923,In_2190,In_2730);
or U6924 (N_6924,In_2540,In_2331);
or U6925 (N_6925,In_1985,In_1995);
and U6926 (N_6926,In_932,In_315);
or U6927 (N_6927,In_2781,In_119);
or U6928 (N_6928,In_689,In_1285);
nand U6929 (N_6929,In_2748,In_2793);
nand U6930 (N_6930,In_1205,In_1974);
nor U6931 (N_6931,In_67,In_1561);
nor U6932 (N_6932,In_1756,In_699);
and U6933 (N_6933,In_1162,In_515);
or U6934 (N_6934,In_1638,In_184);
xor U6935 (N_6935,In_2227,In_271);
and U6936 (N_6936,In_342,In_1041);
nor U6937 (N_6937,In_1850,In_260);
nand U6938 (N_6938,In_693,In_471);
and U6939 (N_6939,In_2291,In_1472);
and U6940 (N_6940,In_1877,In_681);
nor U6941 (N_6941,In_2807,In_2060);
or U6942 (N_6942,In_2738,In_625);
or U6943 (N_6943,In_524,In_2831);
or U6944 (N_6944,In_1995,In_2734);
or U6945 (N_6945,In_1139,In_698);
and U6946 (N_6946,In_2017,In_204);
and U6947 (N_6947,In_1217,In_763);
or U6948 (N_6948,In_2650,In_2055);
nor U6949 (N_6949,In_1828,In_2197);
nor U6950 (N_6950,In_2019,In_2125);
nand U6951 (N_6951,In_1136,In_486);
nand U6952 (N_6952,In_2479,In_2284);
or U6953 (N_6953,In_301,In_236);
nand U6954 (N_6954,In_2252,In_1788);
nor U6955 (N_6955,In_1057,In_2142);
nor U6956 (N_6956,In_2579,In_687);
nand U6957 (N_6957,In_1072,In_283);
nand U6958 (N_6958,In_2845,In_2550);
nor U6959 (N_6959,In_1809,In_1018);
and U6960 (N_6960,In_908,In_206);
nor U6961 (N_6961,In_2731,In_1426);
nand U6962 (N_6962,In_1385,In_2377);
and U6963 (N_6963,In_563,In_1890);
nand U6964 (N_6964,In_1593,In_715);
nor U6965 (N_6965,In_2650,In_1787);
and U6966 (N_6966,In_136,In_2774);
nand U6967 (N_6967,In_2816,In_2153);
nor U6968 (N_6968,In_2231,In_2449);
or U6969 (N_6969,In_601,In_2749);
and U6970 (N_6970,In_1298,In_1813);
or U6971 (N_6971,In_891,In_855);
or U6972 (N_6972,In_2166,In_2081);
nand U6973 (N_6973,In_1926,In_1466);
nand U6974 (N_6974,In_1584,In_2625);
or U6975 (N_6975,In_787,In_124);
nor U6976 (N_6976,In_142,In_2077);
and U6977 (N_6977,In_2996,In_1512);
or U6978 (N_6978,In_2428,In_1498);
nor U6979 (N_6979,In_2854,In_849);
nor U6980 (N_6980,In_1794,In_370);
nor U6981 (N_6981,In_1294,In_783);
nand U6982 (N_6982,In_2783,In_2371);
xor U6983 (N_6983,In_285,In_2794);
and U6984 (N_6984,In_814,In_2167);
or U6985 (N_6985,In_1494,In_2117);
nand U6986 (N_6986,In_2757,In_1982);
nand U6987 (N_6987,In_1784,In_1002);
nor U6988 (N_6988,In_2296,In_808);
nor U6989 (N_6989,In_2911,In_1227);
nor U6990 (N_6990,In_2649,In_1376);
or U6991 (N_6991,In_2812,In_1365);
or U6992 (N_6992,In_722,In_210);
or U6993 (N_6993,In_583,In_130);
nand U6994 (N_6994,In_2438,In_1115);
nor U6995 (N_6995,In_368,In_501);
and U6996 (N_6996,In_467,In_360);
or U6997 (N_6997,In_646,In_7);
nor U6998 (N_6998,In_425,In_781);
nand U6999 (N_6999,In_1825,In_1248);
nor U7000 (N_7000,In_2567,In_484);
nor U7001 (N_7001,In_757,In_2950);
nand U7002 (N_7002,In_1338,In_1551);
and U7003 (N_7003,In_2208,In_354);
and U7004 (N_7004,In_324,In_891);
and U7005 (N_7005,In_1664,In_1022);
and U7006 (N_7006,In_1608,In_1271);
nor U7007 (N_7007,In_2672,In_921);
and U7008 (N_7008,In_1792,In_2580);
nor U7009 (N_7009,In_1735,In_2404);
nor U7010 (N_7010,In_2672,In_1857);
and U7011 (N_7011,In_1241,In_2965);
nor U7012 (N_7012,In_1467,In_587);
nor U7013 (N_7013,In_2462,In_1404);
or U7014 (N_7014,In_497,In_1851);
nand U7015 (N_7015,In_1941,In_1824);
or U7016 (N_7016,In_272,In_2297);
nor U7017 (N_7017,In_162,In_1580);
nand U7018 (N_7018,In_1065,In_2057);
and U7019 (N_7019,In_831,In_2736);
and U7020 (N_7020,In_2546,In_2719);
nand U7021 (N_7021,In_514,In_1258);
nor U7022 (N_7022,In_2557,In_1320);
nand U7023 (N_7023,In_214,In_682);
nand U7024 (N_7024,In_737,In_1041);
and U7025 (N_7025,In_1704,In_867);
nor U7026 (N_7026,In_678,In_1357);
and U7027 (N_7027,In_244,In_590);
and U7028 (N_7028,In_2311,In_672);
nand U7029 (N_7029,In_2222,In_1383);
nor U7030 (N_7030,In_1423,In_1218);
or U7031 (N_7031,In_970,In_1752);
and U7032 (N_7032,In_2390,In_2856);
nor U7033 (N_7033,In_246,In_2593);
nand U7034 (N_7034,In_2886,In_1885);
nor U7035 (N_7035,In_937,In_1419);
nor U7036 (N_7036,In_2388,In_1074);
nor U7037 (N_7037,In_834,In_2410);
and U7038 (N_7038,In_2100,In_1478);
nor U7039 (N_7039,In_122,In_793);
nor U7040 (N_7040,In_638,In_1092);
or U7041 (N_7041,In_2175,In_538);
or U7042 (N_7042,In_2948,In_699);
or U7043 (N_7043,In_2757,In_2278);
nand U7044 (N_7044,In_1421,In_649);
nor U7045 (N_7045,In_2630,In_2598);
or U7046 (N_7046,In_634,In_1780);
nand U7047 (N_7047,In_939,In_2412);
or U7048 (N_7048,In_275,In_1910);
and U7049 (N_7049,In_2459,In_1171);
nor U7050 (N_7050,In_2969,In_1346);
or U7051 (N_7051,In_2816,In_1998);
nor U7052 (N_7052,In_607,In_2145);
and U7053 (N_7053,In_1209,In_648);
nor U7054 (N_7054,In_630,In_1484);
or U7055 (N_7055,In_596,In_1830);
nor U7056 (N_7056,In_1918,In_554);
or U7057 (N_7057,In_271,In_2590);
or U7058 (N_7058,In_1685,In_1556);
nor U7059 (N_7059,In_1059,In_167);
and U7060 (N_7060,In_1331,In_466);
nor U7061 (N_7061,In_1852,In_1295);
or U7062 (N_7062,In_0,In_1471);
nor U7063 (N_7063,In_2711,In_108);
nor U7064 (N_7064,In_716,In_843);
and U7065 (N_7065,In_1003,In_2287);
or U7066 (N_7066,In_2678,In_1160);
nor U7067 (N_7067,In_2906,In_2979);
or U7068 (N_7068,In_2212,In_970);
or U7069 (N_7069,In_427,In_1452);
or U7070 (N_7070,In_848,In_2214);
or U7071 (N_7071,In_2208,In_301);
nand U7072 (N_7072,In_1469,In_1197);
nand U7073 (N_7073,In_2054,In_25);
or U7074 (N_7074,In_2972,In_1269);
or U7075 (N_7075,In_2439,In_1031);
nand U7076 (N_7076,In_1701,In_1152);
nor U7077 (N_7077,In_1476,In_2215);
and U7078 (N_7078,In_739,In_1843);
nor U7079 (N_7079,In_221,In_2945);
or U7080 (N_7080,In_2367,In_2025);
nand U7081 (N_7081,In_1234,In_1111);
nor U7082 (N_7082,In_837,In_391);
or U7083 (N_7083,In_2396,In_1123);
nand U7084 (N_7084,In_777,In_692);
and U7085 (N_7085,In_387,In_2674);
or U7086 (N_7086,In_1801,In_2210);
or U7087 (N_7087,In_2440,In_207);
nand U7088 (N_7088,In_796,In_918);
nand U7089 (N_7089,In_463,In_27);
or U7090 (N_7090,In_546,In_33);
nor U7091 (N_7091,In_28,In_2601);
and U7092 (N_7092,In_714,In_502);
nand U7093 (N_7093,In_1315,In_1030);
and U7094 (N_7094,In_825,In_2838);
nand U7095 (N_7095,In_1245,In_177);
and U7096 (N_7096,In_1632,In_2452);
nand U7097 (N_7097,In_2149,In_1709);
and U7098 (N_7098,In_66,In_428);
nor U7099 (N_7099,In_1440,In_1557);
and U7100 (N_7100,In_322,In_1800);
or U7101 (N_7101,In_1282,In_1244);
and U7102 (N_7102,In_94,In_1441);
and U7103 (N_7103,In_2702,In_2980);
and U7104 (N_7104,In_770,In_2968);
or U7105 (N_7105,In_2309,In_1617);
or U7106 (N_7106,In_2680,In_1536);
or U7107 (N_7107,In_1445,In_279);
nor U7108 (N_7108,In_2586,In_2703);
nor U7109 (N_7109,In_1300,In_2914);
or U7110 (N_7110,In_1607,In_2533);
nand U7111 (N_7111,In_2826,In_2125);
nor U7112 (N_7112,In_1719,In_302);
or U7113 (N_7113,In_1773,In_1032);
and U7114 (N_7114,In_2460,In_1462);
nor U7115 (N_7115,In_1599,In_97);
nand U7116 (N_7116,In_424,In_1419);
nor U7117 (N_7117,In_1493,In_2748);
or U7118 (N_7118,In_2167,In_1583);
nor U7119 (N_7119,In_859,In_479);
or U7120 (N_7120,In_2005,In_1015);
nand U7121 (N_7121,In_2455,In_2080);
and U7122 (N_7122,In_1871,In_2457);
nand U7123 (N_7123,In_524,In_2804);
xor U7124 (N_7124,In_2526,In_147);
nand U7125 (N_7125,In_893,In_771);
and U7126 (N_7126,In_448,In_2539);
nand U7127 (N_7127,In_519,In_22);
or U7128 (N_7128,In_2324,In_2269);
and U7129 (N_7129,In_1999,In_402);
nor U7130 (N_7130,In_2626,In_1867);
nor U7131 (N_7131,In_2199,In_1861);
nor U7132 (N_7132,In_697,In_1293);
nand U7133 (N_7133,In_292,In_1666);
and U7134 (N_7134,In_1746,In_69);
or U7135 (N_7135,In_1395,In_1746);
or U7136 (N_7136,In_2481,In_131);
nand U7137 (N_7137,In_1732,In_791);
nor U7138 (N_7138,In_1446,In_1587);
or U7139 (N_7139,In_2930,In_2373);
and U7140 (N_7140,In_2432,In_1359);
or U7141 (N_7141,In_1995,In_295);
nor U7142 (N_7142,In_2844,In_313);
or U7143 (N_7143,In_774,In_2103);
or U7144 (N_7144,In_2256,In_788);
and U7145 (N_7145,In_2733,In_1116);
or U7146 (N_7146,In_1314,In_1255);
xnor U7147 (N_7147,In_2562,In_969);
and U7148 (N_7148,In_1776,In_2872);
nor U7149 (N_7149,In_286,In_2202);
nand U7150 (N_7150,In_1014,In_2154);
nand U7151 (N_7151,In_1809,In_260);
and U7152 (N_7152,In_1378,In_1857);
nor U7153 (N_7153,In_2880,In_312);
xor U7154 (N_7154,In_35,In_1499);
nor U7155 (N_7155,In_2113,In_109);
or U7156 (N_7156,In_750,In_2667);
or U7157 (N_7157,In_720,In_83);
nand U7158 (N_7158,In_1300,In_818);
nand U7159 (N_7159,In_1304,In_1938);
and U7160 (N_7160,In_1407,In_1697);
nor U7161 (N_7161,In_1015,In_2152);
and U7162 (N_7162,In_1694,In_660);
and U7163 (N_7163,In_2365,In_2498);
nand U7164 (N_7164,In_910,In_2298);
nor U7165 (N_7165,In_1873,In_157);
or U7166 (N_7166,In_876,In_1628);
nor U7167 (N_7167,In_287,In_1377);
nor U7168 (N_7168,In_2590,In_873);
or U7169 (N_7169,In_139,In_2045);
or U7170 (N_7170,In_519,In_2230);
nor U7171 (N_7171,In_1174,In_2123);
nand U7172 (N_7172,In_2729,In_1248);
nand U7173 (N_7173,In_1665,In_751);
or U7174 (N_7174,In_539,In_658);
nor U7175 (N_7175,In_2269,In_877);
nand U7176 (N_7176,In_2514,In_2426);
and U7177 (N_7177,In_416,In_874);
or U7178 (N_7178,In_330,In_16);
nand U7179 (N_7179,In_2670,In_1268);
nand U7180 (N_7180,In_2119,In_1008);
nor U7181 (N_7181,In_1366,In_373);
and U7182 (N_7182,In_2606,In_2617);
or U7183 (N_7183,In_1485,In_2994);
or U7184 (N_7184,In_1187,In_1401);
or U7185 (N_7185,In_2082,In_1707);
or U7186 (N_7186,In_170,In_1547);
nand U7187 (N_7187,In_433,In_603);
nand U7188 (N_7188,In_146,In_1867);
nor U7189 (N_7189,In_1729,In_629);
and U7190 (N_7190,In_2451,In_2356);
or U7191 (N_7191,In_730,In_126);
nand U7192 (N_7192,In_2785,In_331);
and U7193 (N_7193,In_304,In_280);
and U7194 (N_7194,In_880,In_2541);
or U7195 (N_7195,In_2878,In_1031);
nand U7196 (N_7196,In_1003,In_2057);
xnor U7197 (N_7197,In_2033,In_30);
nor U7198 (N_7198,In_1362,In_2028);
and U7199 (N_7199,In_1103,In_1665);
or U7200 (N_7200,In_882,In_2308);
or U7201 (N_7201,In_2040,In_2136);
and U7202 (N_7202,In_1859,In_906);
and U7203 (N_7203,In_150,In_2795);
and U7204 (N_7204,In_748,In_392);
and U7205 (N_7205,In_213,In_1760);
nor U7206 (N_7206,In_2645,In_126);
nand U7207 (N_7207,In_1133,In_165);
nand U7208 (N_7208,In_843,In_2091);
nor U7209 (N_7209,In_2266,In_1230);
nand U7210 (N_7210,In_2571,In_1091);
nor U7211 (N_7211,In_797,In_2051);
nand U7212 (N_7212,In_252,In_2797);
nor U7213 (N_7213,In_2268,In_1883);
or U7214 (N_7214,In_1543,In_2359);
and U7215 (N_7215,In_662,In_2245);
and U7216 (N_7216,In_929,In_1362);
nand U7217 (N_7217,In_218,In_2870);
nor U7218 (N_7218,In_1590,In_2515);
and U7219 (N_7219,In_2630,In_1798);
and U7220 (N_7220,In_1249,In_2762);
or U7221 (N_7221,In_1462,In_2311);
and U7222 (N_7222,In_1827,In_1878);
and U7223 (N_7223,In_2771,In_2696);
nand U7224 (N_7224,In_858,In_333);
nand U7225 (N_7225,In_2105,In_129);
nand U7226 (N_7226,In_1347,In_849);
nor U7227 (N_7227,In_84,In_54);
nand U7228 (N_7228,In_1357,In_1437);
and U7229 (N_7229,In_1910,In_2529);
nor U7230 (N_7230,In_2689,In_1712);
nor U7231 (N_7231,In_2194,In_1352);
and U7232 (N_7232,In_60,In_2501);
and U7233 (N_7233,In_2708,In_1384);
or U7234 (N_7234,In_836,In_1446);
nor U7235 (N_7235,In_229,In_798);
and U7236 (N_7236,In_113,In_2641);
and U7237 (N_7237,In_521,In_1347);
or U7238 (N_7238,In_2518,In_1881);
and U7239 (N_7239,In_502,In_2494);
or U7240 (N_7240,In_1325,In_2940);
or U7241 (N_7241,In_339,In_1619);
nand U7242 (N_7242,In_1638,In_908);
nor U7243 (N_7243,In_2505,In_1974);
and U7244 (N_7244,In_614,In_734);
and U7245 (N_7245,In_171,In_2368);
nand U7246 (N_7246,In_159,In_379);
or U7247 (N_7247,In_1772,In_2725);
nor U7248 (N_7248,In_1259,In_2873);
nor U7249 (N_7249,In_677,In_198);
or U7250 (N_7250,In_1019,In_1720);
nand U7251 (N_7251,In_480,In_1831);
or U7252 (N_7252,In_320,In_1732);
or U7253 (N_7253,In_467,In_2445);
or U7254 (N_7254,In_386,In_1767);
and U7255 (N_7255,In_1167,In_82);
and U7256 (N_7256,In_1553,In_1562);
nor U7257 (N_7257,In_1068,In_1452);
nor U7258 (N_7258,In_1429,In_2924);
nor U7259 (N_7259,In_532,In_2730);
nor U7260 (N_7260,In_1223,In_2830);
or U7261 (N_7261,In_215,In_2185);
and U7262 (N_7262,In_396,In_1804);
or U7263 (N_7263,In_1044,In_2444);
nand U7264 (N_7264,In_2197,In_2453);
or U7265 (N_7265,In_430,In_712);
or U7266 (N_7266,In_1969,In_627);
and U7267 (N_7267,In_657,In_2627);
and U7268 (N_7268,In_792,In_107);
nor U7269 (N_7269,In_1603,In_1412);
nand U7270 (N_7270,In_167,In_1746);
nor U7271 (N_7271,In_128,In_1666);
or U7272 (N_7272,In_1932,In_2386);
or U7273 (N_7273,In_770,In_881);
nor U7274 (N_7274,In_1342,In_2711);
nand U7275 (N_7275,In_693,In_1803);
and U7276 (N_7276,In_1933,In_1629);
and U7277 (N_7277,In_1986,In_1610);
nand U7278 (N_7278,In_1028,In_2935);
nand U7279 (N_7279,In_508,In_180);
or U7280 (N_7280,In_666,In_1564);
or U7281 (N_7281,In_577,In_195);
and U7282 (N_7282,In_1192,In_2541);
nand U7283 (N_7283,In_2690,In_1932);
and U7284 (N_7284,In_975,In_2719);
or U7285 (N_7285,In_1723,In_274);
nand U7286 (N_7286,In_311,In_1);
xor U7287 (N_7287,In_2748,In_1031);
or U7288 (N_7288,In_2431,In_411);
or U7289 (N_7289,In_688,In_1264);
nand U7290 (N_7290,In_2294,In_2524);
or U7291 (N_7291,In_918,In_2560);
nand U7292 (N_7292,In_1684,In_1254);
nor U7293 (N_7293,In_2852,In_395);
and U7294 (N_7294,In_608,In_1110);
nor U7295 (N_7295,In_1351,In_1357);
or U7296 (N_7296,In_403,In_1369);
nand U7297 (N_7297,In_139,In_1393);
or U7298 (N_7298,In_1897,In_727);
nor U7299 (N_7299,In_1666,In_1220);
or U7300 (N_7300,In_2252,In_2095);
nor U7301 (N_7301,In_1394,In_2978);
and U7302 (N_7302,In_2851,In_1518);
or U7303 (N_7303,In_99,In_911);
nand U7304 (N_7304,In_1995,In_801);
and U7305 (N_7305,In_657,In_2378);
and U7306 (N_7306,In_1393,In_1362);
or U7307 (N_7307,In_422,In_983);
or U7308 (N_7308,In_2637,In_2554);
nor U7309 (N_7309,In_2752,In_1201);
nor U7310 (N_7310,In_212,In_2917);
and U7311 (N_7311,In_836,In_1819);
nand U7312 (N_7312,In_1820,In_2176);
nor U7313 (N_7313,In_1651,In_1285);
nor U7314 (N_7314,In_1359,In_2810);
or U7315 (N_7315,In_2201,In_893);
or U7316 (N_7316,In_410,In_478);
or U7317 (N_7317,In_98,In_1241);
nand U7318 (N_7318,In_353,In_2464);
nor U7319 (N_7319,In_2731,In_993);
and U7320 (N_7320,In_2414,In_2273);
and U7321 (N_7321,In_925,In_1771);
and U7322 (N_7322,In_1388,In_1592);
and U7323 (N_7323,In_621,In_2945);
and U7324 (N_7324,In_262,In_751);
or U7325 (N_7325,In_1106,In_1022);
or U7326 (N_7326,In_47,In_1560);
nand U7327 (N_7327,In_1410,In_254);
or U7328 (N_7328,In_2336,In_685);
and U7329 (N_7329,In_2890,In_1456);
and U7330 (N_7330,In_951,In_866);
nor U7331 (N_7331,In_1576,In_2108);
or U7332 (N_7332,In_2275,In_517);
nor U7333 (N_7333,In_297,In_1815);
and U7334 (N_7334,In_459,In_2327);
nand U7335 (N_7335,In_151,In_897);
and U7336 (N_7336,In_1160,In_161);
nor U7337 (N_7337,In_2801,In_2781);
or U7338 (N_7338,In_2863,In_2465);
or U7339 (N_7339,In_2304,In_978);
nand U7340 (N_7340,In_2881,In_1053);
nor U7341 (N_7341,In_2656,In_578);
nor U7342 (N_7342,In_1074,In_131);
or U7343 (N_7343,In_2151,In_1508);
and U7344 (N_7344,In_1149,In_551);
nor U7345 (N_7345,In_976,In_2109);
and U7346 (N_7346,In_574,In_2622);
nor U7347 (N_7347,In_1983,In_1984);
and U7348 (N_7348,In_1490,In_425);
and U7349 (N_7349,In_2454,In_416);
nand U7350 (N_7350,In_2,In_1747);
and U7351 (N_7351,In_310,In_1355);
nand U7352 (N_7352,In_2024,In_1419);
and U7353 (N_7353,In_1857,In_2464);
and U7354 (N_7354,In_2512,In_2190);
and U7355 (N_7355,In_1569,In_1029);
nor U7356 (N_7356,In_401,In_2840);
and U7357 (N_7357,In_519,In_1413);
nor U7358 (N_7358,In_1373,In_1380);
and U7359 (N_7359,In_2737,In_99);
and U7360 (N_7360,In_2265,In_2944);
nand U7361 (N_7361,In_2297,In_626);
and U7362 (N_7362,In_2790,In_883);
and U7363 (N_7363,In_1601,In_946);
nor U7364 (N_7364,In_20,In_2019);
nand U7365 (N_7365,In_419,In_2061);
and U7366 (N_7366,In_352,In_560);
or U7367 (N_7367,In_159,In_1892);
nor U7368 (N_7368,In_533,In_1212);
nor U7369 (N_7369,In_2473,In_248);
and U7370 (N_7370,In_2402,In_726);
or U7371 (N_7371,In_1279,In_2793);
nor U7372 (N_7372,In_455,In_1058);
nor U7373 (N_7373,In_2762,In_2119);
nand U7374 (N_7374,In_1088,In_2016);
or U7375 (N_7375,In_1038,In_323);
and U7376 (N_7376,In_1500,In_936);
or U7377 (N_7377,In_2707,In_2362);
or U7378 (N_7378,In_1462,In_2918);
nor U7379 (N_7379,In_2859,In_2855);
or U7380 (N_7380,In_1499,In_2646);
nor U7381 (N_7381,In_2210,In_1712);
nand U7382 (N_7382,In_888,In_160);
and U7383 (N_7383,In_2687,In_351);
nor U7384 (N_7384,In_2760,In_1703);
nand U7385 (N_7385,In_1400,In_940);
and U7386 (N_7386,In_1997,In_1633);
and U7387 (N_7387,In_1372,In_110);
and U7388 (N_7388,In_2161,In_2382);
or U7389 (N_7389,In_993,In_1509);
nand U7390 (N_7390,In_2837,In_239);
and U7391 (N_7391,In_2249,In_2118);
or U7392 (N_7392,In_360,In_1828);
nand U7393 (N_7393,In_2365,In_1310);
nor U7394 (N_7394,In_159,In_164);
nor U7395 (N_7395,In_913,In_2848);
nand U7396 (N_7396,In_2467,In_112);
nand U7397 (N_7397,In_1690,In_264);
nor U7398 (N_7398,In_359,In_2283);
xnor U7399 (N_7399,In_337,In_737);
or U7400 (N_7400,In_1831,In_2887);
xnor U7401 (N_7401,In_2451,In_1475);
or U7402 (N_7402,In_1224,In_898);
and U7403 (N_7403,In_1269,In_1521);
and U7404 (N_7404,In_1249,In_1536);
or U7405 (N_7405,In_2069,In_981);
nor U7406 (N_7406,In_2440,In_1398);
or U7407 (N_7407,In_1409,In_439);
nand U7408 (N_7408,In_213,In_2635);
nor U7409 (N_7409,In_1341,In_673);
nand U7410 (N_7410,In_2711,In_2843);
or U7411 (N_7411,In_1275,In_2846);
and U7412 (N_7412,In_1678,In_1792);
and U7413 (N_7413,In_2271,In_2592);
nand U7414 (N_7414,In_1248,In_687);
and U7415 (N_7415,In_608,In_287);
or U7416 (N_7416,In_2752,In_987);
nand U7417 (N_7417,In_430,In_610);
or U7418 (N_7418,In_2530,In_498);
or U7419 (N_7419,In_964,In_1017);
nor U7420 (N_7420,In_200,In_1884);
nor U7421 (N_7421,In_564,In_501);
nand U7422 (N_7422,In_2920,In_2338);
nand U7423 (N_7423,In_544,In_1398);
nand U7424 (N_7424,In_466,In_2920);
or U7425 (N_7425,In_1328,In_918);
nor U7426 (N_7426,In_899,In_1704);
nand U7427 (N_7427,In_1690,In_1562);
nor U7428 (N_7428,In_2851,In_1664);
or U7429 (N_7429,In_1794,In_2732);
nor U7430 (N_7430,In_2440,In_1518);
nor U7431 (N_7431,In_1315,In_1182);
xor U7432 (N_7432,In_2374,In_2572);
nor U7433 (N_7433,In_2922,In_312);
and U7434 (N_7434,In_1066,In_810);
and U7435 (N_7435,In_2395,In_1067);
and U7436 (N_7436,In_1302,In_1093);
and U7437 (N_7437,In_1772,In_2283);
nor U7438 (N_7438,In_2301,In_1929);
nor U7439 (N_7439,In_2228,In_1308);
and U7440 (N_7440,In_575,In_1716);
nor U7441 (N_7441,In_234,In_1562);
or U7442 (N_7442,In_2370,In_1206);
nand U7443 (N_7443,In_1959,In_34);
nor U7444 (N_7444,In_449,In_2323);
nor U7445 (N_7445,In_1997,In_1423);
nor U7446 (N_7446,In_1429,In_972);
xnor U7447 (N_7447,In_2119,In_1326);
and U7448 (N_7448,In_2137,In_45);
nor U7449 (N_7449,In_1893,In_1382);
or U7450 (N_7450,In_2543,In_982);
and U7451 (N_7451,In_2192,In_393);
nand U7452 (N_7452,In_53,In_823);
and U7453 (N_7453,In_1277,In_2006);
nor U7454 (N_7454,In_1588,In_2718);
or U7455 (N_7455,In_1058,In_1775);
or U7456 (N_7456,In_2171,In_304);
and U7457 (N_7457,In_2233,In_1936);
nand U7458 (N_7458,In_2131,In_2920);
or U7459 (N_7459,In_630,In_681);
nor U7460 (N_7460,In_520,In_2066);
nand U7461 (N_7461,In_1175,In_789);
nand U7462 (N_7462,In_1864,In_2756);
nor U7463 (N_7463,In_2278,In_882);
or U7464 (N_7464,In_2039,In_1519);
or U7465 (N_7465,In_125,In_1794);
nand U7466 (N_7466,In_617,In_379);
nand U7467 (N_7467,In_72,In_2118);
or U7468 (N_7468,In_1854,In_591);
or U7469 (N_7469,In_2687,In_1406);
or U7470 (N_7470,In_2710,In_1934);
nand U7471 (N_7471,In_1657,In_225);
and U7472 (N_7472,In_1708,In_199);
and U7473 (N_7473,In_2469,In_2753);
and U7474 (N_7474,In_2235,In_2415);
nor U7475 (N_7475,In_2634,In_41);
nor U7476 (N_7476,In_1694,In_1643);
nor U7477 (N_7477,In_100,In_1468);
and U7478 (N_7478,In_1479,In_1489);
or U7479 (N_7479,In_1860,In_456);
or U7480 (N_7480,In_2231,In_462);
or U7481 (N_7481,In_2132,In_2675);
or U7482 (N_7482,In_423,In_2711);
or U7483 (N_7483,In_293,In_2106);
nor U7484 (N_7484,In_1804,In_2251);
and U7485 (N_7485,In_409,In_807);
nor U7486 (N_7486,In_2680,In_2910);
nor U7487 (N_7487,In_1816,In_2429);
nor U7488 (N_7488,In_877,In_734);
nand U7489 (N_7489,In_1822,In_181);
or U7490 (N_7490,In_2366,In_2056);
nand U7491 (N_7491,In_1671,In_1771);
nor U7492 (N_7492,In_1796,In_596);
nand U7493 (N_7493,In_1878,In_546);
nor U7494 (N_7494,In_927,In_2596);
nor U7495 (N_7495,In_910,In_2461);
or U7496 (N_7496,In_1255,In_2944);
nor U7497 (N_7497,In_1028,In_2417);
and U7498 (N_7498,In_1319,In_2777);
and U7499 (N_7499,In_254,In_53);
nand U7500 (N_7500,In_2977,In_649);
and U7501 (N_7501,In_1307,In_2907);
or U7502 (N_7502,In_733,In_1083);
nor U7503 (N_7503,In_1604,In_1623);
nor U7504 (N_7504,In_421,In_0);
or U7505 (N_7505,In_1177,In_2785);
or U7506 (N_7506,In_1528,In_1603);
nor U7507 (N_7507,In_523,In_2810);
nand U7508 (N_7508,In_2726,In_539);
xor U7509 (N_7509,In_2325,In_761);
nand U7510 (N_7510,In_452,In_294);
nand U7511 (N_7511,In_67,In_1065);
and U7512 (N_7512,In_300,In_868);
or U7513 (N_7513,In_1826,In_1018);
xnor U7514 (N_7514,In_2250,In_387);
nor U7515 (N_7515,In_1035,In_1009);
nor U7516 (N_7516,In_629,In_459);
nand U7517 (N_7517,In_1782,In_2157);
or U7518 (N_7518,In_2795,In_2701);
and U7519 (N_7519,In_1440,In_1641);
nor U7520 (N_7520,In_1329,In_535);
or U7521 (N_7521,In_703,In_910);
nor U7522 (N_7522,In_1250,In_250);
and U7523 (N_7523,In_532,In_685);
nor U7524 (N_7524,In_2428,In_2993);
nor U7525 (N_7525,In_523,In_1233);
nor U7526 (N_7526,In_1985,In_2739);
or U7527 (N_7527,In_2452,In_1843);
nor U7528 (N_7528,In_1092,In_600);
nand U7529 (N_7529,In_2464,In_210);
nor U7530 (N_7530,In_729,In_198);
nand U7531 (N_7531,In_2300,In_300);
nor U7532 (N_7532,In_1413,In_1274);
or U7533 (N_7533,In_877,In_2340);
nor U7534 (N_7534,In_2416,In_2883);
xor U7535 (N_7535,In_333,In_2367);
nor U7536 (N_7536,In_2050,In_987);
nand U7537 (N_7537,In_1742,In_1667);
or U7538 (N_7538,In_147,In_448);
nand U7539 (N_7539,In_592,In_913);
or U7540 (N_7540,In_202,In_2783);
nor U7541 (N_7541,In_1858,In_521);
nand U7542 (N_7542,In_847,In_2790);
nand U7543 (N_7543,In_841,In_2728);
and U7544 (N_7544,In_1654,In_167);
nand U7545 (N_7545,In_1217,In_2403);
and U7546 (N_7546,In_1315,In_2323);
nand U7547 (N_7547,In_1136,In_670);
or U7548 (N_7548,In_1588,In_1490);
nor U7549 (N_7549,In_1817,In_2626);
nand U7550 (N_7550,In_39,In_463);
nand U7551 (N_7551,In_623,In_2197);
nor U7552 (N_7552,In_2426,In_2074);
or U7553 (N_7553,In_1849,In_839);
or U7554 (N_7554,In_1453,In_938);
or U7555 (N_7555,In_2445,In_1278);
nand U7556 (N_7556,In_122,In_1474);
nor U7557 (N_7557,In_32,In_2853);
and U7558 (N_7558,In_1292,In_2281);
nand U7559 (N_7559,In_40,In_2492);
nand U7560 (N_7560,In_2122,In_1796);
nand U7561 (N_7561,In_2779,In_1051);
nor U7562 (N_7562,In_1588,In_2141);
nand U7563 (N_7563,In_784,In_1848);
nor U7564 (N_7564,In_2297,In_2287);
or U7565 (N_7565,In_1345,In_2976);
nand U7566 (N_7566,In_1129,In_2706);
nor U7567 (N_7567,In_2797,In_2800);
nand U7568 (N_7568,In_547,In_2487);
xor U7569 (N_7569,In_1787,In_1042);
or U7570 (N_7570,In_1535,In_2743);
nand U7571 (N_7571,In_876,In_2360);
nand U7572 (N_7572,In_1325,In_1902);
and U7573 (N_7573,In_760,In_146);
and U7574 (N_7574,In_777,In_537);
and U7575 (N_7575,In_1767,In_888);
nand U7576 (N_7576,In_572,In_1841);
nand U7577 (N_7577,In_2866,In_1577);
xor U7578 (N_7578,In_235,In_1833);
nand U7579 (N_7579,In_2502,In_2867);
nor U7580 (N_7580,In_470,In_747);
nor U7581 (N_7581,In_1108,In_915);
or U7582 (N_7582,In_2667,In_70);
or U7583 (N_7583,In_1503,In_763);
nor U7584 (N_7584,In_2012,In_39);
or U7585 (N_7585,In_2327,In_725);
nor U7586 (N_7586,In_2439,In_1898);
and U7587 (N_7587,In_1197,In_2509);
or U7588 (N_7588,In_849,In_619);
nand U7589 (N_7589,In_1571,In_1596);
nor U7590 (N_7590,In_2257,In_757);
nand U7591 (N_7591,In_1857,In_668);
nor U7592 (N_7592,In_1773,In_391);
or U7593 (N_7593,In_544,In_348);
and U7594 (N_7594,In_2858,In_975);
and U7595 (N_7595,In_1038,In_2814);
nor U7596 (N_7596,In_120,In_23);
nand U7597 (N_7597,In_2416,In_1844);
nand U7598 (N_7598,In_887,In_388);
and U7599 (N_7599,In_80,In_2811);
nor U7600 (N_7600,In_1148,In_1286);
nand U7601 (N_7601,In_1487,In_2416);
or U7602 (N_7602,In_1082,In_1531);
nand U7603 (N_7603,In_2374,In_2287);
nand U7604 (N_7604,In_2295,In_1925);
and U7605 (N_7605,In_2256,In_2593);
or U7606 (N_7606,In_1730,In_2791);
and U7607 (N_7607,In_1491,In_2925);
and U7608 (N_7608,In_894,In_2951);
and U7609 (N_7609,In_2756,In_34);
nor U7610 (N_7610,In_2010,In_548);
or U7611 (N_7611,In_2029,In_2322);
nor U7612 (N_7612,In_2418,In_937);
nor U7613 (N_7613,In_1840,In_1087);
nand U7614 (N_7614,In_968,In_2400);
nand U7615 (N_7615,In_1840,In_1256);
nor U7616 (N_7616,In_78,In_2378);
nand U7617 (N_7617,In_1611,In_34);
or U7618 (N_7618,In_2680,In_2595);
or U7619 (N_7619,In_2766,In_2449);
and U7620 (N_7620,In_2456,In_1343);
nor U7621 (N_7621,In_1236,In_286);
nand U7622 (N_7622,In_845,In_995);
or U7623 (N_7623,In_1286,In_245);
and U7624 (N_7624,In_657,In_832);
and U7625 (N_7625,In_2965,In_2957);
or U7626 (N_7626,In_1951,In_895);
nor U7627 (N_7627,In_2317,In_2263);
and U7628 (N_7628,In_2042,In_2445);
nor U7629 (N_7629,In_128,In_1821);
or U7630 (N_7630,In_2862,In_1607);
and U7631 (N_7631,In_1431,In_178);
or U7632 (N_7632,In_509,In_947);
or U7633 (N_7633,In_631,In_530);
and U7634 (N_7634,In_2602,In_2033);
nand U7635 (N_7635,In_318,In_1211);
nor U7636 (N_7636,In_2899,In_175);
or U7637 (N_7637,In_2926,In_1663);
nand U7638 (N_7638,In_2539,In_180);
or U7639 (N_7639,In_589,In_502);
or U7640 (N_7640,In_217,In_70);
and U7641 (N_7641,In_1477,In_2978);
or U7642 (N_7642,In_486,In_1573);
nand U7643 (N_7643,In_459,In_1109);
nand U7644 (N_7644,In_1876,In_2115);
nand U7645 (N_7645,In_2767,In_2092);
nor U7646 (N_7646,In_216,In_2352);
nor U7647 (N_7647,In_2415,In_1421);
nand U7648 (N_7648,In_73,In_1022);
or U7649 (N_7649,In_1424,In_570);
and U7650 (N_7650,In_1185,In_1688);
or U7651 (N_7651,In_1542,In_527);
nand U7652 (N_7652,In_2973,In_1788);
nor U7653 (N_7653,In_988,In_2304);
or U7654 (N_7654,In_2791,In_86);
nor U7655 (N_7655,In_1741,In_1765);
and U7656 (N_7656,In_1611,In_457);
nand U7657 (N_7657,In_279,In_2969);
or U7658 (N_7658,In_1081,In_2139);
or U7659 (N_7659,In_658,In_843);
nor U7660 (N_7660,In_2788,In_1332);
nand U7661 (N_7661,In_1920,In_1);
nand U7662 (N_7662,In_1365,In_2366);
nor U7663 (N_7663,In_1009,In_672);
nand U7664 (N_7664,In_2212,In_1415);
or U7665 (N_7665,In_1316,In_750);
nand U7666 (N_7666,In_2671,In_934);
or U7667 (N_7667,In_264,In_2129);
or U7668 (N_7668,In_2034,In_468);
nand U7669 (N_7669,In_2278,In_1994);
and U7670 (N_7670,In_2550,In_2312);
or U7671 (N_7671,In_2724,In_2922);
nand U7672 (N_7672,In_986,In_477);
or U7673 (N_7673,In_2066,In_287);
or U7674 (N_7674,In_2369,In_2987);
and U7675 (N_7675,In_1690,In_1408);
nor U7676 (N_7676,In_2701,In_2063);
and U7677 (N_7677,In_1893,In_307);
and U7678 (N_7678,In_2404,In_2581);
or U7679 (N_7679,In_2617,In_910);
or U7680 (N_7680,In_2137,In_270);
nand U7681 (N_7681,In_242,In_1393);
nor U7682 (N_7682,In_201,In_2388);
or U7683 (N_7683,In_96,In_1504);
and U7684 (N_7684,In_478,In_164);
nand U7685 (N_7685,In_2528,In_1449);
or U7686 (N_7686,In_975,In_2144);
nor U7687 (N_7687,In_781,In_535);
or U7688 (N_7688,In_2851,In_2146);
nor U7689 (N_7689,In_497,In_2303);
nor U7690 (N_7690,In_2381,In_643);
or U7691 (N_7691,In_483,In_2821);
nor U7692 (N_7692,In_1361,In_848);
or U7693 (N_7693,In_1828,In_545);
and U7694 (N_7694,In_889,In_2969);
nor U7695 (N_7695,In_952,In_810);
and U7696 (N_7696,In_465,In_220);
nand U7697 (N_7697,In_315,In_1696);
and U7698 (N_7698,In_1355,In_1247);
and U7699 (N_7699,In_1743,In_1328);
and U7700 (N_7700,In_826,In_2500);
nor U7701 (N_7701,In_1765,In_1791);
nor U7702 (N_7702,In_1509,In_1321);
nor U7703 (N_7703,In_1294,In_820);
nand U7704 (N_7704,In_2167,In_2786);
nand U7705 (N_7705,In_1163,In_2294);
and U7706 (N_7706,In_2550,In_2865);
nand U7707 (N_7707,In_678,In_297);
nor U7708 (N_7708,In_2102,In_2996);
and U7709 (N_7709,In_298,In_1399);
or U7710 (N_7710,In_311,In_1811);
nor U7711 (N_7711,In_1679,In_2471);
or U7712 (N_7712,In_1730,In_2320);
nand U7713 (N_7713,In_205,In_380);
and U7714 (N_7714,In_1268,In_483);
and U7715 (N_7715,In_2376,In_1245);
or U7716 (N_7716,In_1666,In_1322);
nor U7717 (N_7717,In_1970,In_2273);
and U7718 (N_7718,In_696,In_2494);
or U7719 (N_7719,In_1735,In_256);
or U7720 (N_7720,In_831,In_1656);
nor U7721 (N_7721,In_2391,In_1942);
xor U7722 (N_7722,In_372,In_617);
and U7723 (N_7723,In_485,In_1180);
or U7724 (N_7724,In_645,In_2122);
nor U7725 (N_7725,In_2281,In_884);
nor U7726 (N_7726,In_1028,In_2230);
nor U7727 (N_7727,In_1003,In_1344);
nand U7728 (N_7728,In_1648,In_1974);
or U7729 (N_7729,In_2484,In_1503);
and U7730 (N_7730,In_465,In_1387);
nor U7731 (N_7731,In_1303,In_938);
and U7732 (N_7732,In_1007,In_2585);
or U7733 (N_7733,In_1452,In_1278);
nand U7734 (N_7734,In_2357,In_2670);
nand U7735 (N_7735,In_1938,In_1913);
and U7736 (N_7736,In_2240,In_2599);
nor U7737 (N_7737,In_408,In_2407);
and U7738 (N_7738,In_1152,In_2428);
nand U7739 (N_7739,In_94,In_1901);
nand U7740 (N_7740,In_2174,In_1993);
nor U7741 (N_7741,In_2496,In_1702);
and U7742 (N_7742,In_251,In_1572);
or U7743 (N_7743,In_2377,In_2118);
or U7744 (N_7744,In_323,In_2263);
or U7745 (N_7745,In_1990,In_2597);
nor U7746 (N_7746,In_69,In_1776);
and U7747 (N_7747,In_1651,In_446);
nand U7748 (N_7748,In_1471,In_1282);
xnor U7749 (N_7749,In_771,In_2013);
nor U7750 (N_7750,In_1458,In_815);
or U7751 (N_7751,In_240,In_1966);
and U7752 (N_7752,In_255,In_61);
and U7753 (N_7753,In_619,In_1346);
nor U7754 (N_7754,In_2858,In_1748);
or U7755 (N_7755,In_1098,In_11);
nor U7756 (N_7756,In_2210,In_1661);
and U7757 (N_7757,In_2246,In_218);
nor U7758 (N_7758,In_2940,In_434);
nor U7759 (N_7759,In_1210,In_1897);
and U7760 (N_7760,In_2699,In_1034);
nor U7761 (N_7761,In_690,In_2253);
nor U7762 (N_7762,In_2508,In_1209);
nor U7763 (N_7763,In_2123,In_204);
xnor U7764 (N_7764,In_1409,In_685);
nor U7765 (N_7765,In_2127,In_78);
nand U7766 (N_7766,In_739,In_2077);
nor U7767 (N_7767,In_2948,In_2633);
nor U7768 (N_7768,In_2574,In_1228);
nand U7769 (N_7769,In_1806,In_1050);
nand U7770 (N_7770,In_2783,In_2483);
nand U7771 (N_7771,In_2294,In_2772);
nor U7772 (N_7772,In_2884,In_1431);
nand U7773 (N_7773,In_1074,In_1625);
nand U7774 (N_7774,In_2552,In_487);
nand U7775 (N_7775,In_1223,In_254);
nor U7776 (N_7776,In_1647,In_741);
nand U7777 (N_7777,In_1603,In_1202);
and U7778 (N_7778,In_2399,In_2114);
or U7779 (N_7779,In_1741,In_355);
nor U7780 (N_7780,In_1879,In_522);
or U7781 (N_7781,In_1687,In_2492);
and U7782 (N_7782,In_975,In_458);
nand U7783 (N_7783,In_2371,In_2840);
or U7784 (N_7784,In_2820,In_2843);
nor U7785 (N_7785,In_851,In_1599);
nor U7786 (N_7786,In_194,In_131);
nand U7787 (N_7787,In_979,In_2548);
nand U7788 (N_7788,In_957,In_446);
and U7789 (N_7789,In_1620,In_1643);
and U7790 (N_7790,In_1076,In_1302);
nor U7791 (N_7791,In_2229,In_2678);
nand U7792 (N_7792,In_1098,In_2739);
or U7793 (N_7793,In_907,In_1343);
or U7794 (N_7794,In_102,In_1962);
or U7795 (N_7795,In_2242,In_1393);
nand U7796 (N_7796,In_1522,In_161);
or U7797 (N_7797,In_2798,In_240);
nor U7798 (N_7798,In_622,In_2232);
nand U7799 (N_7799,In_1428,In_761);
nor U7800 (N_7800,In_1942,In_970);
and U7801 (N_7801,In_193,In_853);
nand U7802 (N_7802,In_565,In_1770);
or U7803 (N_7803,In_374,In_2535);
nor U7804 (N_7804,In_2991,In_1153);
and U7805 (N_7805,In_1869,In_44);
and U7806 (N_7806,In_1072,In_1865);
nor U7807 (N_7807,In_1757,In_2912);
or U7808 (N_7808,In_1466,In_443);
nand U7809 (N_7809,In_2337,In_2640);
or U7810 (N_7810,In_932,In_2103);
or U7811 (N_7811,In_1420,In_2952);
or U7812 (N_7812,In_2643,In_825);
nand U7813 (N_7813,In_513,In_2676);
xor U7814 (N_7814,In_1474,In_1716);
or U7815 (N_7815,In_2410,In_737);
nor U7816 (N_7816,In_2634,In_2242);
nor U7817 (N_7817,In_390,In_873);
nor U7818 (N_7818,In_2680,In_1278);
nand U7819 (N_7819,In_1441,In_241);
and U7820 (N_7820,In_1755,In_2863);
and U7821 (N_7821,In_1433,In_438);
and U7822 (N_7822,In_1396,In_2855);
and U7823 (N_7823,In_500,In_1845);
and U7824 (N_7824,In_2423,In_2194);
or U7825 (N_7825,In_2733,In_2392);
nor U7826 (N_7826,In_2205,In_1072);
nand U7827 (N_7827,In_2291,In_835);
nor U7828 (N_7828,In_985,In_1486);
or U7829 (N_7829,In_712,In_876);
nor U7830 (N_7830,In_1494,In_1696);
and U7831 (N_7831,In_1815,In_1479);
nand U7832 (N_7832,In_831,In_1615);
nor U7833 (N_7833,In_1188,In_515);
or U7834 (N_7834,In_1769,In_1295);
or U7835 (N_7835,In_1929,In_1173);
nor U7836 (N_7836,In_787,In_741);
nand U7837 (N_7837,In_1091,In_2127);
and U7838 (N_7838,In_1385,In_750);
or U7839 (N_7839,In_176,In_490);
nor U7840 (N_7840,In_637,In_1286);
and U7841 (N_7841,In_2463,In_2823);
nor U7842 (N_7842,In_2758,In_1045);
and U7843 (N_7843,In_2802,In_1967);
or U7844 (N_7844,In_2943,In_1825);
nand U7845 (N_7845,In_1358,In_2502);
and U7846 (N_7846,In_1882,In_2455);
nand U7847 (N_7847,In_2463,In_1749);
and U7848 (N_7848,In_486,In_620);
or U7849 (N_7849,In_920,In_1091);
or U7850 (N_7850,In_1732,In_2714);
or U7851 (N_7851,In_1238,In_2121);
nor U7852 (N_7852,In_1116,In_1064);
nor U7853 (N_7853,In_2309,In_2602);
or U7854 (N_7854,In_2458,In_2372);
nor U7855 (N_7855,In_1701,In_505);
or U7856 (N_7856,In_1500,In_119);
xor U7857 (N_7857,In_1140,In_165);
nand U7858 (N_7858,In_692,In_1907);
nor U7859 (N_7859,In_259,In_541);
or U7860 (N_7860,In_129,In_1213);
nor U7861 (N_7861,In_116,In_524);
nor U7862 (N_7862,In_1538,In_2389);
nor U7863 (N_7863,In_1212,In_37);
or U7864 (N_7864,In_1766,In_2491);
nor U7865 (N_7865,In_774,In_2677);
nor U7866 (N_7866,In_452,In_823);
or U7867 (N_7867,In_273,In_2780);
nor U7868 (N_7868,In_2134,In_2627);
or U7869 (N_7869,In_2360,In_1641);
or U7870 (N_7870,In_1521,In_964);
nor U7871 (N_7871,In_1430,In_2352);
and U7872 (N_7872,In_1913,In_55);
nand U7873 (N_7873,In_2741,In_2988);
nand U7874 (N_7874,In_2505,In_1815);
and U7875 (N_7875,In_996,In_2458);
nand U7876 (N_7876,In_1268,In_2439);
and U7877 (N_7877,In_702,In_1172);
nor U7878 (N_7878,In_1165,In_2818);
or U7879 (N_7879,In_793,In_1548);
nand U7880 (N_7880,In_1830,In_629);
xor U7881 (N_7881,In_2003,In_1938);
or U7882 (N_7882,In_347,In_267);
and U7883 (N_7883,In_180,In_1549);
nor U7884 (N_7884,In_1571,In_967);
nor U7885 (N_7885,In_1889,In_1481);
nand U7886 (N_7886,In_2040,In_1495);
and U7887 (N_7887,In_2444,In_2745);
and U7888 (N_7888,In_201,In_951);
nor U7889 (N_7889,In_545,In_1342);
and U7890 (N_7890,In_2032,In_18);
nor U7891 (N_7891,In_1837,In_877);
or U7892 (N_7892,In_211,In_2000);
and U7893 (N_7893,In_547,In_1090);
nor U7894 (N_7894,In_2662,In_442);
nand U7895 (N_7895,In_2377,In_2510);
nand U7896 (N_7896,In_502,In_1371);
nand U7897 (N_7897,In_1518,In_1994);
or U7898 (N_7898,In_1676,In_2356);
nand U7899 (N_7899,In_2357,In_2482);
nor U7900 (N_7900,In_2650,In_1784);
or U7901 (N_7901,In_556,In_1996);
and U7902 (N_7902,In_253,In_158);
nand U7903 (N_7903,In_351,In_1190);
or U7904 (N_7904,In_252,In_2600);
and U7905 (N_7905,In_2051,In_2709);
nand U7906 (N_7906,In_2497,In_2968);
or U7907 (N_7907,In_1006,In_2880);
nand U7908 (N_7908,In_2219,In_2409);
nand U7909 (N_7909,In_2632,In_2163);
nand U7910 (N_7910,In_1345,In_447);
and U7911 (N_7911,In_2630,In_2901);
nor U7912 (N_7912,In_2824,In_2623);
nand U7913 (N_7913,In_1800,In_421);
or U7914 (N_7914,In_235,In_2327);
and U7915 (N_7915,In_552,In_1819);
or U7916 (N_7916,In_1488,In_2255);
nand U7917 (N_7917,In_822,In_2989);
or U7918 (N_7918,In_2872,In_2735);
nor U7919 (N_7919,In_1642,In_292);
or U7920 (N_7920,In_24,In_1944);
nor U7921 (N_7921,In_523,In_2354);
or U7922 (N_7922,In_2817,In_2856);
or U7923 (N_7923,In_2096,In_673);
and U7924 (N_7924,In_1310,In_1884);
or U7925 (N_7925,In_232,In_390);
and U7926 (N_7926,In_1723,In_202);
nand U7927 (N_7927,In_1798,In_1850);
and U7928 (N_7928,In_844,In_1247);
nand U7929 (N_7929,In_2297,In_1034);
and U7930 (N_7930,In_1578,In_2786);
nor U7931 (N_7931,In_2711,In_968);
or U7932 (N_7932,In_1856,In_1928);
and U7933 (N_7933,In_2416,In_1789);
nor U7934 (N_7934,In_2069,In_113);
or U7935 (N_7935,In_1150,In_1348);
or U7936 (N_7936,In_1177,In_1388);
xor U7937 (N_7937,In_1966,In_1175);
nor U7938 (N_7938,In_1895,In_955);
and U7939 (N_7939,In_547,In_2621);
and U7940 (N_7940,In_1214,In_578);
nand U7941 (N_7941,In_859,In_2863);
and U7942 (N_7942,In_508,In_760);
nand U7943 (N_7943,In_1554,In_1220);
nor U7944 (N_7944,In_1521,In_1342);
nand U7945 (N_7945,In_2672,In_2184);
nor U7946 (N_7946,In_741,In_1877);
nor U7947 (N_7947,In_1752,In_1053);
nor U7948 (N_7948,In_2732,In_146);
or U7949 (N_7949,In_1968,In_1349);
nor U7950 (N_7950,In_2086,In_74);
or U7951 (N_7951,In_1069,In_762);
and U7952 (N_7952,In_540,In_1378);
nand U7953 (N_7953,In_1295,In_1864);
and U7954 (N_7954,In_1732,In_1852);
or U7955 (N_7955,In_379,In_285);
or U7956 (N_7956,In_831,In_2978);
nor U7957 (N_7957,In_2157,In_2564);
nor U7958 (N_7958,In_859,In_16);
nor U7959 (N_7959,In_1226,In_545);
nor U7960 (N_7960,In_1780,In_2464);
nand U7961 (N_7961,In_2601,In_2183);
nand U7962 (N_7962,In_2046,In_445);
or U7963 (N_7963,In_2674,In_21);
nand U7964 (N_7964,In_1176,In_1337);
or U7965 (N_7965,In_284,In_2281);
and U7966 (N_7966,In_471,In_141);
nand U7967 (N_7967,In_2795,In_2926);
and U7968 (N_7968,In_2219,In_1159);
and U7969 (N_7969,In_549,In_2176);
and U7970 (N_7970,In_1846,In_2827);
nand U7971 (N_7971,In_1203,In_2810);
and U7972 (N_7972,In_25,In_1873);
and U7973 (N_7973,In_2408,In_1736);
nor U7974 (N_7974,In_944,In_2350);
nor U7975 (N_7975,In_1860,In_2985);
or U7976 (N_7976,In_846,In_769);
or U7977 (N_7977,In_2814,In_2976);
or U7978 (N_7978,In_479,In_102);
and U7979 (N_7979,In_124,In_619);
nor U7980 (N_7980,In_365,In_1733);
and U7981 (N_7981,In_1314,In_2219);
nor U7982 (N_7982,In_2499,In_558);
nor U7983 (N_7983,In_2287,In_270);
nor U7984 (N_7984,In_1108,In_2282);
or U7985 (N_7985,In_1965,In_483);
and U7986 (N_7986,In_2469,In_19);
or U7987 (N_7987,In_184,In_1235);
or U7988 (N_7988,In_228,In_1126);
or U7989 (N_7989,In_817,In_1302);
or U7990 (N_7990,In_886,In_765);
nor U7991 (N_7991,In_1511,In_2914);
or U7992 (N_7992,In_2987,In_293);
nand U7993 (N_7993,In_1702,In_2917);
or U7994 (N_7994,In_2039,In_2167);
nor U7995 (N_7995,In_1535,In_1297);
nand U7996 (N_7996,In_2107,In_2978);
or U7997 (N_7997,In_1445,In_1148);
nor U7998 (N_7998,In_1407,In_2521);
and U7999 (N_7999,In_62,In_1754);
nor U8000 (N_8000,In_59,In_2497);
xor U8001 (N_8001,In_2503,In_170);
nor U8002 (N_8002,In_262,In_2625);
nand U8003 (N_8003,In_577,In_2874);
nand U8004 (N_8004,In_46,In_276);
and U8005 (N_8005,In_2013,In_2252);
or U8006 (N_8006,In_749,In_303);
nor U8007 (N_8007,In_2465,In_55);
nor U8008 (N_8008,In_532,In_2315);
nor U8009 (N_8009,In_2179,In_1970);
nand U8010 (N_8010,In_680,In_511);
nor U8011 (N_8011,In_327,In_712);
or U8012 (N_8012,In_1055,In_769);
nor U8013 (N_8013,In_569,In_1789);
nor U8014 (N_8014,In_1184,In_1946);
nand U8015 (N_8015,In_2977,In_158);
and U8016 (N_8016,In_1520,In_1159);
or U8017 (N_8017,In_967,In_193);
nor U8018 (N_8018,In_593,In_1915);
or U8019 (N_8019,In_2182,In_2945);
nor U8020 (N_8020,In_436,In_1624);
nand U8021 (N_8021,In_2253,In_1331);
nor U8022 (N_8022,In_2324,In_231);
and U8023 (N_8023,In_377,In_2917);
nand U8024 (N_8024,In_1716,In_2324);
nand U8025 (N_8025,In_918,In_15);
and U8026 (N_8026,In_515,In_2025);
and U8027 (N_8027,In_2178,In_2328);
or U8028 (N_8028,In_2057,In_2017);
nand U8029 (N_8029,In_2534,In_1371);
or U8030 (N_8030,In_1910,In_231);
nand U8031 (N_8031,In_1050,In_2378);
nor U8032 (N_8032,In_1952,In_118);
and U8033 (N_8033,In_2982,In_1253);
nand U8034 (N_8034,In_2819,In_659);
nor U8035 (N_8035,In_1069,In_2213);
and U8036 (N_8036,In_1682,In_2202);
nand U8037 (N_8037,In_1297,In_1880);
and U8038 (N_8038,In_2970,In_632);
nand U8039 (N_8039,In_2160,In_1726);
or U8040 (N_8040,In_1358,In_178);
and U8041 (N_8041,In_1126,In_1440);
and U8042 (N_8042,In_982,In_469);
nand U8043 (N_8043,In_1710,In_846);
nand U8044 (N_8044,In_1598,In_233);
nand U8045 (N_8045,In_46,In_2492);
nor U8046 (N_8046,In_183,In_68);
or U8047 (N_8047,In_794,In_421);
or U8048 (N_8048,In_1909,In_955);
or U8049 (N_8049,In_1323,In_1080);
and U8050 (N_8050,In_2693,In_424);
nand U8051 (N_8051,In_2649,In_2086);
or U8052 (N_8052,In_2464,In_306);
nor U8053 (N_8053,In_1572,In_1230);
nor U8054 (N_8054,In_2523,In_422);
and U8055 (N_8055,In_2050,In_1936);
or U8056 (N_8056,In_2350,In_1832);
nor U8057 (N_8057,In_2868,In_2396);
or U8058 (N_8058,In_840,In_1165);
nor U8059 (N_8059,In_121,In_2604);
or U8060 (N_8060,In_2432,In_1096);
and U8061 (N_8061,In_147,In_1152);
or U8062 (N_8062,In_1232,In_2845);
nand U8063 (N_8063,In_774,In_1200);
nand U8064 (N_8064,In_1868,In_847);
nor U8065 (N_8065,In_2804,In_1467);
or U8066 (N_8066,In_2772,In_2532);
nor U8067 (N_8067,In_2694,In_1850);
nand U8068 (N_8068,In_2863,In_2038);
or U8069 (N_8069,In_2535,In_1846);
or U8070 (N_8070,In_1049,In_930);
nand U8071 (N_8071,In_2301,In_1010);
nor U8072 (N_8072,In_1896,In_1262);
or U8073 (N_8073,In_2272,In_2302);
xnor U8074 (N_8074,In_2887,In_477);
or U8075 (N_8075,In_618,In_1718);
nor U8076 (N_8076,In_1077,In_1460);
nand U8077 (N_8077,In_220,In_79);
or U8078 (N_8078,In_2260,In_294);
nand U8079 (N_8079,In_1213,In_2996);
nor U8080 (N_8080,In_2511,In_386);
nor U8081 (N_8081,In_1540,In_1745);
or U8082 (N_8082,In_775,In_1578);
nand U8083 (N_8083,In_2640,In_456);
nor U8084 (N_8084,In_1999,In_696);
and U8085 (N_8085,In_2875,In_1471);
and U8086 (N_8086,In_752,In_1923);
nor U8087 (N_8087,In_2141,In_556);
nand U8088 (N_8088,In_2866,In_378);
nor U8089 (N_8089,In_187,In_2800);
nand U8090 (N_8090,In_30,In_746);
or U8091 (N_8091,In_2466,In_2166);
or U8092 (N_8092,In_2274,In_914);
or U8093 (N_8093,In_597,In_499);
or U8094 (N_8094,In_268,In_2763);
or U8095 (N_8095,In_1928,In_2441);
nor U8096 (N_8096,In_1818,In_1311);
and U8097 (N_8097,In_683,In_61);
nor U8098 (N_8098,In_436,In_1860);
nor U8099 (N_8099,In_1897,In_1836);
and U8100 (N_8100,In_2188,In_1252);
nor U8101 (N_8101,In_152,In_1336);
nand U8102 (N_8102,In_1853,In_151);
nor U8103 (N_8103,In_1452,In_2556);
nand U8104 (N_8104,In_1504,In_283);
nand U8105 (N_8105,In_2233,In_284);
nand U8106 (N_8106,In_2494,In_2927);
nor U8107 (N_8107,In_2030,In_2571);
nand U8108 (N_8108,In_2171,In_305);
or U8109 (N_8109,In_1837,In_2810);
or U8110 (N_8110,In_160,In_1791);
nor U8111 (N_8111,In_374,In_1937);
and U8112 (N_8112,In_2518,In_2905);
and U8113 (N_8113,In_1103,In_970);
or U8114 (N_8114,In_1948,In_478);
nor U8115 (N_8115,In_168,In_1959);
or U8116 (N_8116,In_1304,In_42);
nor U8117 (N_8117,In_2327,In_2706);
nand U8118 (N_8118,In_529,In_1290);
and U8119 (N_8119,In_1041,In_1808);
and U8120 (N_8120,In_478,In_914);
and U8121 (N_8121,In_331,In_873);
and U8122 (N_8122,In_2129,In_2086);
nand U8123 (N_8123,In_1240,In_2751);
nand U8124 (N_8124,In_2847,In_1309);
nor U8125 (N_8125,In_1997,In_759);
nor U8126 (N_8126,In_2096,In_2731);
nand U8127 (N_8127,In_2171,In_2552);
nand U8128 (N_8128,In_2719,In_1449);
nand U8129 (N_8129,In_135,In_456);
nand U8130 (N_8130,In_2738,In_195);
or U8131 (N_8131,In_1062,In_4);
and U8132 (N_8132,In_940,In_445);
and U8133 (N_8133,In_287,In_1512);
or U8134 (N_8134,In_2926,In_17);
and U8135 (N_8135,In_1477,In_1169);
and U8136 (N_8136,In_1674,In_2092);
nand U8137 (N_8137,In_2908,In_532);
or U8138 (N_8138,In_894,In_1313);
nand U8139 (N_8139,In_1205,In_2935);
nand U8140 (N_8140,In_868,In_819);
and U8141 (N_8141,In_2610,In_2518);
nand U8142 (N_8142,In_1379,In_1126);
nand U8143 (N_8143,In_391,In_1586);
nand U8144 (N_8144,In_1490,In_919);
nand U8145 (N_8145,In_548,In_2453);
nand U8146 (N_8146,In_173,In_1929);
nand U8147 (N_8147,In_401,In_2702);
nand U8148 (N_8148,In_206,In_2273);
or U8149 (N_8149,In_1233,In_1284);
or U8150 (N_8150,In_2832,In_1155);
nand U8151 (N_8151,In_2208,In_1789);
and U8152 (N_8152,In_1355,In_1168);
or U8153 (N_8153,In_2545,In_1743);
and U8154 (N_8154,In_235,In_2594);
and U8155 (N_8155,In_1546,In_1680);
nor U8156 (N_8156,In_58,In_1918);
and U8157 (N_8157,In_1309,In_1172);
and U8158 (N_8158,In_961,In_395);
and U8159 (N_8159,In_691,In_2444);
nor U8160 (N_8160,In_1379,In_1037);
nand U8161 (N_8161,In_2637,In_2615);
nand U8162 (N_8162,In_360,In_1616);
and U8163 (N_8163,In_166,In_679);
or U8164 (N_8164,In_2100,In_814);
nand U8165 (N_8165,In_2493,In_2548);
nand U8166 (N_8166,In_2819,In_1129);
or U8167 (N_8167,In_613,In_1263);
nand U8168 (N_8168,In_1375,In_1754);
nor U8169 (N_8169,In_1476,In_451);
or U8170 (N_8170,In_1454,In_1730);
and U8171 (N_8171,In_1906,In_843);
and U8172 (N_8172,In_2955,In_748);
and U8173 (N_8173,In_1778,In_2275);
nor U8174 (N_8174,In_651,In_1169);
or U8175 (N_8175,In_2370,In_2544);
xor U8176 (N_8176,In_2045,In_2206);
or U8177 (N_8177,In_2200,In_2615);
or U8178 (N_8178,In_2403,In_1054);
or U8179 (N_8179,In_2347,In_2205);
nor U8180 (N_8180,In_1545,In_128);
nand U8181 (N_8181,In_1399,In_1451);
nor U8182 (N_8182,In_2300,In_2957);
nor U8183 (N_8183,In_1726,In_2618);
and U8184 (N_8184,In_1861,In_2402);
and U8185 (N_8185,In_1664,In_2691);
or U8186 (N_8186,In_968,In_1863);
nor U8187 (N_8187,In_837,In_1758);
or U8188 (N_8188,In_1008,In_1780);
or U8189 (N_8189,In_306,In_2058);
nor U8190 (N_8190,In_2123,In_1465);
and U8191 (N_8191,In_2464,In_2802);
nand U8192 (N_8192,In_2604,In_134);
xnor U8193 (N_8193,In_575,In_929);
or U8194 (N_8194,In_2543,In_1635);
nor U8195 (N_8195,In_2770,In_2729);
or U8196 (N_8196,In_647,In_197);
nand U8197 (N_8197,In_1432,In_719);
and U8198 (N_8198,In_967,In_1033);
xor U8199 (N_8199,In_1376,In_1714);
and U8200 (N_8200,In_2922,In_1163);
nor U8201 (N_8201,In_582,In_2035);
or U8202 (N_8202,In_106,In_1886);
nor U8203 (N_8203,In_2175,In_2137);
nand U8204 (N_8204,In_852,In_2007);
or U8205 (N_8205,In_2986,In_2181);
nand U8206 (N_8206,In_1730,In_1131);
nand U8207 (N_8207,In_2641,In_2347);
or U8208 (N_8208,In_1611,In_1258);
or U8209 (N_8209,In_873,In_93);
nand U8210 (N_8210,In_66,In_1558);
nand U8211 (N_8211,In_2123,In_1963);
nor U8212 (N_8212,In_676,In_192);
and U8213 (N_8213,In_1966,In_2874);
or U8214 (N_8214,In_559,In_2763);
nand U8215 (N_8215,In_2760,In_2436);
or U8216 (N_8216,In_2193,In_1684);
nand U8217 (N_8217,In_1282,In_320);
nor U8218 (N_8218,In_1625,In_1981);
nand U8219 (N_8219,In_600,In_898);
nand U8220 (N_8220,In_2241,In_1801);
or U8221 (N_8221,In_1546,In_2092);
nor U8222 (N_8222,In_1167,In_2622);
nand U8223 (N_8223,In_2512,In_2780);
xnor U8224 (N_8224,In_1577,In_2058);
or U8225 (N_8225,In_655,In_2177);
or U8226 (N_8226,In_2931,In_2854);
nand U8227 (N_8227,In_247,In_2120);
nand U8228 (N_8228,In_2123,In_643);
or U8229 (N_8229,In_1168,In_1230);
and U8230 (N_8230,In_1858,In_548);
nor U8231 (N_8231,In_115,In_1592);
and U8232 (N_8232,In_1586,In_1783);
or U8233 (N_8233,In_369,In_2883);
nor U8234 (N_8234,In_2033,In_1449);
or U8235 (N_8235,In_2542,In_1627);
nand U8236 (N_8236,In_871,In_221);
or U8237 (N_8237,In_964,In_1901);
nand U8238 (N_8238,In_2926,In_1968);
or U8239 (N_8239,In_1572,In_2044);
nor U8240 (N_8240,In_2980,In_1273);
and U8241 (N_8241,In_1417,In_2300);
nand U8242 (N_8242,In_2006,In_567);
and U8243 (N_8243,In_1353,In_650);
or U8244 (N_8244,In_2733,In_1113);
nor U8245 (N_8245,In_2605,In_1552);
or U8246 (N_8246,In_2337,In_2044);
or U8247 (N_8247,In_2476,In_865);
nor U8248 (N_8248,In_1566,In_1760);
or U8249 (N_8249,In_495,In_146);
nand U8250 (N_8250,In_2056,In_1011);
and U8251 (N_8251,In_490,In_83);
nor U8252 (N_8252,In_2653,In_1201);
nor U8253 (N_8253,In_2664,In_611);
and U8254 (N_8254,In_727,In_1423);
xor U8255 (N_8255,In_699,In_2700);
and U8256 (N_8256,In_1969,In_2362);
or U8257 (N_8257,In_1823,In_1105);
or U8258 (N_8258,In_838,In_153);
nand U8259 (N_8259,In_1871,In_891);
or U8260 (N_8260,In_2781,In_486);
nand U8261 (N_8261,In_2401,In_2521);
nor U8262 (N_8262,In_852,In_226);
nor U8263 (N_8263,In_1926,In_1689);
nand U8264 (N_8264,In_1251,In_2208);
nor U8265 (N_8265,In_1379,In_985);
nor U8266 (N_8266,In_2245,In_2818);
nand U8267 (N_8267,In_576,In_1529);
nor U8268 (N_8268,In_1322,In_2072);
nor U8269 (N_8269,In_1105,In_1850);
and U8270 (N_8270,In_85,In_1695);
and U8271 (N_8271,In_264,In_122);
nand U8272 (N_8272,In_1228,In_2465);
nor U8273 (N_8273,In_2603,In_2884);
or U8274 (N_8274,In_1581,In_932);
nand U8275 (N_8275,In_756,In_345);
and U8276 (N_8276,In_1470,In_1282);
nand U8277 (N_8277,In_777,In_2334);
nor U8278 (N_8278,In_2099,In_1358);
nand U8279 (N_8279,In_2433,In_979);
and U8280 (N_8280,In_506,In_29);
nor U8281 (N_8281,In_2295,In_2284);
nand U8282 (N_8282,In_996,In_2061);
and U8283 (N_8283,In_987,In_2558);
nor U8284 (N_8284,In_1459,In_1723);
nand U8285 (N_8285,In_1691,In_1976);
and U8286 (N_8286,In_883,In_1407);
nand U8287 (N_8287,In_2009,In_2115);
nor U8288 (N_8288,In_1532,In_705);
and U8289 (N_8289,In_1450,In_1042);
nand U8290 (N_8290,In_336,In_259);
or U8291 (N_8291,In_374,In_1442);
and U8292 (N_8292,In_930,In_2210);
nor U8293 (N_8293,In_1542,In_1832);
or U8294 (N_8294,In_688,In_2151);
and U8295 (N_8295,In_345,In_2514);
or U8296 (N_8296,In_2568,In_2114);
or U8297 (N_8297,In_2192,In_1231);
nand U8298 (N_8298,In_1011,In_5);
nand U8299 (N_8299,In_2760,In_2747);
xor U8300 (N_8300,In_1263,In_2194);
nand U8301 (N_8301,In_2594,In_173);
nand U8302 (N_8302,In_1466,In_1086);
nand U8303 (N_8303,In_2042,In_2177);
nor U8304 (N_8304,In_774,In_881);
or U8305 (N_8305,In_2433,In_1415);
or U8306 (N_8306,In_782,In_670);
nor U8307 (N_8307,In_2187,In_1499);
nor U8308 (N_8308,In_1071,In_162);
nor U8309 (N_8309,In_1526,In_2618);
nand U8310 (N_8310,In_1073,In_942);
and U8311 (N_8311,In_1971,In_426);
nor U8312 (N_8312,In_476,In_369);
or U8313 (N_8313,In_2923,In_2730);
nand U8314 (N_8314,In_2169,In_2921);
and U8315 (N_8315,In_2516,In_989);
nor U8316 (N_8316,In_279,In_1897);
or U8317 (N_8317,In_502,In_2355);
nand U8318 (N_8318,In_585,In_1494);
and U8319 (N_8319,In_928,In_72);
nor U8320 (N_8320,In_2769,In_1868);
and U8321 (N_8321,In_924,In_1986);
or U8322 (N_8322,In_1438,In_953);
and U8323 (N_8323,In_40,In_2419);
nor U8324 (N_8324,In_298,In_2105);
or U8325 (N_8325,In_2100,In_1068);
nand U8326 (N_8326,In_1885,In_2389);
or U8327 (N_8327,In_2158,In_1482);
and U8328 (N_8328,In_1839,In_501);
xnor U8329 (N_8329,In_2969,In_819);
nand U8330 (N_8330,In_1606,In_866);
nand U8331 (N_8331,In_101,In_2272);
or U8332 (N_8332,In_1515,In_605);
nor U8333 (N_8333,In_608,In_1863);
or U8334 (N_8334,In_911,In_395);
nor U8335 (N_8335,In_2006,In_1718);
or U8336 (N_8336,In_1395,In_2355);
nand U8337 (N_8337,In_1714,In_969);
nand U8338 (N_8338,In_390,In_2668);
or U8339 (N_8339,In_1458,In_2785);
nand U8340 (N_8340,In_749,In_1380);
nand U8341 (N_8341,In_2500,In_1077);
nand U8342 (N_8342,In_2215,In_1457);
and U8343 (N_8343,In_2484,In_2912);
and U8344 (N_8344,In_790,In_793);
nand U8345 (N_8345,In_872,In_663);
nor U8346 (N_8346,In_1795,In_1967);
or U8347 (N_8347,In_43,In_2766);
and U8348 (N_8348,In_1215,In_2594);
or U8349 (N_8349,In_637,In_483);
or U8350 (N_8350,In_852,In_2350);
nor U8351 (N_8351,In_2196,In_1516);
nor U8352 (N_8352,In_1772,In_2644);
and U8353 (N_8353,In_1488,In_249);
nand U8354 (N_8354,In_337,In_1786);
or U8355 (N_8355,In_2638,In_1367);
and U8356 (N_8356,In_1426,In_2841);
nor U8357 (N_8357,In_1562,In_2987);
and U8358 (N_8358,In_1974,In_240);
and U8359 (N_8359,In_974,In_41);
and U8360 (N_8360,In_2427,In_2476);
or U8361 (N_8361,In_1595,In_2334);
or U8362 (N_8362,In_1490,In_2793);
nand U8363 (N_8363,In_2128,In_1509);
and U8364 (N_8364,In_2606,In_683);
or U8365 (N_8365,In_1694,In_2521);
or U8366 (N_8366,In_1541,In_1543);
nand U8367 (N_8367,In_1095,In_2858);
nor U8368 (N_8368,In_2495,In_1864);
or U8369 (N_8369,In_2471,In_2853);
nand U8370 (N_8370,In_2535,In_2217);
or U8371 (N_8371,In_99,In_554);
nor U8372 (N_8372,In_1124,In_1787);
nor U8373 (N_8373,In_1473,In_840);
nor U8374 (N_8374,In_302,In_524);
nor U8375 (N_8375,In_2777,In_581);
nand U8376 (N_8376,In_490,In_1276);
or U8377 (N_8377,In_2472,In_2070);
nor U8378 (N_8378,In_788,In_2537);
nand U8379 (N_8379,In_113,In_1419);
and U8380 (N_8380,In_1351,In_1032);
or U8381 (N_8381,In_200,In_2408);
and U8382 (N_8382,In_2758,In_437);
nor U8383 (N_8383,In_263,In_2993);
nand U8384 (N_8384,In_2871,In_1691);
nor U8385 (N_8385,In_41,In_841);
and U8386 (N_8386,In_359,In_2331);
nand U8387 (N_8387,In_2667,In_861);
nand U8388 (N_8388,In_1178,In_2767);
nand U8389 (N_8389,In_838,In_7);
or U8390 (N_8390,In_1271,In_1889);
nor U8391 (N_8391,In_2264,In_1144);
nand U8392 (N_8392,In_2970,In_440);
nor U8393 (N_8393,In_1990,In_1576);
and U8394 (N_8394,In_432,In_1183);
nand U8395 (N_8395,In_2891,In_1414);
xnor U8396 (N_8396,In_1689,In_1331);
nand U8397 (N_8397,In_988,In_1953);
nor U8398 (N_8398,In_331,In_1241);
nor U8399 (N_8399,In_1391,In_1344);
or U8400 (N_8400,In_1971,In_1107);
nor U8401 (N_8401,In_2702,In_2319);
nor U8402 (N_8402,In_16,In_1653);
nor U8403 (N_8403,In_2389,In_1021);
and U8404 (N_8404,In_2633,In_2131);
nor U8405 (N_8405,In_240,In_909);
nor U8406 (N_8406,In_2883,In_2663);
nor U8407 (N_8407,In_1451,In_2794);
and U8408 (N_8408,In_2959,In_2324);
or U8409 (N_8409,In_2517,In_2273);
or U8410 (N_8410,In_445,In_1884);
and U8411 (N_8411,In_950,In_1267);
nand U8412 (N_8412,In_339,In_2329);
nand U8413 (N_8413,In_2937,In_1073);
or U8414 (N_8414,In_2145,In_862);
nand U8415 (N_8415,In_879,In_2153);
or U8416 (N_8416,In_280,In_1595);
and U8417 (N_8417,In_186,In_1314);
and U8418 (N_8418,In_548,In_2847);
nand U8419 (N_8419,In_396,In_984);
and U8420 (N_8420,In_2524,In_1799);
nor U8421 (N_8421,In_1841,In_1853);
nand U8422 (N_8422,In_2713,In_2545);
and U8423 (N_8423,In_2319,In_1358);
nor U8424 (N_8424,In_1392,In_2274);
and U8425 (N_8425,In_1869,In_1497);
or U8426 (N_8426,In_856,In_1591);
or U8427 (N_8427,In_76,In_1538);
and U8428 (N_8428,In_2560,In_2769);
and U8429 (N_8429,In_2169,In_1544);
nor U8430 (N_8430,In_941,In_30);
or U8431 (N_8431,In_1325,In_374);
nand U8432 (N_8432,In_2405,In_2057);
nand U8433 (N_8433,In_2471,In_545);
or U8434 (N_8434,In_1671,In_65);
nand U8435 (N_8435,In_2129,In_541);
nand U8436 (N_8436,In_2724,In_831);
nor U8437 (N_8437,In_2019,In_2924);
nor U8438 (N_8438,In_1504,In_1294);
or U8439 (N_8439,In_1595,In_1455);
nand U8440 (N_8440,In_942,In_2938);
and U8441 (N_8441,In_1995,In_359);
or U8442 (N_8442,In_2503,In_2498);
or U8443 (N_8443,In_629,In_999);
or U8444 (N_8444,In_1920,In_2904);
nor U8445 (N_8445,In_2241,In_1595);
and U8446 (N_8446,In_2939,In_1900);
or U8447 (N_8447,In_2243,In_1363);
nand U8448 (N_8448,In_2707,In_1087);
nor U8449 (N_8449,In_1325,In_23);
nand U8450 (N_8450,In_1101,In_416);
and U8451 (N_8451,In_335,In_49);
and U8452 (N_8452,In_2452,In_1518);
xor U8453 (N_8453,In_1005,In_2778);
and U8454 (N_8454,In_679,In_0);
nor U8455 (N_8455,In_142,In_2049);
nor U8456 (N_8456,In_2629,In_46);
or U8457 (N_8457,In_2261,In_2045);
and U8458 (N_8458,In_173,In_2885);
nand U8459 (N_8459,In_2834,In_1198);
nand U8460 (N_8460,In_1662,In_1710);
or U8461 (N_8461,In_1339,In_1776);
nand U8462 (N_8462,In_2217,In_1388);
or U8463 (N_8463,In_1777,In_1953);
and U8464 (N_8464,In_815,In_2369);
nor U8465 (N_8465,In_2303,In_2795);
nor U8466 (N_8466,In_1335,In_2581);
or U8467 (N_8467,In_26,In_399);
nand U8468 (N_8468,In_2433,In_58);
and U8469 (N_8469,In_2346,In_1489);
or U8470 (N_8470,In_341,In_361);
nor U8471 (N_8471,In_308,In_990);
and U8472 (N_8472,In_1037,In_1113);
nor U8473 (N_8473,In_440,In_2225);
nand U8474 (N_8474,In_1222,In_167);
and U8475 (N_8475,In_785,In_2604);
nor U8476 (N_8476,In_2027,In_1494);
and U8477 (N_8477,In_1102,In_780);
or U8478 (N_8478,In_802,In_348);
nor U8479 (N_8479,In_505,In_1885);
nand U8480 (N_8480,In_180,In_2799);
nand U8481 (N_8481,In_2204,In_2369);
or U8482 (N_8482,In_984,In_2940);
or U8483 (N_8483,In_2149,In_2381);
nor U8484 (N_8484,In_1360,In_337);
nor U8485 (N_8485,In_2338,In_321);
and U8486 (N_8486,In_1010,In_2438);
and U8487 (N_8487,In_1807,In_98);
or U8488 (N_8488,In_2747,In_2821);
nor U8489 (N_8489,In_1004,In_2745);
or U8490 (N_8490,In_2644,In_2726);
and U8491 (N_8491,In_1447,In_560);
or U8492 (N_8492,In_429,In_2381);
nand U8493 (N_8493,In_2994,In_2606);
nor U8494 (N_8494,In_612,In_245);
nand U8495 (N_8495,In_1384,In_344);
and U8496 (N_8496,In_2265,In_1187);
nand U8497 (N_8497,In_1612,In_2992);
nand U8498 (N_8498,In_1860,In_2439);
or U8499 (N_8499,In_2007,In_1797);
nand U8500 (N_8500,In_2226,In_1594);
nand U8501 (N_8501,In_1774,In_1670);
and U8502 (N_8502,In_1965,In_717);
nand U8503 (N_8503,In_1422,In_1485);
or U8504 (N_8504,In_2367,In_2896);
or U8505 (N_8505,In_2507,In_668);
or U8506 (N_8506,In_514,In_1001);
nand U8507 (N_8507,In_650,In_728);
and U8508 (N_8508,In_2609,In_1310);
nand U8509 (N_8509,In_526,In_2850);
nand U8510 (N_8510,In_987,In_1383);
nor U8511 (N_8511,In_951,In_2832);
nand U8512 (N_8512,In_995,In_1954);
or U8513 (N_8513,In_2179,In_2079);
nand U8514 (N_8514,In_1215,In_1919);
nor U8515 (N_8515,In_986,In_2984);
nor U8516 (N_8516,In_685,In_2794);
nor U8517 (N_8517,In_1745,In_389);
and U8518 (N_8518,In_1127,In_2325);
and U8519 (N_8519,In_1767,In_1556);
nand U8520 (N_8520,In_2689,In_542);
or U8521 (N_8521,In_293,In_2532);
and U8522 (N_8522,In_1141,In_2724);
and U8523 (N_8523,In_364,In_765);
or U8524 (N_8524,In_1663,In_877);
and U8525 (N_8525,In_1422,In_384);
and U8526 (N_8526,In_1837,In_2807);
or U8527 (N_8527,In_2140,In_1433);
and U8528 (N_8528,In_599,In_1089);
or U8529 (N_8529,In_2270,In_1845);
and U8530 (N_8530,In_1944,In_1400);
and U8531 (N_8531,In_1457,In_2608);
or U8532 (N_8532,In_1991,In_462);
nor U8533 (N_8533,In_2598,In_1010);
and U8534 (N_8534,In_2105,In_2372);
nor U8535 (N_8535,In_2766,In_2061);
or U8536 (N_8536,In_290,In_2738);
nand U8537 (N_8537,In_2258,In_2403);
and U8538 (N_8538,In_1662,In_1745);
nor U8539 (N_8539,In_2557,In_31);
and U8540 (N_8540,In_2408,In_1367);
nand U8541 (N_8541,In_2596,In_1204);
or U8542 (N_8542,In_966,In_987);
nand U8543 (N_8543,In_2940,In_2012);
and U8544 (N_8544,In_1078,In_240);
nand U8545 (N_8545,In_2116,In_2932);
nor U8546 (N_8546,In_2586,In_2112);
or U8547 (N_8547,In_691,In_1922);
and U8548 (N_8548,In_2738,In_173);
or U8549 (N_8549,In_1261,In_1537);
and U8550 (N_8550,In_2131,In_1523);
and U8551 (N_8551,In_2573,In_2344);
nand U8552 (N_8552,In_2995,In_1261);
nor U8553 (N_8553,In_2089,In_491);
nand U8554 (N_8554,In_1952,In_2168);
or U8555 (N_8555,In_942,In_922);
and U8556 (N_8556,In_2575,In_974);
nor U8557 (N_8557,In_2958,In_2852);
nor U8558 (N_8558,In_2294,In_955);
nand U8559 (N_8559,In_1721,In_1144);
nand U8560 (N_8560,In_1151,In_1737);
or U8561 (N_8561,In_2899,In_588);
nor U8562 (N_8562,In_2811,In_1805);
nand U8563 (N_8563,In_1253,In_2533);
nand U8564 (N_8564,In_267,In_1784);
and U8565 (N_8565,In_2153,In_770);
nand U8566 (N_8566,In_1028,In_202);
nor U8567 (N_8567,In_745,In_1223);
or U8568 (N_8568,In_2582,In_1325);
and U8569 (N_8569,In_779,In_1750);
or U8570 (N_8570,In_706,In_2039);
nand U8571 (N_8571,In_567,In_598);
nor U8572 (N_8572,In_2719,In_2593);
and U8573 (N_8573,In_2043,In_2585);
nand U8574 (N_8574,In_2914,In_2229);
nor U8575 (N_8575,In_447,In_141);
and U8576 (N_8576,In_901,In_2054);
nor U8577 (N_8577,In_869,In_2767);
nor U8578 (N_8578,In_111,In_2035);
and U8579 (N_8579,In_1553,In_1430);
nor U8580 (N_8580,In_2768,In_2209);
or U8581 (N_8581,In_1757,In_2030);
nand U8582 (N_8582,In_986,In_1400);
nor U8583 (N_8583,In_204,In_2327);
and U8584 (N_8584,In_1144,In_1920);
or U8585 (N_8585,In_1865,In_327);
nand U8586 (N_8586,In_2166,In_2956);
or U8587 (N_8587,In_736,In_66);
and U8588 (N_8588,In_1140,In_2824);
and U8589 (N_8589,In_966,In_166);
nor U8590 (N_8590,In_1972,In_133);
and U8591 (N_8591,In_298,In_1499);
nand U8592 (N_8592,In_1458,In_418);
or U8593 (N_8593,In_1600,In_455);
nor U8594 (N_8594,In_1622,In_731);
and U8595 (N_8595,In_2454,In_401);
and U8596 (N_8596,In_2154,In_792);
or U8597 (N_8597,In_2993,In_1161);
or U8598 (N_8598,In_918,In_2178);
and U8599 (N_8599,In_25,In_266);
nand U8600 (N_8600,In_794,In_2628);
or U8601 (N_8601,In_632,In_2999);
or U8602 (N_8602,In_1347,In_120);
and U8603 (N_8603,In_271,In_2363);
xor U8604 (N_8604,In_2704,In_695);
or U8605 (N_8605,In_1923,In_1739);
nor U8606 (N_8606,In_824,In_2741);
nand U8607 (N_8607,In_1796,In_170);
nand U8608 (N_8608,In_1218,In_1028);
nand U8609 (N_8609,In_80,In_126);
nor U8610 (N_8610,In_2991,In_1919);
xor U8611 (N_8611,In_1973,In_1758);
nor U8612 (N_8612,In_467,In_238);
and U8613 (N_8613,In_1435,In_618);
or U8614 (N_8614,In_1678,In_2959);
and U8615 (N_8615,In_1737,In_2039);
or U8616 (N_8616,In_1349,In_1496);
nand U8617 (N_8617,In_893,In_672);
nand U8618 (N_8618,In_2353,In_2866);
nand U8619 (N_8619,In_1862,In_799);
or U8620 (N_8620,In_1460,In_443);
nand U8621 (N_8621,In_2645,In_898);
and U8622 (N_8622,In_193,In_2388);
and U8623 (N_8623,In_784,In_2405);
or U8624 (N_8624,In_2359,In_2815);
or U8625 (N_8625,In_510,In_2449);
nor U8626 (N_8626,In_1421,In_2359);
nand U8627 (N_8627,In_453,In_575);
and U8628 (N_8628,In_1864,In_1599);
nor U8629 (N_8629,In_1757,In_1067);
and U8630 (N_8630,In_1251,In_744);
or U8631 (N_8631,In_2586,In_2696);
nor U8632 (N_8632,In_1937,In_555);
or U8633 (N_8633,In_1136,In_1246);
or U8634 (N_8634,In_1415,In_1864);
or U8635 (N_8635,In_2333,In_432);
or U8636 (N_8636,In_1424,In_637);
and U8637 (N_8637,In_2664,In_1005);
nand U8638 (N_8638,In_2209,In_785);
or U8639 (N_8639,In_831,In_384);
nor U8640 (N_8640,In_420,In_2014);
nand U8641 (N_8641,In_500,In_1085);
or U8642 (N_8642,In_927,In_547);
nor U8643 (N_8643,In_168,In_2591);
nor U8644 (N_8644,In_325,In_1251);
nand U8645 (N_8645,In_422,In_610);
and U8646 (N_8646,In_2889,In_2930);
nand U8647 (N_8647,In_895,In_503);
and U8648 (N_8648,In_2142,In_2083);
nand U8649 (N_8649,In_457,In_1141);
nand U8650 (N_8650,In_1492,In_2361);
nand U8651 (N_8651,In_2562,In_2959);
nor U8652 (N_8652,In_2368,In_1127);
nand U8653 (N_8653,In_2764,In_2144);
nor U8654 (N_8654,In_646,In_2076);
nor U8655 (N_8655,In_1706,In_2361);
nand U8656 (N_8656,In_2140,In_2481);
or U8657 (N_8657,In_1783,In_159);
and U8658 (N_8658,In_916,In_59);
and U8659 (N_8659,In_2960,In_2538);
and U8660 (N_8660,In_910,In_413);
or U8661 (N_8661,In_1087,In_2972);
nor U8662 (N_8662,In_2491,In_1274);
nor U8663 (N_8663,In_840,In_137);
nand U8664 (N_8664,In_2013,In_1294);
or U8665 (N_8665,In_2416,In_544);
nor U8666 (N_8666,In_2085,In_183);
nand U8667 (N_8667,In_1490,In_2403);
and U8668 (N_8668,In_1101,In_2621);
and U8669 (N_8669,In_2054,In_687);
nand U8670 (N_8670,In_507,In_2519);
nand U8671 (N_8671,In_299,In_1744);
and U8672 (N_8672,In_389,In_2892);
and U8673 (N_8673,In_1771,In_1882);
nand U8674 (N_8674,In_100,In_1629);
or U8675 (N_8675,In_2587,In_2795);
nor U8676 (N_8676,In_1380,In_2156);
or U8677 (N_8677,In_1541,In_2837);
nand U8678 (N_8678,In_1809,In_2400);
or U8679 (N_8679,In_639,In_1115);
nand U8680 (N_8680,In_1913,In_1338);
or U8681 (N_8681,In_788,In_2633);
nor U8682 (N_8682,In_1676,In_2733);
nand U8683 (N_8683,In_2298,In_2268);
or U8684 (N_8684,In_1947,In_2604);
nand U8685 (N_8685,In_2447,In_2394);
and U8686 (N_8686,In_1195,In_1878);
nor U8687 (N_8687,In_2865,In_452);
or U8688 (N_8688,In_1062,In_1310);
or U8689 (N_8689,In_990,In_1693);
nor U8690 (N_8690,In_2787,In_604);
and U8691 (N_8691,In_1231,In_2822);
nand U8692 (N_8692,In_609,In_831);
nand U8693 (N_8693,In_1932,In_2979);
nor U8694 (N_8694,In_773,In_2190);
or U8695 (N_8695,In_867,In_1204);
nand U8696 (N_8696,In_2361,In_2635);
or U8697 (N_8697,In_2226,In_174);
xor U8698 (N_8698,In_1271,In_966);
nor U8699 (N_8699,In_2839,In_2804);
and U8700 (N_8700,In_2508,In_1498);
or U8701 (N_8701,In_1804,In_1786);
nor U8702 (N_8702,In_1376,In_399);
or U8703 (N_8703,In_2703,In_1264);
and U8704 (N_8704,In_1715,In_2487);
and U8705 (N_8705,In_335,In_1363);
or U8706 (N_8706,In_1557,In_1812);
and U8707 (N_8707,In_437,In_2616);
or U8708 (N_8708,In_786,In_2577);
or U8709 (N_8709,In_1815,In_2925);
nor U8710 (N_8710,In_2510,In_1843);
nor U8711 (N_8711,In_798,In_2644);
and U8712 (N_8712,In_2761,In_228);
nor U8713 (N_8713,In_826,In_686);
nor U8714 (N_8714,In_2535,In_744);
and U8715 (N_8715,In_1185,In_2747);
nor U8716 (N_8716,In_123,In_929);
nand U8717 (N_8717,In_1815,In_930);
nand U8718 (N_8718,In_1442,In_468);
and U8719 (N_8719,In_263,In_570);
nor U8720 (N_8720,In_2398,In_1360);
nand U8721 (N_8721,In_1115,In_2621);
nor U8722 (N_8722,In_1466,In_2090);
nor U8723 (N_8723,In_1001,In_154);
nor U8724 (N_8724,In_319,In_297);
or U8725 (N_8725,In_2917,In_475);
or U8726 (N_8726,In_968,In_1653);
or U8727 (N_8727,In_2209,In_124);
nor U8728 (N_8728,In_2947,In_2031);
nand U8729 (N_8729,In_1109,In_718);
nand U8730 (N_8730,In_1903,In_344);
or U8731 (N_8731,In_2106,In_453);
or U8732 (N_8732,In_363,In_189);
nand U8733 (N_8733,In_1440,In_629);
and U8734 (N_8734,In_1072,In_1753);
nand U8735 (N_8735,In_2607,In_1384);
or U8736 (N_8736,In_2039,In_1313);
nor U8737 (N_8737,In_2852,In_2211);
and U8738 (N_8738,In_2361,In_526);
and U8739 (N_8739,In_1317,In_132);
or U8740 (N_8740,In_2665,In_1297);
nand U8741 (N_8741,In_1804,In_0);
or U8742 (N_8742,In_1280,In_2035);
or U8743 (N_8743,In_2521,In_1276);
nand U8744 (N_8744,In_114,In_649);
or U8745 (N_8745,In_2722,In_46);
nand U8746 (N_8746,In_143,In_660);
nor U8747 (N_8747,In_98,In_210);
or U8748 (N_8748,In_1564,In_1704);
nand U8749 (N_8749,In_595,In_2210);
and U8750 (N_8750,In_1455,In_754);
nand U8751 (N_8751,In_2554,In_487);
or U8752 (N_8752,In_1958,In_2808);
or U8753 (N_8753,In_2997,In_1576);
nand U8754 (N_8754,In_2359,In_239);
or U8755 (N_8755,In_249,In_29);
and U8756 (N_8756,In_669,In_379);
and U8757 (N_8757,In_1161,In_1145);
nand U8758 (N_8758,In_387,In_744);
or U8759 (N_8759,In_1975,In_2836);
nand U8760 (N_8760,In_2423,In_1450);
and U8761 (N_8761,In_354,In_1467);
or U8762 (N_8762,In_2386,In_630);
and U8763 (N_8763,In_141,In_492);
and U8764 (N_8764,In_1932,In_1767);
or U8765 (N_8765,In_1823,In_1955);
nor U8766 (N_8766,In_95,In_2095);
and U8767 (N_8767,In_409,In_1805);
or U8768 (N_8768,In_2556,In_1860);
nand U8769 (N_8769,In_1389,In_1722);
and U8770 (N_8770,In_1621,In_1561);
nand U8771 (N_8771,In_46,In_1440);
nor U8772 (N_8772,In_1581,In_2158);
nand U8773 (N_8773,In_632,In_686);
nand U8774 (N_8774,In_2202,In_1929);
nor U8775 (N_8775,In_2130,In_2755);
and U8776 (N_8776,In_1714,In_1831);
or U8777 (N_8777,In_2444,In_1647);
nor U8778 (N_8778,In_1782,In_2332);
nand U8779 (N_8779,In_741,In_138);
nor U8780 (N_8780,In_1780,In_2099);
and U8781 (N_8781,In_402,In_2384);
nor U8782 (N_8782,In_1846,In_2722);
and U8783 (N_8783,In_2429,In_1546);
xor U8784 (N_8784,In_429,In_990);
nand U8785 (N_8785,In_199,In_213);
nor U8786 (N_8786,In_2354,In_1701);
nor U8787 (N_8787,In_417,In_710);
and U8788 (N_8788,In_1136,In_19);
nand U8789 (N_8789,In_2088,In_2039);
or U8790 (N_8790,In_1508,In_638);
nor U8791 (N_8791,In_1328,In_1884);
nand U8792 (N_8792,In_2143,In_71);
or U8793 (N_8793,In_455,In_863);
nand U8794 (N_8794,In_1681,In_445);
nand U8795 (N_8795,In_2590,In_1072);
or U8796 (N_8796,In_1441,In_905);
or U8797 (N_8797,In_1015,In_572);
or U8798 (N_8798,In_1145,In_722);
nand U8799 (N_8799,In_2607,In_2453);
nand U8800 (N_8800,In_1433,In_102);
or U8801 (N_8801,In_1899,In_435);
nor U8802 (N_8802,In_2408,In_1242);
or U8803 (N_8803,In_1781,In_2253);
nand U8804 (N_8804,In_2776,In_6);
nor U8805 (N_8805,In_2307,In_2704);
nand U8806 (N_8806,In_1206,In_2017);
xor U8807 (N_8807,In_1642,In_1973);
and U8808 (N_8808,In_2788,In_1229);
or U8809 (N_8809,In_370,In_754);
and U8810 (N_8810,In_1762,In_85);
and U8811 (N_8811,In_130,In_2241);
or U8812 (N_8812,In_198,In_2296);
and U8813 (N_8813,In_1526,In_445);
nand U8814 (N_8814,In_453,In_1871);
and U8815 (N_8815,In_1028,In_1985);
nor U8816 (N_8816,In_1502,In_2389);
nor U8817 (N_8817,In_1278,In_1662);
or U8818 (N_8818,In_1751,In_2926);
or U8819 (N_8819,In_2387,In_96);
nand U8820 (N_8820,In_1962,In_763);
and U8821 (N_8821,In_1650,In_2528);
nand U8822 (N_8822,In_2595,In_114);
nor U8823 (N_8823,In_649,In_1337);
nor U8824 (N_8824,In_25,In_824);
nor U8825 (N_8825,In_911,In_987);
nor U8826 (N_8826,In_1851,In_674);
and U8827 (N_8827,In_2033,In_447);
and U8828 (N_8828,In_1000,In_2983);
or U8829 (N_8829,In_1837,In_269);
and U8830 (N_8830,In_1939,In_310);
and U8831 (N_8831,In_111,In_2642);
or U8832 (N_8832,In_1719,In_2348);
nor U8833 (N_8833,In_435,In_108);
nor U8834 (N_8834,In_2264,In_25);
nor U8835 (N_8835,In_1390,In_953);
nand U8836 (N_8836,In_925,In_1346);
and U8837 (N_8837,In_2770,In_2107);
nor U8838 (N_8838,In_1617,In_2953);
and U8839 (N_8839,In_1113,In_2809);
nand U8840 (N_8840,In_2331,In_275);
and U8841 (N_8841,In_2199,In_1530);
nand U8842 (N_8842,In_1459,In_128);
nor U8843 (N_8843,In_2684,In_1930);
and U8844 (N_8844,In_2516,In_2943);
and U8845 (N_8845,In_1314,In_1291);
or U8846 (N_8846,In_770,In_179);
and U8847 (N_8847,In_760,In_1883);
and U8848 (N_8848,In_982,In_1420);
or U8849 (N_8849,In_256,In_965);
nor U8850 (N_8850,In_1182,In_2406);
or U8851 (N_8851,In_458,In_582);
and U8852 (N_8852,In_2717,In_231);
or U8853 (N_8853,In_2096,In_29);
nand U8854 (N_8854,In_1332,In_2003);
and U8855 (N_8855,In_1647,In_970);
and U8856 (N_8856,In_2027,In_2212);
and U8857 (N_8857,In_1875,In_860);
and U8858 (N_8858,In_1238,In_1230);
and U8859 (N_8859,In_304,In_2703);
nor U8860 (N_8860,In_602,In_138);
nand U8861 (N_8861,In_396,In_1514);
nor U8862 (N_8862,In_1978,In_578);
or U8863 (N_8863,In_1406,In_830);
and U8864 (N_8864,In_963,In_1037);
nand U8865 (N_8865,In_388,In_2851);
and U8866 (N_8866,In_1502,In_2232);
and U8867 (N_8867,In_2144,In_2321);
nand U8868 (N_8868,In_92,In_2627);
or U8869 (N_8869,In_2556,In_1175);
nand U8870 (N_8870,In_686,In_2250);
xnor U8871 (N_8871,In_2741,In_303);
nor U8872 (N_8872,In_2409,In_1194);
nor U8873 (N_8873,In_2626,In_1060);
or U8874 (N_8874,In_1199,In_1818);
and U8875 (N_8875,In_310,In_443);
nand U8876 (N_8876,In_1650,In_966);
nor U8877 (N_8877,In_2918,In_707);
nor U8878 (N_8878,In_371,In_1442);
and U8879 (N_8879,In_937,In_2212);
and U8880 (N_8880,In_527,In_1399);
nor U8881 (N_8881,In_2519,In_1539);
nand U8882 (N_8882,In_1479,In_2070);
or U8883 (N_8883,In_1767,In_937);
or U8884 (N_8884,In_855,In_2982);
nor U8885 (N_8885,In_1226,In_2814);
nor U8886 (N_8886,In_1264,In_1380);
nand U8887 (N_8887,In_1174,In_2803);
nand U8888 (N_8888,In_1132,In_1120);
nand U8889 (N_8889,In_34,In_2534);
or U8890 (N_8890,In_2218,In_748);
and U8891 (N_8891,In_1940,In_1291);
nor U8892 (N_8892,In_2130,In_1453);
and U8893 (N_8893,In_1708,In_418);
or U8894 (N_8894,In_1585,In_917);
nand U8895 (N_8895,In_260,In_734);
nor U8896 (N_8896,In_1372,In_2828);
or U8897 (N_8897,In_2159,In_2183);
nor U8898 (N_8898,In_2415,In_1124);
nand U8899 (N_8899,In_666,In_1519);
and U8900 (N_8900,In_589,In_829);
nor U8901 (N_8901,In_1841,In_1647);
and U8902 (N_8902,In_2970,In_1769);
nor U8903 (N_8903,In_1885,In_2354);
and U8904 (N_8904,In_2106,In_690);
and U8905 (N_8905,In_822,In_1056);
and U8906 (N_8906,In_394,In_1321);
nor U8907 (N_8907,In_2419,In_1618);
nor U8908 (N_8908,In_1980,In_623);
nand U8909 (N_8909,In_1952,In_2188);
nand U8910 (N_8910,In_2940,In_926);
or U8911 (N_8911,In_849,In_1869);
nand U8912 (N_8912,In_1507,In_1577);
nand U8913 (N_8913,In_2208,In_2385);
nor U8914 (N_8914,In_1639,In_1492);
or U8915 (N_8915,In_1092,In_1602);
or U8916 (N_8916,In_1821,In_234);
nand U8917 (N_8917,In_1196,In_933);
or U8918 (N_8918,In_690,In_1171);
nor U8919 (N_8919,In_2187,In_1748);
nor U8920 (N_8920,In_200,In_1285);
and U8921 (N_8921,In_2279,In_2633);
nor U8922 (N_8922,In_2724,In_1126);
nand U8923 (N_8923,In_1606,In_2967);
nand U8924 (N_8924,In_497,In_2894);
or U8925 (N_8925,In_1081,In_1864);
nand U8926 (N_8926,In_2376,In_267);
nand U8927 (N_8927,In_763,In_519);
nor U8928 (N_8928,In_2149,In_1409);
nand U8929 (N_8929,In_2942,In_2975);
or U8930 (N_8930,In_658,In_1381);
nor U8931 (N_8931,In_2810,In_2907);
or U8932 (N_8932,In_2712,In_1352);
nand U8933 (N_8933,In_2677,In_1112);
or U8934 (N_8934,In_338,In_267);
and U8935 (N_8935,In_353,In_2785);
nand U8936 (N_8936,In_2972,In_423);
nor U8937 (N_8937,In_796,In_623);
nor U8938 (N_8938,In_1476,In_2314);
and U8939 (N_8939,In_734,In_2839);
nand U8940 (N_8940,In_526,In_1564);
nor U8941 (N_8941,In_331,In_2832);
or U8942 (N_8942,In_1384,In_1506);
nand U8943 (N_8943,In_2735,In_2527);
or U8944 (N_8944,In_2680,In_454);
nor U8945 (N_8945,In_2097,In_1264);
nor U8946 (N_8946,In_2938,In_472);
and U8947 (N_8947,In_845,In_2530);
and U8948 (N_8948,In_801,In_2713);
nor U8949 (N_8949,In_141,In_2080);
nor U8950 (N_8950,In_1528,In_2791);
and U8951 (N_8951,In_923,In_1335);
and U8952 (N_8952,In_1763,In_1818);
nand U8953 (N_8953,In_641,In_1302);
or U8954 (N_8954,In_2839,In_285);
nor U8955 (N_8955,In_2736,In_1823);
and U8956 (N_8956,In_1641,In_1177);
nor U8957 (N_8957,In_1841,In_1673);
nor U8958 (N_8958,In_2364,In_2367);
nor U8959 (N_8959,In_1948,In_1524);
nor U8960 (N_8960,In_1837,In_452);
nor U8961 (N_8961,In_2403,In_207);
nor U8962 (N_8962,In_1663,In_2904);
nand U8963 (N_8963,In_2593,In_2916);
nand U8964 (N_8964,In_332,In_2675);
and U8965 (N_8965,In_1829,In_82);
nor U8966 (N_8966,In_1817,In_515);
nor U8967 (N_8967,In_2667,In_2469);
or U8968 (N_8968,In_2872,In_481);
nor U8969 (N_8969,In_332,In_1354);
or U8970 (N_8970,In_1897,In_1675);
nor U8971 (N_8971,In_559,In_479);
nand U8972 (N_8972,In_2574,In_2500);
and U8973 (N_8973,In_1959,In_1659);
and U8974 (N_8974,In_1815,In_2841);
and U8975 (N_8975,In_940,In_2782);
or U8976 (N_8976,In_26,In_1638);
or U8977 (N_8977,In_2093,In_2291);
nor U8978 (N_8978,In_2222,In_1477);
nand U8979 (N_8979,In_530,In_2515);
nor U8980 (N_8980,In_1263,In_551);
nand U8981 (N_8981,In_1537,In_1831);
or U8982 (N_8982,In_2384,In_1613);
nand U8983 (N_8983,In_2020,In_233);
and U8984 (N_8984,In_1894,In_404);
and U8985 (N_8985,In_887,In_591);
or U8986 (N_8986,In_197,In_1957);
nor U8987 (N_8987,In_2773,In_2179);
nand U8988 (N_8988,In_2794,In_1455);
nand U8989 (N_8989,In_1564,In_256);
nor U8990 (N_8990,In_2710,In_1417);
nand U8991 (N_8991,In_53,In_1722);
xnor U8992 (N_8992,In_1272,In_532);
or U8993 (N_8993,In_1823,In_93);
nor U8994 (N_8994,In_2935,In_1813);
nor U8995 (N_8995,In_648,In_2849);
and U8996 (N_8996,In_1158,In_1106);
and U8997 (N_8997,In_2071,In_1602);
and U8998 (N_8998,In_1740,In_2461);
nand U8999 (N_8999,In_1285,In_632);
nor U9000 (N_9000,In_508,In_376);
or U9001 (N_9001,In_1002,In_1700);
nand U9002 (N_9002,In_2570,In_1238);
or U9003 (N_9003,In_1939,In_399);
and U9004 (N_9004,In_156,In_2302);
and U9005 (N_9005,In_955,In_2228);
and U9006 (N_9006,In_1643,In_773);
or U9007 (N_9007,In_207,In_327);
and U9008 (N_9008,In_2620,In_2564);
nor U9009 (N_9009,In_2835,In_873);
and U9010 (N_9010,In_2573,In_2123);
nand U9011 (N_9011,In_2994,In_349);
and U9012 (N_9012,In_2756,In_2751);
nor U9013 (N_9013,In_1555,In_460);
nor U9014 (N_9014,In_2454,In_1093);
nor U9015 (N_9015,In_1673,In_1574);
nand U9016 (N_9016,In_879,In_1731);
nor U9017 (N_9017,In_718,In_478);
nor U9018 (N_9018,In_2083,In_1917);
and U9019 (N_9019,In_2958,In_2917);
nand U9020 (N_9020,In_1038,In_1384);
or U9021 (N_9021,In_1675,In_820);
nand U9022 (N_9022,In_372,In_1798);
or U9023 (N_9023,In_783,In_1539);
and U9024 (N_9024,In_2676,In_2807);
or U9025 (N_9025,In_518,In_589);
xnor U9026 (N_9026,In_2595,In_2178);
nand U9027 (N_9027,In_1707,In_881);
or U9028 (N_9028,In_2937,In_1737);
xnor U9029 (N_9029,In_2050,In_1152);
nor U9030 (N_9030,In_834,In_2490);
and U9031 (N_9031,In_2512,In_1700);
nand U9032 (N_9032,In_884,In_1415);
or U9033 (N_9033,In_2982,In_2709);
and U9034 (N_9034,In_1228,In_2129);
nor U9035 (N_9035,In_731,In_53);
nor U9036 (N_9036,In_1839,In_1489);
nor U9037 (N_9037,In_1440,In_660);
nor U9038 (N_9038,In_1596,In_1745);
and U9039 (N_9039,In_926,In_902);
or U9040 (N_9040,In_2743,In_1070);
nor U9041 (N_9041,In_2074,In_2660);
and U9042 (N_9042,In_625,In_2290);
or U9043 (N_9043,In_1365,In_1443);
and U9044 (N_9044,In_1167,In_1161);
nor U9045 (N_9045,In_2345,In_942);
nand U9046 (N_9046,In_1389,In_2587);
nor U9047 (N_9047,In_2638,In_439);
xnor U9048 (N_9048,In_176,In_527);
nand U9049 (N_9049,In_329,In_428);
nor U9050 (N_9050,In_2720,In_1339);
nand U9051 (N_9051,In_239,In_2174);
or U9052 (N_9052,In_801,In_387);
nand U9053 (N_9053,In_201,In_1067);
or U9054 (N_9054,In_2925,In_2674);
nand U9055 (N_9055,In_1253,In_1315);
and U9056 (N_9056,In_1256,In_1536);
nor U9057 (N_9057,In_593,In_1318);
and U9058 (N_9058,In_1851,In_1385);
or U9059 (N_9059,In_2287,In_2334);
and U9060 (N_9060,In_2962,In_944);
or U9061 (N_9061,In_2665,In_1056);
or U9062 (N_9062,In_1183,In_2893);
nor U9063 (N_9063,In_1272,In_514);
or U9064 (N_9064,In_1575,In_279);
and U9065 (N_9065,In_1409,In_70);
or U9066 (N_9066,In_2220,In_714);
nor U9067 (N_9067,In_2447,In_1963);
or U9068 (N_9068,In_111,In_1807);
nand U9069 (N_9069,In_1083,In_1166);
xor U9070 (N_9070,In_2021,In_2648);
nand U9071 (N_9071,In_2884,In_4);
nand U9072 (N_9072,In_2832,In_580);
or U9073 (N_9073,In_2584,In_68);
or U9074 (N_9074,In_18,In_1827);
nand U9075 (N_9075,In_861,In_1099);
and U9076 (N_9076,In_1289,In_2023);
or U9077 (N_9077,In_2454,In_141);
or U9078 (N_9078,In_688,In_386);
and U9079 (N_9079,In_1684,In_1541);
nand U9080 (N_9080,In_2342,In_76);
nand U9081 (N_9081,In_1772,In_41);
or U9082 (N_9082,In_1011,In_2651);
nand U9083 (N_9083,In_569,In_1155);
or U9084 (N_9084,In_1714,In_2353);
and U9085 (N_9085,In_1583,In_1665);
or U9086 (N_9086,In_2562,In_1911);
or U9087 (N_9087,In_1416,In_1639);
or U9088 (N_9088,In_2887,In_1328);
or U9089 (N_9089,In_146,In_1751);
or U9090 (N_9090,In_2326,In_822);
and U9091 (N_9091,In_1061,In_2208);
nor U9092 (N_9092,In_2388,In_1627);
nand U9093 (N_9093,In_2188,In_1043);
nor U9094 (N_9094,In_1476,In_246);
and U9095 (N_9095,In_1216,In_2629);
and U9096 (N_9096,In_320,In_1085);
and U9097 (N_9097,In_1303,In_310);
and U9098 (N_9098,In_827,In_750);
nand U9099 (N_9099,In_1271,In_2197);
or U9100 (N_9100,In_1133,In_1399);
or U9101 (N_9101,In_66,In_1108);
and U9102 (N_9102,In_1598,In_2659);
and U9103 (N_9103,In_2173,In_2243);
or U9104 (N_9104,In_2584,In_430);
nor U9105 (N_9105,In_2064,In_2117);
nor U9106 (N_9106,In_2893,In_893);
nand U9107 (N_9107,In_640,In_1494);
nand U9108 (N_9108,In_1133,In_1624);
nor U9109 (N_9109,In_2080,In_807);
and U9110 (N_9110,In_1851,In_2824);
nor U9111 (N_9111,In_424,In_813);
nor U9112 (N_9112,In_941,In_1286);
nand U9113 (N_9113,In_1503,In_1455);
or U9114 (N_9114,In_2761,In_852);
nor U9115 (N_9115,In_1641,In_283);
nor U9116 (N_9116,In_2388,In_2907);
or U9117 (N_9117,In_339,In_1837);
and U9118 (N_9118,In_2631,In_1915);
nor U9119 (N_9119,In_2762,In_2279);
or U9120 (N_9120,In_953,In_615);
and U9121 (N_9121,In_810,In_1610);
nor U9122 (N_9122,In_2282,In_1302);
nand U9123 (N_9123,In_470,In_398);
nand U9124 (N_9124,In_601,In_617);
or U9125 (N_9125,In_1629,In_2649);
or U9126 (N_9126,In_1625,In_83);
or U9127 (N_9127,In_2794,In_273);
and U9128 (N_9128,In_1838,In_1193);
nor U9129 (N_9129,In_732,In_2045);
nand U9130 (N_9130,In_2535,In_1155);
and U9131 (N_9131,In_2924,In_2432);
and U9132 (N_9132,In_740,In_2185);
nor U9133 (N_9133,In_2768,In_1311);
and U9134 (N_9134,In_2232,In_144);
or U9135 (N_9135,In_342,In_2887);
or U9136 (N_9136,In_2933,In_380);
and U9137 (N_9137,In_711,In_839);
or U9138 (N_9138,In_1952,In_359);
or U9139 (N_9139,In_2730,In_137);
nand U9140 (N_9140,In_7,In_1427);
or U9141 (N_9141,In_1264,In_2711);
or U9142 (N_9142,In_1683,In_362);
and U9143 (N_9143,In_1454,In_1380);
xnor U9144 (N_9144,In_2143,In_534);
nor U9145 (N_9145,In_905,In_1769);
or U9146 (N_9146,In_939,In_1228);
nor U9147 (N_9147,In_721,In_1599);
nor U9148 (N_9148,In_889,In_2173);
or U9149 (N_9149,In_1744,In_2573);
and U9150 (N_9150,In_266,In_1534);
or U9151 (N_9151,In_2101,In_1947);
and U9152 (N_9152,In_2439,In_91);
and U9153 (N_9153,In_1323,In_512);
nor U9154 (N_9154,In_1328,In_2529);
nor U9155 (N_9155,In_328,In_1815);
and U9156 (N_9156,In_1625,In_2985);
nand U9157 (N_9157,In_1882,In_1520);
nand U9158 (N_9158,In_953,In_1511);
or U9159 (N_9159,In_1369,In_2242);
nand U9160 (N_9160,In_2792,In_2302);
nor U9161 (N_9161,In_2487,In_1368);
nand U9162 (N_9162,In_848,In_2639);
and U9163 (N_9163,In_925,In_2604);
and U9164 (N_9164,In_1323,In_2599);
and U9165 (N_9165,In_164,In_2821);
or U9166 (N_9166,In_1756,In_943);
and U9167 (N_9167,In_344,In_60);
or U9168 (N_9168,In_1211,In_1966);
or U9169 (N_9169,In_573,In_1033);
nand U9170 (N_9170,In_2137,In_1193);
nand U9171 (N_9171,In_691,In_178);
nor U9172 (N_9172,In_2600,In_463);
and U9173 (N_9173,In_498,In_2149);
or U9174 (N_9174,In_1321,In_507);
or U9175 (N_9175,In_2191,In_1972);
nor U9176 (N_9176,In_1905,In_2091);
nand U9177 (N_9177,In_1808,In_2869);
and U9178 (N_9178,In_1051,In_574);
and U9179 (N_9179,In_195,In_1070);
or U9180 (N_9180,In_2154,In_1525);
nand U9181 (N_9181,In_2715,In_1468);
xor U9182 (N_9182,In_89,In_878);
and U9183 (N_9183,In_2607,In_2005);
nand U9184 (N_9184,In_980,In_1821);
nand U9185 (N_9185,In_2191,In_619);
nor U9186 (N_9186,In_2494,In_710);
and U9187 (N_9187,In_2048,In_842);
or U9188 (N_9188,In_1598,In_343);
or U9189 (N_9189,In_1774,In_2071);
nor U9190 (N_9190,In_828,In_2136);
or U9191 (N_9191,In_2862,In_2185);
nand U9192 (N_9192,In_905,In_2710);
nand U9193 (N_9193,In_2280,In_2531);
xor U9194 (N_9194,In_2146,In_1515);
and U9195 (N_9195,In_102,In_1294);
nand U9196 (N_9196,In_1432,In_1498);
nor U9197 (N_9197,In_144,In_1232);
or U9198 (N_9198,In_2897,In_656);
and U9199 (N_9199,In_664,In_739);
and U9200 (N_9200,In_2636,In_1515);
and U9201 (N_9201,In_2294,In_952);
and U9202 (N_9202,In_67,In_166);
or U9203 (N_9203,In_2956,In_1066);
and U9204 (N_9204,In_1808,In_2529);
or U9205 (N_9205,In_306,In_2610);
nand U9206 (N_9206,In_2983,In_1588);
nand U9207 (N_9207,In_1500,In_982);
nor U9208 (N_9208,In_238,In_815);
nor U9209 (N_9209,In_407,In_224);
and U9210 (N_9210,In_1084,In_1713);
or U9211 (N_9211,In_1394,In_1405);
and U9212 (N_9212,In_1557,In_305);
nor U9213 (N_9213,In_1793,In_1711);
nor U9214 (N_9214,In_2144,In_2463);
nor U9215 (N_9215,In_2773,In_1023);
or U9216 (N_9216,In_1159,In_2763);
or U9217 (N_9217,In_469,In_691);
nand U9218 (N_9218,In_225,In_2572);
nor U9219 (N_9219,In_2715,In_423);
and U9220 (N_9220,In_1744,In_1842);
nor U9221 (N_9221,In_1276,In_988);
nand U9222 (N_9222,In_2297,In_1542);
nor U9223 (N_9223,In_2444,In_1060);
or U9224 (N_9224,In_1977,In_2541);
and U9225 (N_9225,In_2496,In_1031);
nor U9226 (N_9226,In_2691,In_232);
nor U9227 (N_9227,In_678,In_2875);
nand U9228 (N_9228,In_1847,In_1019);
nand U9229 (N_9229,In_584,In_2941);
or U9230 (N_9230,In_2731,In_1471);
or U9231 (N_9231,In_473,In_2578);
and U9232 (N_9232,In_1028,In_219);
nor U9233 (N_9233,In_2846,In_2777);
nand U9234 (N_9234,In_2416,In_1905);
nand U9235 (N_9235,In_2316,In_656);
or U9236 (N_9236,In_2047,In_1504);
nor U9237 (N_9237,In_307,In_1951);
and U9238 (N_9238,In_77,In_1259);
or U9239 (N_9239,In_2248,In_1699);
or U9240 (N_9240,In_2926,In_2411);
nor U9241 (N_9241,In_1579,In_955);
nor U9242 (N_9242,In_1241,In_2386);
nor U9243 (N_9243,In_1989,In_807);
nand U9244 (N_9244,In_2810,In_1020);
nor U9245 (N_9245,In_771,In_1815);
nor U9246 (N_9246,In_709,In_2661);
or U9247 (N_9247,In_1841,In_1206);
nor U9248 (N_9248,In_41,In_2497);
and U9249 (N_9249,In_1989,In_1006);
nand U9250 (N_9250,In_2307,In_1431);
or U9251 (N_9251,In_2037,In_1933);
or U9252 (N_9252,In_2538,In_477);
or U9253 (N_9253,In_603,In_2317);
and U9254 (N_9254,In_2493,In_1991);
and U9255 (N_9255,In_2968,In_739);
or U9256 (N_9256,In_917,In_1875);
or U9257 (N_9257,In_710,In_1954);
or U9258 (N_9258,In_2519,In_1455);
nand U9259 (N_9259,In_409,In_591);
and U9260 (N_9260,In_1484,In_2449);
and U9261 (N_9261,In_2141,In_2487);
and U9262 (N_9262,In_1761,In_1699);
nand U9263 (N_9263,In_2110,In_1464);
nand U9264 (N_9264,In_182,In_1252);
and U9265 (N_9265,In_1346,In_653);
nor U9266 (N_9266,In_1786,In_1776);
and U9267 (N_9267,In_1198,In_708);
and U9268 (N_9268,In_2909,In_683);
nand U9269 (N_9269,In_970,In_2712);
and U9270 (N_9270,In_2677,In_2044);
and U9271 (N_9271,In_1852,In_1289);
nor U9272 (N_9272,In_2632,In_2799);
or U9273 (N_9273,In_1745,In_1736);
nand U9274 (N_9274,In_146,In_1314);
nand U9275 (N_9275,In_2862,In_626);
and U9276 (N_9276,In_2421,In_1373);
or U9277 (N_9277,In_1916,In_1193);
nor U9278 (N_9278,In_1223,In_679);
and U9279 (N_9279,In_23,In_939);
nand U9280 (N_9280,In_2020,In_1256);
nand U9281 (N_9281,In_2093,In_966);
or U9282 (N_9282,In_2210,In_2786);
nand U9283 (N_9283,In_2716,In_2354);
nor U9284 (N_9284,In_2181,In_898);
nand U9285 (N_9285,In_2182,In_1265);
nand U9286 (N_9286,In_538,In_2205);
nor U9287 (N_9287,In_1189,In_655);
or U9288 (N_9288,In_2394,In_2030);
and U9289 (N_9289,In_1813,In_2368);
and U9290 (N_9290,In_430,In_155);
nor U9291 (N_9291,In_321,In_119);
or U9292 (N_9292,In_2908,In_450);
or U9293 (N_9293,In_1458,In_2062);
nand U9294 (N_9294,In_16,In_2658);
nor U9295 (N_9295,In_2864,In_2872);
or U9296 (N_9296,In_1440,In_2047);
or U9297 (N_9297,In_1638,In_251);
nand U9298 (N_9298,In_1232,In_1079);
and U9299 (N_9299,In_745,In_158);
and U9300 (N_9300,In_1524,In_1353);
or U9301 (N_9301,In_1385,In_279);
nor U9302 (N_9302,In_2055,In_386);
and U9303 (N_9303,In_1518,In_1887);
nand U9304 (N_9304,In_1030,In_148);
nor U9305 (N_9305,In_1436,In_1215);
nand U9306 (N_9306,In_489,In_2232);
nand U9307 (N_9307,In_1066,In_698);
or U9308 (N_9308,In_1676,In_47);
or U9309 (N_9309,In_1793,In_1859);
or U9310 (N_9310,In_1108,In_1985);
nand U9311 (N_9311,In_2902,In_2624);
nand U9312 (N_9312,In_1781,In_431);
and U9313 (N_9313,In_2493,In_434);
and U9314 (N_9314,In_1665,In_2487);
or U9315 (N_9315,In_1264,In_1942);
and U9316 (N_9316,In_1251,In_2607);
nor U9317 (N_9317,In_415,In_2838);
nand U9318 (N_9318,In_2315,In_463);
nor U9319 (N_9319,In_2155,In_2680);
nand U9320 (N_9320,In_5,In_807);
nor U9321 (N_9321,In_1770,In_280);
and U9322 (N_9322,In_206,In_1551);
nand U9323 (N_9323,In_1629,In_748);
nor U9324 (N_9324,In_315,In_924);
or U9325 (N_9325,In_2372,In_2462);
or U9326 (N_9326,In_1461,In_354);
and U9327 (N_9327,In_1660,In_2684);
nand U9328 (N_9328,In_1946,In_2707);
and U9329 (N_9329,In_418,In_1873);
nor U9330 (N_9330,In_1300,In_1638);
nor U9331 (N_9331,In_2832,In_2568);
or U9332 (N_9332,In_1334,In_1860);
or U9333 (N_9333,In_1513,In_479);
nand U9334 (N_9334,In_935,In_1566);
xnor U9335 (N_9335,In_2015,In_7);
and U9336 (N_9336,In_2199,In_2586);
nor U9337 (N_9337,In_2036,In_87);
nor U9338 (N_9338,In_1451,In_1293);
nor U9339 (N_9339,In_2325,In_2990);
and U9340 (N_9340,In_213,In_1073);
nand U9341 (N_9341,In_1764,In_79);
and U9342 (N_9342,In_470,In_894);
nor U9343 (N_9343,In_1102,In_1648);
and U9344 (N_9344,In_1658,In_222);
or U9345 (N_9345,In_626,In_2193);
nand U9346 (N_9346,In_316,In_2314);
or U9347 (N_9347,In_702,In_512);
nand U9348 (N_9348,In_864,In_2526);
nand U9349 (N_9349,In_430,In_42);
nand U9350 (N_9350,In_2134,In_2098);
nor U9351 (N_9351,In_1861,In_2946);
nor U9352 (N_9352,In_564,In_1558);
nand U9353 (N_9353,In_2517,In_475);
nor U9354 (N_9354,In_2387,In_2524);
and U9355 (N_9355,In_980,In_1506);
or U9356 (N_9356,In_2356,In_628);
and U9357 (N_9357,In_2752,In_2079);
nor U9358 (N_9358,In_2593,In_297);
nor U9359 (N_9359,In_61,In_1408);
or U9360 (N_9360,In_2418,In_590);
nor U9361 (N_9361,In_2214,In_2518);
nand U9362 (N_9362,In_650,In_2800);
or U9363 (N_9363,In_2695,In_2154);
nor U9364 (N_9364,In_1124,In_1452);
nand U9365 (N_9365,In_725,In_2348);
nor U9366 (N_9366,In_866,In_2825);
or U9367 (N_9367,In_1555,In_165);
or U9368 (N_9368,In_403,In_86);
or U9369 (N_9369,In_1253,In_2003);
or U9370 (N_9370,In_1125,In_1520);
or U9371 (N_9371,In_1774,In_367);
and U9372 (N_9372,In_1399,In_1812);
or U9373 (N_9373,In_427,In_738);
nor U9374 (N_9374,In_751,In_849);
and U9375 (N_9375,In_595,In_2235);
nand U9376 (N_9376,In_2476,In_1601);
nand U9377 (N_9377,In_43,In_1913);
nand U9378 (N_9378,In_2186,In_930);
and U9379 (N_9379,In_1366,In_2511);
or U9380 (N_9380,In_2255,In_1670);
and U9381 (N_9381,In_112,In_2000);
and U9382 (N_9382,In_1083,In_2940);
nand U9383 (N_9383,In_347,In_598);
nand U9384 (N_9384,In_2999,In_69);
and U9385 (N_9385,In_2796,In_6);
nand U9386 (N_9386,In_2501,In_758);
nand U9387 (N_9387,In_2320,In_2323);
nor U9388 (N_9388,In_2798,In_1055);
nand U9389 (N_9389,In_642,In_1535);
nand U9390 (N_9390,In_1320,In_1741);
and U9391 (N_9391,In_52,In_1853);
nor U9392 (N_9392,In_2072,In_192);
nor U9393 (N_9393,In_2555,In_2762);
and U9394 (N_9394,In_2744,In_614);
and U9395 (N_9395,In_2150,In_2437);
nand U9396 (N_9396,In_2933,In_1676);
and U9397 (N_9397,In_1944,In_1943);
nand U9398 (N_9398,In_696,In_589);
nand U9399 (N_9399,In_2670,In_2905);
nor U9400 (N_9400,In_2909,In_379);
nor U9401 (N_9401,In_105,In_1398);
or U9402 (N_9402,In_1523,In_1293);
and U9403 (N_9403,In_2292,In_1572);
nand U9404 (N_9404,In_256,In_2622);
and U9405 (N_9405,In_24,In_1798);
or U9406 (N_9406,In_1327,In_2430);
and U9407 (N_9407,In_886,In_1263);
nand U9408 (N_9408,In_938,In_1062);
or U9409 (N_9409,In_1589,In_327);
and U9410 (N_9410,In_2637,In_2904);
xor U9411 (N_9411,In_2424,In_670);
or U9412 (N_9412,In_1460,In_1499);
and U9413 (N_9413,In_2948,In_1775);
nor U9414 (N_9414,In_506,In_961);
or U9415 (N_9415,In_590,In_1855);
nand U9416 (N_9416,In_1371,In_1967);
nand U9417 (N_9417,In_1424,In_2930);
nand U9418 (N_9418,In_930,In_854);
or U9419 (N_9419,In_1244,In_2729);
nand U9420 (N_9420,In_1618,In_954);
nand U9421 (N_9421,In_527,In_2571);
nand U9422 (N_9422,In_606,In_1554);
and U9423 (N_9423,In_2179,In_2940);
and U9424 (N_9424,In_1873,In_174);
nand U9425 (N_9425,In_939,In_544);
nor U9426 (N_9426,In_1352,In_103);
or U9427 (N_9427,In_1855,In_1684);
nor U9428 (N_9428,In_2851,In_2434);
and U9429 (N_9429,In_2667,In_2156);
nand U9430 (N_9430,In_1589,In_42);
xor U9431 (N_9431,In_759,In_1413);
and U9432 (N_9432,In_64,In_1017);
nand U9433 (N_9433,In_1563,In_1410);
and U9434 (N_9434,In_2031,In_2099);
and U9435 (N_9435,In_809,In_2806);
or U9436 (N_9436,In_1510,In_2496);
nand U9437 (N_9437,In_2901,In_579);
or U9438 (N_9438,In_1383,In_2888);
and U9439 (N_9439,In_684,In_503);
and U9440 (N_9440,In_1726,In_1888);
and U9441 (N_9441,In_197,In_1959);
and U9442 (N_9442,In_2750,In_2480);
or U9443 (N_9443,In_965,In_54);
nand U9444 (N_9444,In_2974,In_1151);
or U9445 (N_9445,In_2649,In_1265);
and U9446 (N_9446,In_2944,In_2385);
and U9447 (N_9447,In_183,In_788);
or U9448 (N_9448,In_1311,In_1452);
and U9449 (N_9449,In_2312,In_557);
nand U9450 (N_9450,In_2518,In_1824);
nand U9451 (N_9451,In_221,In_494);
and U9452 (N_9452,In_661,In_763);
nand U9453 (N_9453,In_1500,In_2868);
or U9454 (N_9454,In_1878,In_782);
or U9455 (N_9455,In_1025,In_60);
nor U9456 (N_9456,In_769,In_2759);
and U9457 (N_9457,In_1710,In_2817);
nor U9458 (N_9458,In_2771,In_1359);
nor U9459 (N_9459,In_1220,In_282);
or U9460 (N_9460,In_1141,In_1831);
nor U9461 (N_9461,In_270,In_914);
and U9462 (N_9462,In_2441,In_1107);
or U9463 (N_9463,In_1046,In_1727);
nor U9464 (N_9464,In_1053,In_2080);
and U9465 (N_9465,In_2206,In_2350);
nor U9466 (N_9466,In_1468,In_2624);
nand U9467 (N_9467,In_1911,In_270);
or U9468 (N_9468,In_974,In_1313);
nor U9469 (N_9469,In_2481,In_1321);
or U9470 (N_9470,In_1361,In_2416);
and U9471 (N_9471,In_1657,In_428);
nand U9472 (N_9472,In_741,In_2967);
and U9473 (N_9473,In_879,In_2329);
nand U9474 (N_9474,In_479,In_825);
or U9475 (N_9475,In_93,In_1430);
or U9476 (N_9476,In_1307,In_256);
xnor U9477 (N_9477,In_1218,In_1023);
or U9478 (N_9478,In_2957,In_970);
nor U9479 (N_9479,In_2369,In_714);
nand U9480 (N_9480,In_1277,In_1737);
nand U9481 (N_9481,In_894,In_2290);
or U9482 (N_9482,In_1374,In_2312);
and U9483 (N_9483,In_1167,In_1460);
and U9484 (N_9484,In_1790,In_1475);
and U9485 (N_9485,In_1126,In_2816);
nor U9486 (N_9486,In_2114,In_1325);
and U9487 (N_9487,In_1960,In_315);
nor U9488 (N_9488,In_978,In_2559);
nand U9489 (N_9489,In_2071,In_86);
nor U9490 (N_9490,In_2633,In_918);
nor U9491 (N_9491,In_1990,In_8);
and U9492 (N_9492,In_1402,In_2523);
nor U9493 (N_9493,In_2820,In_1861);
and U9494 (N_9494,In_1942,In_2722);
xor U9495 (N_9495,In_543,In_505);
nor U9496 (N_9496,In_228,In_2491);
or U9497 (N_9497,In_2897,In_1225);
nor U9498 (N_9498,In_788,In_2899);
or U9499 (N_9499,In_2658,In_93);
or U9500 (N_9500,In_1933,In_332);
nand U9501 (N_9501,In_322,In_2851);
or U9502 (N_9502,In_618,In_2587);
and U9503 (N_9503,In_2159,In_64);
nor U9504 (N_9504,In_2715,In_562);
nand U9505 (N_9505,In_1119,In_859);
and U9506 (N_9506,In_357,In_180);
or U9507 (N_9507,In_1409,In_1190);
nand U9508 (N_9508,In_553,In_2814);
or U9509 (N_9509,In_1418,In_1883);
nand U9510 (N_9510,In_202,In_2770);
or U9511 (N_9511,In_384,In_260);
nand U9512 (N_9512,In_2443,In_1296);
and U9513 (N_9513,In_2550,In_868);
and U9514 (N_9514,In_983,In_978);
nand U9515 (N_9515,In_1329,In_1656);
and U9516 (N_9516,In_670,In_1380);
nand U9517 (N_9517,In_572,In_1768);
and U9518 (N_9518,In_1283,In_1106);
and U9519 (N_9519,In_2560,In_1058);
nor U9520 (N_9520,In_2626,In_1466);
or U9521 (N_9521,In_1751,In_1267);
nand U9522 (N_9522,In_1037,In_1805);
and U9523 (N_9523,In_1634,In_154);
and U9524 (N_9524,In_1178,In_2500);
nand U9525 (N_9525,In_178,In_1740);
or U9526 (N_9526,In_883,In_1353);
nor U9527 (N_9527,In_2097,In_2059);
or U9528 (N_9528,In_4,In_1235);
nor U9529 (N_9529,In_1121,In_178);
or U9530 (N_9530,In_582,In_824);
nand U9531 (N_9531,In_1120,In_1437);
nor U9532 (N_9532,In_2480,In_2702);
or U9533 (N_9533,In_1428,In_2725);
or U9534 (N_9534,In_2533,In_1015);
nor U9535 (N_9535,In_1081,In_1618);
or U9536 (N_9536,In_1823,In_242);
xor U9537 (N_9537,In_566,In_1493);
or U9538 (N_9538,In_2135,In_114);
nand U9539 (N_9539,In_1761,In_2279);
nand U9540 (N_9540,In_2360,In_171);
or U9541 (N_9541,In_2468,In_2485);
nand U9542 (N_9542,In_1191,In_439);
or U9543 (N_9543,In_2939,In_2138);
nand U9544 (N_9544,In_1768,In_2643);
or U9545 (N_9545,In_24,In_908);
nor U9546 (N_9546,In_2134,In_2138);
nand U9547 (N_9547,In_36,In_583);
nor U9548 (N_9548,In_1403,In_239);
or U9549 (N_9549,In_1929,In_1503);
and U9550 (N_9550,In_1629,In_166);
and U9551 (N_9551,In_2112,In_2097);
nor U9552 (N_9552,In_1050,In_565);
nor U9553 (N_9553,In_337,In_650);
nand U9554 (N_9554,In_1574,In_2834);
nor U9555 (N_9555,In_1451,In_85);
nor U9556 (N_9556,In_2129,In_2672);
nand U9557 (N_9557,In_1029,In_1686);
nand U9558 (N_9558,In_2380,In_140);
nand U9559 (N_9559,In_2100,In_547);
nor U9560 (N_9560,In_951,In_2631);
and U9561 (N_9561,In_475,In_1430);
nand U9562 (N_9562,In_1778,In_1617);
and U9563 (N_9563,In_1829,In_1925);
or U9564 (N_9564,In_1361,In_998);
nor U9565 (N_9565,In_324,In_2800);
nor U9566 (N_9566,In_2676,In_654);
and U9567 (N_9567,In_2198,In_434);
or U9568 (N_9568,In_1538,In_452);
and U9569 (N_9569,In_465,In_718);
xor U9570 (N_9570,In_1263,In_1895);
nor U9571 (N_9571,In_120,In_227);
and U9572 (N_9572,In_2416,In_644);
nor U9573 (N_9573,In_2946,In_1377);
nand U9574 (N_9574,In_95,In_1424);
and U9575 (N_9575,In_7,In_1660);
or U9576 (N_9576,In_1330,In_1304);
or U9577 (N_9577,In_2136,In_90);
nand U9578 (N_9578,In_1066,In_2916);
or U9579 (N_9579,In_1819,In_2999);
or U9580 (N_9580,In_65,In_629);
and U9581 (N_9581,In_2586,In_1429);
nor U9582 (N_9582,In_2458,In_649);
and U9583 (N_9583,In_1993,In_2436);
or U9584 (N_9584,In_882,In_1961);
nand U9585 (N_9585,In_1302,In_1315);
and U9586 (N_9586,In_1719,In_2730);
nand U9587 (N_9587,In_17,In_166);
nor U9588 (N_9588,In_2829,In_2005);
nand U9589 (N_9589,In_1851,In_1443);
nand U9590 (N_9590,In_444,In_2208);
nand U9591 (N_9591,In_80,In_1236);
nand U9592 (N_9592,In_1078,In_482);
and U9593 (N_9593,In_2061,In_1556);
or U9594 (N_9594,In_2416,In_2110);
and U9595 (N_9595,In_1051,In_770);
and U9596 (N_9596,In_655,In_71);
or U9597 (N_9597,In_893,In_757);
nor U9598 (N_9598,In_756,In_152);
nor U9599 (N_9599,In_2955,In_1301);
and U9600 (N_9600,In_142,In_1584);
nor U9601 (N_9601,In_774,In_42);
or U9602 (N_9602,In_2882,In_1887);
nor U9603 (N_9603,In_1760,In_1358);
nand U9604 (N_9604,In_87,In_2382);
and U9605 (N_9605,In_470,In_1292);
and U9606 (N_9606,In_961,In_2400);
and U9607 (N_9607,In_1114,In_1282);
or U9608 (N_9608,In_441,In_1437);
nor U9609 (N_9609,In_340,In_1950);
or U9610 (N_9610,In_2532,In_1568);
or U9611 (N_9611,In_2785,In_810);
and U9612 (N_9612,In_2971,In_1369);
nor U9613 (N_9613,In_925,In_1223);
nor U9614 (N_9614,In_208,In_1177);
nand U9615 (N_9615,In_253,In_1940);
nor U9616 (N_9616,In_502,In_887);
nor U9617 (N_9617,In_2014,In_1744);
nand U9618 (N_9618,In_326,In_2480);
or U9619 (N_9619,In_2433,In_2156);
or U9620 (N_9620,In_1373,In_1050);
and U9621 (N_9621,In_1397,In_355);
nor U9622 (N_9622,In_2474,In_2037);
nor U9623 (N_9623,In_363,In_1920);
or U9624 (N_9624,In_1529,In_114);
or U9625 (N_9625,In_2859,In_2270);
nor U9626 (N_9626,In_588,In_2151);
nor U9627 (N_9627,In_281,In_447);
and U9628 (N_9628,In_578,In_2576);
and U9629 (N_9629,In_1803,In_2881);
and U9630 (N_9630,In_178,In_2624);
and U9631 (N_9631,In_506,In_1031);
nand U9632 (N_9632,In_1648,In_2362);
nand U9633 (N_9633,In_1163,In_55);
and U9634 (N_9634,In_322,In_719);
and U9635 (N_9635,In_489,In_293);
and U9636 (N_9636,In_1054,In_2140);
nand U9637 (N_9637,In_1125,In_1812);
or U9638 (N_9638,In_378,In_699);
and U9639 (N_9639,In_581,In_292);
nand U9640 (N_9640,In_1349,In_1677);
and U9641 (N_9641,In_267,In_1846);
nor U9642 (N_9642,In_2463,In_851);
and U9643 (N_9643,In_493,In_2564);
nor U9644 (N_9644,In_2131,In_2864);
nand U9645 (N_9645,In_2489,In_2029);
nand U9646 (N_9646,In_1813,In_253);
nand U9647 (N_9647,In_170,In_788);
nand U9648 (N_9648,In_1650,In_749);
and U9649 (N_9649,In_2862,In_2542);
nand U9650 (N_9650,In_869,In_2000);
and U9651 (N_9651,In_2652,In_2706);
and U9652 (N_9652,In_678,In_1656);
nor U9653 (N_9653,In_1395,In_174);
or U9654 (N_9654,In_107,In_2298);
nand U9655 (N_9655,In_317,In_2725);
nor U9656 (N_9656,In_396,In_2036);
nor U9657 (N_9657,In_1351,In_1431);
and U9658 (N_9658,In_1756,In_1788);
nor U9659 (N_9659,In_267,In_706);
nand U9660 (N_9660,In_1414,In_447);
and U9661 (N_9661,In_1213,In_843);
and U9662 (N_9662,In_1432,In_1306);
nor U9663 (N_9663,In_875,In_2151);
nor U9664 (N_9664,In_1299,In_2527);
or U9665 (N_9665,In_706,In_814);
and U9666 (N_9666,In_313,In_1205);
and U9667 (N_9667,In_1782,In_47);
nand U9668 (N_9668,In_1437,In_2691);
or U9669 (N_9669,In_1485,In_2085);
nor U9670 (N_9670,In_1645,In_1218);
or U9671 (N_9671,In_1523,In_2338);
or U9672 (N_9672,In_1088,In_34);
or U9673 (N_9673,In_387,In_216);
or U9674 (N_9674,In_1134,In_338);
nor U9675 (N_9675,In_1606,In_2463);
and U9676 (N_9676,In_1626,In_1460);
nand U9677 (N_9677,In_1535,In_729);
and U9678 (N_9678,In_2705,In_1457);
and U9679 (N_9679,In_2713,In_669);
or U9680 (N_9680,In_1115,In_1698);
and U9681 (N_9681,In_2217,In_2203);
nor U9682 (N_9682,In_732,In_1785);
nand U9683 (N_9683,In_2068,In_2335);
or U9684 (N_9684,In_30,In_1886);
or U9685 (N_9685,In_1918,In_1166);
or U9686 (N_9686,In_2,In_2666);
or U9687 (N_9687,In_2238,In_351);
nand U9688 (N_9688,In_1442,In_494);
nor U9689 (N_9689,In_41,In_1203);
nand U9690 (N_9690,In_2414,In_115);
nand U9691 (N_9691,In_2387,In_341);
nand U9692 (N_9692,In_1943,In_2354);
and U9693 (N_9693,In_1826,In_491);
nor U9694 (N_9694,In_768,In_1657);
and U9695 (N_9695,In_1980,In_2211);
nand U9696 (N_9696,In_2,In_898);
or U9697 (N_9697,In_1597,In_387);
nor U9698 (N_9698,In_1397,In_1024);
or U9699 (N_9699,In_1096,In_1605);
or U9700 (N_9700,In_424,In_122);
nor U9701 (N_9701,In_318,In_660);
nor U9702 (N_9702,In_1878,In_2058);
or U9703 (N_9703,In_964,In_565);
nor U9704 (N_9704,In_106,In_467);
nor U9705 (N_9705,In_1419,In_712);
and U9706 (N_9706,In_2410,In_273);
nand U9707 (N_9707,In_2178,In_332);
and U9708 (N_9708,In_1634,In_1501);
or U9709 (N_9709,In_1891,In_1551);
nand U9710 (N_9710,In_1785,In_2821);
and U9711 (N_9711,In_2519,In_717);
or U9712 (N_9712,In_2682,In_2059);
nand U9713 (N_9713,In_1424,In_1456);
nor U9714 (N_9714,In_1494,In_2753);
or U9715 (N_9715,In_2637,In_576);
and U9716 (N_9716,In_533,In_91);
nand U9717 (N_9717,In_439,In_1026);
or U9718 (N_9718,In_1229,In_2834);
and U9719 (N_9719,In_1890,In_1467);
or U9720 (N_9720,In_2849,In_771);
or U9721 (N_9721,In_1421,In_2535);
nand U9722 (N_9722,In_2253,In_1753);
and U9723 (N_9723,In_1588,In_2757);
nand U9724 (N_9724,In_226,In_2290);
nor U9725 (N_9725,In_225,In_2606);
nand U9726 (N_9726,In_662,In_725);
or U9727 (N_9727,In_1282,In_939);
nand U9728 (N_9728,In_326,In_227);
nor U9729 (N_9729,In_1254,In_1455);
or U9730 (N_9730,In_64,In_2513);
nand U9731 (N_9731,In_1589,In_2716);
or U9732 (N_9732,In_927,In_1631);
nand U9733 (N_9733,In_836,In_1521);
and U9734 (N_9734,In_733,In_2124);
or U9735 (N_9735,In_1671,In_1209);
nand U9736 (N_9736,In_1735,In_379);
nand U9737 (N_9737,In_2473,In_1149);
and U9738 (N_9738,In_1599,In_2840);
nor U9739 (N_9739,In_1132,In_458);
nand U9740 (N_9740,In_1864,In_2585);
and U9741 (N_9741,In_2318,In_1702);
or U9742 (N_9742,In_1754,In_507);
and U9743 (N_9743,In_1483,In_1447);
nand U9744 (N_9744,In_296,In_774);
and U9745 (N_9745,In_2836,In_2480);
or U9746 (N_9746,In_477,In_1413);
and U9747 (N_9747,In_2572,In_53);
and U9748 (N_9748,In_2989,In_2362);
nand U9749 (N_9749,In_279,In_464);
or U9750 (N_9750,In_1787,In_1066);
nor U9751 (N_9751,In_1284,In_2658);
or U9752 (N_9752,In_2623,In_2909);
nand U9753 (N_9753,In_1515,In_893);
nand U9754 (N_9754,In_1295,In_2785);
nor U9755 (N_9755,In_1809,In_97);
nor U9756 (N_9756,In_2928,In_2057);
nand U9757 (N_9757,In_1415,In_2775);
nand U9758 (N_9758,In_882,In_199);
or U9759 (N_9759,In_79,In_690);
nand U9760 (N_9760,In_2718,In_2104);
nand U9761 (N_9761,In_2434,In_615);
or U9762 (N_9762,In_1438,In_2413);
or U9763 (N_9763,In_476,In_1552);
and U9764 (N_9764,In_2741,In_1456);
or U9765 (N_9765,In_2658,In_137);
and U9766 (N_9766,In_872,In_360);
or U9767 (N_9767,In_15,In_2673);
and U9768 (N_9768,In_597,In_2382);
and U9769 (N_9769,In_1994,In_1197);
or U9770 (N_9770,In_2021,In_2580);
nand U9771 (N_9771,In_1438,In_1148);
nor U9772 (N_9772,In_1172,In_503);
or U9773 (N_9773,In_1424,In_689);
or U9774 (N_9774,In_2578,In_1918);
nand U9775 (N_9775,In_2665,In_1868);
nand U9776 (N_9776,In_294,In_220);
or U9777 (N_9777,In_1111,In_1697);
xor U9778 (N_9778,In_1359,In_2533);
nor U9779 (N_9779,In_1378,In_940);
nor U9780 (N_9780,In_64,In_1726);
nand U9781 (N_9781,In_1783,In_841);
nor U9782 (N_9782,In_2830,In_2134);
nand U9783 (N_9783,In_2455,In_1483);
or U9784 (N_9784,In_401,In_2156);
and U9785 (N_9785,In_2083,In_130);
nor U9786 (N_9786,In_196,In_732);
or U9787 (N_9787,In_1345,In_519);
nor U9788 (N_9788,In_976,In_2643);
nor U9789 (N_9789,In_200,In_121);
and U9790 (N_9790,In_2621,In_820);
nor U9791 (N_9791,In_1727,In_1698);
or U9792 (N_9792,In_1223,In_2473);
nand U9793 (N_9793,In_2081,In_1120);
nor U9794 (N_9794,In_1369,In_2541);
nor U9795 (N_9795,In_2910,In_2635);
nor U9796 (N_9796,In_769,In_845);
nand U9797 (N_9797,In_1388,In_2495);
nand U9798 (N_9798,In_2770,In_2370);
nor U9799 (N_9799,In_896,In_1500);
nand U9800 (N_9800,In_1957,In_2146);
nand U9801 (N_9801,In_98,In_2211);
and U9802 (N_9802,In_545,In_1230);
and U9803 (N_9803,In_2385,In_553);
or U9804 (N_9804,In_2408,In_519);
nand U9805 (N_9805,In_1746,In_1368);
or U9806 (N_9806,In_1047,In_2129);
and U9807 (N_9807,In_9,In_1767);
and U9808 (N_9808,In_916,In_317);
nor U9809 (N_9809,In_1420,In_1298);
and U9810 (N_9810,In_835,In_1056);
or U9811 (N_9811,In_1197,In_840);
nor U9812 (N_9812,In_2847,In_1345);
nor U9813 (N_9813,In_853,In_2529);
or U9814 (N_9814,In_2229,In_272);
nand U9815 (N_9815,In_233,In_2127);
nor U9816 (N_9816,In_1555,In_2153);
nor U9817 (N_9817,In_1833,In_2564);
nor U9818 (N_9818,In_773,In_1667);
nand U9819 (N_9819,In_2173,In_2197);
nand U9820 (N_9820,In_1283,In_1292);
nor U9821 (N_9821,In_2422,In_2888);
or U9822 (N_9822,In_2501,In_2966);
nand U9823 (N_9823,In_1381,In_1478);
and U9824 (N_9824,In_2989,In_2871);
nor U9825 (N_9825,In_1086,In_2192);
nand U9826 (N_9826,In_409,In_1440);
and U9827 (N_9827,In_2824,In_2194);
or U9828 (N_9828,In_2950,In_2023);
and U9829 (N_9829,In_180,In_503);
and U9830 (N_9830,In_1398,In_1108);
and U9831 (N_9831,In_2873,In_2073);
nor U9832 (N_9832,In_1828,In_1720);
or U9833 (N_9833,In_736,In_2922);
nor U9834 (N_9834,In_613,In_1361);
and U9835 (N_9835,In_69,In_2472);
and U9836 (N_9836,In_754,In_1331);
nor U9837 (N_9837,In_2257,In_788);
nor U9838 (N_9838,In_835,In_2195);
nor U9839 (N_9839,In_781,In_10);
or U9840 (N_9840,In_1429,In_770);
nand U9841 (N_9841,In_485,In_222);
nand U9842 (N_9842,In_2754,In_1876);
nor U9843 (N_9843,In_1946,In_364);
or U9844 (N_9844,In_1004,In_2542);
nand U9845 (N_9845,In_2270,In_726);
nand U9846 (N_9846,In_289,In_936);
and U9847 (N_9847,In_1931,In_1163);
or U9848 (N_9848,In_1223,In_1267);
nand U9849 (N_9849,In_699,In_1276);
and U9850 (N_9850,In_2896,In_2602);
or U9851 (N_9851,In_201,In_1245);
or U9852 (N_9852,In_1949,In_1008);
nand U9853 (N_9853,In_1517,In_371);
and U9854 (N_9854,In_349,In_1188);
and U9855 (N_9855,In_1682,In_2267);
or U9856 (N_9856,In_1152,In_2906);
and U9857 (N_9857,In_940,In_350);
or U9858 (N_9858,In_2951,In_293);
or U9859 (N_9859,In_2031,In_1292);
nand U9860 (N_9860,In_2715,In_1088);
nor U9861 (N_9861,In_613,In_2671);
nand U9862 (N_9862,In_2187,In_2633);
nor U9863 (N_9863,In_514,In_2867);
nand U9864 (N_9864,In_1766,In_838);
and U9865 (N_9865,In_119,In_1033);
or U9866 (N_9866,In_572,In_1997);
nand U9867 (N_9867,In_1119,In_235);
and U9868 (N_9868,In_2568,In_2365);
nand U9869 (N_9869,In_1389,In_2614);
and U9870 (N_9870,In_1236,In_1705);
nor U9871 (N_9871,In_290,In_2205);
and U9872 (N_9872,In_731,In_1831);
nor U9873 (N_9873,In_143,In_362);
or U9874 (N_9874,In_2662,In_2668);
nor U9875 (N_9875,In_189,In_1497);
or U9876 (N_9876,In_1301,In_1471);
and U9877 (N_9877,In_1247,In_936);
nor U9878 (N_9878,In_574,In_691);
xnor U9879 (N_9879,In_2301,In_2508);
or U9880 (N_9880,In_1136,In_234);
or U9881 (N_9881,In_1555,In_567);
nor U9882 (N_9882,In_1821,In_2532);
nor U9883 (N_9883,In_308,In_1515);
and U9884 (N_9884,In_2936,In_249);
and U9885 (N_9885,In_1716,In_1541);
or U9886 (N_9886,In_1292,In_620);
or U9887 (N_9887,In_1190,In_1500);
and U9888 (N_9888,In_268,In_2962);
nor U9889 (N_9889,In_922,In_487);
nor U9890 (N_9890,In_1171,In_707);
nor U9891 (N_9891,In_2515,In_1835);
nor U9892 (N_9892,In_1503,In_1257);
and U9893 (N_9893,In_1161,In_2382);
and U9894 (N_9894,In_618,In_1512);
nand U9895 (N_9895,In_2119,In_2794);
or U9896 (N_9896,In_1788,In_939);
nor U9897 (N_9897,In_2615,In_983);
nand U9898 (N_9898,In_2688,In_2690);
or U9899 (N_9899,In_1840,In_557);
or U9900 (N_9900,In_1741,In_2388);
xor U9901 (N_9901,In_851,In_1226);
or U9902 (N_9902,In_550,In_2787);
or U9903 (N_9903,In_2140,In_2603);
nor U9904 (N_9904,In_1544,In_981);
and U9905 (N_9905,In_1494,In_841);
or U9906 (N_9906,In_2998,In_731);
nor U9907 (N_9907,In_219,In_506);
or U9908 (N_9908,In_2733,In_889);
nand U9909 (N_9909,In_1595,In_1276);
or U9910 (N_9910,In_454,In_266);
nor U9911 (N_9911,In_1868,In_2895);
nor U9912 (N_9912,In_2990,In_182);
nand U9913 (N_9913,In_232,In_2334);
nor U9914 (N_9914,In_1728,In_1084);
nand U9915 (N_9915,In_513,In_1691);
or U9916 (N_9916,In_2848,In_1678);
nand U9917 (N_9917,In_1078,In_2166);
or U9918 (N_9918,In_1203,In_718);
nor U9919 (N_9919,In_1066,In_944);
or U9920 (N_9920,In_402,In_193);
nand U9921 (N_9921,In_2777,In_1160);
nand U9922 (N_9922,In_2526,In_929);
nand U9923 (N_9923,In_2975,In_2609);
nand U9924 (N_9924,In_1146,In_1562);
nor U9925 (N_9925,In_2478,In_1088);
nand U9926 (N_9926,In_97,In_1794);
nor U9927 (N_9927,In_1071,In_2753);
and U9928 (N_9928,In_2017,In_2661);
nand U9929 (N_9929,In_2990,In_1274);
or U9930 (N_9930,In_186,In_2014);
or U9931 (N_9931,In_1956,In_2489);
and U9932 (N_9932,In_64,In_2403);
and U9933 (N_9933,In_1706,In_2177);
nand U9934 (N_9934,In_546,In_1726);
and U9935 (N_9935,In_1543,In_2979);
or U9936 (N_9936,In_2840,In_1410);
nand U9937 (N_9937,In_1028,In_2598);
or U9938 (N_9938,In_1260,In_31);
and U9939 (N_9939,In_901,In_1962);
nand U9940 (N_9940,In_2716,In_2150);
nor U9941 (N_9941,In_2595,In_519);
nand U9942 (N_9942,In_2893,In_273);
and U9943 (N_9943,In_667,In_685);
nor U9944 (N_9944,In_2471,In_893);
nand U9945 (N_9945,In_1807,In_1117);
and U9946 (N_9946,In_135,In_2098);
nor U9947 (N_9947,In_831,In_1839);
nor U9948 (N_9948,In_2529,In_459);
and U9949 (N_9949,In_255,In_1946);
or U9950 (N_9950,In_1460,In_2497);
or U9951 (N_9951,In_2876,In_1076);
xnor U9952 (N_9952,In_1878,In_467);
or U9953 (N_9953,In_1642,In_481);
and U9954 (N_9954,In_1050,In_1795);
nor U9955 (N_9955,In_2548,In_1930);
and U9956 (N_9956,In_2842,In_619);
nor U9957 (N_9957,In_1450,In_1749);
nand U9958 (N_9958,In_2206,In_2393);
nor U9959 (N_9959,In_579,In_64);
or U9960 (N_9960,In_2250,In_1912);
and U9961 (N_9961,In_1951,In_1723);
and U9962 (N_9962,In_92,In_2452);
or U9963 (N_9963,In_2309,In_1198);
nand U9964 (N_9964,In_1931,In_647);
and U9965 (N_9965,In_244,In_2878);
nand U9966 (N_9966,In_1282,In_1916);
or U9967 (N_9967,In_980,In_1231);
nand U9968 (N_9968,In_1098,In_2812);
and U9969 (N_9969,In_2006,In_2194);
or U9970 (N_9970,In_442,In_86);
nand U9971 (N_9971,In_1901,In_617);
nor U9972 (N_9972,In_427,In_2628);
nor U9973 (N_9973,In_2693,In_2784);
or U9974 (N_9974,In_971,In_1175);
and U9975 (N_9975,In_2832,In_598);
nand U9976 (N_9976,In_1020,In_2232);
nor U9977 (N_9977,In_1459,In_1932);
and U9978 (N_9978,In_384,In_1609);
nand U9979 (N_9979,In_702,In_1641);
and U9980 (N_9980,In_2795,In_908);
or U9981 (N_9981,In_699,In_2544);
nor U9982 (N_9982,In_276,In_2875);
nand U9983 (N_9983,In_701,In_2990);
and U9984 (N_9984,In_81,In_529);
or U9985 (N_9985,In_212,In_349);
or U9986 (N_9986,In_1151,In_1265);
xor U9987 (N_9987,In_2697,In_869);
nand U9988 (N_9988,In_80,In_2344);
or U9989 (N_9989,In_879,In_2469);
and U9990 (N_9990,In_403,In_1098);
and U9991 (N_9991,In_71,In_2273);
or U9992 (N_9992,In_725,In_1782);
nor U9993 (N_9993,In_1497,In_2005);
nor U9994 (N_9994,In_2360,In_621);
nand U9995 (N_9995,In_2465,In_414);
nand U9996 (N_9996,In_2165,In_646);
nand U9997 (N_9997,In_2715,In_2499);
or U9998 (N_9998,In_2195,In_757);
and U9999 (N_9999,In_2057,In_138);
nand U10000 (N_10000,N_2700,N_2916);
or U10001 (N_10001,N_9698,N_2580);
nor U10002 (N_10002,N_3787,N_3992);
or U10003 (N_10003,N_6742,N_140);
nand U10004 (N_10004,N_2088,N_7879);
and U10005 (N_10005,N_6774,N_9404);
nand U10006 (N_10006,N_6151,N_520);
nor U10007 (N_10007,N_9344,N_2646);
or U10008 (N_10008,N_648,N_4225);
nor U10009 (N_10009,N_5866,N_8349);
nand U10010 (N_10010,N_1309,N_3591);
or U10011 (N_10011,N_1914,N_5540);
nand U10012 (N_10012,N_9573,N_5971);
nand U10013 (N_10013,N_7523,N_8244);
or U10014 (N_10014,N_8202,N_713);
or U10015 (N_10015,N_6492,N_3994);
nand U10016 (N_10016,N_9565,N_7071);
and U10017 (N_10017,N_381,N_7790);
nor U10018 (N_10018,N_9209,N_6285);
or U10019 (N_10019,N_9729,N_6510);
and U10020 (N_10020,N_4954,N_8576);
nor U10021 (N_10021,N_6807,N_6697);
or U10022 (N_10022,N_5995,N_6192);
and U10023 (N_10023,N_639,N_8800);
nand U10024 (N_10024,N_502,N_5180);
or U10025 (N_10025,N_9616,N_7875);
nor U10026 (N_10026,N_8520,N_6638);
and U10027 (N_10027,N_4023,N_324);
and U10028 (N_10028,N_6511,N_8342);
nand U10029 (N_10029,N_8986,N_5408);
nand U10030 (N_10030,N_4646,N_9882);
nor U10031 (N_10031,N_6760,N_489);
nand U10032 (N_10032,N_8731,N_8238);
or U10033 (N_10033,N_3716,N_4893);
or U10034 (N_10034,N_9776,N_7270);
or U10035 (N_10035,N_6162,N_7215);
nor U10036 (N_10036,N_1066,N_4339);
or U10037 (N_10037,N_9241,N_7479);
and U10038 (N_10038,N_3327,N_8114);
nor U10039 (N_10039,N_3764,N_1496);
and U10040 (N_10040,N_112,N_3410);
and U10041 (N_10041,N_6475,N_5535);
nor U10042 (N_10042,N_123,N_7385);
and U10043 (N_10043,N_3199,N_7932);
and U10044 (N_10044,N_8968,N_9387);
and U10045 (N_10045,N_9763,N_3677);
and U10046 (N_10046,N_79,N_6999);
nand U10047 (N_10047,N_396,N_8888);
and U10048 (N_10048,N_8209,N_6332);
and U10049 (N_10049,N_4425,N_6426);
nor U10050 (N_10050,N_2972,N_4113);
nand U10051 (N_10051,N_2125,N_8214);
or U10052 (N_10052,N_7151,N_40);
and U10053 (N_10053,N_8021,N_6878);
nor U10054 (N_10054,N_5359,N_2904);
nand U10055 (N_10055,N_3974,N_542);
or U10056 (N_10056,N_1673,N_7955);
nor U10057 (N_10057,N_3499,N_2309);
nor U10058 (N_10058,N_1121,N_3569);
nand U10059 (N_10059,N_6272,N_8460);
nor U10060 (N_10060,N_4866,N_6078);
or U10061 (N_10061,N_6199,N_1377);
nand U10062 (N_10062,N_2147,N_5494);
nor U10063 (N_10063,N_3283,N_5178);
nor U10064 (N_10064,N_5271,N_7830);
xnor U10065 (N_10065,N_5794,N_793);
nand U10066 (N_10066,N_5083,N_8502);
and U10067 (N_10067,N_1549,N_9701);
nor U10068 (N_10068,N_1832,N_8675);
nor U10069 (N_10069,N_6471,N_7319);
nand U10070 (N_10070,N_7450,N_6743);
nor U10071 (N_10071,N_4544,N_113);
or U10072 (N_10072,N_3048,N_3537);
nand U10073 (N_10073,N_1768,N_5331);
nor U10074 (N_10074,N_4024,N_3091);
or U10075 (N_10075,N_217,N_9984);
nor U10076 (N_10076,N_9694,N_8756);
and U10077 (N_10077,N_7880,N_6991);
nand U10078 (N_10078,N_4914,N_2883);
and U10079 (N_10079,N_5816,N_9875);
and U10080 (N_10080,N_775,N_6083);
nand U10081 (N_10081,N_2713,N_8147);
or U10082 (N_10082,N_5886,N_4801);
or U10083 (N_10083,N_3206,N_6022);
or U10084 (N_10084,N_6893,N_7108);
nor U10085 (N_10085,N_3865,N_8057);
or U10086 (N_10086,N_825,N_1636);
and U10087 (N_10087,N_4230,N_5952);
or U10088 (N_10088,N_4970,N_23);
nor U10089 (N_10089,N_951,N_6944);
or U10090 (N_10090,N_3980,N_1823);
nand U10091 (N_10091,N_1846,N_2599);
nor U10092 (N_10092,N_7914,N_1761);
nand U10093 (N_10093,N_2668,N_5675);
and U10094 (N_10094,N_4399,N_3768);
nand U10095 (N_10095,N_9775,N_9700);
nand U10096 (N_10096,N_5486,N_3093);
nor U10097 (N_10097,N_8016,N_9655);
nor U10098 (N_10098,N_322,N_3495);
and U10099 (N_10099,N_2430,N_4788);
nand U10100 (N_10100,N_9915,N_3377);
and U10101 (N_10101,N_4580,N_1555);
or U10102 (N_10102,N_9502,N_2057);
or U10103 (N_10103,N_1136,N_8055);
and U10104 (N_10104,N_8599,N_9372);
nor U10105 (N_10105,N_8827,N_7553);
or U10106 (N_10106,N_6861,N_4984);
nand U10107 (N_10107,N_496,N_9738);
nand U10108 (N_10108,N_8984,N_3727);
nand U10109 (N_10109,N_629,N_7721);
nand U10110 (N_10110,N_9708,N_2681);
or U10111 (N_10111,N_6460,N_2334);
and U10112 (N_10112,N_514,N_9749);
and U10113 (N_10113,N_6675,N_5517);
nor U10114 (N_10114,N_1610,N_4329);
and U10115 (N_10115,N_4175,N_2265);
nand U10116 (N_10116,N_9699,N_7736);
nor U10117 (N_10117,N_1539,N_854);
or U10118 (N_10118,N_7083,N_1645);
and U10119 (N_10119,N_4516,N_220);
and U10120 (N_10120,N_9881,N_5684);
or U10121 (N_10121,N_546,N_2472);
and U10122 (N_10122,N_9453,N_6410);
and U10123 (N_10123,N_1639,N_3270);
nor U10124 (N_10124,N_7172,N_9692);
or U10125 (N_10125,N_8645,N_8755);
nor U10126 (N_10126,N_1347,N_253);
nor U10127 (N_10127,N_9594,N_6731);
and U10128 (N_10128,N_273,N_1877);
nand U10129 (N_10129,N_4563,N_4238);
nand U10130 (N_10130,N_4409,N_4129);
nor U10131 (N_10131,N_6916,N_6322);
and U10132 (N_10132,N_5537,N_3651);
nand U10133 (N_10133,N_2453,N_7930);
nor U10134 (N_10134,N_3058,N_8039);
nand U10135 (N_10135,N_245,N_5039);
nor U10136 (N_10136,N_92,N_5880);
or U10137 (N_10137,N_4081,N_7009);
nor U10138 (N_10138,N_2263,N_5367);
or U10139 (N_10139,N_4445,N_5227);
and U10140 (N_10140,N_7053,N_8097);
nand U10141 (N_10141,N_557,N_4868);
nor U10142 (N_10142,N_7217,N_9173);
nor U10143 (N_10143,N_8913,N_3018);
xor U10144 (N_10144,N_3408,N_5115);
nor U10145 (N_10145,N_8562,N_6993);
nor U10146 (N_10146,N_2281,N_8668);
or U10147 (N_10147,N_4297,N_8872);
nor U10148 (N_10148,N_3543,N_8243);
or U10149 (N_10149,N_7119,N_7084);
and U10150 (N_10150,N_7923,N_3274);
or U10151 (N_10151,N_8464,N_2830);
nand U10152 (N_10152,N_5177,N_3471);
nor U10153 (N_10153,N_6350,N_1518);
or U10154 (N_10154,N_647,N_9551);
and U10155 (N_10155,N_8720,N_3373);
and U10156 (N_10156,N_6565,N_7670);
nor U10157 (N_10157,N_3067,N_5104);
nand U10158 (N_10158,N_5048,N_6722);
or U10159 (N_10159,N_4256,N_7289);
nand U10160 (N_10160,N_7438,N_2186);
and U10161 (N_10161,N_4761,N_677);
and U10162 (N_10162,N_8279,N_2261);
xor U10163 (N_10163,N_1769,N_3040);
nand U10164 (N_10164,N_3039,N_7537);
nor U10165 (N_10165,N_4688,N_884);
and U10166 (N_10166,N_4228,N_3717);
nor U10167 (N_10167,N_415,N_2441);
nand U10168 (N_10168,N_3969,N_4483);
nor U10169 (N_10169,N_650,N_3724);
and U10170 (N_10170,N_4180,N_2802);
or U10171 (N_10171,N_4921,N_2040);
nor U10172 (N_10172,N_2950,N_6023);
nand U10173 (N_10173,N_9552,N_3350);
and U10174 (N_10174,N_3598,N_5895);
or U10175 (N_10175,N_8833,N_3117);
and U10176 (N_10176,N_9941,N_4524);
nor U10177 (N_10177,N_9707,N_4336);
nor U10178 (N_10178,N_2491,N_9617);
or U10179 (N_10179,N_7744,N_5824);
and U10180 (N_10180,N_53,N_6099);
and U10181 (N_10181,N_303,N_4201);
or U10182 (N_10182,N_9156,N_3671);
xor U10183 (N_10183,N_4433,N_9505);
or U10184 (N_10184,N_1640,N_6113);
nor U10185 (N_10185,N_5449,N_495);
and U10186 (N_10186,N_3406,N_7219);
nand U10187 (N_10187,N_5044,N_686);
nand U10188 (N_10188,N_1473,N_8068);
or U10189 (N_10189,N_1429,N_1354);
or U10190 (N_10190,N_4928,N_9789);
nor U10191 (N_10191,N_1678,N_8127);
and U10192 (N_10192,N_3482,N_529);
or U10193 (N_10193,N_7858,N_5365);
nand U10194 (N_10194,N_8108,N_5043);
and U10195 (N_10195,N_4440,N_7019);
and U10196 (N_10196,N_4387,N_9538);
and U10197 (N_10197,N_4839,N_9382);
and U10198 (N_10198,N_4161,N_687);
nand U10199 (N_10199,N_7961,N_1974);
nand U10200 (N_10200,N_7771,N_3933);
nor U10201 (N_10201,N_1861,N_4687);
and U10202 (N_10202,N_8273,N_9019);
nand U10203 (N_10203,N_465,N_3839);
nor U10204 (N_10204,N_642,N_1030);
nor U10205 (N_10205,N_8171,N_5953);
nor U10206 (N_10206,N_5396,N_4089);
and U10207 (N_10207,N_3934,N_8894);
or U10208 (N_10208,N_5021,N_8981);
xor U10209 (N_10209,N_8960,N_3281);
or U10210 (N_10210,N_290,N_8264);
nor U10211 (N_10211,N_2322,N_3621);
and U10212 (N_10212,N_9548,N_1698);
or U10213 (N_10213,N_9049,N_6280);
nand U10214 (N_10214,N_1318,N_755);
or U10215 (N_10215,N_6705,N_5761);
nor U10216 (N_10216,N_836,N_9026);
nor U10217 (N_10217,N_9774,N_1452);
or U10218 (N_10218,N_100,N_4541);
nand U10219 (N_10219,N_8671,N_788);
or U10220 (N_10220,N_5395,N_6971);
nand U10221 (N_10221,N_2406,N_2448);
nor U10222 (N_10222,N_4488,N_816);
and U10223 (N_10223,N_8155,N_6803);
or U10224 (N_10224,N_987,N_2409);
xor U10225 (N_10225,N_6937,N_4342);
nand U10226 (N_10226,N_1020,N_726);
and U10227 (N_10227,N_9831,N_1023);
nand U10228 (N_10228,N_3036,N_990);
and U10229 (N_10229,N_1274,N_1133);
and U10230 (N_10230,N_6771,N_3129);
nand U10231 (N_10231,N_8431,N_7892);
nand U10232 (N_10232,N_785,N_3595);
nor U10233 (N_10233,N_3095,N_8775);
nand U10234 (N_10234,N_7872,N_2079);
or U10235 (N_10235,N_2195,N_916);
nor U10236 (N_10236,N_19,N_1268);
or U10237 (N_10237,N_8507,N_8985);
nand U10238 (N_10238,N_7052,N_6551);
and U10239 (N_10239,N_5538,N_9528);
and U10240 (N_10240,N_7583,N_919);
and U10241 (N_10241,N_5234,N_9833);
or U10242 (N_10242,N_292,N_314);
or U10243 (N_10243,N_447,N_924);
nand U10244 (N_10244,N_1538,N_2690);
nor U10245 (N_10245,N_6139,N_4739);
and U10246 (N_10246,N_2731,N_843);
nand U10247 (N_10247,N_76,N_414);
and U10248 (N_10248,N_9613,N_5727);
nor U10249 (N_10249,N_2848,N_5410);
xnor U10250 (N_10250,N_1467,N_662);
or U10251 (N_10251,N_638,N_5691);
and U10252 (N_10252,N_2849,N_9371);
nand U10253 (N_10253,N_8667,N_4527);
nor U10254 (N_10254,N_5547,N_6820);
nand U10255 (N_10255,N_8956,N_171);
and U10256 (N_10256,N_9444,N_5913);
nor U10257 (N_10257,N_519,N_7012);
nor U10258 (N_10258,N_3114,N_6300);
nor U10259 (N_10259,N_700,N_7336);
nor U10260 (N_10260,N_5798,N_7718);
xor U10261 (N_10261,N_8803,N_7051);
and U10262 (N_10262,N_9992,N_6919);
nor U10263 (N_10263,N_740,N_5503);
or U10264 (N_10264,N_3896,N_8063);
nor U10265 (N_10265,N_6443,N_3664);
nand U10266 (N_10266,N_1873,N_9126);
and U10267 (N_10267,N_8383,N_6571);
and U10268 (N_10268,N_5189,N_5338);
nand U10269 (N_10269,N_8194,N_6028);
nor U10270 (N_10270,N_5671,N_1000);
and U10271 (N_10271,N_7032,N_6415);
or U10272 (N_10272,N_5676,N_9290);
nor U10273 (N_10273,N_8554,N_5735);
or U10274 (N_10274,N_4709,N_5041);
nand U10275 (N_10275,N_7206,N_4345);
nor U10276 (N_10276,N_4176,N_9358);
nor U10277 (N_10277,N_5124,N_2412);
and U10278 (N_10278,N_1383,N_733);
nand U10279 (N_10279,N_2636,N_346);
nor U10280 (N_10280,N_6337,N_3593);
xnor U10281 (N_10281,N_5652,N_705);
nand U10282 (N_10282,N_5533,N_6989);
and U10283 (N_10283,N_663,N_7777);
or U10284 (N_10284,N_9213,N_3506);
or U10285 (N_10285,N_43,N_9033);
and U10286 (N_10286,N_4572,N_9540);
or U10287 (N_10287,N_9943,N_1232);
nor U10288 (N_10288,N_1852,N_9687);
and U10289 (N_10289,N_3294,N_3486);
xor U10290 (N_10290,N_4263,N_3968);
nand U10291 (N_10291,N_9711,N_6456);
nor U10292 (N_10292,N_3207,N_5448);
nor U10293 (N_10293,N_9479,N_8817);
nand U10294 (N_10294,N_2576,N_1128);
nand U10295 (N_10295,N_2685,N_4075);
nand U10296 (N_10296,N_7432,N_8966);
or U10297 (N_10297,N_8205,N_1917);
or U10298 (N_10298,N_1457,N_1629);
nor U10299 (N_10299,N_7495,N_3260);
and U10300 (N_10300,N_5069,N_3087);
nor U10301 (N_10301,N_8659,N_7317);
nor U10302 (N_10302,N_7035,N_3265);
nor U10303 (N_10303,N_2374,N_8796);
nand U10304 (N_10304,N_7784,N_8565);
and U10305 (N_10305,N_7047,N_758);
nor U10306 (N_10306,N_3005,N_1421);
and U10307 (N_10307,N_7348,N_1126);
nand U10308 (N_10308,N_2129,N_6140);
and U10309 (N_10309,N_6035,N_4466);
or U10310 (N_10310,N_961,N_1267);
nand U10311 (N_10311,N_5551,N_1864);
and U10312 (N_10312,N_9798,N_1893);
nor U10313 (N_10313,N_6775,N_1311);
or U10314 (N_10314,N_2965,N_6513);
or U10315 (N_10315,N_6871,N_5808);
and U10316 (N_10316,N_8010,N_3920);
nor U10317 (N_10317,N_5525,N_5889);
or U10318 (N_10318,N_7242,N_8864);
and U10319 (N_10319,N_7689,N_852);
nand U10320 (N_10320,N_5141,N_8597);
or U10321 (N_10321,N_4054,N_8271);
nand U10322 (N_10322,N_5768,N_4553);
nand U10323 (N_10323,N_3835,N_5101);
or U10324 (N_10324,N_618,N_517);
and U10325 (N_10325,N_9500,N_9236);
nand U10326 (N_10326,N_7680,N_7732);
or U10327 (N_10327,N_9248,N_1038);
nand U10328 (N_10328,N_6933,N_9690);
and U10329 (N_10329,N_8902,N_5781);
nor U10330 (N_10330,N_7696,N_7541);
and U10331 (N_10331,N_3193,N_5831);
or U10332 (N_10332,N_878,N_4923);
nand U10333 (N_10333,N_2898,N_128);
and U10334 (N_10334,N_1447,N_5660);
nor U10335 (N_10335,N_8609,N_3403);
and U10336 (N_10336,N_1369,N_3785);
nor U10337 (N_10337,N_269,N_7650);
nor U10338 (N_10338,N_7294,N_4063);
or U10339 (N_10339,N_9265,N_5976);
nand U10340 (N_10340,N_9920,N_6464);
nor U10341 (N_10341,N_5878,N_4745);
nor U10342 (N_10342,N_1446,N_3726);
nand U10343 (N_10343,N_617,N_2829);
nand U10344 (N_10344,N_820,N_9979);
and U10345 (N_10345,N_1899,N_6902);
or U10346 (N_10346,N_7086,N_4212);
and U10347 (N_10347,N_6290,N_289);
nand U10348 (N_10348,N_3171,N_1305);
nor U10349 (N_10349,N_7692,N_4406);
nand U10350 (N_10350,N_1749,N_3352);
nor U10351 (N_10351,N_6884,N_4105);
or U10352 (N_10352,N_1194,N_7210);
and U10353 (N_10353,N_1477,N_2456);
nand U10354 (N_10354,N_7895,N_931);
or U10355 (N_10355,N_3478,N_4033);
or U10356 (N_10356,N_8240,N_6527);
and U10357 (N_10357,N_3590,N_3083);
nor U10358 (N_10358,N_4738,N_8983);
nand U10359 (N_10359,N_4790,N_2171);
and U10360 (N_10360,N_4755,N_7153);
and U10361 (N_10361,N_6433,N_4640);
nand U10362 (N_10362,N_9588,N_4925);
nor U10363 (N_10363,N_7156,N_5349);
or U10364 (N_10364,N_5053,N_5931);
or U10365 (N_10365,N_7524,N_9272);
nand U10366 (N_10366,N_248,N_373);
nand U10367 (N_10367,N_298,N_973);
nand U10368 (N_10368,N_4767,N_6348);
and U10369 (N_10369,N_6185,N_1826);
nor U10370 (N_10370,N_1179,N_494);
nand U10371 (N_10371,N_885,N_4955);
nor U10372 (N_10372,N_5149,N_9499);
nor U10373 (N_10373,N_8514,N_4814);
nor U10374 (N_10374,N_6547,N_5625);
or U10375 (N_10375,N_5063,N_7936);
nand U10376 (N_10376,N_3552,N_1443);
nor U10377 (N_10377,N_4463,N_9419);
nor U10378 (N_10378,N_681,N_6112);
or U10379 (N_10379,N_9360,N_8611);
and U10380 (N_10380,N_7379,N_1881);
nand U10381 (N_10381,N_8718,N_2126);
and U10382 (N_10382,N_1079,N_2332);
and U10383 (N_10383,N_1871,N_6194);
nor U10384 (N_10384,N_7257,N_5457);
and U10385 (N_10385,N_724,N_9099);
and U10386 (N_10386,N_1257,N_7446);
or U10387 (N_10387,N_1743,N_9312);
nand U10388 (N_10388,N_410,N_1760);
nand U10389 (N_10389,N_9061,N_4945);
nor U10390 (N_10390,N_1970,N_867);
and U10391 (N_10391,N_7478,N_4286);
nor U10392 (N_10392,N_9309,N_3588);
nand U10393 (N_10393,N_9119,N_5644);
nor U10394 (N_10394,N_7843,N_4775);
and U10395 (N_10395,N_6680,N_2467);
and U10396 (N_10396,N_3563,N_5392);
nor U10397 (N_10397,N_4253,N_3277);
nor U10398 (N_10398,N_5161,N_3230);
nand U10399 (N_10399,N_5065,N_471);
nor U10400 (N_10400,N_5212,N_6381);
and U10401 (N_10401,N_6744,N_6549);
or U10402 (N_10402,N_1392,N_6636);
nor U10403 (N_10403,N_7128,N_6397);
nor U10404 (N_10404,N_6073,N_7397);
nor U10405 (N_10405,N_9206,N_4543);
nand U10406 (N_10406,N_7102,N_4910);
nor U10407 (N_10407,N_8741,N_8862);
nor U10408 (N_10408,N_5918,N_7421);
and U10409 (N_10409,N_2672,N_2891);
nand U10410 (N_10410,N_7525,N_6717);
nand U10411 (N_10411,N_8435,N_5283);
or U10412 (N_10412,N_2561,N_6845);
nand U10413 (N_10413,N_8256,N_7829);
nor U10414 (N_10414,N_7402,N_6687);
nor U10415 (N_10415,N_938,N_2205);
nor U10416 (N_10416,N_2476,N_94);
nand U10417 (N_10417,N_6425,N_7138);
and U10418 (N_10418,N_4402,N_2046);
and U10419 (N_10419,N_7236,N_3520);
nand U10420 (N_10420,N_7863,N_6345);
nor U10421 (N_10421,N_4264,N_5370);
and U10422 (N_10422,N_9826,N_4148);
and U10423 (N_10423,N_4015,N_5344);
nand U10424 (N_10424,N_5582,N_2020);
or U10425 (N_10425,N_160,N_4638);
and U10426 (N_10426,N_3155,N_727);
and U10427 (N_10427,N_2922,N_6400);
nor U10428 (N_10428,N_9703,N_1765);
or U10429 (N_10429,N_1434,N_2372);
and U10430 (N_10430,N_470,N_8289);
nand U10431 (N_10431,N_107,N_6106);
nor U10432 (N_10432,N_8144,N_7503);
nand U10433 (N_10433,N_6776,N_2792);
and U10434 (N_10434,N_125,N_8679);
and U10435 (N_10435,N_4116,N_4571);
nand U10436 (N_10436,N_2940,N_9630);
nor U10437 (N_10437,N_809,N_1817);
or U10438 (N_10438,N_6044,N_9037);
or U10439 (N_10439,N_7116,N_2073);
nor U10440 (N_10440,N_8737,N_1073);
nand U10441 (N_10441,N_4107,N_6664);
or U10442 (N_10442,N_369,N_2710);
nor U10443 (N_10443,N_8575,N_8587);
nor U10444 (N_10444,N_8959,N_8103);
or U10445 (N_10445,N_8628,N_6158);
and U10446 (N_10446,N_4375,N_329);
nor U10447 (N_10447,N_9696,N_9152);
nor U10448 (N_10448,N_4403,N_3956);
and U10449 (N_10449,N_7970,N_1780);
and U10450 (N_10450,N_3614,N_623);
nand U10451 (N_10451,N_8525,N_2019);
nor U10452 (N_10452,N_9392,N_5012);
or U10453 (N_10453,N_6439,N_2966);
and U10454 (N_10454,N_960,N_1512);
nor U10455 (N_10455,N_7701,N_4272);
or U10456 (N_10456,N_8823,N_2927);
nand U10457 (N_10457,N_7034,N_2942);
or U10458 (N_10458,N_7021,N_7975);
nand U10459 (N_10459,N_9714,N_22);
nor U10460 (N_10460,N_9051,N_9086);
nand U10461 (N_10461,N_2596,N_8694);
and U10462 (N_10462,N_7756,N_6030);
or U10463 (N_10463,N_2715,N_8007);
and U10464 (N_10464,N_6907,N_388);
nor U10465 (N_10465,N_3108,N_2844);
and U10466 (N_10466,N_4090,N_9989);
nand U10467 (N_10467,N_6545,N_4777);
nand U10468 (N_10468,N_7033,N_4762);
nor U10469 (N_10469,N_7468,N_1460);
nand U10470 (N_10470,N_4992,N_8539);
nand U10471 (N_10471,N_4785,N_6132);
nand U10472 (N_10472,N_974,N_3784);
nand U10473 (N_10473,N_5749,N_964);
nand U10474 (N_10474,N_7315,N_1657);
or U10475 (N_10475,N_4848,N_4897);
nand U10476 (N_10476,N_7061,N_9125);
xnor U10477 (N_10477,N_7926,N_9651);
or U10478 (N_10478,N_6765,N_7905);
and U10479 (N_10479,N_7551,N_4467);
xor U10480 (N_10480,N_6404,N_8974);
and U10481 (N_10481,N_2648,N_3741);
nor U10482 (N_10482,N_3594,N_2252);
nor U10483 (N_10483,N_9462,N_4325);
nor U10484 (N_10484,N_3703,N_8762);
nand U10485 (N_10485,N_7601,N_3013);
and U10486 (N_10486,N_7423,N_208);
or U10487 (N_10487,N_8170,N_7207);
and U10488 (N_10488,N_2273,N_9919);
nand U10489 (N_10489,N_4960,N_3582);
nor U10490 (N_10490,N_7469,N_1068);
nor U10491 (N_10491,N_8360,N_4670);
nor U10492 (N_10492,N_1674,N_1520);
nand U10493 (N_10493,N_9103,N_6550);
and U10494 (N_10494,N_5734,N_1468);
nand U10495 (N_10495,N_8850,N_3172);
nand U10496 (N_10496,N_6681,N_9496);
or U10497 (N_10497,N_5470,N_1025);
or U10498 (N_10498,N_2568,N_5692);
nand U10499 (N_10499,N_1588,N_343);
and U10500 (N_10500,N_4784,N_9169);
or U10501 (N_10501,N_957,N_8162);
xnor U10502 (N_10502,N_2845,N_9283);
nor U10503 (N_10503,N_4899,N_6922);
nor U10504 (N_10504,N_9179,N_9408);
nand U10505 (N_10505,N_8607,N_5243);
nand U10506 (N_10506,N_115,N_5513);
and U10507 (N_10507,N_6941,N_2719);
nor U10508 (N_10508,N_4340,N_2324);
and U10509 (N_10509,N_61,N_7072);
nand U10510 (N_10510,N_5292,N_3395);
or U10511 (N_10511,N_3789,N_9250);
nor U10512 (N_10512,N_9182,N_8638);
or U10513 (N_10513,N_9207,N_287);
and U10514 (N_10514,N_3580,N_7890);
and U10515 (N_10515,N_6446,N_3140);
nand U10516 (N_10516,N_4528,N_8941);
or U10517 (N_10517,N_8182,N_8557);
nor U10518 (N_10518,N_6522,N_266);
and U10519 (N_10519,N_6234,N_1323);
and U10520 (N_10520,N_3947,N_4172);
nor U10521 (N_10521,N_7586,N_3423);
and U10522 (N_10522,N_8138,N_3376);
or U10523 (N_10523,N_7806,N_5121);
nor U10524 (N_10524,N_4258,N_656);
or U10525 (N_10525,N_274,N_12);
and U10526 (N_10526,N_3906,N_2030);
and U10527 (N_10527,N_7383,N_2039);
or U10528 (N_10528,N_2928,N_8125);
or U10529 (N_10529,N_1004,N_6912);
nand U10530 (N_10530,N_5740,N_7231);
nand U10531 (N_10531,N_5957,N_1422);
or U10532 (N_10532,N_1003,N_4482);
nand U10533 (N_10533,N_8865,N_1951);
nand U10534 (N_10534,N_3313,N_1173);
nor U10535 (N_10535,N_5111,N_301);
and U10536 (N_10536,N_2331,N_104);
and U10537 (N_10537,N_3760,N_9802);
and U10538 (N_10538,N_2455,N_9464);
nand U10539 (N_10539,N_4496,N_9286);
or U10540 (N_10540,N_4880,N_9968);
and U10541 (N_10541,N_1730,N_584);
and U10542 (N_10542,N_9672,N_1012);
and U10543 (N_10543,N_814,N_1391);
nor U10544 (N_10544,N_7309,N_5265);
and U10545 (N_10545,N_730,N_7493);
and U10546 (N_10546,N_7595,N_8037);
or U10547 (N_10547,N_5220,N_2274);
or U10548 (N_10548,N_2156,N_1902);
nor U10549 (N_10549,N_2475,N_8534);
nand U10550 (N_10550,N_5126,N_4053);
nand U10551 (N_10551,N_1719,N_4676);
and U10552 (N_10552,N_6913,N_7591);
and U10553 (N_10553,N_7191,N_4026);
and U10554 (N_10554,N_5184,N_682);
or U10555 (N_10555,N_3264,N_9321);
and U10556 (N_10556,N_6378,N_6874);
nor U10557 (N_10557,N_8361,N_6490);
or U10558 (N_10558,N_6377,N_3324);
or U10559 (N_10559,N_2155,N_992);
nor U10560 (N_10560,N_4803,N_5667);
nor U10561 (N_10561,N_1397,N_483);
nor U10562 (N_10562,N_8302,N_7668);
nor U10563 (N_10563,N_3330,N_5862);
nor U10564 (N_10564,N_6063,N_3769);
or U10565 (N_10565,N_6894,N_1284);
and U10566 (N_10566,N_2123,N_8511);
nand U10567 (N_10567,N_224,N_3924);
or U10568 (N_10568,N_8386,N_9063);
nor U10569 (N_10569,N_7888,N_7173);
nand U10570 (N_10570,N_8608,N_2502);
nor U10571 (N_10571,N_3672,N_9740);
or U10572 (N_10572,N_8591,N_6782);
nor U10573 (N_10573,N_6835,N_4713);
nand U10574 (N_10574,N_64,N_8826);
or U10575 (N_10575,N_2678,N_9847);
nand U10576 (N_10576,N_3970,N_7535);
nand U10577 (N_10577,N_2833,N_9602);
nand U10578 (N_10578,N_9577,N_1611);
and U10579 (N_10579,N_4120,N_5516);
or U10580 (N_10580,N_4617,N_7947);
nor U10581 (N_10581,N_7202,N_8433);
and U10582 (N_10582,N_4014,N_606);
nor U10583 (N_10583,N_1651,N_8695);
nand U10584 (N_10584,N_6660,N_2651);
or U10585 (N_10585,N_2508,N_7821);
or U10586 (N_10586,N_2996,N_7200);
nand U10587 (N_10587,N_7564,N_7780);
and U10588 (N_10588,N_1291,N_4892);
or U10589 (N_10589,N_3551,N_1277);
nor U10590 (N_10590,N_5894,N_1906);
nor U10591 (N_10591,N_2338,N_8757);
nand U10592 (N_10592,N_6892,N_5597);
nor U10593 (N_10593,N_8670,N_7725);
and U10594 (N_10594,N_5253,N_8920);
nor U10595 (N_10595,N_8141,N_6659);
nor U10596 (N_10596,N_4509,N_1110);
or U10597 (N_10597,N_2603,N_5760);
or U10598 (N_10598,N_8485,N_347);
or U10599 (N_10599,N_6152,N_4294);
or U10600 (N_10600,N_9004,N_2828);
nand U10601 (N_10601,N_7655,N_9411);
nor U10602 (N_10602,N_1758,N_3900);
nand U10603 (N_10603,N_4760,N_491);
nand U10604 (N_10604,N_156,N_5);
nor U10605 (N_10605,N_6560,N_3394);
and U10606 (N_10606,N_8190,N_8293);
nor U10607 (N_10607,N_2018,N_4614);
nand U10608 (N_10608,N_9071,N_6581);
or U10609 (N_10609,N_6533,N_5656);
nor U10610 (N_10610,N_3450,N_321);
or U10611 (N_10611,N_6141,N_5681);
or U10612 (N_10612,N_2569,N_920);
and U10613 (N_10613,N_9878,N_7966);
nor U10614 (N_10614,N_9027,N_7550);
nand U10615 (N_10615,N_7007,N_8142);
and U10616 (N_10616,N_940,N_1335);
nand U10617 (N_10617,N_2283,N_1218);
nor U10618 (N_10618,N_9549,N_3660);
nand U10619 (N_10619,N_9014,N_2975);
nand U10620 (N_10620,N_3119,N_2243);
and U10621 (N_10621,N_6877,N_1247);
and U10622 (N_10622,N_6619,N_3032);
or U10623 (N_10623,N_2705,N_3624);
nor U10624 (N_10624,N_645,N_5007);
and U10625 (N_10625,N_1793,N_1887);
nand U10626 (N_10626,N_4743,N_6773);
nand U10627 (N_10627,N_1524,N_9334);
nor U10628 (N_10628,N_5884,N_8931);
nand U10629 (N_10629,N_9897,N_7229);
xnor U10630 (N_10630,N_3386,N_1045);
and U10631 (N_10631,N_2169,N_5811);
or U10632 (N_10632,N_2451,N_82);
nand U10633 (N_10633,N_9192,N_6001);
and U10634 (N_10634,N_7855,N_3561);
and U10635 (N_10635,N_3761,N_9974);
or U10636 (N_10636,N_3491,N_3068);
and U10637 (N_10637,N_172,N_9751);
and U10638 (N_10638,N_614,N_4683);
nor U10639 (N_10639,N_8768,N_6186);
nor U10640 (N_10640,N_8674,N_1568);
and U10641 (N_10641,N_9395,N_1269);
xor U10642 (N_10642,N_4595,N_3744);
nand U10643 (N_10643,N_891,N_7927);
nor U10644 (N_10644,N_2325,N_5505);
xor U10645 (N_10645,N_2794,N_1227);
nand U10646 (N_10646,N_6211,N_4404);
nor U10647 (N_10647,N_5881,N_3272);
and U10648 (N_10648,N_4031,N_2092);
and U10649 (N_10649,N_2798,N_1181);
and U10650 (N_10650,N_236,N_2145);
nand U10651 (N_10651,N_7358,N_5140);
nand U10652 (N_10652,N_1774,N_5869);
or U10653 (N_10653,N_9535,N_8031);
or U10654 (N_10654,N_563,N_880);
and U10655 (N_10655,N_8518,N_808);
nand U10656 (N_10656,N_1818,N_1159);
nand U10657 (N_10657,N_7850,N_8301);
and U10658 (N_10658,N_6357,N_2774);
nor U10659 (N_10659,N_9723,N_7730);
nor U10660 (N_10660,N_5793,N_5250);
or U10661 (N_10661,N_7112,N_2288);
or U10662 (N_10662,N_1129,N_5295);
nor U10663 (N_10663,N_4020,N_1116);
nand U10664 (N_10664,N_6585,N_9050);
nand U10665 (N_10665,N_7611,N_2431);
nor U10666 (N_10666,N_7506,N_8029);
and U10667 (N_10667,N_2284,N_1195);
or U10668 (N_10668,N_3960,N_4797);
nor U10669 (N_10669,N_5591,N_4536);
nor U10670 (N_10670,N_2684,N_567);
or U10671 (N_10671,N_5710,N_8310);
or U10672 (N_10672,N_4146,N_8200);
nand U10673 (N_10673,N_2861,N_3174);
nand U10674 (N_10674,N_6834,N_7254);
or U10675 (N_10675,N_7406,N_2017);
and U10676 (N_10676,N_2723,N_3869);
nor U10677 (N_10677,N_1829,N_3778);
and U10678 (N_10678,N_1016,N_728);
and U10679 (N_10679,N_6244,N_9870);
or U10680 (N_10680,N_4578,N_3825);
nor U10681 (N_10681,N_6324,N_1506);
or U10682 (N_10682,N_732,N_7059);
nand U10683 (N_10683,N_4080,N_2742);
nor U10684 (N_10684,N_1693,N_6333);
xnor U10685 (N_10685,N_7709,N_5443);
nand U10686 (N_10686,N_4426,N_5416);
nand U10687 (N_10687,N_6153,N_3023);
and U10688 (N_10688,N_4168,N_5491);
nand U10689 (N_10689,N_6256,N_8483);
or U10690 (N_10690,N_5753,N_9351);
and U10691 (N_10691,N_5242,N_1880);
nor U10692 (N_10692,N_2490,N_1930);
and U10693 (N_10693,N_6354,N_1196);
nand U10694 (N_10694,N_7934,N_7750);
nand U10695 (N_10695,N_4703,N_2085);
nor U10696 (N_10696,N_1620,N_8548);
nor U10697 (N_10697,N_4641,N_3041);
nor U10698 (N_10698,N_1428,N_1807);
and U10699 (N_10699,N_2353,N_1385);
nand U10700 (N_10700,N_5746,N_3198);
and U10701 (N_10701,N_2076,N_5281);
or U10702 (N_10702,N_6491,N_9226);
or U10703 (N_10703,N_9041,N_2873);
or U10704 (N_10704,N_5228,N_8236);
nand U10705 (N_10705,N_7043,N_385);
nor U10706 (N_10706,N_5045,N_4235);
nor U10707 (N_10707,N_9454,N_1455);
nand U10708 (N_10708,N_3780,N_4163);
nor U10709 (N_10709,N_7861,N_51);
and U10710 (N_10710,N_212,N_3164);
or U10711 (N_10711,N_4898,N_9914);
nor U10712 (N_10712,N_1485,N_7919);
or U10713 (N_10713,N_9777,N_4042);
or U10714 (N_10714,N_2408,N_6707);
and U10715 (N_10715,N_6447,N_8745);
or U10716 (N_10716,N_5536,N_5060);
and U10717 (N_10717,N_6694,N_6281);
and U10718 (N_10718,N_9385,N_3470);
nor U10719 (N_10719,N_9726,N_678);
nand U10720 (N_10720,N_4448,N_9966);
and U10721 (N_10721,N_2669,N_4937);
nor U10722 (N_10722,N_7628,N_6116);
and U10723 (N_10723,N_3154,N_2810);
or U10724 (N_10724,N_1008,N_6810);
or U10725 (N_10725,N_7263,N_555);
nand U10726 (N_10726,N_4355,N_8592);
and U10727 (N_10727,N_7765,N_2276);
and U10728 (N_10728,N_7455,N_4711);
nor U10729 (N_10729,N_7704,N_7620);
and U10730 (N_10730,N_9410,N_7266);
and U10731 (N_10731,N_8971,N_14);
and U10732 (N_10732,N_3467,N_201);
nand U10733 (N_10733,N_3142,N_7090);
and U10734 (N_10734,N_7101,N_8276);
and U10735 (N_10735,N_1442,N_2158);
nor U10736 (N_10736,N_8743,N_1590);
or U10737 (N_10737,N_2851,N_3679);
nand U10738 (N_10738,N_6724,N_6650);
nor U10739 (N_10739,N_3527,N_1417);
nand U10740 (N_10740,N_8975,N_2984);
nand U10741 (N_10741,N_6201,N_1950);
nor U10742 (N_10742,N_8385,N_3369);
or U10743 (N_10743,N_6268,N_4194);
nor U10744 (N_10744,N_4187,N_3818);
and U10745 (N_10745,N_9839,N_4096);
nand U10746 (N_10746,N_9463,N_2376);
nand U10747 (N_10747,N_6175,N_6095);
nor U10748 (N_10748,N_8430,N_6863);
and U10749 (N_10749,N_2788,N_234);
and U10750 (N_10750,N_2172,N_3697);
and U10751 (N_10751,N_863,N_1217);
nor U10752 (N_10752,N_7482,N_530);
and U10753 (N_10753,N_868,N_6146);
and U10754 (N_10754,N_4747,N_378);
nor U10755 (N_10755,N_219,N_6356);
nor U10756 (N_10756,N_2834,N_5695);
or U10757 (N_10757,N_6349,N_2977);
nor U10758 (N_10758,N_2791,N_5226);
nand U10759 (N_10759,N_9812,N_4444);
and U10760 (N_10760,N_5278,N_6482);
and U10761 (N_10761,N_2237,N_8336);
and U10762 (N_10762,N_5636,N_9459);
and U10763 (N_10763,N_1259,N_7920);
nand U10764 (N_10764,N_8723,N_7441);
nand U10765 (N_10765,N_3454,N_5802);
or U10766 (N_10766,N_3229,N_8786);
nor U10767 (N_10767,N_6239,N_4408);
or U10768 (N_10768,N_4849,N_7133);
and U10769 (N_10769,N_5599,N_8115);
nand U10770 (N_10770,N_3524,N_2783);
nor U10771 (N_10771,N_572,N_894);
or U10772 (N_10772,N_4099,N_3565);
and U10773 (N_10773,N_4245,N_5908);
and U10774 (N_10774,N_6520,N_1550);
or U10775 (N_10775,N_9853,N_738);
and U10776 (N_10776,N_8779,N_2677);
and U10777 (N_10777,N_3156,N_2607);
or U10778 (N_10778,N_9401,N_6860);
and U10779 (N_10779,N_9541,N_699);
and U10780 (N_10780,N_7373,N_2212);
and U10781 (N_10781,N_6413,N_9543);
nand U10782 (N_10782,N_9811,N_3965);
and U10783 (N_10783,N_2207,N_5251);
and U10784 (N_10784,N_9023,N_4724);
nand U10785 (N_10785,N_7769,N_6405);
nor U10786 (N_10786,N_6069,N_8239);
nand U10787 (N_10787,N_8707,N_5680);
or U10788 (N_10788,N_440,N_4521);
or U10789 (N_10789,N_1119,N_4596);
and U10790 (N_10790,N_7442,N_4786);
nor U10791 (N_10791,N_2343,N_5308);
or U10792 (N_10792,N_3271,N_249);
nand U10793 (N_10793,N_1988,N_691);
nand U10794 (N_10794,N_5257,N_4262);
nor U10795 (N_10795,N_7448,N_4922);
or U10796 (N_10796,N_6219,N_2356);
or U10797 (N_10797,N_4661,N_7416);
and U10798 (N_10798,N_9925,N_7954);
or U10799 (N_10799,N_8545,N_3516);
and U10800 (N_10800,N_2464,N_4526);
or U10801 (N_10801,N_7994,N_3421);
nor U10802 (N_10802,N_3261,N_2167);
and U10803 (N_10803,N_9838,N_7456);
and U10804 (N_10804,N_1345,N_8663);
and U10805 (N_10805,N_3750,N_4827);
and U10806 (N_10806,N_7181,N_9139);
or U10807 (N_10807,N_1155,N_3182);
and U10808 (N_10808,N_3705,N_5473);
or U10809 (N_10809,N_978,N_2777);
nor U10810 (N_10810,N_4706,N_4322);
nor U10811 (N_10811,N_2667,N_8306);
nand U10812 (N_10812,N_4232,N_6319);
nor U10813 (N_10813,N_3384,N_2986);
and U10814 (N_10814,N_995,N_769);
and U10815 (N_10815,N_1384,N_3978);
and U10816 (N_10816,N_4733,N_8542);
nor U10817 (N_10817,N_5403,N_1071);
nand U10818 (N_10818,N_8152,N_6947);
or U10819 (N_10819,N_8690,N_8424);
nand U10820 (N_10820,N_4574,N_895);
or U10821 (N_10821,N_9895,N_3425);
nor U10822 (N_10822,N_5666,N_4494);
nand U10823 (N_10823,N_8399,N_1890);
and U10824 (N_10824,N_760,N_8651);
or U10825 (N_10825,N_317,N_431);
or U10826 (N_10826,N_9623,N_2062);
nor U10827 (N_10827,N_1297,N_5334);
and U10828 (N_10828,N_3233,N_4009);
or U10829 (N_10829,N_7260,N_4289);
or U10830 (N_10830,N_1612,N_7758);
or U10831 (N_10831,N_3308,N_8569);
nor U10832 (N_10832,N_4846,N_9135);
and U10833 (N_10833,N_1936,N_4453);
nand U10834 (N_10834,N_8896,N_8305);
nor U10835 (N_10835,N_5890,N_3460);
and U10836 (N_10836,N_5986,N_2793);
nand U10837 (N_10837,N_105,N_6238);
nand U10838 (N_10838,N_7328,N_8555);
nor U10839 (N_10839,N_937,N_1165);
nor U10840 (N_10840,N_7570,N_6133);
or U10841 (N_10841,N_1860,N_2894);
and U10842 (N_10842,N_7723,N_4592);
nor U10843 (N_10843,N_3284,N_800);
and U10844 (N_10844,N_1533,N_7427);
nand U10845 (N_10845,N_6122,N_6019);
nor U10846 (N_10846,N_4963,N_3278);
nand U10847 (N_10847,N_3881,N_9380);
or U10848 (N_10848,N_5422,N_9261);
nor U10849 (N_10849,N_7657,N_3959);
and U10850 (N_10850,N_1088,N_8325);
or U10851 (N_10851,N_1011,N_1676);
nand U10852 (N_10852,N_16,N_9378);
nor U10853 (N_10853,N_8149,N_9960);
nor U10854 (N_10854,N_7995,N_680);
nor U10855 (N_10855,N_7589,N_4823);
nor U10856 (N_10856,N_173,N_5398);
and U10857 (N_10857,N_4844,N_2468);
or U10858 (N_10858,N_3890,N_2142);
or U10859 (N_10859,N_2529,N_3871);
nor U10860 (N_10860,N_2881,N_3700);
and U10861 (N_10861,N_3722,N_5247);
nand U10862 (N_10862,N_6007,N_9057);
nor U10863 (N_10863,N_2647,N_1592);
or U10864 (N_10864,N_8268,N_3584);
nand U10865 (N_10865,N_6004,N_8749);
or U10866 (N_10866,N_3713,N_1941);
nor U10867 (N_10867,N_1925,N_6881);
nand U10868 (N_10868,N_8673,N_4067);
nor U10869 (N_10869,N_8283,N_3139);
and U10870 (N_10870,N_3942,N_8612);
or U10871 (N_10871,N_3922,N_9268);
nand U10872 (N_10872,N_2595,N_6957);
nand U10873 (N_10873,N_3531,N_8198);
nand U10874 (N_10874,N_860,N_1557);
or U10875 (N_10875,N_657,N_792);
nor U10876 (N_10876,N_4214,N_9932);
nand U10877 (N_10877,N_8314,N_8078);
or U10878 (N_10878,N_7074,N_1414);
and U10879 (N_10879,N_7004,N_6293);
nor U10880 (N_10880,N_5488,N_4074);
or U10881 (N_10881,N_3383,N_8778);
nand U10882 (N_10882,N_6737,N_811);
nor U10883 (N_10883,N_4499,N_2297);
nand U10884 (N_10884,N_424,N_6111);
and U10885 (N_10885,N_6736,N_2806);
nor U10886 (N_10886,N_4410,N_2385);
or U10887 (N_10887,N_7248,N_9075);
nand U10888 (N_10888,N_6229,N_6396);
and U10889 (N_10889,N_6005,N_2826);
nand U10890 (N_10890,N_2176,N_1961);
and U10891 (N_10891,N_2724,N_4667);
or U10892 (N_10892,N_9359,N_1853);
or U10893 (N_10893,N_8047,N_6025);
and U10894 (N_10894,N_6709,N_379);
and U10895 (N_10895,N_3134,N_8879);
nand U10896 (N_10896,N_4307,N_9736);
and U10897 (N_10897,N_8364,N_579);
nand U10898 (N_10898,N_114,N_9197);
or U10899 (N_10899,N_2757,N_5329);
and U10900 (N_10900,N_136,N_3519);
and U10901 (N_10901,N_1147,N_4392);
xnor U10902 (N_10902,N_7759,N_8024);
nand U10903 (N_10903,N_8134,N_1789);
nor U10904 (N_10904,N_2188,N_5452);
and U10905 (N_10905,N_6109,N_7556);
or U10906 (N_10906,N_8649,N_6657);
and U10907 (N_10907,N_7147,N_3512);
or U10908 (N_10908,N_8881,N_7845);
or U10909 (N_10909,N_5674,N_2862);
nand U10910 (N_10910,N_271,N_3607);
and U10911 (N_10911,N_2541,N_9466);
or U10912 (N_10912,N_4860,N_4435);
nand U10913 (N_10913,N_1794,N_5301);
nor U10914 (N_10914,N_6176,N_5497);
or U10915 (N_10915,N_8522,N_1190);
and U10916 (N_10916,N_4774,N_9631);
and U10917 (N_10917,N_1085,N_7578);
xor U10918 (N_10918,N_5097,N_8877);
nor U10919 (N_10919,N_4851,N_2230);
or U10920 (N_10920,N_9081,N_4057);
or U10921 (N_10921,N_226,N_1798);
or U10922 (N_10922,N_9773,N_5279);
nor U10923 (N_10923,N_8228,N_7302);
nand U10924 (N_10924,N_1816,N_7604);
nor U10925 (N_10925,N_1061,N_157);
or U10926 (N_10926,N_3323,N_9430);
or U10927 (N_10927,N_1990,N_3566);
and U10928 (N_10928,N_7337,N_4674);
and U10929 (N_10929,N_7621,N_1234);
and U10930 (N_10930,N_3322,N_4792);
or U10931 (N_10931,N_5444,N_2389);
nor U10932 (N_10932,N_151,N_2056);
and U10933 (N_10933,N_7395,N_210);
and U10934 (N_10934,N_1876,N_8897);
nand U10935 (N_10935,N_5464,N_9217);
nor U10936 (N_10936,N_5595,N_4729);
nor U10937 (N_10937,N_1584,N_6984);
nor U10938 (N_10938,N_4476,N_4045);
and U10939 (N_10939,N_8925,N_9011);
and U10940 (N_10940,N_6953,N_6537);
or U10941 (N_10941,N_3197,N_5888);
nor U10942 (N_10942,N_9418,N_8381);
nor U10943 (N_10943,N_1252,N_2823);
or U10944 (N_10944,N_5380,N_1614);
nor U10945 (N_10945,N_9525,N_5554);
and U10946 (N_10946,N_8023,N_915);
nand U10947 (N_10947,N_7027,N_9007);
nand U10948 (N_10948,N_2285,N_3932);
nand U10949 (N_10949,N_4291,N_4003);
nand U10950 (N_10950,N_4904,N_7637);
or U10951 (N_10951,N_9815,N_1525);
nand U10952 (N_10952,N_7582,N_8372);
nor U10953 (N_10953,N_3504,N_5107);
or U10954 (N_10954,N_7558,N_666);
and U10955 (N_10955,N_7447,N_4139);
or U10956 (N_10956,N_3034,N_901);
or U10957 (N_10957,N_4736,N_9439);
nand U10958 (N_10958,N_3781,N_8121);
and U10959 (N_10959,N_1435,N_5098);
nor U10960 (N_10960,N_3694,N_2355);
or U10961 (N_10961,N_6828,N_1208);
or U10962 (N_10962,N_7244,N_8475);
or U10963 (N_10963,N_9953,N_9854);
or U10964 (N_10964,N_9567,N_858);
or U10965 (N_10965,N_7946,N_2027);
or U10966 (N_10966,N_232,N_2381);
nand U10967 (N_10967,N_3641,N_9614);
and U10968 (N_10968,N_6483,N_7795);
nand U10969 (N_10969,N_3100,N_4847);
nand U10970 (N_10970,N_4025,N_6163);
and U10971 (N_10971,N_7238,N_7470);
nand U10972 (N_10972,N_8393,N_6805);
or U10973 (N_10973,N_4659,N_2546);
xor U10974 (N_10974,N_1834,N_9313);
nor U10975 (N_10975,N_2657,N_8567);
and U10976 (N_10976,N_7433,N_4579);
and U10977 (N_10977,N_8523,N_9524);
or U10978 (N_10978,N_7548,N_7891);
nor U10979 (N_10979,N_9291,N_568);
nor U10980 (N_10980,N_9142,N_3437);
nand U10981 (N_10981,N_405,N_5272);
and U10982 (N_10982,N_8400,N_6395);
or U10983 (N_10983,N_3338,N_4331);
and U10984 (N_10984,N_463,N_7008);
or U10985 (N_10985,N_9376,N_9480);
and U10986 (N_10986,N_1575,N_5728);
nor U10987 (N_10987,N_9884,N_8835);
and U10988 (N_10988,N_6986,N_7196);
nand U10989 (N_10989,N_8185,N_627);
or U10990 (N_10990,N_3609,N_4489);
nand U10991 (N_10991,N_6448,N_2217);
nand U10992 (N_10992,N_5330,N_3521);
or U10993 (N_10993,N_764,N_6382);
and U10994 (N_10994,N_7796,N_6600);
and U10995 (N_10995,N_7836,N_3355);
nand U10996 (N_10996,N_4712,N_4292);
nand U10997 (N_10997,N_3997,N_635);
nand U10998 (N_10998,N_9680,N_641);
nor U10999 (N_10999,N_4400,N_9422);
nor U11000 (N_11000,N_2183,N_5241);
and U11001 (N_11001,N_4385,N_7807);
nand U11002 (N_11002,N_6120,N_9328);
or U11003 (N_11003,N_3792,N_2269);
or U11004 (N_11004,N_280,N_8951);
nor U11005 (N_11005,N_9778,N_5179);
and U11006 (N_11006,N_5752,N_4030);
nor U11007 (N_11007,N_3431,N_2712);
nand U11008 (N_11008,N_6243,N_5756);
or U11009 (N_11009,N_9388,N_6391);
nand U11010 (N_11010,N_6173,N_823);
and U11011 (N_11011,N_8546,N_1006);
nor U11012 (N_11012,N_5051,N_2368);
and U11013 (N_11013,N_1992,N_7259);
and U11014 (N_11014,N_8801,N_1288);
or U11015 (N_11015,N_1666,N_988);
nand U11016 (N_11016,N_8861,N_9306);
nand U11017 (N_11017,N_5934,N_3245);
or U11018 (N_11018,N_7815,N_5920);
nor U11019 (N_11019,N_9132,N_8206);
or U11020 (N_11020,N_4005,N_9846);
or U11021 (N_11021,N_4123,N_5418);
and U11022 (N_11022,N_3966,N_6003);
and U11023 (N_11023,N_6963,N_8631);
nor U11024 (N_11024,N_9221,N_8080);
nand U11025 (N_11025,N_9367,N_4227);
or U11026 (N_11026,N_4637,N_2148);
and U11027 (N_11027,N_2658,N_95);
and U11028 (N_11028,N_1364,N_4497);
and U11029 (N_11029,N_1296,N_1256);
xnor U11030 (N_11030,N_790,N_4604);
and U11031 (N_11031,N_270,N_3873);
nand U11032 (N_11032,N_8451,N_779);
nor U11033 (N_11033,N_5154,N_5099);
nor U11034 (N_11034,N_7355,N_5487);
nand U11035 (N_11035,N_9899,N_9461);
or U11036 (N_11036,N_6427,N_8627);
and U11037 (N_11037,N_196,N_3575);
nand U11038 (N_11038,N_511,N_1359);
nand U11039 (N_11039,N_3634,N_7820);
nor U11040 (N_11040,N_2619,N_5714);
and U11041 (N_11041,N_3640,N_8193);
or U11042 (N_11042,N_6691,N_8445);
nand U11043 (N_11043,N_7296,N_3885);
nand U11044 (N_11044,N_4383,N_9818);
or U11045 (N_11045,N_6751,N_9095);
or U11046 (N_11046,N_9149,N_6720);
nor U11047 (N_11047,N_3256,N_1532);
nor U11048 (N_11048,N_2329,N_4302);
and U11049 (N_11049,N_8637,N_673);
and U11050 (N_11050,N_3733,N_2366);
nand U11051 (N_11051,N_2421,N_4062);
nand U11052 (N_11052,N_1642,N_364);
nor U11053 (N_11053,N_7399,N_6070);
or U11054 (N_11054,N_9905,N_3685);
nor U11055 (N_11055,N_5829,N_8000);
nand U11056 (N_11056,N_946,N_2175);
nor U11057 (N_11057,N_6309,N_8515);
or U11058 (N_11058,N_1042,N_2443);
nand U11059 (N_11059,N_4461,N_9803);
or U11060 (N_11060,N_6529,N_8571);
nor U11061 (N_11061,N_4798,N_4815);
nand U11062 (N_11062,N_1909,N_5366);
or U11063 (N_11063,N_4171,N_6384);
and U11064 (N_11064,N_1105,N_9621);
and U11065 (N_11065,N_1643,N_1800);
or U11066 (N_11066,N_9918,N_7234);
nor U11067 (N_11067,N_7720,N_5635);
nor U11068 (N_11068,N_8,N_4916);
nor U11069 (N_11069,N_2162,N_998);
and U11070 (N_11070,N_6075,N_9731);
nand U11071 (N_11071,N_835,N_4918);
or U11072 (N_11072,N_8341,N_6692);
nand U11073 (N_11073,N_6516,N_1432);
nand U11074 (N_11074,N_6943,N_8488);
nor U11075 (N_11075,N_4842,N_6221);
or U11076 (N_11076,N_5198,N_3078);
nor U11077 (N_11077,N_7943,N_6002);
nand U11078 (N_11078,N_719,N_2253);
nand U11079 (N_11079,N_6642,N_6499);
nand U11080 (N_11080,N_5568,N_4889);
or U11081 (N_11081,N_448,N_4312);
nor U11082 (N_11082,N_5984,N_4246);
nor U11083 (N_11083,N_2817,N_9111);
or U11084 (N_11084,N_2318,N_3014);
or U11085 (N_11085,N_6034,N_8910);
and U11086 (N_11086,N_7278,N_6833);
and U11087 (N_11087,N_518,N_2305);
and U11088 (N_11088,N_7776,N_5804);
and U11089 (N_11089,N_4649,N_2775);
or U11090 (N_11090,N_9532,N_2812);
or U11091 (N_11091,N_906,N_2038);
nand U11092 (N_11092,N_4064,N_4236);
and U11093 (N_11093,N_240,N_7949);
or U11094 (N_11094,N_2417,N_2540);
nor U11095 (N_11095,N_8120,N_4095);
nand U11096 (N_11096,N_7318,N_9356);
nand U11097 (N_11097,N_7786,N_6506);
and U11098 (N_11098,N_7638,N_1837);
or U11099 (N_11099,N_2052,N_5639);
or U11100 (N_11100,N_7942,N_7372);
and U11101 (N_11101,N_2543,N_1519);
or U11102 (N_11102,N_9603,N_7099);
or U11103 (N_11103,N_2888,N_4352);
nand U11104 (N_11104,N_8330,N_7676);
nor U11105 (N_11105,N_4993,N_9759);
and U11106 (N_11106,N_111,N_2197);
or U11107 (N_11107,N_3476,N_3046);
and U11108 (N_11108,N_9589,N_707);
or U11109 (N_11109,N_844,N_7477);
and U11110 (N_11110,N_1795,N_1874);
nor U11111 (N_11111,N_8374,N_1582);
or U11112 (N_11112,N_8498,N_3783);
or U11113 (N_11113,N_9012,N_7169);
and U11114 (N_11114,N_631,N_9214);
nand U11115 (N_11115,N_2360,N_1728);
nor U11116 (N_11116,N_5172,N_1790);
or U11117 (N_11117,N_7343,N_4396);
nand U11118 (N_11118,N_3573,N_8280);
nand U11119 (N_11119,N_9861,N_8493);
or U11120 (N_11120,N_3490,N_7106);
nand U11121 (N_11121,N_445,N_5912);
or U11122 (N_11122,N_1975,N_8561);
nand U11123 (N_11123,N_4932,N_9653);
or U11124 (N_11124,N_4092,N_4582);
nand U11125 (N_11125,N_8836,N_159);
xor U11126 (N_11126,N_8815,N_7623);
and U11127 (N_11127,N_2799,N_2729);
or U11128 (N_11128,N_3077,N_4293);
or U11129 (N_11129,N_8763,N_6126);
nor U11130 (N_11130,N_3712,N_7262);
nor U11131 (N_11131,N_2250,N_7011);
nand U11132 (N_11132,N_3951,N_7220);
nand U11133 (N_11133,N_6327,N_9144);
and U11134 (N_11134,N_8822,N_9730);
or U11135 (N_11135,N_5983,N_1782);
or U11136 (N_11136,N_4906,N_2901);
or U11137 (N_11137,N_8787,N_6453);
and U11138 (N_11138,N_7362,N_5442);
or U11139 (N_11139,N_4973,N_5381);
or U11140 (N_11140,N_8949,N_2364);
and U11141 (N_11141,N_1048,N_8477);
or U11142 (N_11142,N_5096,N_6449);
and U11143 (N_11143,N_2565,N_1034);
or U11144 (N_11144,N_3877,N_430);
nor U11145 (N_11145,N_7568,N_7697);
and U11146 (N_11146,N_6917,N_574);
and U11147 (N_11147,N_6622,N_9715);
nor U11148 (N_11148,N_7187,N_3192);
and U11149 (N_11149,N_2407,N_3585);
nor U11150 (N_11150,N_9995,N_8972);
nor U11151 (N_11151,N_8740,N_857);
nand U11152 (N_11152,N_5672,N_3205);
nand U11153 (N_11153,N_2605,N_4867);
nor U11154 (N_11154,N_6224,N_1193);
nor U11155 (N_11155,N_9416,N_5026);
nor U11156 (N_11156,N_3866,N_772);
nand U11157 (N_11157,N_9470,N_9901);
or U11158 (N_11158,N_893,N_6323);
nor U11159 (N_11159,N_564,N_6738);
nor U11160 (N_11160,N_5987,N_9186);
nand U11161 (N_11161,N_239,N_950);
and U11162 (N_11162,N_2330,N_3816);
and U11163 (N_11163,N_4768,N_5508);
nor U11164 (N_11164,N_9587,N_5303);
and U11165 (N_11165,N_6866,N_2921);
or U11166 (N_11166,N_8429,N_1844);
nand U11167 (N_11167,N_6470,N_6463);
and U11168 (N_11168,N_9427,N_7794);
and U11169 (N_11169,N_634,N_4311);
nor U11170 (N_11170,N_167,N_4840);
nor U11171 (N_11171,N_6882,N_5989);
nand U11172 (N_11172,N_8272,N_5846);
and U11173 (N_11173,N_1857,N_3979);
nor U11174 (N_11174,N_4112,N_6847);
nand U11175 (N_11175,N_9316,N_3247);
or U11176 (N_11176,N_4517,N_6127);
nand U11177 (N_11177,N_7481,N_7339);
and U11178 (N_11178,N_3084,N_7606);
or U11179 (N_11179,N_6455,N_7006);
and U11180 (N_11180,N_7673,N_8167);
and U11181 (N_11181,N_6899,N_8924);
and U11182 (N_11182,N_6667,N_9816);
nor U11183 (N_11183,N_6609,N_6849);
nor U11184 (N_11184,N_2173,N_5837);
nand U11185 (N_11185,N_9062,N_416);
nor U11186 (N_11186,N_6230,N_3907);
or U11187 (N_11187,N_8187,N_3004);
or U11188 (N_11188,N_9262,N_3916);
and U11189 (N_11189,N_1290,N_6380);
xor U11190 (N_11190,N_9638,N_2641);
nor U11191 (N_11191,N_6159,N_8616);
nand U11192 (N_11192,N_5634,N_1107);
and U11193 (N_11193,N_1842,N_789);
nand U11194 (N_11194,N_3365,N_4217);
nor U11195 (N_11195,N_5199,N_5697);
or U11196 (N_11196,N_1830,N_2836);
nand U11197 (N_11197,N_9559,N_5696);
or U11198 (N_11198,N_3794,N_1145);
or U11199 (N_11199,N_4737,N_263);
nand U11200 (N_11200,N_5004,N_1514);
or U11201 (N_11201,N_162,N_5483);
nor U11202 (N_11202,N_4654,N_7430);
and U11203 (N_11203,N_879,N_7988);
and U11204 (N_11204,N_6105,N_4723);
and U11205 (N_11205,N_7860,N_7782);
and U11206 (N_11206,N_3303,N_7092);
and U11207 (N_11207,N_3532,N_6837);
nand U11208 (N_11208,N_2182,N_6383);
nand U11209 (N_11209,N_5478,N_1060);
nor U11210 (N_11210,N_6274,N_831);
and U11211 (N_11211,N_7078,N_1481);
nor U11212 (N_11212,N_5414,N_4470);
nand U11213 (N_11213,N_7539,N_4947);
nor U11214 (N_11214,N_8299,N_8662);
nor U11215 (N_11215,N_2686,N_1799);
nand U11216 (N_11216,N_3829,N_6064);
nor U11217 (N_11217,N_1497,N_8437);
nor U11218 (N_11218,N_1723,N_5834);
nand U11219 (N_11219,N_9157,N_1969);
or U11220 (N_11220,N_1652,N_7110);
or U11221 (N_11221,N_6205,N_1938);
or U11222 (N_11222,N_5621,N_3187);
and U11223 (N_11223,N_9490,N_4939);
or U11224 (N_11224,N_6568,N_4721);
nor U11225 (N_11225,N_778,N_9647);
and U11226 (N_11226,N_7808,N_1069);
nand U11227 (N_11227,N_2444,N_5851);
or U11228 (N_11228,N_1622,N_3208);
nand U11229 (N_11229,N_7852,N_3334);
or U11230 (N_11230,N_5818,N_4237);
nand U11231 (N_11231,N_6467,N_7908);
nor U11232 (N_11232,N_1413,N_1515);
nor U11233 (N_11233,N_7857,N_2131);
nand U11234 (N_11234,N_4055,N_9397);
xor U11235 (N_11235,N_5729,N_3767);
or U11236 (N_11236,N_6867,N_9693);
nor U11237 (N_11237,N_6335,N_2920);
nor U11238 (N_11238,N_4835,N_8260);
nor U11239 (N_11239,N_1956,N_1228);
nand U11240 (N_11240,N_9440,N_2931);
and U11241 (N_11241,N_4837,N_1445);
or U11242 (N_11242,N_1405,N_8315);
or U11243 (N_11243,N_742,N_1937);
or U11244 (N_11244,N_8819,N_7249);
nand U11245 (N_11245,N_2786,N_9481);
nand U11246 (N_11246,N_6087,N_4305);
or U11247 (N_11247,N_1720,N_2438);
or U11248 (N_11248,N_6081,N_8586);
or U11249 (N_11249,N_3106,N_2292);
nor U11250 (N_11250,N_3838,N_5393);
or U11251 (N_11251,N_1808,N_5219);
and U11252 (N_11252,N_9564,N_1096);
nor U11253 (N_11253,N_4505,N_2221);
and U11254 (N_11254,N_5796,N_8699);
nand U11255 (N_11255,N_8231,N_813);
nor U11256 (N_11256,N_5468,N_9330);
and U11257 (N_11257,N_8553,N_8770);
nand U11258 (N_11258,N_762,N_4660);
nor U11259 (N_11259,N_158,N_5375);
and U11260 (N_11260,N_4953,N_8163);
or U11261 (N_11261,N_1912,N_8573);
and U11262 (N_11262,N_7554,N_5456);
nor U11263 (N_11263,N_5930,N_4279);
nor U11264 (N_11264,N_137,N_6554);
nand U11265 (N_11265,N_4708,N_2919);
nor U11266 (N_11266,N_6909,N_1669);
nand U11267 (N_11267,N_9790,N_6972);
nand U11268 (N_11268,N_1386,N_6183);
nor U11269 (N_11269,N_2630,N_7303);
nand U11270 (N_11270,N_8105,N_652);
or U11271 (N_11271,N_5213,N_8806);
nand U11272 (N_11272,N_7557,N_7694);
and U11273 (N_11273,N_1249,N_6237);
and U11274 (N_11274,N_8067,N_9830);
nand U11275 (N_11275,N_1680,N_7884);
or U11276 (N_11276,N_955,N_5287);
nor U11277 (N_11277,N_9643,N_533);
xor U11278 (N_11278,N_9607,N_3810);
and U11279 (N_11279,N_2294,N_3430);
and U11280 (N_11280,N_9432,N_442);
and U11281 (N_11281,N_2051,N_178);
nor U11282 (N_11282,N_9593,N_4145);
nand U11283 (N_11283,N_6257,N_4730);
nor U11284 (N_11284,N_3254,N_3353);
or U11285 (N_11285,N_2991,N_5010);
nand U11286 (N_11286,N_1833,N_3238);
or U11287 (N_11287,N_7370,N_9166);
xor U11288 (N_11288,N_6379,N_194);
nor U11289 (N_11289,N_423,N_8042);
or U11290 (N_11290,N_6869,N_8932);
or U11291 (N_11291,N_8832,N_2948);
nand U11292 (N_11292,N_4111,N_7212);
nor U11293 (N_11293,N_1489,N_3827);
nor U11294 (N_11294,N_8600,N_4853);
nor U11295 (N_11295,N_3913,N_488);
and U11296 (N_11296,N_8964,N_4118);
or U11297 (N_11297,N_9746,N_4450);
or U11298 (N_11298,N_5411,N_4994);
nor U11299 (N_11299,N_5311,N_9632);
xor U11300 (N_11300,N_7264,N_8750);
or U11301 (N_11301,N_5707,N_6686);
nor U11302 (N_11302,N_3124,N_9596);
and U11303 (N_11303,N_4215,N_8876);
nand U11304 (N_11304,N_5557,N_6684);
and U11305 (N_11305,N_3686,N_8721);
or U11306 (N_11306,N_5118,N_8119);
and U11307 (N_11307,N_9370,N_6310);
nand U11308 (N_11308,N_8211,N_2762);
or U11309 (N_11309,N_9107,N_7062);
nor U11310 (N_11310,N_3928,N_4354);
nor U11311 (N_11311,N_971,N_4793);
nor U11312 (N_11312,N_3185,N_2717);
and U11313 (N_11313,N_7028,N_8390);
or U11314 (N_11314,N_4398,N_2196);
nand U11315 (N_11315,N_218,N_8653);
nand U11316 (N_11316,N_7143,N_595);
and U11317 (N_11317,N_7854,N_560);
or U11318 (N_11318,N_9122,N_9233);
or U11319 (N_11319,N_7079,N_1398);
and U11320 (N_11320,N_7703,N_4845);
or U11321 (N_11321,N_5476,N_341);
nand U11322 (N_11322,N_5183,N_4878);
xor U11323 (N_11323,N_3862,N_2573);
nand U11324 (N_11324,N_2380,N_2822);
nand U11325 (N_11325,N_1764,N_9684);
or U11326 (N_11326,N_9667,N_7804);
nand U11327 (N_11327,N_7361,N_25);
nand U11328 (N_11328,N_4913,N_1027);
nor U11329 (N_11329,N_7480,N_2009);
nor U11330 (N_11330,N_6862,N_4032);
xor U11331 (N_11331,N_7894,N_5572);
and U11332 (N_11332,N_7365,N_6236);
and U11333 (N_11333,N_8124,N_1632);
or U11334 (N_11334,N_9158,N_8320);
and U11335 (N_11335,N_8635,N_1438);
nand U11336 (N_11336,N_8224,N_709);
nand U11337 (N_11337,N_3088,N_5914);
and U11338 (N_11338,N_4565,N_9364);
or U11339 (N_11339,N_2112,N_180);
nand U11340 (N_11340,N_2933,N_259);
nor U11341 (N_11341,N_8487,N_1815);
nand U11342 (N_11342,N_845,N_413);
nand U11343 (N_11343,N_8842,N_5006);
xor U11344 (N_11344,N_3707,N_7968);
nor U11345 (N_11345,N_4326,N_9181);
and U11346 (N_11346,N_4719,N_7048);
nand U11347 (N_11347,N_407,N_2241);
and U11348 (N_11348,N_8472,N_3362);
and U11349 (N_11349,N_9827,N_1149);
nand U11350 (N_11350,N_2618,N_1041);
and U11351 (N_11351,N_747,N_4367);
or U11352 (N_11352,N_2936,N_7547);
nor U11353 (N_11353,N_202,N_7653);
or U11354 (N_11354,N_8952,N_5294);
and U11355 (N_11355,N_8478,N_8622);
and U11356 (N_11356,N_3173,N_1092);
or U11357 (N_11357,N_2391,N_7614);
and U11358 (N_11358,N_9922,N_8443);
nand U11359 (N_11359,N_2871,N_3950);
nor U11360 (N_11360,N_2457,N_1737);
and U11361 (N_11361,N_7377,N_7293);
and U11362 (N_11362,N_1402,N_4861);
or U11363 (N_11363,N_716,N_3466);
and U11364 (N_11364,N_8077,N_1602);
or U11365 (N_11365,N_1502,N_5777);
nor U11366 (N_11366,N_943,N_3442);
and U11367 (N_11367,N_5030,N_2365);
and U11368 (N_11368,N_5200,N_3648);
nand U11369 (N_11369,N_8890,N_255);
nand U11370 (N_11370,N_1600,N_7960);
and U11371 (N_11371,N_8156,N_7561);
and U11372 (N_11372,N_9468,N_3657);
or U11373 (N_11373,N_6809,N_4990);
and U11374 (N_11374,N_4393,N_8049);
and U11375 (N_11375,N_5848,N_6401);
nand U11376 (N_11376,N_3227,N_1486);
nor U11377 (N_11377,N_5321,N_4468);
nor U11378 (N_11378,N_6282,N_4930);
and U11379 (N_11379,N_5980,N_6969);
nor U11380 (N_11380,N_7755,N_5561);
nor U11381 (N_11381,N_1355,N_1083);
nand U11382 (N_11382,N_5541,N_8991);
or U11383 (N_11383,N_1399,N_1403);
nor U11384 (N_11384,N_6602,N_2093);
and U11385 (N_11385,N_45,N_4811);
or U11386 (N_11386,N_6301,N_4965);
nor U11387 (N_11387,N_8168,N_6767);
nand U11388 (N_11388,N_4363,N_5900);
and U11389 (N_11389,N_6287,N_1859);
nor U11390 (N_11390,N_4679,N_9465);
and U11391 (N_11391,N_6231,N_7889);
and U11392 (N_11392,N_443,N_9866);
nor U11393 (N_11393,N_5040,N_420);
or U11394 (N_11394,N_2789,N_5325);
nor U11395 (N_11395,N_9615,N_3401);
or U11396 (N_11396,N_1585,N_3497);
and U11397 (N_11397,N_5699,N_4018);
and U11398 (N_11398,N_4696,N_3445);
nor U11399 (N_11399,N_3891,N_6294);
nor U11400 (N_11400,N_911,N_3578);
nor U11401 (N_11401,N_7241,N_1976);
nand U11402 (N_11402,N_103,N_9270);
nand U11403 (N_11403,N_8139,N_5929);
nor U11404 (N_11404,N_9355,N_3986);
or U11405 (N_11405,N_7418,N_4138);
or U11406 (N_11406,N_6039,N_5108);
nor U11407 (N_11407,N_601,N_1574);
and U11408 (N_11408,N_7618,N_3070);
nor U11409 (N_11409,N_815,N_1948);
nor U11410 (N_11410,N_7460,N_5797);
or U11411 (N_11411,N_6735,N_4441);
and U11412 (N_11412,N_124,N_117);
nor U11413 (N_11413,N_4222,N_7388);
and U11414 (N_11414,N_8137,N_3426);
or U11415 (N_11415,N_862,N_1634);
nor U11416 (N_11416,N_1616,N_3748);
and U11417 (N_11417,N_6747,N_3424);
and U11418 (N_11418,N_8107,N_1885);
and U11419 (N_11419,N_3762,N_5095);
nor U11420 (N_11420,N_6789,N_9492);
and U11421 (N_11421,N_7813,N_8791);
nand U11422 (N_11422,N_8022,N_3414);
nand U11423 (N_11423,N_1381,N_8666);
nor U11424 (N_11424,N_1499,N_3791);
or U11425 (N_11425,N_7768,N_846);
nand U11426 (N_11426,N_698,N_509);
and U11427 (N_11427,N_493,N_4401);
or U11428 (N_11428,N_4126,N_3440);
nand U11429 (N_11429,N_615,N_7598);
or U11430 (N_11430,N_8263,N_8685);
or U11431 (N_11431,N_1401,N_9292);
or U11432 (N_11432,N_8081,N_306);
nand U11433 (N_11433,N_2346,N_7877);
and U11434 (N_11434,N_2682,N_7375);
nand U11435 (N_11435,N_2486,N_7391);
nor U11436 (N_11436,N_7724,N_602);
and U11437 (N_11437,N_9626,N_1281);
nand U11438 (N_11438,N_9147,N_6888);
nor U11439 (N_11439,N_8730,N_3122);
nor U11440 (N_11440,N_3250,N_3459);
and U11441 (N_11441,N_1285,N_3699);
and U11442 (N_11442,N_5379,N_6588);
nand U11443 (N_11443,N_8711,N_1444);
or U11444 (N_11444,N_1721,N_6177);
nand U11445 (N_11445,N_9450,N_4876);
nor U11446 (N_11446,N_7656,N_2497);
and U11447 (N_11447,N_2617,N_6361);
nor U11448 (N_11448,N_9951,N_4780);
or U11449 (N_11449,N_8241,N_5820);
or U11450 (N_11450,N_1572,N_1546);
or U11451 (N_11451,N_3774,N_765);
nand U11452 (N_11452,N_4303,N_4725);
or U11453 (N_11453,N_1475,N_2982);
nor U11454 (N_11454,N_9825,N_8759);
nand U11455 (N_11455,N_7710,N_576);
nand U11456 (N_11456,N_429,N_5612);
or U11457 (N_11457,N_3773,N_5049);
and U11458 (N_11458,N_2047,N_2575);
or U11459 (N_11459,N_1848,N_8978);
nand U11460 (N_11460,N_8814,N_9760);
nor U11461 (N_11461,N_4987,N_1360);
or U11462 (N_11462,N_7024,N_5080);
nand U11463 (N_11463,N_9720,N_8935);
nor U11464 (N_11464,N_3777,N_7733);
nand U11465 (N_11465,N_6626,N_6998);
nand U11466 (N_11466,N_9637,N_1665);
nor U11467 (N_11467,N_4437,N_5389);
and U11468 (N_11468,N_7512,N_1307);
or U11469 (N_11469,N_8489,N_5262);
nand U11470 (N_11470,N_7711,N_910);
and U11471 (N_11471,N_7644,N_9753);
and U11472 (N_11472,N_1854,N_7114);
and U11473 (N_11473,N_7973,N_3847);
or U11474 (N_11474,N_2024,N_6647);
nor U11475 (N_11475,N_8585,N_5316);
nand U11476 (N_11476,N_4069,N_2231);
nand U11477 (N_11477,N_367,N_8192);
or U11478 (N_11478,N_3333,N_3446);
and U11479 (N_11479,N_2606,N_4986);
nand U11480 (N_11480,N_2487,N_8747);
and U11481 (N_11481,N_580,N_6115);
nor U11482 (N_11482,N_9933,N_6843);
nor U11483 (N_11483,N_5318,N_6607);
nand U11484 (N_11484,N_7748,N_2910);
or U11485 (N_11485,N_8317,N_7100);
or U11486 (N_11486,N_3448,N_138);
and U11487 (N_11487,N_9445,N_7897);
or U11488 (N_11488,N_4142,N_8043);
or U11489 (N_11489,N_3654,N_4309);
nand U11490 (N_11490,N_4338,N_5382);
nor U11491 (N_11491,N_972,N_9879);
nor U11492 (N_11492,N_4799,N_1253);
nor U11493 (N_11493,N_3479,N_3803);
xnor U11494 (N_11494,N_2247,N_1869);
nand U11495 (N_11495,N_2973,N_2533);
nand U11496 (N_11496,N_1394,N_5481);
and U11497 (N_11497,N_4419,N_9349);
and U11498 (N_11498,N_7349,N_4905);
or U11499 (N_11499,N_7575,N_229);
nand U11500 (N_11500,N_9553,N_7674);
and U11501 (N_11501,N_2116,N_8961);
nor U11502 (N_11502,N_8146,N_6200);
or U11503 (N_11503,N_909,N_5011);
and U11504 (N_11504,N_8676,N_714);
nand U11505 (N_11505,N_1358,N_4334);
nor U11506 (N_11506,N_970,N_4710);
and U11507 (N_11507,N_9780,N_3349);
or U11508 (N_11508,N_6108,N_3073);
nor U11509 (N_11509,N_433,N_7111);
nand U11510 (N_11510,N_9859,N_5565);
or U11511 (N_11511,N_3788,N_7144);
nor U11512 (N_11512,N_896,N_3289);
nor U11513 (N_11513,N_633,N_9204);
or U11514 (N_11514,N_9817,N_2474);
nand U11515 (N_11515,N_3213,N_7613);
nand U11516 (N_11516,N_7831,N_4088);
nor U11517 (N_11517,N_4934,N_7904);
or U11518 (N_11518,N_9580,N_6255);
nor U11519 (N_11519,N_8632,N_9043);
or U11520 (N_11520,N_3195,N_3927);
and U11521 (N_11521,N_5472,N_1319);
or U11522 (N_11522,N_7839,N_8914);
or U11523 (N_11523,N_3190,N_2785);
or U11524 (N_11524,N_1503,N_8442);
nand U11525 (N_11525,N_177,N_649);
nand U11526 (N_11526,N_85,N_9820);
nor U11527 (N_11527,N_5249,N_9323);
nand U11528 (N_11528,N_5474,N_4298);
nor U11529 (N_11529,N_9377,N_7799);
and U11530 (N_11530,N_6756,N_383);
and U11531 (N_11531,N_664,N_9129);
nor U11532 (N_11532,N_5100,N_2917);
and U11533 (N_11533,N_4783,N_6465);
nand U11534 (N_11534,N_9504,N_3215);
and U11535 (N_11535,N_9318,N_1545);
nand U11536 (N_11536,N_8401,N_9074);
and U11537 (N_11537,N_888,N_8903);
nor U11538 (N_11538,N_7814,N_3026);
and U11539 (N_11539,N_6649,N_1047);
nand U11540 (N_11540,N_9476,N_2012);
or U11541 (N_11541,N_8003,N_8230);
nor U11542 (N_11542,N_3045,N_9220);
nand U11543 (N_11543,N_5447,N_8875);
nand U11544 (N_11544,N_6320,N_182);
and U11545 (N_11545,N_3152,N_8886);
or U11546 (N_11546,N_5922,N_3054);
nor U11547 (N_11547,N_254,N_2577);
nor U11548 (N_11548,N_1646,N_8533);
nand U11549 (N_11549,N_8922,N_1341);
and U11550 (N_11550,N_9891,N_4364);
and U11551 (N_11551,N_8870,N_6223);
or U11552 (N_11552,N_5662,N_6050);
or U11553 (N_11553,N_8096,N_2772);
nor U11554 (N_11554,N_2944,N_3631);
nor U11555 (N_11555,N_3111,N_2321);
or U11556 (N_11556,N_2045,N_6065);
and U11557 (N_11557,N_6387,N_3887);
nand U11558 (N_11558,N_7617,N_293);
or U11559 (N_11559,N_2279,N_3200);
and U11560 (N_11560,N_7389,N_1138);
and U11561 (N_11561,N_6526,N_1022);
nand U11562 (N_11562,N_2632,N_6374);
nor U11563 (N_11563,N_3999,N_5231);
and U11564 (N_11564,N_4029,N_8328);
or U11565 (N_11565,N_6572,N_4874);
or U11566 (N_11566,N_2896,N_8500);
and U11567 (N_11567,N_1480,N_9971);
nor U11568 (N_11568,N_5061,N_9098);
nand U11569 (N_11569,N_1254,N_510);
nor U11570 (N_11570,N_9526,N_1856);
nand U11571 (N_11571,N_8560,N_5937);
or U11572 (N_11572,N_2314,N_139);
or U11573 (N_11573,N_5789,N_4972);
nor U11574 (N_11574,N_4556,N_56);
nand U11575 (N_11575,N_8258,N_7290);
xor U11576 (N_11576,N_3957,N_1981);
nor U11577 (N_11577,N_9761,N_48);
or U11578 (N_11578,N_2025,N_5629);
or U11579 (N_11579,N_5602,N_6472);
nor U11580 (N_11580,N_4485,N_7491);
and U11581 (N_11581,N_7522,N_6623);
nand U11582 (N_11582,N_7251,N_3880);
nor U11583 (N_11583,N_6474,N_310);
or U11584 (N_11584,N_6032,N_6597);
nor U11585 (N_11585,N_8062,N_3850);
and U11586 (N_11586,N_9471,N_268);
nor U11587 (N_11587,N_4140,N_449);
and U11588 (N_11588,N_5056,N_3347);
nor U11589 (N_11589,N_1863,N_4124);
nand U11590 (N_11590,N_7616,N_9787);
nand U11591 (N_11591,N_7517,N_5974);
nand U11592 (N_11592,N_5428,N_7403);
nand U11593 (N_11593,N_6924,N_5686);
or U11594 (N_11594,N_966,N_5436);
nand U11595 (N_11595,N_6189,N_4622);
nor U11596 (N_11596,N_9571,N_1523);
nor U11597 (N_11597,N_5429,N_587);
nor U11598 (N_11598,N_6946,N_9258);
and U11599 (N_11599,N_801,N_6363);
and U11600 (N_11600,N_7344,N_2741);
nor U11601 (N_11601,N_7608,N_6566);
nor U11602 (N_11602,N_2855,N_3320);
or U11603 (N_11603,N_9563,N_7492);
nand U11604 (N_11604,N_1260,N_1589);
or U11605 (N_11605,N_3465,N_2642);
and U11606 (N_11606,N_1203,N_5355);
nand U11607 (N_11607,N_6247,N_8736);
nand U11608 (N_11608,N_4701,N_6246);
and U11609 (N_11609,N_4503,N_5188);
nor U11610 (N_11610,N_712,N_6840);
or U11611 (N_11611,N_370,N_8919);
or U11612 (N_11612,N_2482,N_646);
or U11613 (N_11613,N_9601,N_5658);
nor U11614 (N_11614,N_6276,N_1819);
nand U11615 (N_11615,N_1177,N_6299);
and U11616 (N_11616,N_4872,N_432);
nand U11617 (N_11617,N_1017,N_9341);
nor U11618 (N_11618,N_7937,N_8732);
nor U11619 (N_11619,N_9664,N_9200);
nand U11620 (N_11620,N_2402,N_1104);
nor U11621 (N_11621,N_8075,N_3800);
and U11622 (N_11622,N_2003,N_4532);
and U11623 (N_11623,N_2248,N_8681);
nand U11624 (N_11624,N_537,N_4078);
nor U11625 (N_11625,N_2280,N_644);
or U11626 (N_11626,N_8714,N_1583);
nor U11627 (N_11627,N_7165,N_409);
or U11628 (N_11628,N_702,N_6051);
nand U11629 (N_11629,N_3809,N_4663);
or U11630 (N_11630,N_6495,N_4668);
or U11631 (N_11631,N_5374,N_9624);
nand U11632 (N_11632,N_5129,N_5125);
and U11633 (N_11633,N_8943,N_715);
or U11634 (N_11634,N_8851,N_6213);
nor U11635 (N_11635,N_5025,N_8541);
and U11636 (N_11636,N_7098,N_7366);
and U11637 (N_11637,N_6784,N_230);
or U11638 (N_11638,N_927,N_8867);
nand U11639 (N_11639,N_706,N_7310);
or U11640 (N_11640,N_3101,N_4635);
and U11641 (N_11641,N_185,N_7058);
nand U11642 (N_11642,N_6150,N_5299);
and U11643 (N_11643,N_1649,N_1624);
nand U11644 (N_11644,N_3031,N_2549);
and U11645 (N_11645,N_6090,N_5207);
and U11646 (N_11646,N_3930,N_8338);
or U11647 (N_11647,N_2939,N_767);
nor U11648 (N_11648,N_9544,N_5270);
nor U11649 (N_11649,N_4662,N_1641);
and U11650 (N_11650,N_5872,N_3834);
nand U11651 (N_11651,N_8332,N_4490);
and U11652 (N_11652,N_9828,N_7651);
or U11653 (N_11653,N_4546,N_7610);
nand U11654 (N_11654,N_1370,N_8413);
nor U11655 (N_11655,N_384,N_4251);
nor U11656 (N_11656,N_1601,N_1416);
nand U11657 (N_11657,N_4202,N_4181);
nand U11658 (N_11658,N_7118,N_8860);
xnor U11659 (N_11659,N_1214,N_9913);
or U11660 (N_11660,N_6258,N_6806);
or U11661 (N_11661,N_1091,N_2460);
or U11662 (N_11662,N_8510,N_2080);
or U11663 (N_11663,N_4942,N_9491);
and U11664 (N_11664,N_3556,N_2763);
nor U11665 (N_11665,N_91,N_3633);
nor U11666 (N_11666,N_6045,N_5091);
and U11667 (N_11667,N_6770,N_9082);
nor U11668 (N_11668,N_9741,N_4750);
nor U11669 (N_11669,N_3496,N_2102);
nand U11670 (N_11670,N_9509,N_1586);
nand U11671 (N_11671,N_5350,N_1140);
and U11672 (N_11672,N_9120,N_3841);
nor U11673 (N_11673,N_6494,N_7409);
or U11674 (N_11674,N_2209,N_1233);
nand U11675 (N_11675,N_9136,N_7700);
or U11676 (N_11676,N_8072,N_918);
and U11677 (N_11677,N_739,N_3655);
xnor U11678 (N_11678,N_5388,N_7044);
or U11679 (N_11679,N_7393,N_4644);
nor U11680 (N_11680,N_8871,N_7282);
or U11681 (N_11681,N_225,N_6673);
or U11682 (N_11682,N_1757,N_73);
nor U11683 (N_11683,N_4717,N_9649);
nand U11684 (N_11684,N_3153,N_8353);
and U11685 (N_11685,N_2581,N_2534);
and U11686 (N_11686,N_1463,N_8418);
nor U11687 (N_11687,N_756,N_4156);
nor U11688 (N_11688,N_4821,N_2286);
nor U11689 (N_11689,N_1971,N_5590);
or U11690 (N_11690,N_3043,N_4313);
nand U11691 (N_11691,N_1922,N_5210);
and U11692 (N_11692,N_75,N_2725);
or U11693 (N_11693,N_5741,N_7527);
and U11694 (N_11694,N_2518,N_3220);
or U11695 (N_11695,N_8040,N_2929);
xor U11696 (N_11696,N_6121,N_8849);
nor U11697 (N_11697,N_6061,N_3618);
nand U11698 (N_11698,N_4522,N_2864);
and U11699 (N_11699,N_9785,N_6102);
or U11700 (N_11700,N_8053,N_8729);
or U11701 (N_11701,N_607,N_7708);
nand U11702 (N_11702,N_8917,N_1137);
nor U11703 (N_11703,N_7532,N_3540);
and U11704 (N_11704,N_6517,N_8291);
xor U11705 (N_11705,N_2307,N_7931);
or U11706 (N_11706,N_8652,N_4515);
and U11707 (N_11707,N_9254,N_1325);
and U11708 (N_11708,N_5454,N_4749);
nand U11709 (N_11709,N_5601,N_1120);
or U11710 (N_11710,N_3453,N_3557);
nand U11711 (N_11711,N_7661,N_5939);
or U11712 (N_11712,N_3002,N_9542);
or U11713 (N_11713,N_4603,N_6000);
or U11714 (N_11714,N_8287,N_74);
nor U11715 (N_11715,N_8898,N_1505);
nor U11716 (N_11716,N_3239,N_7198);
nor U11717 (N_11717,N_1849,N_8700);
nor U11718 (N_11718,N_275,N_3861);
nor U11719 (N_11719,N_8996,N_2805);
xnor U11720 (N_11720,N_559,N_6755);
nor U11721 (N_11721,N_2895,N_3846);
and U11722 (N_11722,N_7633,N_2582);
or U11723 (N_11723,N_8249,N_544);
and U11724 (N_11724,N_3396,N_4561);
xnor U11725 (N_11725,N_6538,N_5893);
nand U11726 (N_11726,N_9611,N_2278);
and U11727 (N_11727,N_9482,N_345);
or U11728 (N_11728,N_499,N_4671);
and U11729 (N_11729,N_5357,N_1057);
or U11730 (N_11730,N_3127,N_7847);
nor U11731 (N_11731,N_3910,N_1072);
nand U11732 (N_11732,N_237,N_9338);
nor U11733 (N_11733,N_4613,N_3288);
and U11734 (N_11734,N_9177,N_8191);
nand U11735 (N_11735,N_9455,N_9190);
and U11736 (N_11736,N_9029,N_311);
nor U11737 (N_11737,N_2863,N_947);
nor U11738 (N_11738,N_9956,N_1637);
and U11739 (N_11739,N_9493,N_5204);
nand U11740 (N_11740,N_2949,N_366);
and U11741 (N_11741,N_6783,N_9627);
nor U11742 (N_11742,N_8036,N_3253);
or U11743 (N_11743,N_334,N_4475);
nor U11744 (N_11744,N_8219,N_8509);
nand U11745 (N_11745,N_4672,N_7298);
or U11746 (N_11746,N_818,N_8154);
or U11747 (N_11747,N_7883,N_7002);
nand U11748 (N_11748,N_2399,N_7679);
nand U11749 (N_11749,N_4469,N_3180);
or U11750 (N_11750,N_9008,N_8131);
or U11751 (N_11751,N_8458,N_1565);
nor U11752 (N_11752,N_2153,N_4199);
and U11753 (N_11753,N_426,N_7042);
nand U11754 (N_11754,N_1164,N_6772);
nor U11755 (N_11755,N_2191,N_1796);
nor U11756 (N_11756,N_7594,N_276);
or U11757 (N_11757,N_8368,N_9331);
or U11758 (N_11758,N_7464,N_3397);
and U11759 (N_11759,N_6417,N_5524);
and U11760 (N_11760,N_4066,N_480);
nor U11761 (N_11761,N_8958,N_2101);
nand U11762 (N_11762,N_3175,N_1544);
or U11763 (N_11763,N_211,N_2660);
or U11764 (N_11764,N_986,N_5412);
nand U11765 (N_11765,N_6168,N_5648);
or U11766 (N_11766,N_1671,N_8973);
and U11767 (N_11767,N_1724,N_6366);
nor U11768 (N_11768,N_6553,N_3276);
nor U11769 (N_11769,N_2726,N_4411);
xnor U11770 (N_11770,N_5562,N_5814);
nand U11771 (N_11771,N_2104,N_4241);
nand U11772 (N_11772,N_8713,N_8382);
or U11773 (N_11773,N_4852,N_630);
and U11774 (N_11774,N_1153,N_2656);
nand U11775 (N_11775,N_5574,N_9791);
nor U11776 (N_11776,N_9118,N_620);
and U11777 (N_11777,N_1436,N_353);
nand U11778 (N_11778,N_9523,N_397);
and U11779 (N_11779,N_5084,N_38);
and U11780 (N_11780,N_6434,N_2226);
nand U11781 (N_11781,N_5801,N_692);
nand U11782 (N_11782,N_4618,N_3989);
and U11783 (N_11783,N_2349,N_5322);
and U11784 (N_11784,N_6629,N_487);
and U11785 (N_11785,N_5907,N_9917);
and U11786 (N_11786,N_9153,N_5014);
nor U11787 (N_11787,N_7394,N_610);
nand U11788 (N_11788,N_9456,N_4838);
nand U11789 (N_11789,N_4183,N_4144);
nand U11790 (N_11790,N_7986,N_2889);
nor U11791 (N_11791,N_3967,N_4530);
nor U11792 (N_11792,N_8969,N_9597);
nand U11793 (N_11793,N_1862,N_1779);
nor U11794 (N_11794,N_6076,N_4863);
and U11795 (N_11795,N_5751,N_72);
or U11796 (N_11796,N_2229,N_1638);
or U11797 (N_11797,N_7903,N_2004);
nand U11798 (N_11798,N_7851,N_5208);
and U11799 (N_11799,N_1894,N_5836);
nor U11800 (N_11800,N_2937,N_3390);
nor U11801 (N_11801,N_3456,N_8333);
xor U11802 (N_11802,N_9020,N_5333);
or U11803 (N_11803,N_594,N_1224);
nand U11804 (N_11804,N_3463,N_9507);
nor U11805 (N_11805,N_3063,N_9691);
nor U11806 (N_11806,N_3735,N_9997);
nand U11807 (N_11807,N_7345,N_1690);
or U11808 (N_11808,N_8395,N_2960);
and U11809 (N_11809,N_1415,N_6056);
nor U11810 (N_11810,N_4699,N_753);
nand U11811 (N_11811,N_1967,N_2752);
nor U11812 (N_11812,N_8858,N_9665);
nand U11813 (N_11813,N_5534,N_9909);
nand U11814 (N_11814,N_1904,N_8322);
nor U11815 (N_11815,N_6528,N_2852);
xor U11816 (N_11816,N_7734,N_5132);
nor U11817 (N_11817,N_3316,N_734);
or U11818 (N_11818,N_8285,N_2236);
nand U11819 (N_11819,N_1905,N_1400);
nor U11820 (N_11820,N_2693,N_624);
and U11821 (N_11821,N_8728,N_2587);
and U11822 (N_11822,N_3315,N_5343);
nand U11823 (N_11823,N_166,N_6763);
and U11824 (N_11824,N_1040,N_9092);
nor U11825 (N_11825,N_671,N_7842);
or U11826 (N_11826,N_5642,N_6563);
nor U11827 (N_11827,N_7015,N_360);
nand U11828 (N_11828,N_1996,N_4948);
or U11829 (N_11829,N_6072,N_7330);
nand U11830 (N_11830,N_3112,N_1161);
and U11831 (N_11831,N_6315,N_9474);
nand U11832 (N_11832,N_6678,N_4362);
and U11833 (N_11833,N_4605,N_4252);
or U11834 (N_11834,N_6868,N_5022);
or U11835 (N_11835,N_821,N_5587);
and U11836 (N_11836,N_8428,N_6209);
nor U11837 (N_11837,N_1802,N_4177);
nand U11838 (N_11838,N_6440,N_8051);
or U11839 (N_11839,N_1705,N_444);
or U11840 (N_11840,N_2519,N_9354);
nor U11841 (N_11841,N_3675,N_3806);
or U11842 (N_11842,N_5577,N_3680);
nand U11843 (N_11843,N_5936,N_7360);
nor U11844 (N_11844,N_309,N_5620);
nor U11845 (N_11845,N_3935,N_5910);
or U11846 (N_11846,N_6469,N_9769);
nand U11847 (N_11847,N_832,N_5081);
and U11848 (N_11848,N_2594,N_8708);
nand U11849 (N_11849,N_1508,N_637);
and U11850 (N_11850,N_5853,N_1143);
and U11851 (N_11851,N_722,N_5263);
nor U11852 (N_11852,N_6155,N_3492);
nand U11853 (N_11853,N_3118,N_7005);
nand U11854 (N_11854,N_3335,N_9150);
or U11855 (N_11855,N_2390,N_1411);
nor U11856 (N_11856,N_3507,N_9398);
nor U11857 (N_11857,N_2363,N_4554);
and U11858 (N_11858,N_6815,N_8421);
nor U11859 (N_11859,N_8449,N_7162);
or U11860 (N_11860,N_1139,N_1094);
nand U11861 (N_11861,N_203,N_9018);
and U11862 (N_11862,N_3751,N_5134);
nand U11863 (N_11863,N_948,N_7881);
or U11864 (N_11864,N_4356,N_8613);
and U11865 (N_11865,N_2903,N_4836);
and U11866 (N_11866,N_184,N_8887);
nor U11867 (N_11867,N_6212,N_4691);
and U11868 (N_11868,N_8006,N_2547);
nor U11869 (N_11869,N_3902,N_9963);
nand U11870 (N_11870,N_5175,N_1542);
nor U11871 (N_11871,N_8809,N_3183);
and U11872 (N_11872,N_8456,N_5606);
or U11873 (N_11873,N_1656,N_3632);
and U11874 (N_11874,N_5206,N_8403);
and U11875 (N_11875,N_8416,N_1191);
or U11876 (N_11876,N_2733,N_5237);
or U11877 (N_11877,N_1087,N_6325);
and U11878 (N_11878,N_54,N_7166);
and U11879 (N_11879,N_9002,N_7487);
nand U11880 (N_11880,N_3643,N_2000);
nor U11881 (N_11881,N_7354,N_3678);
or U11882 (N_11882,N_2445,N_6424);
and U11883 (N_11883,N_8069,N_5033);
nand U11884 (N_11884,N_4430,N_5948);
nand U11885 (N_11885,N_4283,N_5352);
or U11886 (N_11886,N_7224,N_4625);
and U11887 (N_11887,N_8076,N_581);
nand U11888 (N_11888,N_6824,N_5947);
and U11889 (N_11889,N_2485,N_8377);
or U11890 (N_11890,N_3505,N_5792);
nor U11891 (N_11891,N_7199,N_8020);
nor U11892 (N_11892,N_2803,N_2107);
nor U11893 (N_11893,N_3688,N_1113);
and U11894 (N_11894,N_7727,N_777);
nor U11895 (N_11895,N_525,N_7602);
or U11896 (N_11896,N_3457,N_553);
and U11897 (N_11897,N_737,N_8118);
and U11898 (N_11898,N_3681,N_6466);
nand U11899 (N_11899,N_7120,N_7816);
and U11900 (N_11900,N_5902,N_6399);
and U11901 (N_11901,N_3547,N_5275);
or U11902 (N_11902,N_3296,N_7929);
nand U11903 (N_11903,N_8995,N_5348);
or U11904 (N_11904,N_6458,N_6148);
nor U11905 (N_11905,N_1786,N_1681);
nand U11906 (N_11906,N_6225,N_9230);
or U11907 (N_11907,N_6901,N_3529);
and U11908 (N_11908,N_7333,N_976);
nor U11909 (N_11909,N_2537,N_9732);
nor U11910 (N_11910,N_8180,N_8639);
nand U11911 (N_11911,N_6286,N_7486);
and U11912 (N_11912,N_3336,N_3876);
nand U11913 (N_11913,N_5339,N_7245);
nand U11914 (N_11914,N_1573,N_2572);
nor U11915 (N_11915,N_2449,N_6787);
nand U11916 (N_11916,N_827,N_8580);
nor U11917 (N_11917,N_9994,N_7307);
and U11918 (N_11918,N_7095,N_8048);
and U11919 (N_11919,N_5110,N_7378);
nand U11920 (N_11920,N_335,N_497);
or U11921 (N_11921,N_4381,N_3518);
and U11922 (N_11922,N_5152,N_2902);
and U11923 (N_11923,N_6037,N_1543);
or U11924 (N_11924,N_3782,N_1562);
and U11925 (N_11925,N_4149,N_9373);
nand U11926 (N_11926,N_351,N_4772);
nand U11927 (N_11927,N_9501,N_9944);
or U11928 (N_11928,N_395,N_865);
xnor U11929 (N_11929,N_548,N_3988);
or U11930 (N_11930,N_1979,N_2501);
nand U11931 (N_11931,N_3541,N_6875);
or U11932 (N_11932,N_1363,N_5156);
and U11933 (N_11933,N_7369,N_8203);
nand U11934 (N_11934,N_7148,N_2592);
nor U11935 (N_11935,N_6682,N_708);
nand U11936 (N_11936,N_1762,N_8178);
and U11937 (N_11937,N_4771,N_9755);
and U11938 (N_11938,N_5089,N_1896);
nor U11939 (N_11939,N_9719,N_5860);
nor U11940 (N_11940,N_8089,N_4382);
or U11941 (N_11941,N_3589,N_2847);
or U11942 (N_11942,N_214,N_8626);
and U11943 (N_11943,N_9685,N_6555);
or U11944 (N_11944,N_6981,N_6618);
and U11945 (N_11945,N_9654,N_2146);
and U11946 (N_11946,N_7555,N_4917);
nor U11947 (N_11947,N_5337,N_3993);
or U11948 (N_11948,N_4247,N_4100);
nand U11949 (N_11949,N_9116,N_2493);
nand U11950 (N_11950,N_999,N_5688);
nor U11951 (N_11951,N_6641,N_9296);
and U11952 (N_11952,N_8884,N_1230);
or U11953 (N_11953,N_8593,N_5750);
and U11954 (N_11954,N_757,N_2523);
nand U11955 (N_11955,N_9786,N_4357);
and U11956 (N_11956,N_9216,N_3961);
nor U11957 (N_11957,N_3931,N_1201);
nand U11958 (N_11958,N_6733,N_7023);
nor U11959 (N_11959,N_3480,N_3851);
nand U11960 (N_11960,N_3009,N_604);
or U11961 (N_11961,N_4397,N_9224);
nor U11962 (N_11962,N_4773,N_8159);
nor U11963 (N_11963,N_2084,N_453);
and U11964 (N_11964,N_1855,N_4349);
or U11965 (N_11965,N_2255,N_1198);
nand U11966 (N_11966,N_2608,N_6573);
and U11967 (N_11967,N_5094,N_5928);
nor U11968 (N_11968,N_9604,N_7669);
or U11969 (N_11969,N_8496,N_2718);
and U11970 (N_11970,N_6442,N_4151);
and U11971 (N_11971,N_7823,N_1957);
or U11972 (N_11972,N_8073,N_3170);
nor U11973 (N_11973,N_9375,N_812);
or U11974 (N_11974,N_9508,N_3603);
and U11975 (N_11975,N_1722,N_5446);
nor U11976 (N_11976,N_993,N_5373);
nand U11977 (N_11977,N_3683,N_5260);
or U11978 (N_11978,N_8764,N_1308);
nor U11979 (N_11979,N_7459,N_8177);
or U11980 (N_11980,N_6988,N_7865);
nand U11981 (N_11981,N_806,N_6879);
nor U11982 (N_11982,N_1114,N_5399);
nand U11983 (N_11983,N_3202,N_4210);
or U11984 (N_11984,N_5384,N_3656);
and U11985 (N_11985,N_349,N_1875);
nand U11986 (N_11986,N_1647,N_7649);
and U11987 (N_11987,N_2117,N_5972);
or U11988 (N_11988,N_6646,N_7916);
nand U11989 (N_11989,N_7176,N_4590);
or U11990 (N_11990,N_887,N_2239);
or U11991 (N_11991,N_3962,N_3549);
nand U11992 (N_11992,N_3444,N_6461);
nand U11993 (N_11993,N_2354,N_7581);
and U11994 (N_11994,N_5112,N_1273);
and U11995 (N_11995,N_8186,N_7565);
nand U11996 (N_11996,N_300,N_9188);
and U11997 (N_11997,N_2222,N_7466);
nor U11998 (N_11998,N_4013,N_4900);
nand U11999 (N_11999,N_8344,N_1587);
nor U12000 (N_12000,N_6872,N_7571);
nor U12001 (N_12001,N_7713,N_4940);
or U12002 (N_12002,N_2957,N_4794);
nand U12003 (N_12003,N_8133,N_3099);
nor U12004 (N_12004,N_6519,N_7140);
or U12005 (N_12005,N_8905,N_5849);
or U12006 (N_12006,N_6398,N_2120);
or U12007 (N_12007,N_1526,N_3089);
nor U12008 (N_12008,N_6788,N_3766);
nand U12009 (N_12009,N_1021,N_6749);
and U12010 (N_12010,N_6103,N_5415);
or U12011 (N_12011,N_4615,N_3592);
and U12012 (N_12012,N_9046,N_7800);
nand U12013 (N_12013,N_4525,N_1010);
nor U12014 (N_12014,N_675,N_3514);
nand U12015 (N_12015,N_5963,N_5778);
nor U12016 (N_12016,N_1708,N_5453);
nor U12017 (N_12017,N_5068,N_9572);
and U12018 (N_12018,N_348,N_9560);
and U12019 (N_12019,N_3028,N_5614);
nor U12020 (N_12020,N_1685,N_2926);
nor U12021 (N_12021,N_590,N_3564);
or U12022 (N_12022,N_3901,N_1965);
nand U12023 (N_12023,N_9843,N_9282);
nand U12024 (N_12024,N_7472,N_7992);
and U12025 (N_12025,N_4086,N_3151);
nand U12026 (N_12026,N_9053,N_7483);
nand U12027 (N_12027,N_9872,N_5016);
or U12028 (N_12028,N_8901,N_2143);
or U12029 (N_12029,N_3555,N_9449);
nand U12030 (N_12030,N_8825,N_549);
nor U12031 (N_12031,N_3169,N_8490);
nor U12032 (N_12032,N_6292,N_8270);
and U12033 (N_12033,N_2947,N_68);
nor U12034 (N_12034,N_3085,N_6096);
nor U12035 (N_12035,N_4678,N_9764);
nor U12036 (N_12036,N_4669,N_9137);
and U12037 (N_12037,N_9325,N_8857);
or U12038 (N_12038,N_7049,N_2082);
nor U12039 (N_12039,N_5996,N_368);
nand U12040 (N_12040,N_3626,N_5082);
or U12041 (N_12041,N_3179,N_7170);
nand U12042 (N_12042,N_4680,N_1739);
and U12043 (N_12043,N_8878,N_1581);
nor U12044 (N_12044,N_4261,N_7549);
and U12045 (N_12045,N_55,N_5610);
nor U12046 (N_12046,N_3081,N_612);
and U12047 (N_12047,N_2483,N_3357);
nor U12048 (N_12048,N_9938,N_9424);
nand U12049 (N_12049,N_1295,N_4328);
or U12050 (N_12050,N_3427,N_8369);
nand U12051 (N_12051,N_3110,N_2301);
or U12052 (N_12052,N_1692,N_5160);
nand U12053 (N_12053,N_2629,N_5905);
nand U12054 (N_12054,N_5903,N_1567);
nor U12055 (N_12055,N_8583,N_6008);
or U12056 (N_12056,N_244,N_9280);
and U12057 (N_12057,N_7274,N_7675);
or U12058 (N_12058,N_8623,N_1716);
or U12059 (N_12059,N_4324,N_1064);
nor U12060 (N_12060,N_8227,N_9210);
and U12061 (N_12061,N_8892,N_9689);
nor U12062 (N_12062,N_6823,N_565);
or U12063 (N_12063,N_9641,N_7737);
nand U12064 (N_12064,N_9289,N_1102);
nor U12065 (N_12065,N_7283,N_7864);
xnor U12066 (N_12066,N_3652,N_9557);
or U12067 (N_12067,N_6266,N_3691);
nand U12068 (N_12068,N_1440,N_5607);
or U12069 (N_12069,N_9606,N_1977);
or U12070 (N_12070,N_450,N_6757);
nand U12071 (N_12071,N_6801,N_2065);
and U12072 (N_12072,N_7105,N_6699);
nand U12073 (N_12073,N_5057,N_7825);
or U12074 (N_12074,N_2031,N_1778);
or U12075 (N_12075,N_4414,N_2041);
and U12076 (N_12076,N_6024,N_6215);
or U12077 (N_12077,N_9383,N_2998);
or U12078 (N_12078,N_9514,N_7250);
nor U12079 (N_12079,N_7125,N_5305);
nor U12080 (N_12080,N_4508,N_9413);
and U12081 (N_12081,N_6696,N_3053);
xor U12082 (N_12082,N_8222,N_5171);
nand U12083 (N_12083,N_3836,N_4050);
nor U12084 (N_12084,N_7746,N_718);
or U12085 (N_12085,N_2118,N_7629);
and U12086 (N_12086,N_2958,N_4520);
and U12087 (N_12087,N_7501,N_3059);
nor U12088 (N_12088,N_5578,N_5153);
and U12089 (N_12089,N_3756,N_9985);
nor U12090 (N_12090,N_6376,N_8603);
or U12091 (N_12091,N_1240,N_6026);
or U12092 (N_12092,N_1124,N_2181);
nand U12093 (N_12093,N_2734,N_7444);
nand U12094 (N_12094,N_3807,N_3094);
nand U12095 (N_12095,N_8615,N_2328);
xor U12096 (N_12096,N_9284,N_6480);
xnor U12097 (N_12097,N_1623,N_9434);
nor U12098 (N_12098,N_198,N_5921);
nand U12099 (N_12099,N_5619,N_8038);
and U12100 (N_12100,N_9094,N_3553);
or U12101 (N_12101,N_6362,N_1393);
and U12102 (N_12102,N_1154,N_589);
and U12103 (N_12103,N_3128,N_3399);
or U12104 (N_12104,N_8277,N_4551);
or U12105 (N_12105,N_3012,N_7978);
and U12106 (N_12106,N_3189,N_8197);
nor U12107 (N_12107,N_741,N_8636);
nand U12108 (N_12108,N_1250,N_7959);
nand U12109 (N_12109,N_1108,N_4164);
nand U12110 (N_12110,N_4454,N_9702);
or U12111 (N_12111,N_2340,N_1667);
nand U12112 (N_12112,N_761,N_3344);
and U12113 (N_12113,N_1679,N_354);
nand U12114 (N_12114,N_9352,N_5146);
nand U12115 (N_12115,N_4196,N_2981);
or U12116 (N_12116,N_7612,N_3060);
and U12117 (N_12117,N_1013,N_7287);
nand U12118 (N_12118,N_1376,N_1466);
and U12119 (N_12119,N_3461,N_2178);
and U12120 (N_12120,N_4479,N_5609);
or U12121 (N_12121,N_8688,N_9072);
and U12122 (N_12122,N_768,N_766);
and U12123 (N_12123,N_838,N_5451);
and U12124 (N_12124,N_6854,N_1280);
nor U12125 (N_12125,N_7876,N_3708);
and U12126 (N_12126,N_9912,N_7347);
or U12127 (N_12127,N_4967,N_9335);
and U12128 (N_12128,N_1746,N_8771);
nand U12129 (N_12129,N_1357,N_4931);
nor U12130 (N_12130,N_3130,N_586);
nand U12131 (N_12131,N_8617,N_8444);
or U12132 (N_12132,N_9347,N_6084);
and U12133 (N_12133,N_8702,N_161);
nand U12134 (N_12134,N_2075,N_5312);
xor U12135 (N_12135,N_2578,N_3955);
nor U12136 (N_12136,N_3181,N_5899);
nand U12137 (N_12137,N_5550,N_3388);
or U12138 (N_12138,N_1740,N_4962);
and U12139 (N_12139,N_3695,N_4513);
and U12140 (N_12140,N_7928,N_688);
nor U12141 (N_12141,N_923,N_9844);
nand U12142 (N_12142,N_6188,N_6811);
and U12143 (N_12143,N_7453,N_2692);
xnor U12144 (N_12144,N_7186,N_4991);
nor U12145 (N_12145,N_8698,N_4834);
or U12146 (N_12146,N_7188,N_4988);
nand U12147 (N_12147,N_1464,N_5378);
or U12148 (N_12148,N_60,N_1185);
or U12149 (N_12149,N_9044,N_4665);
nand U12150 (N_12150,N_9443,N_2511);
nand U12151 (N_12151,N_6329,N_4152);
nand U12152 (N_12152,N_6898,N_8470);
nand U12153 (N_12153,N_284,N_6612);
and U12154 (N_12154,N_4961,N_1836);
or U12155 (N_12155,N_3799,N_4857);
nor U12156 (N_12156,N_6386,N_8229);
and U12157 (N_12157,N_119,N_8099);
and U12158 (N_12158,N_4285,N_472);
nor U12159 (N_12159,N_3941,N_7484);
and U12160 (N_12160,N_711,N_6956);
and U12161 (N_12161,N_3982,N_830);
and U12162 (N_12162,N_315,N_7271);
and U12163 (N_12163,N_428,N_8284);
nand U12164 (N_12164,N_4653,N_5489);
nor U12165 (N_12165,N_6603,N_9123);
nand U12166 (N_12166,N_4828,N_435);
nand U12167 (N_12167,N_8517,N_6429);
nor U12168 (N_12168,N_8150,N_4843);
nor U12169 (N_12169,N_8987,N_7738);
or U12170 (N_12170,N_6454,N_3511);
and U12171 (N_12171,N_3044,N_93);
nand U12172 (N_12172,N_2643,N_9644);
or U12173 (N_12173,N_0,N_2335);
and U12174 (N_12174,N_2553,N_5064);
nand U12175 (N_12175,N_5871,N_4985);
and U12176 (N_12176,N_3441,N_7201);
and U12177 (N_12177,N_2795,N_8440);
and U12178 (N_12178,N_7363,N_4833);
or U12179 (N_12179,N_7001,N_2738);
or U12180 (N_12180,N_9666,N_1745);
nor U12181 (N_12181,N_8543,N_8199);
nor U12182 (N_12182,N_9084,N_7678);
nand U12183 (N_12183,N_8028,N_46);
or U12184 (N_12184,N_2154,N_512);
and U12185 (N_12185,N_6180,N_9678);
and U12186 (N_12186,N_9510,N_4234);
or U12187 (N_12187,N_411,N_3898);
nor U12188 (N_12188,N_6669,N_3331);
or U12189 (N_12189,N_34,N_3226);
nor U12190 (N_12190,N_5981,N_1781);
or U12191 (N_12191,N_6038,N_2839);
nor U12192 (N_12192,N_3212,N_4606);
or U12193 (N_12193,N_2094,N_446);
nand U12194 (N_12194,N_902,N_5031);
or U12195 (N_12195,N_3533,N_4203);
nand U12196 (N_12196,N_9274,N_7387);
nand U12197 (N_12197,N_1607,N_9391);
nand U12198 (N_12198,N_3061,N_8012);
or U12199 (N_12199,N_2633,N_6402);
and U12200 (N_12200,N_2177,N_2317);
nor U12201 (N_12201,N_3899,N_6328);
nor U12202 (N_12202,N_6071,N_7917);
and U12203 (N_12203,N_3567,N_2064);
nor U12204 (N_12204,N_9010,N_2913);
or U12205 (N_12205,N_9924,N_4301);
or U12206 (N_12206,N_1334,N_500);
and U12207 (N_12207,N_9590,N_6307);
nor U12208 (N_12208,N_1534,N_4464);
and U12209 (N_12209,N_8746,N_3370);
nand U12210 (N_12210,N_9539,N_5072);
nand U12211 (N_12211,N_4185,N_2218);
and U12212 (N_12212,N_4700,N_4971);
nor U12213 (N_12213,N_8054,N_1483);
or U12214 (N_12214,N_6006,N_7476);
nand U12215 (N_12215,N_4567,N_5552);
and U12216 (N_12216,N_9267,N_7805);
nand U12217 (N_12217,N_5763,N_286);
nand U12218 (N_12218,N_1729,N_5267);
nor U12219 (N_12219,N_2348,N_325);
or U12220 (N_12220,N_3299,N_5584);
and U12221 (N_12221,N_9300,N_3282);
nand U12222 (N_12222,N_1299,N_1395);
or U12223 (N_12223,N_4951,N_4978);
and U12224 (N_12224,N_6147,N_9980);
nor U12225 (N_12225,N_1283,N_3576);
nor U12226 (N_12226,N_7957,N_8552);
nor U12227 (N_12227,N_1420,N_8091);
or U12228 (N_12228,N_3372,N_6939);
or U12229 (N_12229,N_4021,N_2313);
and U12230 (N_12230,N_282,N_3339);
nor U12231 (N_12231,N_5927,N_3135);
nand U12232 (N_12232,N_9357,N_7392);
nor U12233 (N_12233,N_6793,N_833);
and U12234 (N_12234,N_327,N_5694);
nand U12235 (N_12235,N_9890,N_6358);
and U12236 (N_12236,N_7055,N_8348);
nor U12237 (N_12237,N_4016,N_6713);
and U12238 (N_12238,N_1098,N_6570);
and U12239 (N_12239,N_3925,N_3984);
and U12240 (N_12240,N_2695,N_6799);
nand U12241 (N_12241,N_3462,N_3025);
xnor U12242 (N_12242,N_2008,N_5812);
or U12243 (N_12243,N_6955,N_9163);
and U12244 (N_12244,N_5290,N_5248);
nor U12245 (N_12245,N_8847,N_7764);
nand U12246 (N_12246,N_5588,N_5546);
nor U12247 (N_12247,N_7056,N_4421);
nor U12248 (N_12248,N_8854,N_3770);
nand U12249 (N_12249,N_6754,N_3796);
and U12250 (N_12250,N_7454,N_7146);
nor U12251 (N_12251,N_1603,N_3911);
and U12252 (N_12252,N_2911,N_7087);
or U12253 (N_12253,N_3730,N_1032);
nand U12254 (N_12254,N_3650,N_3452);
or U12255 (N_12255,N_543,N_8064);
or U12256 (N_12256,N_7440,N_7096);
or U12257 (N_12257,N_8033,N_9996);
and U12258 (N_12258,N_8594,N_7435);
or U12259 (N_12259,N_2007,N_3473);
or U12260 (N_12260,N_6114,N_1146);
nor U12261 (N_12261,N_5819,N_5130);
nand U12262 (N_12262,N_3739,N_840);
and U12263 (N_12263,N_9078,N_2227);
or U12264 (N_12264,N_1916,N_8657);
nand U12265 (N_12265,N_876,N_6593);
nor U12266 (N_12266,N_9494,N_6856);
nand U12267 (N_12267,N_3743,N_1579);
and U12268 (N_12268,N_7536,N_6226);
or U12269 (N_12269,N_5145,N_6920);
nor U12270 (N_12270,N_969,N_7157);
and U12271 (N_12271,N_7022,N_2691);
and U12272 (N_12272,N_143,N_6457);
or U12273 (N_12273,N_8447,N_7870);
nand U12274 (N_12274,N_1148,N_9805);
nor U12275 (N_12275,N_2424,N_2905);
and U12276 (N_12276,N_8722,N_2386);
or U12277 (N_12277,N_2469,N_3165);
nand U12278 (N_12278,N_2032,N_9056);
or U12279 (N_12279,N_4388,N_8643);
and U12280 (N_12280,N_2095,N_5637);
xnor U12281 (N_12281,N_4439,N_4158);
and U12282 (N_12282,N_6701,N_8630);
nand U12283 (N_12283,N_1755,N_3001);
nor U12284 (N_12284,N_2160,N_6409);
nand U12285 (N_12285,N_9363,N_1697);
nand U12286 (N_12286,N_934,N_8660);
nor U12287 (N_12287,N_7134,N_6662);
or U12288 (N_12288,N_5722,N_2538);
nand U12289 (N_12289,N_2971,N_5788);
and U12290 (N_12290,N_6966,N_4192);
nand U12291 (N_12291,N_6858,N_1686);
and U12292 (N_12292,N_3684,N_7993);
and U12293 (N_12293,N_6508,N_3019);
nand U12294 (N_12294,N_2141,N_9959);
nor U12295 (N_12295,N_2140,N_9117);
and U12296 (N_12296,N_227,N_1293);
nor U12297 (N_12297,N_256,N_3801);
nor U12298 (N_12298,N_577,N_3184);
nor U12299 (N_12299,N_2645,N_5863);
or U12300 (N_12300,N_2983,N_2601);
nand U12301 (N_12301,N_3833,N_3166);
and U12302 (N_12302,N_216,N_4447);
nor U12303 (N_12303,N_1984,N_8100);
and U12304 (N_12304,N_3817,N_6959);
and U12305 (N_12305,N_8292,N_456);
or U12306 (N_12306,N_541,N_7273);
and U12307 (N_12307,N_5854,N_8384);
nor U12308 (N_12308,N_6117,N_5090);
nor U12309 (N_12309,N_4996,N_5277);
or U12310 (N_12310,N_2109,N_8065);
nor U12311 (N_12311,N_7625,N_8165);
nand U12312 (N_12312,N_47,N_5371);
nor U12313 (N_12313,N_1479,N_2397);
or U12314 (N_12314,N_6058,N_6208);
nor U12315 (N_12315,N_7364,N_4278);
or U12316 (N_12316,N_3964,N_9814);
or U12317 (N_12317,N_1163,N_4267);
xnor U12318 (N_12318,N_265,N_4549);
or U12319 (N_12319,N_6781,N_4611);
or U12320 (N_12320,N_6883,N_4135);
nand U12321 (N_12321,N_2527,N_1086);
or U12322 (N_12322,N_1966,N_3599);
nand U12323 (N_12323,N_1127,N_221);
and U12324 (N_12324,N_9964,N_6304);
nand U12325 (N_12325,N_2414,N_5623);
or U12326 (N_12326,N_1650,N_3105);
and U12327 (N_12327,N_4165,N_2477);
nand U12328 (N_12328,N_744,N_5661);
and U12329 (N_12329,N_1476,N_7646);
or U12330 (N_12330,N_754,N_1074);
and U12331 (N_12331,N_7422,N_6651);
and U12332 (N_12332,N_9556,N_2515);
nor U12333 (N_12333,N_5236,N_277);
and U12334 (N_12334,N_6342,N_9170);
and U12335 (N_12335,N_3312,N_1330);
nand U12336 (N_12336,N_9796,N_2761);
nor U12337 (N_12337,N_7801,N_2384);
nand U12338 (N_12338,N_1522,N_8715);
nand U12339 (N_12339,N_5743,N_7205);
or U12340 (N_12340,N_8765,N_4330);
or U12341 (N_12341,N_9832,N_8195);
nand U12342 (N_12342,N_9888,N_2439);
or U12343 (N_12343,N_9835,N_9162);
nand U12344 (N_12344,N_6497,N_9436);
nor U12345 (N_12345,N_3022,N_2670);
or U12346 (N_12346,N_8965,N_5158);
and U12347 (N_12347,N_5641,N_4936);
nor U12348 (N_12348,N_6317,N_9115);
or U12349 (N_12349,N_9175,N_20);
or U12350 (N_12350,N_5437,N_4957);
and U12351 (N_12351,N_6846,N_5982);
nor U12352 (N_12352,N_5549,N_4609);
or U12353 (N_12353,N_3888,N_1029);
nor U12354 (N_12354,N_2800,N_4405);
nor U12355 (N_12355,N_1210,N_4035);
nand U12356 (N_12356,N_850,N_8484);
nor U12357 (N_12357,N_5276,N_2707);
or U12358 (N_12358,N_9857,N_5341);
nand U12359 (N_12359,N_1459,N_9340);
nand U12360 (N_12360,N_5755,N_1156);
nor U12361 (N_12361,N_1851,N_6009);
nor U12362 (N_12362,N_7909,N_8365);
nor U12363 (N_12363,N_2784,N_1998);
and U12364 (N_12364,N_6165,N_2967);
nand U12365 (N_12365,N_9639,N_1872);
nand U12366 (N_12366,N_540,N_8866);
nor U12367 (N_12367,N_6726,N_6639);
or U12368 (N_12368,N_9661,N_925);
nor U12369 (N_12369,N_4384,N_5770);
and U12370 (N_12370,N_7754,N_6013);
nand U12371 (N_12371,N_8684,N_6702);
and U12372 (N_12372,N_7849,N_4887);
and U12373 (N_12373,N_7605,N_3341);
or U12374 (N_12374,N_3030,N_6251);
and U12375 (N_12375,N_8584,N_2968);
nand U12376 (N_12376,N_1596,N_3468);
or U12377 (N_12377,N_9521,N_5223);
or U12378 (N_12378,N_9990,N_6269);
and U12379 (N_12379,N_7896,N_5000);
nand U12380 (N_12380,N_782,N_9841);
and U12381 (N_12381,N_8950,N_4776);
nor U12382 (N_12382,N_2918,N_6509);
nand U12383 (N_12383,N_1014,N_6277);
nand U12384 (N_12384,N_8183,N_3035);
nor U12385 (N_12385,N_4981,N_9620);
nand U12386 (N_12386,N_336,N_2953);
and U12387 (N_12387,N_9610,N_6822);
or U12388 (N_12388,N_7145,N_2198);
and U12389 (N_12389,N_4770,N_3275);
and U12390 (N_12390,N_4060,N_1962);
and U12391 (N_12391,N_6728,N_7269);
nor U12392 (N_12392,N_4871,N_3157);
or U12393 (N_12393,N_7677,N_1374);
and U12394 (N_12394,N_9675,N_454);
and U12395 (N_12395,N_9140,N_8739);
xor U12396 (N_12396,N_3038,N_2808);
nand U12397 (N_12397,N_7067,N_4920);
and U12398 (N_12398,N_8766,N_9681);
or U12399 (N_12399,N_1202,N_1216);
and U12400 (N_12400,N_2326,N_5495);
nand U12401 (N_12401,N_5484,N_1644);
nand U12402 (N_12402,N_1759,N_1465);
and U12403 (N_12403,N_7445,N_9174);
or U12404 (N_12404,N_1599,N_4817);
or U12405 (N_12405,N_7853,N_6048);
or U12406 (N_12406,N_7965,N_875);
and U12407 (N_12407,N_357,N_1615);
nor U12408 (N_12408,N_4909,N_9420);
and U12409 (N_12409,N_4555,N_7045);
nor U12410 (N_12410,N_6761,N_1454);
or U12411 (N_12411,N_6210,N_2213);
nor U12412 (N_12412,N_2835,N_302);
and U12413 (N_12413,N_7451,N_8821);
and U12414 (N_12414,N_3,N_5951);
nor U12415 (N_12415,N_9783,N_7474);
and U12416 (N_12416,N_7778,N_7425);
nor U12417 (N_12417,N_4274,N_1606);
nand U12418 (N_12418,N_6992,N_8173);
nand U12419 (N_12419,N_7507,N_9421);
and U12420 (N_12420,N_1262,N_9622);
and U12421 (N_12421,N_5822,N_5240);
or U12422 (N_12422,N_4167,N_3814);
or U12423 (N_12423,N_2586,N_6715);
nor U12424 (N_12424,N_8453,N_7530);
and U12425 (N_12425,N_1327,N_4449);
nand U12426 (N_12426,N_7867,N_6740);
and U12427 (N_12427,N_1655,N_5323);
nand U12428 (N_12428,N_5521,N_6932);
nand U12429 (N_12429,N_7359,N_3872);
nand U12430 (N_12430,N_7743,N_9141);
and U12431 (N_12431,N_6248,N_4027);
or U12432 (N_12432,N_6643,N_6610);
nor U12433 (N_12433,N_473,N_4059);
or U12434 (N_12434,N_451,N_4714);
or U12435 (N_12435,N_984,N_6752);
nor U12436 (N_12436,N_2584,N_5037);
and U12437 (N_12437,N_1897,N_7779);
and U12438 (N_12438,N_8820,N_5579);
and U12439 (N_12439,N_4125,N_3422);
and U12440 (N_12440,N_5631,N_5423);
and U12441 (N_12441,N_7803,N_8558);
nand U12442 (N_12442,N_4769,N_9851);
or U12443 (N_12443,N_4121,N_2151);
or U12444 (N_12444,N_2768,N_3306);
or U12445 (N_12445,N_981,N_4281);
nor U12446 (N_12446,N_8019,N_7531);
nor U12447 (N_12447,N_4869,N_7761);
and U12448 (N_12448,N_9568,N_3894);
and U12449 (N_12449,N_2134,N_907);
and U12450 (N_12450,N_99,N_7434);
or U12451 (N_12451,N_5358,N_2049);
nor U12452 (N_12452,N_7722,N_1924);
and U12453 (N_12453,N_7576,N_3304);
or U12454 (N_12454,N_6695,N_967);
or U12455 (N_12455,N_4097,N_1750);
and U12456 (N_12456,N_7076,N_8015);
or U12457 (N_12457,N_7915,N_5733);
and U12458 (N_12458,N_4046,N_3860);
nand U12459 (N_12459,N_77,N_4534);
and U12460 (N_12460,N_2906,N_7467);
or U12461 (N_12461,N_9045,N_200);
and U12462 (N_12462,N_6748,N_4153);
or U12463 (N_12463,N_7025,N_3374);
nand U12464 (N_12464,N_4456,N_6086);
or U12465 (N_12465,N_6552,N_3845);
or U12466 (N_12466,N_4502,N_4657);
nor U12467 (N_12467,N_8680,N_5961);
or U12468 (N_12468,N_3725,N_418);
nand U12469 (N_12469,N_866,N_1339);
nand U12470 (N_12470,N_1504,N_8471);
nand U12471 (N_12471,N_4593,N_3293);
and U12472 (N_12472,N_6927,N_6614);
or U12473 (N_12473,N_5990,N_6887);
nor U12474 (N_12474,N_5876,N_3194);
xor U12475 (N_12475,N_3309,N_8136);
nor U12476 (N_12476,N_7334,N_5782);
and U12477 (N_12477,N_7313,N_5868);
or U12478 (N_12478,N_5998,N_3436);
nand U12479 (N_12479,N_1321,N_4372);
or U12480 (N_12480,N_1553,N_7967);
nor U12481 (N_12481,N_5956,N_1482);
and U12482 (N_12482,N_482,N_3755);
or U12483 (N_12483,N_5019,N_506);
and U12484 (N_12484,N_2589,N_5490);
or U12485 (N_12485,N_3513,N_1683);
or U12486 (N_12486,N_8143,N_222);
nor U12487 (N_12487,N_979,N_8436);
nand U12488 (N_12488,N_4929,N_848);
nand U12489 (N_12489,N_9981,N_1344);
or U12490 (N_12490,N_260,N_8412);
or U12491 (N_12491,N_7989,N_4702);
or U12492 (N_12492,N_6976,N_4751);
and U12493 (N_12493,N_6481,N_8841);
and U12494 (N_12494,N_4601,N_3016);
and U12495 (N_12495,N_2042,N_359);
nand U12496 (N_12496,N_5589,N_4583);
nand U12497 (N_12497,N_6561,N_1985);
nor U12498 (N_12498,N_619,N_5896);
nand U12499 (N_12499,N_9067,N_9298);
and U12500 (N_12500,N_2166,N_6711);
or U12501 (N_12501,N_1426,N_2769);
and U12502 (N_12502,N_1215,N_7939);
and U12503 (N_12503,N_2819,N_6596);
and U12504 (N_12504,N_1493,N_204);
nand U12505 (N_12505,N_8101,N_4722);
nand U12506 (N_12506,N_7753,N_7211);
nand U12507 (N_12507,N_2703,N_5356);
and U12508 (N_12508,N_1462,N_9109);
nand U12509 (N_12509,N_839,N_5909);
or U12510 (N_12510,N_7980,N_2345);
and U12511 (N_12511,N_4308,N_8446);
or U12512 (N_12512,N_3568,N_7910);
nand U12513 (N_12513,N_8423,N_8041);
nand U12514 (N_12514,N_2621,N_4147);
and U12515 (N_12515,N_2875,N_3998);
nand U12516 (N_12516,N_4188,N_1287);
nor U12517 (N_12517,N_2400,N_1653);
nand U12518 (N_12518,N_2615,N_296);
nand U12519 (N_12519,N_1540,N_8434);
or U12520 (N_12520,N_4968,N_2600);
and U12521 (N_12521,N_109,N_251);
or U12522 (N_12522,N_9970,N_5038);
nor U12523 (N_12523,N_9127,N_874);
nor U12524 (N_12524,N_1044,N_3909);
or U12525 (N_12525,N_3052,N_84);
or U12526 (N_12526,N_817,N_6498);
and U12527 (N_12527,N_4886,N_841);
or U12528 (N_12528,N_9293,N_6166);
nand U12529 (N_12529,N_1879,N_5480);
nand U12530 (N_12530,N_897,N_1425);
nor U12531 (N_12531,N_8840,N_3610);
nor U12532 (N_12532,N_1430,N_1888);
nor U12533 (N_12533,N_8419,N_4106);
nor U12534 (N_12534,N_4473,N_829);
and U12535 (N_12535,N_2535,N_3613);
or U12536 (N_12536,N_6355,N_6326);
and U12537 (N_12537,N_13,N_9257);
or U12538 (N_12538,N_2924,N_5823);
and U12539 (N_12539,N_6535,N_7521);
nand U12540 (N_12540,N_3662,N_31);
and U12541 (N_12541,N_9695,N_6074);
xnor U12542 (N_12542,N_524,N_2558);
and U12543 (N_12543,N_6918,N_6589);
or U12544 (N_12544,N_2892,N_6870);
or U12545 (N_12545,N_4073,N_9976);
nor U12546 (N_12546,N_4465,N_3915);
or U12547 (N_12547,N_4629,N_3501);
nor U12548 (N_12548,N_5563,N_9868);
or U12549 (N_12549,N_89,N_195);
and U12550 (N_12550,N_7026,N_7630);
nor U12551 (N_12551,N_2461,N_8432);
or U12552 (N_12552,N_7976,N_4591);
and U12553 (N_12553,N_936,N_7757);
or U12554 (N_12554,N_6745,N_154);
and U12555 (N_12555,N_5604,N_7463);
nand U12556 (N_12556,N_2466,N_611);
nor U12557 (N_12557,N_9788,N_8479);
nor U12558 (N_12558,N_7770,N_7417);
and U12559 (N_12559,N_3090,N_1237);
or U12560 (N_12560,N_4529,N_1510);
and U12561 (N_12561,N_1470,N_743);
or U12562 (N_12562,N_8112,N_4395);
or U12563 (N_12563,N_1352,N_2108);
and U12564 (N_12564,N_8963,N_7115);
nor U12565 (N_12565,N_7010,N_877);
or U12566 (N_12566,N_6818,N_810);
or U12567 (N_12567,N_7216,N_2499);
nor U12568 (N_12568,N_5076,N_6830);
nor U12569 (N_12569,N_1942,N_864);
or U12570 (N_12570,N_6178,N_5523);
nand U12571 (N_12571,N_2245,N_1882);
or U12572 (N_12572,N_9756,N_8844);
nand U12573 (N_12573,N_3522,N_1243);
xor U12574 (N_12574,N_1944,N_3855);
or U12575 (N_12575,N_583,N_8116);
nor U12576 (N_12576,N_1390,N_2275);
nand U12577 (N_12577,N_7835,N_9229);
or U12578 (N_12578,N_8321,N_7907);
nor U12579 (N_12579,N_1521,N_2454);
nand U12580 (N_12580,N_8677,N_828);
and U12581 (N_12581,N_8337,N_3647);
nand U12582 (N_12582,N_7252,N_1167);
and U12583 (N_12583,N_4417,N_683);
nor U12584 (N_12584,N_3469,N_183);
nand U12585 (N_12585,N_8980,N_2666);
nor U12586 (N_12586,N_3098,N_2459);
nor U12587 (N_12587,N_2420,N_188);
or U12588 (N_12588,N_2139,N_7619);
nand U12589 (N_12589,N_3234,N_1412);
and U12590 (N_12590,N_8610,N_4977);
or U12591 (N_12591,N_6321,N_582);
nor U12592 (N_12592,N_7542,N_8093);
nor U12593 (N_12593,N_5970,N_8529);
nor U12594 (N_12594,N_4209,N_9108);
nand U12595 (N_12595,N_1814,N_5718);
nand U12596 (N_12596,N_8706,N_2860);
nor U12597 (N_12597,N_3487,N_8226);
or U12598 (N_12598,N_6036,N_5477);
nor U12599 (N_12599,N_4726,N_6800);
and U12600 (N_12600,N_6970,N_7887);
and U12601 (N_12601,N_929,N_5832);
xnor U12602 (N_12602,N_1168,N_1209);
nand U12603 (N_12603,N_8304,N_3661);
nor U12604 (N_12604,N_1809,N_1300);
nand U12605 (N_12605,N_5332,N_1186);
or U12606 (N_12606,N_7747,N_3458);
and U12607 (N_12607,N_1820,N_371);
or U12608 (N_12608,N_9670,N_5291);
nor U12609 (N_12609,N_4883,N_1918);
and U12610 (N_12610,N_5736,N_6621);
or U12611 (N_12611,N_1991,N_6403);
and U12612 (N_12612,N_6558,N_6367);
nor U12613 (N_12613,N_5657,N_3223);
or U12614 (N_12614,N_588,N_2687);
nor U12615 (N_12615,N_6144,N_6974);
nor U12616 (N_12616,N_7340,N_5360);
or U12617 (N_12617,N_9353,N_1840);
nand U12618 (N_12618,N_7593,N_6303);
or U12619 (N_12619,N_363,N_8992);
nand U12620 (N_12620,N_7664,N_3015);
nor U12621 (N_12621,N_5857,N_9900);
nor U12622 (N_12622,N_2022,N_5509);
or U12623 (N_12623,N_6011,N_5002);
nor U12624 (N_12624,N_5531,N_4619);
and U12625 (N_12625,N_6331,N_4079);
nand U12626 (N_12626,N_1248,N_6343);
nor U12627 (N_12627,N_8761,N_5815);
nor U12628 (N_12628,N_1935,N_1892);
or U12629 (N_12629,N_2204,N_2985);
nor U12630 (N_12630,N_3665,N_4757);
nand U12631 (N_12631,N_9569,N_5813);
nand U12632 (N_12632,N_9561,N_4829);
nand U12633 (N_12633,N_7132,N_9864);
nor U12634 (N_12634,N_6389,N_9266);
and U12635 (N_12635,N_1577,N_8359);
and U12636 (N_12636,N_3351,N_1082);
nor U12637 (N_12637,N_7401,N_7276);
nand U12638 (N_12638,N_2130,N_2701);
nor U12639 (N_12639,N_3995,N_1838);
nand U12640 (N_12640,N_2925,N_9503);
nand U12641 (N_12641,N_7921,N_262);
nand U12642 (N_12642,N_6312,N_3011);
and U12643 (N_12643,N_9784,N_3472);
and U12644 (N_12644,N_2416,N_3071);
or U12645 (N_12645,N_1409,N_7922);
and U12646 (N_12646,N_1627,N_1725);
nor U12647 (N_12647,N_5581,N_5372);
or U12648 (N_12648,N_9394,N_5461);
and U12649 (N_12649,N_6599,N_7243);
xnor U12650 (N_12650,N_539,N_6385);
nand U12651 (N_12651,N_4455,N_6341);
or U12652 (N_12652,N_8046,N_9658);
nor U12653 (N_12653,N_659,N_1810);
nand U12654 (N_12654,N_751,N_6360);
nand U12655 (N_12655,N_1070,N_1380);
and U12656 (N_12656,N_6586,N_5391);
nor U12657 (N_12657,N_6940,N_5803);
nor U12658 (N_12658,N_3136,N_4022);
or U12659 (N_12659,N_5633,N_3554);
and U12660 (N_12660,N_4756,N_5113);
xnor U12661 (N_12661,N_1994,N_4);
or U12662 (N_12662,N_3843,N_7580);
xnor U12663 (N_12663,N_1682,N_2513);
or U12664 (N_12664,N_8058,N_2388);
or U12665 (N_12665,N_890,N_9402);
or U12666 (N_12666,N_1736,N_4652);
and U12667 (N_12667,N_3107,N_3790);
and U12668 (N_12668,N_5510,N_3754);
nand U12669 (N_12669,N_1404,N_2699);
or U12670 (N_12670,N_1811,N_279);
nor U12671 (N_12671,N_9208,N_6187);
or U12672 (N_12672,N_7149,N_1329);
or U12673 (N_12673,N_1418,N_8094);
nor U12674 (N_12674,N_5507,N_4875);
nor U12675 (N_12675,N_2425,N_2091);
nand U12676 (N_12676,N_2727,N_2465);
and U12677 (N_12677,N_4500,N_7197);
or U12678 (N_12678,N_5545,N_8846);
nor U12679 (N_12679,N_9842,N_2133);
nor U12680 (N_12680,N_3912,N_8893);
nor U12681 (N_12681,N_3132,N_4380);
or U12682 (N_12682,N_7981,N_1058);
and U12683 (N_12683,N_8405,N_9036);
or U12684 (N_12684,N_3732,N_6452);
nand U12685 (N_12685,N_2071,N_6207);
or U12686 (N_12686,N_2790,N_632);
and U12687 (N_12687,N_803,N_9448);
nor U12688 (N_12688,N_3718,N_9039);
or U12689 (N_12689,N_2168,N_6990);
or U12690 (N_12690,N_7573,N_6053);
nand U12691 (N_12691,N_313,N_9618);
nand U12692 (N_12692,N_5435,N_9836);
and U12693 (N_12693,N_5222,N_2882);
and U12694 (N_12694,N_2106,N_6906);
and U12695 (N_12695,N_8863,N_1495);
nand U12696 (N_12696,N_8788,N_8710);
nor U12697 (N_12697,N_5703,N_3167);
or U12698 (N_12698,N_5015,N_4243);
and U12699 (N_12699,N_8928,N_4001);
and U12700 (N_12700,N_1172,N_609);
nor U12701 (N_12701,N_6451,N_1753);
xnor U12702 (N_12702,N_2333,N_382);
and U12703 (N_12703,N_6576,N_1776);
nor U12704 (N_12704,N_2506,N_6145);
nand U12705 (N_12705,N_8544,N_1067);
and U12706 (N_12706,N_9911,N_8955);
or U12707 (N_12707,N_5943,N_5433);
nor U12708 (N_12708,N_1886,N_3258);
nor U12709 (N_12709,N_3673,N_1763);
or U12710 (N_12710,N_1554,N_7990);
or U12711 (N_12711,N_8748,N_980);
and U12712 (N_12712,N_596,N_6852);
nor U12713 (N_12713,N_3973,N_7404);
nor U12714 (N_12714,N_6406,N_4540);
nand U12715 (N_12715,N_4862,N_8130);
or U12716 (N_12716,N_8563,N_651);
and U12717 (N_12717,N_5571,N_9782);
and U12718 (N_12718,N_5288,N_8391);
nand U12719 (N_12719,N_8818,N_6423);
nand U12720 (N_12720,N_5944,N_4137);
and U12721 (N_12721,N_130,N_1707);
nor U12722 (N_12722,N_2121,N_1770);
nand U12723 (N_12723,N_5109,N_8908);
nor U12724 (N_12724,N_4296,N_2815);
and U12725 (N_12725,N_7351,N_6548);
or U12726 (N_12726,N_5839,N_770);
and U12727 (N_12727,N_8188,N_5455);
or U12728 (N_12728,N_6925,N_2524);
nor U12729 (N_12729,N_6577,N_7520);
and U12730 (N_12730,N_1353,N_3805);
nand U12731 (N_12731,N_3612,N_6079);
nand U12732 (N_12732,N_5511,N_3163);
and U12733 (N_12733,N_6066,N_8282);
nor U12734 (N_12734,N_8792,N_5499);
nor U12735 (N_12735,N_8415,N_4620);
and U12736 (N_12736,N_1213,N_7514);
nor U12737 (N_12737,N_2428,N_2721);
or U12738 (N_12738,N_4407,N_4753);
nand U12739 (N_12739,N_4810,N_6929);
and U12740 (N_12740,N_5702,N_1118);
nor U12741 (N_12741,N_1158,N_7054);
and U12742 (N_12742,N_7963,N_1033);
or U12743 (N_12743,N_5683,N_1282);
or U12744 (N_12744,N_3137,N_9288);
or U12745 (N_12745,N_6842,N_9498);
or U12746 (N_12746,N_3772,N_6488);
nor U12747 (N_12747,N_2522,N_7982);
nand U12748 (N_12748,N_7094,N_1356);
or U12749 (N_12749,N_1031,N_5843);
nor U12750 (N_12750,N_6437,N_7272);
nand U12751 (N_12751,N_4812,N_921);
nand U12752 (N_12752,N_1943,N_6313);
nand U12753 (N_12753,N_8812,N_6136);
and U12754 (N_12754,N_8784,N_3321);
or U12755 (N_12755,N_436,N_5024);
nor U12756 (N_12756,N_1275,N_1578);
nand U12757 (N_12757,N_5190,N_2811);
nand U12758 (N_12758,N_7972,N_3393);
nor U12759 (N_12759,N_2563,N_228);
or U12760 (N_12760,N_5630,N_9739);
and U12761 (N_12761,N_7322,N_7018);
nor U12762 (N_12762,N_5706,N_8060);
nor U12763 (N_12763,N_2709,N_6973);
or U12764 (N_12764,N_536,N_5594);
and U12765 (N_12765,N_4870,N_8454);
nand U12766 (N_12766,N_6938,N_4127);
and U12767 (N_12767,N_8102,N_6797);
and U12768 (N_12768,N_1972,N_5058);
and U12769 (N_12769,N_9452,N_4412);
nand U12770 (N_12770,N_2370,N_2516);
nor U12771 (N_12771,N_2480,N_9735);
or U12772 (N_12772,N_5576,N_2435);
and U12773 (N_12773,N_7374,N_5608);
nor U12774 (N_12774,N_1002,N_8461);
nand U12775 (N_12775,N_278,N_2479);
nand U12776 (N_12776,N_5800,N_8217);
and U12777 (N_12777,N_4157,N_9663);
and U12778 (N_12778,N_4763,N_2759);
nor U12779 (N_12779,N_5028,N_1788);
nor U12780 (N_12780,N_5779,N_6054);
and U12781 (N_12781,N_930,N_3936);
or U12782 (N_12782,N_9801,N_3939);
and U12783 (N_12783,N_320,N_1);
and U12784 (N_12784,N_8811,N_9529);
or U12785 (N_12785,N_1772,N_9892);
nor U12786 (N_12786,N_6010,N_490);
and U12787 (N_12787,N_7329,N_5835);
and U12788 (N_12788,N_9721,N_372);
or U12789 (N_12789,N_7031,N_5784);
nor U12790 (N_12790,N_3658,N_9533);
nand U12791 (N_12791,N_4284,N_4195);
nand U12792 (N_12792,N_2562,N_1053);
and U12793 (N_12793,N_5475,N_8248);
nand U12794 (N_12794,N_9530,N_6314);
and U12795 (N_12795,N_3158,N_5528);
or U12796 (N_12796,N_2315,N_7408);
or U12797 (N_12797,N_243,N_4512);
nor U12798 (N_12798,N_997,N_6948);
nand U12799 (N_12799,N_2688,N_4795);
nor U12800 (N_12800,N_528,N_8406);
nand U12801 (N_12801,N_4130,N_3297);
or U12802 (N_12802,N_7626,N_4204);
or U12803 (N_12803,N_3736,N_2539);
nor U12804 (N_12804,N_5320,N_3121);
or U12805 (N_12805,N_1831,N_6958);
nor U12806 (N_12806,N_78,N_704);
and U12807 (N_12807,N_3494,N_5850);
nand U12808 (N_12808,N_4778,N_29);
and U12809 (N_12809,N_6130,N_2780);
and U12810 (N_12810,N_6688,N_8252);
and U12811 (N_12811,N_5139,N_3758);
and U12812 (N_12812,N_3653,N_6698);
or U12813 (N_12813,N_9600,N_9860);
or U12814 (N_12814,N_2077,N_9898);
and U12815 (N_12815,N_5842,N_3360);
nand U12816 (N_12816,N_9060,N_2067);
or U12817 (N_12817,N_9942,N_5901);
nand U12818 (N_12818,N_7636,N_5670);
and U12819 (N_12819,N_6302,N_1558);
nor U12820 (N_12820,N_5238,N_7235);
or U12821 (N_12821,N_4056,N_679);
nand U12822 (N_12822,N_8373,N_8957);
or U12823 (N_12823,N_3214,N_5754);
nand U12824 (N_12824,N_6430,N_247);
or U12825 (N_12825,N_8082,N_5724);
nand U12826 (N_12826,N_2081,N_5362);
nand U12827 (N_12827,N_6289,N_1710);
or U12828 (N_12828,N_9113,N_9937);
or U12829 (N_12829,N_9311,N_1396);
and U12830 (N_12830,N_5440,N_9017);
or U12831 (N_12831,N_6505,N_9035);
nor U12832 (N_12832,N_9821,N_5289);
or U12833 (N_12833,N_9447,N_759);
or U12834 (N_12834,N_9329,N_7962);
nor U12835 (N_12835,N_797,N_3325);
and U12836 (N_12836,N_6780,N_8640);
and U12837 (N_12837,N_5527,N_5310);
and U12838 (N_12838,N_6880,N_6445);
nand U12839 (N_12839,N_6665,N_7465);
nand U12840 (N_12840,N_1953,N_6093);
and U12841 (N_12841,N_3546,N_9295);
nand U12842 (N_12842,N_8648,N_7899);
or U12843 (N_12843,N_5390,N_7352);
nor U12844 (N_12844,N_5445,N_9478);
or U12845 (N_12845,N_4221,N_9431);
nand U12846 (N_12846,N_3498,N_6104);
and U12847 (N_12847,N_8417,N_8551);
nor U12848 (N_12848,N_1608,N_6206);
or U12849 (N_12849,N_2214,N_8056);
nand U12850 (N_12850,N_3483,N_8309);
nand U12851 (N_12851,N_5035,N_3037);
nor U12852 (N_12852,N_3619,N_1993);
or U12853 (N_12853,N_8181,N_643);
or U12854 (N_12854,N_6203,N_8528);
nand U12855 (N_12855,N_8160,N_1812);
nand U12856 (N_12856,N_1580,N_5769);
nor U12857 (N_12857,N_935,N_4282);
or U12858 (N_12858,N_9406,N_2930);
or U12859 (N_12859,N_6468,N_6435);
or U12860 (N_12860,N_685,N_2086);
nand U12861 (N_12861,N_7597,N_8210);
and U12862 (N_12862,N_2637,N_122);
nand U12863 (N_12863,N_5841,N_2840);
nand U12864 (N_12864,N_8911,N_1026);
nor U12865 (N_12865,N_7000,N_9064);
nand U12866 (N_12866,N_7826,N_3332);
and U12867 (N_12867,N_3292,N_2938);
or U12868 (N_12868,N_8678,N_9143);
nand U12869 (N_12869,N_3241,N_8619);
and U12870 (N_12870,N_965,N_7300);
or U12871 (N_12871,N_6616,N_9957);
and U12872 (N_12872,N_1211,N_9303);
or U12873 (N_12873,N_5345,N_1103);
nor U12874 (N_12874,N_2598,N_9088);
nand U12875 (N_12875,N_2856,N_7436);
nand U12876 (N_12876,N_1664,N_5967);
or U12877 (N_12877,N_7998,N_9148);
nor U12878 (N_12878,N_6635,N_8410);
nor U12879 (N_12879,N_2551,N_774);
nor U12880 (N_12880,N_8793,N_4720);
or U12881 (N_12881,N_5492,N_319);
nand U12882 (N_12882,N_6584,N_8550);
xnor U12883 (N_12883,N_6029,N_9251);
nor U12884 (N_12884,N_5336,N_1689);
or U12885 (N_12885,N_7225,N_5123);
nand U12886 (N_12886,N_65,N_2429);
nand U12887 (N_12887,N_7874,N_7368);
nand U12888 (N_12888,N_2999,N_1278);
nand U12889 (N_12889,N_7175,N_1631);
nand U12890 (N_12890,N_8404,N_498);
nor U12891 (N_12891,N_7856,N_5720);
and U12892 (N_12892,N_3823,N_2415);
nor U12893 (N_12893,N_8098,N_697);
nand U12894 (N_12894,N_9332,N_2886);
nand U12895 (N_12895,N_3489,N_2765);
and U12896 (N_12896,N_8086,N_7511);
nor U12897 (N_12897,N_1316,N_9893);
and U12898 (N_12898,N_8936,N_3990);
nor U12899 (N_12899,N_5066,N_96);
nand U12900 (N_12900,N_4273,N_7357);
or U12901 (N_12901,N_6590,N_9240);
nand U12902 (N_12902,N_6170,N_7439);
and U12903 (N_12903,N_3340,N_2300);
or U12904 (N_12904,N_3819,N_1223);
nand U12905 (N_12905,N_3109,N_5162);
nand U12906 (N_12906,N_3000,N_6479);
and U12907 (N_12907,N_1824,N_1099);
and U12908 (N_12908,N_6364,N_9952);
nor U12909 (N_12909,N_4982,N_7985);
or U12910 (N_12910,N_1478,N_3617);
nor U12911 (N_12911,N_2739,N_9752);
and U12912 (N_12912,N_605,N_6580);
or U12913 (N_12913,N_1968,N_1903);
and U12914 (N_12914,N_4545,N_9608);
nor U12915 (N_12915,N_3065,N_7654);
nand U12916 (N_12916,N_8148,N_7510);
and U12917 (N_12917,N_1734,N_9305);
nor U12918 (N_12918,N_522,N_7592);
nor U12919 (N_12919,N_8387,N_8883);
nor U12920 (N_12920,N_1511,N_6677);
nand U12921 (N_12921,N_7607,N_4566);
and U12922 (N_12922,N_3314,N_8389);
or U12923 (N_12923,N_1303,N_5726);
or U12924 (N_12924,N_9635,N_7135);
and U12925 (N_12925,N_3405,N_7324);
nand U12926 (N_12926,N_7500,N_2653);
or U12927 (N_12927,N_5791,N_7577);
nor U12928 (N_12928,N_9369,N_7070);
or U12929 (N_12929,N_2899,N_3635);
and U12930 (N_12930,N_8704,N_6690);
nand U12931 (N_12931,N_7840,N_859);
or U12932 (N_12932,N_8050,N_4085);
nor U12933 (N_12933,N_5685,N_2870);
nor U12934 (N_12934,N_8259,N_3337);
and U12935 (N_12935,N_6125,N_1451);
or U12936 (N_12936,N_6813,N_1298);
and U12937 (N_12937,N_6574,N_2382);
and U12938 (N_12938,N_9013,N_5600);
nor U12939 (N_12939,N_6204,N_9381);
nor U12940 (N_12940,N_7382,N_4260);
nor U12941 (N_12941,N_2362,N_9934);
and U12942 (N_12942,N_9412,N_7634);
or U12943 (N_12943,N_3559,N_7174);
and U12944 (N_12944,N_1805,N_2234);
nand U12945 (N_12945,N_4211,N_5747);
or U12946 (N_12946,N_9910,N_7226);
and U12947 (N_12947,N_6693,N_7085);
or U12948 (N_12948,N_7193,N_9252);
and U12949 (N_12949,N_6791,N_458);
nand U12950 (N_12950,N_9304,N_3358);
or U12951 (N_12951,N_2369,N_2495);
nand U12952 (N_12952,N_7918,N_1748);
nor U12953 (N_12953,N_8752,N_1313);
and U12954 (N_12954,N_3417,N_9425);
nand U12955 (N_12955,N_49,N_4718);
nor U12956 (N_12956,N_8916,N_9161);
nor U12957 (N_12957,N_6077,N_8297);
nand U12958 (N_12958,N_1310,N_6967);
or U12959 (N_12959,N_7911,N_7342);
nand U12960 (N_12960,N_1453,N_4365);
nand U12961 (N_12961,N_2190,N_2375);
nand U12962 (N_12962,N_338,N_696);
or U12963 (N_12963,N_953,N_6067);
nor U12964 (N_12964,N_7811,N_2915);
and U12965 (N_12965,N_3991,N_7566);
and U12966 (N_12966,N_7141,N_7846);
or U12967 (N_12967,N_5479,N_2846);
nor U12968 (N_12968,N_4216,N_9299);
or U12969 (N_12969,N_7707,N_9151);
and U12970 (N_12970,N_9000,N_1699);
or U12971 (N_12971,N_6359,N_505);
or U12972 (N_12972,N_242,N_9201);
nand U12973 (N_12973,N_752,N_9907);
or U12974 (N_12974,N_6291,N_8030);
nand U12975 (N_12975,N_837,N_417);
nor U12976 (N_12976,N_8109,N_6252);
nand U12977 (N_12977,N_5077,N_8904);
and U12978 (N_12978,N_4949,N_2532);
nand U12979 (N_12979,N_1843,N_628);
or U12980 (N_12980,N_8506,N_5462);
nor U12981 (N_12981,N_9069,N_8473);
nor U12982 (N_12982,N_8531,N_842);
or U12983 (N_12983,N_7885,N_6644);
or U12984 (N_12984,N_1822,N_2697);
and U12985 (N_12985,N_4855,N_7258);
nor U12986 (N_12986,N_7246,N_9748);
nor U12987 (N_12987,N_944,N_3752);
nand U12988 (N_12988,N_3428,N_1379);
nor U12989 (N_12989,N_4731,N_4472);
nor U12990 (N_12990,N_7367,N_2964);
or U12991 (N_12991,N_2422,N_8066);
or U12992 (N_12992,N_2825,N_1078);
nor U12993 (N_12993,N_3080,N_1207);
or U12994 (N_12994,N_3131,N_9085);
nand U12995 (N_12995,N_7124,N_1331);
and U12996 (N_12996,N_3485,N_88);
and U12997 (N_12997,N_213,N_7203);
nor U12998 (N_12998,N_7818,N_5185);
nand U12999 (N_12999,N_6218,N_7684);
and U13000 (N_13000,N_3033,N_5005);
nand U13001 (N_13001,N_1018,N_4896);
or U13002 (N_13002,N_8970,N_1362);
nand U13003 (N_13003,N_2216,N_9168);
nand U13004 (N_13004,N_7221,N_4995);
nor U13005 (N_13005,N_7123,N_2548);
or U13006 (N_13006,N_9215,N_6923);
nand U13007 (N_13007,N_4879,N_9025);
or U13008 (N_13008,N_8782,N_2481);
nand U13009 (N_13009,N_1952,N_2809);
nor U13010 (N_13010,N_3451,N_8997);
and U13011 (N_13011,N_2675,N_5892);
nor U13012 (N_13012,N_7599,N_6942);
nor U13013 (N_13013,N_6928,N_5583);
or U13014 (N_13014,N_6567,N_2650);
and U13015 (N_13015,N_9733,N_9591);
or U13016 (N_13016,N_4877,N_4207);
and U13017 (N_13017,N_2098,N_261);
and U13018 (N_13018,N_2398,N_9562);
nand U13019 (N_13019,N_164,N_33);
nand U13020 (N_13020,N_1312,N_9520);
nand U13021 (N_13021,N_8934,N_9038);
or U13022 (N_13022,N_824,N_5512);
nor U13023 (N_13023,N_153,N_8059);
and U13024 (N_13024,N_3882,N_3858);
or U13025 (N_13025,N_2323,N_9485);
or U13026 (N_13026,N_7706,N_6962);
and U13027 (N_13027,N_6534,N_2377);
nor U13028 (N_13028,N_6848,N_9263);
nor U13029 (N_13029,N_6031,N_7809);
and U13030 (N_13030,N_2818,N_8658);
xnor U13031 (N_13031,N_2228,N_9668);
nor U13032 (N_13032,N_7529,N_1986);
or U13033 (N_13033,N_4040,N_1317);
and U13034 (N_13034,N_5906,N_7179);
nor U13035 (N_13035,N_8319,N_295);
or U13036 (N_13036,N_516,N_7037);
nand U13037 (N_13037,N_900,N_5187);
nand U13038 (N_13038,N_6531,N_945);
or U13039 (N_13039,N_4389,N_2492);
nor U13040 (N_13040,N_3544,N_3055);
nand U13041 (N_13041,N_7288,N_5086);
nand U13042 (N_13042,N_3203,N_8469);
nand U13043 (N_13043,N_535,N_7775);
nand U13044 (N_13044,N_8242,N_3731);
or U13045 (N_13045,N_9850,N_4248);
or U13046 (N_13046,N_7150,N_6601);
or U13047 (N_13047,N_7693,N_8174);
or U13048 (N_13048,N_5235,N_8129);
or U13049 (N_13049,N_1242,N_7063);
or U13050 (N_13050,N_1051,N_9058);
or U13051 (N_13051,N_8641,N_8371);
or U13052 (N_13052,N_7792,N_7584);
and U13053 (N_13053,N_6987,N_8669);
nor U13054 (N_13054,N_6351,N_186);
or U13055 (N_13055,N_6484,N_2945);
nor U13056 (N_13056,N_8536,N_526);
nand U13057 (N_13057,N_1265,N_3523);
and U13058 (N_13058,N_7983,N_552);
and U13059 (N_13059,N_7240,N_6829);
and U13060 (N_13060,N_9091,N_6196);
or U13061 (N_13061,N_2661,N_6502);
or U13062 (N_13062,N_7699,N_7662);
and U13063 (N_13063,N_6982,N_7256);
or U13064 (N_13064,N_17,N_2747);
or U13065 (N_13065,N_8938,N_3889);
and U13066 (N_13066,N_4182,N_7773);
and U13067 (N_13067,N_5485,N_2320);
nand U13068 (N_13068,N_9327,N_9955);
nand U13069 (N_13069,N_478,N_3926);
or U13070 (N_13070,N_7237,N_4824);
or U13071 (N_13071,N_2029,N_5062);
nor U13072 (N_13072,N_9977,N_2043);
nor U13073 (N_13073,N_170,N_8128);
nand U13074 (N_13074,N_3439,N_6450);
nand U13075 (N_13075,N_8999,N_4133);
nand U13076 (N_13076,N_9800,N_4642);
nand U13077 (N_13077,N_5215,N_231);
nor U13078 (N_13078,N_2528,N_3908);
and U13079 (N_13079,N_6408,N_7742);
nand U13080 (N_13080,N_9652,N_2773);
or U13081 (N_13081,N_2044,N_3236);
nor U13082 (N_13082,N_3104,N_5564);
and U13083 (N_13083,N_9322,N_3075);
nand U13084 (N_13084,N_7752,N_2246);
or U13085 (N_13085,N_6512,N_2437);
and U13086 (N_13086,N_1777,N_2536);
and U13087 (N_13087,N_4600,N_4633);
nand U13088 (N_13088,N_6796,N_8654);
and U13089 (N_13089,N_3159,N_8946);
nor U13090 (N_13090,N_2771,N_7545);
nand U13091 (N_13091,N_5555,N_5142);
nand U13092 (N_13092,N_5645,N_4128);
nand U13093 (N_13093,N_1597,N_2755);
nand U13094 (N_13094,N_1900,N_4677);
or U13095 (N_13095,N_6014,N_6098);
and U13096 (N_13096,N_2290,N_1372);
nor U13097 (N_13097,N_795,N_4117);
nor U13098 (N_13098,N_5173,N_3515);
nand U13099 (N_13099,N_1261,N_4716);
nand U13100 (N_13100,N_2295,N_8027);
xnor U13101 (N_13101,N_8508,N_4271);
nand U13102 (N_13102,N_3007,N_4630);
nor U13103 (N_13103,N_3923,N_1731);
nand U13104 (N_13104,N_2163,N_4394);
or U13105 (N_13105,N_3812,N_7912);
and U13106 (N_13106,N_5882,N_4457);
and U13107 (N_13107,N_926,N_9765);
nor U13108 (N_13108,N_2748,N_4727);
xnor U13109 (N_13109,N_9172,N_5887);
nor U13110 (N_13110,N_2722,N_7882);
or U13111 (N_13111,N_886,N_8459);
nor U13112 (N_13112,N_4155,N_849);
or U13113 (N_13113,N_3645,N_1151);
nor U13114 (N_13114,N_1804,N_101);
nand U13115 (N_13115,N_2507,N_4159);
and U13116 (N_13116,N_8945,N_4424);
or U13117 (N_13117,N_2005,N_4608);
nor U13118 (N_13118,N_2674,N_7091);
nand U13119 (N_13119,N_5397,N_5654);
or U13120 (N_13120,N_5020,N_2256);
and U13121 (N_13121,N_4481,N_3225);
or U13122 (N_13122,N_8032,N_2946);
or U13123 (N_13123,N_892,N_9873);
nor U13124 (N_13124,N_174,N_3346);
nor U13125 (N_13125,N_5911,N_2588);
nor U13126 (N_13126,N_2857,N_9581);
or U13127 (N_13127,N_6543,N_7490);
or U13128 (N_13128,N_6296,N_7230);
and U13129 (N_13129,N_2078,N_2934);
nand U13130 (N_13130,N_1123,N_9710);
or U13131 (N_13131,N_3382,N_7039);
nor U13132 (N_13132,N_8982,N_3574);
or U13133 (N_13133,N_4559,N_8070);
xnor U13134 (N_13134,N_3977,N_8705);
nor U13135 (N_13135,N_6802,N_3579);
nand U13136 (N_13136,N_6216,N_7953);
and U13137 (N_13137,N_8257,N_9865);
nand U13138 (N_13138,N_4533,N_4950);
nand U13139 (N_13139,N_90,N_6421);
and U13140 (N_13140,N_2979,N_2610);
and U13141 (N_13141,N_2750,N_5556);
and U13142 (N_13142,N_5128,N_5828);
or U13143 (N_13143,N_3943,N_8933);
nand U13144 (N_13144,N_9225,N_5193);
or U13145 (N_13145,N_8744,N_2530);
nand U13146 (N_13146,N_6704,N_3723);
or U13147 (N_13147,N_4832,N_1059);
nor U13148 (N_13148,N_1983,N_5463);
or U13149 (N_13149,N_4076,N_4186);
nor U13150 (N_13150,N_8848,N_97);
nor U13151 (N_13151,N_8556,N_3905);
and U13152 (N_13152,N_4789,N_6712);
nand U13153 (N_13153,N_1751,N_6741);
nor U13154 (N_13154,N_6804,N_2941);
nand U13155 (N_13155,N_2194,N_2014);
nand U13156 (N_13156,N_9506,N_672);
nand U13157 (N_13157,N_7969,N_2746);
nor U13158 (N_13158,N_7081,N_1691);
and U13159 (N_13159,N_5404,N_6808);
nor U13160 (N_13160,N_3049,N_7751);
nand U13161 (N_13161,N_439,N_5689);
or U13162 (N_13162,N_28,N_66);
nor U13163 (N_13163,N_3536,N_3601);
and U13164 (N_13164,N_1365,N_6041);
and U13165 (N_13165,N_9066,N_8111);
and U13166 (N_13166,N_3646,N_358);
and U13167 (N_13167,N_7695,N_7991);
or U13168 (N_13168,N_1304,N_1713);
or U13169 (N_13169,N_4132,N_9187);
nor U13170 (N_13170,N_780,N_6015);
nand U13171 (N_13171,N_7609,N_7533);
and U13172 (N_13172,N_1621,N_2289);
nand U13173 (N_13173,N_1498,N_2418);
nor U13174 (N_13174,N_6191,N_6306);
nor U13175 (N_13175,N_9212,N_2152);
or U13176 (N_13176,N_7528,N_5427);
nand U13177 (N_13177,N_2122,N_6968);
nor U13178 (N_13178,N_8686,N_1302);
nor U13179 (N_13179,N_2613,N_551);
and U13180 (N_13180,N_8953,N_8572);
or U13181 (N_13181,N_7817,N_1999);
nor U13182 (N_13182,N_5401,N_5515);
or U13183 (N_13183,N_8754,N_8312);
nand U13184 (N_13184,N_3945,N_5938);
or U13185 (N_13185,N_5844,N_1973);
and U13186 (N_13186,N_4087,N_6725);
nand U13187 (N_13187,N_4315,N_3763);
or U13188 (N_13188,N_1847,N_2033);
nor U13189 (N_13189,N_6864,N_9645);
nand U13190 (N_13190,N_5259,N_4416);
or U13191 (N_13191,N_5170,N_4704);
and U13192 (N_13192,N_1169,N_5520);
nor U13193 (N_13193,N_2144,N_5870);
nor U13194 (N_13194,N_328,N_8274);
or U13195 (N_13195,N_7588,N_2854);
or U13196 (N_13196,N_2310,N_9415);
or U13197 (N_13197,N_6245,N_3364);
and U13198 (N_13198,N_1246,N_6631);
nor U13199 (N_13199,N_5959,N_3248);
or U13200 (N_13200,N_9595,N_5054);
nor U13201 (N_13201,N_8566,N_7036);
nand U13202 (N_13202,N_8286,N_626);
and U13203 (N_13203,N_7223,N_5933);
nand U13204 (N_13204,N_7540,N_8692);
nand U13205 (N_13205,N_9314,N_6049);
or U13206 (N_13206,N_1423,N_6347);
nor U13207 (N_13207,N_3069,N_5059);
nor U13208 (N_13208,N_4816,N_5659);
or U13209 (N_13209,N_4564,N_425);
nor U13210 (N_13210,N_9950,N_7209);
or U13211 (N_13211,N_4881,N_9003);
and U13212 (N_13212,N_1197,N_4675);
nand U13213 (N_13213,N_485,N_6785);
and U13214 (N_13214,N_6407,N_235);
or U13215 (N_13215,N_7977,N_6950);
nand U13216 (N_13216,N_1160,N_1500);
and U13217 (N_13217,N_3702,N_3745);
nor U13218 (N_13218,N_5302,N_2419);
nand U13219 (N_13219,N_7766,N_3776);
or U13220 (N_13220,N_291,N_8885);
and U13221 (N_13221,N_5616,N_6504);
nand U13222 (N_13222,N_7164,N_7688);
nor U13223 (N_13223,N_6795,N_7712);
and U13224 (N_13224,N_1388,N_6524);
and U13225 (N_13225,N_9301,N_8465);
nand U13226 (N_13226,N_9662,N_3096);
nor U13227 (N_13227,N_9829,N_3317);
or U13228 (N_13228,N_9242,N_6181);
or U13229 (N_13229,N_4011,N_7080);
nor U13230 (N_13230,N_3017,N_7508);
nor U13231 (N_13231,N_3251,N_3176);
or U13232 (N_13232,N_5855,N_1564);
or U13233 (N_13233,N_5407,N_7332);
nand U13234 (N_13234,N_1702,N_3826);
nand U13235 (N_13235,N_4378,N_3892);
or U13236 (N_13236,N_2187,N_6676);
nand U13237 (N_13237,N_783,N_1663);
and U13238 (N_13238,N_5434,N_9682);
and U13239 (N_13239,N_5795,N_1361);
and U13240 (N_13240,N_6241,N_7093);
nand U13241 (N_13241,N_4765,N_9487);
or U13242 (N_13242,N_1131,N_8590);
or U13243 (N_13243,N_5214,N_4935);
or U13244 (N_13244,N_5431,N_6975);
nand U13245 (N_13245,N_3638,N_4681);
nand U13246 (N_13246,N_3728,N_2395);
nand U13247 (N_13247,N_7279,N_2427);
and U13248 (N_13248,N_2988,N_6368);
and U13249 (N_13249,N_7567,N_9570);
nor U13250 (N_13250,N_1315,N_3262);
nand U13251 (N_13251,N_8356,N_2525);
nor U13252 (N_13252,N_3477,N_8092);
nand U13253 (N_13253,N_4084,N_4019);
nand U13254 (N_13254,N_50,N_6656);
or U13255 (N_13255,N_1130,N_8547);
nor U13256 (N_13256,N_9040,N_2337);
nor U13257 (N_13257,N_3538,N_5119);
nand U13258 (N_13258,N_5592,N_5482);
nor U13259 (N_13259,N_5317,N_8396);
and U13260 (N_13260,N_3228,N_3815);
nor U13261 (N_13261,N_4974,N_1001);
nand U13262 (N_13262,N_9259,N_4748);
nand U13263 (N_13263,N_3412,N_6536);
nand U13264 (N_13264,N_2202,N_9180);
and U13265 (N_13265,N_8220,N_2764);
nor U13266 (N_13266,N_2517,N_899);
and U13267 (N_13267,N_7400,N_9779);
nand U13268 (N_13268,N_3144,N_8990);
and U13269 (N_13269,N_7579,N_9336);
nor U13270 (N_13270,N_5502,N_4004);
nor U13271 (N_13271,N_3696,N_215);
nand U13272 (N_13272,N_9717,N_1056);
or U13273 (N_13273,N_6496,N_288);
nand U13274 (N_13274,N_9032,N_7906);
nor U13275 (N_13275,N_6336,N_7420);
or U13276 (N_13276,N_6663,N_7866);
nor U13277 (N_13277,N_312,N_8829);
nor U13278 (N_13278,N_4070,N_8530);
or U13279 (N_13279,N_9070,N_3047);
or U13280 (N_13280,N_5737,N_2296);
or U13281 (N_13281,N_8455,N_3074);
or U13282 (N_13282,N_6365,N_8370);
nor U13283 (N_13283,N_8998,N_4368);
or U13284 (N_13284,N_5677,N_6267);
nor U13285 (N_13285,N_9194,N_21);
or U13286 (N_13286,N_4569,N_1456);
or U13287 (N_13287,N_6930,N_2735);
nand U13288 (N_13288,N_1507,N_9586);
or U13289 (N_13289,N_8450,N_6503);
and U13290 (N_13290,N_8379,N_2379);
or U13291 (N_13291,N_5466,N_5307);
nor U13292 (N_13292,N_4376,N_8824);
nand U13293 (N_13293,N_6441,N_7265);
nand U13294 (N_13294,N_636,N_4208);
nand U13295 (N_13295,N_3307,N_2099);
and U13296 (N_13296,N_9837,N_3644);
or U13297 (N_13297,N_7526,N_4908);
nor U13298 (N_13298,N_7194,N_457);
or U13299 (N_13299,N_9237,N_2211);
nor U13300 (N_13300,N_6716,N_7139);
nand U13301 (N_13301,N_83,N_8398);
and U13302 (N_13302,N_6088,N_9106);
or U13303 (N_13303,N_1552,N_9555);
nand U13304 (N_13304,N_2932,N_6710);
or U13305 (N_13305,N_8873,N_4627);
or U13306 (N_13306,N_1946,N_116);
and U13307 (N_13307,N_4219,N_6559);
nand U13308 (N_13308,N_7812,N_4486);
or U13309 (N_13309,N_1955,N_8300);
and U13310 (N_13310,N_3837,N_6895);
nand U13311 (N_13311,N_942,N_4200);
nand U13312 (N_13312,N_3620,N_9767);
or U13313 (N_13313,N_3291,N_8574);
or U13314 (N_13314,N_9642,N_4436);
nor U13315 (N_13315,N_8234,N_4858);
nand U13316 (N_13316,N_1431,N_1200);
nor U13317 (N_13317,N_5309,N_3642);
nor U13318 (N_13318,N_6934,N_7698);
nand U13319 (N_13319,N_903,N_1741);
nand U13320 (N_13320,N_9433,N_4010);
nor U13321 (N_13321,N_2180,N_4471);
or U13322 (N_13322,N_8438,N_2066);
or U13323 (N_13323,N_977,N_8889);
nand U13324 (N_13324,N_6844,N_6569);
nand U13325 (N_13325,N_2978,N_7560);
and U13326 (N_13326,N_7587,N_9068);
nor U13327 (N_13327,N_5400,N_6182);
and U13328 (N_13328,N_4819,N_3857);
xor U13329 (N_13329,N_9,N_1204);
or U13330 (N_13330,N_6595,N_8294);
nor U13331 (N_13331,N_763,N_8266);
nand U13332 (N_13332,N_1270,N_1178);
nand U13333 (N_13333,N_9393,N_2509);
or U13334 (N_13334,N_8535,N_6977);
and U13335 (N_13335,N_1827,N_4451);
or U13336 (N_13336,N_7666,N_856);
nor U13337 (N_13337,N_7868,N_57);
or U13338 (N_13338,N_5723,N_7232);
or U13339 (N_13339,N_4938,N_4290);
nand U13340 (N_13340,N_2935,N_3709);
or U13341 (N_13341,N_1530,N_1199);
or U13342 (N_13342,N_5514,N_145);
and U13343 (N_13343,N_6160,N_8308);
nor U13344 (N_13344,N_4998,N_264);
xor U13345 (N_13345,N_7635,N_991);
nor U13346 (N_13346,N_1387,N_1605);
nand U13347 (N_13347,N_1609,N_748);
and U13348 (N_13348,N_4370,N_1100);
and U13349 (N_13349,N_4655,N_7335);
nand U13350 (N_13350,N_2689,N_6997);
or U13351 (N_13351,N_8948,N_6851);
nor U13352 (N_13352,N_5245,N_2266);
and U13353 (N_13353,N_3356,N_2193);
xor U13354 (N_13354,N_9819,N_8002);
or U13355 (N_13355,N_2327,N_4429);
nor U13356 (N_13356,N_9131,N_2890);
and U13357 (N_13357,N_4259,N_7797);
or U13358 (N_13358,N_6670,N_1995);
nor U13359 (N_13359,N_8895,N_7652);
or U13360 (N_13360,N_9688,N_3326);
or U13361 (N_13361,N_9326,N_3301);
or U13362 (N_13362,N_5137,N_7585);
nor U13363 (N_13363,N_6615,N_532);
nand U13364 (N_13364,N_8290,N_4323);
nand U13365 (N_13365,N_4859,N_5852);
and U13366 (N_13366,N_9199,N_4782);
nor U13367 (N_13367,N_2254,N_1791);
or U13368 (N_13368,N_9238,N_8110);
nand U13369 (N_13369,N_4813,N_3433);
nor U13370 (N_13370,N_1717,N_9469);
nand U13371 (N_13371,N_3615,N_5861);
nor U13372 (N_13372,N_7020,N_9518);
nand U13373 (N_13373,N_8906,N_4850);
nand U13374 (N_13374,N_1373,N_9024);
nor U13375 (N_13375,N_3875,N_8495);
nor U13376 (N_13376,N_4976,N_8701);
nor U13377 (N_13377,N_4443,N_3737);
nor U13378 (N_13378,N_9972,N_6628);
or U13379 (N_13379,N_4223,N_1152);
nand U13380 (N_13380,N_318,N_7414);
nand U13381 (N_13381,N_2350,N_4754);
nor U13382 (N_13382,N_106,N_4964);
nor U13383 (N_13383,N_7154,N_4041);
or U13384 (N_13384,N_7933,N_7412);
and U13385 (N_13385,N_7788,N_8926);
or U13386 (N_13386,N_9519,N_9015);
nor U13387 (N_13387,N_9945,N_4058);
nand U13388 (N_13388,N_8394,N_1292);
nand U13389 (N_13389,N_9114,N_5916);
nand U13390 (N_13390,N_7869,N_5201);
nand U13391 (N_13391,N_1626,N_8869);
nand U13392 (N_13392,N_7222,N_1926);
nand U13393 (N_13393,N_5693,N_1593);
and U13394 (N_13394,N_1658,N_8795);
nand U13395 (N_13395,N_1747,N_356);
or U13396 (N_13396,N_9435,N_2070);
and U13397 (N_13397,N_2403,N_2570);
and U13398 (N_13398,N_6814,N_4523);
or U13399 (N_13399,N_6812,N_7682);
or U13400 (N_13400,N_4110,N_8988);
nor U13401 (N_13401,N_69,N_6608);
nand U13402 (N_13402,N_2680,N_3534);
nor U13403 (N_13403,N_2271,N_7685);
and U13404 (N_13404,N_6184,N_9090);
or U13405 (N_13405,N_3191,N_9921);
nand U13406 (N_13406,N_1756,N_3367);
xnor U13407 (N_13407,N_120,N_9034);
or U13408 (N_13408,N_9205,N_6047);
nand U13409 (N_13409,N_4423,N_7648);
or U13410 (N_13410,N_9546,N_5075);
and U13411 (N_13411,N_3345,N_6873);
or U13412 (N_13412,N_241,N_6792);
and U13413 (N_13413,N_7774,N_9403);
and U13414 (N_13414,N_3392,N_593);
nor U13415 (N_13415,N_15,N_1141);
nor U13416 (N_13416,N_6721,N_4552);
or U13417 (N_13417,N_5176,N_8856);
or U13418 (N_13418,N_299,N_3056);
nor U13419 (N_13419,N_5364,N_8831);
nand U13420 (N_13420,N_7603,N_4350);
nand U13421 (N_13421,N_7407,N_2897);
and U13422 (N_13422,N_1090,N_3572);
and U13423 (N_13423,N_2622,N_5678);
and U13424 (N_13424,N_7996,N_272);
or U13425 (N_13425,N_8620,N_6914);
nor U13426 (N_13426,N_1910,N_7924);
and U13427 (N_13427,N_5941,N_8785);
or U13428 (N_13428,N_1366,N_9634);
and U13429 (N_13429,N_9983,N_8853);
or U13430 (N_13430,N_1712,N_331);
or U13431 (N_13431,N_5712,N_4568);
or U13432 (N_13432,N_403,N_2210);
and U13433 (N_13433,N_9822,N_2500);
and U13434 (N_13434,N_155,N_9285);
or U13435 (N_13435,N_4335,N_1675);
or U13436 (N_13436,N_3418,N_7155);
or U13437 (N_13437,N_2624,N_2639);
nor U13438 (N_13438,N_2028,N_4373);
nand U13439 (N_13439,N_3359,N_7050);
or U13440 (N_13440,N_4902,N_1541);
and U13441 (N_13441,N_1306,N_2011);
nor U13442 (N_13442,N_2732,N_8303);
nor U13443 (N_13443,N_1695,N_4169);
nand U13444 (N_13444,N_9982,N_9808);
and U13445 (N_13445,N_8225,N_1244);
and U13446 (N_13446,N_2203,N_9134);
nor U13447 (N_13447,N_4037,N_2760);
nor U13448 (N_13448,N_1469,N_5269);
or U13449 (N_13449,N_3361,N_3481);
and U13450 (N_13450,N_9633,N_7350);
or U13451 (N_13451,N_8751,N_150);
nand U13452 (N_13452,N_503,N_8855);
xnor U13453 (N_13453,N_7950,N_6827);
nand U13454 (N_13454,N_2473,N_7902);
and U13455 (N_13455,N_4346,N_4734);
nor U13456 (N_13456,N_8491,N_9973);
and U13457 (N_13457,N_7596,N_2623);
nand U13458 (N_13458,N_1797,N_1783);
or U13459 (N_13459,N_4537,N_4093);
nor U13460 (N_13460,N_3255,N_8691);
and U13461 (N_13461,N_3893,N_5055);
and U13462 (N_13462,N_6620,N_7285);
nand U13463 (N_13463,N_5192,N_9754);
and U13464 (N_13464,N_2956,N_7152);
or U13465 (N_13465,N_1915,N_3062);
nor U13466 (N_13466,N_8427,N_912);
and U13467 (N_13467,N_6283,N_129);
and U13468 (N_13468,N_5593,N_5114);
or U13469 (N_13469,N_8397,N_350);
and U13470 (N_13470,N_9253,N_1458);
and U13471 (N_13471,N_8527,N_9451);
and U13472 (N_13472,N_9722,N_3627);
and U13473 (N_13473,N_1535,N_6865);
nand U13474 (N_13474,N_3474,N_4299);
and U13475 (N_13475,N_3550,N_5994);
and U13476 (N_13476,N_8810,N_819);
or U13477 (N_13477,N_6891,N_5071);
nand U13478 (N_13478,N_7381,N_5500);
and U13479 (N_13479,N_1787,N_7538);
and U13480 (N_13480,N_1617,N_4377);
nand U13481 (N_13481,N_8457,N_3235);
nor U13482 (N_13482,N_7195,N_3419);
or U13483 (N_13483,N_4804,N_2110);
or U13484 (N_13484,N_527,N_4686);
nor U13485 (N_13485,N_2571,N_308);
nor U13486 (N_13486,N_6334,N_5441);
nor U13487 (N_13487,N_2298,N_24);
nor U13488 (N_13488,N_98,N_2200);
nor U13489 (N_13489,N_7177,N_8570);
nor U13490 (N_13490,N_6486,N_6995);
or U13491 (N_13491,N_881,N_4314);
and U13492 (N_13492,N_1927,N_7190);
nor U13493 (N_13493,N_5709,N_6723);
nand U13494 (N_13494,N_8624,N_5042);
nor U13495 (N_13495,N_8235,N_8717);
nand U13496 (N_13496,N_8802,N_7284);
and U13497 (N_13497,N_4268,N_5833);
and U13498 (N_13498,N_3721,N_7627);
nand U13499 (N_13499,N_419,N_8474);
or U13500 (N_13500,N_7308,N_5405);
nor U13501 (N_13501,N_6089,N_7104);
nand U13502 (N_13502,N_3884,N_5539);
or U13503 (N_13503,N_7136,N_7213);
nand U13504 (N_13504,N_2879,N_847);
nor U13505 (N_13505,N_1142,N_6525);
or U13506 (N_13506,N_3429,N_1569);
and U13507 (N_13507,N_603,N_2702);
nor U13508 (N_13508,N_8001,N_8804);
nor U13509 (N_13509,N_5935,N_7749);
or U13510 (N_13510,N_7311,N_3953);
and U13511 (N_13511,N_8117,N_8772);
nor U13512 (N_13512,N_5255,N_2914);
nor U13513 (N_13513,N_3670,N_3698);
and U13514 (N_13514,N_6931,N_4244);
nor U13515 (N_13515,N_9164,N_399);
and U13516 (N_13516,N_9657,N_5191);
nor U13517 (N_13517,N_5705,N_2923);
nor U13518 (N_13518,N_4682,N_5504);
nand U13519 (N_13519,N_62,N_8661);
and U13520 (N_13520,N_1052,N_6605);
nand U13521 (N_13521,N_4705,N_5013);
nor U13522 (N_13522,N_7641,N_2068);
nand U13523 (N_13523,N_4715,N_597);
or U13524 (N_13524,N_4562,N_5144);
nand U13525 (N_13525,N_6259,N_3602);
nand U13526 (N_13526,N_6131,N_2396);
and U13527 (N_13527,N_1449,N_7475);
nor U13528 (N_13528,N_2303,N_6438);
or U13529 (N_13529,N_7772,N_5598);
nor U13530 (N_13530,N_1850,N_7496);
nor U13531 (N_13531,N_9869,N_9022);
nand U13532 (N_13532,N_8735,N_2520);
nand U13533 (N_13533,N_6514,N_994);
or U13534 (N_13534,N_8921,N_8977);
and U13535 (N_13535,N_2351,N_3874);
nand U13536 (N_13536,N_2868,N_2159);
nand U13537 (N_13537,N_550,N_7505);
and U13538 (N_13538,N_3449,N_2232);
nand U13539 (N_13539,N_6020,N_1043);
or U13540 (N_13540,N_5569,N_2664);
and U13541 (N_13541,N_3210,N_3570);
and U13542 (N_13542,N_2192,N_7316);
and U13543 (N_13543,N_9047,N_658);
or U13544 (N_13544,N_668,N_8018);
or U13545 (N_13545,N_6768,N_59);
or U13546 (N_13546,N_1046,N_952);
and U13547 (N_13547,N_4666,N_5078);
nor U13548 (N_13548,N_6515,N_2087);
nor U13549 (N_13549,N_4504,N_2874);
nor U13550 (N_13550,N_4581,N_2638);
nor U13551 (N_13551,N_2458,N_1773);
or U13552 (N_13552,N_2361,N_1813);
nand U13553 (N_13553,N_968,N_5805);
or U13554 (N_13554,N_3628,N_5542);
and U13555 (N_13555,N_3749,N_4796);
nor U13556 (N_13556,N_8578,N_5147);
or U13557 (N_13557,N_5268,N_9400);
and U13558 (N_13558,N_6298,N_4966);
nor U13559 (N_13559,N_5926,N_8346);
or U13560 (N_13560,N_561,N_1294);
nand U13561 (N_13561,N_6485,N_5810);
or U13562 (N_13562,N_9522,N_2813);
nor U13563 (N_13563,N_7075,N_5949);
nor U13564 (N_13564,N_6624,N_6222);
nand U13565 (N_13565,N_4645,N_5284);
or U13566 (N_13566,N_6633,N_5859);
nand U13567 (N_13567,N_4689,N_1279);
and U13568 (N_13568,N_5469,N_2510);
nor U13569 (N_13569,N_3123,N_8278);
or U13570 (N_13570,N_3287,N_1035);
or U13571 (N_13571,N_5773,N_6271);
and U13572 (N_13572,N_8868,N_6339);
nor U13573 (N_13573,N_323,N_10);
and U13574 (N_13574,N_6857,N_2740);
nand U13575 (N_13575,N_342,N_4547);
nor U13576 (N_13576,N_5073,N_791);
or U13577 (N_13577,N_5197,N_4487);
nor U13578 (N_13578,N_8216,N_3759);
or U13579 (N_13579,N_2801,N_571);
nor U13580 (N_13580,N_2900,N_653);
or U13581 (N_13581,N_2796,N_1080);
nor U13582 (N_13582,N_5116,N_8017);
nor U13583 (N_13583,N_776,N_7341);
nor U13584 (N_13584,N_7301,N_4077);
and U13585 (N_13585,N_7068,N_5701);
nand U13586 (N_13586,N_9460,N_5573);
or U13587 (N_13587,N_6655,N_9154);
nor U13588 (N_13588,N_2611,N_1371);
or U13589 (N_13589,N_8233,N_9757);
and U13590 (N_13590,N_4098,N_6232);
nand U13591 (N_13591,N_5168,N_2496);
or U13592 (N_13592,N_4002,N_721);
and U13593 (N_13593,N_4044,N_6249);
or U13594 (N_13594,N_5264,N_191);
or U13595 (N_13595,N_1939,N_4648);
nor U13596 (N_13596,N_9489,N_7739);
and U13597 (N_13597,N_6161,N_3493);
or U13598 (N_13598,N_7502,N_3895);
or U13599 (N_13599,N_7645,N_1084);
nor U13600 (N_13600,N_5787,N_8318);
and U13601 (N_13601,N_5543,N_2378);
and U13602 (N_13602,N_6936,N_5046);
and U13603 (N_13603,N_855,N_6786);
or U13604 (N_13604,N_5874,N_8169);
nand U13605 (N_13605,N_2620,N_5340);
nor U13606 (N_13606,N_8151,N_2544);
nand U13607 (N_13607,N_9368,N_5008);
nor U13608 (N_13608,N_3066,N_9871);
nor U13609 (N_13609,N_8900,N_9405);
and U13610 (N_13610,N_1670,N_6217);
or U13611 (N_13611,N_5651,N_2521);
nand U13612 (N_13612,N_949,N_2659);
nand U13613 (N_13613,N_7832,N_4341);
nor U13614 (N_13614,N_477,N_4316);
or U13615 (N_13615,N_3921,N_9310);
and U13616 (N_13616,N_2450,N_4983);
or U13617 (N_13617,N_8712,N_4698);
nand U13618 (N_13618,N_1009,N_7519);
nor U13619 (N_13619,N_2235,N_3740);
or U13620 (N_13620,N_8452,N_392);
and U13621 (N_13621,N_667,N_6911);
or U13622 (N_13622,N_1222,N_3051);
and U13623 (N_13623,N_4632,N_86);
nor U13624 (N_13624,N_8246,N_9537);
nor U13625 (N_13625,N_8079,N_6983);
nor U13626 (N_13626,N_1189,N_3133);
nor U13627 (N_13627,N_8492,N_3447);
nor U13628 (N_13628,N_1598,N_9486);
or U13629 (N_13629,N_2001,N_882);
and U13630 (N_13630,N_7658,N_5708);
nand U13631 (N_13631,N_736,N_3268);
or U13632 (N_13632,N_6980,N_1019);
and U13633 (N_13633,N_305,N_3734);
and U13634 (N_13634,N_8409,N_9612);
and U13635 (N_13635,N_9512,N_6012);
nand U13636 (N_13636,N_5501,N_3402);
or U13637 (N_13637,N_5335,N_6652);
nor U13638 (N_13638,N_6264,N_3510);
nor U13639 (N_13639,N_9130,N_5745);
nand U13640 (N_13640,N_1389,N_1235);
nor U13641 (N_13641,N_1050,N_9228);
xnor U13642 (N_13642,N_8503,N_9762);
nand U13643 (N_13643,N_8184,N_5838);
or U13644 (N_13644,N_2128,N_8085);
nor U13645 (N_13645,N_4999,N_7741);
or U13646 (N_13646,N_3186,N_2201);
and U13647 (N_13647,N_6428,N_9350);
nand U13648 (N_13648,N_3302,N_9442);
nor U13649 (N_13649,N_2452,N_4885);
nand U13650 (N_13650,N_1180,N_4418);
or U13651 (N_13651,N_2089,N_983);
nand U13652 (N_13652,N_982,N_6369);
and U13653 (N_13653,N_2268,N_2220);
and U13654 (N_13654,N_9713,N_746);
nor U13655 (N_13655,N_9598,N_5891);
and U13656 (N_13656,N_1913,N_7384);
and U13657 (N_13657,N_7268,N_4103);
or U13658 (N_13658,N_2446,N_2015);
and U13659 (N_13659,N_4360,N_1144);
nor U13660 (N_13660,N_6174,N_5506);
or U13661 (N_13661,N_4759,N_1251);
and U13662 (N_13662,N_6370,N_7003);
or U13663 (N_13663,N_6838,N_1784);
or U13664 (N_13664,N_7999,N_5575);
nor U13665 (N_13665,N_4946,N_693);
nor U13666 (N_13666,N_3218,N_2909);
nor U13667 (N_13667,N_4956,N_1494);
nand U13668 (N_13668,N_7228,N_6101);
nand U13669 (N_13669,N_4369,N_7862);
and U13670 (N_13670,N_1775,N_2069);
nor U13671 (N_13671,N_9874,N_4198);
nor U13672 (N_13672,N_4506,N_9659);
nor U13673 (N_13673,N_8034,N_7280);
nand U13674 (N_13674,N_4690,N_7944);
or U13675 (N_13675,N_1931,N_1989);
or U13676 (N_13676,N_9745,N_1949);
nand U13677 (N_13677,N_7499,N_5827);
or U13678 (N_13678,N_2138,N_2189);
and U13679 (N_13679,N_375,N_7690);
or U13680 (N_13680,N_1062,N_1484);
or U13681 (N_13681,N_9536,N_7356);
nand U13682 (N_13682,N_6613,N_3318);
and U13683 (N_13683,N_5817,N_4650);
and U13684 (N_13684,N_4495,N_4626);
nand U13685 (N_13685,N_469,N_7956);
and U13686 (N_13686,N_3020,N_41);
or U13687 (N_13687,N_9472,N_2758);
nor U13688 (N_13688,N_1726,N_3625);
and U13689 (N_13689,N_4820,N_3249);
and U13690 (N_13690,N_2240,N_5103);
nor U13691 (N_13691,N_2359,N_8501);
nand U13692 (N_13692,N_2058,N_6961);
nor U13693 (N_13693,N_4320,N_6671);
nand U13694 (N_13694,N_6392,N_9235);
or U13695 (N_13695,N_387,N_7113);
nand U13696 (N_13696,N_2597,N_6910);
or U13697 (N_13697,N_3010,N_1958);
nand U13698 (N_13698,N_193,N_8307);
nor U13699 (N_13699,N_1668,N_4673);
nor U13700 (N_13700,N_8513,N_9016);
nor U13701 (N_13701,N_1895,N_2105);
nor U13702 (N_13702,N_8179,N_6859);
and U13703 (N_13703,N_7834,N_2352);
and U13704 (N_13704,N_8025,N_750);
nor U13705 (N_13705,N_6978,N_8882);
nor U13706 (N_13706,N_4141,N_4173);
or U13707 (N_13707,N_6137,N_6764);
nand U13708 (N_13708,N_7126,N_4493);
nand U13709 (N_13709,N_3870,N_5611);
nor U13710 (N_13710,N_771,N_333);
and U13711 (N_13711,N_8967,N_3231);
nor U13712 (N_13712,N_670,N_2706);
nor U13713 (N_13713,N_5626,N_9264);
nor U13714 (N_13714,N_6778,N_2841);
nor U13715 (N_13715,N_7461,N_8512);
or U13716 (N_13716,N_2671,N_9345);
or U13717 (N_13717,N_2550,N_8035);
nand U13718 (N_13718,N_110,N_889);
and U13719 (N_13719,N_989,N_7745);
or U13720 (N_13720,N_2560,N_9102);
and U13721 (N_13721,N_3904,N_1427);
nand U13722 (N_13722,N_7552,N_5764);
or U13723 (N_13723,N_4240,N_4431);
and U13724 (N_13724,N_717,N_7208);
nor U13725 (N_13725,N_3006,N_5421);
or U13726 (N_13726,N_1206,N_3150);
nand U13727 (N_13727,N_5406,N_592);
nand U13728 (N_13728,N_1448,N_1752);
or U13729 (N_13729,N_1221,N_2526);
or U13730 (N_13730,N_4344,N_5968);
or U13731 (N_13731,N_5001,N_7515);
and U13732 (N_13732,N_4800,N_1054);
or U13733 (N_13733,N_4597,N_4589);
nand U13734 (N_13734,N_8577,N_1754);
nor U13735 (N_13735,N_8172,N_4651);
or U13736 (N_13736,N_5992,N_9527);
nor U13737 (N_13737,N_5458,N_6284);
and U13738 (N_13738,N_8331,N_3667);
and U13739 (N_13739,N_5985,N_7760);
or U13740 (N_13740,N_3222,N_8044);
and U13741 (N_13741,N_3669,N_3630);
nand U13742 (N_13742,N_7935,N_621);
and U13743 (N_13743,N_807,N_7762);
or U13744 (N_13744,N_7785,N_1320);
or U13745 (N_13745,N_4826,N_8994);
nor U13746 (N_13746,N_1028,N_5715);
nand U13747 (N_13747,N_8773,N_9346);
and U13748 (N_13748,N_6683,N_9880);
nand U13749 (N_13749,N_7871,N_9718);
nand U13750 (N_13750,N_294,N_2842);
nor U13751 (N_13751,N_8923,N_2059);
nand U13752 (N_13752,N_1212,N_660);
nor U13753 (N_13753,N_6903,N_8004);
or U13754 (N_13754,N_8013,N_9795);
nor U13755 (N_13755,N_9744,N_6227);
nand U13756 (N_13756,N_6055,N_4288);
or U13757 (N_13757,N_4166,N_5955);
nand U13758 (N_13758,N_4856,N_2824);
or U13759 (N_13759,N_6172,N_6422);
nand U13760 (N_13760,N_7227,N_2556);
and U13761 (N_13761,N_7431,N_8564);
and U13762 (N_13762,N_9676,N_3639);
nand U13763 (N_13763,N_9967,N_7371);
or U13764 (N_13764,N_4822,N_8084);
nand U13765 (N_13765,N_6591,N_9896);
nor U13766 (N_13766,N_4498,N_8838);
or U13767 (N_13767,N_8153,N_1513);
nor U13768 (N_13768,N_6068,N_4332);
nor U13769 (N_13769,N_873,N_1176);
nor U13770 (N_13770,N_1576,N_8375);
or U13771 (N_13771,N_5377,N_1547);
or U13772 (N_13772,N_7160,N_9889);
and U13773 (N_13773,N_4213,N_5460);
and U13774 (N_13774,N_5036,N_2962);
nand U13775 (N_13775,N_6908,N_8061);
or U13776 (N_13776,N_466,N_7275);
or U13777 (N_13777,N_7819,N_7793);
nor U13778 (N_13778,N_4432,N_798);
and U13779 (N_13779,N_3209,N_2238);
nand U13780 (N_13780,N_6951,N_455);
and U13781 (N_13781,N_1767,N_1461);
nor U13782 (N_13782,N_462,N_2604);
nor U13783 (N_13783,N_3793,N_4514);
nor U13784 (N_13784,N_9239,N_5306);
and U13785 (N_13785,N_4104,N_2612);
or U13786 (N_13786,N_6556,N_9379);
and U13787 (N_13787,N_5027,N_1908);
or U13788 (N_13788,N_6825,N_4538);
nor U13789 (N_13789,N_7346,N_9648);
nor U13790 (N_13790,N_1322,N_4621);
nand U13791 (N_13791,N_6876,N_8734);
nand U13792 (N_13792,N_566,N_5628);
and U13793 (N_13793,N_8606,N_9834);
nor U13794 (N_13794,N_933,N_4732);
and U13795 (N_13795,N_1771,N_3525);
and U13796 (N_13796,N_2728,N_5232);
nand U13797 (N_13797,N_3949,N_9176);
nor U13798 (N_13798,N_4903,N_4136);
nand U13799 (N_13799,N_1982,N_5221);
nand U13800 (N_13800,N_479,N_7802);
nand U13801 (N_13801,N_9605,N_7509);
or U13802 (N_13802,N_2635,N_941);
or U13803 (N_13803,N_1433,N_6412);
and U13804 (N_13804,N_6582,N_1548);
nand U13805 (N_13805,N_1182,N_2208);
nand U13806 (N_13806,N_6905,N_9232);
nand U13807 (N_13807,N_5079,N_3290);
or U13808 (N_13808,N_1571,N_467);
and U13809 (N_13809,N_3849,N_3280);
nand U13810 (N_13810,N_784,N_7419);
or U13811 (N_13811,N_2970,N_9426);
and U13812 (N_13812,N_6143,N_3464);
nand U13813 (N_13813,N_1024,N_3116);
or U13814 (N_13814,N_9902,N_3269);
nand U13815 (N_13815,N_8366,N_5167);
nand U13816 (N_13816,N_7951,N_2504);
nand U13817 (N_13817,N_1613,N_8196);
nor U13818 (N_13818,N_1340,N_2564);
or U13819 (N_13819,N_6233,N_4744);
nand U13820 (N_13820,N_9218,N_9096);
nor U13821 (N_13821,N_8014,N_9414);
or U13822 (N_13822,N_4082,N_9904);
or U13823 (N_13823,N_2593,N_556);
or U13824 (N_13824,N_36,N_2302);
or U13825 (N_13825,N_7184,N_4134);
or U13826 (N_13826,N_2954,N_9852);
and U13827 (N_13827,N_7789,N_3779);
nor U13828 (N_13828,N_861,N_4501);
and U13829 (N_13829,N_6214,N_3079);
nor U13830 (N_13830,N_4154,N_8650);
nor U13831 (N_13831,N_9055,N_7898);
and U13832 (N_13832,N_7137,N_9686);
and U13833 (N_13833,N_1081,N_9550);
and U13834 (N_13834,N_9671,N_9438);
nand U13835 (N_13835,N_5624,N_8724);
nor U13836 (N_13836,N_3329,N_2371);
or U13837 (N_13837,N_9986,N_7437);
nand U13838 (N_13838,N_6583,N_501);
nand U13839 (N_13839,N_165,N_3535);
nand U13840 (N_13840,N_9030,N_4193);
nor U13841 (N_13841,N_1192,N_9885);
and U13842 (N_13842,N_7331,N_8132);
nand U13843 (N_13843,N_870,N_1701);
nand U13844 (N_13844,N_6270,N_3263);
or U13845 (N_13845,N_1907,N_2100);
and U13846 (N_13846,N_461,N_5679);
nand U13847 (N_13847,N_2676,N_9386);
or U13848 (N_13848,N_6540,N_5877);
nor U13849 (N_13849,N_6762,N_2021);
nand U13850 (N_13850,N_8261,N_9077);
and U13851 (N_13851,N_7997,N_3958);
and U13852 (N_13852,N_9926,N_2304);
nand U13853 (N_13853,N_5465,N_684);
and U13854 (N_13854,N_3771,N_6832);
nand U13855 (N_13855,N_4071,N_5687);
and U13856 (N_13856,N_9458,N_1410);
nand U13857 (N_13857,N_3526,N_187);
and U13858 (N_13858,N_8697,N_1529);
and U13859 (N_13859,N_4697,N_6718);
or U13860 (N_13860,N_6419,N_3711);
and U13861 (N_13861,N_3863,N_2698);
nor U13862 (N_13862,N_4531,N_238);
nor U13863 (N_13863,N_6253,N_70);
nor U13864 (N_13864,N_8135,N_7041);
nor U13865 (N_13865,N_4191,N_2053);
nor U13866 (N_13866,N_7214,N_9052);
nand U13867 (N_13867,N_5194,N_4623);
and U13868 (N_13868,N_3411,N_9576);
nand U13869 (N_13869,N_869,N_3972);
and U13870 (N_13870,N_4585,N_7130);
nand U13871 (N_13871,N_2267,N_5050);
nor U13872 (N_13872,N_3311,N_7255);
nor U13873 (N_13873,N_2878,N_5739);
or U13874 (N_13874,N_5704,N_2714);
nor U13875 (N_13875,N_9390,N_3381);
nor U13876 (N_13876,N_2392,N_2048);
nor U13877 (N_13877,N_2872,N_5669);
or U13878 (N_13878,N_4511,N_8899);
nor U13879 (N_13879,N_4366,N_2869);
or U13880 (N_13880,N_6658,N_5772);
or U13881 (N_13881,N_8767,N_6021);
and U13882 (N_13882,N_6949,N_9669);
and U13883 (N_13883,N_5919,N_4560);
nand U13884 (N_13884,N_1835,N_5845);
nor U13885 (N_13885,N_7964,N_30);
or U13886 (N_13886,N_1537,N_2270);
nand U13887 (N_13887,N_5254,N_9771);
nand U13888 (N_13888,N_6018,N_4319);
and U13889 (N_13889,N_7325,N_6729);
nor U13890 (N_13890,N_7952,N_7504);
or U13891 (N_13891,N_2206,N_8221);
nand U13892 (N_13892,N_192,N_8742);
nand U13893 (N_13893,N_5314,N_5567);
nand U13894 (N_13894,N_8329,N_3147);
nor U13895 (N_13895,N_5324,N_5122);
nand U13896 (N_13896,N_297,N_6904);
nand U13897 (N_13897,N_9297,N_9582);
xor U13898 (N_13898,N_5297,N_9276);
nand U13899 (N_13899,N_1919,N_1694);
nand U13900 (N_13900,N_1618,N_9766);
nand U13901 (N_13901,N_8937,N_1509);
nor U13902 (N_13902,N_9583,N_332);
or U13903 (N_13903,N_6530,N_3746);
nor U13904 (N_13904,N_1828,N_1007);
nand U13905 (N_13905,N_2293,N_4927);
nand U13906 (N_13906,N_3488,N_8223);
or U13907 (N_13907,N_3160,N_5439);
and U13908 (N_13908,N_1407,N_5304);
and U13909 (N_13909,N_8323,N_7415);
nand U13910 (N_13910,N_3509,N_9277);
nand U13911 (N_13911,N_2804,N_2976);
nand U13912 (N_13912,N_4122,N_9965);
nand U13913 (N_13913,N_9858,N_7546);
or U13914 (N_13914,N_9697,N_6979);
or U13915 (N_13915,N_2061,N_1929);
nor U13916 (N_13916,N_7900,N_749);
and U13917 (N_13917,N_1350,N_2943);
or U13918 (N_13918,N_985,N_6416);
or U13919 (N_13919,N_6092,N_7791);
or U13920 (N_13920,N_2184,N_9991);
or U13921 (N_13921,N_4343,N_8880);
nand U13922 (N_13922,N_9457,N_5459);
nor U13923 (N_13923,N_9807,N_3689);
nand U13924 (N_13924,N_4008,N_8339);
nand U13925 (N_13925,N_5771,N_4102);
nand U13926 (N_13926,N_5622,N_6110);
or U13927 (N_13927,N_5313,N_8497);
nand U13928 (N_13928,N_2778,N_2737);
nor U13929 (N_13929,N_8716,N_9823);
nor U13930 (N_13930,N_932,N_9929);
nor U13931 (N_13931,N_1883,N_6418);
or U13932 (N_13932,N_8354,N_7958);
nand U13933 (N_13933,N_5825,N_6952);
nand U13934 (N_13934,N_3416,N_9348);
or U13935 (N_13935,N_2952,N_2843);
and U13936 (N_13936,N_3714,N_9275);
nor U13937 (N_13937,N_4634,N_391);
nor U13938 (N_13938,N_2262,N_6487);
and U13939 (N_13939,N_7299,N_3259);
nor U13940 (N_13940,N_5387,N_3221);
nor U13941 (N_13941,N_2401,N_9848);
nand U13942 (N_13942,N_7183,N_3438);
and U13943 (N_13943,N_4160,N_8559);
and U13944 (N_13944,N_2554,N_3813);
nor U13945 (N_13945,N_5991,N_1351);
and U13946 (N_13946,N_2264,N_5432);
nor U13947 (N_13947,N_5450,N_9706);
nor U13948 (N_13948,N_3868,N_8482);
and U13949 (N_13949,N_8683,N_3237);
nand U13950 (N_13950,N_5744,N_3571);
or U13951 (N_13951,N_9246,N_2199);
and U13952 (N_13952,N_5085,N_6279);
and U13953 (N_13953,N_9155,N_1960);
nor U13954 (N_13954,N_1570,N_2566);
nor U13955 (N_13955,N_5665,N_7411);
or U13956 (N_13956,N_1492,N_2787);
or U13957 (N_13957,N_6420,N_4265);
and U13958 (N_13958,N_2955,N_1595);
nand U13959 (N_13959,N_8411,N_7686);
and U13960 (N_13960,N_4474,N_9734);
nand U13961 (N_13961,N_4108,N_7735);
xnor U13962 (N_13962,N_1696,N_8296);
xor U13963 (N_13963,N_5653,N_6473);
or U13964 (N_13964,N_735,N_1187);
xor U13965 (N_13965,N_2090,N_422);
nand U13966 (N_13966,N_4548,N_2311);
and U13967 (N_13967,N_9940,N_2137);
and U13968 (N_13968,N_2694,N_883);
nand U13969 (N_13969,N_2853,N_1063);
and U13970 (N_13970,N_6193,N_6625);
nor U13971 (N_13971,N_2113,N_258);
nor U13972 (N_13972,N_365,N_3008);
and U13973 (N_13973,N_2531,N_4915);
or U13974 (N_13974,N_1406,N_9428);
or U13975 (N_13975,N_5785,N_8324);
nand U13976 (N_13976,N_9768,N_720);
nor U13977 (N_13977,N_5286,N_1238);
nand U13978 (N_13978,N_7663,N_786);
nand U13979 (N_13979,N_2807,N_9677);
or U13980 (N_13980,N_3616,N_4379);
nand U13981 (N_13981,N_917,N_2471);
and U13982 (N_13982,N_8581,N_7163);
or U13983 (N_13983,N_3545,N_4636);
nor U13984 (N_13984,N_8340,N_8316);
nand U13985 (N_13985,N_1039,N_616);
or U13986 (N_13986,N_223,N_2736);
nand U13987 (N_13987,N_6648,N_1594);
nand U13988 (N_13988,N_2754,N_2097);
nor U13989 (N_13989,N_6346,N_205);
nand U13990 (N_13990,N_3897,N_8912);
or U13991 (N_13991,N_3103,N_5586);
or U13992 (N_13992,N_3852,N_4588);
nand U13993 (N_13993,N_3434,N_8126);
or U13994 (N_13994,N_6135,N_1898);
or U13995 (N_13995,N_5731,N_7029);
nor U13996 (N_13996,N_5105,N_2503);
or U13997 (N_13997,N_2249,N_1625);
or U13998 (N_13998,N_2590,N_7485);
or U13999 (N_13999,N_4894,N_1531);
or U14000 (N_14000,N_9121,N_5070);
nor U14001 (N_14001,N_2404,N_9923);
nor U14002 (N_14002,N_9856,N_2858);
and U14003 (N_14003,N_8232,N_7660);
and U14004 (N_14004,N_9609,N_3987);
or U14005 (N_14005,N_3948,N_3484);
nand U14006 (N_14006,N_3232,N_4643);
or U14007 (N_14007,N_1865,N_8090);
and U14008 (N_14008,N_6340,N_2498);
nand U14009 (N_14009,N_591,N_9906);
and U14010 (N_14010,N_3775,N_9704);
nand U14011 (N_14011,N_9619,N_3097);
and U14012 (N_14012,N_8088,N_2756);
nor U14013 (N_14013,N_3092,N_531);
nand U14014 (N_14014,N_8656,N_7691);
or U14015 (N_14015,N_781,N_326);
and U14016 (N_14016,N_6594,N_9862);
nor U14017 (N_14017,N_4353,N_9916);
nand U14018 (N_14018,N_8733,N_7312);
nor U14019 (N_14019,N_4162,N_3115);
nand U14020 (N_14020,N_2339,N_2552);
nor U14021 (N_14021,N_108,N_2514);
nor U14022 (N_14022,N_538,N_8726);
nand U14023 (N_14023,N_7261,N_5605);
or U14024 (N_14024,N_6732,N_2832);
nor U14025 (N_14025,N_1920,N_3983);
nand U14026 (N_14026,N_695,N_5759);
or U14027 (N_14027,N_7671,N_8481);
nor U14028 (N_14028,N_4249,N_7974);
or U14029 (N_14029,N_3715,N_7878);
nor U14030 (N_14030,N_9128,N_1517);
nand U14031 (N_14031,N_871,N_3606);
and U14032 (N_14032,N_339,N_3738);
nand U14033 (N_14033,N_2114,N_6411);
nand U14034 (N_14034,N_1978,N_8807);
or U14035 (N_14035,N_8425,N_9558);
nand U14036 (N_14036,N_8189,N_4458);
or U14037 (N_14037,N_6016,N_8122);
and U14038 (N_14038,N_1556,N_7449);
nor U14039 (N_14039,N_1959,N_5174);
or U14040 (N_14040,N_6330,N_8378);
nor U14041 (N_14041,N_7600,N_1744);
or U14042 (N_14042,N_1801,N_1889);
and U14043 (N_14043,N_996,N_4975);
and U14044 (N_14044,N_5266,N_8087);
nand U14045 (N_14045,N_1336,N_2383);
or U14046 (N_14046,N_2743,N_9396);
or U14047 (N_14047,N_8245,N_5806);
nand U14048 (N_14048,N_9097,N_5965);
nor U14049 (N_14049,N_2663,N_6645);
and U14050 (N_14050,N_5166,N_5585);
nor U14051 (N_14051,N_4028,N_7687);
nand U14052 (N_14052,N_5135,N_9101);
nor U14053 (N_14053,N_8237,N_6414);
or U14054 (N_14054,N_4854,N_8859);
or U14055 (N_14055,N_7828,N_622);
and U14056 (N_14056,N_5711,N_8644);
nor U14057 (N_14057,N_9554,N_58);
or U14058 (N_14058,N_2083,N_7639);
and U14059 (N_14059,N_4519,N_9517);
and U14060 (N_14060,N_6617,N_1231);
nor U14061 (N_14061,N_6564,N_3146);
or U14062 (N_14062,N_9724,N_5518);
or U14063 (N_14063,N_1015,N_9483);
and U14064 (N_14064,N_4764,N_412);
nor U14065 (N_14065,N_9758,N_390);
and U14066 (N_14066,N_4174,N_5430);
and U14067 (N_14067,N_7180,N_3257);
and U14068 (N_14068,N_7327,N_9515);
or U14069 (N_14069,N_7726,N_9281);
nor U14070 (N_14070,N_3050,N_2258);
nor U14071 (N_14071,N_4206,N_4276);
and U14072 (N_14072,N_6734,N_6085);
and U14073 (N_14073,N_3963,N_1338);
nand U14074 (N_14074,N_5873,N_8466);
nand U14075 (N_14075,N_492,N_5940);
nand U14076 (N_14076,N_5394,N_3674);
nor U14077 (N_14077,N_2557,N_585);
nand U14078 (N_14078,N_1239,N_6263);
nor U14079 (N_14079,N_8929,N_6390);
nand U14080 (N_14080,N_898,N_8601);
nand U14081 (N_14081,N_67,N_9958);
nand U14082 (N_14082,N_4348,N_5315);
nand U14083 (N_14083,N_2223,N_4109);
and U14084 (N_14084,N_8776,N_578);
or U14085 (N_14085,N_2357,N_5643);
or U14086 (N_14086,N_2393,N_9167);
nand U14087 (N_14087,N_2880,N_1157);
nand U14088 (N_14088,N_9806,N_2831);
nor U14089 (N_14089,N_6501,N_3328);
or U14090 (N_14090,N_2559,N_8758);
nand U14091 (N_14091,N_9566,N_3919);
nand U14092 (N_14092,N_1076,N_2866);
nand U14093 (N_14093,N_5923,N_5885);
nor U14094 (N_14094,N_6900,N_3798);
nand U14095 (N_14095,N_9315,N_2994);
or U14096 (N_14096,N_9133,N_7291);
or U14097 (N_14097,N_5917,N_4550);
or U14098 (N_14098,N_8422,N_4452);
and U14099 (N_14099,N_5717,N_7457);
nand U14100 (N_14100,N_3704,N_6853);
or U14101 (N_14101,N_504,N_599);
nand U14102 (N_14102,N_3102,N_4269);
nand U14103 (N_14103,N_6964,N_9278);
nor U14104 (N_14104,N_6198,N_3581);
or U14105 (N_14105,N_7103,N_4427);
nand U14106 (N_14106,N_710,N_9185);
or U14107 (N_14107,N_5256,N_6171);
and U14108 (N_14108,N_8045,N_853);
and U14109 (N_14109,N_4742,N_4888);
nor U14110 (N_14110,N_9429,N_5925);
or U14111 (N_14111,N_5603,N_904);
nand U14112 (N_14112,N_6521,N_9629);
or U14113 (N_14113,N_8621,N_6592);
nand U14114 (N_14114,N_3125,N_4557);
and U14115 (N_14115,N_5087,N_7462);
nor U14116 (N_14116,N_5682,N_3918);
or U14117 (N_14117,N_7728,N_7060);
nand U14118 (N_14118,N_7642,N_8414);
nor U14119 (N_14119,N_7443,N_404);
nor U14120 (N_14120,N_2827,N_1619);
and U14121 (N_14121,N_4101,N_959);
or U14122 (N_14122,N_3797,N_141);
and U14123 (N_14123,N_3528,N_6156);
and U14124 (N_14124,N_7306,N_2987);
nand U14125 (N_14125,N_7893,N_4371);
and U14126 (N_14126,N_6082,N_8672);
or U14127 (N_14127,N_6278,N_5830);
nand U14128 (N_14128,N_7562,N_6261);
and U14129 (N_14129,N_8808,N_5774);
nor U14130 (N_14130,N_3649,N_2745);
and U14131 (N_14131,N_6091,N_8774);
and U14132 (N_14132,N_5790,N_8596);
nor U14133 (N_14133,N_6960,N_3729);
nor U14134 (N_14134,N_6046,N_7837);
or U14135 (N_14135,N_8979,N_9222);
and U14136 (N_14136,N_5052,N_6753);
or U14137 (N_14137,N_9998,N_3542);
xor U14138 (N_14138,N_8845,N_2990);
or U14139 (N_14139,N_9260,N_7040);
nand U14140 (N_14140,N_7615,N_1437);
and U14141 (N_14141,N_1677,N_9362);
nor U14142 (N_14142,N_2993,N_9146);
and U14143 (N_14143,N_608,N_9339);
nor U14144 (N_14144,N_1125,N_4462);
nand U14145 (N_14145,N_3831,N_9656);
nor U14146 (N_14146,N_1367,N_6128);
nor U14147 (N_14147,N_2997,N_1109);
nor U14148 (N_14148,N_7984,N_661);
or U14149 (N_14149,N_5426,N_3196);
or U14150 (N_14150,N_7848,N_6254);
nor U14151 (N_14151,N_5420,N_4624);
nand U14152 (N_14152,N_8664,N_9513);
or U14153 (N_14153,N_1928,N_4224);
nand U14154 (N_14154,N_4901,N_3003);
nand U14155 (N_14155,N_2626,N_4610);
or U14156 (N_14156,N_3242,N_4420);
nand U14157 (N_14157,N_5954,N_4048);
and U14158 (N_14158,N_4658,N_149);
nor U14159 (N_14159,N_6632,N_4068);
or U14160 (N_14160,N_4584,N_3380);
or U14161 (N_14161,N_102,N_5946);
and U14162 (N_14162,N_206,N_1093);
or U14163 (N_14163,N_5328,N_3539);
and U14164 (N_14164,N_5776,N_2776);
or U14165 (N_14165,N_1878,N_4818);
nand U14166 (N_14166,N_731,N_5821);
nor U14167 (N_14167,N_1964,N_1241);
nor U14168 (N_14168,N_794,N_5647);
nor U14169 (N_14169,N_9903,N_3240);
or U14170 (N_14170,N_3828,N_3342);
and U14171 (N_14171,N_9407,N_6994);
nand U14172 (N_14172,N_5067,N_1932);
nor U14173 (N_14173,N_5017,N_6262);
and U14174 (N_14174,N_6316,N_6935);
nor U14175 (N_14175,N_2074,N_2908);
nor U14176 (N_14176,N_9545,N_7767);
or U14177 (N_14177,N_4318,N_4131);
or U14178 (N_14178,N_7295,N_1055);
nand U14179 (N_14179,N_8166,N_4575);
and U14180 (N_14180,N_7286,N_6124);
and U14181 (N_14181,N_5293,N_3944);
nor U14182 (N_14182,N_4233,N_6393);
nand U14183 (N_14183,N_4631,N_3042);
nand U14184 (N_14184,N_4825,N_7013);
or U14185 (N_14185,N_3848,N_4907);
nor U14186 (N_14186,N_5757,N_3379);
nor U14187 (N_14187,N_9076,N_3623);
or U14188 (N_14188,N_7945,N_9674);
or U14189 (N_14189,N_3757,N_826);
and U14190 (N_14190,N_2165,N_6052);
nand U14191 (N_14191,N_6817,N_5904);
nor U14192 (N_14192,N_3400,N_2585);
nor U14193 (N_14193,N_434,N_6739);
and U14194 (N_14194,N_5875,N_4295);
nor U14195 (N_14195,N_8769,N_5239);
or U14196 (N_14196,N_4205,N_5690);
or U14197 (N_14197,N_1346,N_2609);
or U14198 (N_14198,N_7665,N_9249);
nor U14199 (N_14199,N_1225,N_475);
or U14200 (N_14200,N_6352,N_4576);
nor U14201 (N_14201,N_9894,N_3937);
nor U14202 (N_14202,N_9792,N_521);
and U14203 (N_14203,N_6836,N_2484);
and U14204 (N_14204,N_8253,N_132);
or U14205 (N_14205,N_4997,N_9495);
nor U14206 (N_14206,N_8362,N_1419);
or U14207 (N_14207,N_2749,N_3145);
and U14208 (N_14208,N_5363,N_1821);
or U14209 (N_14209,N_6790,N_3663);
nor U14210 (N_14210,N_4656,N_562);
nand U14211 (N_14211,N_6462,N_3853);
and U14212 (N_14212,N_2488,N_4507);
and U14213 (N_14213,N_2730,N_7781);
or U14214 (N_14214,N_2665,N_4197);
nor U14215 (N_14215,N_2885,N_1688);
nor U14216 (N_14216,N_3701,N_7131);
and U14217 (N_14217,N_9975,N_8629);
and U14218 (N_14218,N_4491,N_4781);
or U14219 (N_14219,N_6539,N_9770);
or U14220 (N_14220,N_4250,N_7218);
nor U14221 (N_14221,N_8161,N_3387);
or U14222 (N_14222,N_3432,N_1742);
nor U14223 (N_14223,N_3517,N_9497);
nor U14224 (N_14224,N_6027,N_118);
nor U14225 (N_14225,N_4242,N_8083);
and U14226 (N_14226,N_3844,N_8789);
and U14227 (N_14227,N_6338,N_2410);
nor U14228 (N_14228,N_8347,N_2683);
and U14229 (N_14229,N_7913,N_9317);
or U14230 (N_14230,N_1660,N_3267);
nor U14231 (N_14231,N_7247,N_9679);
or U14232 (N_14232,N_7640,N_1841);
nor U14233 (N_14233,N_3952,N_6157);
or U14234 (N_14234,N_5613,N_963);
and U14235 (N_14235,N_1945,N_4359);
nand U14236 (N_14236,N_337,N_3113);
and U14237 (N_14237,N_3824,N_6242);
nor U14238 (N_14238,N_2708,N_9287);
or U14239 (N_14239,N_3854,N_1134);
or U14240 (N_14240,N_5282,N_5780);
nor U14241 (N_14241,N_9809,N_8262);
nor U14242 (N_14242,N_6123,N_9145);
nor U14243 (N_14243,N_3363,N_1727);
and U14244 (N_14244,N_3867,N_1923);
nand U14245 (N_14245,N_7353,N_4477);
or U14246 (N_14246,N_9931,N_2006);
or U14247 (N_14247,N_5233,N_8537);
nor U14248 (N_14248,N_2164,N_2489);
nor U14249 (N_14249,N_6344,N_4043);
or U14250 (N_14250,N_2837,N_6890);
and U14251 (N_14251,N_1604,N_6578);
nor U14252 (N_14252,N_281,N_5353);
nor U14253 (N_14253,N_575,N_5993);
or U14254 (N_14254,N_8907,N_6546);
or U14255 (N_14255,N_8176,N_9195);
nand U14256 (N_14256,N_1150,N_8420);
or U14257 (N_14257,N_355,N_4805);
and U14258 (N_14258,N_6674,N_5165);
nor U14259 (N_14259,N_1271,N_5117);
and U14260 (N_14260,N_7277,N_1825);
or U14261 (N_14261,N_1333,N_5950);
nor U14262 (N_14262,N_1258,N_3886);
and U14263 (N_14263,N_468,N_9845);
or U14264 (N_14264,N_233,N_2767);
and U14265 (N_14265,N_376,N_5762);
nor U14266 (N_14266,N_5999,N_3502);
or U14267 (N_14267,N_4006,N_5960);
nand U14268 (N_14268,N_600,N_5847);
xnor U14269 (N_14269,N_9928,N_135);
or U14270 (N_14270,N_796,N_9599);
nor U14271 (N_14271,N_913,N_142);
nand U14272 (N_14272,N_9578,N_1684);
nor U14273 (N_14273,N_4766,N_8311);
and U14274 (N_14274,N_2319,N_5997);
and U14275 (N_14275,N_9511,N_5386);
nor U14276 (N_14276,N_7590,N_2037);
nand U14277 (N_14277,N_6816,N_956);
nor U14278 (N_14278,N_9384,N_872);
nor U14279 (N_14279,N_5596,N_3162);
and U14280 (N_14280,N_5018,N_486);
or U14281 (N_14281,N_1106,N_570);
and U14282 (N_14282,N_3577,N_8504);
nand U14283 (N_14283,N_1375,N_6305);
nand U14284 (N_14284,N_7064,N_7077);
nand U14285 (N_14285,N_5029,N_7127);
nand U14286 (N_14286,N_8799,N_8589);
nor U14287 (N_14287,N_5150,N_9234);
nor U14288 (N_14288,N_8295,N_6634);
and U14289 (N_14289,N_3971,N_4361);
nor U14290 (N_14290,N_2821,N_799);
or U14291 (N_14291,N_5225,N_3596);
and U14292 (N_14292,N_2644,N_2980);
nand U14293 (N_14293,N_5224,N_9516);
nand U14294 (N_14294,N_8602,N_8760);
and U14295 (N_14295,N_8805,N_5120);
nor U14296 (N_14296,N_3348,N_8915);
nand U14297 (N_14297,N_3057,N_7297);
or U14298 (N_14298,N_2050,N_5655);
nand U14299 (N_14299,N_723,N_4428);
nor U14300 (N_14300,N_146,N_4989);
nand U14301 (N_14301,N_7314,N_406);
nor U14302 (N_14302,N_1328,N_3216);
or U14303 (N_14303,N_8357,N_6273);
nand U14304 (N_14304,N_6250,N_2797);
or U14305 (N_14305,N_2157,N_2426);
and U14306 (N_14306,N_8201,N_9100);
and U14307 (N_14307,N_8813,N_8402);
and U14308 (N_14308,N_8830,N_1785);
nand U14309 (N_14309,N_7410,N_5807);
nor U14310 (N_14310,N_7428,N_8250);
and U14311 (N_14311,N_6703,N_5383);
and U14312 (N_14312,N_7940,N_2224);
or U14313 (N_14313,N_1408,N_3562);
nand U14314 (N_14314,N_1718,N_3710);
nand U14315 (N_14315,N_8247,N_8345);
nor U14316 (N_14316,N_6798,N_3219);
nand U14317 (N_14317,N_9584,N_6627);
or U14318 (N_14318,N_5544,N_5203);
or U14319 (N_14319,N_5942,N_7925);
or U14320 (N_14320,N_9954,N_2010);
xnor U14321 (N_14321,N_6921,N_4841);
xor U14322 (N_14322,N_6476,N_3682);
nor U14323 (N_14323,N_1220,N_3021);
nor U14324 (N_14324,N_6885,N_9389);
or U14325 (N_14325,N_4831,N_2816);
nor U14326 (N_14326,N_725,N_6388);
nand U14327 (N_14327,N_3178,N_7161);
nor U14328 (N_14328,N_9488,N_9534);
and U14329 (N_14329,N_5209,N_8588);
nand U14330 (N_14330,N_9333,N_5732);
nand U14331 (N_14331,N_2545,N_80);
and U14332 (N_14332,N_402,N_9083);
nor U14333 (N_14333,N_9273,N_547);
and U14334 (N_14334,N_8494,N_8634);
and U14335 (N_14335,N_4695,N_6839);
nand U14336 (N_14336,N_6598,N_9855);
nand U14337 (N_14337,N_2662,N_4327);
nand U14338 (N_14338,N_7518,N_9441);
or U14339 (N_14339,N_4758,N_5261);
or U14340 (N_14340,N_1635,N_1324);
nand U14341 (N_14341,N_2820,N_2);
and U14342 (N_14342,N_6821,N_9104);
nor U14343 (N_14343,N_9628,N_3300);
nor U14344 (N_14344,N_1792,N_1115);
and U14345 (N_14345,N_9307,N_1901);
nand U14346 (N_14346,N_2567,N_6727);
and U14347 (N_14347,N_8269,N_1236);
nand U14348 (N_14348,N_7647,N_8604);
or U14349 (N_14349,N_9728,N_8426);
and U14350 (N_14350,N_9048,N_7167);
nor U14351 (N_14351,N_1940,N_4143);
or U14352 (N_14352,N_9005,N_1132);
nor U14353 (N_14353,N_8579,N_8655);
or U14354 (N_14354,N_5559,N_1005);
and U14355 (N_14355,N_9021,N_1715);
nand U14356 (N_14356,N_4647,N_5663);
and U14357 (N_14357,N_787,N_2161);
and U14358 (N_14358,N_5719,N_6489);
nor U14359 (N_14359,N_5966,N_1868);
nand U14360 (N_14360,N_9446,N_958);
and U14361 (N_14361,N_5438,N_4808);
nor U14362 (N_14362,N_4884,N_4012);
nand U14363 (N_14363,N_4333,N_398);
or U14364 (N_14364,N_3285,N_9876);
and U14365 (N_14365,N_374,N_6042);
and U14366 (N_14366,N_6604,N_5361);
and U14367 (N_14367,N_8703,N_6672);
and U14368 (N_14368,N_441,N_694);
nand U14369 (N_14369,N_5424,N_3820);
nor U14370 (N_14370,N_2016,N_1870);
or U14371 (N_14371,N_2628,N_8738);
nor U14372 (N_14372,N_5865,N_1229);
or U14373 (N_14373,N_6926,N_1368);
nand U14374 (N_14374,N_1263,N_9437);
nand U14375 (N_14375,N_3530,N_176);
nand U14376 (N_14376,N_1711,N_5858);
nor U14377 (N_14377,N_4178,N_8976);
and U14378 (N_14378,N_9962,N_1117);
and U14379 (N_14379,N_8463,N_3690);
nor U14380 (N_14380,N_35,N_2055);
nor U14381 (N_14381,N_2974,N_9747);
nand U14382 (N_14382,N_5826,N_5467);
nor U14383 (N_14383,N_121,N_9279);
and U14384 (N_14384,N_1342,N_4300);
nand U14385 (N_14385,N_625,N_1551);
and U14386 (N_14386,N_1934,N_63);
nor U14387 (N_14387,N_9374,N_5924);
nand U14388 (N_14388,N_5285,N_9961);
and U14389 (N_14389,N_6100,N_6661);
and U14390 (N_14390,N_197,N_802);
and U14391 (N_14391,N_8113,N_6040);
nor U14392 (N_14392,N_2432,N_460);
nand U14393 (N_14393,N_7681,N_9245);
and U14394 (N_14394,N_8439,N_3138);
nand U14395 (N_14395,N_4911,N_8828);
and U14396 (N_14396,N_6719,N_7142);
and U14397 (N_14397,N_5673,N_4959);
nor U14398 (N_14398,N_1112,N_3597);
or U14399 (N_14399,N_7426,N_5009);
or U14400 (N_14400,N_5529,N_9793);
and U14401 (N_14401,N_8486,N_6855);
or U14402 (N_14402,N_515,N_5023);
and U14403 (N_14403,N_1566,N_3676);
nand U14404 (N_14404,N_2434,N_7338);
nor U14405 (N_14405,N_3586,N_8392);
and U14406 (N_14406,N_8074,N_2260);
nand U14407 (N_14407,N_1286,N_7178);
nand U14408 (N_14408,N_3413,N_6758);
nand U14409 (N_14409,N_7159,N_3811);
nor U14410 (N_14410,N_914,N_6240);
nor U14411 (N_14411,N_5106,N_5217);
and U14412 (N_14412,N_9949,N_3029);
and U14413 (N_14413,N_8930,N_7783);
and U14414 (N_14414,N_6889,N_3802);
and U14415 (N_14415,N_8582,N_5296);
or U14416 (N_14416,N_2555,N_7624);
nor U14417 (N_14417,N_573,N_4806);
nand U14418 (N_14418,N_9467,N_1528);
nand U14419 (N_14419,N_2115,N_4039);
nor U14420 (N_14420,N_81,N_9184);
or U14421 (N_14421,N_7740,N_5915);
nor U14422 (N_14422,N_484,N_1714);
nor U14423 (N_14423,N_4190,N_1472);
or U14424 (N_14424,N_7396,N_2244);
nand U14425 (N_14425,N_6518,N_4391);
nor U14426 (N_14426,N_8363,N_5274);
nor U14427 (N_14427,N_8480,N_4422);
or U14428 (N_14428,N_5047,N_7066);
or U14429 (N_14429,N_569,N_2054);
and U14430 (N_14430,N_7321,N_2995);
or U14431 (N_14431,N_4587,N_8476);
nand U14432 (N_14432,N_2413,N_9159);
and U14433 (N_14433,N_6630,N_3217);
or U14434 (N_14434,N_2579,N_9223);
or U14435 (N_14435,N_6831,N_9196);
and U14436 (N_14436,N_3409,N_5640);
nor U14437 (N_14437,N_2850,N_2149);
nor U14438 (N_14438,N_1289,N_1738);
nand U14439 (N_14439,N_1591,N_1077);
and U14440 (N_14440,N_4438,N_9105);
nor U14441 (N_14441,N_7971,N_2876);
and U14442 (N_14442,N_9473,N_209);
or U14443 (N_14443,N_2512,N_654);
and U14444 (N_14444,N_8834,N_44);
nand U14445 (N_14445,N_7729,N_3064);
or U14446 (N_14446,N_8505,N_1559);
nor U14447 (N_14447,N_9243,N_4170);
nor U14448 (N_14448,N_3455,N_4280);
nand U14449 (N_14449,N_4434,N_9342);
nor U14450 (N_14450,N_3668,N_6544);
or U14451 (N_14451,N_5385,N_421);
or U14452 (N_14452,N_7405,N_8005);
nor U14453 (N_14453,N_131,N_2751);
or U14454 (N_14454,N_8642,N_2440);
nand U14455 (N_14455,N_3765,N_7787);
or U14456 (N_14456,N_2627,N_7948);
or U14457 (N_14457,N_9804,N_148);
and U14458 (N_14458,N_9006,N_1891);
nand U14459 (N_14459,N_169,N_5258);
nor U14460 (N_14460,N_9705,N_2257);
nand U14461 (N_14461,N_3636,N_3883);
or U14462 (N_14462,N_481,N_5617);
and U14463 (N_14463,N_6779,N_3878);
and U14464 (N_14464,N_1845,N_1264);
nand U14465 (N_14465,N_389,N_2179);
nor U14466 (N_14466,N_7886,N_199);
xor U14467 (N_14467,N_1884,N_6149);
or U14468 (N_14468,N_4150,N_4602);
or U14469 (N_14469,N_7763,N_3375);
or U14470 (N_14470,N_9813,N_9423);
nand U14471 (N_14471,N_1491,N_9271);
nand U14472 (N_14472,N_3141,N_8633);
nand U14473 (N_14473,N_6308,N_7659);
or U14474 (N_14474,N_5767,N_6714);
or U14475 (N_14475,N_4115,N_9080);
and U14476 (N_14476,N_5558,N_3508);
or U14477 (N_14477,N_377,N_9203);
and U14478 (N_14478,N_2060,N_922);
and U14479 (N_14479,N_4598,N_9054);
and U14480 (N_14480,N_5646,N_2111);
and U14481 (N_14481,N_3385,N_5368);
or U14482 (N_14482,N_9939,N_5522);
xor U14483 (N_14483,N_4484,N_2387);
nor U14484 (N_14484,N_9343,N_7030);
nand U14485 (N_14485,N_5195,N_2225);
nand U14486 (N_14486,N_1326,N_5351);
and U14487 (N_14487,N_4270,N_9867);
nor U14488 (N_14488,N_9781,N_3415);
nor U14489 (N_14489,N_6557,N_523);
or U14490 (N_14490,N_9477,N_5300);
or U14491 (N_14491,N_1349,N_1382);
nor U14492 (N_14492,N_9824,N_2865);
and U14493 (N_14493,N_4607,N_3148);
and U14494 (N_14494,N_7810,N_4741);
or U14495 (N_14495,N_9742,N_5163);
xnor U14496 (N_14496,N_7129,N_8326);
or U14497 (N_14497,N_6220,N_1709);
and U14498 (N_14498,N_6311,N_5742);
nand U14499 (N_14499,N_267,N_1245);
and U14500 (N_14500,N_9683,N_6142);
nor U14501 (N_14501,N_8123,N_598);
nand U14502 (N_14502,N_5879,N_8521);
nand U14503 (N_14503,N_4830,N_474);
nand U14504 (N_14504,N_6190,N_330);
and U14505 (N_14505,N_9320,N_8993);
nand U14506 (N_14506,N_5155,N_3842);
nor U14507 (N_14507,N_3600,N_6372);
nor U14508 (N_14508,N_2277,N_2963);
and U14509 (N_14509,N_8689,N_1527);
or U14510 (N_14510,N_9725,N_2649);
nor U14511 (N_14511,N_508,N_7046);
nor U14512 (N_14512,N_2574,N_9574);
or U14513 (N_14513,N_3404,N_8212);
nor U14514 (N_14514,N_4189,N_2036);
nand U14515 (N_14515,N_1171,N_8682);
nor U14516 (N_14516,N_3319,N_5244);
nor U14517 (N_14517,N_1450,N_5417);
or U14518 (N_14518,N_9365,N_6059);
nor U14519 (N_14519,N_8204,N_7979);
and U14520 (N_14520,N_8797,N_189);
or U14521 (N_14521,N_4072,N_6769);
or U14522 (N_14522,N_2505,N_4735);
nor U14523 (N_14523,N_152,N_2103);
nand U14524 (N_14524,N_4692,N_6060);
nand U14525 (N_14525,N_7702,N_3914);
or U14526 (N_14526,N_5765,N_7489);
or U14527 (N_14527,N_1866,N_2282);
xnor U14528 (N_14528,N_4119,N_8524);
or U14529 (N_14529,N_1706,N_6679);
and U14530 (N_14530,N_5138,N_8255);
or U14531 (N_14531,N_52,N_1174);
nand U14532 (N_14532,N_7719,N_3719);
nor U14533 (N_14533,N_9009,N_6730);
or U14534 (N_14534,N_6275,N_5182);
or U14535 (N_14535,N_6850,N_7516);
and U14536 (N_14536,N_3378,N_9930);
or U14537 (N_14537,N_6766,N_7192);
and U14538 (N_14538,N_7631,N_8343);
or U14539 (N_14539,N_3637,N_5783);
nand U14540 (N_14540,N_4599,N_6169);
nor U14541 (N_14541,N_2132,N_3659);
and U14542 (N_14542,N_4034,N_2423);
and U14543 (N_14543,N_2654,N_7452);
or U14544 (N_14544,N_5425,N_7471);
and U14545 (N_14545,N_9165,N_8568);
and U14546 (N_14546,N_6288,N_4628);
nand U14547 (N_14547,N_5945,N_9124);
and U14548 (N_14548,N_4746,N_3120);
or U14549 (N_14549,N_1441,N_6708);
or U14550 (N_14550,N_6477,N_4304);
and U14551 (N_14551,N_4266,N_1516);
nor U14552 (N_14552,N_1921,N_5978);
nand U14553 (N_14553,N_4065,N_1037);
or U14554 (N_14554,N_7824,N_3830);
nand U14555 (N_14555,N_8358,N_5668);
nor U14556 (N_14556,N_4478,N_7717);
and U14557 (N_14557,N_6228,N_4386);
nand U14558 (N_14558,N_2631,N_3024);
and U14559 (N_14559,N_9946,N_9409);
nor U14560 (N_14560,N_7643,N_1205);
or U14561 (N_14561,N_9202,N_2127);
nand U14562 (N_14562,N_7714,N_3560);
and U14563 (N_14563,N_6841,N_126);
and U14564 (N_14564,N_8618,N_2470);
and U14565 (N_14565,N_4460,N_2959);
and U14566 (N_14566,N_362,N_9087);
nor U14567 (N_14567,N_5369,N_2135);
nor U14568 (N_14568,N_9673,N_3622);
and U14569 (N_14569,N_11,N_9484);
nor U14570 (N_14570,N_127,N_1700);
nand U14571 (N_14571,N_5092,N_6654);
nor U14572 (N_14572,N_5969,N_4912);
nor U14573 (N_14573,N_7267,N_4639);
nand U14574 (N_14574,N_7014,N_8499);
nand U14575 (N_14575,N_7320,N_4779);
and U14576 (N_14576,N_8839,N_2989);
and U14577 (N_14577,N_1490,N_8944);
or U14578 (N_14578,N_4229,N_7038);
nand U14579 (N_14579,N_1672,N_1343);
nor U14580 (N_14580,N_1101,N_393);
or U14581 (N_14581,N_6996,N_4616);
nor U14582 (N_14582,N_7122,N_5809);
or U14583 (N_14583,N_2720,N_8441);
and U14584 (N_14584,N_9193,N_4255);
nand U14585 (N_14585,N_26,N_1255);
and U14586 (N_14586,N_1933,N_3822);
and U14587 (N_14587,N_304,N_6062);
or U14588 (N_14588,N_5700,N_7715);
or U14589 (N_14589,N_9399,N_3371);
nand U14590 (N_14590,N_316,N_1704);
nand U14591 (N_14591,N_3976,N_8388);
nand U14592 (N_14592,N_4926,N_8407);
nand U14593 (N_14593,N_7292,N_3126);
or U14594 (N_14594,N_3587,N_1166);
nand U14595 (N_14595,N_5883,N_8164);
nor U14596 (N_14596,N_6915,N_2233);
or U14597 (N_14597,N_6431,N_5725);
nor U14598 (N_14598,N_9065,N_9089);
nand U14599 (N_14599,N_3295,N_1301);
nand U14600 (N_14600,N_5840,N_7380);
or U14601 (N_14601,N_6685,N_3298);
nor U14602 (N_14602,N_4539,N_8780);
nand U14603 (N_14603,N_6459,N_8288);
nand U14604 (N_14604,N_4239,N_8350);
nor U14605 (N_14605,N_1661,N_5638);
nand U14606 (N_14606,N_27,N_3859);
nand U14607 (N_14607,N_4612,N_4740);
nand U14608 (N_14608,N_476,N_168);
or U14609 (N_14609,N_2312,N_4791);
nor U14610 (N_14610,N_2591,N_7498);
or U14611 (N_14611,N_8874,N_7326);
or U14612 (N_14612,N_8989,N_3903);
nand U14613 (N_14613,N_5216,N_4980);
and U14614 (N_14614,N_8267,N_7304);
nor U14615 (N_14615,N_3443,N_133);
or U14616 (N_14616,N_8939,N_8843);
and U14617 (N_14617,N_9908,N_1633);
and U14618 (N_14618,N_4231,N_4049);
nor U14619 (N_14619,N_6353,N_3940);
nor U14620 (N_14620,N_7859,N_4787);
and U14621 (N_14621,N_6080,N_1170);
xnor U14622 (N_14622,N_4358,N_3503);
or U14623 (N_14623,N_8467,N_5560);
nor U14624 (N_14624,N_5530,N_134);
nor U14625 (N_14625,N_1095,N_3027);
xor U14626 (N_14626,N_7069,N_6666);
nor U14627 (N_14627,N_8207,N_452);
nand U14628 (N_14628,N_2394,N_3840);
nand U14629 (N_14629,N_4446,N_9650);
nand U14630 (N_14630,N_5032,N_3879);
and U14631 (N_14631,N_4317,N_4184);
or U14632 (N_14632,N_7543,N_285);
or U14633 (N_14633,N_9073,N_9319);
nand U14634 (N_14634,N_6134,N_6197);
and U14635 (N_14635,N_4809,N_1732);
nor U14636 (N_14636,N_7667,N_437);
nand U14637 (N_14637,N_4306,N_1049);
or U14638 (N_14638,N_908,N_4752);
and U14639 (N_14639,N_834,N_8709);
nor U14640 (N_14640,N_8208,N_3692);
nor U14641 (N_14641,N_5088,N_9059);
nand U14642 (N_14642,N_7844,N_8519);
nand U14643 (N_14643,N_2185,N_4707);
nor U14644 (N_14644,N_8646,N_6587);
nand U14645 (N_14645,N_1911,N_2893);
nor U14646 (N_14646,N_9079,N_7574);
and U14647 (N_14647,N_4321,N_4492);
or U14648 (N_14648,N_6689,N_3929);
nor U14649 (N_14649,N_2494,N_8909);
or U14650 (N_14650,N_361,N_175);
and U14651 (N_14651,N_7097,N_3149);
nand U14652 (N_14652,N_5766,N_3558);
or U14653 (N_14653,N_6033,N_4374);
and U14654 (N_14654,N_2583,N_3753);
nor U14655 (N_14655,N_822,N_3938);
nor U14656 (N_14656,N_3201,N_640);
nand U14657 (N_14657,N_7672,N_5319);
nor U14658 (N_14658,N_8106,N_5169);
nand U14659 (N_14659,N_7239,N_8816);
nor U14660 (N_14660,N_8540,N_5326);
and U14661 (N_14661,N_5775,N_2026);
or U14662 (N_14662,N_5548,N_3985);
nand U14663 (N_14663,N_1659,N_2436);
nor U14664 (N_14664,N_5196,N_2704);
or U14665 (N_14665,N_1947,N_805);
nand U14666 (N_14666,N_9189,N_71);
nand U14667 (N_14667,N_6436,N_9646);
nand U14668 (N_14668,N_9191,N_9772);
or U14669 (N_14669,N_6295,N_147);
and U14670 (N_14670,N_427,N_5713);
and U14671 (N_14671,N_2136,N_2779);
and U14672 (N_14672,N_3629,N_8218);
nor U14673 (N_14673,N_5202,N_9636);
and U14674 (N_14674,N_669,N_7833);
or U14675 (N_14675,N_8313,N_9709);
nand U14676 (N_14676,N_5898,N_400);
and U14677 (N_14677,N_5650,N_250);
nand U14678 (N_14678,N_401,N_9324);
or U14679 (N_14679,N_6017,N_7716);
nand U14680 (N_14680,N_5964,N_5342);
nand U14681 (N_14681,N_5975,N_9028);
nor U14682 (N_14682,N_2411,N_8687);
nor U14683 (N_14683,N_9660,N_7622);
or U14684 (N_14684,N_7089,N_2884);
nand U14685 (N_14685,N_7189,N_6541);
nand U14686 (N_14686,N_3996,N_9575);
nor U14687 (N_14687,N_4882,N_257);
or U14688 (N_14688,N_4952,N_4802);
or U14689 (N_14689,N_6750,N_7073);
nor U14690 (N_14690,N_2907,N_3161);
nand U14691 (N_14691,N_5246,N_5409);
nor U14692 (N_14692,N_8009,N_2951);
or U14693 (N_14693,N_2306,N_3273);
and U14694 (N_14694,N_2696,N_1036);
nor U14695 (N_14695,N_6965,N_2124);
nor U14696 (N_14696,N_9727,N_6202);
or U14697 (N_14697,N_3832,N_4000);
nand U14698 (N_14698,N_8798,N_4047);
and U14699 (N_14699,N_8790,N_6819);
nand U14700 (N_14700,N_5864,N_1272);
nor U14701 (N_14701,N_7534,N_7121);
and U14702 (N_14702,N_7171,N_6373);
and U14703 (N_14703,N_4036,N_3720);
or U14704 (N_14704,N_3693,N_804);
or U14705 (N_14705,N_1654,N_4535);
nand U14706 (N_14706,N_5664,N_2308);
nor U14707 (N_14707,N_4890,N_3224);
nand U14708 (N_14708,N_8408,N_4017);
nor U14709 (N_14709,N_1332,N_9887);
and U14710 (N_14710,N_283,N_7413);
or U14711 (N_14711,N_4518,N_8954);
nand U14712 (N_14712,N_2119,N_558);
nor U14713 (N_14713,N_181,N_5164);
nor U14714 (N_14714,N_1501,N_9886);
nor U14715 (N_14715,N_8140,N_513);
and U14716 (N_14716,N_4941,N_4083);
and U14717 (N_14717,N_8011,N_1987);
nand U14718 (N_14718,N_2770,N_6265);
nor U14719 (N_14719,N_5136,N_554);
nor U14720 (N_14720,N_6954,N_4257);
nor U14721 (N_14721,N_1858,N_3305);
nor U14722 (N_14722,N_394,N_2034);
and U14723 (N_14723,N_438,N_5127);
or U14724 (N_14724,N_7838,N_7182);
and U14725 (N_14725,N_2023,N_7376);
nor U14726 (N_14726,N_8783,N_9211);
nand U14727 (N_14727,N_6562,N_7107);
nor U14728 (N_14728,N_7168,N_4114);
or U14729 (N_14729,N_5580,N_3366);
nand U14730 (N_14730,N_3804,N_2442);
nor U14731 (N_14731,N_8008,N_4415);
or U14732 (N_14732,N_7827,N_8605);
and U14733 (N_14733,N_8265,N_7569);
or U14734 (N_14734,N_2433,N_4958);
and U14735 (N_14735,N_8781,N_2961);
nor U14736 (N_14736,N_5298,N_9969);
or U14737 (N_14737,N_2462,N_5205);
nand U14738 (N_14738,N_8468,N_1183);
nand U14739 (N_14739,N_4728,N_9750);
nor U14740 (N_14740,N_8538,N_1474);
xnor U14741 (N_14741,N_2063,N_1488);
nor U14742 (N_14742,N_5962,N_8158);
nor U14743 (N_14743,N_3211,N_9936);
nand U14744 (N_14744,N_1536,N_5618);
and U14745 (N_14745,N_6118,N_2766);
nor U14746 (N_14746,N_4413,N_4864);
or U14747 (N_14747,N_2287,N_8693);
or U14748 (N_14748,N_9227,N_2358);
and U14749 (N_14749,N_4693,N_9797);
or U14750 (N_14750,N_32,N_2344);
or U14751 (N_14751,N_507,N_3086);
nand U14752 (N_14752,N_2912,N_9877);
or U14753 (N_14753,N_4310,N_9531);
nor U14754 (N_14754,N_3177,N_6542);
nor U14755 (N_14755,N_7798,N_8254);
nor U14756 (N_14756,N_9987,N_7841);
nand U14757 (N_14757,N_9547,N_1337);
nand U14758 (N_14758,N_1219,N_2782);
or U14759 (N_14759,N_2859,N_2640);
and U14760 (N_14760,N_9256,N_939);
xor U14761 (N_14761,N_1378,N_7987);
or U14762 (N_14762,N_1563,N_8942);
and U14763 (N_14763,N_352,N_5102);
and U14764 (N_14764,N_2336,N_2867);
or U14765 (N_14765,N_5716,N_8175);
nor U14766 (N_14766,N_4051,N_4287);
nor U14767 (N_14767,N_4873,N_9001);
or U14768 (N_14768,N_4480,N_3143);
nand U14769 (N_14769,N_8665,N_6107);
nor U14770 (N_14770,N_7544,N_729);
and U14771 (N_14771,N_8549,N_5496);
or U14772 (N_14772,N_7088,N_9138);
or U14773 (N_14773,N_534,N_252);
nand U14774 (N_14774,N_6432,N_2838);
nand U14775 (N_14775,N_4510,N_7683);
or U14776 (N_14776,N_4442,N_8794);
nand U14777 (N_14777,N_9799,N_689);
nor U14778 (N_14778,N_5977,N_9743);
or U14779 (N_14779,N_8355,N_7572);
nor U14780 (N_14780,N_676,N_5273);
nand U14781 (N_14781,N_8614,N_3747);
or U14782 (N_14782,N_3864,N_4459);
nand U14783 (N_14783,N_163,N_5553);
nand U14784 (N_14784,N_6260,N_2219);
nand U14785 (N_14785,N_975,N_8448);
or U14786 (N_14786,N_1733,N_6375);
nand U14787 (N_14787,N_7822,N_9302);
or U14788 (N_14788,N_2170,N_1735);
nand U14789 (N_14789,N_386,N_9308);
nor U14790 (N_14790,N_4807,N_144);
xnor U14791 (N_14791,N_1662,N_2242);
and U14792 (N_14792,N_7,N_1560);
and U14793 (N_14793,N_8352,N_3946);
or U14794 (N_14794,N_3548,N_3076);
nor U14795 (N_14795,N_928,N_2602);
xor U14796 (N_14796,N_4038,N_6706);
and U14797 (N_14797,N_1135,N_8281);
or U14798 (N_14798,N_7731,N_701);
and U14799 (N_14799,N_2072,N_2992);
or U14800 (N_14800,N_9978,N_4220);
and U14801 (N_14801,N_9840,N_9927);
nor U14802 (N_14802,N_8462,N_4979);
or U14803 (N_14803,N_1997,N_5738);
or U14804 (N_14804,N_2634,N_8327);
or U14805 (N_14805,N_6195,N_8532);
or U14806 (N_14806,N_6493,N_851);
nand U14807 (N_14807,N_1276,N_3435);
and U14808 (N_14808,N_1963,N_3821);
and U14809 (N_14809,N_9883,N_6235);
and U14810 (N_14810,N_5151,N_4275);
nand U14811 (N_14811,N_6154,N_2614);
and U14812 (N_14812,N_5148,N_4277);
and U14813 (N_14813,N_3611,N_6668);
nor U14814 (N_14814,N_2625,N_8927);
nand U14815 (N_14815,N_9160,N_2542);
nor U14816 (N_14816,N_703,N_3252);
nand U14817 (N_14817,N_9579,N_9935);
nand U14818 (N_14818,N_3500,N_4218);
nand U14819 (N_14819,N_3808,N_8947);
nand U14820 (N_14820,N_42,N_1184);
and U14821 (N_14821,N_6097,N_8298);
or U14822 (N_14822,N_9640,N_2342);
and U14823 (N_14823,N_3204,N_5498);
nand U14824 (N_14824,N_6138,N_3368);
nand U14825 (N_14825,N_3244,N_408);
nor U14826 (N_14826,N_2673,N_9625);
or U14827 (N_14827,N_6532,N_4684);
nor U14828 (N_14828,N_4061,N_1630);
nand U14829 (N_14829,N_5570,N_9294);
nand U14830 (N_14830,N_773,N_6606);
or U14831 (N_14831,N_4933,N_3795);
and U14832 (N_14832,N_7424,N_3605);
and U14833 (N_14833,N_5748,N_7398);
or U14834 (N_14834,N_5218,N_7488);
nand U14835 (N_14835,N_9366,N_655);
and U14836 (N_14836,N_9988,N_9031);
nor U14837 (N_14837,N_5211,N_6746);
or U14838 (N_14838,N_6653,N_4685);
nand U14839 (N_14839,N_1226,N_8962);
or U14840 (N_14840,N_6500,N_6611);
nand U14841 (N_14841,N_6164,N_380);
nand U14842 (N_14842,N_2373,N_8251);
and U14843 (N_14843,N_6826,N_8380);
and U14844 (N_14844,N_8696,N_4007);
and U14845 (N_14845,N_9947,N_7386);
nor U14846 (N_14846,N_3604,N_6394);
and U14847 (N_14847,N_2096,N_1980);
and U14848 (N_14848,N_3266,N_8595);
and U14849 (N_14849,N_7253,N_3279);
xor U14850 (N_14850,N_3786,N_9093);
nor U14851 (N_14851,N_8275,N_1075);
or U14852 (N_14852,N_954,N_5131);
or U14853 (N_14853,N_8376,N_5979);
nor U14854 (N_14854,N_9794,N_9585);
nor U14855 (N_14855,N_5627,N_5730);
nand U14856 (N_14856,N_4573,N_7941);
nand U14857 (N_14857,N_5034,N_179);
or U14858 (N_14858,N_9231,N_6637);
nor U14859 (N_14859,N_7563,N_6896);
nand U14860 (N_14860,N_7559,N_6318);
nor U14861 (N_14861,N_1471,N_2814);
nand U14862 (N_14862,N_9948,N_1628);
nand U14863 (N_14863,N_4969,N_5786);
or U14864 (N_14864,N_1111,N_8625);
and U14865 (N_14865,N_7158,N_6119);
nand U14866 (N_14866,N_8052,N_5133);
and U14867 (N_14867,N_7938,N_5143);
or U14868 (N_14868,N_4558,N_9255);
and U14869 (N_14869,N_1162,N_6759);
nor U14870 (N_14870,N_459,N_7233);
or U14871 (N_14871,N_5230,N_8940);
nor U14872 (N_14872,N_340,N_3687);
and U14873 (N_14873,N_8516,N_4052);
nand U14874 (N_14874,N_3975,N_3917);
nor U14875 (N_14875,N_8213,N_1487);
and U14876 (N_14876,N_1687,N_8777);
or U14877 (N_14877,N_7117,N_1561);
nand U14878 (N_14878,N_9712,N_3354);
nor U14879 (N_14879,N_6371,N_5402);
nor U14880 (N_14880,N_8215,N_9183);
and U14881 (N_14881,N_6575,N_1188);
and U14882 (N_14882,N_2272,N_5493);
nand U14883 (N_14883,N_674,N_9737);
nor U14884 (N_14884,N_4094,N_3475);
or U14885 (N_14885,N_2341,N_9198);
and U14886 (N_14886,N_2478,N_3666);
and U14887 (N_14887,N_7497,N_7323);
nor U14888 (N_14888,N_8526,N_5347);
xnor U14889 (N_14889,N_6444,N_5698);
nor U14890 (N_14890,N_7513,N_1766);
or U14891 (N_14891,N_7016,N_4542);
nand U14892 (N_14892,N_690,N_9219);
nor U14893 (N_14893,N_7281,N_9244);
and U14894 (N_14894,N_4351,N_9810);
and U14895 (N_14895,N_1439,N_5229);
xor U14896 (N_14896,N_18,N_6886);
nand U14897 (N_14897,N_1089,N_1803);
or U14898 (N_14898,N_2969,N_7390);
and U14899 (N_14899,N_5327,N_545);
nand U14900 (N_14900,N_8145,N_6043);
nand U14901 (N_14901,N_6897,N_2150);
or U14902 (N_14902,N_2616,N_2679);
and U14903 (N_14903,N_4891,N_2744);
nor U14904 (N_14904,N_6179,N_2002);
nand U14905 (N_14905,N_1703,N_7065);
or U14906 (N_14906,N_9178,N_1648);
nand U14907 (N_14907,N_3082,N_5649);
nor U14908 (N_14908,N_9993,N_9716);
or U14909 (N_14909,N_4390,N_6640);
or U14910 (N_14910,N_2652,N_2367);
or U14911 (N_14911,N_4924,N_5252);
and U14912 (N_14912,N_8647,N_6297);
nand U14913 (N_14913,N_7473,N_5532);
nand U14914 (N_14914,N_7429,N_5157);
and U14915 (N_14915,N_7204,N_87);
or U14916 (N_14916,N_3856,N_5856);
or U14917 (N_14917,N_2447,N_5632);
nand U14918 (N_14918,N_6507,N_6579);
nand U14919 (N_14919,N_3742,N_5346);
nor U14920 (N_14920,N_2215,N_4919);
nor U14921 (N_14921,N_1122,N_7305);
or U14922 (N_14922,N_3391,N_2251);
or U14923 (N_14923,N_3343,N_5419);
nor U14924 (N_14924,N_5413,N_7705);
nor U14925 (N_14925,N_7082,N_7109);
nor U14926 (N_14926,N_6985,N_6794);
or U14927 (N_14927,N_2316,N_2716);
and U14928 (N_14928,N_1839,N_8753);
nor U14929 (N_14929,N_1954,N_5721);
nand U14930 (N_14930,N_3608,N_3072);
nor U14931 (N_14931,N_7458,N_8598);
or U14932 (N_14932,N_6167,N_3407);
nand U14933 (N_14933,N_5519,N_5376);
and U14934 (N_14934,N_6945,N_8157);
nor U14935 (N_14935,N_8918,N_9269);
nor U14936 (N_14936,N_4254,N_7494);
nor U14937 (N_14937,N_4570,N_7185);
or U14938 (N_14938,N_962,N_5003);
or U14939 (N_14939,N_9592,N_5181);
nor U14940 (N_14940,N_3706,N_6700);
nor U14941 (N_14941,N_5280,N_5159);
nand U14942 (N_14942,N_8837,N_207);
and U14943 (N_14943,N_5799,N_6057);
and U14944 (N_14944,N_9337,N_8026);
nand U14945 (N_14945,N_8334,N_4179);
nand U14946 (N_14946,N_8104,N_5186);
and U14947 (N_14947,N_4226,N_4577);
nand U14948 (N_14948,N_1867,N_5932);
or U14949 (N_14949,N_6478,N_7632);
nand U14950 (N_14950,N_464,N_3389);
nand U14951 (N_14951,N_1348,N_4091);
nand U14952 (N_14952,N_4586,N_7873);
xor U14953 (N_14953,N_2887,N_9475);
nand U14954 (N_14954,N_2259,N_1806);
nand U14955 (N_14955,N_190,N_5093);
nand U14956 (N_14956,N_3981,N_3188);
or U14957 (N_14957,N_5354,N_5526);
nor U14958 (N_14958,N_37,N_745);
or U14959 (N_14959,N_5958,N_3286);
nor U14960 (N_14960,N_9171,N_5973);
and U14961 (N_14961,N_5566,N_3246);
nand U14962 (N_14962,N_4337,N_5615);
or U14963 (N_14963,N_3168,N_7901);
and U14964 (N_14964,N_1065,N_1097);
or U14965 (N_14965,N_2463,N_9361);
or U14966 (N_14966,N_9112,N_5867);
nand U14967 (N_14967,N_9849,N_1424);
or U14968 (N_14968,N_4347,N_4664);
and U14969 (N_14969,N_9042,N_1314);
or U14970 (N_14970,N_246,N_5758);
or U14971 (N_14971,N_9863,N_2655);
or U14972 (N_14972,N_39,N_8719);
nor U14973 (N_14973,N_3398,N_6523);
nand U14974 (N_14974,N_2405,N_6094);
nor U14975 (N_14975,N_3583,N_8367);
nor U14976 (N_14976,N_8725,N_7057);
nand U14977 (N_14977,N_613,N_9417);
nand U14978 (N_14978,N_4865,N_344);
or U14979 (N_14979,N_9247,N_8071);
nand U14980 (N_14980,N_3954,N_9999);
nand U14981 (N_14981,N_2711,N_5897);
and U14982 (N_14982,N_3243,N_2347);
nand U14983 (N_14983,N_2174,N_8727);
nand U14984 (N_14984,N_8351,N_4694);
nor U14985 (N_14985,N_4895,N_1175);
nand U14986 (N_14986,N_5988,N_7017);
nand U14987 (N_14987,N_2291,N_2753);
or U14988 (N_14988,N_2013,N_5471);
nor U14989 (N_14989,N_2035,N_8095);
or U14990 (N_14990,N_4594,N_3420);
nand U14991 (N_14991,N_8335,N_9110);
and U14992 (N_14992,N_8891,N_1266);
nand U14993 (N_14993,N_6,N_2299);
nor U14994 (N_14994,N_8852,N_4944);
nor U14995 (N_14995,N_665,N_307);
or U14996 (N_14996,N_3310,N_905);
or U14997 (N_14997,N_6777,N_4943);
or U14998 (N_14998,N_6129,N_2781);
nand U14999 (N_14999,N_5074,N_2877);
and U15000 (N_15000,N_2595,N_9472);
or U15001 (N_15001,N_3642,N_524);
nor U15002 (N_15002,N_7962,N_2283);
and U15003 (N_15003,N_8990,N_1746);
and U15004 (N_15004,N_4786,N_9062);
or U15005 (N_15005,N_4953,N_1189);
nor U15006 (N_15006,N_3106,N_7326);
nor U15007 (N_15007,N_5633,N_1808);
nor U15008 (N_15008,N_5230,N_1254);
nand U15009 (N_15009,N_1200,N_7829);
and U15010 (N_15010,N_7640,N_8840);
or U15011 (N_15011,N_3281,N_2686);
and U15012 (N_15012,N_8274,N_8470);
nand U15013 (N_15013,N_6550,N_8429);
nor U15014 (N_15014,N_5110,N_2803);
or U15015 (N_15015,N_1667,N_9107);
and U15016 (N_15016,N_835,N_6065);
nor U15017 (N_15017,N_9432,N_3812);
or U15018 (N_15018,N_36,N_6179);
and U15019 (N_15019,N_1068,N_1563);
or U15020 (N_15020,N_4528,N_8533);
nor U15021 (N_15021,N_3918,N_4730);
and U15022 (N_15022,N_4,N_6547);
nand U15023 (N_15023,N_8447,N_9863);
and U15024 (N_15024,N_8134,N_2299);
or U15025 (N_15025,N_5120,N_4408);
nor U15026 (N_15026,N_7823,N_1097);
and U15027 (N_15027,N_2550,N_1107);
nand U15028 (N_15028,N_3302,N_943);
nor U15029 (N_15029,N_3363,N_7018);
nand U15030 (N_15030,N_5709,N_9535);
nand U15031 (N_15031,N_8616,N_5523);
or U15032 (N_15032,N_6013,N_9128);
nor U15033 (N_15033,N_6330,N_6615);
nand U15034 (N_15034,N_5874,N_3732);
nor U15035 (N_15035,N_2571,N_1073);
and U15036 (N_15036,N_4525,N_1799);
or U15037 (N_15037,N_6229,N_3134);
or U15038 (N_15038,N_6481,N_3398);
or U15039 (N_15039,N_1545,N_7137);
nand U15040 (N_15040,N_996,N_1735);
nand U15041 (N_15041,N_3771,N_1534);
or U15042 (N_15042,N_4225,N_6114);
or U15043 (N_15043,N_4150,N_1543);
and U15044 (N_15044,N_2268,N_2922);
nand U15045 (N_15045,N_7356,N_8075);
nand U15046 (N_15046,N_6189,N_9658);
nor U15047 (N_15047,N_4627,N_340);
or U15048 (N_15048,N_6022,N_2604);
nor U15049 (N_15049,N_2241,N_9967);
nor U15050 (N_15050,N_7174,N_8553);
nor U15051 (N_15051,N_9594,N_8184);
nand U15052 (N_15052,N_6823,N_9379);
nand U15053 (N_15053,N_7002,N_5792);
and U15054 (N_15054,N_2359,N_5013);
or U15055 (N_15055,N_9367,N_3459);
nor U15056 (N_15056,N_7869,N_8593);
and U15057 (N_15057,N_313,N_7717);
and U15058 (N_15058,N_3123,N_5309);
nor U15059 (N_15059,N_1527,N_1424);
nand U15060 (N_15060,N_6505,N_9989);
and U15061 (N_15061,N_1224,N_6002);
nor U15062 (N_15062,N_7370,N_4192);
nand U15063 (N_15063,N_7314,N_5050);
and U15064 (N_15064,N_7901,N_9464);
nand U15065 (N_15065,N_1142,N_5796);
nor U15066 (N_15066,N_8187,N_5145);
or U15067 (N_15067,N_2793,N_5493);
nor U15068 (N_15068,N_6994,N_5723);
nand U15069 (N_15069,N_4238,N_5817);
and U15070 (N_15070,N_8963,N_108);
or U15071 (N_15071,N_5033,N_1647);
and U15072 (N_15072,N_567,N_2201);
and U15073 (N_15073,N_6441,N_6143);
or U15074 (N_15074,N_5465,N_6511);
nand U15075 (N_15075,N_5890,N_7726);
nand U15076 (N_15076,N_9416,N_2084);
nand U15077 (N_15077,N_2450,N_767);
nand U15078 (N_15078,N_5006,N_6895);
nor U15079 (N_15079,N_9998,N_8304);
or U15080 (N_15080,N_4248,N_4854);
nand U15081 (N_15081,N_5736,N_8869);
nand U15082 (N_15082,N_3974,N_5688);
nand U15083 (N_15083,N_5603,N_9160);
and U15084 (N_15084,N_1112,N_5555);
and U15085 (N_15085,N_6635,N_682);
and U15086 (N_15086,N_1133,N_2647);
and U15087 (N_15087,N_5979,N_29);
or U15088 (N_15088,N_4470,N_928);
nand U15089 (N_15089,N_3272,N_356);
nor U15090 (N_15090,N_663,N_8052);
or U15091 (N_15091,N_6757,N_8638);
nor U15092 (N_15092,N_4075,N_7187);
or U15093 (N_15093,N_6381,N_3764);
nand U15094 (N_15094,N_9362,N_6690);
nor U15095 (N_15095,N_3975,N_6527);
and U15096 (N_15096,N_8052,N_4619);
and U15097 (N_15097,N_7615,N_7658);
or U15098 (N_15098,N_5394,N_833);
nor U15099 (N_15099,N_8764,N_3101);
and U15100 (N_15100,N_9715,N_6766);
or U15101 (N_15101,N_9747,N_8797);
or U15102 (N_15102,N_9182,N_5555);
or U15103 (N_15103,N_7103,N_2060);
and U15104 (N_15104,N_9411,N_9109);
and U15105 (N_15105,N_7554,N_1175);
nor U15106 (N_15106,N_9843,N_9135);
nand U15107 (N_15107,N_3071,N_1976);
nor U15108 (N_15108,N_4012,N_8806);
nor U15109 (N_15109,N_9264,N_3326);
and U15110 (N_15110,N_1900,N_5989);
or U15111 (N_15111,N_236,N_3445);
or U15112 (N_15112,N_7521,N_7722);
nor U15113 (N_15113,N_1604,N_4583);
nand U15114 (N_15114,N_9778,N_9286);
or U15115 (N_15115,N_1942,N_3887);
nor U15116 (N_15116,N_9504,N_54);
nand U15117 (N_15117,N_4909,N_87);
nor U15118 (N_15118,N_3329,N_7514);
or U15119 (N_15119,N_9267,N_8047);
or U15120 (N_15120,N_4893,N_7441);
nor U15121 (N_15121,N_9303,N_1366);
and U15122 (N_15122,N_4007,N_9120);
nand U15123 (N_15123,N_4819,N_2149);
or U15124 (N_15124,N_7288,N_2061);
nor U15125 (N_15125,N_4912,N_7185);
nor U15126 (N_15126,N_7225,N_9873);
nand U15127 (N_15127,N_8876,N_8418);
and U15128 (N_15128,N_8443,N_9497);
or U15129 (N_15129,N_3739,N_4707);
and U15130 (N_15130,N_3646,N_7950);
and U15131 (N_15131,N_1943,N_843);
nor U15132 (N_15132,N_5107,N_3913);
or U15133 (N_15133,N_9286,N_6139);
nor U15134 (N_15134,N_6773,N_3197);
or U15135 (N_15135,N_8515,N_6746);
and U15136 (N_15136,N_7686,N_691);
nand U15137 (N_15137,N_361,N_9478);
nor U15138 (N_15138,N_3675,N_5816);
nor U15139 (N_15139,N_1030,N_2727);
nand U15140 (N_15140,N_251,N_7559);
and U15141 (N_15141,N_8911,N_2716);
and U15142 (N_15142,N_4269,N_5624);
and U15143 (N_15143,N_4232,N_9600);
nand U15144 (N_15144,N_9578,N_5734);
and U15145 (N_15145,N_4110,N_3731);
nor U15146 (N_15146,N_6703,N_5744);
and U15147 (N_15147,N_3294,N_9448);
nand U15148 (N_15148,N_543,N_1195);
nor U15149 (N_15149,N_9346,N_6994);
nand U15150 (N_15150,N_2087,N_6627);
and U15151 (N_15151,N_878,N_1164);
and U15152 (N_15152,N_6257,N_8263);
nor U15153 (N_15153,N_7603,N_5023);
or U15154 (N_15154,N_7010,N_9257);
or U15155 (N_15155,N_3197,N_8775);
and U15156 (N_15156,N_5434,N_3064);
nand U15157 (N_15157,N_6097,N_2698);
or U15158 (N_15158,N_3619,N_9787);
or U15159 (N_15159,N_6841,N_9984);
nor U15160 (N_15160,N_9231,N_982);
nand U15161 (N_15161,N_5317,N_8606);
nand U15162 (N_15162,N_7903,N_8467);
or U15163 (N_15163,N_5454,N_4440);
or U15164 (N_15164,N_7658,N_949);
nand U15165 (N_15165,N_5219,N_6057);
or U15166 (N_15166,N_6973,N_4261);
nor U15167 (N_15167,N_6938,N_168);
nand U15168 (N_15168,N_8498,N_7285);
and U15169 (N_15169,N_3091,N_1797);
nand U15170 (N_15170,N_6125,N_2183);
or U15171 (N_15171,N_4684,N_6253);
nand U15172 (N_15172,N_5481,N_8024);
nor U15173 (N_15173,N_1879,N_8057);
or U15174 (N_15174,N_9691,N_3428);
nor U15175 (N_15175,N_5414,N_8101);
or U15176 (N_15176,N_7464,N_1541);
or U15177 (N_15177,N_9961,N_6349);
and U15178 (N_15178,N_4864,N_3004);
xor U15179 (N_15179,N_4040,N_7179);
and U15180 (N_15180,N_9074,N_7629);
nand U15181 (N_15181,N_5441,N_1688);
and U15182 (N_15182,N_5715,N_4363);
and U15183 (N_15183,N_1359,N_5587);
nand U15184 (N_15184,N_9498,N_5295);
nand U15185 (N_15185,N_3001,N_934);
and U15186 (N_15186,N_673,N_3104);
and U15187 (N_15187,N_7128,N_5155);
nor U15188 (N_15188,N_4188,N_3410);
or U15189 (N_15189,N_8349,N_7336);
nor U15190 (N_15190,N_2940,N_9923);
or U15191 (N_15191,N_2543,N_2515);
nand U15192 (N_15192,N_9670,N_4319);
or U15193 (N_15193,N_8399,N_160);
nor U15194 (N_15194,N_4374,N_1955);
nor U15195 (N_15195,N_6010,N_7263);
nand U15196 (N_15196,N_2800,N_9714);
or U15197 (N_15197,N_1739,N_3936);
nand U15198 (N_15198,N_6622,N_4974);
nand U15199 (N_15199,N_4772,N_4221);
nor U15200 (N_15200,N_8867,N_3168);
nand U15201 (N_15201,N_5903,N_1080);
nand U15202 (N_15202,N_1090,N_6409);
nand U15203 (N_15203,N_5412,N_6332);
nor U15204 (N_15204,N_4840,N_1783);
or U15205 (N_15205,N_6081,N_331);
nand U15206 (N_15206,N_9374,N_8236);
or U15207 (N_15207,N_1736,N_9177);
nand U15208 (N_15208,N_3612,N_9693);
nor U15209 (N_15209,N_9418,N_6013);
and U15210 (N_15210,N_1437,N_295);
or U15211 (N_15211,N_5329,N_2525);
or U15212 (N_15212,N_822,N_6048);
nand U15213 (N_15213,N_5132,N_2871);
and U15214 (N_15214,N_634,N_685);
and U15215 (N_15215,N_7090,N_4546);
nor U15216 (N_15216,N_5134,N_1359);
or U15217 (N_15217,N_7582,N_7624);
and U15218 (N_15218,N_8756,N_3629);
or U15219 (N_15219,N_1445,N_9922);
and U15220 (N_15220,N_1898,N_453);
or U15221 (N_15221,N_7779,N_1006);
nor U15222 (N_15222,N_166,N_9309);
and U15223 (N_15223,N_8272,N_8143);
and U15224 (N_15224,N_9477,N_3599);
nand U15225 (N_15225,N_3292,N_9076);
and U15226 (N_15226,N_7210,N_9063);
nor U15227 (N_15227,N_9243,N_4413);
nor U15228 (N_15228,N_6994,N_4778);
nand U15229 (N_15229,N_7092,N_7599);
nor U15230 (N_15230,N_6974,N_6561);
or U15231 (N_15231,N_928,N_417);
nor U15232 (N_15232,N_235,N_8351);
nor U15233 (N_15233,N_162,N_8685);
nand U15234 (N_15234,N_5096,N_5175);
or U15235 (N_15235,N_9851,N_5065);
and U15236 (N_15236,N_629,N_9782);
nor U15237 (N_15237,N_638,N_7519);
nor U15238 (N_15238,N_7841,N_8638);
and U15239 (N_15239,N_9665,N_8723);
nand U15240 (N_15240,N_7930,N_1668);
and U15241 (N_15241,N_4591,N_1632);
or U15242 (N_15242,N_8626,N_4212);
and U15243 (N_15243,N_8405,N_8204);
or U15244 (N_15244,N_9346,N_1124);
nor U15245 (N_15245,N_6851,N_7743);
nand U15246 (N_15246,N_4480,N_312);
and U15247 (N_15247,N_7469,N_2996);
nor U15248 (N_15248,N_4182,N_2448);
nand U15249 (N_15249,N_2053,N_7898);
nor U15250 (N_15250,N_4985,N_5258);
nor U15251 (N_15251,N_9897,N_1040);
or U15252 (N_15252,N_6180,N_6802);
and U15253 (N_15253,N_6485,N_5419);
nor U15254 (N_15254,N_3394,N_1204);
nand U15255 (N_15255,N_4361,N_2173);
nand U15256 (N_15256,N_392,N_3012);
nand U15257 (N_15257,N_871,N_3464);
and U15258 (N_15258,N_7962,N_3017);
nor U15259 (N_15259,N_6595,N_9565);
nor U15260 (N_15260,N_2495,N_5584);
nor U15261 (N_15261,N_4738,N_1649);
and U15262 (N_15262,N_4420,N_6377);
nand U15263 (N_15263,N_7323,N_3251);
or U15264 (N_15264,N_8451,N_3513);
and U15265 (N_15265,N_8706,N_7524);
or U15266 (N_15266,N_9768,N_8778);
nand U15267 (N_15267,N_7550,N_1602);
and U15268 (N_15268,N_6227,N_9000);
and U15269 (N_15269,N_446,N_4365);
or U15270 (N_15270,N_5590,N_3018);
nor U15271 (N_15271,N_8003,N_241);
or U15272 (N_15272,N_5172,N_2216);
nor U15273 (N_15273,N_3758,N_5060);
nand U15274 (N_15274,N_2449,N_4296);
nand U15275 (N_15275,N_7521,N_4293);
and U15276 (N_15276,N_4339,N_6300);
nand U15277 (N_15277,N_7933,N_1886);
nand U15278 (N_15278,N_8706,N_1579);
nand U15279 (N_15279,N_6353,N_6618);
and U15280 (N_15280,N_1611,N_7054);
and U15281 (N_15281,N_5964,N_4310);
nand U15282 (N_15282,N_9436,N_6885);
and U15283 (N_15283,N_4677,N_6008);
or U15284 (N_15284,N_4413,N_1666);
or U15285 (N_15285,N_8841,N_4233);
nor U15286 (N_15286,N_844,N_384);
nor U15287 (N_15287,N_4144,N_6089);
nor U15288 (N_15288,N_8277,N_4544);
or U15289 (N_15289,N_4673,N_9959);
nor U15290 (N_15290,N_9802,N_6115);
and U15291 (N_15291,N_421,N_5920);
nor U15292 (N_15292,N_136,N_2433);
nand U15293 (N_15293,N_9379,N_8791);
and U15294 (N_15294,N_7707,N_3193);
and U15295 (N_15295,N_7233,N_9408);
or U15296 (N_15296,N_7492,N_2025);
and U15297 (N_15297,N_8826,N_2630);
nor U15298 (N_15298,N_1297,N_9183);
and U15299 (N_15299,N_448,N_2031);
and U15300 (N_15300,N_7539,N_3264);
nor U15301 (N_15301,N_8213,N_5689);
or U15302 (N_15302,N_5909,N_3106);
and U15303 (N_15303,N_1077,N_3661);
and U15304 (N_15304,N_2107,N_223);
or U15305 (N_15305,N_1741,N_2220);
nor U15306 (N_15306,N_3758,N_6099);
nor U15307 (N_15307,N_7180,N_9312);
or U15308 (N_15308,N_3438,N_8225);
or U15309 (N_15309,N_1614,N_1146);
or U15310 (N_15310,N_4473,N_6315);
or U15311 (N_15311,N_1652,N_3329);
or U15312 (N_15312,N_8816,N_5900);
and U15313 (N_15313,N_6083,N_1126);
nor U15314 (N_15314,N_2826,N_5469);
nand U15315 (N_15315,N_7578,N_2288);
nor U15316 (N_15316,N_356,N_559);
and U15317 (N_15317,N_8978,N_9575);
nand U15318 (N_15318,N_7919,N_2564);
or U15319 (N_15319,N_9622,N_3713);
or U15320 (N_15320,N_2209,N_2608);
or U15321 (N_15321,N_4691,N_6939);
and U15322 (N_15322,N_1486,N_4805);
nor U15323 (N_15323,N_2520,N_7804);
or U15324 (N_15324,N_7506,N_4473);
nand U15325 (N_15325,N_4740,N_1577);
and U15326 (N_15326,N_9284,N_5871);
or U15327 (N_15327,N_9119,N_5837);
or U15328 (N_15328,N_3681,N_1011);
or U15329 (N_15329,N_7585,N_4409);
or U15330 (N_15330,N_5076,N_3047);
and U15331 (N_15331,N_6238,N_9026);
nand U15332 (N_15332,N_2890,N_3256);
or U15333 (N_15333,N_5791,N_883);
or U15334 (N_15334,N_1769,N_1087);
nand U15335 (N_15335,N_1771,N_6339);
or U15336 (N_15336,N_2147,N_2109);
nor U15337 (N_15337,N_2746,N_6787);
and U15338 (N_15338,N_7719,N_6304);
and U15339 (N_15339,N_8709,N_7289);
nand U15340 (N_15340,N_9641,N_6803);
or U15341 (N_15341,N_9760,N_1257);
nand U15342 (N_15342,N_2054,N_9140);
nor U15343 (N_15343,N_1615,N_2076);
nor U15344 (N_15344,N_5414,N_8895);
or U15345 (N_15345,N_5788,N_2932);
nor U15346 (N_15346,N_2008,N_6830);
or U15347 (N_15347,N_5635,N_2498);
nor U15348 (N_15348,N_9252,N_9725);
nand U15349 (N_15349,N_1474,N_357);
nand U15350 (N_15350,N_2131,N_4285);
and U15351 (N_15351,N_8933,N_9251);
xor U15352 (N_15352,N_8199,N_2259);
nor U15353 (N_15353,N_1089,N_2642);
and U15354 (N_15354,N_5005,N_5673);
nand U15355 (N_15355,N_7236,N_2311);
nor U15356 (N_15356,N_5269,N_9731);
nand U15357 (N_15357,N_5220,N_3806);
nand U15358 (N_15358,N_5035,N_8355);
or U15359 (N_15359,N_4180,N_8129);
or U15360 (N_15360,N_8182,N_6079);
nand U15361 (N_15361,N_8105,N_4689);
or U15362 (N_15362,N_7365,N_8399);
nor U15363 (N_15363,N_9203,N_8744);
nor U15364 (N_15364,N_4650,N_2657);
and U15365 (N_15365,N_7466,N_3657);
nor U15366 (N_15366,N_5727,N_4642);
and U15367 (N_15367,N_7793,N_40);
or U15368 (N_15368,N_4424,N_402);
nor U15369 (N_15369,N_994,N_2543);
nor U15370 (N_15370,N_3296,N_3652);
nand U15371 (N_15371,N_8099,N_8463);
nor U15372 (N_15372,N_4139,N_8684);
or U15373 (N_15373,N_1790,N_1618);
nand U15374 (N_15374,N_3696,N_1547);
or U15375 (N_15375,N_2706,N_4783);
or U15376 (N_15376,N_4702,N_8287);
or U15377 (N_15377,N_907,N_6905);
nor U15378 (N_15378,N_4164,N_9364);
or U15379 (N_15379,N_6141,N_3427);
and U15380 (N_15380,N_3344,N_4904);
nand U15381 (N_15381,N_8014,N_7390);
and U15382 (N_15382,N_2346,N_9858);
and U15383 (N_15383,N_5688,N_3981);
or U15384 (N_15384,N_5550,N_1969);
or U15385 (N_15385,N_2313,N_4053);
or U15386 (N_15386,N_6301,N_2844);
nor U15387 (N_15387,N_7888,N_3585);
nand U15388 (N_15388,N_6072,N_2901);
and U15389 (N_15389,N_3525,N_5069);
nor U15390 (N_15390,N_3793,N_6531);
or U15391 (N_15391,N_8440,N_74);
xnor U15392 (N_15392,N_2787,N_4401);
nor U15393 (N_15393,N_1144,N_936);
nand U15394 (N_15394,N_7131,N_1697);
or U15395 (N_15395,N_6262,N_277);
and U15396 (N_15396,N_7808,N_2756);
and U15397 (N_15397,N_7433,N_8278);
or U15398 (N_15398,N_2509,N_6403);
nor U15399 (N_15399,N_1276,N_4062);
nor U15400 (N_15400,N_7253,N_8203);
or U15401 (N_15401,N_8116,N_2338);
xor U15402 (N_15402,N_5190,N_7936);
nor U15403 (N_15403,N_1393,N_423);
nand U15404 (N_15404,N_4355,N_703);
nor U15405 (N_15405,N_5811,N_2862);
nand U15406 (N_15406,N_2395,N_2908);
nand U15407 (N_15407,N_8742,N_2840);
or U15408 (N_15408,N_3438,N_8261);
or U15409 (N_15409,N_5077,N_8377);
nor U15410 (N_15410,N_3260,N_4488);
or U15411 (N_15411,N_5662,N_3380);
or U15412 (N_15412,N_4131,N_342);
nand U15413 (N_15413,N_9578,N_4873);
and U15414 (N_15414,N_9508,N_2824);
or U15415 (N_15415,N_1381,N_2300);
and U15416 (N_15416,N_1511,N_6008);
and U15417 (N_15417,N_7798,N_1170);
or U15418 (N_15418,N_1131,N_7700);
nand U15419 (N_15419,N_1047,N_5122);
or U15420 (N_15420,N_3114,N_5980);
nand U15421 (N_15421,N_5185,N_3815);
and U15422 (N_15422,N_8777,N_4029);
nand U15423 (N_15423,N_6452,N_5625);
or U15424 (N_15424,N_4198,N_8371);
nand U15425 (N_15425,N_2478,N_9950);
nor U15426 (N_15426,N_5452,N_7167);
nand U15427 (N_15427,N_7989,N_1386);
and U15428 (N_15428,N_2523,N_3600);
or U15429 (N_15429,N_2106,N_704);
nand U15430 (N_15430,N_561,N_9635);
nand U15431 (N_15431,N_673,N_5043);
nor U15432 (N_15432,N_5573,N_613);
or U15433 (N_15433,N_1061,N_150);
nand U15434 (N_15434,N_8265,N_3449);
nor U15435 (N_15435,N_7597,N_3532);
nand U15436 (N_15436,N_9148,N_886);
or U15437 (N_15437,N_558,N_5273);
and U15438 (N_15438,N_5314,N_5371);
or U15439 (N_15439,N_5121,N_600);
and U15440 (N_15440,N_8500,N_8326);
or U15441 (N_15441,N_4434,N_5482);
or U15442 (N_15442,N_7315,N_2755);
nor U15443 (N_15443,N_8008,N_7466);
nor U15444 (N_15444,N_7880,N_8339);
nor U15445 (N_15445,N_9967,N_4221);
xor U15446 (N_15446,N_5033,N_7958);
and U15447 (N_15447,N_9822,N_3280);
nor U15448 (N_15448,N_6076,N_1692);
and U15449 (N_15449,N_6420,N_7392);
and U15450 (N_15450,N_3321,N_7701);
nor U15451 (N_15451,N_5923,N_8318);
or U15452 (N_15452,N_6849,N_2462);
and U15453 (N_15453,N_1479,N_6299);
nand U15454 (N_15454,N_3798,N_396);
nand U15455 (N_15455,N_4360,N_4144);
or U15456 (N_15456,N_7895,N_8452);
and U15457 (N_15457,N_9558,N_2384);
nor U15458 (N_15458,N_805,N_9652);
nand U15459 (N_15459,N_969,N_4335);
and U15460 (N_15460,N_1018,N_6026);
nor U15461 (N_15461,N_2857,N_4597);
or U15462 (N_15462,N_5962,N_9754);
or U15463 (N_15463,N_3231,N_8593);
nor U15464 (N_15464,N_3120,N_3647);
or U15465 (N_15465,N_6489,N_8649);
nand U15466 (N_15466,N_5499,N_2065);
or U15467 (N_15467,N_4176,N_1480);
nor U15468 (N_15468,N_179,N_8592);
and U15469 (N_15469,N_1763,N_3612);
or U15470 (N_15470,N_6446,N_2466);
nor U15471 (N_15471,N_128,N_7468);
nor U15472 (N_15472,N_905,N_3173);
nor U15473 (N_15473,N_4713,N_7619);
and U15474 (N_15474,N_9821,N_6254);
nand U15475 (N_15475,N_1418,N_1652);
nand U15476 (N_15476,N_571,N_6136);
and U15477 (N_15477,N_7061,N_5391);
and U15478 (N_15478,N_5073,N_1398);
nor U15479 (N_15479,N_5033,N_1946);
and U15480 (N_15480,N_5675,N_2524);
or U15481 (N_15481,N_9418,N_5452);
or U15482 (N_15482,N_410,N_2305);
and U15483 (N_15483,N_3030,N_3752);
and U15484 (N_15484,N_9361,N_3550);
or U15485 (N_15485,N_3860,N_4689);
nand U15486 (N_15486,N_9473,N_870);
or U15487 (N_15487,N_4930,N_549);
or U15488 (N_15488,N_9833,N_1159);
and U15489 (N_15489,N_1603,N_7219);
nand U15490 (N_15490,N_7525,N_6255);
nand U15491 (N_15491,N_3683,N_7039);
or U15492 (N_15492,N_3371,N_2046);
or U15493 (N_15493,N_7760,N_5653);
nand U15494 (N_15494,N_4075,N_6359);
nand U15495 (N_15495,N_487,N_1473);
or U15496 (N_15496,N_7423,N_9441);
nand U15497 (N_15497,N_5002,N_6358);
nand U15498 (N_15498,N_9326,N_3241);
nand U15499 (N_15499,N_4389,N_356);
nor U15500 (N_15500,N_6871,N_9803);
or U15501 (N_15501,N_2168,N_3508);
nor U15502 (N_15502,N_9492,N_9545);
and U15503 (N_15503,N_8234,N_3183);
nor U15504 (N_15504,N_7593,N_6306);
and U15505 (N_15505,N_5946,N_6358);
or U15506 (N_15506,N_5779,N_7266);
or U15507 (N_15507,N_9150,N_7999);
and U15508 (N_15508,N_5301,N_6445);
nor U15509 (N_15509,N_598,N_6798);
nand U15510 (N_15510,N_782,N_2667);
nor U15511 (N_15511,N_1218,N_5270);
and U15512 (N_15512,N_311,N_2114);
and U15513 (N_15513,N_7015,N_7866);
nand U15514 (N_15514,N_931,N_7398);
nand U15515 (N_15515,N_8731,N_5413);
nand U15516 (N_15516,N_5236,N_5012);
nor U15517 (N_15517,N_734,N_8477);
and U15518 (N_15518,N_2233,N_3899);
nand U15519 (N_15519,N_4809,N_124);
and U15520 (N_15520,N_8038,N_9906);
or U15521 (N_15521,N_9149,N_4738);
or U15522 (N_15522,N_7840,N_4733);
nor U15523 (N_15523,N_5784,N_1100);
or U15524 (N_15524,N_1088,N_8226);
or U15525 (N_15525,N_1585,N_9790);
nand U15526 (N_15526,N_7551,N_9793);
and U15527 (N_15527,N_1122,N_3917);
and U15528 (N_15528,N_9798,N_6217);
nor U15529 (N_15529,N_8701,N_2626);
nand U15530 (N_15530,N_6068,N_2867);
nor U15531 (N_15531,N_5175,N_8178);
and U15532 (N_15532,N_6044,N_3953);
nand U15533 (N_15533,N_9945,N_1810);
or U15534 (N_15534,N_3624,N_4898);
and U15535 (N_15535,N_6220,N_6650);
nand U15536 (N_15536,N_7149,N_5970);
nor U15537 (N_15537,N_868,N_7443);
nor U15538 (N_15538,N_7664,N_6316);
and U15539 (N_15539,N_9558,N_8121);
nor U15540 (N_15540,N_1460,N_2666);
nor U15541 (N_15541,N_9928,N_5340);
and U15542 (N_15542,N_7264,N_2129);
nand U15543 (N_15543,N_7919,N_909);
nand U15544 (N_15544,N_2637,N_3305);
or U15545 (N_15545,N_8081,N_6149);
nand U15546 (N_15546,N_7894,N_9870);
and U15547 (N_15547,N_1410,N_4258);
nor U15548 (N_15548,N_4902,N_534);
and U15549 (N_15549,N_1521,N_2299);
and U15550 (N_15550,N_789,N_924);
and U15551 (N_15551,N_2537,N_4855);
nand U15552 (N_15552,N_9502,N_3079);
and U15553 (N_15553,N_5224,N_676);
nand U15554 (N_15554,N_9422,N_466);
or U15555 (N_15555,N_7526,N_9720);
nor U15556 (N_15556,N_446,N_5979);
nand U15557 (N_15557,N_5185,N_1823);
and U15558 (N_15558,N_8560,N_2740);
nor U15559 (N_15559,N_9085,N_5870);
or U15560 (N_15560,N_8068,N_4392);
and U15561 (N_15561,N_5411,N_1081);
or U15562 (N_15562,N_9348,N_6013);
nor U15563 (N_15563,N_9067,N_6854);
and U15564 (N_15564,N_3986,N_6317);
or U15565 (N_15565,N_9718,N_7007);
nor U15566 (N_15566,N_412,N_2166);
and U15567 (N_15567,N_7378,N_2237);
or U15568 (N_15568,N_7005,N_9785);
nand U15569 (N_15569,N_284,N_4627);
and U15570 (N_15570,N_8792,N_1207);
or U15571 (N_15571,N_9758,N_1737);
nand U15572 (N_15572,N_8087,N_6194);
or U15573 (N_15573,N_2959,N_1203);
nand U15574 (N_15574,N_8699,N_1432);
nand U15575 (N_15575,N_6464,N_4088);
nor U15576 (N_15576,N_3445,N_1921);
nand U15577 (N_15577,N_9575,N_9697);
nor U15578 (N_15578,N_5771,N_9124);
nor U15579 (N_15579,N_341,N_7443);
nor U15580 (N_15580,N_492,N_6636);
nand U15581 (N_15581,N_306,N_824);
nand U15582 (N_15582,N_356,N_4220);
and U15583 (N_15583,N_7710,N_4577);
nor U15584 (N_15584,N_7594,N_2810);
nor U15585 (N_15585,N_1856,N_2137);
or U15586 (N_15586,N_3035,N_9616);
nor U15587 (N_15587,N_3194,N_5026);
nand U15588 (N_15588,N_147,N_5698);
nor U15589 (N_15589,N_3232,N_6776);
nor U15590 (N_15590,N_3078,N_2251);
or U15591 (N_15591,N_329,N_7445);
or U15592 (N_15592,N_1241,N_4880);
nor U15593 (N_15593,N_1909,N_1947);
nor U15594 (N_15594,N_5917,N_8440);
or U15595 (N_15595,N_2464,N_5479);
nor U15596 (N_15596,N_9706,N_5922);
or U15597 (N_15597,N_5954,N_8747);
nor U15598 (N_15598,N_3762,N_8433);
nor U15599 (N_15599,N_8068,N_1678);
or U15600 (N_15600,N_252,N_7039);
nor U15601 (N_15601,N_5766,N_2035);
or U15602 (N_15602,N_7935,N_814);
nand U15603 (N_15603,N_3715,N_8489);
nand U15604 (N_15604,N_2848,N_8690);
and U15605 (N_15605,N_2539,N_3626);
or U15606 (N_15606,N_5131,N_5498);
or U15607 (N_15607,N_8470,N_8540);
or U15608 (N_15608,N_3701,N_3783);
or U15609 (N_15609,N_6546,N_4841);
and U15610 (N_15610,N_373,N_5580);
nand U15611 (N_15611,N_9297,N_8123);
nor U15612 (N_15612,N_7285,N_5419);
nor U15613 (N_15613,N_9450,N_8052);
or U15614 (N_15614,N_1679,N_8469);
and U15615 (N_15615,N_6664,N_6603);
and U15616 (N_15616,N_687,N_7251);
or U15617 (N_15617,N_5292,N_3220);
or U15618 (N_15618,N_3203,N_7182);
and U15619 (N_15619,N_7133,N_7911);
and U15620 (N_15620,N_3421,N_4721);
xnor U15621 (N_15621,N_4250,N_3375);
nor U15622 (N_15622,N_5897,N_4762);
and U15623 (N_15623,N_5165,N_6272);
nand U15624 (N_15624,N_4828,N_4631);
or U15625 (N_15625,N_5221,N_3358);
nor U15626 (N_15626,N_6920,N_5033);
nor U15627 (N_15627,N_6060,N_9926);
nand U15628 (N_15628,N_9355,N_3247);
or U15629 (N_15629,N_1821,N_278);
nor U15630 (N_15630,N_7603,N_2694);
or U15631 (N_15631,N_1871,N_2165);
and U15632 (N_15632,N_6628,N_475);
and U15633 (N_15633,N_8472,N_4877);
nor U15634 (N_15634,N_5420,N_6213);
or U15635 (N_15635,N_3769,N_2130);
or U15636 (N_15636,N_4114,N_4019);
nand U15637 (N_15637,N_4115,N_385);
nor U15638 (N_15638,N_2132,N_7777);
and U15639 (N_15639,N_286,N_3112);
or U15640 (N_15640,N_2788,N_202);
nand U15641 (N_15641,N_716,N_7361);
or U15642 (N_15642,N_4366,N_8239);
nand U15643 (N_15643,N_8528,N_8085);
or U15644 (N_15644,N_3693,N_6478);
nand U15645 (N_15645,N_3162,N_5125);
nor U15646 (N_15646,N_4472,N_4816);
nand U15647 (N_15647,N_3368,N_457);
nor U15648 (N_15648,N_4808,N_6127);
or U15649 (N_15649,N_9947,N_7220);
nand U15650 (N_15650,N_1207,N_8757);
and U15651 (N_15651,N_9305,N_1505);
nand U15652 (N_15652,N_5644,N_8568);
nor U15653 (N_15653,N_9959,N_5958);
or U15654 (N_15654,N_1381,N_2642);
or U15655 (N_15655,N_5916,N_1000);
and U15656 (N_15656,N_310,N_9567);
or U15657 (N_15657,N_4168,N_7181);
nand U15658 (N_15658,N_1834,N_169);
nand U15659 (N_15659,N_3127,N_5566);
and U15660 (N_15660,N_7263,N_1024);
and U15661 (N_15661,N_4475,N_3452);
or U15662 (N_15662,N_9794,N_5763);
or U15663 (N_15663,N_3637,N_9451);
and U15664 (N_15664,N_9528,N_7533);
nor U15665 (N_15665,N_5938,N_9936);
nor U15666 (N_15666,N_2809,N_9876);
nor U15667 (N_15667,N_8033,N_9952);
or U15668 (N_15668,N_4346,N_6848);
and U15669 (N_15669,N_2024,N_8613);
nor U15670 (N_15670,N_7066,N_5290);
nor U15671 (N_15671,N_5533,N_6394);
and U15672 (N_15672,N_8927,N_3150);
nor U15673 (N_15673,N_8875,N_6552);
nor U15674 (N_15674,N_1767,N_8119);
or U15675 (N_15675,N_7678,N_9042);
and U15676 (N_15676,N_1145,N_1224);
and U15677 (N_15677,N_3985,N_7055);
nor U15678 (N_15678,N_3422,N_3918);
and U15679 (N_15679,N_9663,N_3991);
nand U15680 (N_15680,N_3182,N_2421);
and U15681 (N_15681,N_5917,N_2102);
or U15682 (N_15682,N_8211,N_2013);
or U15683 (N_15683,N_9501,N_5826);
nor U15684 (N_15684,N_4782,N_2566);
and U15685 (N_15685,N_5663,N_1497);
nor U15686 (N_15686,N_6907,N_1724);
and U15687 (N_15687,N_8670,N_8417);
or U15688 (N_15688,N_928,N_5925);
or U15689 (N_15689,N_5275,N_3673);
or U15690 (N_15690,N_8903,N_4483);
or U15691 (N_15691,N_897,N_3011);
nor U15692 (N_15692,N_1990,N_8932);
and U15693 (N_15693,N_6159,N_8777);
or U15694 (N_15694,N_7406,N_4621);
or U15695 (N_15695,N_1364,N_8515);
or U15696 (N_15696,N_9053,N_3018);
nor U15697 (N_15697,N_7587,N_9297);
nor U15698 (N_15698,N_1996,N_4312);
xor U15699 (N_15699,N_9588,N_2511);
nor U15700 (N_15700,N_1597,N_8380);
or U15701 (N_15701,N_9034,N_8793);
nor U15702 (N_15702,N_7237,N_4329);
nand U15703 (N_15703,N_6064,N_4991);
or U15704 (N_15704,N_9970,N_8055);
or U15705 (N_15705,N_8700,N_9359);
or U15706 (N_15706,N_3748,N_5937);
or U15707 (N_15707,N_7039,N_1740);
nand U15708 (N_15708,N_8833,N_8275);
and U15709 (N_15709,N_34,N_5993);
xnor U15710 (N_15710,N_9695,N_6838);
and U15711 (N_15711,N_4464,N_5743);
nand U15712 (N_15712,N_3232,N_2438);
and U15713 (N_15713,N_6833,N_1227);
nand U15714 (N_15714,N_228,N_7904);
or U15715 (N_15715,N_6550,N_8254);
nand U15716 (N_15716,N_1735,N_3405);
nand U15717 (N_15717,N_1848,N_2754);
nand U15718 (N_15718,N_1514,N_969);
and U15719 (N_15719,N_6377,N_2835);
nand U15720 (N_15720,N_4418,N_1839);
or U15721 (N_15721,N_5686,N_9103);
and U15722 (N_15722,N_6135,N_7624);
nand U15723 (N_15723,N_4449,N_6917);
nand U15724 (N_15724,N_3390,N_3213);
or U15725 (N_15725,N_401,N_5619);
nor U15726 (N_15726,N_5197,N_7868);
nor U15727 (N_15727,N_8907,N_209);
or U15728 (N_15728,N_3345,N_1442);
and U15729 (N_15729,N_5567,N_4671);
and U15730 (N_15730,N_38,N_6379);
or U15731 (N_15731,N_4195,N_2070);
or U15732 (N_15732,N_3397,N_9229);
or U15733 (N_15733,N_2726,N_7578);
nand U15734 (N_15734,N_211,N_7839);
nor U15735 (N_15735,N_6479,N_831);
nand U15736 (N_15736,N_7566,N_4939);
nand U15737 (N_15737,N_1291,N_5625);
nand U15738 (N_15738,N_6104,N_7909);
nand U15739 (N_15739,N_4502,N_6707);
nand U15740 (N_15740,N_6414,N_965);
nand U15741 (N_15741,N_4864,N_310);
nor U15742 (N_15742,N_6109,N_9427);
nor U15743 (N_15743,N_2731,N_8330);
nand U15744 (N_15744,N_9752,N_5348);
nor U15745 (N_15745,N_6583,N_563);
nor U15746 (N_15746,N_6861,N_4733);
nor U15747 (N_15747,N_4575,N_6186);
or U15748 (N_15748,N_8981,N_6411);
or U15749 (N_15749,N_5777,N_9334);
and U15750 (N_15750,N_5010,N_7607);
nand U15751 (N_15751,N_8536,N_1435);
or U15752 (N_15752,N_4427,N_7565);
nand U15753 (N_15753,N_8668,N_5188);
xnor U15754 (N_15754,N_8046,N_7543);
xor U15755 (N_15755,N_795,N_5542);
nand U15756 (N_15756,N_4061,N_2010);
nand U15757 (N_15757,N_6642,N_1970);
nand U15758 (N_15758,N_9077,N_6135);
nand U15759 (N_15759,N_6307,N_9263);
or U15760 (N_15760,N_4905,N_6581);
or U15761 (N_15761,N_8964,N_5325);
and U15762 (N_15762,N_3630,N_4392);
xor U15763 (N_15763,N_3404,N_6780);
nand U15764 (N_15764,N_9959,N_8211);
nor U15765 (N_15765,N_4126,N_2019);
nor U15766 (N_15766,N_5551,N_9782);
nor U15767 (N_15767,N_8031,N_6227);
nor U15768 (N_15768,N_9949,N_5117);
and U15769 (N_15769,N_4126,N_9047);
and U15770 (N_15770,N_1100,N_2430);
and U15771 (N_15771,N_7273,N_664);
or U15772 (N_15772,N_6694,N_4260);
and U15773 (N_15773,N_4546,N_8629);
nor U15774 (N_15774,N_2901,N_2625);
and U15775 (N_15775,N_9716,N_3088);
and U15776 (N_15776,N_6654,N_7526);
nand U15777 (N_15777,N_5341,N_8962);
or U15778 (N_15778,N_5350,N_2475);
nand U15779 (N_15779,N_6749,N_1185);
nor U15780 (N_15780,N_1610,N_9443);
nand U15781 (N_15781,N_7659,N_9133);
or U15782 (N_15782,N_2010,N_6222);
nand U15783 (N_15783,N_2419,N_9546);
nand U15784 (N_15784,N_4700,N_4650);
nor U15785 (N_15785,N_5382,N_5887);
or U15786 (N_15786,N_7572,N_1209);
or U15787 (N_15787,N_8019,N_1734);
or U15788 (N_15788,N_6323,N_5148);
and U15789 (N_15789,N_1696,N_5040);
nand U15790 (N_15790,N_4584,N_4901);
and U15791 (N_15791,N_9581,N_8703);
and U15792 (N_15792,N_8127,N_1362);
and U15793 (N_15793,N_8927,N_4288);
nand U15794 (N_15794,N_4630,N_7402);
or U15795 (N_15795,N_7468,N_4065);
or U15796 (N_15796,N_3823,N_3273);
or U15797 (N_15797,N_5067,N_6071);
or U15798 (N_15798,N_8619,N_4058);
nand U15799 (N_15799,N_1327,N_593);
and U15800 (N_15800,N_2142,N_1173);
nor U15801 (N_15801,N_2201,N_9315);
nor U15802 (N_15802,N_5264,N_6575);
nor U15803 (N_15803,N_9877,N_9645);
nand U15804 (N_15804,N_8236,N_6429);
nand U15805 (N_15805,N_8955,N_3642);
and U15806 (N_15806,N_7954,N_5807);
xor U15807 (N_15807,N_9492,N_4423);
nor U15808 (N_15808,N_5143,N_5309);
nor U15809 (N_15809,N_5920,N_3666);
nor U15810 (N_15810,N_8516,N_9289);
nor U15811 (N_15811,N_510,N_8666);
nand U15812 (N_15812,N_8307,N_9001);
nand U15813 (N_15813,N_8823,N_4449);
nand U15814 (N_15814,N_9718,N_5495);
nand U15815 (N_15815,N_643,N_5465);
nand U15816 (N_15816,N_3422,N_6548);
or U15817 (N_15817,N_39,N_8375);
and U15818 (N_15818,N_9766,N_9786);
nor U15819 (N_15819,N_1234,N_5515);
and U15820 (N_15820,N_6630,N_9707);
and U15821 (N_15821,N_5446,N_3208);
and U15822 (N_15822,N_3900,N_5562);
nor U15823 (N_15823,N_9396,N_9558);
or U15824 (N_15824,N_4846,N_3565);
nand U15825 (N_15825,N_9380,N_2516);
and U15826 (N_15826,N_303,N_3024);
and U15827 (N_15827,N_621,N_7542);
nor U15828 (N_15828,N_3099,N_2513);
nor U15829 (N_15829,N_2421,N_797);
nand U15830 (N_15830,N_696,N_4062);
or U15831 (N_15831,N_840,N_3891);
nand U15832 (N_15832,N_1050,N_1335);
nand U15833 (N_15833,N_9632,N_3144);
nor U15834 (N_15834,N_9069,N_8172);
and U15835 (N_15835,N_3735,N_9049);
nand U15836 (N_15836,N_7552,N_5513);
nand U15837 (N_15837,N_7977,N_9935);
nand U15838 (N_15838,N_3387,N_3367);
and U15839 (N_15839,N_3953,N_9365);
and U15840 (N_15840,N_382,N_128);
or U15841 (N_15841,N_4362,N_1760);
nor U15842 (N_15842,N_5413,N_5857);
nor U15843 (N_15843,N_2175,N_7872);
nand U15844 (N_15844,N_3249,N_5355);
and U15845 (N_15845,N_1113,N_622);
nor U15846 (N_15846,N_4483,N_9493);
or U15847 (N_15847,N_2290,N_6278);
nand U15848 (N_15848,N_4301,N_7327);
or U15849 (N_15849,N_5587,N_8865);
nand U15850 (N_15850,N_5915,N_9956);
nand U15851 (N_15851,N_4124,N_6235);
and U15852 (N_15852,N_7051,N_8300);
or U15853 (N_15853,N_4819,N_4429);
nor U15854 (N_15854,N_6855,N_9013);
and U15855 (N_15855,N_5978,N_4611);
and U15856 (N_15856,N_1036,N_3389);
or U15857 (N_15857,N_59,N_9765);
nand U15858 (N_15858,N_4770,N_762);
nor U15859 (N_15859,N_4521,N_1955);
or U15860 (N_15860,N_306,N_3973);
and U15861 (N_15861,N_4652,N_7420);
and U15862 (N_15862,N_132,N_699);
nor U15863 (N_15863,N_3683,N_4383);
nand U15864 (N_15864,N_4765,N_2329);
nand U15865 (N_15865,N_5002,N_4125);
nor U15866 (N_15866,N_8302,N_9092);
nor U15867 (N_15867,N_3754,N_4434);
and U15868 (N_15868,N_6623,N_8058);
and U15869 (N_15869,N_4149,N_4726);
nand U15870 (N_15870,N_358,N_9401);
nand U15871 (N_15871,N_1001,N_3288);
and U15872 (N_15872,N_974,N_1193);
and U15873 (N_15873,N_1947,N_3609);
and U15874 (N_15874,N_6963,N_4847);
or U15875 (N_15875,N_8166,N_5018);
or U15876 (N_15876,N_7627,N_3595);
nor U15877 (N_15877,N_3201,N_8504);
and U15878 (N_15878,N_9081,N_4065);
nor U15879 (N_15879,N_9025,N_2639);
or U15880 (N_15880,N_7085,N_103);
nor U15881 (N_15881,N_3544,N_1922);
nand U15882 (N_15882,N_5966,N_5979);
nor U15883 (N_15883,N_1998,N_7867);
and U15884 (N_15884,N_5452,N_3926);
and U15885 (N_15885,N_2775,N_5372);
nand U15886 (N_15886,N_7979,N_1259);
nor U15887 (N_15887,N_9739,N_6259);
and U15888 (N_15888,N_3558,N_2430);
nor U15889 (N_15889,N_2709,N_2662);
nor U15890 (N_15890,N_8792,N_2084);
nor U15891 (N_15891,N_7080,N_161);
nand U15892 (N_15892,N_1878,N_6308);
and U15893 (N_15893,N_758,N_7595);
or U15894 (N_15894,N_6685,N_676);
nor U15895 (N_15895,N_8161,N_4068);
or U15896 (N_15896,N_8662,N_3360);
nor U15897 (N_15897,N_450,N_3940);
nand U15898 (N_15898,N_6491,N_2827);
and U15899 (N_15899,N_4245,N_4559);
or U15900 (N_15900,N_2206,N_4914);
or U15901 (N_15901,N_4468,N_7294);
nand U15902 (N_15902,N_6621,N_412);
nand U15903 (N_15903,N_5629,N_3530);
and U15904 (N_15904,N_5926,N_6080);
or U15905 (N_15905,N_7132,N_9840);
or U15906 (N_15906,N_8904,N_7718);
or U15907 (N_15907,N_3598,N_1187);
or U15908 (N_15908,N_126,N_8056);
nand U15909 (N_15909,N_4395,N_3637);
nor U15910 (N_15910,N_2745,N_1365);
nor U15911 (N_15911,N_3988,N_6326);
nand U15912 (N_15912,N_6855,N_4976);
and U15913 (N_15913,N_9327,N_2388);
or U15914 (N_15914,N_9060,N_4153);
or U15915 (N_15915,N_2735,N_845);
and U15916 (N_15916,N_7102,N_6308);
nand U15917 (N_15917,N_1796,N_7984);
and U15918 (N_15918,N_6139,N_2816);
or U15919 (N_15919,N_7809,N_6748);
or U15920 (N_15920,N_8969,N_5633);
nand U15921 (N_15921,N_3327,N_4753);
nor U15922 (N_15922,N_4581,N_9443);
or U15923 (N_15923,N_2402,N_2516);
and U15924 (N_15924,N_3252,N_1068);
nand U15925 (N_15925,N_1958,N_9441);
nor U15926 (N_15926,N_5825,N_896);
nor U15927 (N_15927,N_4938,N_7615);
nand U15928 (N_15928,N_7457,N_6889);
nand U15929 (N_15929,N_6006,N_2122);
nand U15930 (N_15930,N_1159,N_2518);
and U15931 (N_15931,N_7041,N_2718);
nand U15932 (N_15932,N_2583,N_2906);
nor U15933 (N_15933,N_9197,N_3276);
nor U15934 (N_15934,N_6692,N_1772);
and U15935 (N_15935,N_6331,N_5723);
nand U15936 (N_15936,N_9716,N_1131);
or U15937 (N_15937,N_1310,N_1176);
and U15938 (N_15938,N_3683,N_4960);
and U15939 (N_15939,N_6685,N_572);
or U15940 (N_15940,N_227,N_1993);
nor U15941 (N_15941,N_3411,N_7196);
nand U15942 (N_15942,N_7194,N_1841);
nand U15943 (N_15943,N_8845,N_9823);
nand U15944 (N_15944,N_3220,N_2817);
nor U15945 (N_15945,N_4908,N_3968);
or U15946 (N_15946,N_2262,N_6368);
nor U15947 (N_15947,N_6339,N_4189);
and U15948 (N_15948,N_9716,N_4619);
or U15949 (N_15949,N_8784,N_93);
nand U15950 (N_15950,N_5168,N_6349);
nor U15951 (N_15951,N_1559,N_8467);
and U15952 (N_15952,N_5061,N_3968);
and U15953 (N_15953,N_4949,N_123);
or U15954 (N_15954,N_9946,N_9362);
nand U15955 (N_15955,N_6319,N_8239);
nor U15956 (N_15956,N_9013,N_6671);
or U15957 (N_15957,N_6897,N_7011);
or U15958 (N_15958,N_2171,N_7753);
nand U15959 (N_15959,N_1588,N_7524);
nand U15960 (N_15960,N_5787,N_1877);
and U15961 (N_15961,N_3515,N_5782);
and U15962 (N_15962,N_3299,N_8119);
or U15963 (N_15963,N_6548,N_2857);
and U15964 (N_15964,N_6952,N_5401);
nor U15965 (N_15965,N_3336,N_8634);
and U15966 (N_15966,N_2763,N_5045);
or U15967 (N_15967,N_646,N_7946);
or U15968 (N_15968,N_2478,N_3799);
nor U15969 (N_15969,N_3577,N_2855);
nor U15970 (N_15970,N_1703,N_5197);
or U15971 (N_15971,N_8338,N_5046);
and U15972 (N_15972,N_8534,N_2946);
and U15973 (N_15973,N_5959,N_3543);
nor U15974 (N_15974,N_9200,N_1182);
and U15975 (N_15975,N_4593,N_9016);
xnor U15976 (N_15976,N_4340,N_7127);
and U15977 (N_15977,N_6052,N_2618);
nand U15978 (N_15978,N_7455,N_3757);
or U15979 (N_15979,N_6074,N_1288);
or U15980 (N_15980,N_550,N_6695);
and U15981 (N_15981,N_590,N_414);
and U15982 (N_15982,N_1789,N_7734);
or U15983 (N_15983,N_1513,N_497);
or U15984 (N_15984,N_4575,N_2455);
or U15985 (N_15985,N_2860,N_6166);
nand U15986 (N_15986,N_5314,N_475);
nand U15987 (N_15987,N_4434,N_7869);
or U15988 (N_15988,N_6053,N_197);
nand U15989 (N_15989,N_676,N_3123);
and U15990 (N_15990,N_6436,N_9416);
nand U15991 (N_15991,N_4627,N_8733);
or U15992 (N_15992,N_1134,N_9091);
nor U15993 (N_15993,N_9299,N_344);
nor U15994 (N_15994,N_7349,N_6516);
nand U15995 (N_15995,N_382,N_6700);
nand U15996 (N_15996,N_8287,N_2789);
and U15997 (N_15997,N_5622,N_1613);
nand U15998 (N_15998,N_862,N_834);
and U15999 (N_15999,N_9404,N_5597);
and U16000 (N_16000,N_2718,N_2903);
nor U16001 (N_16001,N_4088,N_8353);
or U16002 (N_16002,N_4061,N_5947);
and U16003 (N_16003,N_418,N_9053);
nor U16004 (N_16004,N_8129,N_7953);
nor U16005 (N_16005,N_7772,N_2499);
and U16006 (N_16006,N_171,N_2562);
or U16007 (N_16007,N_4914,N_3227);
nand U16008 (N_16008,N_6980,N_2838);
or U16009 (N_16009,N_3514,N_7929);
nor U16010 (N_16010,N_7978,N_5448);
nor U16011 (N_16011,N_6733,N_6580);
nand U16012 (N_16012,N_9403,N_4670);
nand U16013 (N_16013,N_8331,N_198);
and U16014 (N_16014,N_45,N_9644);
nor U16015 (N_16015,N_9632,N_104);
nor U16016 (N_16016,N_7198,N_557);
or U16017 (N_16017,N_3489,N_3334);
or U16018 (N_16018,N_5862,N_1455);
nand U16019 (N_16019,N_2559,N_6290);
and U16020 (N_16020,N_6541,N_6982);
or U16021 (N_16021,N_5400,N_1648);
nand U16022 (N_16022,N_3667,N_9352);
nor U16023 (N_16023,N_8358,N_3302);
nand U16024 (N_16024,N_2592,N_4068);
nand U16025 (N_16025,N_8503,N_8819);
nor U16026 (N_16026,N_4924,N_4909);
nand U16027 (N_16027,N_2425,N_232);
and U16028 (N_16028,N_1678,N_8324);
or U16029 (N_16029,N_7022,N_5199);
or U16030 (N_16030,N_8619,N_4301);
and U16031 (N_16031,N_8411,N_9094);
and U16032 (N_16032,N_9635,N_4899);
or U16033 (N_16033,N_5676,N_7272);
and U16034 (N_16034,N_6967,N_631);
or U16035 (N_16035,N_2613,N_6153);
nor U16036 (N_16036,N_6677,N_6470);
or U16037 (N_16037,N_6490,N_9524);
xor U16038 (N_16038,N_8477,N_8637);
or U16039 (N_16039,N_9862,N_1802);
nand U16040 (N_16040,N_694,N_4982);
and U16041 (N_16041,N_1437,N_7594);
and U16042 (N_16042,N_2898,N_798);
and U16043 (N_16043,N_167,N_40);
nand U16044 (N_16044,N_6478,N_1864);
and U16045 (N_16045,N_896,N_3668);
nor U16046 (N_16046,N_2526,N_3470);
and U16047 (N_16047,N_901,N_840);
or U16048 (N_16048,N_1997,N_1534);
or U16049 (N_16049,N_8990,N_5400);
nor U16050 (N_16050,N_53,N_8291);
or U16051 (N_16051,N_4935,N_9443);
nor U16052 (N_16052,N_6836,N_5478);
nor U16053 (N_16053,N_8625,N_6350);
nor U16054 (N_16054,N_9090,N_7721);
nor U16055 (N_16055,N_1503,N_3704);
and U16056 (N_16056,N_1732,N_1875);
or U16057 (N_16057,N_1832,N_176);
or U16058 (N_16058,N_7561,N_2888);
nand U16059 (N_16059,N_12,N_304);
or U16060 (N_16060,N_8205,N_2270);
and U16061 (N_16061,N_9116,N_3558);
nor U16062 (N_16062,N_8590,N_7483);
nand U16063 (N_16063,N_8598,N_7653);
nor U16064 (N_16064,N_1040,N_6902);
nor U16065 (N_16065,N_3786,N_933);
nand U16066 (N_16066,N_8281,N_1626);
and U16067 (N_16067,N_1544,N_2807);
or U16068 (N_16068,N_1231,N_3024);
nand U16069 (N_16069,N_3855,N_2219);
or U16070 (N_16070,N_6127,N_4148);
nand U16071 (N_16071,N_6881,N_763);
nand U16072 (N_16072,N_1360,N_6711);
nand U16073 (N_16073,N_606,N_3115);
nand U16074 (N_16074,N_4466,N_1152);
nand U16075 (N_16075,N_36,N_6479);
nor U16076 (N_16076,N_9128,N_3063);
xnor U16077 (N_16077,N_6004,N_1305);
and U16078 (N_16078,N_8430,N_9948);
nand U16079 (N_16079,N_3690,N_396);
nor U16080 (N_16080,N_7021,N_5365);
or U16081 (N_16081,N_2102,N_5843);
or U16082 (N_16082,N_3389,N_7925);
or U16083 (N_16083,N_9637,N_2473);
nand U16084 (N_16084,N_2408,N_3991);
nor U16085 (N_16085,N_3062,N_1631);
and U16086 (N_16086,N_2624,N_5816);
nand U16087 (N_16087,N_3027,N_3508);
nand U16088 (N_16088,N_6003,N_8485);
or U16089 (N_16089,N_4319,N_9293);
or U16090 (N_16090,N_6106,N_296);
or U16091 (N_16091,N_5346,N_5974);
or U16092 (N_16092,N_2922,N_6488);
nor U16093 (N_16093,N_7485,N_3658);
or U16094 (N_16094,N_7848,N_6295);
or U16095 (N_16095,N_5887,N_925);
nand U16096 (N_16096,N_5532,N_7706);
nor U16097 (N_16097,N_6426,N_9522);
nand U16098 (N_16098,N_3497,N_8218);
nand U16099 (N_16099,N_7467,N_2902);
nand U16100 (N_16100,N_2918,N_4830);
and U16101 (N_16101,N_4452,N_3387);
nand U16102 (N_16102,N_2444,N_3005);
or U16103 (N_16103,N_6139,N_9989);
or U16104 (N_16104,N_8604,N_5231);
nand U16105 (N_16105,N_5858,N_2198);
and U16106 (N_16106,N_5947,N_4739);
nor U16107 (N_16107,N_6951,N_3545);
nor U16108 (N_16108,N_5276,N_8981);
or U16109 (N_16109,N_4467,N_4317);
or U16110 (N_16110,N_7471,N_5583);
nor U16111 (N_16111,N_3679,N_8119);
nor U16112 (N_16112,N_85,N_4011);
or U16113 (N_16113,N_236,N_8066);
and U16114 (N_16114,N_2549,N_4277);
nor U16115 (N_16115,N_5998,N_5297);
nor U16116 (N_16116,N_1869,N_9004);
nor U16117 (N_16117,N_161,N_929);
and U16118 (N_16118,N_4064,N_8795);
nand U16119 (N_16119,N_6473,N_6485);
nand U16120 (N_16120,N_8893,N_2748);
or U16121 (N_16121,N_3445,N_7643);
nand U16122 (N_16122,N_9168,N_6931);
and U16123 (N_16123,N_2442,N_707);
and U16124 (N_16124,N_9604,N_7065);
nor U16125 (N_16125,N_3341,N_856);
nor U16126 (N_16126,N_6684,N_278);
nand U16127 (N_16127,N_3270,N_804);
nand U16128 (N_16128,N_4172,N_8765);
xnor U16129 (N_16129,N_6484,N_5034);
or U16130 (N_16130,N_353,N_9425);
nor U16131 (N_16131,N_1735,N_3325);
nand U16132 (N_16132,N_3558,N_6804);
nor U16133 (N_16133,N_1201,N_3764);
nand U16134 (N_16134,N_3382,N_4745);
nor U16135 (N_16135,N_4922,N_8671);
or U16136 (N_16136,N_3525,N_4774);
or U16137 (N_16137,N_9085,N_9210);
or U16138 (N_16138,N_6631,N_7897);
nand U16139 (N_16139,N_1407,N_7730);
or U16140 (N_16140,N_7740,N_4809);
nor U16141 (N_16141,N_8485,N_7455);
nor U16142 (N_16142,N_6741,N_4724);
nand U16143 (N_16143,N_6678,N_7795);
nand U16144 (N_16144,N_2808,N_7085);
nand U16145 (N_16145,N_6606,N_8273);
and U16146 (N_16146,N_1161,N_2837);
nor U16147 (N_16147,N_8132,N_3280);
nor U16148 (N_16148,N_7675,N_1776);
nand U16149 (N_16149,N_9470,N_5184);
nand U16150 (N_16150,N_5368,N_9464);
nand U16151 (N_16151,N_7532,N_3486);
nor U16152 (N_16152,N_1356,N_5748);
or U16153 (N_16153,N_627,N_5854);
and U16154 (N_16154,N_1832,N_4227);
nand U16155 (N_16155,N_2608,N_3586);
nor U16156 (N_16156,N_3677,N_7862);
nand U16157 (N_16157,N_1085,N_4876);
nor U16158 (N_16158,N_8313,N_8799);
and U16159 (N_16159,N_3989,N_2830);
or U16160 (N_16160,N_1797,N_8439);
or U16161 (N_16161,N_4917,N_2171);
and U16162 (N_16162,N_1550,N_6898);
nor U16163 (N_16163,N_7891,N_6854);
or U16164 (N_16164,N_6718,N_6572);
nor U16165 (N_16165,N_5179,N_8121);
and U16166 (N_16166,N_4167,N_4260);
or U16167 (N_16167,N_2610,N_4726);
nor U16168 (N_16168,N_749,N_9445);
and U16169 (N_16169,N_6210,N_4990);
nand U16170 (N_16170,N_6044,N_8644);
or U16171 (N_16171,N_4433,N_969);
nor U16172 (N_16172,N_9884,N_8792);
and U16173 (N_16173,N_5265,N_939);
and U16174 (N_16174,N_1448,N_314);
or U16175 (N_16175,N_8767,N_3227);
and U16176 (N_16176,N_7713,N_8961);
or U16177 (N_16177,N_8516,N_7253);
and U16178 (N_16178,N_2783,N_3094);
and U16179 (N_16179,N_5020,N_3402);
xnor U16180 (N_16180,N_2363,N_3659);
and U16181 (N_16181,N_1849,N_1148);
nand U16182 (N_16182,N_2566,N_6985);
nand U16183 (N_16183,N_6450,N_6468);
or U16184 (N_16184,N_6270,N_4539);
or U16185 (N_16185,N_5141,N_2142);
and U16186 (N_16186,N_3799,N_6478);
or U16187 (N_16187,N_4338,N_4466);
nor U16188 (N_16188,N_7770,N_8163);
or U16189 (N_16189,N_7042,N_5977);
or U16190 (N_16190,N_9961,N_740);
or U16191 (N_16191,N_7593,N_7906);
and U16192 (N_16192,N_6716,N_137);
nand U16193 (N_16193,N_237,N_2374);
nor U16194 (N_16194,N_9498,N_4506);
nand U16195 (N_16195,N_5618,N_6338);
or U16196 (N_16196,N_1080,N_7690);
and U16197 (N_16197,N_4185,N_2400);
nor U16198 (N_16198,N_1355,N_7320);
and U16199 (N_16199,N_3065,N_9993);
nand U16200 (N_16200,N_1804,N_473);
and U16201 (N_16201,N_2052,N_3073);
nor U16202 (N_16202,N_6471,N_5484);
or U16203 (N_16203,N_4875,N_5782);
and U16204 (N_16204,N_6459,N_9641);
or U16205 (N_16205,N_5808,N_2392);
and U16206 (N_16206,N_9906,N_8422);
nor U16207 (N_16207,N_6691,N_3632);
nand U16208 (N_16208,N_179,N_7720);
nor U16209 (N_16209,N_8848,N_6631);
and U16210 (N_16210,N_4181,N_2739);
nand U16211 (N_16211,N_6788,N_9709);
or U16212 (N_16212,N_9199,N_3414);
nor U16213 (N_16213,N_9304,N_3970);
and U16214 (N_16214,N_8137,N_5732);
nor U16215 (N_16215,N_5784,N_3723);
or U16216 (N_16216,N_1342,N_3971);
or U16217 (N_16217,N_7914,N_7192);
nor U16218 (N_16218,N_6726,N_2491);
or U16219 (N_16219,N_9855,N_309);
or U16220 (N_16220,N_4276,N_4137);
or U16221 (N_16221,N_1559,N_5644);
nand U16222 (N_16222,N_5312,N_9090);
and U16223 (N_16223,N_9009,N_6977);
and U16224 (N_16224,N_4937,N_5804);
and U16225 (N_16225,N_1273,N_9129);
nor U16226 (N_16226,N_9360,N_1945);
nor U16227 (N_16227,N_7674,N_4946);
and U16228 (N_16228,N_465,N_5317);
or U16229 (N_16229,N_5977,N_5875);
nand U16230 (N_16230,N_2350,N_3722);
nor U16231 (N_16231,N_3552,N_4697);
nand U16232 (N_16232,N_5936,N_4910);
or U16233 (N_16233,N_586,N_4087);
and U16234 (N_16234,N_4041,N_3927);
nor U16235 (N_16235,N_1993,N_6862);
nand U16236 (N_16236,N_3642,N_4418);
and U16237 (N_16237,N_1578,N_4498);
nand U16238 (N_16238,N_3189,N_286);
and U16239 (N_16239,N_494,N_9060);
nand U16240 (N_16240,N_170,N_7655);
nand U16241 (N_16241,N_6006,N_5037);
nor U16242 (N_16242,N_2150,N_9187);
and U16243 (N_16243,N_5177,N_3621);
nor U16244 (N_16244,N_8262,N_9882);
and U16245 (N_16245,N_6551,N_1232);
and U16246 (N_16246,N_84,N_3514);
or U16247 (N_16247,N_2775,N_3041);
or U16248 (N_16248,N_6344,N_1813);
nor U16249 (N_16249,N_3688,N_4540);
nand U16250 (N_16250,N_9320,N_1343);
and U16251 (N_16251,N_1406,N_8240);
and U16252 (N_16252,N_2520,N_4865);
nand U16253 (N_16253,N_4112,N_9253);
nand U16254 (N_16254,N_7905,N_4925);
nor U16255 (N_16255,N_3103,N_1154);
xor U16256 (N_16256,N_7276,N_2930);
or U16257 (N_16257,N_2188,N_9772);
or U16258 (N_16258,N_3116,N_6494);
and U16259 (N_16259,N_1845,N_7679);
and U16260 (N_16260,N_2181,N_3963);
and U16261 (N_16261,N_2264,N_6372);
or U16262 (N_16262,N_4793,N_1522);
xor U16263 (N_16263,N_9221,N_6432);
nand U16264 (N_16264,N_565,N_3718);
nand U16265 (N_16265,N_5602,N_6577);
and U16266 (N_16266,N_9198,N_5044);
nor U16267 (N_16267,N_7164,N_9768);
nor U16268 (N_16268,N_4101,N_5583);
or U16269 (N_16269,N_1794,N_6576);
nor U16270 (N_16270,N_5232,N_7732);
or U16271 (N_16271,N_5164,N_9927);
and U16272 (N_16272,N_8291,N_7415);
nand U16273 (N_16273,N_3286,N_1210);
or U16274 (N_16274,N_8482,N_6920);
or U16275 (N_16275,N_5693,N_2501);
nor U16276 (N_16276,N_6162,N_2605);
nor U16277 (N_16277,N_8685,N_5701);
nand U16278 (N_16278,N_3285,N_5447);
or U16279 (N_16279,N_535,N_7415);
nand U16280 (N_16280,N_9448,N_1131);
nor U16281 (N_16281,N_2478,N_6245);
nand U16282 (N_16282,N_9435,N_5487);
nor U16283 (N_16283,N_9628,N_6168);
and U16284 (N_16284,N_9790,N_437);
and U16285 (N_16285,N_4891,N_8219);
or U16286 (N_16286,N_8878,N_4986);
and U16287 (N_16287,N_8922,N_8437);
nand U16288 (N_16288,N_6661,N_9250);
and U16289 (N_16289,N_2643,N_3015);
and U16290 (N_16290,N_47,N_6588);
nand U16291 (N_16291,N_6556,N_9528);
or U16292 (N_16292,N_5880,N_6568);
or U16293 (N_16293,N_8608,N_7748);
or U16294 (N_16294,N_9384,N_5963);
and U16295 (N_16295,N_4053,N_2063);
nor U16296 (N_16296,N_6733,N_3976);
nor U16297 (N_16297,N_3938,N_5662);
nor U16298 (N_16298,N_769,N_6002);
or U16299 (N_16299,N_8513,N_3874);
nand U16300 (N_16300,N_5779,N_6527);
and U16301 (N_16301,N_1615,N_420);
and U16302 (N_16302,N_4917,N_6305);
or U16303 (N_16303,N_8544,N_3461);
nor U16304 (N_16304,N_969,N_857);
or U16305 (N_16305,N_49,N_484);
or U16306 (N_16306,N_4255,N_1965);
nand U16307 (N_16307,N_2742,N_4345);
nor U16308 (N_16308,N_6939,N_3355);
and U16309 (N_16309,N_5793,N_9669);
nand U16310 (N_16310,N_3914,N_671);
nor U16311 (N_16311,N_3747,N_9353);
nor U16312 (N_16312,N_576,N_4016);
nor U16313 (N_16313,N_8404,N_3220);
nor U16314 (N_16314,N_4632,N_650);
or U16315 (N_16315,N_3727,N_5007);
nand U16316 (N_16316,N_5083,N_4034);
or U16317 (N_16317,N_8962,N_4314);
nand U16318 (N_16318,N_7452,N_6650);
or U16319 (N_16319,N_2894,N_1740);
and U16320 (N_16320,N_4741,N_7756);
and U16321 (N_16321,N_8008,N_4120);
or U16322 (N_16322,N_1168,N_663);
or U16323 (N_16323,N_1338,N_8836);
and U16324 (N_16324,N_882,N_2839);
and U16325 (N_16325,N_7399,N_2500);
nand U16326 (N_16326,N_15,N_3350);
nor U16327 (N_16327,N_6436,N_1813);
nand U16328 (N_16328,N_9384,N_5947);
or U16329 (N_16329,N_2967,N_9917);
nand U16330 (N_16330,N_7979,N_3521);
and U16331 (N_16331,N_8334,N_4726);
or U16332 (N_16332,N_7992,N_9116);
or U16333 (N_16333,N_5126,N_3108);
nor U16334 (N_16334,N_62,N_2559);
nor U16335 (N_16335,N_5379,N_8895);
and U16336 (N_16336,N_7823,N_1179);
or U16337 (N_16337,N_8401,N_8927);
nand U16338 (N_16338,N_5665,N_998);
and U16339 (N_16339,N_1885,N_6965);
and U16340 (N_16340,N_9576,N_7174);
or U16341 (N_16341,N_5266,N_7237);
nor U16342 (N_16342,N_3604,N_499);
and U16343 (N_16343,N_1987,N_7629);
nand U16344 (N_16344,N_2668,N_8601);
and U16345 (N_16345,N_820,N_806);
or U16346 (N_16346,N_8625,N_3047);
or U16347 (N_16347,N_4699,N_8685);
and U16348 (N_16348,N_7576,N_6350);
and U16349 (N_16349,N_172,N_8253);
or U16350 (N_16350,N_4377,N_5895);
nand U16351 (N_16351,N_9589,N_5269);
nor U16352 (N_16352,N_964,N_3089);
and U16353 (N_16353,N_1496,N_5362);
or U16354 (N_16354,N_8458,N_8139);
or U16355 (N_16355,N_4612,N_7242);
or U16356 (N_16356,N_6990,N_9754);
and U16357 (N_16357,N_2283,N_5113);
or U16358 (N_16358,N_4120,N_9190);
and U16359 (N_16359,N_861,N_1661);
nor U16360 (N_16360,N_7998,N_2585);
nor U16361 (N_16361,N_6121,N_9777);
nor U16362 (N_16362,N_9699,N_3940);
and U16363 (N_16363,N_2923,N_5295);
nor U16364 (N_16364,N_1372,N_3873);
nor U16365 (N_16365,N_5408,N_1778);
nor U16366 (N_16366,N_1601,N_6757);
and U16367 (N_16367,N_2039,N_6567);
nand U16368 (N_16368,N_3585,N_2718);
or U16369 (N_16369,N_9565,N_2267);
or U16370 (N_16370,N_277,N_7000);
and U16371 (N_16371,N_3639,N_7896);
nand U16372 (N_16372,N_6845,N_5341);
nor U16373 (N_16373,N_5139,N_2566);
nor U16374 (N_16374,N_723,N_3379);
nand U16375 (N_16375,N_3428,N_8070);
xor U16376 (N_16376,N_7903,N_2035);
or U16377 (N_16377,N_4386,N_4832);
nand U16378 (N_16378,N_5817,N_1974);
nand U16379 (N_16379,N_5063,N_9440);
and U16380 (N_16380,N_3995,N_8517);
and U16381 (N_16381,N_888,N_1262);
nor U16382 (N_16382,N_1669,N_2704);
and U16383 (N_16383,N_2976,N_3359);
and U16384 (N_16384,N_485,N_5406);
and U16385 (N_16385,N_7612,N_867);
and U16386 (N_16386,N_1544,N_1886);
nor U16387 (N_16387,N_8678,N_158);
or U16388 (N_16388,N_4729,N_5959);
or U16389 (N_16389,N_6345,N_5232);
and U16390 (N_16390,N_6992,N_1461);
nor U16391 (N_16391,N_7748,N_7411);
nor U16392 (N_16392,N_7273,N_2212);
and U16393 (N_16393,N_7835,N_347);
or U16394 (N_16394,N_7431,N_1119);
nand U16395 (N_16395,N_6619,N_7646);
nor U16396 (N_16396,N_7620,N_4083);
and U16397 (N_16397,N_2830,N_2077);
xor U16398 (N_16398,N_4779,N_6121);
and U16399 (N_16399,N_7042,N_6983);
nand U16400 (N_16400,N_9824,N_7698);
nand U16401 (N_16401,N_7492,N_8329);
nand U16402 (N_16402,N_8606,N_6238);
xnor U16403 (N_16403,N_146,N_5931);
and U16404 (N_16404,N_8446,N_3335);
nand U16405 (N_16405,N_5034,N_6465);
nand U16406 (N_16406,N_1019,N_4961);
nor U16407 (N_16407,N_3535,N_4468);
nand U16408 (N_16408,N_8875,N_4751);
or U16409 (N_16409,N_5476,N_920);
nor U16410 (N_16410,N_1805,N_9140);
nand U16411 (N_16411,N_1484,N_6957);
nor U16412 (N_16412,N_1944,N_8553);
and U16413 (N_16413,N_1077,N_123);
nor U16414 (N_16414,N_9162,N_2172);
and U16415 (N_16415,N_8903,N_8315);
nor U16416 (N_16416,N_2904,N_8597);
or U16417 (N_16417,N_4447,N_7778);
and U16418 (N_16418,N_6979,N_803);
nand U16419 (N_16419,N_8998,N_8914);
or U16420 (N_16420,N_7981,N_1580);
and U16421 (N_16421,N_8659,N_8986);
nand U16422 (N_16422,N_8843,N_3760);
nor U16423 (N_16423,N_3749,N_9709);
nand U16424 (N_16424,N_1848,N_7405);
and U16425 (N_16425,N_1868,N_7857);
or U16426 (N_16426,N_4639,N_3607);
or U16427 (N_16427,N_8282,N_3559);
or U16428 (N_16428,N_6981,N_9166);
and U16429 (N_16429,N_7346,N_3382);
nor U16430 (N_16430,N_8530,N_2073);
nand U16431 (N_16431,N_9943,N_6053);
nor U16432 (N_16432,N_3563,N_7328);
and U16433 (N_16433,N_7855,N_2128);
nor U16434 (N_16434,N_7870,N_2973);
nand U16435 (N_16435,N_1844,N_354);
or U16436 (N_16436,N_8041,N_7071);
or U16437 (N_16437,N_6662,N_8606);
nor U16438 (N_16438,N_1661,N_1577);
and U16439 (N_16439,N_4429,N_6526);
nor U16440 (N_16440,N_4027,N_9864);
nand U16441 (N_16441,N_7857,N_7016);
nor U16442 (N_16442,N_5656,N_9465);
or U16443 (N_16443,N_8531,N_1947);
nand U16444 (N_16444,N_2444,N_8800);
nand U16445 (N_16445,N_2344,N_3843);
nor U16446 (N_16446,N_3537,N_8684);
or U16447 (N_16447,N_4497,N_1084);
nand U16448 (N_16448,N_4176,N_3261);
or U16449 (N_16449,N_5981,N_8598);
nor U16450 (N_16450,N_2919,N_3475);
nand U16451 (N_16451,N_7821,N_6096);
xnor U16452 (N_16452,N_8669,N_7008);
and U16453 (N_16453,N_4318,N_7343);
and U16454 (N_16454,N_7852,N_3090);
and U16455 (N_16455,N_3412,N_3682);
or U16456 (N_16456,N_2696,N_2653);
and U16457 (N_16457,N_4018,N_6440);
or U16458 (N_16458,N_8655,N_9614);
nand U16459 (N_16459,N_443,N_9719);
or U16460 (N_16460,N_3675,N_5065);
and U16461 (N_16461,N_30,N_9117);
nand U16462 (N_16462,N_1554,N_6997);
nand U16463 (N_16463,N_6358,N_6649);
xor U16464 (N_16464,N_2647,N_1922);
and U16465 (N_16465,N_9832,N_7611);
nor U16466 (N_16466,N_3667,N_2428);
and U16467 (N_16467,N_149,N_795);
nor U16468 (N_16468,N_3599,N_9829);
nor U16469 (N_16469,N_2996,N_7650);
and U16470 (N_16470,N_3168,N_7075);
nand U16471 (N_16471,N_3428,N_6758);
nor U16472 (N_16472,N_4041,N_8779);
and U16473 (N_16473,N_4817,N_6127);
and U16474 (N_16474,N_822,N_4586);
nand U16475 (N_16475,N_3822,N_7784);
nand U16476 (N_16476,N_3831,N_3132);
nor U16477 (N_16477,N_2045,N_4777);
nand U16478 (N_16478,N_2189,N_2085);
and U16479 (N_16479,N_4008,N_5546);
or U16480 (N_16480,N_3618,N_9142);
nand U16481 (N_16481,N_6507,N_6641);
nor U16482 (N_16482,N_7582,N_5625);
or U16483 (N_16483,N_7,N_9281);
nor U16484 (N_16484,N_6466,N_7001);
nor U16485 (N_16485,N_9951,N_5596);
nand U16486 (N_16486,N_9557,N_3484);
nor U16487 (N_16487,N_5751,N_1248);
or U16488 (N_16488,N_7878,N_4429);
or U16489 (N_16489,N_9918,N_9803);
and U16490 (N_16490,N_7276,N_3685);
and U16491 (N_16491,N_3710,N_831);
nor U16492 (N_16492,N_7294,N_5725);
or U16493 (N_16493,N_6790,N_8675);
nand U16494 (N_16494,N_6628,N_9659);
nor U16495 (N_16495,N_2627,N_9594);
nand U16496 (N_16496,N_8757,N_5762);
nand U16497 (N_16497,N_5421,N_3017);
and U16498 (N_16498,N_9527,N_8552);
nor U16499 (N_16499,N_2778,N_3317);
and U16500 (N_16500,N_4255,N_2889);
nor U16501 (N_16501,N_6275,N_145);
or U16502 (N_16502,N_5391,N_9307);
or U16503 (N_16503,N_6938,N_4511);
or U16504 (N_16504,N_4695,N_4147);
and U16505 (N_16505,N_7355,N_3000);
nor U16506 (N_16506,N_369,N_8135);
nand U16507 (N_16507,N_102,N_1751);
nor U16508 (N_16508,N_3757,N_9403);
nor U16509 (N_16509,N_9551,N_9339);
nand U16510 (N_16510,N_1520,N_9897);
nand U16511 (N_16511,N_9169,N_2189);
and U16512 (N_16512,N_6998,N_9180);
or U16513 (N_16513,N_8020,N_6664);
or U16514 (N_16514,N_5067,N_9336);
and U16515 (N_16515,N_1981,N_1399);
or U16516 (N_16516,N_3149,N_3161);
and U16517 (N_16517,N_308,N_4928);
or U16518 (N_16518,N_5295,N_3717);
nor U16519 (N_16519,N_8538,N_6958);
nand U16520 (N_16520,N_3722,N_2007);
or U16521 (N_16521,N_2634,N_1689);
nand U16522 (N_16522,N_1269,N_4240);
nor U16523 (N_16523,N_4729,N_5488);
and U16524 (N_16524,N_666,N_5979);
or U16525 (N_16525,N_7139,N_65);
nand U16526 (N_16526,N_2725,N_5143);
and U16527 (N_16527,N_7507,N_603);
nor U16528 (N_16528,N_3497,N_1796);
and U16529 (N_16529,N_6718,N_9132);
nor U16530 (N_16530,N_562,N_2202);
and U16531 (N_16531,N_7810,N_8276);
and U16532 (N_16532,N_1082,N_9807);
nor U16533 (N_16533,N_8808,N_137);
nor U16534 (N_16534,N_456,N_7879);
and U16535 (N_16535,N_3762,N_6671);
or U16536 (N_16536,N_7309,N_2227);
and U16537 (N_16537,N_7735,N_5616);
nor U16538 (N_16538,N_4573,N_6825);
nor U16539 (N_16539,N_7890,N_6530);
nor U16540 (N_16540,N_4100,N_1669);
nand U16541 (N_16541,N_6968,N_856);
nor U16542 (N_16542,N_9737,N_5767);
nand U16543 (N_16543,N_946,N_667);
nand U16544 (N_16544,N_680,N_3024);
or U16545 (N_16545,N_8683,N_7383);
nand U16546 (N_16546,N_7508,N_8796);
or U16547 (N_16547,N_7955,N_6408);
nor U16548 (N_16548,N_6308,N_1089);
nor U16549 (N_16549,N_9146,N_1299);
nand U16550 (N_16550,N_7120,N_6272);
nand U16551 (N_16551,N_6060,N_8522);
and U16552 (N_16552,N_864,N_7598);
nand U16553 (N_16553,N_3605,N_8124);
and U16554 (N_16554,N_8951,N_922);
nand U16555 (N_16555,N_7393,N_1988);
or U16556 (N_16556,N_7022,N_3476);
nor U16557 (N_16557,N_8762,N_8674);
nor U16558 (N_16558,N_2179,N_1715);
nor U16559 (N_16559,N_6301,N_2397);
nor U16560 (N_16560,N_3186,N_146);
and U16561 (N_16561,N_2658,N_7963);
nor U16562 (N_16562,N_8774,N_7112);
nor U16563 (N_16563,N_3730,N_8109);
nand U16564 (N_16564,N_9219,N_6666);
nand U16565 (N_16565,N_1757,N_2911);
nand U16566 (N_16566,N_7083,N_8796);
and U16567 (N_16567,N_1578,N_6982);
nor U16568 (N_16568,N_7768,N_1069);
nand U16569 (N_16569,N_4740,N_1785);
and U16570 (N_16570,N_4292,N_24);
nand U16571 (N_16571,N_7647,N_8240);
nor U16572 (N_16572,N_5542,N_5744);
nor U16573 (N_16573,N_8962,N_2709);
and U16574 (N_16574,N_1469,N_2069);
or U16575 (N_16575,N_6480,N_4217);
nand U16576 (N_16576,N_9104,N_6165);
or U16577 (N_16577,N_9106,N_7625);
nor U16578 (N_16578,N_877,N_2457);
or U16579 (N_16579,N_4517,N_9774);
and U16580 (N_16580,N_6173,N_832);
or U16581 (N_16581,N_3227,N_7428);
or U16582 (N_16582,N_4294,N_4895);
and U16583 (N_16583,N_4104,N_4809);
nor U16584 (N_16584,N_4750,N_752);
nor U16585 (N_16585,N_2156,N_9697);
nor U16586 (N_16586,N_6439,N_5521);
nand U16587 (N_16587,N_5467,N_7475);
or U16588 (N_16588,N_3015,N_446);
or U16589 (N_16589,N_6043,N_3639);
and U16590 (N_16590,N_7526,N_4781);
nor U16591 (N_16591,N_6141,N_4910);
and U16592 (N_16592,N_3879,N_3256);
and U16593 (N_16593,N_9790,N_2583);
nand U16594 (N_16594,N_1379,N_5216);
nand U16595 (N_16595,N_864,N_8094);
or U16596 (N_16596,N_2169,N_3940);
or U16597 (N_16597,N_5448,N_2946);
nor U16598 (N_16598,N_1194,N_5161);
nand U16599 (N_16599,N_5391,N_2702);
or U16600 (N_16600,N_1020,N_3086);
and U16601 (N_16601,N_4445,N_406);
nor U16602 (N_16602,N_9568,N_7140);
and U16603 (N_16603,N_7394,N_745);
or U16604 (N_16604,N_9027,N_3733);
and U16605 (N_16605,N_6905,N_8930);
nand U16606 (N_16606,N_8772,N_7828);
nand U16607 (N_16607,N_2974,N_7137);
nand U16608 (N_16608,N_1405,N_33);
and U16609 (N_16609,N_8241,N_3137);
nand U16610 (N_16610,N_6228,N_8722);
nand U16611 (N_16611,N_1765,N_3946);
and U16612 (N_16612,N_3348,N_3182);
nand U16613 (N_16613,N_5173,N_7900);
nand U16614 (N_16614,N_8604,N_881);
or U16615 (N_16615,N_2844,N_7862);
or U16616 (N_16616,N_4131,N_2360);
and U16617 (N_16617,N_1607,N_1139);
nor U16618 (N_16618,N_1044,N_9893);
and U16619 (N_16619,N_7632,N_9933);
nor U16620 (N_16620,N_5176,N_5521);
nand U16621 (N_16621,N_3758,N_1029);
or U16622 (N_16622,N_5287,N_651);
or U16623 (N_16623,N_199,N_4236);
nand U16624 (N_16624,N_7263,N_5679);
nor U16625 (N_16625,N_2742,N_6463);
and U16626 (N_16626,N_96,N_1713);
or U16627 (N_16627,N_9135,N_633);
nand U16628 (N_16628,N_1954,N_2308);
or U16629 (N_16629,N_4359,N_7372);
nand U16630 (N_16630,N_9256,N_2569);
or U16631 (N_16631,N_3918,N_2055);
or U16632 (N_16632,N_1621,N_1780);
and U16633 (N_16633,N_5983,N_1872);
nor U16634 (N_16634,N_7451,N_9124);
and U16635 (N_16635,N_8875,N_6139);
nor U16636 (N_16636,N_3640,N_8294);
and U16637 (N_16637,N_8511,N_7201);
or U16638 (N_16638,N_8479,N_1647);
nor U16639 (N_16639,N_9990,N_9873);
nor U16640 (N_16640,N_4158,N_6377);
and U16641 (N_16641,N_4792,N_6579);
and U16642 (N_16642,N_9853,N_6077);
nor U16643 (N_16643,N_8174,N_9378);
and U16644 (N_16644,N_1836,N_4356);
and U16645 (N_16645,N_3056,N_182);
nor U16646 (N_16646,N_3937,N_8044);
nand U16647 (N_16647,N_5362,N_4899);
or U16648 (N_16648,N_927,N_7076);
nor U16649 (N_16649,N_309,N_1421);
and U16650 (N_16650,N_6257,N_4602);
or U16651 (N_16651,N_424,N_4460);
nand U16652 (N_16652,N_4111,N_3803);
and U16653 (N_16653,N_5682,N_4290);
nand U16654 (N_16654,N_7140,N_2256);
or U16655 (N_16655,N_9013,N_2578);
or U16656 (N_16656,N_6426,N_7754);
nand U16657 (N_16657,N_6321,N_8140);
nand U16658 (N_16658,N_6308,N_4233);
or U16659 (N_16659,N_639,N_5805);
or U16660 (N_16660,N_6196,N_4106);
nand U16661 (N_16661,N_3921,N_6586);
or U16662 (N_16662,N_7955,N_2840);
and U16663 (N_16663,N_7520,N_9071);
or U16664 (N_16664,N_168,N_3214);
nor U16665 (N_16665,N_3732,N_4641);
nor U16666 (N_16666,N_7623,N_6553);
and U16667 (N_16667,N_5323,N_3767);
or U16668 (N_16668,N_4465,N_7206);
and U16669 (N_16669,N_9739,N_1758);
or U16670 (N_16670,N_6569,N_6231);
and U16671 (N_16671,N_9509,N_8065);
nand U16672 (N_16672,N_9820,N_8035);
nor U16673 (N_16673,N_7092,N_4867);
and U16674 (N_16674,N_1584,N_1821);
or U16675 (N_16675,N_2298,N_1487);
nand U16676 (N_16676,N_1150,N_3456);
nor U16677 (N_16677,N_7043,N_4419);
or U16678 (N_16678,N_4359,N_6834);
nor U16679 (N_16679,N_1756,N_4613);
and U16680 (N_16680,N_6607,N_3287);
or U16681 (N_16681,N_5566,N_1485);
or U16682 (N_16682,N_174,N_5908);
xnor U16683 (N_16683,N_6430,N_8296);
and U16684 (N_16684,N_9756,N_575);
nor U16685 (N_16685,N_3527,N_6676);
nor U16686 (N_16686,N_8581,N_8028);
nand U16687 (N_16687,N_7936,N_8397);
or U16688 (N_16688,N_1876,N_3420);
or U16689 (N_16689,N_3974,N_6053);
or U16690 (N_16690,N_7944,N_9122);
nor U16691 (N_16691,N_94,N_8037);
and U16692 (N_16692,N_9613,N_3611);
nand U16693 (N_16693,N_5401,N_8755);
nor U16694 (N_16694,N_3041,N_482);
nand U16695 (N_16695,N_9456,N_7187);
nand U16696 (N_16696,N_2347,N_1189);
and U16697 (N_16697,N_6390,N_188);
or U16698 (N_16698,N_62,N_7810);
nand U16699 (N_16699,N_9651,N_4551);
and U16700 (N_16700,N_7976,N_2742);
or U16701 (N_16701,N_4389,N_9491);
nor U16702 (N_16702,N_9325,N_5797);
nor U16703 (N_16703,N_2634,N_7151);
and U16704 (N_16704,N_3371,N_375);
nand U16705 (N_16705,N_2954,N_6631);
or U16706 (N_16706,N_6428,N_8234);
nand U16707 (N_16707,N_9129,N_1031);
or U16708 (N_16708,N_5672,N_1602);
and U16709 (N_16709,N_5485,N_2300);
nand U16710 (N_16710,N_7934,N_4327);
or U16711 (N_16711,N_5235,N_3138);
and U16712 (N_16712,N_5496,N_9324);
nand U16713 (N_16713,N_3881,N_9815);
nand U16714 (N_16714,N_7902,N_8868);
and U16715 (N_16715,N_2817,N_8763);
nand U16716 (N_16716,N_5690,N_4219);
or U16717 (N_16717,N_6127,N_5571);
nor U16718 (N_16718,N_405,N_4443);
or U16719 (N_16719,N_3857,N_7589);
or U16720 (N_16720,N_368,N_7881);
nor U16721 (N_16721,N_7668,N_2770);
and U16722 (N_16722,N_9004,N_2803);
nor U16723 (N_16723,N_8241,N_3507);
and U16724 (N_16724,N_3934,N_2400);
or U16725 (N_16725,N_2210,N_1853);
nor U16726 (N_16726,N_9164,N_9031);
and U16727 (N_16727,N_4244,N_1856);
nor U16728 (N_16728,N_8012,N_7962);
nor U16729 (N_16729,N_9869,N_9334);
and U16730 (N_16730,N_9234,N_791);
nor U16731 (N_16731,N_2381,N_4449);
nor U16732 (N_16732,N_8110,N_6974);
and U16733 (N_16733,N_8180,N_7979);
nor U16734 (N_16734,N_4524,N_5145);
nand U16735 (N_16735,N_4352,N_7893);
nand U16736 (N_16736,N_1621,N_694);
nand U16737 (N_16737,N_5535,N_4323);
or U16738 (N_16738,N_8419,N_9840);
and U16739 (N_16739,N_1226,N_2037);
and U16740 (N_16740,N_3598,N_5873);
and U16741 (N_16741,N_6967,N_5723);
or U16742 (N_16742,N_5746,N_3137);
nand U16743 (N_16743,N_5826,N_8257);
nand U16744 (N_16744,N_4932,N_5713);
nand U16745 (N_16745,N_2011,N_1618);
nand U16746 (N_16746,N_4948,N_8911);
nand U16747 (N_16747,N_6622,N_3602);
and U16748 (N_16748,N_6690,N_7676);
nor U16749 (N_16749,N_7917,N_1970);
nor U16750 (N_16750,N_7677,N_1470);
nand U16751 (N_16751,N_1762,N_2714);
and U16752 (N_16752,N_2105,N_5775);
or U16753 (N_16753,N_9497,N_8703);
and U16754 (N_16754,N_4529,N_4394);
or U16755 (N_16755,N_9875,N_872);
and U16756 (N_16756,N_5008,N_2305);
or U16757 (N_16757,N_7003,N_3944);
nor U16758 (N_16758,N_8047,N_6475);
or U16759 (N_16759,N_9721,N_7758);
nor U16760 (N_16760,N_996,N_9510);
nand U16761 (N_16761,N_9322,N_9789);
xnor U16762 (N_16762,N_6741,N_8461);
or U16763 (N_16763,N_3559,N_9584);
and U16764 (N_16764,N_6305,N_3741);
nor U16765 (N_16765,N_1419,N_5228);
or U16766 (N_16766,N_4025,N_372);
nor U16767 (N_16767,N_8751,N_7690);
or U16768 (N_16768,N_2496,N_548);
and U16769 (N_16769,N_8486,N_3011);
nand U16770 (N_16770,N_7462,N_8310);
and U16771 (N_16771,N_500,N_1541);
nor U16772 (N_16772,N_9682,N_6793);
and U16773 (N_16773,N_2968,N_1031);
nor U16774 (N_16774,N_3781,N_8566);
nor U16775 (N_16775,N_7858,N_2742);
nand U16776 (N_16776,N_7523,N_8097);
nor U16777 (N_16777,N_9157,N_6826);
and U16778 (N_16778,N_691,N_4137);
nor U16779 (N_16779,N_6178,N_1634);
nor U16780 (N_16780,N_6720,N_3830);
or U16781 (N_16781,N_4824,N_8124);
or U16782 (N_16782,N_6723,N_5462);
nand U16783 (N_16783,N_1281,N_6176);
and U16784 (N_16784,N_5418,N_7105);
or U16785 (N_16785,N_5645,N_4432);
or U16786 (N_16786,N_8158,N_1385);
nor U16787 (N_16787,N_2585,N_1875);
and U16788 (N_16788,N_5830,N_6778);
nor U16789 (N_16789,N_283,N_9278);
or U16790 (N_16790,N_6726,N_6343);
and U16791 (N_16791,N_8489,N_7441);
nor U16792 (N_16792,N_4687,N_8526);
nor U16793 (N_16793,N_7309,N_804);
nor U16794 (N_16794,N_7293,N_6492);
and U16795 (N_16795,N_5996,N_6770);
and U16796 (N_16796,N_5547,N_6330);
nand U16797 (N_16797,N_7221,N_1964);
and U16798 (N_16798,N_6160,N_5622);
nor U16799 (N_16799,N_986,N_6917);
nor U16800 (N_16800,N_3301,N_6703);
nand U16801 (N_16801,N_1939,N_4191);
nor U16802 (N_16802,N_9322,N_8783);
nor U16803 (N_16803,N_1780,N_5743);
nor U16804 (N_16804,N_2772,N_6497);
nor U16805 (N_16805,N_9509,N_9445);
nand U16806 (N_16806,N_3212,N_4697);
nor U16807 (N_16807,N_5528,N_2172);
or U16808 (N_16808,N_7130,N_7935);
nand U16809 (N_16809,N_1662,N_7448);
nand U16810 (N_16810,N_7851,N_2247);
or U16811 (N_16811,N_842,N_4542);
and U16812 (N_16812,N_2341,N_6901);
and U16813 (N_16813,N_5875,N_9376);
and U16814 (N_16814,N_3495,N_4733);
and U16815 (N_16815,N_5796,N_2187);
nand U16816 (N_16816,N_4511,N_4549);
nand U16817 (N_16817,N_5942,N_8815);
nor U16818 (N_16818,N_6648,N_6228);
nand U16819 (N_16819,N_7953,N_483);
nor U16820 (N_16820,N_3870,N_5242);
nor U16821 (N_16821,N_7933,N_7627);
and U16822 (N_16822,N_8159,N_6471);
nand U16823 (N_16823,N_7312,N_7048);
and U16824 (N_16824,N_7691,N_7235);
xor U16825 (N_16825,N_6324,N_4057);
and U16826 (N_16826,N_2906,N_9711);
nor U16827 (N_16827,N_1229,N_3299);
and U16828 (N_16828,N_6290,N_5523);
nand U16829 (N_16829,N_7085,N_7201);
nor U16830 (N_16830,N_2902,N_851);
nand U16831 (N_16831,N_570,N_6723);
nor U16832 (N_16832,N_1459,N_2628);
nor U16833 (N_16833,N_318,N_9692);
nor U16834 (N_16834,N_8843,N_8011);
nand U16835 (N_16835,N_217,N_9910);
nand U16836 (N_16836,N_7754,N_4591);
nor U16837 (N_16837,N_4962,N_401);
and U16838 (N_16838,N_2096,N_5869);
and U16839 (N_16839,N_5016,N_2159);
and U16840 (N_16840,N_9969,N_3364);
nand U16841 (N_16841,N_703,N_7450);
and U16842 (N_16842,N_4,N_7791);
nor U16843 (N_16843,N_4984,N_6768);
nor U16844 (N_16844,N_5678,N_1763);
nor U16845 (N_16845,N_8654,N_4305);
or U16846 (N_16846,N_3936,N_3487);
nor U16847 (N_16847,N_6250,N_1003);
nand U16848 (N_16848,N_3065,N_6582);
nor U16849 (N_16849,N_3593,N_4793);
or U16850 (N_16850,N_8101,N_46);
nor U16851 (N_16851,N_3487,N_8697);
nor U16852 (N_16852,N_2254,N_5783);
nor U16853 (N_16853,N_4590,N_1244);
nand U16854 (N_16854,N_7713,N_8386);
nand U16855 (N_16855,N_3510,N_3);
or U16856 (N_16856,N_1725,N_6248);
or U16857 (N_16857,N_5515,N_7014);
or U16858 (N_16858,N_2373,N_2317);
nor U16859 (N_16859,N_7314,N_6884);
nand U16860 (N_16860,N_3073,N_6868);
nor U16861 (N_16861,N_7926,N_319);
or U16862 (N_16862,N_1933,N_5612);
nor U16863 (N_16863,N_1074,N_7908);
nor U16864 (N_16864,N_9363,N_9524);
or U16865 (N_16865,N_6071,N_9476);
and U16866 (N_16866,N_9226,N_7296);
and U16867 (N_16867,N_1419,N_2013);
and U16868 (N_16868,N_8366,N_9412);
or U16869 (N_16869,N_5042,N_3925);
and U16870 (N_16870,N_2478,N_5726);
nand U16871 (N_16871,N_6930,N_6811);
and U16872 (N_16872,N_3239,N_2463);
and U16873 (N_16873,N_1365,N_4669);
and U16874 (N_16874,N_8952,N_3421);
nand U16875 (N_16875,N_3891,N_5382);
nand U16876 (N_16876,N_2685,N_3777);
or U16877 (N_16877,N_5464,N_159);
nor U16878 (N_16878,N_2885,N_6982);
nor U16879 (N_16879,N_3266,N_5200);
and U16880 (N_16880,N_8953,N_6793);
nand U16881 (N_16881,N_5228,N_2351);
nand U16882 (N_16882,N_5131,N_5624);
nand U16883 (N_16883,N_4620,N_8820);
and U16884 (N_16884,N_445,N_9221);
nor U16885 (N_16885,N_3821,N_9422);
nor U16886 (N_16886,N_1,N_5973);
nand U16887 (N_16887,N_3539,N_7693);
or U16888 (N_16888,N_648,N_8169);
nor U16889 (N_16889,N_5465,N_524);
nand U16890 (N_16890,N_932,N_4509);
nand U16891 (N_16891,N_6392,N_2871);
and U16892 (N_16892,N_6561,N_8032);
nor U16893 (N_16893,N_6542,N_3170);
or U16894 (N_16894,N_8405,N_3141);
nand U16895 (N_16895,N_1278,N_6586);
nor U16896 (N_16896,N_6107,N_311);
nor U16897 (N_16897,N_5151,N_297);
and U16898 (N_16898,N_6117,N_6422);
nand U16899 (N_16899,N_6540,N_8468);
and U16900 (N_16900,N_1365,N_4788);
nand U16901 (N_16901,N_5619,N_3780);
or U16902 (N_16902,N_5516,N_1274);
or U16903 (N_16903,N_4338,N_3099);
and U16904 (N_16904,N_3198,N_7432);
or U16905 (N_16905,N_4202,N_5918);
and U16906 (N_16906,N_292,N_4197);
nor U16907 (N_16907,N_4360,N_1245);
or U16908 (N_16908,N_6170,N_9511);
nand U16909 (N_16909,N_6116,N_292);
nor U16910 (N_16910,N_436,N_7268);
or U16911 (N_16911,N_7139,N_3804);
nand U16912 (N_16912,N_1797,N_1589);
nor U16913 (N_16913,N_3847,N_9249);
and U16914 (N_16914,N_9480,N_4404);
or U16915 (N_16915,N_9061,N_7739);
nand U16916 (N_16916,N_9697,N_5061);
nand U16917 (N_16917,N_6424,N_7367);
nand U16918 (N_16918,N_2024,N_8883);
nor U16919 (N_16919,N_449,N_2135);
or U16920 (N_16920,N_2477,N_1899);
or U16921 (N_16921,N_6621,N_1722);
and U16922 (N_16922,N_1753,N_7918);
nand U16923 (N_16923,N_4945,N_9812);
and U16924 (N_16924,N_8092,N_8402);
nor U16925 (N_16925,N_5207,N_683);
and U16926 (N_16926,N_4172,N_9033);
nor U16927 (N_16927,N_1919,N_8822);
or U16928 (N_16928,N_4401,N_765);
or U16929 (N_16929,N_3570,N_7063);
and U16930 (N_16930,N_600,N_3516);
nand U16931 (N_16931,N_4299,N_5903);
and U16932 (N_16932,N_7041,N_5105);
and U16933 (N_16933,N_5143,N_5868);
nor U16934 (N_16934,N_7571,N_4438);
nand U16935 (N_16935,N_5759,N_3411);
nand U16936 (N_16936,N_4624,N_6296);
nand U16937 (N_16937,N_6644,N_2211);
and U16938 (N_16938,N_1613,N_500);
nor U16939 (N_16939,N_727,N_723);
and U16940 (N_16940,N_897,N_834);
and U16941 (N_16941,N_4823,N_7123);
nand U16942 (N_16942,N_1157,N_3251);
nor U16943 (N_16943,N_4849,N_1930);
and U16944 (N_16944,N_3095,N_7216);
nor U16945 (N_16945,N_3805,N_304);
and U16946 (N_16946,N_2960,N_2046);
nor U16947 (N_16947,N_2680,N_8360);
or U16948 (N_16948,N_1204,N_7130);
nand U16949 (N_16949,N_9342,N_773);
or U16950 (N_16950,N_6913,N_9778);
or U16951 (N_16951,N_1965,N_5770);
or U16952 (N_16952,N_4545,N_3953);
nand U16953 (N_16953,N_2790,N_3909);
nor U16954 (N_16954,N_2449,N_4738);
nand U16955 (N_16955,N_2491,N_278);
nor U16956 (N_16956,N_5650,N_9094);
nor U16957 (N_16957,N_8412,N_9763);
xnor U16958 (N_16958,N_2659,N_5274);
nor U16959 (N_16959,N_4378,N_3026);
nand U16960 (N_16960,N_6870,N_7493);
and U16961 (N_16961,N_3476,N_9466);
or U16962 (N_16962,N_7888,N_8611);
or U16963 (N_16963,N_8876,N_2741);
nand U16964 (N_16964,N_5656,N_8698);
nor U16965 (N_16965,N_8990,N_6326);
or U16966 (N_16966,N_1778,N_6691);
nand U16967 (N_16967,N_4994,N_9595);
nand U16968 (N_16968,N_2847,N_12);
nor U16969 (N_16969,N_4529,N_3810);
nor U16970 (N_16970,N_2102,N_2295);
nor U16971 (N_16971,N_4539,N_7378);
and U16972 (N_16972,N_4078,N_1222);
nand U16973 (N_16973,N_3272,N_4774);
nand U16974 (N_16974,N_525,N_8574);
and U16975 (N_16975,N_3948,N_9060);
nor U16976 (N_16976,N_5949,N_604);
nor U16977 (N_16977,N_2300,N_3845);
nor U16978 (N_16978,N_1102,N_1370);
nand U16979 (N_16979,N_5811,N_2578);
and U16980 (N_16980,N_6501,N_7859);
or U16981 (N_16981,N_2058,N_1121);
nand U16982 (N_16982,N_5848,N_103);
or U16983 (N_16983,N_7087,N_9894);
or U16984 (N_16984,N_7295,N_5391);
and U16985 (N_16985,N_5800,N_3259);
nor U16986 (N_16986,N_7461,N_2174);
or U16987 (N_16987,N_4893,N_6864);
and U16988 (N_16988,N_1041,N_9712);
or U16989 (N_16989,N_4828,N_574);
and U16990 (N_16990,N_9553,N_1314);
and U16991 (N_16991,N_8248,N_9446);
xnor U16992 (N_16992,N_5015,N_7072);
nand U16993 (N_16993,N_5217,N_533);
nand U16994 (N_16994,N_5470,N_2550);
nand U16995 (N_16995,N_2927,N_7633);
or U16996 (N_16996,N_4130,N_74);
or U16997 (N_16997,N_8829,N_5199);
or U16998 (N_16998,N_6328,N_7630);
nor U16999 (N_16999,N_4047,N_715);
nand U17000 (N_17000,N_9957,N_9265);
nor U17001 (N_17001,N_6027,N_2326);
nor U17002 (N_17002,N_897,N_2218);
or U17003 (N_17003,N_4352,N_6526);
and U17004 (N_17004,N_2394,N_5408);
nor U17005 (N_17005,N_5350,N_381);
or U17006 (N_17006,N_6282,N_1234);
and U17007 (N_17007,N_6202,N_4604);
or U17008 (N_17008,N_6550,N_7564);
nand U17009 (N_17009,N_1525,N_8247);
nor U17010 (N_17010,N_606,N_7884);
nor U17011 (N_17011,N_1243,N_6669);
nand U17012 (N_17012,N_5956,N_2295);
nand U17013 (N_17013,N_8079,N_6723);
and U17014 (N_17014,N_7231,N_8277);
and U17015 (N_17015,N_7971,N_2318);
nor U17016 (N_17016,N_8495,N_2826);
nand U17017 (N_17017,N_6729,N_2186);
and U17018 (N_17018,N_2960,N_6556);
nor U17019 (N_17019,N_4203,N_6113);
nand U17020 (N_17020,N_2621,N_6739);
nand U17021 (N_17021,N_9716,N_8607);
nor U17022 (N_17022,N_9479,N_3916);
nand U17023 (N_17023,N_9313,N_7408);
or U17024 (N_17024,N_197,N_5937);
nor U17025 (N_17025,N_5170,N_1152);
and U17026 (N_17026,N_3231,N_6750);
nor U17027 (N_17027,N_5541,N_8097);
or U17028 (N_17028,N_1755,N_1113);
or U17029 (N_17029,N_2484,N_7961);
nor U17030 (N_17030,N_8715,N_1693);
nor U17031 (N_17031,N_9817,N_5480);
or U17032 (N_17032,N_5005,N_9456);
nand U17033 (N_17033,N_4663,N_7608);
nor U17034 (N_17034,N_2375,N_2567);
or U17035 (N_17035,N_6281,N_3646);
and U17036 (N_17036,N_8097,N_8929);
and U17037 (N_17037,N_4917,N_1767);
nand U17038 (N_17038,N_3239,N_628);
and U17039 (N_17039,N_6048,N_2883);
nor U17040 (N_17040,N_8499,N_5159);
xnor U17041 (N_17041,N_9143,N_3894);
nand U17042 (N_17042,N_387,N_5408);
and U17043 (N_17043,N_2695,N_1571);
nand U17044 (N_17044,N_88,N_9593);
and U17045 (N_17045,N_7201,N_1051);
or U17046 (N_17046,N_5720,N_3865);
nor U17047 (N_17047,N_9599,N_3744);
and U17048 (N_17048,N_1500,N_3102);
and U17049 (N_17049,N_3790,N_6576);
nor U17050 (N_17050,N_1479,N_8016);
nor U17051 (N_17051,N_3478,N_7954);
nand U17052 (N_17052,N_6612,N_1070);
and U17053 (N_17053,N_2484,N_2321);
and U17054 (N_17054,N_1216,N_3562);
or U17055 (N_17055,N_4569,N_703);
nor U17056 (N_17056,N_9505,N_9719);
nor U17057 (N_17057,N_9051,N_1437);
nor U17058 (N_17058,N_6419,N_5168);
nand U17059 (N_17059,N_6800,N_9070);
xnor U17060 (N_17060,N_7720,N_3472);
nand U17061 (N_17061,N_8462,N_5274);
and U17062 (N_17062,N_4046,N_6544);
nand U17063 (N_17063,N_9395,N_1266);
and U17064 (N_17064,N_3059,N_7290);
or U17065 (N_17065,N_2513,N_8883);
nor U17066 (N_17066,N_7986,N_5451);
nand U17067 (N_17067,N_9112,N_5994);
or U17068 (N_17068,N_2983,N_7498);
or U17069 (N_17069,N_662,N_2997);
and U17070 (N_17070,N_8870,N_5107);
or U17071 (N_17071,N_369,N_3885);
xor U17072 (N_17072,N_3042,N_8351);
or U17073 (N_17073,N_4398,N_997);
nand U17074 (N_17074,N_7816,N_7935);
or U17075 (N_17075,N_365,N_5691);
and U17076 (N_17076,N_6146,N_3174);
or U17077 (N_17077,N_2255,N_1721);
nor U17078 (N_17078,N_8618,N_8383);
or U17079 (N_17079,N_9568,N_5522);
nand U17080 (N_17080,N_4991,N_6533);
or U17081 (N_17081,N_8921,N_3449);
or U17082 (N_17082,N_2142,N_7078);
nand U17083 (N_17083,N_1282,N_3820);
or U17084 (N_17084,N_2483,N_3072);
nand U17085 (N_17085,N_1955,N_468);
nand U17086 (N_17086,N_1561,N_3273);
and U17087 (N_17087,N_9610,N_8135);
nand U17088 (N_17088,N_504,N_3980);
and U17089 (N_17089,N_6078,N_4510);
nor U17090 (N_17090,N_2842,N_3918);
or U17091 (N_17091,N_4937,N_1797);
nor U17092 (N_17092,N_854,N_8019);
nor U17093 (N_17093,N_3902,N_1960);
and U17094 (N_17094,N_8661,N_4691);
and U17095 (N_17095,N_334,N_8736);
nand U17096 (N_17096,N_7417,N_5487);
or U17097 (N_17097,N_5630,N_8731);
and U17098 (N_17098,N_3005,N_3460);
nor U17099 (N_17099,N_5293,N_8250);
nor U17100 (N_17100,N_5392,N_2079);
nand U17101 (N_17101,N_8885,N_7018);
or U17102 (N_17102,N_8979,N_6494);
or U17103 (N_17103,N_1618,N_1651);
and U17104 (N_17104,N_5172,N_5072);
nor U17105 (N_17105,N_5144,N_6061);
and U17106 (N_17106,N_1123,N_1763);
and U17107 (N_17107,N_1740,N_7773);
or U17108 (N_17108,N_6555,N_4868);
nor U17109 (N_17109,N_2703,N_5510);
or U17110 (N_17110,N_2851,N_9009);
nor U17111 (N_17111,N_1460,N_5398);
xnor U17112 (N_17112,N_1529,N_2826);
nor U17113 (N_17113,N_7992,N_1294);
or U17114 (N_17114,N_142,N_4286);
or U17115 (N_17115,N_1677,N_6158);
nor U17116 (N_17116,N_7197,N_5137);
nand U17117 (N_17117,N_2149,N_2818);
nand U17118 (N_17118,N_1564,N_4692);
and U17119 (N_17119,N_7211,N_5235);
nand U17120 (N_17120,N_4172,N_8989);
or U17121 (N_17121,N_2874,N_1315);
nor U17122 (N_17122,N_8517,N_2515);
or U17123 (N_17123,N_3767,N_5815);
nor U17124 (N_17124,N_8010,N_7895);
nor U17125 (N_17125,N_5425,N_9837);
or U17126 (N_17126,N_2938,N_8327);
and U17127 (N_17127,N_2713,N_4879);
and U17128 (N_17128,N_9898,N_7700);
nand U17129 (N_17129,N_8846,N_6424);
nand U17130 (N_17130,N_1435,N_4888);
or U17131 (N_17131,N_3763,N_7094);
nor U17132 (N_17132,N_8038,N_6518);
or U17133 (N_17133,N_8358,N_9161);
nor U17134 (N_17134,N_58,N_7673);
nand U17135 (N_17135,N_8347,N_7529);
nor U17136 (N_17136,N_1573,N_6215);
and U17137 (N_17137,N_9373,N_4180);
nor U17138 (N_17138,N_7549,N_5823);
or U17139 (N_17139,N_6337,N_8283);
nand U17140 (N_17140,N_8368,N_6168);
nor U17141 (N_17141,N_3454,N_4435);
nand U17142 (N_17142,N_901,N_4290);
nor U17143 (N_17143,N_1979,N_6424);
nand U17144 (N_17144,N_7396,N_9030);
or U17145 (N_17145,N_5226,N_9393);
nor U17146 (N_17146,N_7683,N_3254);
nand U17147 (N_17147,N_416,N_479);
and U17148 (N_17148,N_8374,N_4442);
or U17149 (N_17149,N_7328,N_625);
nor U17150 (N_17150,N_5023,N_2398);
nor U17151 (N_17151,N_8018,N_1916);
and U17152 (N_17152,N_1556,N_1059);
or U17153 (N_17153,N_479,N_2988);
and U17154 (N_17154,N_6646,N_3526);
nand U17155 (N_17155,N_7439,N_5046);
nor U17156 (N_17156,N_9874,N_9009);
or U17157 (N_17157,N_2805,N_348);
or U17158 (N_17158,N_3934,N_3077);
nor U17159 (N_17159,N_2346,N_3430);
nor U17160 (N_17160,N_8185,N_5993);
and U17161 (N_17161,N_3978,N_5566);
or U17162 (N_17162,N_8188,N_1087);
or U17163 (N_17163,N_123,N_6320);
nor U17164 (N_17164,N_1359,N_8524);
or U17165 (N_17165,N_5470,N_8855);
or U17166 (N_17166,N_6226,N_3095);
and U17167 (N_17167,N_9530,N_6310);
nor U17168 (N_17168,N_1313,N_7930);
or U17169 (N_17169,N_6177,N_9270);
nor U17170 (N_17170,N_7492,N_308);
and U17171 (N_17171,N_1425,N_3190);
nand U17172 (N_17172,N_1141,N_7912);
nand U17173 (N_17173,N_4838,N_1288);
nor U17174 (N_17174,N_1588,N_429);
nand U17175 (N_17175,N_4527,N_5845);
or U17176 (N_17176,N_4371,N_1554);
nand U17177 (N_17177,N_8713,N_7882);
and U17178 (N_17178,N_5999,N_6633);
nand U17179 (N_17179,N_8274,N_389);
nand U17180 (N_17180,N_7252,N_2822);
or U17181 (N_17181,N_4012,N_8694);
nor U17182 (N_17182,N_4547,N_1742);
nand U17183 (N_17183,N_4166,N_9885);
and U17184 (N_17184,N_8231,N_2285);
nor U17185 (N_17185,N_1663,N_1343);
nand U17186 (N_17186,N_4149,N_7479);
and U17187 (N_17187,N_6506,N_255);
nand U17188 (N_17188,N_8756,N_3761);
nor U17189 (N_17189,N_3115,N_2866);
or U17190 (N_17190,N_553,N_9104);
nand U17191 (N_17191,N_6300,N_7735);
or U17192 (N_17192,N_9363,N_4579);
or U17193 (N_17193,N_7112,N_2072);
nand U17194 (N_17194,N_9960,N_7462);
nor U17195 (N_17195,N_1153,N_8575);
or U17196 (N_17196,N_9251,N_7744);
nor U17197 (N_17197,N_659,N_520);
nor U17198 (N_17198,N_8201,N_7868);
and U17199 (N_17199,N_5654,N_5666);
nor U17200 (N_17200,N_5036,N_5113);
nand U17201 (N_17201,N_40,N_6049);
and U17202 (N_17202,N_3653,N_2819);
nand U17203 (N_17203,N_8758,N_4386);
or U17204 (N_17204,N_3784,N_4738);
or U17205 (N_17205,N_1991,N_4498);
nor U17206 (N_17206,N_3905,N_4456);
or U17207 (N_17207,N_9562,N_5245);
and U17208 (N_17208,N_2821,N_7502);
and U17209 (N_17209,N_6927,N_617);
nor U17210 (N_17210,N_386,N_8620);
and U17211 (N_17211,N_2838,N_8702);
nand U17212 (N_17212,N_1306,N_7863);
and U17213 (N_17213,N_5320,N_8786);
or U17214 (N_17214,N_4435,N_6629);
nor U17215 (N_17215,N_5157,N_763);
and U17216 (N_17216,N_5571,N_2593);
or U17217 (N_17217,N_1695,N_7531);
nor U17218 (N_17218,N_5370,N_8395);
nor U17219 (N_17219,N_381,N_6336);
nand U17220 (N_17220,N_1432,N_5302);
nor U17221 (N_17221,N_3812,N_9855);
nor U17222 (N_17222,N_9296,N_2200);
and U17223 (N_17223,N_6296,N_5632);
and U17224 (N_17224,N_9883,N_6143);
or U17225 (N_17225,N_9599,N_8201);
or U17226 (N_17226,N_7857,N_958);
nor U17227 (N_17227,N_6610,N_90);
and U17228 (N_17228,N_8001,N_2769);
and U17229 (N_17229,N_8991,N_7507);
and U17230 (N_17230,N_8037,N_8302);
or U17231 (N_17231,N_6756,N_4517);
nor U17232 (N_17232,N_6760,N_3013);
nor U17233 (N_17233,N_6326,N_7378);
nand U17234 (N_17234,N_4984,N_8197);
or U17235 (N_17235,N_4795,N_3042);
nor U17236 (N_17236,N_1082,N_5673);
nand U17237 (N_17237,N_9914,N_4119);
or U17238 (N_17238,N_7680,N_3828);
nand U17239 (N_17239,N_8798,N_6563);
and U17240 (N_17240,N_5786,N_9795);
and U17241 (N_17241,N_3789,N_1001);
or U17242 (N_17242,N_2508,N_1426);
and U17243 (N_17243,N_5444,N_7993);
and U17244 (N_17244,N_6147,N_4907);
or U17245 (N_17245,N_1067,N_1690);
or U17246 (N_17246,N_1675,N_6936);
nand U17247 (N_17247,N_9631,N_7466);
or U17248 (N_17248,N_1342,N_9542);
or U17249 (N_17249,N_3981,N_1905);
and U17250 (N_17250,N_4690,N_3330);
nand U17251 (N_17251,N_557,N_9640);
nor U17252 (N_17252,N_318,N_7520);
nor U17253 (N_17253,N_32,N_4918);
xor U17254 (N_17254,N_3320,N_6497);
nand U17255 (N_17255,N_4245,N_7378);
nor U17256 (N_17256,N_971,N_9443);
or U17257 (N_17257,N_6428,N_249);
nand U17258 (N_17258,N_4515,N_4885);
nand U17259 (N_17259,N_155,N_8997);
nor U17260 (N_17260,N_3367,N_1708);
nand U17261 (N_17261,N_1055,N_5402);
and U17262 (N_17262,N_3582,N_4042);
and U17263 (N_17263,N_3766,N_2746);
nand U17264 (N_17264,N_3429,N_9377);
nor U17265 (N_17265,N_924,N_8665);
or U17266 (N_17266,N_4087,N_9252);
nor U17267 (N_17267,N_4309,N_891);
nor U17268 (N_17268,N_2908,N_7110);
nand U17269 (N_17269,N_5976,N_7001);
nand U17270 (N_17270,N_4902,N_7702);
and U17271 (N_17271,N_2009,N_9532);
or U17272 (N_17272,N_2788,N_4121);
nand U17273 (N_17273,N_3025,N_5088);
nand U17274 (N_17274,N_5160,N_3514);
nor U17275 (N_17275,N_8679,N_1563);
or U17276 (N_17276,N_6242,N_5948);
or U17277 (N_17277,N_5633,N_6040);
nand U17278 (N_17278,N_8448,N_3113);
nor U17279 (N_17279,N_4887,N_6685);
nor U17280 (N_17280,N_8119,N_3544);
nor U17281 (N_17281,N_1587,N_4022);
and U17282 (N_17282,N_9931,N_3912);
or U17283 (N_17283,N_6897,N_8627);
and U17284 (N_17284,N_961,N_6079);
nand U17285 (N_17285,N_9271,N_3308);
and U17286 (N_17286,N_3642,N_568);
and U17287 (N_17287,N_1456,N_3003);
nor U17288 (N_17288,N_6764,N_2213);
or U17289 (N_17289,N_1832,N_4427);
nand U17290 (N_17290,N_5256,N_6856);
or U17291 (N_17291,N_5470,N_52);
and U17292 (N_17292,N_4153,N_9690);
and U17293 (N_17293,N_157,N_1264);
or U17294 (N_17294,N_2460,N_7938);
or U17295 (N_17295,N_9836,N_8521);
nor U17296 (N_17296,N_9968,N_3722);
or U17297 (N_17297,N_4699,N_6989);
nor U17298 (N_17298,N_5549,N_5916);
or U17299 (N_17299,N_8521,N_1824);
nand U17300 (N_17300,N_517,N_9827);
nand U17301 (N_17301,N_7939,N_9233);
or U17302 (N_17302,N_8388,N_1208);
or U17303 (N_17303,N_8745,N_6866);
nor U17304 (N_17304,N_7512,N_3699);
xor U17305 (N_17305,N_8184,N_4833);
nand U17306 (N_17306,N_4052,N_8874);
nand U17307 (N_17307,N_6138,N_1201);
or U17308 (N_17308,N_2926,N_4004);
or U17309 (N_17309,N_28,N_9776);
nor U17310 (N_17310,N_7003,N_2735);
nand U17311 (N_17311,N_1146,N_5502);
nand U17312 (N_17312,N_7784,N_5226);
nor U17313 (N_17313,N_5088,N_3234);
nand U17314 (N_17314,N_3024,N_6842);
or U17315 (N_17315,N_7289,N_7419);
or U17316 (N_17316,N_2654,N_2364);
nor U17317 (N_17317,N_4886,N_6411);
nor U17318 (N_17318,N_6352,N_3205);
or U17319 (N_17319,N_1525,N_9773);
or U17320 (N_17320,N_9122,N_819);
nand U17321 (N_17321,N_8050,N_5375);
xor U17322 (N_17322,N_6037,N_2128);
or U17323 (N_17323,N_4363,N_2369);
nand U17324 (N_17324,N_2258,N_5305);
nand U17325 (N_17325,N_9974,N_1313);
nand U17326 (N_17326,N_3606,N_9232);
or U17327 (N_17327,N_2879,N_7164);
and U17328 (N_17328,N_2608,N_1883);
and U17329 (N_17329,N_7441,N_7813);
nand U17330 (N_17330,N_5185,N_6756);
nand U17331 (N_17331,N_146,N_8979);
and U17332 (N_17332,N_8693,N_4999);
nor U17333 (N_17333,N_4318,N_2122);
nor U17334 (N_17334,N_5371,N_1054);
nor U17335 (N_17335,N_6048,N_9821);
xnor U17336 (N_17336,N_753,N_3477);
and U17337 (N_17337,N_9737,N_2762);
or U17338 (N_17338,N_2130,N_653);
and U17339 (N_17339,N_1568,N_7794);
or U17340 (N_17340,N_7418,N_2428);
and U17341 (N_17341,N_6546,N_5985);
nor U17342 (N_17342,N_5697,N_2242);
nand U17343 (N_17343,N_854,N_2622);
or U17344 (N_17344,N_2817,N_8638);
nor U17345 (N_17345,N_3699,N_1826);
nor U17346 (N_17346,N_6001,N_8897);
nand U17347 (N_17347,N_1002,N_424);
and U17348 (N_17348,N_5250,N_3554);
nor U17349 (N_17349,N_3310,N_1699);
or U17350 (N_17350,N_9407,N_9547);
nor U17351 (N_17351,N_640,N_5586);
nor U17352 (N_17352,N_3282,N_1096);
nand U17353 (N_17353,N_2536,N_3345);
or U17354 (N_17354,N_2732,N_2856);
or U17355 (N_17355,N_947,N_5465);
nor U17356 (N_17356,N_9422,N_8248);
nand U17357 (N_17357,N_7194,N_1246);
and U17358 (N_17358,N_6117,N_4894);
or U17359 (N_17359,N_3541,N_8962);
or U17360 (N_17360,N_3702,N_792);
or U17361 (N_17361,N_6904,N_532);
nor U17362 (N_17362,N_5895,N_2053);
nand U17363 (N_17363,N_8428,N_8717);
and U17364 (N_17364,N_9997,N_3298);
and U17365 (N_17365,N_5917,N_563);
nand U17366 (N_17366,N_365,N_4265);
or U17367 (N_17367,N_926,N_8794);
or U17368 (N_17368,N_4523,N_9344);
nand U17369 (N_17369,N_1034,N_2554);
nand U17370 (N_17370,N_705,N_4029);
nand U17371 (N_17371,N_7408,N_3137);
and U17372 (N_17372,N_1728,N_1597);
nand U17373 (N_17373,N_3658,N_3131);
and U17374 (N_17374,N_6704,N_9904);
nand U17375 (N_17375,N_1796,N_6780);
nor U17376 (N_17376,N_108,N_3262);
nand U17377 (N_17377,N_1376,N_6053);
or U17378 (N_17378,N_376,N_7102);
nand U17379 (N_17379,N_2849,N_769);
nand U17380 (N_17380,N_4428,N_289);
or U17381 (N_17381,N_3303,N_1666);
or U17382 (N_17382,N_3404,N_9668);
nor U17383 (N_17383,N_7672,N_3738);
or U17384 (N_17384,N_9920,N_9415);
nor U17385 (N_17385,N_8908,N_8922);
or U17386 (N_17386,N_5214,N_2091);
nand U17387 (N_17387,N_6713,N_4228);
or U17388 (N_17388,N_723,N_5129);
nor U17389 (N_17389,N_8212,N_9247);
and U17390 (N_17390,N_9092,N_6256);
and U17391 (N_17391,N_4352,N_9104);
or U17392 (N_17392,N_7969,N_3068);
or U17393 (N_17393,N_3604,N_8076);
and U17394 (N_17394,N_9636,N_5727);
and U17395 (N_17395,N_6800,N_6724);
nand U17396 (N_17396,N_9124,N_2263);
and U17397 (N_17397,N_4650,N_1769);
nand U17398 (N_17398,N_6778,N_3841);
nand U17399 (N_17399,N_3955,N_7730);
nand U17400 (N_17400,N_9339,N_3679);
and U17401 (N_17401,N_2342,N_2842);
or U17402 (N_17402,N_7174,N_3325);
nor U17403 (N_17403,N_3989,N_6242);
nor U17404 (N_17404,N_2920,N_694);
or U17405 (N_17405,N_6978,N_3892);
nor U17406 (N_17406,N_3740,N_3103);
and U17407 (N_17407,N_4942,N_2739);
or U17408 (N_17408,N_7013,N_2959);
and U17409 (N_17409,N_3603,N_2125);
nand U17410 (N_17410,N_8298,N_6464);
nand U17411 (N_17411,N_8376,N_9685);
nand U17412 (N_17412,N_2255,N_4881);
nor U17413 (N_17413,N_7112,N_8366);
and U17414 (N_17414,N_4893,N_858);
nand U17415 (N_17415,N_7017,N_627);
nor U17416 (N_17416,N_6636,N_1902);
and U17417 (N_17417,N_468,N_3062);
nand U17418 (N_17418,N_7849,N_2480);
nor U17419 (N_17419,N_2343,N_9460);
nor U17420 (N_17420,N_3253,N_410);
nor U17421 (N_17421,N_8581,N_7931);
nand U17422 (N_17422,N_2905,N_1417);
nor U17423 (N_17423,N_2857,N_8706);
or U17424 (N_17424,N_6411,N_6994);
nor U17425 (N_17425,N_2141,N_4759);
or U17426 (N_17426,N_7287,N_533);
nor U17427 (N_17427,N_3715,N_776);
nand U17428 (N_17428,N_7099,N_169);
nor U17429 (N_17429,N_60,N_7294);
or U17430 (N_17430,N_5360,N_7577);
or U17431 (N_17431,N_7416,N_9461);
nor U17432 (N_17432,N_4984,N_4543);
and U17433 (N_17433,N_6193,N_6656);
or U17434 (N_17434,N_498,N_1187);
and U17435 (N_17435,N_3523,N_8785);
xnor U17436 (N_17436,N_9835,N_2313);
nor U17437 (N_17437,N_9479,N_6023);
and U17438 (N_17438,N_5775,N_8337);
or U17439 (N_17439,N_7517,N_8334);
nand U17440 (N_17440,N_9877,N_4830);
nor U17441 (N_17441,N_6551,N_7162);
or U17442 (N_17442,N_6367,N_894);
and U17443 (N_17443,N_1279,N_7772);
or U17444 (N_17444,N_6221,N_3218);
nor U17445 (N_17445,N_4214,N_7531);
nor U17446 (N_17446,N_2209,N_4694);
and U17447 (N_17447,N_9018,N_9135);
nor U17448 (N_17448,N_4744,N_1292);
and U17449 (N_17449,N_9027,N_6088);
nor U17450 (N_17450,N_9786,N_3093);
or U17451 (N_17451,N_242,N_9094);
nor U17452 (N_17452,N_9272,N_1531);
nor U17453 (N_17453,N_9032,N_3102);
nor U17454 (N_17454,N_7961,N_6170);
nor U17455 (N_17455,N_5224,N_152);
and U17456 (N_17456,N_8481,N_3993);
and U17457 (N_17457,N_4611,N_9520);
and U17458 (N_17458,N_6089,N_6486);
or U17459 (N_17459,N_9847,N_2925);
and U17460 (N_17460,N_7423,N_9993);
nand U17461 (N_17461,N_5560,N_2441);
nor U17462 (N_17462,N_9303,N_9223);
nor U17463 (N_17463,N_7862,N_1814);
and U17464 (N_17464,N_1023,N_6525);
nand U17465 (N_17465,N_8338,N_3865);
nor U17466 (N_17466,N_5674,N_3329);
or U17467 (N_17467,N_8867,N_1835);
nand U17468 (N_17468,N_8861,N_9998);
nor U17469 (N_17469,N_2848,N_8011);
and U17470 (N_17470,N_2060,N_718);
or U17471 (N_17471,N_6435,N_6004);
nor U17472 (N_17472,N_2053,N_2676);
or U17473 (N_17473,N_733,N_6911);
nand U17474 (N_17474,N_5084,N_8991);
nand U17475 (N_17475,N_2168,N_6211);
and U17476 (N_17476,N_9621,N_9390);
nand U17477 (N_17477,N_4100,N_8921);
nand U17478 (N_17478,N_5432,N_1078);
nand U17479 (N_17479,N_9401,N_8051);
and U17480 (N_17480,N_9517,N_5368);
nor U17481 (N_17481,N_234,N_194);
nor U17482 (N_17482,N_9847,N_1254);
and U17483 (N_17483,N_7890,N_7389);
and U17484 (N_17484,N_1450,N_7105);
nor U17485 (N_17485,N_684,N_6711);
or U17486 (N_17486,N_2427,N_752);
nor U17487 (N_17487,N_8040,N_6092);
nor U17488 (N_17488,N_2732,N_9509);
nand U17489 (N_17489,N_8611,N_2760);
or U17490 (N_17490,N_5790,N_3138);
nand U17491 (N_17491,N_2331,N_2254);
and U17492 (N_17492,N_5823,N_6433);
nor U17493 (N_17493,N_3556,N_4484);
nand U17494 (N_17494,N_7039,N_3161);
or U17495 (N_17495,N_225,N_7101);
and U17496 (N_17496,N_542,N_9826);
and U17497 (N_17497,N_2485,N_6143);
and U17498 (N_17498,N_2389,N_9913);
and U17499 (N_17499,N_9526,N_5294);
nor U17500 (N_17500,N_6923,N_8218);
or U17501 (N_17501,N_7965,N_2356);
nor U17502 (N_17502,N_7995,N_2146);
nand U17503 (N_17503,N_4750,N_5797);
nand U17504 (N_17504,N_5774,N_1662);
or U17505 (N_17505,N_2176,N_7135);
nand U17506 (N_17506,N_2494,N_9480);
or U17507 (N_17507,N_8033,N_2864);
or U17508 (N_17508,N_8931,N_6470);
and U17509 (N_17509,N_877,N_7981);
nor U17510 (N_17510,N_689,N_6884);
nand U17511 (N_17511,N_6695,N_9898);
and U17512 (N_17512,N_4795,N_7799);
and U17513 (N_17513,N_3108,N_1377);
nor U17514 (N_17514,N_1845,N_9210);
and U17515 (N_17515,N_370,N_3870);
nor U17516 (N_17516,N_8298,N_6947);
nand U17517 (N_17517,N_1485,N_7139);
or U17518 (N_17518,N_297,N_4312);
nor U17519 (N_17519,N_2815,N_8280);
nor U17520 (N_17520,N_9301,N_632);
or U17521 (N_17521,N_5315,N_2947);
nand U17522 (N_17522,N_2485,N_1947);
nor U17523 (N_17523,N_5020,N_5054);
and U17524 (N_17524,N_470,N_4729);
nand U17525 (N_17525,N_115,N_5658);
nand U17526 (N_17526,N_5760,N_1115);
or U17527 (N_17527,N_1461,N_9996);
or U17528 (N_17528,N_8396,N_2133);
nand U17529 (N_17529,N_4451,N_6262);
and U17530 (N_17530,N_9263,N_8502);
and U17531 (N_17531,N_2775,N_2784);
and U17532 (N_17532,N_9352,N_8564);
or U17533 (N_17533,N_4165,N_1936);
or U17534 (N_17534,N_9852,N_1481);
nand U17535 (N_17535,N_8753,N_4587);
nor U17536 (N_17536,N_1891,N_724);
and U17537 (N_17537,N_9741,N_5210);
nor U17538 (N_17538,N_8176,N_664);
nor U17539 (N_17539,N_3651,N_336);
nand U17540 (N_17540,N_7936,N_592);
xor U17541 (N_17541,N_5326,N_6931);
nor U17542 (N_17542,N_6518,N_5125);
or U17543 (N_17543,N_2092,N_5930);
or U17544 (N_17544,N_5759,N_2664);
nand U17545 (N_17545,N_1896,N_2636);
or U17546 (N_17546,N_4297,N_2179);
or U17547 (N_17547,N_1754,N_2010);
and U17548 (N_17548,N_8836,N_8436);
nor U17549 (N_17549,N_8920,N_1336);
and U17550 (N_17550,N_7961,N_8129);
and U17551 (N_17551,N_5149,N_9102);
and U17552 (N_17552,N_2180,N_3460);
nand U17553 (N_17553,N_4514,N_3095);
or U17554 (N_17554,N_9359,N_9501);
or U17555 (N_17555,N_2763,N_3907);
and U17556 (N_17556,N_2508,N_1461);
or U17557 (N_17557,N_1835,N_3131);
nor U17558 (N_17558,N_2412,N_2075);
nand U17559 (N_17559,N_3878,N_8043);
or U17560 (N_17560,N_2894,N_7535);
nor U17561 (N_17561,N_1191,N_2971);
nor U17562 (N_17562,N_9209,N_9308);
and U17563 (N_17563,N_8717,N_1749);
or U17564 (N_17564,N_7116,N_8551);
and U17565 (N_17565,N_7345,N_1212);
nor U17566 (N_17566,N_5063,N_1586);
nor U17567 (N_17567,N_4640,N_8977);
nand U17568 (N_17568,N_3256,N_4144);
nor U17569 (N_17569,N_3331,N_528);
nor U17570 (N_17570,N_6470,N_3450);
or U17571 (N_17571,N_856,N_8773);
nand U17572 (N_17572,N_3067,N_5462);
nand U17573 (N_17573,N_1408,N_3483);
or U17574 (N_17574,N_3536,N_8498);
nand U17575 (N_17575,N_8137,N_7359);
or U17576 (N_17576,N_2222,N_901);
or U17577 (N_17577,N_3055,N_7433);
nor U17578 (N_17578,N_135,N_4039);
nand U17579 (N_17579,N_2491,N_645);
nor U17580 (N_17580,N_5496,N_9011);
nand U17581 (N_17581,N_3078,N_4521);
and U17582 (N_17582,N_3059,N_7302);
nand U17583 (N_17583,N_6650,N_2463);
or U17584 (N_17584,N_7890,N_3768);
nor U17585 (N_17585,N_744,N_6787);
and U17586 (N_17586,N_2652,N_3999);
nor U17587 (N_17587,N_7603,N_9367);
nand U17588 (N_17588,N_8272,N_7780);
and U17589 (N_17589,N_2654,N_1622);
nor U17590 (N_17590,N_1880,N_2039);
and U17591 (N_17591,N_2634,N_3641);
or U17592 (N_17592,N_2795,N_7204);
nand U17593 (N_17593,N_905,N_8023);
nand U17594 (N_17594,N_1479,N_1142);
nor U17595 (N_17595,N_9494,N_3874);
nor U17596 (N_17596,N_6404,N_4341);
and U17597 (N_17597,N_5271,N_886);
nor U17598 (N_17598,N_2172,N_5361);
nand U17599 (N_17599,N_13,N_7371);
nand U17600 (N_17600,N_1308,N_7853);
and U17601 (N_17601,N_7443,N_1938);
nor U17602 (N_17602,N_592,N_375);
nor U17603 (N_17603,N_9669,N_6921);
nand U17604 (N_17604,N_9944,N_1750);
and U17605 (N_17605,N_2935,N_6605);
nor U17606 (N_17606,N_9006,N_1633);
nor U17607 (N_17607,N_3593,N_8075);
and U17608 (N_17608,N_500,N_1670);
nor U17609 (N_17609,N_5503,N_2626);
nand U17610 (N_17610,N_6061,N_9820);
nand U17611 (N_17611,N_9252,N_3964);
and U17612 (N_17612,N_6166,N_7303);
nand U17613 (N_17613,N_6745,N_4843);
nand U17614 (N_17614,N_2071,N_3382);
nand U17615 (N_17615,N_3388,N_9035);
or U17616 (N_17616,N_6434,N_6029);
and U17617 (N_17617,N_8825,N_4399);
nor U17618 (N_17618,N_7118,N_5431);
and U17619 (N_17619,N_3317,N_5941);
and U17620 (N_17620,N_3404,N_6656);
nor U17621 (N_17621,N_5347,N_9022);
or U17622 (N_17622,N_831,N_424);
nor U17623 (N_17623,N_8080,N_5360);
nand U17624 (N_17624,N_8127,N_3792);
nand U17625 (N_17625,N_3437,N_7232);
nor U17626 (N_17626,N_3778,N_8506);
and U17627 (N_17627,N_3906,N_361);
and U17628 (N_17628,N_1374,N_5213);
and U17629 (N_17629,N_924,N_9706);
nand U17630 (N_17630,N_1945,N_6946);
nand U17631 (N_17631,N_1725,N_195);
or U17632 (N_17632,N_6503,N_9411);
or U17633 (N_17633,N_1139,N_651);
nand U17634 (N_17634,N_5111,N_4480);
nor U17635 (N_17635,N_7912,N_6481);
nor U17636 (N_17636,N_5500,N_6665);
nor U17637 (N_17637,N_9578,N_2654);
and U17638 (N_17638,N_1922,N_3806);
nor U17639 (N_17639,N_7370,N_2626);
nand U17640 (N_17640,N_4833,N_3769);
or U17641 (N_17641,N_8462,N_6215);
or U17642 (N_17642,N_3351,N_4312);
or U17643 (N_17643,N_8130,N_4937);
nor U17644 (N_17644,N_1930,N_8463);
nor U17645 (N_17645,N_7099,N_3378);
xnor U17646 (N_17646,N_4050,N_2606);
or U17647 (N_17647,N_1712,N_373);
or U17648 (N_17648,N_4222,N_1854);
nor U17649 (N_17649,N_9454,N_6818);
nand U17650 (N_17650,N_4665,N_6672);
nor U17651 (N_17651,N_6354,N_9525);
nand U17652 (N_17652,N_1237,N_6502);
nor U17653 (N_17653,N_828,N_6883);
nand U17654 (N_17654,N_5129,N_2997);
nor U17655 (N_17655,N_7646,N_7752);
nor U17656 (N_17656,N_9952,N_3879);
nand U17657 (N_17657,N_7884,N_7035);
nand U17658 (N_17658,N_9735,N_1538);
nand U17659 (N_17659,N_7503,N_2558);
or U17660 (N_17660,N_1305,N_2543);
and U17661 (N_17661,N_2919,N_2101);
nand U17662 (N_17662,N_6445,N_2363);
and U17663 (N_17663,N_5712,N_9466);
or U17664 (N_17664,N_9264,N_2350);
and U17665 (N_17665,N_7964,N_2497);
nand U17666 (N_17666,N_4659,N_6415);
nand U17667 (N_17667,N_7450,N_1056);
and U17668 (N_17668,N_2606,N_5580);
and U17669 (N_17669,N_6988,N_6335);
or U17670 (N_17670,N_4727,N_4202);
nor U17671 (N_17671,N_8938,N_9423);
nand U17672 (N_17672,N_8581,N_877);
or U17673 (N_17673,N_5766,N_9885);
and U17674 (N_17674,N_4530,N_1202);
nand U17675 (N_17675,N_7519,N_941);
or U17676 (N_17676,N_6911,N_9972);
or U17677 (N_17677,N_7005,N_6973);
and U17678 (N_17678,N_8262,N_4234);
nand U17679 (N_17679,N_6349,N_693);
nand U17680 (N_17680,N_1816,N_2719);
nor U17681 (N_17681,N_2448,N_6672);
or U17682 (N_17682,N_7975,N_5947);
or U17683 (N_17683,N_7649,N_9432);
nor U17684 (N_17684,N_3397,N_6943);
nand U17685 (N_17685,N_6143,N_21);
nand U17686 (N_17686,N_936,N_1589);
nand U17687 (N_17687,N_7244,N_7679);
or U17688 (N_17688,N_3411,N_6245);
and U17689 (N_17689,N_1990,N_4461);
nor U17690 (N_17690,N_7065,N_625);
and U17691 (N_17691,N_3779,N_2382);
or U17692 (N_17692,N_3006,N_6462);
or U17693 (N_17693,N_7867,N_5631);
and U17694 (N_17694,N_387,N_2582);
or U17695 (N_17695,N_5593,N_8481);
or U17696 (N_17696,N_2255,N_4648);
nor U17697 (N_17697,N_2777,N_3202);
nand U17698 (N_17698,N_8840,N_4908);
and U17699 (N_17699,N_1152,N_7250);
xor U17700 (N_17700,N_9109,N_9843);
nand U17701 (N_17701,N_1420,N_48);
nand U17702 (N_17702,N_2053,N_2745);
nor U17703 (N_17703,N_4493,N_7651);
or U17704 (N_17704,N_1342,N_3707);
nor U17705 (N_17705,N_5747,N_4592);
or U17706 (N_17706,N_5402,N_1567);
or U17707 (N_17707,N_2529,N_5819);
nor U17708 (N_17708,N_9317,N_4984);
and U17709 (N_17709,N_2384,N_3065);
and U17710 (N_17710,N_8059,N_9203);
or U17711 (N_17711,N_6358,N_7286);
nor U17712 (N_17712,N_8653,N_4590);
or U17713 (N_17713,N_6284,N_5187);
nor U17714 (N_17714,N_2016,N_9794);
nor U17715 (N_17715,N_4436,N_5421);
or U17716 (N_17716,N_6581,N_2552);
nor U17717 (N_17717,N_9016,N_1476);
and U17718 (N_17718,N_4499,N_424);
and U17719 (N_17719,N_2889,N_7285);
nor U17720 (N_17720,N_2343,N_7535);
nand U17721 (N_17721,N_7246,N_4978);
nor U17722 (N_17722,N_8243,N_6360);
nor U17723 (N_17723,N_9450,N_2716);
nor U17724 (N_17724,N_6140,N_2655);
or U17725 (N_17725,N_8293,N_1178);
and U17726 (N_17726,N_8765,N_4375);
nand U17727 (N_17727,N_6642,N_9603);
nor U17728 (N_17728,N_6003,N_7886);
nand U17729 (N_17729,N_4914,N_5892);
nand U17730 (N_17730,N_6695,N_1553);
nand U17731 (N_17731,N_154,N_4569);
or U17732 (N_17732,N_2329,N_5812);
nand U17733 (N_17733,N_7448,N_4558);
or U17734 (N_17734,N_6674,N_7737);
nand U17735 (N_17735,N_3491,N_8841);
nor U17736 (N_17736,N_8459,N_742);
nand U17737 (N_17737,N_7795,N_9147);
and U17738 (N_17738,N_4687,N_5799);
nand U17739 (N_17739,N_671,N_8922);
or U17740 (N_17740,N_366,N_3408);
nand U17741 (N_17741,N_9824,N_3020);
nand U17742 (N_17742,N_9702,N_1139);
nand U17743 (N_17743,N_6577,N_351);
nand U17744 (N_17744,N_5919,N_4922);
nand U17745 (N_17745,N_7639,N_6497);
and U17746 (N_17746,N_1910,N_1413);
nor U17747 (N_17747,N_8366,N_4279);
or U17748 (N_17748,N_8184,N_1716);
or U17749 (N_17749,N_7419,N_82);
or U17750 (N_17750,N_4751,N_5818);
or U17751 (N_17751,N_3473,N_6460);
nor U17752 (N_17752,N_7323,N_9306);
and U17753 (N_17753,N_6742,N_3546);
nor U17754 (N_17754,N_8255,N_8627);
and U17755 (N_17755,N_1298,N_8098);
or U17756 (N_17756,N_4816,N_5643);
or U17757 (N_17757,N_9230,N_7891);
and U17758 (N_17758,N_5534,N_5941);
nand U17759 (N_17759,N_5651,N_9503);
and U17760 (N_17760,N_3364,N_7363);
nand U17761 (N_17761,N_3015,N_9647);
and U17762 (N_17762,N_9410,N_5006);
or U17763 (N_17763,N_4134,N_4150);
nand U17764 (N_17764,N_9799,N_5972);
nor U17765 (N_17765,N_5479,N_407);
and U17766 (N_17766,N_1744,N_4529);
nand U17767 (N_17767,N_2340,N_1828);
nor U17768 (N_17768,N_4229,N_7846);
nor U17769 (N_17769,N_3258,N_3091);
and U17770 (N_17770,N_6141,N_3323);
or U17771 (N_17771,N_9849,N_8303);
or U17772 (N_17772,N_7461,N_1865);
nor U17773 (N_17773,N_4700,N_2334);
and U17774 (N_17774,N_7986,N_3419);
nand U17775 (N_17775,N_3576,N_4978);
and U17776 (N_17776,N_8858,N_7496);
nor U17777 (N_17777,N_1712,N_6177);
or U17778 (N_17778,N_6232,N_2174);
or U17779 (N_17779,N_7507,N_3944);
or U17780 (N_17780,N_448,N_1320);
and U17781 (N_17781,N_2437,N_7530);
or U17782 (N_17782,N_399,N_2876);
nand U17783 (N_17783,N_4943,N_8046);
nand U17784 (N_17784,N_7380,N_4229);
nand U17785 (N_17785,N_8665,N_5234);
nand U17786 (N_17786,N_6761,N_9410);
nand U17787 (N_17787,N_3249,N_6786);
and U17788 (N_17788,N_2483,N_3891);
or U17789 (N_17789,N_6099,N_1902);
or U17790 (N_17790,N_4389,N_403);
nand U17791 (N_17791,N_4754,N_2664);
or U17792 (N_17792,N_2427,N_4044);
nand U17793 (N_17793,N_8231,N_8252);
nor U17794 (N_17794,N_9722,N_6174);
or U17795 (N_17795,N_5089,N_8016);
or U17796 (N_17796,N_7372,N_5774);
and U17797 (N_17797,N_8525,N_280);
and U17798 (N_17798,N_4660,N_9176);
nor U17799 (N_17799,N_2008,N_1522);
nand U17800 (N_17800,N_7946,N_9488);
or U17801 (N_17801,N_2030,N_7703);
nand U17802 (N_17802,N_7532,N_9705);
and U17803 (N_17803,N_4207,N_3007);
nor U17804 (N_17804,N_3763,N_9801);
nand U17805 (N_17805,N_6618,N_7571);
or U17806 (N_17806,N_2413,N_3171);
nand U17807 (N_17807,N_7123,N_6172);
nor U17808 (N_17808,N_6441,N_1340);
nand U17809 (N_17809,N_7629,N_7426);
or U17810 (N_17810,N_3603,N_2178);
and U17811 (N_17811,N_5935,N_4718);
nor U17812 (N_17812,N_1794,N_7285);
or U17813 (N_17813,N_7561,N_6155);
nor U17814 (N_17814,N_8924,N_2436);
nor U17815 (N_17815,N_6459,N_8471);
nand U17816 (N_17816,N_7792,N_5974);
nand U17817 (N_17817,N_948,N_6853);
or U17818 (N_17818,N_4895,N_5326);
or U17819 (N_17819,N_2333,N_3322);
nor U17820 (N_17820,N_4138,N_4739);
nor U17821 (N_17821,N_5600,N_4943);
or U17822 (N_17822,N_4293,N_1136);
and U17823 (N_17823,N_9215,N_9361);
nor U17824 (N_17824,N_5879,N_2419);
nor U17825 (N_17825,N_8632,N_1911);
nor U17826 (N_17826,N_6216,N_2584);
or U17827 (N_17827,N_8901,N_8363);
nor U17828 (N_17828,N_920,N_679);
nand U17829 (N_17829,N_1863,N_3650);
or U17830 (N_17830,N_6658,N_3914);
or U17831 (N_17831,N_9916,N_4771);
nor U17832 (N_17832,N_3105,N_9196);
or U17833 (N_17833,N_9630,N_9196);
nor U17834 (N_17834,N_6545,N_4992);
xor U17835 (N_17835,N_8210,N_8966);
and U17836 (N_17836,N_410,N_5748);
and U17837 (N_17837,N_7179,N_2695);
nand U17838 (N_17838,N_7397,N_5231);
nor U17839 (N_17839,N_4846,N_8184);
nor U17840 (N_17840,N_159,N_9695);
or U17841 (N_17841,N_3470,N_3284);
or U17842 (N_17842,N_4693,N_9226);
nand U17843 (N_17843,N_4352,N_3054);
nor U17844 (N_17844,N_2614,N_4477);
or U17845 (N_17845,N_7966,N_8171);
nor U17846 (N_17846,N_2891,N_3398);
nor U17847 (N_17847,N_5691,N_1375);
and U17848 (N_17848,N_1468,N_875);
and U17849 (N_17849,N_4098,N_5792);
nand U17850 (N_17850,N_9804,N_3924);
xnor U17851 (N_17851,N_5013,N_7639);
nand U17852 (N_17852,N_3320,N_6650);
nand U17853 (N_17853,N_3551,N_1300);
nand U17854 (N_17854,N_4770,N_7105);
nor U17855 (N_17855,N_428,N_8649);
nor U17856 (N_17856,N_8792,N_2224);
nand U17857 (N_17857,N_2744,N_3391);
and U17858 (N_17858,N_1466,N_9983);
and U17859 (N_17859,N_6271,N_1188);
nand U17860 (N_17860,N_5682,N_5767);
and U17861 (N_17861,N_5227,N_5064);
nor U17862 (N_17862,N_9556,N_9939);
nand U17863 (N_17863,N_176,N_540);
and U17864 (N_17864,N_3416,N_2100);
xnor U17865 (N_17865,N_7391,N_8874);
nor U17866 (N_17866,N_8040,N_618);
and U17867 (N_17867,N_5641,N_1547);
nor U17868 (N_17868,N_8777,N_5995);
and U17869 (N_17869,N_7540,N_8208);
nor U17870 (N_17870,N_2849,N_6382);
or U17871 (N_17871,N_5667,N_8795);
and U17872 (N_17872,N_6339,N_1894);
or U17873 (N_17873,N_9474,N_9367);
or U17874 (N_17874,N_4349,N_1645);
nand U17875 (N_17875,N_7302,N_8781);
or U17876 (N_17876,N_9105,N_8909);
xnor U17877 (N_17877,N_5818,N_4046);
nand U17878 (N_17878,N_2585,N_9498);
or U17879 (N_17879,N_211,N_7979);
nor U17880 (N_17880,N_5738,N_9042);
nand U17881 (N_17881,N_6033,N_442);
nor U17882 (N_17882,N_899,N_55);
or U17883 (N_17883,N_8951,N_3118);
and U17884 (N_17884,N_6936,N_8921);
or U17885 (N_17885,N_7243,N_9500);
and U17886 (N_17886,N_4451,N_5192);
or U17887 (N_17887,N_7821,N_91);
and U17888 (N_17888,N_3189,N_4947);
nand U17889 (N_17889,N_1283,N_39);
xnor U17890 (N_17890,N_2196,N_8875);
nand U17891 (N_17891,N_2286,N_3402);
nand U17892 (N_17892,N_5725,N_6767);
or U17893 (N_17893,N_5680,N_6723);
or U17894 (N_17894,N_2553,N_9585);
and U17895 (N_17895,N_2768,N_5034);
nand U17896 (N_17896,N_2962,N_6232);
or U17897 (N_17897,N_5648,N_8248);
nand U17898 (N_17898,N_6485,N_6229);
nand U17899 (N_17899,N_3305,N_3601);
and U17900 (N_17900,N_8495,N_3485);
nor U17901 (N_17901,N_7985,N_7891);
nor U17902 (N_17902,N_7518,N_6418);
or U17903 (N_17903,N_9991,N_2812);
nand U17904 (N_17904,N_2232,N_477);
nand U17905 (N_17905,N_7285,N_1038);
nor U17906 (N_17906,N_1830,N_5221);
or U17907 (N_17907,N_6192,N_8735);
nand U17908 (N_17908,N_5046,N_4338);
nor U17909 (N_17909,N_6916,N_1645);
nor U17910 (N_17910,N_9073,N_5399);
nor U17911 (N_17911,N_8706,N_1375);
or U17912 (N_17912,N_6173,N_2823);
and U17913 (N_17913,N_5929,N_1400);
and U17914 (N_17914,N_1136,N_2521);
nor U17915 (N_17915,N_60,N_8041);
or U17916 (N_17916,N_4932,N_4740);
or U17917 (N_17917,N_1322,N_329);
and U17918 (N_17918,N_6862,N_1468);
and U17919 (N_17919,N_7950,N_2108);
xnor U17920 (N_17920,N_1475,N_5227);
or U17921 (N_17921,N_4511,N_8006);
nor U17922 (N_17922,N_1500,N_5054);
xor U17923 (N_17923,N_3512,N_3663);
or U17924 (N_17924,N_4209,N_4900);
nor U17925 (N_17925,N_7534,N_225);
or U17926 (N_17926,N_4773,N_23);
nand U17927 (N_17927,N_5465,N_7642);
nor U17928 (N_17928,N_2028,N_645);
and U17929 (N_17929,N_5723,N_4174);
nor U17930 (N_17930,N_3245,N_4402);
nand U17931 (N_17931,N_1785,N_1645);
nor U17932 (N_17932,N_9761,N_5387);
nand U17933 (N_17933,N_1153,N_7173);
nand U17934 (N_17934,N_5909,N_9742);
or U17935 (N_17935,N_5611,N_6059);
nor U17936 (N_17936,N_1913,N_5872);
and U17937 (N_17937,N_9581,N_6312);
nor U17938 (N_17938,N_5505,N_9996);
or U17939 (N_17939,N_3194,N_5202);
and U17940 (N_17940,N_1015,N_7548);
or U17941 (N_17941,N_7667,N_6218);
nor U17942 (N_17942,N_1242,N_6855);
nand U17943 (N_17943,N_3123,N_3187);
nor U17944 (N_17944,N_6285,N_4125);
and U17945 (N_17945,N_310,N_7865);
and U17946 (N_17946,N_4,N_212);
or U17947 (N_17947,N_8175,N_485);
or U17948 (N_17948,N_8287,N_9456);
nand U17949 (N_17949,N_6509,N_8392);
and U17950 (N_17950,N_2359,N_1877);
and U17951 (N_17951,N_9416,N_2338);
nand U17952 (N_17952,N_9480,N_4013);
or U17953 (N_17953,N_5060,N_3057);
nand U17954 (N_17954,N_3570,N_3864);
nand U17955 (N_17955,N_2799,N_5791);
nand U17956 (N_17956,N_5344,N_2908);
nand U17957 (N_17957,N_4440,N_5231);
nand U17958 (N_17958,N_6890,N_3691);
nand U17959 (N_17959,N_9488,N_5255);
and U17960 (N_17960,N_5055,N_7642);
nand U17961 (N_17961,N_201,N_8804);
xnor U17962 (N_17962,N_3376,N_3625);
nand U17963 (N_17963,N_9531,N_4447);
or U17964 (N_17964,N_7829,N_5087);
nor U17965 (N_17965,N_515,N_2703);
nor U17966 (N_17966,N_2465,N_8300);
and U17967 (N_17967,N_2026,N_807);
and U17968 (N_17968,N_5178,N_941);
and U17969 (N_17969,N_1067,N_5185);
nand U17970 (N_17970,N_5454,N_5869);
or U17971 (N_17971,N_1364,N_5617);
nand U17972 (N_17972,N_5414,N_9401);
or U17973 (N_17973,N_4217,N_4876);
nand U17974 (N_17974,N_3452,N_9433);
nor U17975 (N_17975,N_5097,N_5576);
and U17976 (N_17976,N_2557,N_9364);
nand U17977 (N_17977,N_9012,N_2716);
nand U17978 (N_17978,N_3732,N_6399);
and U17979 (N_17979,N_8261,N_69);
and U17980 (N_17980,N_2744,N_9471);
nand U17981 (N_17981,N_6120,N_854);
nor U17982 (N_17982,N_3757,N_314);
nor U17983 (N_17983,N_5696,N_1553);
and U17984 (N_17984,N_8818,N_587);
or U17985 (N_17985,N_5798,N_5969);
nor U17986 (N_17986,N_4946,N_3286);
nor U17987 (N_17987,N_3875,N_7202);
and U17988 (N_17988,N_8222,N_4933);
nor U17989 (N_17989,N_670,N_7929);
nand U17990 (N_17990,N_6633,N_4857);
nor U17991 (N_17991,N_7718,N_671);
nand U17992 (N_17992,N_5520,N_3300);
nand U17993 (N_17993,N_7722,N_3858);
nor U17994 (N_17994,N_6793,N_1589);
and U17995 (N_17995,N_5490,N_6663);
or U17996 (N_17996,N_2876,N_1501);
or U17997 (N_17997,N_1155,N_3158);
nor U17998 (N_17998,N_6005,N_2294);
nand U17999 (N_17999,N_9068,N_8137);
and U18000 (N_18000,N_5478,N_2227);
nand U18001 (N_18001,N_5511,N_5996);
nor U18002 (N_18002,N_1932,N_2648);
or U18003 (N_18003,N_1904,N_1886);
nand U18004 (N_18004,N_7056,N_2747);
nor U18005 (N_18005,N_3962,N_233);
nor U18006 (N_18006,N_3068,N_8863);
nor U18007 (N_18007,N_1096,N_3440);
nor U18008 (N_18008,N_4676,N_5223);
and U18009 (N_18009,N_7409,N_2843);
nor U18010 (N_18010,N_8558,N_3745);
nor U18011 (N_18011,N_8397,N_7350);
or U18012 (N_18012,N_8792,N_4973);
nand U18013 (N_18013,N_8916,N_596);
nor U18014 (N_18014,N_6389,N_1289);
nor U18015 (N_18015,N_4210,N_3700);
nand U18016 (N_18016,N_6313,N_4264);
nor U18017 (N_18017,N_7214,N_4806);
or U18018 (N_18018,N_2989,N_3171);
or U18019 (N_18019,N_4184,N_4253);
or U18020 (N_18020,N_8515,N_3906);
nor U18021 (N_18021,N_7013,N_1735);
and U18022 (N_18022,N_8884,N_3648);
nand U18023 (N_18023,N_8365,N_2719);
nand U18024 (N_18024,N_1474,N_8489);
nand U18025 (N_18025,N_9618,N_9959);
or U18026 (N_18026,N_8981,N_515);
nor U18027 (N_18027,N_839,N_902);
nor U18028 (N_18028,N_5439,N_9926);
nand U18029 (N_18029,N_9017,N_8785);
and U18030 (N_18030,N_432,N_8463);
and U18031 (N_18031,N_3051,N_8545);
or U18032 (N_18032,N_441,N_4300);
nand U18033 (N_18033,N_1495,N_6984);
nor U18034 (N_18034,N_1814,N_9473);
or U18035 (N_18035,N_3428,N_9536);
nor U18036 (N_18036,N_335,N_6846);
nor U18037 (N_18037,N_131,N_6868);
or U18038 (N_18038,N_4467,N_2999);
nand U18039 (N_18039,N_5062,N_4207);
nand U18040 (N_18040,N_9288,N_5055);
nor U18041 (N_18041,N_2716,N_3923);
nor U18042 (N_18042,N_6316,N_8617);
nand U18043 (N_18043,N_5907,N_6244);
nor U18044 (N_18044,N_67,N_8678);
or U18045 (N_18045,N_6051,N_9591);
nand U18046 (N_18046,N_2587,N_4397);
or U18047 (N_18047,N_7132,N_622);
nor U18048 (N_18048,N_493,N_710);
nand U18049 (N_18049,N_5094,N_4444);
nand U18050 (N_18050,N_9205,N_3603);
nor U18051 (N_18051,N_5215,N_1689);
nand U18052 (N_18052,N_6435,N_1560);
nor U18053 (N_18053,N_1959,N_9636);
or U18054 (N_18054,N_9855,N_6808);
and U18055 (N_18055,N_3100,N_8357);
or U18056 (N_18056,N_4114,N_2273);
and U18057 (N_18057,N_9817,N_3580);
or U18058 (N_18058,N_2152,N_6365);
and U18059 (N_18059,N_5766,N_3187);
nand U18060 (N_18060,N_3836,N_3762);
or U18061 (N_18061,N_7167,N_6035);
and U18062 (N_18062,N_1842,N_4828);
or U18063 (N_18063,N_6248,N_4929);
and U18064 (N_18064,N_4232,N_4431);
or U18065 (N_18065,N_335,N_110);
or U18066 (N_18066,N_4775,N_5927);
nor U18067 (N_18067,N_8585,N_3539);
and U18068 (N_18068,N_6247,N_8381);
nand U18069 (N_18069,N_5264,N_3316);
nor U18070 (N_18070,N_35,N_9226);
nor U18071 (N_18071,N_812,N_220);
or U18072 (N_18072,N_5220,N_9720);
nor U18073 (N_18073,N_4682,N_4060);
nor U18074 (N_18074,N_8118,N_9563);
and U18075 (N_18075,N_7466,N_8099);
and U18076 (N_18076,N_5231,N_7166);
nand U18077 (N_18077,N_8618,N_489);
or U18078 (N_18078,N_4547,N_3525);
and U18079 (N_18079,N_5798,N_9330);
nor U18080 (N_18080,N_7999,N_2583);
and U18081 (N_18081,N_5050,N_4333);
nand U18082 (N_18082,N_980,N_8188);
or U18083 (N_18083,N_3054,N_5413);
nor U18084 (N_18084,N_1788,N_8165);
nand U18085 (N_18085,N_8586,N_2361);
and U18086 (N_18086,N_627,N_9634);
nor U18087 (N_18087,N_8237,N_7260);
nand U18088 (N_18088,N_5059,N_3434);
nor U18089 (N_18089,N_4682,N_1986);
or U18090 (N_18090,N_7791,N_4860);
nand U18091 (N_18091,N_9491,N_991);
nand U18092 (N_18092,N_1276,N_8335);
nand U18093 (N_18093,N_340,N_236);
or U18094 (N_18094,N_8736,N_6222);
nand U18095 (N_18095,N_472,N_6939);
nor U18096 (N_18096,N_1772,N_2563);
and U18097 (N_18097,N_6151,N_2708);
and U18098 (N_18098,N_1604,N_5495);
or U18099 (N_18099,N_9541,N_9693);
or U18100 (N_18100,N_8890,N_3225);
or U18101 (N_18101,N_6029,N_7720);
nor U18102 (N_18102,N_8086,N_2866);
nor U18103 (N_18103,N_2933,N_4046);
nor U18104 (N_18104,N_1940,N_4495);
or U18105 (N_18105,N_9098,N_1203);
or U18106 (N_18106,N_1330,N_6999);
nand U18107 (N_18107,N_1619,N_6826);
and U18108 (N_18108,N_4174,N_266);
nor U18109 (N_18109,N_7037,N_4914);
and U18110 (N_18110,N_5287,N_5317);
and U18111 (N_18111,N_8612,N_1221);
and U18112 (N_18112,N_1861,N_9872);
nor U18113 (N_18113,N_1856,N_5123);
and U18114 (N_18114,N_5065,N_8373);
nor U18115 (N_18115,N_6926,N_2740);
nor U18116 (N_18116,N_4986,N_8576);
nor U18117 (N_18117,N_7322,N_3871);
or U18118 (N_18118,N_1971,N_5060);
and U18119 (N_18119,N_5322,N_2373);
or U18120 (N_18120,N_7758,N_3360);
and U18121 (N_18121,N_3095,N_1567);
or U18122 (N_18122,N_9232,N_650);
nand U18123 (N_18123,N_8036,N_1158);
and U18124 (N_18124,N_2474,N_7349);
nand U18125 (N_18125,N_3453,N_9896);
nand U18126 (N_18126,N_4573,N_4097);
nor U18127 (N_18127,N_6941,N_1372);
nand U18128 (N_18128,N_881,N_3481);
or U18129 (N_18129,N_7610,N_9223);
and U18130 (N_18130,N_5927,N_8654);
nand U18131 (N_18131,N_6124,N_7726);
and U18132 (N_18132,N_951,N_1616);
and U18133 (N_18133,N_4188,N_2827);
and U18134 (N_18134,N_9788,N_1855);
nor U18135 (N_18135,N_5216,N_6090);
nor U18136 (N_18136,N_955,N_3671);
or U18137 (N_18137,N_8141,N_5202);
or U18138 (N_18138,N_294,N_5850);
nor U18139 (N_18139,N_9444,N_6057);
nand U18140 (N_18140,N_4712,N_7545);
and U18141 (N_18141,N_3639,N_4370);
nor U18142 (N_18142,N_9565,N_8046);
and U18143 (N_18143,N_5092,N_7356);
nor U18144 (N_18144,N_1422,N_6358);
and U18145 (N_18145,N_6711,N_9587);
or U18146 (N_18146,N_2379,N_8688);
nand U18147 (N_18147,N_6970,N_4590);
and U18148 (N_18148,N_5187,N_2776);
and U18149 (N_18149,N_9319,N_169);
or U18150 (N_18150,N_5023,N_60);
and U18151 (N_18151,N_7516,N_7152);
nor U18152 (N_18152,N_4615,N_5997);
nor U18153 (N_18153,N_6407,N_4704);
or U18154 (N_18154,N_1016,N_8280);
nor U18155 (N_18155,N_8945,N_9893);
or U18156 (N_18156,N_1325,N_3439);
or U18157 (N_18157,N_545,N_7668);
nor U18158 (N_18158,N_4786,N_8817);
or U18159 (N_18159,N_5272,N_4315);
or U18160 (N_18160,N_6871,N_385);
and U18161 (N_18161,N_9572,N_7474);
nand U18162 (N_18162,N_2878,N_8093);
nand U18163 (N_18163,N_1413,N_1288);
and U18164 (N_18164,N_7409,N_3327);
nor U18165 (N_18165,N_9452,N_8161);
or U18166 (N_18166,N_9324,N_758);
nand U18167 (N_18167,N_5725,N_190);
or U18168 (N_18168,N_1891,N_5490);
or U18169 (N_18169,N_2546,N_2832);
nand U18170 (N_18170,N_8905,N_9047);
nor U18171 (N_18171,N_6405,N_199);
and U18172 (N_18172,N_5499,N_9195);
nand U18173 (N_18173,N_3735,N_7544);
nor U18174 (N_18174,N_9153,N_5441);
nor U18175 (N_18175,N_5518,N_3354);
nor U18176 (N_18176,N_9714,N_2732);
nor U18177 (N_18177,N_311,N_1525);
nor U18178 (N_18178,N_1636,N_6117);
nor U18179 (N_18179,N_8247,N_1999);
nand U18180 (N_18180,N_170,N_314);
nand U18181 (N_18181,N_2972,N_6973);
nand U18182 (N_18182,N_9641,N_8017);
and U18183 (N_18183,N_1652,N_4767);
and U18184 (N_18184,N_4708,N_1862);
or U18185 (N_18185,N_1946,N_6777);
nor U18186 (N_18186,N_3411,N_7371);
and U18187 (N_18187,N_5984,N_6252);
or U18188 (N_18188,N_5613,N_3653);
nand U18189 (N_18189,N_7786,N_2367);
nand U18190 (N_18190,N_5758,N_8638);
or U18191 (N_18191,N_6950,N_6120);
and U18192 (N_18192,N_8921,N_1614);
nor U18193 (N_18193,N_4670,N_6947);
nor U18194 (N_18194,N_1820,N_8241);
xor U18195 (N_18195,N_736,N_5621);
and U18196 (N_18196,N_4601,N_4772);
or U18197 (N_18197,N_1408,N_5516);
nor U18198 (N_18198,N_7544,N_4999);
and U18199 (N_18199,N_9768,N_6973);
nand U18200 (N_18200,N_969,N_9090);
or U18201 (N_18201,N_8906,N_6449);
nand U18202 (N_18202,N_3100,N_1107);
and U18203 (N_18203,N_5804,N_751);
or U18204 (N_18204,N_3156,N_9840);
nor U18205 (N_18205,N_3180,N_177);
nor U18206 (N_18206,N_5712,N_2338);
nand U18207 (N_18207,N_6654,N_7365);
nor U18208 (N_18208,N_8895,N_9492);
nor U18209 (N_18209,N_6334,N_2349);
nand U18210 (N_18210,N_3181,N_2769);
nand U18211 (N_18211,N_1395,N_4591);
nand U18212 (N_18212,N_6438,N_2992);
and U18213 (N_18213,N_2743,N_1753);
nand U18214 (N_18214,N_4958,N_9151);
nor U18215 (N_18215,N_3606,N_2907);
or U18216 (N_18216,N_4849,N_7034);
nand U18217 (N_18217,N_3197,N_6721);
nor U18218 (N_18218,N_3406,N_7029);
nand U18219 (N_18219,N_957,N_8526);
nor U18220 (N_18220,N_8053,N_4466);
nor U18221 (N_18221,N_1807,N_8368);
and U18222 (N_18222,N_377,N_1595);
or U18223 (N_18223,N_5503,N_1763);
or U18224 (N_18224,N_4461,N_9827);
nand U18225 (N_18225,N_959,N_2432);
or U18226 (N_18226,N_8341,N_9026);
or U18227 (N_18227,N_4279,N_8412);
nand U18228 (N_18228,N_7140,N_2164);
xnor U18229 (N_18229,N_6814,N_9409);
and U18230 (N_18230,N_8711,N_1911);
nand U18231 (N_18231,N_5817,N_7943);
and U18232 (N_18232,N_2788,N_7595);
or U18233 (N_18233,N_8560,N_1039);
nor U18234 (N_18234,N_5070,N_6193);
nand U18235 (N_18235,N_1769,N_7417);
nand U18236 (N_18236,N_2683,N_2173);
and U18237 (N_18237,N_4990,N_4061);
nor U18238 (N_18238,N_7876,N_8133);
nand U18239 (N_18239,N_5778,N_4630);
nand U18240 (N_18240,N_1201,N_4797);
or U18241 (N_18241,N_2217,N_7653);
and U18242 (N_18242,N_7304,N_3986);
nand U18243 (N_18243,N_6152,N_1136);
nand U18244 (N_18244,N_475,N_3716);
and U18245 (N_18245,N_4201,N_4460);
or U18246 (N_18246,N_3422,N_1954);
and U18247 (N_18247,N_7864,N_302);
nand U18248 (N_18248,N_4057,N_8397);
nand U18249 (N_18249,N_9177,N_9247);
and U18250 (N_18250,N_9480,N_4335);
and U18251 (N_18251,N_587,N_2071);
and U18252 (N_18252,N_6746,N_4635);
nand U18253 (N_18253,N_3748,N_5518);
nor U18254 (N_18254,N_8889,N_1357);
nor U18255 (N_18255,N_1163,N_9);
or U18256 (N_18256,N_1769,N_504);
nand U18257 (N_18257,N_9764,N_2520);
nand U18258 (N_18258,N_6828,N_7444);
and U18259 (N_18259,N_1613,N_1516);
nand U18260 (N_18260,N_2,N_2235);
nor U18261 (N_18261,N_4731,N_4671);
and U18262 (N_18262,N_6835,N_1114);
or U18263 (N_18263,N_6979,N_9054);
nand U18264 (N_18264,N_1143,N_7671);
nor U18265 (N_18265,N_7157,N_7788);
nor U18266 (N_18266,N_8174,N_1824);
nand U18267 (N_18267,N_5924,N_4618);
or U18268 (N_18268,N_6711,N_5166);
and U18269 (N_18269,N_4225,N_1906);
nand U18270 (N_18270,N_4477,N_2467);
or U18271 (N_18271,N_5628,N_5106);
nand U18272 (N_18272,N_3211,N_5185);
or U18273 (N_18273,N_5692,N_2133);
and U18274 (N_18274,N_2410,N_583);
nor U18275 (N_18275,N_5794,N_5644);
and U18276 (N_18276,N_8012,N_517);
nand U18277 (N_18277,N_5952,N_6726);
nand U18278 (N_18278,N_9528,N_5398);
nor U18279 (N_18279,N_5226,N_3199);
nand U18280 (N_18280,N_8814,N_6541);
nor U18281 (N_18281,N_7424,N_1924);
nor U18282 (N_18282,N_7530,N_5289);
nand U18283 (N_18283,N_1617,N_8870);
or U18284 (N_18284,N_5395,N_1881);
or U18285 (N_18285,N_6352,N_9132);
and U18286 (N_18286,N_4586,N_1547);
nor U18287 (N_18287,N_3935,N_5031);
and U18288 (N_18288,N_8670,N_1330);
or U18289 (N_18289,N_4012,N_4765);
and U18290 (N_18290,N_1796,N_8599);
or U18291 (N_18291,N_1185,N_8202);
nor U18292 (N_18292,N_416,N_8981);
nor U18293 (N_18293,N_5744,N_230);
or U18294 (N_18294,N_2108,N_4330);
nor U18295 (N_18295,N_9204,N_2848);
and U18296 (N_18296,N_7729,N_1331);
or U18297 (N_18297,N_3735,N_8489);
nor U18298 (N_18298,N_5150,N_4818);
nor U18299 (N_18299,N_69,N_4986);
nand U18300 (N_18300,N_4064,N_6829);
nor U18301 (N_18301,N_2063,N_1851);
or U18302 (N_18302,N_7895,N_3674);
nor U18303 (N_18303,N_4143,N_8699);
nand U18304 (N_18304,N_8013,N_938);
and U18305 (N_18305,N_7127,N_8431);
nand U18306 (N_18306,N_1941,N_491);
and U18307 (N_18307,N_589,N_7125);
xnor U18308 (N_18308,N_7065,N_7907);
nor U18309 (N_18309,N_1701,N_517);
nor U18310 (N_18310,N_1176,N_6476);
nand U18311 (N_18311,N_8656,N_530);
or U18312 (N_18312,N_4742,N_7555);
or U18313 (N_18313,N_5388,N_4095);
and U18314 (N_18314,N_2540,N_6657);
or U18315 (N_18315,N_7179,N_7317);
nor U18316 (N_18316,N_1494,N_2178);
nor U18317 (N_18317,N_8372,N_8739);
or U18318 (N_18318,N_3965,N_8991);
nor U18319 (N_18319,N_142,N_2749);
nand U18320 (N_18320,N_220,N_9371);
nor U18321 (N_18321,N_6977,N_2157);
nand U18322 (N_18322,N_5981,N_4831);
nor U18323 (N_18323,N_6190,N_6004);
nand U18324 (N_18324,N_271,N_3020);
and U18325 (N_18325,N_3493,N_4247);
nor U18326 (N_18326,N_1394,N_1890);
or U18327 (N_18327,N_2272,N_188);
and U18328 (N_18328,N_1171,N_5587);
and U18329 (N_18329,N_8692,N_4366);
nor U18330 (N_18330,N_3373,N_5249);
nor U18331 (N_18331,N_4161,N_5287);
and U18332 (N_18332,N_8617,N_5654);
and U18333 (N_18333,N_2333,N_1840);
and U18334 (N_18334,N_2698,N_5080);
or U18335 (N_18335,N_8948,N_2559);
or U18336 (N_18336,N_3296,N_1648);
and U18337 (N_18337,N_8533,N_2263);
or U18338 (N_18338,N_6179,N_2327);
or U18339 (N_18339,N_1110,N_8139);
and U18340 (N_18340,N_9318,N_5072);
or U18341 (N_18341,N_1904,N_1166);
and U18342 (N_18342,N_9858,N_4915);
nand U18343 (N_18343,N_7692,N_8230);
nor U18344 (N_18344,N_4199,N_8910);
and U18345 (N_18345,N_3565,N_7495);
or U18346 (N_18346,N_3671,N_8517);
nand U18347 (N_18347,N_3062,N_6047);
nand U18348 (N_18348,N_8847,N_4820);
nor U18349 (N_18349,N_4634,N_5886);
nand U18350 (N_18350,N_3321,N_2610);
or U18351 (N_18351,N_2531,N_9320);
or U18352 (N_18352,N_6592,N_2526);
nand U18353 (N_18353,N_5769,N_2834);
nand U18354 (N_18354,N_6459,N_1365);
or U18355 (N_18355,N_9542,N_2144);
or U18356 (N_18356,N_903,N_1390);
or U18357 (N_18357,N_6336,N_6657);
and U18358 (N_18358,N_4265,N_4861);
nand U18359 (N_18359,N_2115,N_6923);
and U18360 (N_18360,N_9363,N_6416);
nor U18361 (N_18361,N_9425,N_9226);
nand U18362 (N_18362,N_8796,N_6872);
nor U18363 (N_18363,N_2881,N_241);
or U18364 (N_18364,N_5744,N_2808);
nor U18365 (N_18365,N_2369,N_7669);
and U18366 (N_18366,N_3101,N_3765);
nor U18367 (N_18367,N_6157,N_5665);
nand U18368 (N_18368,N_8680,N_7515);
and U18369 (N_18369,N_5234,N_4223);
and U18370 (N_18370,N_5442,N_5976);
xnor U18371 (N_18371,N_7323,N_2482);
and U18372 (N_18372,N_2819,N_6774);
or U18373 (N_18373,N_7282,N_94);
or U18374 (N_18374,N_8949,N_1059);
nor U18375 (N_18375,N_6574,N_3018);
or U18376 (N_18376,N_8562,N_5414);
or U18377 (N_18377,N_3130,N_226);
nand U18378 (N_18378,N_3123,N_7132);
or U18379 (N_18379,N_1229,N_8418);
or U18380 (N_18380,N_4129,N_4355);
nor U18381 (N_18381,N_110,N_7157);
and U18382 (N_18382,N_3245,N_8324);
nor U18383 (N_18383,N_123,N_741);
and U18384 (N_18384,N_8310,N_2210);
and U18385 (N_18385,N_9980,N_1278);
nand U18386 (N_18386,N_9355,N_3203);
nor U18387 (N_18387,N_7417,N_5940);
or U18388 (N_18388,N_1590,N_5252);
or U18389 (N_18389,N_9095,N_4963);
nor U18390 (N_18390,N_9453,N_5174);
nor U18391 (N_18391,N_9211,N_723);
nor U18392 (N_18392,N_5088,N_1275);
or U18393 (N_18393,N_2063,N_5345);
or U18394 (N_18394,N_4713,N_4847);
or U18395 (N_18395,N_7022,N_7137);
nor U18396 (N_18396,N_6987,N_9602);
or U18397 (N_18397,N_6029,N_5408);
and U18398 (N_18398,N_7306,N_820);
nand U18399 (N_18399,N_8592,N_5186);
nand U18400 (N_18400,N_8782,N_5706);
or U18401 (N_18401,N_352,N_3208);
nand U18402 (N_18402,N_6036,N_9473);
nor U18403 (N_18403,N_6394,N_7496);
nand U18404 (N_18404,N_3458,N_1906);
nand U18405 (N_18405,N_6159,N_9854);
nand U18406 (N_18406,N_5719,N_1031);
and U18407 (N_18407,N_8357,N_6662);
and U18408 (N_18408,N_3398,N_823);
and U18409 (N_18409,N_3772,N_31);
nor U18410 (N_18410,N_479,N_5507);
nor U18411 (N_18411,N_4819,N_1421);
and U18412 (N_18412,N_9410,N_4396);
nor U18413 (N_18413,N_7354,N_9854);
nor U18414 (N_18414,N_4965,N_8173);
nor U18415 (N_18415,N_2003,N_6719);
or U18416 (N_18416,N_7643,N_8726);
nand U18417 (N_18417,N_4305,N_5869);
nor U18418 (N_18418,N_9488,N_9691);
and U18419 (N_18419,N_8132,N_2785);
nor U18420 (N_18420,N_3666,N_9849);
nor U18421 (N_18421,N_4495,N_6747);
nand U18422 (N_18422,N_5041,N_5155);
nor U18423 (N_18423,N_9100,N_4762);
nor U18424 (N_18424,N_5939,N_4333);
nand U18425 (N_18425,N_5457,N_3256);
or U18426 (N_18426,N_3146,N_9481);
nand U18427 (N_18427,N_3012,N_959);
or U18428 (N_18428,N_2693,N_9918);
nor U18429 (N_18429,N_9328,N_2585);
or U18430 (N_18430,N_947,N_129);
or U18431 (N_18431,N_8962,N_4512);
nor U18432 (N_18432,N_8820,N_6175);
or U18433 (N_18433,N_3827,N_8590);
nand U18434 (N_18434,N_524,N_9525);
nor U18435 (N_18435,N_9351,N_1601);
nor U18436 (N_18436,N_3634,N_3384);
nand U18437 (N_18437,N_6011,N_3966);
and U18438 (N_18438,N_557,N_2602);
or U18439 (N_18439,N_7325,N_1313);
or U18440 (N_18440,N_2070,N_8468);
and U18441 (N_18441,N_6605,N_153);
nor U18442 (N_18442,N_168,N_4977);
nor U18443 (N_18443,N_5798,N_6445);
and U18444 (N_18444,N_2485,N_4891);
or U18445 (N_18445,N_2538,N_8299);
nand U18446 (N_18446,N_578,N_2016);
or U18447 (N_18447,N_7134,N_5539);
nor U18448 (N_18448,N_5252,N_5405);
nor U18449 (N_18449,N_8755,N_3495);
nand U18450 (N_18450,N_1601,N_7443);
nand U18451 (N_18451,N_9343,N_3211);
nand U18452 (N_18452,N_8728,N_5072);
nor U18453 (N_18453,N_1071,N_6652);
or U18454 (N_18454,N_4084,N_1581);
nand U18455 (N_18455,N_9506,N_4777);
or U18456 (N_18456,N_7625,N_9687);
or U18457 (N_18457,N_2410,N_9125);
nor U18458 (N_18458,N_2679,N_4143);
and U18459 (N_18459,N_3750,N_9151);
or U18460 (N_18460,N_9597,N_9479);
or U18461 (N_18461,N_9567,N_1496);
nor U18462 (N_18462,N_1313,N_270);
nor U18463 (N_18463,N_5318,N_5276);
and U18464 (N_18464,N_6331,N_9074);
or U18465 (N_18465,N_8527,N_4191);
and U18466 (N_18466,N_2263,N_9639);
and U18467 (N_18467,N_6054,N_2908);
nor U18468 (N_18468,N_9528,N_2179);
nand U18469 (N_18469,N_21,N_1414);
nand U18470 (N_18470,N_4828,N_9199);
nand U18471 (N_18471,N_5085,N_6168);
nand U18472 (N_18472,N_5171,N_3250);
xnor U18473 (N_18473,N_9812,N_8738);
nor U18474 (N_18474,N_8825,N_6351);
or U18475 (N_18475,N_5160,N_5055);
and U18476 (N_18476,N_9035,N_3490);
nand U18477 (N_18477,N_1421,N_3248);
or U18478 (N_18478,N_8144,N_9594);
nor U18479 (N_18479,N_1773,N_9866);
nand U18480 (N_18480,N_1649,N_785);
nand U18481 (N_18481,N_4517,N_6064);
nor U18482 (N_18482,N_6109,N_946);
and U18483 (N_18483,N_3719,N_6352);
or U18484 (N_18484,N_3338,N_2102);
and U18485 (N_18485,N_8575,N_7163);
or U18486 (N_18486,N_3325,N_7290);
nand U18487 (N_18487,N_7211,N_6519);
nand U18488 (N_18488,N_9271,N_2007);
nor U18489 (N_18489,N_373,N_3788);
nor U18490 (N_18490,N_1610,N_3060);
nor U18491 (N_18491,N_1503,N_5143);
nor U18492 (N_18492,N_5136,N_3015);
and U18493 (N_18493,N_3304,N_3357);
and U18494 (N_18494,N_70,N_9474);
or U18495 (N_18495,N_6574,N_3780);
and U18496 (N_18496,N_1767,N_8974);
nand U18497 (N_18497,N_742,N_3760);
and U18498 (N_18498,N_2689,N_7860);
nand U18499 (N_18499,N_9262,N_7194);
and U18500 (N_18500,N_4080,N_1966);
and U18501 (N_18501,N_1568,N_7183);
nand U18502 (N_18502,N_8787,N_2960);
nand U18503 (N_18503,N_2639,N_6578);
and U18504 (N_18504,N_225,N_5360);
nand U18505 (N_18505,N_4147,N_9790);
nand U18506 (N_18506,N_2419,N_4756);
nor U18507 (N_18507,N_1130,N_1403);
or U18508 (N_18508,N_1738,N_4583);
xor U18509 (N_18509,N_1133,N_255);
and U18510 (N_18510,N_6430,N_1821);
or U18511 (N_18511,N_5107,N_8038);
and U18512 (N_18512,N_8701,N_4550);
or U18513 (N_18513,N_8023,N_9366);
nor U18514 (N_18514,N_8173,N_2487);
and U18515 (N_18515,N_9594,N_7287);
or U18516 (N_18516,N_2266,N_7374);
or U18517 (N_18517,N_4263,N_7665);
and U18518 (N_18518,N_150,N_7524);
nor U18519 (N_18519,N_9921,N_1561);
or U18520 (N_18520,N_6059,N_6816);
and U18521 (N_18521,N_804,N_7331);
or U18522 (N_18522,N_3062,N_7075);
nor U18523 (N_18523,N_7614,N_6839);
and U18524 (N_18524,N_2297,N_9277);
nor U18525 (N_18525,N_8933,N_871);
and U18526 (N_18526,N_2713,N_8925);
or U18527 (N_18527,N_741,N_5009);
nand U18528 (N_18528,N_2008,N_8713);
and U18529 (N_18529,N_8757,N_6934);
or U18530 (N_18530,N_2091,N_732);
nor U18531 (N_18531,N_5969,N_2632);
or U18532 (N_18532,N_6725,N_4633);
nor U18533 (N_18533,N_3307,N_1624);
nand U18534 (N_18534,N_719,N_9045);
nand U18535 (N_18535,N_4313,N_1171);
or U18536 (N_18536,N_1914,N_6323);
or U18537 (N_18537,N_956,N_2736);
nand U18538 (N_18538,N_7366,N_1696);
and U18539 (N_18539,N_5397,N_2975);
nor U18540 (N_18540,N_3632,N_1788);
nand U18541 (N_18541,N_6776,N_6084);
nor U18542 (N_18542,N_1024,N_528);
nand U18543 (N_18543,N_6297,N_9862);
xnor U18544 (N_18544,N_2973,N_1172);
and U18545 (N_18545,N_8569,N_5365);
nor U18546 (N_18546,N_487,N_6174);
and U18547 (N_18547,N_3312,N_8507);
or U18548 (N_18548,N_7497,N_3175);
nor U18549 (N_18549,N_6368,N_8914);
nand U18550 (N_18550,N_8675,N_8442);
and U18551 (N_18551,N_1370,N_9772);
and U18552 (N_18552,N_9605,N_3001);
nor U18553 (N_18553,N_9155,N_1449);
nand U18554 (N_18554,N_6799,N_5879);
and U18555 (N_18555,N_9440,N_3207);
nand U18556 (N_18556,N_4486,N_3922);
nand U18557 (N_18557,N_34,N_9230);
nand U18558 (N_18558,N_4431,N_6556);
nor U18559 (N_18559,N_24,N_6471);
xor U18560 (N_18560,N_9518,N_277);
and U18561 (N_18561,N_9886,N_5273);
or U18562 (N_18562,N_5073,N_5723);
nor U18563 (N_18563,N_3382,N_1721);
and U18564 (N_18564,N_1643,N_390);
and U18565 (N_18565,N_8993,N_8681);
nor U18566 (N_18566,N_9833,N_9641);
or U18567 (N_18567,N_3266,N_4838);
nor U18568 (N_18568,N_7716,N_8936);
nand U18569 (N_18569,N_6932,N_1839);
and U18570 (N_18570,N_3509,N_2542);
nand U18571 (N_18571,N_8827,N_8472);
and U18572 (N_18572,N_6714,N_4966);
nand U18573 (N_18573,N_7840,N_3359);
nor U18574 (N_18574,N_5984,N_7476);
nor U18575 (N_18575,N_2448,N_6060);
nor U18576 (N_18576,N_1722,N_2982);
nor U18577 (N_18577,N_2782,N_9898);
or U18578 (N_18578,N_7397,N_6567);
nor U18579 (N_18579,N_8288,N_7565);
nand U18580 (N_18580,N_7874,N_8408);
nor U18581 (N_18581,N_6005,N_2130);
nor U18582 (N_18582,N_9846,N_7365);
or U18583 (N_18583,N_6527,N_6484);
nand U18584 (N_18584,N_5711,N_1062);
and U18585 (N_18585,N_5626,N_7999);
nand U18586 (N_18586,N_9332,N_5433);
nand U18587 (N_18587,N_4541,N_6261);
nor U18588 (N_18588,N_311,N_2068);
and U18589 (N_18589,N_2935,N_5203);
nor U18590 (N_18590,N_1864,N_5661);
nor U18591 (N_18591,N_7106,N_1389);
or U18592 (N_18592,N_5870,N_9503);
and U18593 (N_18593,N_1916,N_1760);
nor U18594 (N_18594,N_1366,N_7261);
nand U18595 (N_18595,N_4512,N_8091);
and U18596 (N_18596,N_1129,N_5361);
nand U18597 (N_18597,N_1596,N_4439);
or U18598 (N_18598,N_170,N_5932);
nor U18599 (N_18599,N_6374,N_228);
nor U18600 (N_18600,N_8320,N_490);
nand U18601 (N_18601,N_4098,N_8812);
nor U18602 (N_18602,N_1726,N_5408);
and U18603 (N_18603,N_1316,N_717);
or U18604 (N_18604,N_7534,N_5101);
or U18605 (N_18605,N_9071,N_7420);
nor U18606 (N_18606,N_3909,N_7894);
or U18607 (N_18607,N_1129,N_9807);
nor U18608 (N_18608,N_6070,N_1756);
nand U18609 (N_18609,N_5885,N_2988);
nand U18610 (N_18610,N_9958,N_4299);
nand U18611 (N_18611,N_6222,N_6181);
nand U18612 (N_18612,N_505,N_5455);
nor U18613 (N_18613,N_3736,N_5900);
nor U18614 (N_18614,N_7276,N_2702);
nor U18615 (N_18615,N_8761,N_5352);
and U18616 (N_18616,N_534,N_4648);
nand U18617 (N_18617,N_5878,N_1902);
or U18618 (N_18618,N_4542,N_4352);
or U18619 (N_18619,N_273,N_7517);
or U18620 (N_18620,N_2631,N_1477);
and U18621 (N_18621,N_6034,N_6936);
or U18622 (N_18622,N_3946,N_9665);
nor U18623 (N_18623,N_4674,N_8087);
or U18624 (N_18624,N_873,N_6488);
nand U18625 (N_18625,N_6309,N_3255);
and U18626 (N_18626,N_5015,N_9836);
or U18627 (N_18627,N_2809,N_4270);
or U18628 (N_18628,N_6619,N_8602);
nand U18629 (N_18629,N_8919,N_8085);
or U18630 (N_18630,N_5351,N_1123);
xnor U18631 (N_18631,N_2015,N_8300);
nand U18632 (N_18632,N_3137,N_5544);
nor U18633 (N_18633,N_6701,N_4706);
and U18634 (N_18634,N_2546,N_5993);
or U18635 (N_18635,N_7003,N_7102);
nand U18636 (N_18636,N_5879,N_5924);
nor U18637 (N_18637,N_5307,N_3741);
nor U18638 (N_18638,N_927,N_3547);
xor U18639 (N_18639,N_2485,N_7256);
and U18640 (N_18640,N_5547,N_3497);
nand U18641 (N_18641,N_3868,N_6672);
nor U18642 (N_18642,N_9375,N_4142);
and U18643 (N_18643,N_8069,N_7667);
or U18644 (N_18644,N_3066,N_6753);
or U18645 (N_18645,N_153,N_4345);
or U18646 (N_18646,N_902,N_7093);
nand U18647 (N_18647,N_5152,N_1320);
and U18648 (N_18648,N_3755,N_3758);
nor U18649 (N_18649,N_9486,N_2258);
and U18650 (N_18650,N_485,N_6988);
nor U18651 (N_18651,N_534,N_2872);
or U18652 (N_18652,N_272,N_4964);
or U18653 (N_18653,N_582,N_7514);
nand U18654 (N_18654,N_9213,N_4368);
nor U18655 (N_18655,N_312,N_3405);
and U18656 (N_18656,N_1442,N_8048);
nor U18657 (N_18657,N_2989,N_178);
nand U18658 (N_18658,N_6252,N_4964);
and U18659 (N_18659,N_6255,N_6846);
and U18660 (N_18660,N_9117,N_4023);
or U18661 (N_18661,N_1563,N_3419);
or U18662 (N_18662,N_951,N_2173);
and U18663 (N_18663,N_1014,N_6573);
and U18664 (N_18664,N_6143,N_1760);
and U18665 (N_18665,N_7025,N_3992);
nor U18666 (N_18666,N_8013,N_5919);
and U18667 (N_18667,N_1184,N_5797);
nand U18668 (N_18668,N_4685,N_6574);
nor U18669 (N_18669,N_9272,N_5694);
nor U18670 (N_18670,N_5013,N_8330);
nor U18671 (N_18671,N_5236,N_6160);
nand U18672 (N_18672,N_1349,N_951);
and U18673 (N_18673,N_3647,N_6356);
nor U18674 (N_18674,N_118,N_5123);
nor U18675 (N_18675,N_9715,N_7085);
nand U18676 (N_18676,N_3306,N_7759);
nand U18677 (N_18677,N_1232,N_3636);
or U18678 (N_18678,N_9185,N_9918);
or U18679 (N_18679,N_3309,N_2101);
or U18680 (N_18680,N_8571,N_9321);
nor U18681 (N_18681,N_1428,N_8804);
nand U18682 (N_18682,N_2850,N_2225);
nand U18683 (N_18683,N_4599,N_8011);
or U18684 (N_18684,N_6684,N_5826);
nor U18685 (N_18685,N_9132,N_4960);
nor U18686 (N_18686,N_314,N_4864);
or U18687 (N_18687,N_5326,N_6136);
and U18688 (N_18688,N_9548,N_8783);
and U18689 (N_18689,N_8574,N_3409);
or U18690 (N_18690,N_195,N_7621);
nor U18691 (N_18691,N_3948,N_8600);
nor U18692 (N_18692,N_4838,N_3723);
nand U18693 (N_18693,N_7120,N_7740);
xor U18694 (N_18694,N_3130,N_3589);
or U18695 (N_18695,N_579,N_5348);
nor U18696 (N_18696,N_4946,N_236);
or U18697 (N_18697,N_5833,N_4764);
nor U18698 (N_18698,N_9104,N_1846);
or U18699 (N_18699,N_5991,N_8400);
nor U18700 (N_18700,N_2110,N_140);
nor U18701 (N_18701,N_9801,N_9059);
nand U18702 (N_18702,N_5194,N_9930);
or U18703 (N_18703,N_9727,N_9768);
or U18704 (N_18704,N_2412,N_5571);
nand U18705 (N_18705,N_4238,N_4763);
nor U18706 (N_18706,N_2296,N_2494);
nor U18707 (N_18707,N_2915,N_2894);
nand U18708 (N_18708,N_8695,N_1707);
and U18709 (N_18709,N_1980,N_8738);
xor U18710 (N_18710,N_5751,N_415);
or U18711 (N_18711,N_4513,N_6900);
and U18712 (N_18712,N_4939,N_6014);
nor U18713 (N_18713,N_6960,N_2765);
or U18714 (N_18714,N_6998,N_8118);
nor U18715 (N_18715,N_5797,N_443);
or U18716 (N_18716,N_3478,N_5637);
xnor U18717 (N_18717,N_622,N_8906);
and U18718 (N_18718,N_9711,N_895);
nand U18719 (N_18719,N_5795,N_671);
and U18720 (N_18720,N_7488,N_316);
nor U18721 (N_18721,N_9494,N_6551);
nand U18722 (N_18722,N_9674,N_3056);
and U18723 (N_18723,N_7818,N_4515);
or U18724 (N_18724,N_1288,N_1746);
nand U18725 (N_18725,N_9641,N_9984);
nand U18726 (N_18726,N_6497,N_8267);
or U18727 (N_18727,N_7797,N_4117);
or U18728 (N_18728,N_7672,N_7045);
and U18729 (N_18729,N_4519,N_3040);
or U18730 (N_18730,N_7935,N_8397);
and U18731 (N_18731,N_358,N_9439);
nor U18732 (N_18732,N_8370,N_402);
and U18733 (N_18733,N_2456,N_9913);
and U18734 (N_18734,N_8406,N_6981);
and U18735 (N_18735,N_9706,N_6286);
nor U18736 (N_18736,N_5098,N_5309);
nor U18737 (N_18737,N_2595,N_7587);
and U18738 (N_18738,N_9311,N_6791);
nor U18739 (N_18739,N_1492,N_8413);
or U18740 (N_18740,N_9515,N_1768);
and U18741 (N_18741,N_7336,N_5025);
nor U18742 (N_18742,N_1067,N_3743);
or U18743 (N_18743,N_4928,N_8371);
and U18744 (N_18744,N_3891,N_610);
and U18745 (N_18745,N_8245,N_5529);
and U18746 (N_18746,N_1116,N_6163);
nand U18747 (N_18747,N_5273,N_2194);
nand U18748 (N_18748,N_1148,N_4086);
and U18749 (N_18749,N_9955,N_4930);
and U18750 (N_18750,N_2449,N_7298);
nor U18751 (N_18751,N_3813,N_9495);
nand U18752 (N_18752,N_2221,N_1334);
nand U18753 (N_18753,N_5926,N_9662);
and U18754 (N_18754,N_9359,N_3464);
nand U18755 (N_18755,N_5251,N_2050);
nor U18756 (N_18756,N_6024,N_7366);
and U18757 (N_18757,N_4005,N_4479);
nand U18758 (N_18758,N_4164,N_3946);
nor U18759 (N_18759,N_8697,N_557);
and U18760 (N_18760,N_7292,N_2911);
or U18761 (N_18761,N_1919,N_1845);
nor U18762 (N_18762,N_8795,N_831);
and U18763 (N_18763,N_7254,N_9579);
or U18764 (N_18764,N_8588,N_4466);
and U18765 (N_18765,N_8084,N_4823);
or U18766 (N_18766,N_1222,N_3460);
nor U18767 (N_18767,N_6305,N_1209);
nor U18768 (N_18768,N_5086,N_2690);
nand U18769 (N_18769,N_4644,N_2280);
nor U18770 (N_18770,N_777,N_1208);
or U18771 (N_18771,N_7815,N_6755);
nand U18772 (N_18772,N_9726,N_6884);
nand U18773 (N_18773,N_3145,N_2150);
xor U18774 (N_18774,N_1074,N_8487);
and U18775 (N_18775,N_369,N_7208);
or U18776 (N_18776,N_4116,N_4668);
or U18777 (N_18777,N_197,N_1873);
and U18778 (N_18778,N_9954,N_8788);
xor U18779 (N_18779,N_2993,N_565);
nor U18780 (N_18780,N_4026,N_1784);
and U18781 (N_18781,N_2654,N_3383);
or U18782 (N_18782,N_2721,N_467);
nor U18783 (N_18783,N_5964,N_1183);
or U18784 (N_18784,N_6960,N_3497);
or U18785 (N_18785,N_9358,N_7736);
and U18786 (N_18786,N_3382,N_499);
or U18787 (N_18787,N_3586,N_818);
or U18788 (N_18788,N_215,N_8740);
or U18789 (N_18789,N_7990,N_6682);
nand U18790 (N_18790,N_751,N_7535);
and U18791 (N_18791,N_3900,N_2889);
nor U18792 (N_18792,N_2939,N_7055);
and U18793 (N_18793,N_9886,N_5962);
nand U18794 (N_18794,N_1711,N_5746);
and U18795 (N_18795,N_6719,N_8932);
nor U18796 (N_18796,N_8492,N_4912);
or U18797 (N_18797,N_7984,N_3581);
or U18798 (N_18798,N_7974,N_6766);
or U18799 (N_18799,N_9255,N_1019);
nand U18800 (N_18800,N_9705,N_3445);
nand U18801 (N_18801,N_4836,N_339);
or U18802 (N_18802,N_4166,N_2081);
nand U18803 (N_18803,N_7270,N_4726);
nor U18804 (N_18804,N_967,N_1284);
and U18805 (N_18805,N_3899,N_5202);
nand U18806 (N_18806,N_342,N_1472);
or U18807 (N_18807,N_1898,N_4063);
and U18808 (N_18808,N_1939,N_8868);
nand U18809 (N_18809,N_8912,N_2763);
nor U18810 (N_18810,N_1692,N_5220);
and U18811 (N_18811,N_2346,N_3353);
and U18812 (N_18812,N_6958,N_2519);
or U18813 (N_18813,N_1065,N_5373);
or U18814 (N_18814,N_7812,N_9922);
and U18815 (N_18815,N_1763,N_1908);
and U18816 (N_18816,N_4582,N_8489);
and U18817 (N_18817,N_6292,N_6455);
nand U18818 (N_18818,N_1068,N_7053);
and U18819 (N_18819,N_4053,N_9507);
or U18820 (N_18820,N_5736,N_9352);
or U18821 (N_18821,N_6585,N_1113);
or U18822 (N_18822,N_8586,N_5798);
or U18823 (N_18823,N_9473,N_4083);
or U18824 (N_18824,N_1298,N_1829);
or U18825 (N_18825,N_1556,N_6919);
and U18826 (N_18826,N_9584,N_2105);
or U18827 (N_18827,N_1210,N_1031);
and U18828 (N_18828,N_5013,N_8139);
or U18829 (N_18829,N_9419,N_3497);
nand U18830 (N_18830,N_7287,N_8874);
nor U18831 (N_18831,N_5137,N_2838);
nor U18832 (N_18832,N_7685,N_9102);
nor U18833 (N_18833,N_143,N_8006);
and U18834 (N_18834,N_6967,N_5845);
and U18835 (N_18835,N_3883,N_2359);
nor U18836 (N_18836,N_4033,N_2617);
or U18837 (N_18837,N_2621,N_2645);
or U18838 (N_18838,N_3176,N_1211);
nand U18839 (N_18839,N_7293,N_9900);
nand U18840 (N_18840,N_5437,N_8465);
or U18841 (N_18841,N_2400,N_7688);
nor U18842 (N_18842,N_1551,N_7108);
or U18843 (N_18843,N_4715,N_718);
nand U18844 (N_18844,N_7468,N_7276);
nor U18845 (N_18845,N_7098,N_7243);
and U18846 (N_18846,N_3578,N_5838);
nand U18847 (N_18847,N_8559,N_8819);
or U18848 (N_18848,N_458,N_1711);
or U18849 (N_18849,N_73,N_8288);
nand U18850 (N_18850,N_7482,N_9928);
nor U18851 (N_18851,N_3652,N_698);
and U18852 (N_18852,N_4747,N_3064);
or U18853 (N_18853,N_1943,N_5268);
nor U18854 (N_18854,N_9687,N_7955);
nor U18855 (N_18855,N_2818,N_2667);
nor U18856 (N_18856,N_9517,N_2049);
and U18857 (N_18857,N_1936,N_3134);
nor U18858 (N_18858,N_5713,N_5440);
or U18859 (N_18859,N_6980,N_6793);
or U18860 (N_18860,N_4417,N_9664);
or U18861 (N_18861,N_7966,N_1153);
and U18862 (N_18862,N_6926,N_5662);
nor U18863 (N_18863,N_2878,N_5479);
and U18864 (N_18864,N_5525,N_1892);
nor U18865 (N_18865,N_2991,N_4986);
and U18866 (N_18866,N_1243,N_1455);
nand U18867 (N_18867,N_6691,N_4092);
or U18868 (N_18868,N_5942,N_9652);
nand U18869 (N_18869,N_8747,N_8842);
nor U18870 (N_18870,N_3058,N_5080);
and U18871 (N_18871,N_5446,N_780);
nand U18872 (N_18872,N_8607,N_6829);
and U18873 (N_18873,N_4703,N_6798);
nand U18874 (N_18874,N_4593,N_98);
nor U18875 (N_18875,N_8419,N_9355);
and U18876 (N_18876,N_5036,N_5179);
and U18877 (N_18877,N_8396,N_4002);
nor U18878 (N_18878,N_9280,N_8385);
nor U18879 (N_18879,N_9035,N_4693);
nor U18880 (N_18880,N_1562,N_7241);
or U18881 (N_18881,N_5982,N_8773);
nand U18882 (N_18882,N_3126,N_4742);
nor U18883 (N_18883,N_5650,N_1846);
nor U18884 (N_18884,N_3254,N_2992);
nor U18885 (N_18885,N_7464,N_4402);
nor U18886 (N_18886,N_510,N_9643);
nand U18887 (N_18887,N_6117,N_1018);
nand U18888 (N_18888,N_4638,N_9182);
nor U18889 (N_18889,N_3760,N_8499);
or U18890 (N_18890,N_548,N_3371);
and U18891 (N_18891,N_5225,N_8174);
and U18892 (N_18892,N_5134,N_5818);
nor U18893 (N_18893,N_2823,N_5807);
and U18894 (N_18894,N_3741,N_608);
or U18895 (N_18895,N_6823,N_8603);
nor U18896 (N_18896,N_559,N_442);
and U18897 (N_18897,N_455,N_9450);
or U18898 (N_18898,N_4727,N_6007);
or U18899 (N_18899,N_7973,N_8540);
nand U18900 (N_18900,N_3834,N_3496);
or U18901 (N_18901,N_1831,N_9506);
nand U18902 (N_18902,N_3289,N_5081);
nand U18903 (N_18903,N_4676,N_8551);
nand U18904 (N_18904,N_5524,N_1470);
nor U18905 (N_18905,N_634,N_7701);
xnor U18906 (N_18906,N_3443,N_3890);
nand U18907 (N_18907,N_1867,N_2365);
and U18908 (N_18908,N_5038,N_9310);
nand U18909 (N_18909,N_3168,N_9693);
and U18910 (N_18910,N_2822,N_8872);
nand U18911 (N_18911,N_7869,N_8172);
nand U18912 (N_18912,N_6895,N_2173);
and U18913 (N_18913,N_1414,N_6893);
and U18914 (N_18914,N_9861,N_6687);
nor U18915 (N_18915,N_5482,N_5217);
nor U18916 (N_18916,N_2783,N_8403);
or U18917 (N_18917,N_1013,N_4095);
or U18918 (N_18918,N_2004,N_9150);
and U18919 (N_18919,N_8830,N_4341);
and U18920 (N_18920,N_4038,N_1965);
and U18921 (N_18921,N_9264,N_6458);
xnor U18922 (N_18922,N_9564,N_9095);
and U18923 (N_18923,N_376,N_584);
or U18924 (N_18924,N_6333,N_6149);
nand U18925 (N_18925,N_5852,N_2960);
and U18926 (N_18926,N_7255,N_2627);
or U18927 (N_18927,N_4346,N_7507);
nand U18928 (N_18928,N_5860,N_1361);
nand U18929 (N_18929,N_3189,N_9093);
nor U18930 (N_18930,N_4672,N_4194);
or U18931 (N_18931,N_7273,N_2711);
nand U18932 (N_18932,N_4159,N_8193);
nand U18933 (N_18933,N_5372,N_3588);
nand U18934 (N_18934,N_7134,N_8483);
nor U18935 (N_18935,N_2267,N_5833);
nand U18936 (N_18936,N_8342,N_7887);
or U18937 (N_18937,N_2771,N_4000);
and U18938 (N_18938,N_2964,N_3517);
nor U18939 (N_18939,N_8101,N_1958);
or U18940 (N_18940,N_7111,N_1692);
or U18941 (N_18941,N_4991,N_592);
or U18942 (N_18942,N_7580,N_4366);
or U18943 (N_18943,N_5779,N_8334);
nand U18944 (N_18944,N_6112,N_7448);
or U18945 (N_18945,N_2706,N_8686);
or U18946 (N_18946,N_872,N_825);
nor U18947 (N_18947,N_8342,N_3712);
nand U18948 (N_18948,N_6329,N_2745);
or U18949 (N_18949,N_3934,N_5408);
and U18950 (N_18950,N_5812,N_7170);
nand U18951 (N_18951,N_2827,N_8823);
nor U18952 (N_18952,N_2817,N_2021);
or U18953 (N_18953,N_3398,N_3619);
nor U18954 (N_18954,N_8861,N_1165);
xnor U18955 (N_18955,N_7926,N_5421);
nand U18956 (N_18956,N_6126,N_7731);
and U18957 (N_18957,N_1445,N_360);
and U18958 (N_18958,N_5840,N_8846);
nor U18959 (N_18959,N_6497,N_3486);
nor U18960 (N_18960,N_2928,N_550);
and U18961 (N_18961,N_4272,N_5522);
or U18962 (N_18962,N_161,N_7553);
nand U18963 (N_18963,N_3334,N_1755);
nor U18964 (N_18964,N_6968,N_3802);
nor U18965 (N_18965,N_7534,N_1034);
nand U18966 (N_18966,N_6690,N_3480);
nand U18967 (N_18967,N_5702,N_9251);
nor U18968 (N_18968,N_5277,N_323);
or U18969 (N_18969,N_2185,N_5052);
nand U18970 (N_18970,N_8990,N_3419);
or U18971 (N_18971,N_623,N_6802);
or U18972 (N_18972,N_684,N_1609);
and U18973 (N_18973,N_1578,N_5967);
or U18974 (N_18974,N_8676,N_7250);
nor U18975 (N_18975,N_2618,N_1442);
and U18976 (N_18976,N_2705,N_6664);
and U18977 (N_18977,N_7835,N_771);
or U18978 (N_18978,N_5371,N_7942);
nand U18979 (N_18979,N_4844,N_2843);
nor U18980 (N_18980,N_6213,N_5088);
and U18981 (N_18981,N_7369,N_9094);
nand U18982 (N_18982,N_2355,N_2593);
nand U18983 (N_18983,N_5732,N_7721);
nand U18984 (N_18984,N_3282,N_7752);
and U18985 (N_18985,N_9386,N_3796);
or U18986 (N_18986,N_7431,N_8461);
and U18987 (N_18987,N_1717,N_1879);
or U18988 (N_18988,N_4848,N_9606);
nand U18989 (N_18989,N_829,N_4229);
nand U18990 (N_18990,N_3617,N_9578);
and U18991 (N_18991,N_9833,N_4720);
or U18992 (N_18992,N_6861,N_869);
or U18993 (N_18993,N_6900,N_6508);
nand U18994 (N_18994,N_1791,N_4203);
nor U18995 (N_18995,N_7073,N_741);
or U18996 (N_18996,N_3432,N_4013);
nor U18997 (N_18997,N_635,N_595);
nor U18998 (N_18998,N_6550,N_4507);
or U18999 (N_18999,N_1272,N_3264);
nor U19000 (N_19000,N_1524,N_1073);
nor U19001 (N_19001,N_7992,N_9762);
or U19002 (N_19002,N_889,N_2118);
and U19003 (N_19003,N_4710,N_4551);
nor U19004 (N_19004,N_4089,N_9413);
xor U19005 (N_19005,N_1614,N_1134);
or U19006 (N_19006,N_6409,N_2050);
and U19007 (N_19007,N_2255,N_6595);
nand U19008 (N_19008,N_3825,N_2393);
nor U19009 (N_19009,N_4662,N_1975);
and U19010 (N_19010,N_6870,N_7901);
nor U19011 (N_19011,N_7269,N_2627);
or U19012 (N_19012,N_4422,N_4083);
nand U19013 (N_19013,N_4207,N_9851);
nor U19014 (N_19014,N_8222,N_404);
nand U19015 (N_19015,N_6401,N_4843);
nand U19016 (N_19016,N_6972,N_8415);
or U19017 (N_19017,N_1869,N_2436);
nand U19018 (N_19018,N_8726,N_6861);
nor U19019 (N_19019,N_950,N_6961);
nand U19020 (N_19020,N_2412,N_8743);
nor U19021 (N_19021,N_4928,N_2722);
nand U19022 (N_19022,N_4114,N_3361);
or U19023 (N_19023,N_4226,N_6835);
nor U19024 (N_19024,N_3470,N_800);
nand U19025 (N_19025,N_9136,N_7693);
nand U19026 (N_19026,N_5378,N_4238);
and U19027 (N_19027,N_258,N_609);
and U19028 (N_19028,N_9067,N_3500);
or U19029 (N_19029,N_6953,N_3618);
and U19030 (N_19030,N_3309,N_3190);
or U19031 (N_19031,N_9116,N_5181);
nand U19032 (N_19032,N_4402,N_1915);
and U19033 (N_19033,N_4518,N_653);
nor U19034 (N_19034,N_2714,N_8014);
nand U19035 (N_19035,N_8336,N_7279);
nor U19036 (N_19036,N_6318,N_4725);
or U19037 (N_19037,N_5062,N_5480);
nand U19038 (N_19038,N_2699,N_4863);
nor U19039 (N_19039,N_1921,N_2968);
and U19040 (N_19040,N_4437,N_8577);
or U19041 (N_19041,N_2528,N_226);
or U19042 (N_19042,N_1258,N_2903);
nand U19043 (N_19043,N_2830,N_4647);
and U19044 (N_19044,N_6845,N_5964);
nand U19045 (N_19045,N_9278,N_6944);
or U19046 (N_19046,N_4336,N_3859);
and U19047 (N_19047,N_1483,N_9696);
or U19048 (N_19048,N_5474,N_425);
nand U19049 (N_19049,N_7128,N_6897);
and U19050 (N_19050,N_1393,N_549);
nor U19051 (N_19051,N_9659,N_2536);
nor U19052 (N_19052,N_9479,N_4837);
nand U19053 (N_19053,N_4330,N_2851);
or U19054 (N_19054,N_5841,N_122);
or U19055 (N_19055,N_9859,N_5152);
and U19056 (N_19056,N_8672,N_8807);
and U19057 (N_19057,N_2630,N_19);
nand U19058 (N_19058,N_6927,N_3276);
nand U19059 (N_19059,N_3515,N_1976);
nand U19060 (N_19060,N_2726,N_8962);
or U19061 (N_19061,N_7754,N_1282);
nor U19062 (N_19062,N_371,N_5404);
and U19063 (N_19063,N_7812,N_2756);
nand U19064 (N_19064,N_6856,N_7177);
and U19065 (N_19065,N_4065,N_6201);
nor U19066 (N_19066,N_7837,N_6952);
and U19067 (N_19067,N_5322,N_9026);
nor U19068 (N_19068,N_3288,N_8867);
and U19069 (N_19069,N_5050,N_8855);
nor U19070 (N_19070,N_5202,N_8731);
nor U19071 (N_19071,N_4566,N_8281);
nor U19072 (N_19072,N_5091,N_6112);
nand U19073 (N_19073,N_2317,N_1454);
or U19074 (N_19074,N_3694,N_6113);
or U19075 (N_19075,N_2837,N_8128);
nor U19076 (N_19076,N_6537,N_2262);
or U19077 (N_19077,N_7773,N_6868);
and U19078 (N_19078,N_6657,N_115);
nor U19079 (N_19079,N_870,N_1936);
nor U19080 (N_19080,N_9018,N_2144);
nand U19081 (N_19081,N_915,N_8486);
and U19082 (N_19082,N_6070,N_5404);
or U19083 (N_19083,N_8045,N_4806);
or U19084 (N_19084,N_7074,N_8442);
and U19085 (N_19085,N_6639,N_7717);
or U19086 (N_19086,N_7362,N_6188);
and U19087 (N_19087,N_6518,N_3204);
nand U19088 (N_19088,N_8249,N_9449);
xor U19089 (N_19089,N_2523,N_607);
nand U19090 (N_19090,N_14,N_8789);
or U19091 (N_19091,N_9014,N_1840);
nor U19092 (N_19092,N_6293,N_140);
or U19093 (N_19093,N_3900,N_2330);
nor U19094 (N_19094,N_2797,N_6272);
and U19095 (N_19095,N_2314,N_689);
nand U19096 (N_19096,N_2619,N_8591);
nand U19097 (N_19097,N_4025,N_2953);
nand U19098 (N_19098,N_7502,N_4348);
and U19099 (N_19099,N_6950,N_4365);
and U19100 (N_19100,N_7101,N_5713);
nand U19101 (N_19101,N_9484,N_8055);
and U19102 (N_19102,N_6692,N_5655);
nand U19103 (N_19103,N_8638,N_2844);
nand U19104 (N_19104,N_9755,N_5662);
nand U19105 (N_19105,N_9304,N_1348);
nor U19106 (N_19106,N_1185,N_5629);
or U19107 (N_19107,N_3200,N_4276);
nor U19108 (N_19108,N_7527,N_1996);
nand U19109 (N_19109,N_4919,N_1080);
nor U19110 (N_19110,N_1910,N_5687);
or U19111 (N_19111,N_6798,N_8803);
nor U19112 (N_19112,N_8350,N_3798);
nor U19113 (N_19113,N_1100,N_862);
nand U19114 (N_19114,N_7685,N_7748);
or U19115 (N_19115,N_65,N_9931);
nand U19116 (N_19116,N_2420,N_5139);
nor U19117 (N_19117,N_9745,N_2313);
nor U19118 (N_19118,N_1891,N_7819);
nand U19119 (N_19119,N_7924,N_9739);
and U19120 (N_19120,N_293,N_5271);
or U19121 (N_19121,N_1987,N_8807);
and U19122 (N_19122,N_5164,N_1210);
nand U19123 (N_19123,N_2985,N_4594);
xor U19124 (N_19124,N_4155,N_2386);
nand U19125 (N_19125,N_6260,N_3996);
or U19126 (N_19126,N_4502,N_6680);
or U19127 (N_19127,N_1788,N_4117);
nor U19128 (N_19128,N_7846,N_3754);
and U19129 (N_19129,N_9732,N_5538);
or U19130 (N_19130,N_4206,N_1030);
or U19131 (N_19131,N_7746,N_2428);
and U19132 (N_19132,N_1072,N_1512);
and U19133 (N_19133,N_3333,N_2318);
nand U19134 (N_19134,N_6023,N_8743);
nand U19135 (N_19135,N_4592,N_7213);
nor U19136 (N_19136,N_7131,N_8251);
or U19137 (N_19137,N_6813,N_4977);
nand U19138 (N_19138,N_6140,N_8662);
nand U19139 (N_19139,N_7223,N_2954);
or U19140 (N_19140,N_6952,N_8664);
nand U19141 (N_19141,N_4793,N_9040);
nand U19142 (N_19142,N_8767,N_6658);
or U19143 (N_19143,N_1341,N_2523);
nand U19144 (N_19144,N_4486,N_6795);
nand U19145 (N_19145,N_9638,N_2484);
nor U19146 (N_19146,N_1257,N_2014);
nor U19147 (N_19147,N_3510,N_6261);
or U19148 (N_19148,N_5063,N_5270);
nor U19149 (N_19149,N_8418,N_6002);
or U19150 (N_19150,N_5322,N_3824);
and U19151 (N_19151,N_1727,N_2852);
and U19152 (N_19152,N_3955,N_1753);
nor U19153 (N_19153,N_7613,N_6142);
or U19154 (N_19154,N_9068,N_6460);
or U19155 (N_19155,N_6319,N_6101);
nor U19156 (N_19156,N_9061,N_469);
nand U19157 (N_19157,N_9910,N_2048);
or U19158 (N_19158,N_455,N_6493);
nor U19159 (N_19159,N_5658,N_3205);
and U19160 (N_19160,N_2020,N_5160);
and U19161 (N_19161,N_6940,N_7535);
nand U19162 (N_19162,N_1033,N_6971);
or U19163 (N_19163,N_3924,N_5473);
and U19164 (N_19164,N_9504,N_1254);
and U19165 (N_19165,N_9537,N_2823);
nand U19166 (N_19166,N_788,N_5680);
nand U19167 (N_19167,N_6624,N_5296);
and U19168 (N_19168,N_1542,N_2061);
or U19169 (N_19169,N_1716,N_2688);
or U19170 (N_19170,N_8642,N_619);
nor U19171 (N_19171,N_982,N_1335);
nand U19172 (N_19172,N_7698,N_9454);
nand U19173 (N_19173,N_410,N_7394);
nand U19174 (N_19174,N_2475,N_9512);
and U19175 (N_19175,N_8022,N_7800);
nor U19176 (N_19176,N_1177,N_3702);
nor U19177 (N_19177,N_3715,N_7045);
and U19178 (N_19178,N_1474,N_9041);
nor U19179 (N_19179,N_7851,N_4457);
or U19180 (N_19180,N_8791,N_3130);
or U19181 (N_19181,N_1605,N_7227);
nor U19182 (N_19182,N_3025,N_1790);
and U19183 (N_19183,N_7577,N_3206);
and U19184 (N_19184,N_660,N_1573);
or U19185 (N_19185,N_9934,N_7825);
nand U19186 (N_19186,N_4091,N_758);
or U19187 (N_19187,N_8843,N_2971);
nor U19188 (N_19188,N_4979,N_2291);
or U19189 (N_19189,N_8025,N_2981);
nand U19190 (N_19190,N_8899,N_2823);
and U19191 (N_19191,N_3349,N_4557);
nor U19192 (N_19192,N_7544,N_3774);
or U19193 (N_19193,N_671,N_3941);
nand U19194 (N_19194,N_4383,N_5610);
nand U19195 (N_19195,N_3185,N_1652);
nand U19196 (N_19196,N_3786,N_4883);
nand U19197 (N_19197,N_2292,N_4399);
and U19198 (N_19198,N_4592,N_7234);
or U19199 (N_19199,N_5856,N_7576);
and U19200 (N_19200,N_5195,N_3992);
xor U19201 (N_19201,N_3864,N_6975);
or U19202 (N_19202,N_9153,N_7744);
nor U19203 (N_19203,N_5693,N_446);
or U19204 (N_19204,N_6296,N_8080);
or U19205 (N_19205,N_9367,N_7722);
or U19206 (N_19206,N_769,N_5162);
or U19207 (N_19207,N_4681,N_5990);
nand U19208 (N_19208,N_8885,N_2005);
and U19209 (N_19209,N_3826,N_8266);
nand U19210 (N_19210,N_7826,N_8877);
nand U19211 (N_19211,N_2558,N_3045);
nor U19212 (N_19212,N_8094,N_1084);
and U19213 (N_19213,N_5668,N_3494);
nand U19214 (N_19214,N_8075,N_7728);
nor U19215 (N_19215,N_3559,N_7145);
xnor U19216 (N_19216,N_4013,N_8518);
or U19217 (N_19217,N_5055,N_6494);
nand U19218 (N_19218,N_2241,N_9123);
nand U19219 (N_19219,N_6714,N_2725);
and U19220 (N_19220,N_1111,N_8666);
nand U19221 (N_19221,N_8840,N_8463);
nand U19222 (N_19222,N_9275,N_7626);
nor U19223 (N_19223,N_7558,N_1995);
or U19224 (N_19224,N_1687,N_556);
or U19225 (N_19225,N_1502,N_6286);
or U19226 (N_19226,N_52,N_9646);
and U19227 (N_19227,N_9466,N_4762);
or U19228 (N_19228,N_4161,N_778);
nor U19229 (N_19229,N_7925,N_1931);
nor U19230 (N_19230,N_625,N_1936);
nor U19231 (N_19231,N_701,N_5243);
and U19232 (N_19232,N_2165,N_5071);
and U19233 (N_19233,N_9917,N_6578);
and U19234 (N_19234,N_3012,N_4305);
xnor U19235 (N_19235,N_5649,N_3385);
nand U19236 (N_19236,N_6558,N_1207);
nor U19237 (N_19237,N_316,N_2080);
or U19238 (N_19238,N_2279,N_7202);
nand U19239 (N_19239,N_2670,N_3405);
nand U19240 (N_19240,N_5831,N_3362);
and U19241 (N_19241,N_5359,N_1346);
nand U19242 (N_19242,N_6648,N_8283);
and U19243 (N_19243,N_9045,N_1250);
or U19244 (N_19244,N_3807,N_1065);
nor U19245 (N_19245,N_185,N_8383);
or U19246 (N_19246,N_639,N_5015);
nor U19247 (N_19247,N_3528,N_8790);
or U19248 (N_19248,N_9804,N_9571);
nor U19249 (N_19249,N_5019,N_1546);
nor U19250 (N_19250,N_2364,N_53);
and U19251 (N_19251,N_5265,N_5170);
and U19252 (N_19252,N_186,N_4443);
nand U19253 (N_19253,N_264,N_475);
nand U19254 (N_19254,N_7946,N_2987);
and U19255 (N_19255,N_5009,N_9800);
nand U19256 (N_19256,N_7748,N_6237);
or U19257 (N_19257,N_3861,N_347);
or U19258 (N_19258,N_3926,N_8747);
or U19259 (N_19259,N_9428,N_7422);
nand U19260 (N_19260,N_4772,N_4327);
or U19261 (N_19261,N_1049,N_2310);
or U19262 (N_19262,N_6489,N_3887);
and U19263 (N_19263,N_8889,N_6501);
or U19264 (N_19264,N_5180,N_9935);
or U19265 (N_19265,N_2998,N_6471);
nor U19266 (N_19266,N_9411,N_3394);
and U19267 (N_19267,N_4861,N_4162);
or U19268 (N_19268,N_8312,N_5862);
or U19269 (N_19269,N_8500,N_2561);
nor U19270 (N_19270,N_3054,N_4022);
nor U19271 (N_19271,N_5381,N_3376);
nor U19272 (N_19272,N_5562,N_9426);
and U19273 (N_19273,N_6787,N_5183);
and U19274 (N_19274,N_8231,N_4502);
nor U19275 (N_19275,N_3623,N_5849);
and U19276 (N_19276,N_9518,N_2131);
nor U19277 (N_19277,N_9826,N_7975);
or U19278 (N_19278,N_9064,N_7661);
nor U19279 (N_19279,N_4788,N_9817);
nor U19280 (N_19280,N_202,N_8908);
or U19281 (N_19281,N_2573,N_143);
nor U19282 (N_19282,N_1189,N_9343);
or U19283 (N_19283,N_9512,N_7805);
or U19284 (N_19284,N_503,N_388);
nor U19285 (N_19285,N_4430,N_6129);
nand U19286 (N_19286,N_1463,N_5246);
or U19287 (N_19287,N_6049,N_3883);
and U19288 (N_19288,N_466,N_368);
and U19289 (N_19289,N_2354,N_7198);
and U19290 (N_19290,N_9820,N_5013);
nand U19291 (N_19291,N_780,N_5696);
or U19292 (N_19292,N_7297,N_4233);
nand U19293 (N_19293,N_4381,N_8605);
and U19294 (N_19294,N_4154,N_3015);
or U19295 (N_19295,N_2204,N_1101);
nor U19296 (N_19296,N_9635,N_5605);
or U19297 (N_19297,N_3549,N_6108);
nand U19298 (N_19298,N_3653,N_6866);
xor U19299 (N_19299,N_9028,N_1593);
or U19300 (N_19300,N_6991,N_8410);
or U19301 (N_19301,N_5058,N_6490);
nand U19302 (N_19302,N_9609,N_5363);
or U19303 (N_19303,N_9623,N_8080);
or U19304 (N_19304,N_6268,N_7966);
nor U19305 (N_19305,N_1331,N_6268);
or U19306 (N_19306,N_5420,N_1657);
nand U19307 (N_19307,N_1233,N_3608);
and U19308 (N_19308,N_6403,N_3729);
nand U19309 (N_19309,N_3057,N_9172);
or U19310 (N_19310,N_2494,N_9815);
and U19311 (N_19311,N_1602,N_4091);
and U19312 (N_19312,N_9376,N_511);
nand U19313 (N_19313,N_6471,N_2337);
nand U19314 (N_19314,N_3867,N_2979);
nand U19315 (N_19315,N_2711,N_3723);
or U19316 (N_19316,N_7429,N_3203);
nand U19317 (N_19317,N_8111,N_271);
and U19318 (N_19318,N_5102,N_7193);
or U19319 (N_19319,N_1315,N_4543);
or U19320 (N_19320,N_639,N_5704);
nand U19321 (N_19321,N_8811,N_6601);
nor U19322 (N_19322,N_2838,N_7725);
and U19323 (N_19323,N_5194,N_5568);
nor U19324 (N_19324,N_2853,N_9718);
or U19325 (N_19325,N_3232,N_6251);
nand U19326 (N_19326,N_8935,N_923);
nor U19327 (N_19327,N_3463,N_9484);
nand U19328 (N_19328,N_1802,N_561);
or U19329 (N_19329,N_8120,N_1941);
and U19330 (N_19330,N_9538,N_1868);
and U19331 (N_19331,N_6803,N_7668);
nor U19332 (N_19332,N_4394,N_7773);
and U19333 (N_19333,N_2899,N_2532);
and U19334 (N_19334,N_3911,N_2506);
or U19335 (N_19335,N_5627,N_8080);
or U19336 (N_19336,N_4524,N_9715);
nor U19337 (N_19337,N_9731,N_6299);
nor U19338 (N_19338,N_7228,N_12);
nand U19339 (N_19339,N_9411,N_8989);
or U19340 (N_19340,N_5351,N_6229);
nand U19341 (N_19341,N_8845,N_2921);
or U19342 (N_19342,N_1989,N_8996);
nand U19343 (N_19343,N_9636,N_5387);
nor U19344 (N_19344,N_9886,N_4177);
nand U19345 (N_19345,N_9486,N_7691);
nor U19346 (N_19346,N_2724,N_4460);
nor U19347 (N_19347,N_3036,N_3525);
xor U19348 (N_19348,N_2708,N_3024);
nand U19349 (N_19349,N_2026,N_2910);
nor U19350 (N_19350,N_4768,N_676);
and U19351 (N_19351,N_7735,N_9452);
or U19352 (N_19352,N_175,N_9378);
nand U19353 (N_19353,N_6740,N_5726);
nor U19354 (N_19354,N_9632,N_2726);
nand U19355 (N_19355,N_2017,N_1302);
nand U19356 (N_19356,N_2434,N_5806);
or U19357 (N_19357,N_2099,N_5379);
and U19358 (N_19358,N_7057,N_9541);
or U19359 (N_19359,N_5598,N_3250);
nand U19360 (N_19360,N_1186,N_1109);
and U19361 (N_19361,N_8737,N_8924);
nor U19362 (N_19362,N_6083,N_6992);
nor U19363 (N_19363,N_3061,N_3456);
or U19364 (N_19364,N_8789,N_3221);
nor U19365 (N_19365,N_6235,N_2613);
nand U19366 (N_19366,N_2435,N_1622);
or U19367 (N_19367,N_9619,N_1469);
nand U19368 (N_19368,N_9526,N_7999);
or U19369 (N_19369,N_8115,N_8350);
nand U19370 (N_19370,N_5222,N_7199);
nand U19371 (N_19371,N_6461,N_458);
xnor U19372 (N_19372,N_1394,N_9286);
nand U19373 (N_19373,N_354,N_3068);
nand U19374 (N_19374,N_1254,N_93);
nand U19375 (N_19375,N_4709,N_5805);
and U19376 (N_19376,N_4452,N_1724);
nor U19377 (N_19377,N_2904,N_7743);
nor U19378 (N_19378,N_2059,N_7087);
and U19379 (N_19379,N_1246,N_8083);
nor U19380 (N_19380,N_1675,N_9858);
or U19381 (N_19381,N_5816,N_2101);
nor U19382 (N_19382,N_9618,N_4688);
nand U19383 (N_19383,N_7157,N_3897);
nor U19384 (N_19384,N_5643,N_5389);
nand U19385 (N_19385,N_4716,N_2965);
or U19386 (N_19386,N_9804,N_5602);
or U19387 (N_19387,N_7916,N_4154);
nand U19388 (N_19388,N_4548,N_936);
or U19389 (N_19389,N_4872,N_3823);
or U19390 (N_19390,N_242,N_8081);
or U19391 (N_19391,N_1422,N_6291);
nand U19392 (N_19392,N_184,N_5994);
and U19393 (N_19393,N_7953,N_757);
nor U19394 (N_19394,N_6887,N_2233);
or U19395 (N_19395,N_9617,N_8943);
or U19396 (N_19396,N_9159,N_175);
nor U19397 (N_19397,N_3817,N_4780);
nor U19398 (N_19398,N_9014,N_1838);
xnor U19399 (N_19399,N_9538,N_5160);
nor U19400 (N_19400,N_8025,N_7421);
nor U19401 (N_19401,N_5030,N_1936);
nor U19402 (N_19402,N_5660,N_2096);
and U19403 (N_19403,N_6791,N_2299);
nor U19404 (N_19404,N_3157,N_7764);
and U19405 (N_19405,N_8733,N_358);
nand U19406 (N_19406,N_8047,N_6119);
nor U19407 (N_19407,N_1207,N_8271);
nor U19408 (N_19408,N_5704,N_7077);
nor U19409 (N_19409,N_8169,N_5093);
and U19410 (N_19410,N_4574,N_6253);
or U19411 (N_19411,N_2164,N_4033);
nand U19412 (N_19412,N_3343,N_2895);
and U19413 (N_19413,N_8112,N_244);
nand U19414 (N_19414,N_6476,N_4181);
nor U19415 (N_19415,N_1877,N_8942);
or U19416 (N_19416,N_9268,N_1230);
or U19417 (N_19417,N_6976,N_5406);
xor U19418 (N_19418,N_3248,N_881);
nor U19419 (N_19419,N_6697,N_6493);
nand U19420 (N_19420,N_2500,N_3906);
and U19421 (N_19421,N_4269,N_8412);
and U19422 (N_19422,N_3553,N_6741);
or U19423 (N_19423,N_8277,N_5423);
or U19424 (N_19424,N_8636,N_2267);
nor U19425 (N_19425,N_2760,N_6112);
or U19426 (N_19426,N_4536,N_4502);
or U19427 (N_19427,N_7817,N_1012);
nand U19428 (N_19428,N_1488,N_6802);
nand U19429 (N_19429,N_4440,N_9869);
or U19430 (N_19430,N_1120,N_6457);
nor U19431 (N_19431,N_3089,N_8816);
xnor U19432 (N_19432,N_4073,N_6936);
nand U19433 (N_19433,N_6467,N_3595);
nor U19434 (N_19434,N_2793,N_5116);
and U19435 (N_19435,N_1017,N_8902);
xnor U19436 (N_19436,N_1616,N_2434);
or U19437 (N_19437,N_9526,N_1835);
nor U19438 (N_19438,N_5994,N_9876);
nand U19439 (N_19439,N_9145,N_9225);
or U19440 (N_19440,N_6594,N_2114);
nand U19441 (N_19441,N_1134,N_7154);
nand U19442 (N_19442,N_9018,N_4845);
nor U19443 (N_19443,N_6717,N_8441);
xor U19444 (N_19444,N_5159,N_1240);
and U19445 (N_19445,N_6920,N_6245);
or U19446 (N_19446,N_3114,N_3401);
or U19447 (N_19447,N_3199,N_1675);
nor U19448 (N_19448,N_9499,N_6557);
and U19449 (N_19449,N_3207,N_4967);
nand U19450 (N_19450,N_6620,N_6972);
nor U19451 (N_19451,N_5308,N_3622);
or U19452 (N_19452,N_2567,N_9430);
nand U19453 (N_19453,N_8338,N_7924);
nor U19454 (N_19454,N_2010,N_6623);
nor U19455 (N_19455,N_9303,N_7388);
or U19456 (N_19456,N_4903,N_8936);
and U19457 (N_19457,N_7480,N_2058);
nand U19458 (N_19458,N_273,N_7217);
xor U19459 (N_19459,N_8313,N_2998);
nor U19460 (N_19460,N_2228,N_2429);
nand U19461 (N_19461,N_9884,N_1405);
nand U19462 (N_19462,N_3976,N_8474);
nand U19463 (N_19463,N_2648,N_3279);
nand U19464 (N_19464,N_1467,N_637);
nor U19465 (N_19465,N_1449,N_2617);
or U19466 (N_19466,N_9445,N_5849);
xor U19467 (N_19467,N_4142,N_8666);
nor U19468 (N_19468,N_7534,N_8107);
or U19469 (N_19469,N_4065,N_1929);
and U19470 (N_19470,N_2039,N_2272);
and U19471 (N_19471,N_1015,N_444);
nand U19472 (N_19472,N_651,N_1428);
and U19473 (N_19473,N_4672,N_817);
and U19474 (N_19474,N_9177,N_7420);
or U19475 (N_19475,N_6296,N_1773);
nor U19476 (N_19476,N_9134,N_8384);
and U19477 (N_19477,N_8088,N_8664);
nor U19478 (N_19478,N_8240,N_7701);
and U19479 (N_19479,N_880,N_136);
nand U19480 (N_19480,N_7163,N_4306);
and U19481 (N_19481,N_800,N_9442);
nor U19482 (N_19482,N_9801,N_8047);
xnor U19483 (N_19483,N_7082,N_5686);
and U19484 (N_19484,N_6015,N_3223);
nor U19485 (N_19485,N_6667,N_3190);
and U19486 (N_19486,N_281,N_5970);
or U19487 (N_19487,N_6472,N_4888);
and U19488 (N_19488,N_6265,N_8112);
nor U19489 (N_19489,N_9008,N_7405);
nor U19490 (N_19490,N_4369,N_8804);
nor U19491 (N_19491,N_4247,N_8011);
nand U19492 (N_19492,N_1129,N_1200);
nand U19493 (N_19493,N_2445,N_228);
nor U19494 (N_19494,N_6168,N_355);
and U19495 (N_19495,N_4502,N_3478);
and U19496 (N_19496,N_1815,N_5294);
or U19497 (N_19497,N_8532,N_3036);
or U19498 (N_19498,N_3951,N_3536);
and U19499 (N_19499,N_562,N_1952);
or U19500 (N_19500,N_3237,N_1443);
and U19501 (N_19501,N_4760,N_9251);
nor U19502 (N_19502,N_2015,N_45);
or U19503 (N_19503,N_507,N_7266);
nor U19504 (N_19504,N_7836,N_2026);
nor U19505 (N_19505,N_47,N_3335);
nor U19506 (N_19506,N_3134,N_4315);
and U19507 (N_19507,N_1119,N_5575);
and U19508 (N_19508,N_8253,N_3676);
nand U19509 (N_19509,N_2121,N_6157);
and U19510 (N_19510,N_5718,N_7788);
nand U19511 (N_19511,N_2184,N_4034);
and U19512 (N_19512,N_5181,N_9620);
nand U19513 (N_19513,N_8307,N_9554);
or U19514 (N_19514,N_3864,N_7474);
or U19515 (N_19515,N_8300,N_5204);
nand U19516 (N_19516,N_2061,N_1035);
and U19517 (N_19517,N_2997,N_7733);
nand U19518 (N_19518,N_6152,N_3058);
nand U19519 (N_19519,N_7218,N_7826);
nand U19520 (N_19520,N_2155,N_8441);
or U19521 (N_19521,N_8381,N_5153);
nand U19522 (N_19522,N_7257,N_5466);
nor U19523 (N_19523,N_6905,N_8285);
or U19524 (N_19524,N_3836,N_8849);
nand U19525 (N_19525,N_3169,N_4472);
or U19526 (N_19526,N_498,N_8072);
nand U19527 (N_19527,N_9795,N_9708);
nor U19528 (N_19528,N_4443,N_6693);
nand U19529 (N_19529,N_2765,N_6654);
nand U19530 (N_19530,N_248,N_4841);
or U19531 (N_19531,N_9883,N_9797);
or U19532 (N_19532,N_3196,N_3033);
or U19533 (N_19533,N_6496,N_2232);
nand U19534 (N_19534,N_6976,N_9205);
nand U19535 (N_19535,N_1373,N_8793);
or U19536 (N_19536,N_3999,N_6744);
nor U19537 (N_19537,N_5896,N_3495);
or U19538 (N_19538,N_9896,N_5697);
nand U19539 (N_19539,N_2340,N_3629);
and U19540 (N_19540,N_5846,N_7171);
nand U19541 (N_19541,N_6590,N_5607);
nand U19542 (N_19542,N_7894,N_7380);
nand U19543 (N_19543,N_7432,N_7732);
nor U19544 (N_19544,N_6518,N_7349);
or U19545 (N_19545,N_8229,N_9437);
nor U19546 (N_19546,N_5129,N_1011);
nor U19547 (N_19547,N_3013,N_5572);
and U19548 (N_19548,N_3764,N_3506);
and U19549 (N_19549,N_2480,N_1455);
or U19550 (N_19550,N_1532,N_4416);
or U19551 (N_19551,N_6042,N_6058);
nor U19552 (N_19552,N_1639,N_1065);
or U19553 (N_19553,N_236,N_5708);
nor U19554 (N_19554,N_7740,N_3011);
nor U19555 (N_19555,N_4953,N_2347);
nor U19556 (N_19556,N_691,N_2497);
nor U19557 (N_19557,N_3504,N_9437);
nor U19558 (N_19558,N_1262,N_8854);
nand U19559 (N_19559,N_6921,N_2684);
nand U19560 (N_19560,N_4314,N_5192);
nand U19561 (N_19561,N_970,N_6593);
or U19562 (N_19562,N_1453,N_7810);
nand U19563 (N_19563,N_376,N_5571);
nand U19564 (N_19564,N_3149,N_9404);
nand U19565 (N_19565,N_19,N_9254);
nand U19566 (N_19566,N_5127,N_6177);
nand U19567 (N_19567,N_6501,N_3295);
nand U19568 (N_19568,N_7593,N_5798);
and U19569 (N_19569,N_3037,N_7734);
or U19570 (N_19570,N_9110,N_1196);
or U19571 (N_19571,N_6271,N_7288);
nand U19572 (N_19572,N_3780,N_2688);
nand U19573 (N_19573,N_5807,N_6880);
nand U19574 (N_19574,N_5023,N_6174);
nor U19575 (N_19575,N_6083,N_308);
or U19576 (N_19576,N_3293,N_2216);
nand U19577 (N_19577,N_6978,N_8871);
nor U19578 (N_19578,N_9158,N_1456);
or U19579 (N_19579,N_1139,N_8636);
nor U19580 (N_19580,N_238,N_2181);
nor U19581 (N_19581,N_7889,N_9590);
nand U19582 (N_19582,N_6915,N_9870);
and U19583 (N_19583,N_7599,N_1041);
nand U19584 (N_19584,N_4045,N_8157);
nand U19585 (N_19585,N_4352,N_651);
and U19586 (N_19586,N_3079,N_5997);
xor U19587 (N_19587,N_4380,N_5165);
nand U19588 (N_19588,N_6870,N_4071);
and U19589 (N_19589,N_5867,N_3096);
and U19590 (N_19590,N_5954,N_6981);
nor U19591 (N_19591,N_1537,N_2999);
nor U19592 (N_19592,N_3576,N_279);
nor U19593 (N_19593,N_6350,N_9934);
or U19594 (N_19594,N_6005,N_7392);
or U19595 (N_19595,N_8206,N_3767);
nor U19596 (N_19596,N_1098,N_6359);
nand U19597 (N_19597,N_3998,N_6522);
or U19598 (N_19598,N_8429,N_4096);
nand U19599 (N_19599,N_2436,N_4461);
nand U19600 (N_19600,N_6091,N_6509);
nand U19601 (N_19601,N_4537,N_2757);
or U19602 (N_19602,N_6807,N_9078);
or U19603 (N_19603,N_446,N_5761);
or U19604 (N_19604,N_5678,N_8454);
or U19605 (N_19605,N_1786,N_1362);
nand U19606 (N_19606,N_3593,N_3066);
or U19607 (N_19607,N_514,N_3015);
or U19608 (N_19608,N_9783,N_2525);
nor U19609 (N_19609,N_2586,N_5541);
nor U19610 (N_19610,N_5485,N_7752);
nor U19611 (N_19611,N_8899,N_808);
nand U19612 (N_19612,N_480,N_2763);
or U19613 (N_19613,N_4950,N_4839);
and U19614 (N_19614,N_3632,N_8110);
nor U19615 (N_19615,N_675,N_7617);
nand U19616 (N_19616,N_748,N_7658);
or U19617 (N_19617,N_6815,N_1722);
and U19618 (N_19618,N_4510,N_5373);
or U19619 (N_19619,N_6354,N_8105);
and U19620 (N_19620,N_4236,N_4283);
and U19621 (N_19621,N_692,N_7311);
or U19622 (N_19622,N_9496,N_4943);
xnor U19623 (N_19623,N_8696,N_431);
xnor U19624 (N_19624,N_8320,N_4326);
or U19625 (N_19625,N_3856,N_9436);
nor U19626 (N_19626,N_3224,N_6558);
nand U19627 (N_19627,N_1647,N_6350);
and U19628 (N_19628,N_2726,N_3662);
nor U19629 (N_19629,N_7277,N_9434);
nand U19630 (N_19630,N_3272,N_2467);
nand U19631 (N_19631,N_5040,N_5604);
nor U19632 (N_19632,N_9026,N_4648);
or U19633 (N_19633,N_4765,N_4262);
nor U19634 (N_19634,N_966,N_6452);
or U19635 (N_19635,N_2869,N_5544);
nand U19636 (N_19636,N_4597,N_8243);
and U19637 (N_19637,N_8219,N_1411);
or U19638 (N_19638,N_2250,N_859);
nor U19639 (N_19639,N_6333,N_3852);
or U19640 (N_19640,N_6138,N_4292);
nor U19641 (N_19641,N_6554,N_7676);
nand U19642 (N_19642,N_8672,N_5607);
or U19643 (N_19643,N_4743,N_2149);
nand U19644 (N_19644,N_6203,N_310);
or U19645 (N_19645,N_2778,N_9207);
and U19646 (N_19646,N_6264,N_3221);
or U19647 (N_19647,N_8725,N_2017);
and U19648 (N_19648,N_9085,N_4661);
nor U19649 (N_19649,N_635,N_9855);
and U19650 (N_19650,N_3096,N_5359);
nor U19651 (N_19651,N_9351,N_9247);
nand U19652 (N_19652,N_943,N_8543);
nor U19653 (N_19653,N_3856,N_539);
nand U19654 (N_19654,N_8365,N_1143);
nand U19655 (N_19655,N_1172,N_493);
or U19656 (N_19656,N_595,N_4846);
or U19657 (N_19657,N_6816,N_8309);
nor U19658 (N_19658,N_6880,N_8325);
nor U19659 (N_19659,N_5421,N_8427);
nor U19660 (N_19660,N_5140,N_5137);
nand U19661 (N_19661,N_5415,N_6539);
or U19662 (N_19662,N_4383,N_2433);
or U19663 (N_19663,N_3225,N_5480);
and U19664 (N_19664,N_8053,N_9627);
nor U19665 (N_19665,N_8300,N_2198);
and U19666 (N_19666,N_5200,N_2192);
and U19667 (N_19667,N_6241,N_1603);
nand U19668 (N_19668,N_9384,N_2749);
nor U19669 (N_19669,N_8917,N_7607);
or U19670 (N_19670,N_5800,N_9119);
and U19671 (N_19671,N_9647,N_7040);
nand U19672 (N_19672,N_4547,N_8414);
or U19673 (N_19673,N_4440,N_2826);
nor U19674 (N_19674,N_2689,N_3927);
nor U19675 (N_19675,N_1955,N_4236);
or U19676 (N_19676,N_1972,N_571);
and U19677 (N_19677,N_4570,N_6476);
and U19678 (N_19678,N_4136,N_8275);
xnor U19679 (N_19679,N_7332,N_1670);
and U19680 (N_19680,N_4736,N_9046);
nor U19681 (N_19681,N_4336,N_976);
nor U19682 (N_19682,N_3458,N_9887);
nand U19683 (N_19683,N_212,N_2202);
and U19684 (N_19684,N_9415,N_9080);
nor U19685 (N_19685,N_9359,N_8139);
and U19686 (N_19686,N_6798,N_8143);
nand U19687 (N_19687,N_8838,N_4482);
nand U19688 (N_19688,N_9137,N_339);
nand U19689 (N_19689,N_9363,N_2335);
nand U19690 (N_19690,N_4046,N_9015);
nand U19691 (N_19691,N_7123,N_5602);
and U19692 (N_19692,N_6632,N_8042);
nand U19693 (N_19693,N_1897,N_4299);
and U19694 (N_19694,N_6698,N_3097);
and U19695 (N_19695,N_6947,N_569);
nand U19696 (N_19696,N_6823,N_4603);
or U19697 (N_19697,N_3713,N_5286);
or U19698 (N_19698,N_2189,N_1075);
and U19699 (N_19699,N_1966,N_5470);
nor U19700 (N_19700,N_7519,N_5513);
nor U19701 (N_19701,N_9197,N_8639);
and U19702 (N_19702,N_7124,N_683);
and U19703 (N_19703,N_3916,N_875);
or U19704 (N_19704,N_2712,N_5223);
and U19705 (N_19705,N_2558,N_2124);
nand U19706 (N_19706,N_7242,N_7279);
and U19707 (N_19707,N_7882,N_359);
nand U19708 (N_19708,N_8098,N_7919);
and U19709 (N_19709,N_4848,N_7904);
and U19710 (N_19710,N_9584,N_4891);
and U19711 (N_19711,N_3683,N_5851);
and U19712 (N_19712,N_9596,N_8187);
or U19713 (N_19713,N_9920,N_7934);
nor U19714 (N_19714,N_6802,N_4166);
or U19715 (N_19715,N_6677,N_8609);
nor U19716 (N_19716,N_1065,N_2292);
and U19717 (N_19717,N_2339,N_8008);
or U19718 (N_19718,N_9490,N_6474);
xnor U19719 (N_19719,N_6379,N_8085);
nand U19720 (N_19720,N_8602,N_991);
nand U19721 (N_19721,N_2386,N_6769);
nand U19722 (N_19722,N_229,N_3012);
or U19723 (N_19723,N_2384,N_34);
nor U19724 (N_19724,N_5744,N_868);
and U19725 (N_19725,N_6952,N_9386);
nor U19726 (N_19726,N_8104,N_2175);
nor U19727 (N_19727,N_6097,N_6992);
or U19728 (N_19728,N_5038,N_7771);
and U19729 (N_19729,N_6525,N_389);
and U19730 (N_19730,N_751,N_7541);
or U19731 (N_19731,N_503,N_33);
and U19732 (N_19732,N_700,N_1206);
or U19733 (N_19733,N_7673,N_7652);
nor U19734 (N_19734,N_5442,N_9903);
nor U19735 (N_19735,N_9859,N_6714);
nor U19736 (N_19736,N_2682,N_8760);
nor U19737 (N_19737,N_3481,N_6146);
nand U19738 (N_19738,N_2860,N_7477);
or U19739 (N_19739,N_7360,N_8978);
and U19740 (N_19740,N_9031,N_3485);
nor U19741 (N_19741,N_9373,N_1266);
nand U19742 (N_19742,N_2952,N_9248);
xor U19743 (N_19743,N_8139,N_6763);
nor U19744 (N_19744,N_8066,N_8629);
nand U19745 (N_19745,N_5870,N_6856);
or U19746 (N_19746,N_5881,N_4685);
and U19747 (N_19747,N_3083,N_8425);
nor U19748 (N_19748,N_7025,N_4042);
or U19749 (N_19749,N_6702,N_7542);
or U19750 (N_19750,N_6670,N_4845);
nand U19751 (N_19751,N_3472,N_3058);
nor U19752 (N_19752,N_2504,N_4783);
and U19753 (N_19753,N_4891,N_560);
nand U19754 (N_19754,N_850,N_8989);
nor U19755 (N_19755,N_7933,N_3934);
and U19756 (N_19756,N_651,N_9011);
nor U19757 (N_19757,N_5888,N_2666);
and U19758 (N_19758,N_9893,N_2716);
or U19759 (N_19759,N_838,N_1300);
nand U19760 (N_19760,N_3898,N_774);
nand U19761 (N_19761,N_130,N_1888);
nand U19762 (N_19762,N_9430,N_670);
nor U19763 (N_19763,N_2575,N_5500);
nor U19764 (N_19764,N_8958,N_4067);
and U19765 (N_19765,N_4227,N_1590);
or U19766 (N_19766,N_6018,N_3103);
and U19767 (N_19767,N_4129,N_1154);
or U19768 (N_19768,N_9314,N_4635);
or U19769 (N_19769,N_4334,N_6555);
nor U19770 (N_19770,N_5823,N_3515);
nand U19771 (N_19771,N_2304,N_1536);
and U19772 (N_19772,N_8162,N_8297);
nor U19773 (N_19773,N_1883,N_2115);
or U19774 (N_19774,N_4841,N_3692);
nand U19775 (N_19775,N_1309,N_1252);
nor U19776 (N_19776,N_9382,N_8509);
or U19777 (N_19777,N_5634,N_9223);
and U19778 (N_19778,N_973,N_5190);
or U19779 (N_19779,N_6448,N_1778);
or U19780 (N_19780,N_8498,N_7173);
nor U19781 (N_19781,N_5589,N_8344);
and U19782 (N_19782,N_781,N_3961);
and U19783 (N_19783,N_2952,N_5169);
nor U19784 (N_19784,N_2143,N_5299);
and U19785 (N_19785,N_4836,N_9893);
nor U19786 (N_19786,N_9816,N_8693);
nor U19787 (N_19787,N_5527,N_5654);
nor U19788 (N_19788,N_3232,N_7092);
or U19789 (N_19789,N_14,N_1937);
nand U19790 (N_19790,N_3430,N_2604);
nor U19791 (N_19791,N_9842,N_8288);
or U19792 (N_19792,N_8046,N_560);
nand U19793 (N_19793,N_9135,N_8031);
nand U19794 (N_19794,N_1951,N_5522);
or U19795 (N_19795,N_7904,N_8092);
nand U19796 (N_19796,N_3868,N_6303);
nor U19797 (N_19797,N_529,N_1116);
or U19798 (N_19798,N_3573,N_621);
nor U19799 (N_19799,N_3060,N_3859);
or U19800 (N_19800,N_2345,N_6434);
nor U19801 (N_19801,N_8192,N_9807);
nand U19802 (N_19802,N_2940,N_8019);
nor U19803 (N_19803,N_6494,N_6149);
nor U19804 (N_19804,N_6712,N_8808);
or U19805 (N_19805,N_4345,N_7709);
and U19806 (N_19806,N_7738,N_4610);
or U19807 (N_19807,N_3292,N_9185);
and U19808 (N_19808,N_6715,N_1676);
or U19809 (N_19809,N_278,N_155);
or U19810 (N_19810,N_407,N_9509);
and U19811 (N_19811,N_4725,N_9333);
nand U19812 (N_19812,N_9155,N_5358);
or U19813 (N_19813,N_8425,N_7352);
or U19814 (N_19814,N_8730,N_6451);
and U19815 (N_19815,N_8070,N_951);
nor U19816 (N_19816,N_7232,N_186);
nor U19817 (N_19817,N_6723,N_3782);
or U19818 (N_19818,N_388,N_8146);
nand U19819 (N_19819,N_9701,N_7355);
nor U19820 (N_19820,N_4658,N_2140);
and U19821 (N_19821,N_9459,N_6330);
nand U19822 (N_19822,N_6164,N_1758);
or U19823 (N_19823,N_9504,N_7567);
nand U19824 (N_19824,N_3742,N_7892);
xnor U19825 (N_19825,N_6035,N_7242);
nor U19826 (N_19826,N_2585,N_1248);
nand U19827 (N_19827,N_5354,N_8137);
and U19828 (N_19828,N_3196,N_4536);
nand U19829 (N_19829,N_9790,N_2684);
nand U19830 (N_19830,N_7226,N_878);
and U19831 (N_19831,N_2940,N_5330);
and U19832 (N_19832,N_8268,N_8264);
or U19833 (N_19833,N_4900,N_6138);
or U19834 (N_19834,N_1188,N_5291);
and U19835 (N_19835,N_1047,N_6791);
or U19836 (N_19836,N_8847,N_6035);
nor U19837 (N_19837,N_7759,N_4519);
nor U19838 (N_19838,N_795,N_486);
nand U19839 (N_19839,N_4161,N_3325);
nor U19840 (N_19840,N_1127,N_2544);
or U19841 (N_19841,N_7747,N_9604);
or U19842 (N_19842,N_5089,N_189);
nor U19843 (N_19843,N_9598,N_9670);
or U19844 (N_19844,N_6850,N_4711);
xor U19845 (N_19845,N_3789,N_3430);
and U19846 (N_19846,N_278,N_9716);
and U19847 (N_19847,N_2694,N_1676);
nor U19848 (N_19848,N_6323,N_480);
or U19849 (N_19849,N_7812,N_6932);
nor U19850 (N_19850,N_3154,N_2980);
and U19851 (N_19851,N_8847,N_7798);
and U19852 (N_19852,N_1199,N_7731);
and U19853 (N_19853,N_7902,N_9061);
or U19854 (N_19854,N_62,N_9244);
nor U19855 (N_19855,N_1407,N_4082);
nand U19856 (N_19856,N_1422,N_8746);
nand U19857 (N_19857,N_3927,N_1030);
or U19858 (N_19858,N_2650,N_5659);
and U19859 (N_19859,N_9456,N_7969);
or U19860 (N_19860,N_8589,N_8321);
and U19861 (N_19861,N_8076,N_9875);
and U19862 (N_19862,N_1062,N_2534);
nand U19863 (N_19863,N_3801,N_6223);
nor U19864 (N_19864,N_5576,N_3728);
nand U19865 (N_19865,N_3736,N_2573);
or U19866 (N_19866,N_1426,N_2828);
or U19867 (N_19867,N_4118,N_4930);
and U19868 (N_19868,N_1471,N_2775);
nand U19869 (N_19869,N_2012,N_899);
or U19870 (N_19870,N_8709,N_7146);
xnor U19871 (N_19871,N_6349,N_5584);
or U19872 (N_19872,N_7681,N_799);
nor U19873 (N_19873,N_145,N_3925);
nand U19874 (N_19874,N_741,N_8687);
nor U19875 (N_19875,N_2461,N_1462);
nand U19876 (N_19876,N_6410,N_8677);
and U19877 (N_19877,N_1845,N_8561);
nand U19878 (N_19878,N_4249,N_9352);
nor U19879 (N_19879,N_5491,N_8027);
and U19880 (N_19880,N_3006,N_3361);
and U19881 (N_19881,N_7094,N_9230);
and U19882 (N_19882,N_8252,N_3881);
and U19883 (N_19883,N_8815,N_8573);
nor U19884 (N_19884,N_2433,N_1308);
or U19885 (N_19885,N_3229,N_2921);
nand U19886 (N_19886,N_9950,N_7532);
nand U19887 (N_19887,N_8225,N_3529);
nor U19888 (N_19888,N_5393,N_6932);
and U19889 (N_19889,N_9874,N_2240);
nor U19890 (N_19890,N_8,N_8452);
nor U19891 (N_19891,N_4164,N_1745);
or U19892 (N_19892,N_7101,N_3426);
and U19893 (N_19893,N_3340,N_1403);
or U19894 (N_19894,N_6948,N_3459);
nor U19895 (N_19895,N_9273,N_6733);
and U19896 (N_19896,N_6629,N_9991);
and U19897 (N_19897,N_1516,N_9592);
or U19898 (N_19898,N_8785,N_4280);
or U19899 (N_19899,N_6512,N_6270);
and U19900 (N_19900,N_3971,N_5494);
nand U19901 (N_19901,N_5239,N_3233);
nor U19902 (N_19902,N_1147,N_9806);
or U19903 (N_19903,N_7644,N_5529);
nor U19904 (N_19904,N_2564,N_7295);
nand U19905 (N_19905,N_8802,N_2928);
nor U19906 (N_19906,N_4806,N_5069);
nor U19907 (N_19907,N_5823,N_8396);
nor U19908 (N_19908,N_3047,N_873);
or U19909 (N_19909,N_7129,N_163);
nor U19910 (N_19910,N_995,N_8761);
nand U19911 (N_19911,N_4611,N_9400);
and U19912 (N_19912,N_1320,N_6497);
nor U19913 (N_19913,N_3684,N_1558);
nand U19914 (N_19914,N_4615,N_1399);
nor U19915 (N_19915,N_1916,N_938);
nand U19916 (N_19916,N_2373,N_3690);
nand U19917 (N_19917,N_7928,N_7623);
nor U19918 (N_19918,N_8699,N_9494);
and U19919 (N_19919,N_7508,N_4640);
and U19920 (N_19920,N_104,N_861);
nand U19921 (N_19921,N_2790,N_4331);
nor U19922 (N_19922,N_602,N_7222);
nor U19923 (N_19923,N_7427,N_9966);
nand U19924 (N_19924,N_9397,N_1434);
and U19925 (N_19925,N_3055,N_8642);
nand U19926 (N_19926,N_4474,N_4207);
nand U19927 (N_19927,N_3971,N_3855);
nor U19928 (N_19928,N_3869,N_2575);
and U19929 (N_19929,N_3483,N_4858);
nand U19930 (N_19930,N_5955,N_8943);
nand U19931 (N_19931,N_9922,N_6989);
nor U19932 (N_19932,N_280,N_535);
and U19933 (N_19933,N_4921,N_736);
and U19934 (N_19934,N_1478,N_5117);
nor U19935 (N_19935,N_4988,N_4367);
nor U19936 (N_19936,N_4129,N_8479);
and U19937 (N_19937,N_4773,N_9958);
and U19938 (N_19938,N_2392,N_3257);
nor U19939 (N_19939,N_5689,N_496);
xnor U19940 (N_19940,N_9330,N_790);
or U19941 (N_19941,N_3015,N_9646);
nor U19942 (N_19942,N_1182,N_92);
nor U19943 (N_19943,N_8463,N_5538);
nor U19944 (N_19944,N_8426,N_9788);
or U19945 (N_19945,N_544,N_8474);
nor U19946 (N_19946,N_5810,N_4944);
nand U19947 (N_19947,N_9875,N_7101);
and U19948 (N_19948,N_9102,N_7523);
nor U19949 (N_19949,N_4687,N_5975);
or U19950 (N_19950,N_2542,N_4436);
nand U19951 (N_19951,N_8728,N_9258);
or U19952 (N_19952,N_7853,N_7400);
nor U19953 (N_19953,N_2024,N_2498);
and U19954 (N_19954,N_2958,N_2712);
and U19955 (N_19955,N_812,N_7153);
nor U19956 (N_19956,N_9294,N_8338);
and U19957 (N_19957,N_5825,N_3636);
nor U19958 (N_19958,N_7318,N_3100);
nand U19959 (N_19959,N_9547,N_3024);
and U19960 (N_19960,N_3900,N_3004);
or U19961 (N_19961,N_2506,N_2907);
and U19962 (N_19962,N_1970,N_6291);
and U19963 (N_19963,N_595,N_1673);
or U19964 (N_19964,N_2192,N_1889);
and U19965 (N_19965,N_6791,N_9339);
nand U19966 (N_19966,N_7826,N_9831);
nor U19967 (N_19967,N_311,N_5267);
nor U19968 (N_19968,N_7316,N_9694);
and U19969 (N_19969,N_2993,N_4500);
or U19970 (N_19970,N_2680,N_3499);
and U19971 (N_19971,N_5214,N_7432);
nand U19972 (N_19972,N_2893,N_6861);
and U19973 (N_19973,N_1953,N_2851);
or U19974 (N_19974,N_7823,N_477);
nand U19975 (N_19975,N_3652,N_34);
nand U19976 (N_19976,N_7753,N_6552);
nor U19977 (N_19977,N_1773,N_8934);
and U19978 (N_19978,N_2932,N_6230);
nand U19979 (N_19979,N_221,N_6932);
or U19980 (N_19980,N_3904,N_4871);
nand U19981 (N_19981,N_5482,N_1225);
nand U19982 (N_19982,N_1792,N_4299);
nor U19983 (N_19983,N_6385,N_6181);
or U19984 (N_19984,N_57,N_6642);
or U19985 (N_19985,N_4100,N_6653);
nand U19986 (N_19986,N_4121,N_7793);
nand U19987 (N_19987,N_5683,N_2027);
nand U19988 (N_19988,N_3453,N_9429);
and U19989 (N_19989,N_4641,N_8447);
nand U19990 (N_19990,N_61,N_5007);
and U19991 (N_19991,N_5661,N_5767);
or U19992 (N_19992,N_9837,N_3943);
or U19993 (N_19993,N_7339,N_9846);
and U19994 (N_19994,N_3905,N_1636);
nor U19995 (N_19995,N_7803,N_3452);
nand U19996 (N_19996,N_9678,N_3469);
nand U19997 (N_19997,N_9935,N_3296);
and U19998 (N_19998,N_480,N_8198);
nor U19999 (N_19999,N_221,N_7146);
nand U20000 (N_20000,N_12137,N_13595);
or U20001 (N_20001,N_14694,N_15144);
or U20002 (N_20002,N_15224,N_16130);
nor U20003 (N_20003,N_15041,N_17246);
and U20004 (N_20004,N_18936,N_15243);
nor U20005 (N_20005,N_11744,N_19756);
nor U20006 (N_20006,N_18039,N_18652);
nand U20007 (N_20007,N_13467,N_10726);
nand U20008 (N_20008,N_13038,N_12613);
or U20009 (N_20009,N_14248,N_13210);
nor U20010 (N_20010,N_16291,N_12851);
or U20011 (N_20011,N_15109,N_11139);
or U20012 (N_20012,N_12487,N_16231);
or U20013 (N_20013,N_12964,N_18741);
nand U20014 (N_20014,N_11125,N_19595);
nand U20015 (N_20015,N_15546,N_19402);
and U20016 (N_20016,N_17967,N_14152);
or U20017 (N_20017,N_18236,N_16634);
or U20018 (N_20018,N_18851,N_16373);
and U20019 (N_20019,N_16612,N_14031);
and U20020 (N_20020,N_11629,N_17468);
and U20021 (N_20021,N_16013,N_18161);
nand U20022 (N_20022,N_11817,N_13458);
or U20023 (N_20023,N_14830,N_17323);
or U20024 (N_20024,N_16700,N_14590);
nand U20025 (N_20025,N_10320,N_12539);
nor U20026 (N_20026,N_18891,N_10224);
nor U20027 (N_20027,N_19236,N_11997);
nor U20028 (N_20028,N_10333,N_17187);
and U20029 (N_20029,N_18769,N_19390);
nor U20030 (N_20030,N_19108,N_19344);
nand U20031 (N_20031,N_10542,N_19971);
and U20032 (N_20032,N_13295,N_19730);
nand U20033 (N_20033,N_15641,N_16591);
xnor U20034 (N_20034,N_16303,N_14892);
nand U20035 (N_20035,N_12824,N_13422);
nand U20036 (N_20036,N_11952,N_12109);
and U20037 (N_20037,N_13963,N_18075);
or U20038 (N_20038,N_13378,N_15296);
or U20039 (N_20039,N_11084,N_17055);
nand U20040 (N_20040,N_19984,N_12517);
or U20041 (N_20041,N_18433,N_19070);
or U20042 (N_20042,N_10339,N_17998);
nand U20043 (N_20043,N_12268,N_15187);
and U20044 (N_20044,N_16405,N_10172);
nand U20045 (N_20045,N_13681,N_11825);
or U20046 (N_20046,N_13465,N_19016);
nor U20047 (N_20047,N_14887,N_11552);
nor U20048 (N_20048,N_12233,N_18377);
nand U20049 (N_20049,N_11649,N_17926);
and U20050 (N_20050,N_18867,N_13875);
and U20051 (N_20051,N_19962,N_10665);
nor U20052 (N_20052,N_16768,N_12110);
nand U20053 (N_20053,N_14500,N_11726);
and U20054 (N_20054,N_12407,N_15951);
or U20055 (N_20055,N_17106,N_11079);
or U20056 (N_20056,N_18342,N_12205);
or U20057 (N_20057,N_17892,N_11562);
or U20058 (N_20058,N_17980,N_12956);
nor U20059 (N_20059,N_11209,N_11239);
nor U20060 (N_20060,N_19780,N_14310);
and U20061 (N_20061,N_13810,N_12275);
nor U20062 (N_20062,N_14909,N_15826);
nor U20063 (N_20063,N_10119,N_19943);
nand U20064 (N_20064,N_10911,N_14692);
nor U20065 (N_20065,N_18220,N_18362);
or U20066 (N_20066,N_11994,N_12133);
or U20067 (N_20067,N_11648,N_13518);
nand U20068 (N_20068,N_16128,N_13568);
or U20069 (N_20069,N_15181,N_11222);
nand U20070 (N_20070,N_14176,N_12253);
nor U20071 (N_20071,N_14577,N_12269);
or U20072 (N_20072,N_10104,N_11859);
and U20073 (N_20073,N_13744,N_12601);
nor U20074 (N_20074,N_17612,N_18458);
nor U20075 (N_20075,N_16605,N_10718);
nand U20076 (N_20076,N_19471,N_12913);
nand U20077 (N_20077,N_12043,N_11001);
and U20078 (N_20078,N_17464,N_10652);
nor U20079 (N_20079,N_18750,N_18809);
or U20080 (N_20080,N_19221,N_19209);
and U20081 (N_20081,N_14959,N_10567);
and U20082 (N_20082,N_19431,N_16032);
nand U20083 (N_20083,N_13028,N_16949);
or U20084 (N_20084,N_13361,N_12095);
and U20085 (N_20085,N_16520,N_16814);
nand U20086 (N_20086,N_13989,N_15804);
or U20087 (N_20087,N_16261,N_10288);
xor U20088 (N_20088,N_13775,N_12583);
or U20089 (N_20089,N_15568,N_19718);
nor U20090 (N_20090,N_17823,N_16567);
and U20091 (N_20091,N_17152,N_14274);
nand U20092 (N_20092,N_15777,N_10977);
or U20093 (N_20093,N_19151,N_11325);
nand U20094 (N_20094,N_19452,N_13443);
nor U20095 (N_20095,N_18666,N_11512);
and U20096 (N_20096,N_15721,N_18719);
nor U20097 (N_20097,N_14113,N_16580);
xor U20098 (N_20098,N_16937,N_18005);
nor U20099 (N_20099,N_11220,N_12370);
and U20100 (N_20100,N_10532,N_11176);
nor U20101 (N_20101,N_13202,N_10502);
or U20102 (N_20102,N_11033,N_12187);
nor U20103 (N_20103,N_12970,N_10360);
nor U20104 (N_20104,N_10185,N_19442);
or U20105 (N_20105,N_17010,N_15082);
nor U20106 (N_20106,N_11959,N_16452);
and U20107 (N_20107,N_13799,N_11097);
nor U20108 (N_20108,N_16907,N_14174);
nand U20109 (N_20109,N_18691,N_19583);
and U20110 (N_20110,N_16073,N_12162);
or U20111 (N_20111,N_10160,N_11123);
nor U20112 (N_20112,N_12068,N_10703);
nor U20113 (N_20113,N_13303,N_13979);
nand U20114 (N_20114,N_13608,N_15027);
and U20115 (N_20115,N_18307,N_19034);
and U20116 (N_20116,N_13504,N_10755);
nor U20117 (N_20117,N_18873,N_14187);
and U20118 (N_20118,N_16687,N_18462);
nand U20119 (N_20119,N_10489,N_15774);
or U20120 (N_20120,N_19739,N_12936);
and U20121 (N_20121,N_17493,N_18281);
and U20122 (N_20122,N_14369,N_13476);
nor U20123 (N_20123,N_18733,N_10423);
or U20124 (N_20124,N_12156,N_15998);
nor U20125 (N_20125,N_17052,N_17377);
nand U20126 (N_20126,N_17525,N_15387);
and U20127 (N_20127,N_16354,N_13659);
nand U20128 (N_20128,N_16667,N_13734);
and U20129 (N_20129,N_16964,N_19251);
and U20130 (N_20130,N_10910,N_14855);
nor U20131 (N_20131,N_12121,N_19046);
and U20132 (N_20132,N_18519,N_14184);
or U20133 (N_20133,N_14664,N_16944);
and U20134 (N_20134,N_16828,N_18509);
nand U20135 (N_20135,N_11761,N_10709);
or U20136 (N_20136,N_12607,N_16871);
nand U20137 (N_20137,N_11835,N_19698);
nor U20138 (N_20138,N_14936,N_17869);
or U20139 (N_20139,N_10457,N_11993);
nand U20140 (N_20140,N_16169,N_12429);
nor U20141 (N_20141,N_13635,N_18793);
nand U20142 (N_20142,N_15415,N_11856);
nor U20143 (N_20143,N_18522,N_17291);
nand U20144 (N_20144,N_19256,N_14092);
nor U20145 (N_20145,N_16263,N_12488);
or U20146 (N_20146,N_13528,N_13582);
and U20147 (N_20147,N_14685,N_12695);
and U20148 (N_20148,N_17144,N_14493);
or U20149 (N_20149,N_12518,N_13732);
nor U20150 (N_20150,N_16272,N_13245);
nor U20151 (N_20151,N_12317,N_17366);
or U20152 (N_20152,N_19872,N_18246);
nand U20153 (N_20153,N_18909,N_19915);
nor U20154 (N_20154,N_11180,N_17994);
or U20155 (N_20155,N_19412,N_18243);
or U20156 (N_20156,N_17518,N_15791);
or U20157 (N_20157,N_12919,N_15557);
and U20158 (N_20158,N_16306,N_10663);
nor U20159 (N_20159,N_16463,N_19287);
and U20160 (N_20160,N_11102,N_10302);
nor U20161 (N_20161,N_15884,N_12418);
or U20162 (N_20162,N_12852,N_19688);
nor U20163 (N_20163,N_17629,N_16923);
and U20164 (N_20164,N_15202,N_13594);
or U20165 (N_20165,N_12290,N_10516);
nand U20166 (N_20166,N_16668,N_11367);
nor U20167 (N_20167,N_17127,N_12528);
and U20168 (N_20168,N_14464,N_15107);
nor U20169 (N_20169,N_16382,N_19793);
nor U20170 (N_20170,N_11638,N_14134);
nor U20171 (N_20171,N_16080,N_19916);
or U20172 (N_20172,N_13764,N_15106);
or U20173 (N_20173,N_17541,N_18613);
nor U20174 (N_20174,N_13238,N_12107);
and U20175 (N_20175,N_18860,N_15069);
or U20176 (N_20176,N_19634,N_16853);
and U20177 (N_20177,N_14436,N_16656);
or U20178 (N_20178,N_15469,N_15234);
nor U20179 (N_20179,N_10710,N_11331);
and U20180 (N_20180,N_18600,N_13018);
nor U20181 (N_20181,N_12765,N_18013);
nor U20182 (N_20182,N_11599,N_16832);
nand U20183 (N_20183,N_11685,N_11315);
nand U20184 (N_20184,N_12425,N_13633);
or U20185 (N_20185,N_11731,N_13144);
nand U20186 (N_20186,N_18847,N_12368);
nand U20187 (N_20187,N_12141,N_16782);
nand U20188 (N_20188,N_10705,N_17704);
nor U20189 (N_20189,N_15662,N_13816);
nand U20190 (N_20190,N_14489,N_17416);
and U20191 (N_20191,N_18024,N_11313);
and U20192 (N_20192,N_15821,N_17070);
nand U20193 (N_20193,N_15708,N_14398);
or U20194 (N_20194,N_19667,N_13736);
or U20195 (N_20195,N_17007,N_12566);
nand U20196 (N_20196,N_13501,N_11736);
nor U20197 (N_20197,N_14346,N_17725);
and U20198 (N_20198,N_19605,N_10589);
nor U20199 (N_20199,N_14713,N_14714);
nand U20200 (N_20200,N_14110,N_11434);
or U20201 (N_20201,N_19677,N_14632);
and U20202 (N_20202,N_12255,N_15205);
and U20203 (N_20203,N_18446,N_12892);
or U20204 (N_20204,N_17972,N_12018);
or U20205 (N_20205,N_19656,N_11181);
or U20206 (N_20206,N_17181,N_13027);
or U20207 (N_20207,N_12449,N_18440);
nand U20208 (N_20208,N_18837,N_11839);
and U20209 (N_20209,N_13226,N_18435);
nor U20210 (N_20210,N_10049,N_18604);
nand U20211 (N_20211,N_19042,N_10157);
or U20212 (N_20212,N_15006,N_13793);
nand U20213 (N_20213,N_16517,N_10308);
and U20214 (N_20214,N_14601,N_17941);
and U20215 (N_20215,N_12663,N_11378);
nor U20216 (N_20216,N_11285,N_17078);
or U20217 (N_20217,N_13461,N_17263);
nor U20218 (N_20218,N_19642,N_12232);
or U20219 (N_20219,N_17299,N_12432);
nor U20220 (N_20220,N_11692,N_15459);
nor U20221 (N_20221,N_13575,N_12013);
or U20222 (N_20222,N_11483,N_11364);
or U20223 (N_20223,N_16985,N_18850);
nand U20224 (N_20224,N_19906,N_10252);
and U20225 (N_20225,N_13511,N_13407);
nor U20226 (N_20226,N_16812,N_11444);
nor U20227 (N_20227,N_19530,N_18050);
and U20228 (N_20228,N_15214,N_13142);
or U20229 (N_20229,N_16010,N_11404);
or U20230 (N_20230,N_16242,N_12041);
nor U20231 (N_20231,N_13817,N_16495);
or U20232 (N_20232,N_19000,N_17064);
nor U20233 (N_20233,N_14704,N_10978);
and U20234 (N_20234,N_12788,N_10635);
and U20235 (N_20235,N_16062,N_14381);
nand U20236 (N_20236,N_19839,N_11980);
nor U20237 (N_20237,N_19982,N_18423);
or U20238 (N_20238,N_18137,N_13923);
nand U20239 (N_20239,N_16037,N_18306);
nand U20240 (N_20240,N_15577,N_12206);
nand U20241 (N_20241,N_16608,N_13348);
nor U20242 (N_20242,N_10646,N_15925);
nand U20243 (N_20243,N_13921,N_16981);
nand U20244 (N_20244,N_15513,N_14103);
or U20245 (N_20245,N_13399,N_18735);
nand U20246 (N_20246,N_11152,N_11253);
nand U20247 (N_20247,N_17765,N_19222);
and U20248 (N_20248,N_18193,N_18726);
and U20249 (N_20249,N_18263,N_15710);
nand U20250 (N_20250,N_15968,N_13757);
nand U20251 (N_20251,N_16940,N_16643);
or U20252 (N_20252,N_13743,N_19959);
nand U20253 (N_20253,N_10855,N_18775);
nor U20254 (N_20254,N_10420,N_18004);
and U20255 (N_20255,N_19666,N_10056);
nand U20256 (N_20256,N_17460,N_15455);
and U20257 (N_20257,N_15248,N_17895);
nor U20258 (N_20258,N_14677,N_13918);
nand U20259 (N_20259,N_19711,N_19383);
nor U20260 (N_20260,N_12748,N_12330);
or U20261 (N_20261,N_16683,N_11979);
and U20262 (N_20262,N_14011,N_10244);
or U20263 (N_20263,N_11850,N_10373);
nor U20264 (N_20264,N_13095,N_11436);
and U20265 (N_20265,N_13400,N_14856);
nor U20266 (N_20266,N_19162,N_11082);
or U20267 (N_20267,N_17017,N_14827);
and U20268 (N_20268,N_15518,N_19717);
and U20269 (N_20269,N_13163,N_10968);
nor U20270 (N_20270,N_10928,N_13972);
or U20271 (N_20271,N_14296,N_12096);
nand U20272 (N_20272,N_17424,N_13909);
and U20273 (N_20273,N_15651,N_19701);
xnor U20274 (N_20274,N_19296,N_19012);
nor U20275 (N_20275,N_18504,N_18833);
and U20276 (N_20276,N_17203,N_17953);
and U20277 (N_20277,N_16222,N_15948);
nand U20278 (N_20278,N_11073,N_12988);
nor U20279 (N_20279,N_14298,N_12951);
nand U20280 (N_20280,N_19650,N_17741);
nor U20281 (N_20281,N_18403,N_13453);
or U20282 (N_20282,N_11866,N_10437);
or U20283 (N_20283,N_15343,N_13859);
and U20284 (N_20284,N_14434,N_18674);
and U20285 (N_20285,N_13089,N_11245);
nor U20286 (N_20286,N_11138,N_16575);
or U20287 (N_20287,N_11504,N_15898);
and U20288 (N_20288,N_15918,N_14233);
or U20289 (N_20289,N_13887,N_16809);
or U20290 (N_20290,N_14029,N_19842);
nand U20291 (N_20291,N_13956,N_10095);
nor U20292 (N_20292,N_11153,N_10925);
nor U20293 (N_20293,N_18250,N_18607);
nor U20294 (N_20294,N_18799,N_17983);
and U20295 (N_20295,N_11957,N_15696);
nand U20296 (N_20296,N_19752,N_12085);
xor U20297 (N_20297,N_19153,N_13546);
nand U20298 (N_20298,N_12501,N_12863);
and U20299 (N_20299,N_12003,N_14263);
and U20300 (N_20300,N_18372,N_17217);
nand U20301 (N_20301,N_17485,N_10883);
nor U20302 (N_20302,N_14875,N_12752);
and U20303 (N_20303,N_13865,N_15330);
and U20304 (N_20304,N_18126,N_10544);
and U20305 (N_20305,N_10527,N_10551);
nand U20306 (N_20306,N_16323,N_16191);
and U20307 (N_20307,N_16371,N_14156);
nor U20308 (N_20308,N_15299,N_15342);
or U20309 (N_20309,N_15039,N_15920);
nand U20310 (N_20310,N_17531,N_15160);
nor U20311 (N_20311,N_10303,N_11007);
nand U20312 (N_20312,N_11203,N_10430);
or U20313 (N_20313,N_12777,N_13081);
nor U20314 (N_20314,N_16682,N_14358);
nor U20315 (N_20315,N_16255,N_18595);
nor U20316 (N_20316,N_15258,N_15716);
or U20317 (N_20317,N_12022,N_18664);
nand U20318 (N_20318,N_19481,N_10972);
nand U20319 (N_20319,N_13746,N_19898);
nand U20320 (N_20320,N_10281,N_16283);
nor U20321 (N_20321,N_10083,N_10647);
and U20322 (N_20322,N_11738,N_11252);
or U20323 (N_20323,N_17829,N_19294);
and U20324 (N_20324,N_14277,N_18027);
nor U20325 (N_20325,N_17922,N_17790);
nand U20326 (N_20326,N_11494,N_14882);
or U20327 (N_20327,N_14040,N_12912);
nand U20328 (N_20328,N_14534,N_19806);
or U20329 (N_20329,N_13408,N_19206);
or U20330 (N_20330,N_12670,N_18701);
nand U20331 (N_20331,N_16094,N_12678);
or U20332 (N_20332,N_16796,N_14622);
or U20333 (N_20333,N_15910,N_17326);
and U20334 (N_20334,N_12124,N_18185);
nand U20335 (N_20335,N_19630,N_18935);
nor U20336 (N_20336,N_12393,N_19434);
nor U20337 (N_20337,N_15573,N_14799);
and U20338 (N_20338,N_16176,N_13688);
or U20339 (N_20339,N_13165,N_14597);
nand U20340 (N_20340,N_13680,N_15403);
nor U20341 (N_20341,N_19304,N_12421);
or U20342 (N_20342,N_10720,N_14286);
nor U20343 (N_20343,N_16095,N_19678);
and U20344 (N_20344,N_15003,N_18951);
xor U20345 (N_20345,N_14897,N_18612);
and U20346 (N_20346,N_19154,N_10068);
and U20347 (N_20347,N_12885,N_11934);
and U20348 (N_20348,N_15864,N_18222);
and U20349 (N_20349,N_11016,N_18336);
nand U20350 (N_20350,N_13882,N_15575);
nor U20351 (N_20351,N_13969,N_10934);
and U20352 (N_20352,N_11336,N_16144);
nor U20353 (N_20353,N_10965,N_18728);
nand U20354 (N_20354,N_17774,N_12431);
and U20355 (N_20355,N_18532,N_11670);
and U20356 (N_20356,N_18670,N_16519);
nor U20357 (N_20357,N_18110,N_14266);
nand U20358 (N_20358,N_11144,N_10372);
nor U20359 (N_20359,N_10241,N_14846);
and U20360 (N_20360,N_11415,N_17315);
and U20361 (N_20361,N_18881,N_11184);
and U20362 (N_20362,N_15283,N_17373);
nand U20363 (N_20363,N_11855,N_16815);
and U20364 (N_20364,N_11191,N_19719);
or U20365 (N_20365,N_10467,N_12219);
nor U20366 (N_20366,N_12448,N_16802);
nor U20367 (N_20367,N_19449,N_10295);
nor U20368 (N_20368,N_10454,N_10594);
and U20369 (N_20369,N_19527,N_11369);
or U20370 (N_20370,N_16670,N_13225);
nor U20371 (N_20371,N_18197,N_11476);
and U20372 (N_20372,N_17176,N_19500);
nand U20373 (N_20373,N_19263,N_14899);
nand U20374 (N_20374,N_19243,N_14292);
or U20375 (N_20375,N_15508,N_18894);
and U20376 (N_20376,N_12231,N_15988);
nor U20377 (N_20377,N_12942,N_13006);
nand U20378 (N_20378,N_13751,N_15528);
nand U20379 (N_20379,N_18730,N_14302);
nor U20380 (N_20380,N_10315,N_16837);
xnor U20381 (N_20381,N_11889,N_18940);
or U20382 (N_20382,N_13493,N_16948);
nand U20383 (N_20383,N_15409,N_14129);
nor U20384 (N_20384,N_12955,N_16320);
nor U20385 (N_20385,N_12415,N_15657);
nand U20386 (N_20386,N_11339,N_10108);
and U20387 (N_20387,N_15043,N_17784);
nor U20388 (N_20388,N_15261,N_10109);
nor U20389 (N_20389,N_18716,N_14935);
and U20390 (N_20390,N_13778,N_12716);
and U20391 (N_20391,N_10679,N_14680);
or U20392 (N_20392,N_10946,N_12135);
nand U20393 (N_20393,N_14442,N_12900);
nand U20394 (N_20394,N_13088,N_15799);
or U20395 (N_20395,N_19712,N_13357);
and U20396 (N_20396,N_16705,N_15776);
or U20397 (N_20397,N_10908,N_13349);
and U20398 (N_20398,N_13730,N_19036);
nor U20399 (N_20399,N_15801,N_18541);
xnor U20400 (N_20400,N_11400,N_15077);
and U20401 (N_20401,N_15534,N_19413);
and U20402 (N_20402,N_17193,N_12559);
and U20403 (N_20403,N_19974,N_16841);
nand U20404 (N_20404,N_16881,N_12782);
nor U20405 (N_20405,N_12465,N_14874);
nand U20406 (N_20406,N_19241,N_19435);
nor U20407 (N_20407,N_19836,N_12014);
and U20408 (N_20408,N_11608,N_10633);
nor U20409 (N_20409,N_12651,N_13779);
nand U20410 (N_20410,N_11255,N_17896);
or U20411 (N_20411,N_17305,N_11732);
nand U20412 (N_20412,N_14318,N_16984);
nor U20413 (N_20413,N_18605,N_13428);
and U20414 (N_20414,N_12247,N_13665);
nand U20415 (N_20415,N_16436,N_15159);
or U20416 (N_20416,N_13061,N_10634);
nand U20417 (N_20417,N_11657,N_15896);
and U20418 (N_20418,N_16071,N_12949);
nor U20419 (N_20419,N_10677,N_12277);
nor U20420 (N_20420,N_13241,N_12481);
and U20421 (N_20421,N_17242,N_17839);
nand U20422 (N_20422,N_18035,N_14140);
nor U20423 (N_20423,N_12442,N_15808);
or U20424 (N_20424,N_18866,N_10260);
nand U20425 (N_20425,N_11679,N_17380);
and U20426 (N_20426,N_10917,N_13919);
or U20427 (N_20427,N_14957,N_19182);
nor U20428 (N_20428,N_17686,N_13391);
or U20429 (N_20429,N_17944,N_13851);
nor U20430 (N_20430,N_14484,N_17251);
nand U20431 (N_20431,N_16297,N_19416);
nor U20432 (N_20432,N_11585,N_19592);
and U20433 (N_20433,N_16978,N_13913);
or U20434 (N_20434,N_16322,N_18025);
nand U20435 (N_20435,N_10477,N_16686);
or U20436 (N_20436,N_11143,N_14056);
nand U20437 (N_20437,N_13090,N_12971);
or U20438 (N_20438,N_15763,N_13403);
and U20439 (N_20439,N_11517,N_17183);
and U20440 (N_20440,N_17477,N_18157);
and U20441 (N_20441,N_13544,N_15288);
nand U20442 (N_20442,N_13886,N_16794);
nor U20443 (N_20443,N_12379,N_13469);
or U20444 (N_20444,N_10803,N_17474);
nor U20445 (N_20445,N_10630,N_13074);
nor U20446 (N_20446,N_14256,N_16501);
nor U20447 (N_20447,N_11307,N_10022);
or U20448 (N_20448,N_10044,N_11019);
and U20449 (N_20449,N_18817,N_17247);
nor U20450 (N_20450,N_14421,N_17337);
nand U20451 (N_20451,N_10047,N_11495);
nor U20452 (N_20452,N_12193,N_18871);
and U20453 (N_20453,N_17509,N_15530);
or U20454 (N_20454,N_15357,N_10074);
and U20455 (N_20455,N_13950,N_19053);
nand U20456 (N_20456,N_15157,N_13647);
and U20457 (N_20457,N_18655,N_18346);
nor U20458 (N_20458,N_19059,N_16123);
or U20459 (N_20459,N_10541,N_16883);
or U20460 (N_20460,N_14842,N_15210);
nor U20461 (N_20461,N_14463,N_10576);
and U20462 (N_20462,N_14071,N_10891);
and U20463 (N_20463,N_11514,N_12775);
or U20464 (N_20464,N_10903,N_17256);
nor U20465 (N_20465,N_13794,N_13726);
or U20466 (N_20466,N_17693,N_15828);
or U20467 (N_20467,N_15450,N_19320);
and U20468 (N_20468,N_16108,N_10818);
nor U20469 (N_20469,N_12471,N_15670);
and U20470 (N_20470,N_14787,N_14996);
nor U20471 (N_20471,N_18695,N_13797);
nor U20472 (N_20472,N_11049,N_10805);
nand U20473 (N_20473,N_11845,N_12024);
nand U20474 (N_20474,N_16831,N_17554);
nand U20475 (N_20475,N_16084,N_19186);
nor U20476 (N_20476,N_16976,N_16471);
and U20477 (N_20477,N_19691,N_16906);
nor U20478 (N_20478,N_18191,N_19755);
xor U20479 (N_20479,N_13611,N_17018);
or U20480 (N_20480,N_12020,N_17559);
and U20481 (N_20481,N_12793,N_19208);
nand U20482 (N_20482,N_16989,N_15977);
and U20483 (N_20483,N_17746,N_12300);
or U20484 (N_20484,N_18428,N_13293);
nand U20485 (N_20485,N_10788,N_18152);
nand U20486 (N_20486,N_14451,N_12577);
and U20487 (N_20487,N_12893,N_17089);
or U20488 (N_20488,N_19450,N_18389);
nand U20489 (N_20489,N_18888,N_16661);
or U20490 (N_20490,N_19710,N_15348);
nor U20491 (N_20491,N_17884,N_13227);
or U20492 (N_20492,N_13836,N_15772);
nand U20493 (N_20493,N_14759,N_11626);
and U20494 (N_20494,N_18105,N_12183);
nand U20495 (N_20495,N_14158,N_18966);
or U20496 (N_20496,N_19043,N_17919);
nand U20497 (N_20497,N_12688,N_15426);
or U20498 (N_20498,N_13415,N_11801);
nor U20499 (N_20499,N_16194,N_13526);
or U20500 (N_20500,N_10649,N_16170);
or U20501 (N_20501,N_15973,N_19664);
nor U20502 (N_20502,N_13618,N_19851);
nor U20503 (N_20503,N_19968,N_10490);
and U20504 (N_20504,N_15011,N_12204);
or U20505 (N_20505,N_13555,N_17549);
or U20506 (N_20506,N_18396,N_18070);
or U20507 (N_20507,N_19545,N_10696);
or U20508 (N_20508,N_16380,N_15295);
and U20509 (N_20509,N_17874,N_13041);
and U20510 (N_20510,N_16206,N_13500);
nor U20511 (N_20511,N_10379,N_18079);
and U20512 (N_20512,N_18536,N_14976);
and U20513 (N_20513,N_12426,N_11916);
xnor U20514 (N_20514,N_15743,N_14417);
nand U20515 (N_20515,N_13749,N_18348);
or U20516 (N_20516,N_18308,N_10833);
nor U20517 (N_20517,N_13248,N_10382);
or U20518 (N_20518,N_16227,N_19703);
nor U20519 (N_20519,N_13801,N_13845);
xor U20520 (N_20520,N_11396,N_12932);
nand U20521 (N_20521,N_13976,N_12721);
nor U20522 (N_20522,N_12582,N_14516);
and U20523 (N_20523,N_10800,N_18777);
nand U20524 (N_20524,N_11273,N_19185);
nand U20525 (N_20525,N_10470,N_19461);
nor U20526 (N_20526,N_13644,N_15349);
nor U20527 (N_20527,N_14299,N_17899);
nor U20528 (N_20528,N_13258,N_10539);
or U20529 (N_20529,N_10632,N_10948);
nor U20530 (N_20530,N_17066,N_17755);
or U20531 (N_20531,N_10767,N_19069);
nand U20532 (N_20532,N_15803,N_18326);
nor U20533 (N_20533,N_11527,N_14797);
nor U20534 (N_20534,N_14425,N_13529);
nor U20535 (N_20535,N_12858,N_13143);
and U20536 (N_20536,N_12147,N_19290);
and U20537 (N_20537,N_11070,N_14430);
or U20538 (N_20538,N_18477,N_10258);
or U20539 (N_20539,N_18554,N_16641);
nor U20540 (N_20540,N_14845,N_12647);
nor U20541 (N_20541,N_11256,N_14760);
or U20542 (N_20542,N_14626,N_14227);
and U20543 (N_20543,N_16811,N_19991);
or U20544 (N_20544,N_18514,N_12485);
nand U20545 (N_20545,N_17513,N_10954);
nand U20546 (N_20546,N_15779,N_14331);
nor U20547 (N_20547,N_12336,N_14699);
nor U20548 (N_20548,N_16134,N_14885);
nand U20549 (N_20549,N_17471,N_17840);
nor U20550 (N_20550,N_17616,N_12922);
nor U20551 (N_20551,N_13628,N_13970);
and U20552 (N_20552,N_19098,N_18333);
nand U20553 (N_20553,N_19697,N_19265);
nand U20554 (N_20554,N_10535,N_19096);
nor U20555 (N_20555,N_15219,N_10992);
or U20556 (N_20556,N_14209,N_14046);
and U20557 (N_20557,N_11428,N_19179);
nor U20558 (N_20558,N_15474,N_13748);
nand U20559 (N_20559,N_11793,N_15916);
nand U20560 (N_20560,N_15223,N_10105);
or U20561 (N_20561,N_17696,N_18919);
and U20562 (N_20562,N_16168,N_10272);
nand U20563 (N_20563,N_11593,N_19727);
or U20564 (N_20564,N_11235,N_18097);
or U20565 (N_20565,N_18767,N_16783);
nand U20566 (N_20566,N_14039,N_13048);
or U20567 (N_20567,N_18366,N_14988);
or U20568 (N_20568,N_17602,N_11217);
or U20569 (N_20569,N_10424,N_13747);
nand U20570 (N_20570,N_12700,N_12258);
nor U20571 (N_20571,N_14416,N_13233);
or U20572 (N_20572,N_16639,N_19557);
nor U20573 (N_20573,N_13934,N_18190);
and U20574 (N_20574,N_17348,N_18374);
or U20575 (N_20575,N_19498,N_17885);
or U20576 (N_20576,N_17766,N_16711);
or U20577 (N_20577,N_16307,N_16792);
and U20578 (N_20578,N_10672,N_15752);
or U20579 (N_20579,N_18155,N_12004);
or U20580 (N_20580,N_11680,N_13944);
or U20581 (N_20581,N_15890,N_17621);
or U20582 (N_20582,N_18911,N_17752);
nand U20583 (N_20583,N_17800,N_16963);
nand U20584 (N_20584,N_18581,N_14775);
nor U20585 (N_20585,N_14940,N_10826);
and U20586 (N_20586,N_19829,N_12769);
nand U20587 (N_20587,N_17325,N_13581);
nor U20588 (N_20588,N_13650,N_16779);
and U20589 (N_20589,N_17274,N_15026);
nor U20590 (N_20590,N_17608,N_14678);
nor U20591 (N_20591,N_13080,N_16150);
or U20592 (N_20592,N_10257,N_15682);
nor U20593 (N_20593,N_17981,N_18165);
or U20594 (N_20594,N_13452,N_13494);
nand U20595 (N_20595,N_18801,N_14053);
nor U20596 (N_20596,N_16561,N_14244);
or U20597 (N_20597,N_11357,N_16087);
and U20598 (N_20598,N_12920,N_14530);
nand U20599 (N_20599,N_16726,N_14089);
or U20600 (N_20600,N_17657,N_13762);
and U20601 (N_20601,N_17003,N_15341);
and U20602 (N_20602,N_15639,N_18186);
and U20603 (N_20603,N_14225,N_17259);
nand U20604 (N_20604,N_12238,N_12962);
and U20605 (N_20605,N_18009,N_11529);
nand U20606 (N_20606,N_17226,N_17041);
nand U20607 (N_20607,N_15883,N_15231);
and U20608 (N_20608,N_11709,N_10361);
or U20609 (N_20609,N_15758,N_17792);
nand U20610 (N_20610,N_14947,N_12221);
nor U20611 (N_20611,N_10892,N_19031);
nand U20612 (N_20612,N_16339,N_12184);
and U20613 (N_20613,N_19216,N_13496);
nand U20614 (N_20614,N_10897,N_18431);
and U20615 (N_20615,N_15183,N_15386);
and U20616 (N_20616,N_11885,N_16347);
nand U20617 (N_20617,N_14171,N_17042);
nand U20618 (N_20618,N_10919,N_13521);
and U20619 (N_20619,N_15561,N_10953);
or U20620 (N_20620,N_14117,N_16910);
nor U20621 (N_20621,N_12470,N_15631);
and U20622 (N_20622,N_11725,N_11412);
and U20623 (N_20623,N_10760,N_18018);
and U20624 (N_20624,N_19879,N_18773);
and U20625 (N_20625,N_10132,N_18912);
nor U20626 (N_20626,N_12409,N_10650);
nor U20627 (N_20627,N_17768,N_19888);
and U20628 (N_20628,N_18011,N_10124);
nor U20629 (N_20629,N_11609,N_17143);
and U20630 (N_20630,N_14456,N_13375);
nand U20631 (N_20631,N_10553,N_16935);
or U20632 (N_20632,N_16763,N_12977);
and U20633 (N_20633,N_15212,N_10827);
nand U20634 (N_20634,N_13002,N_15309);
and U20635 (N_20635,N_10114,N_14466);
or U20636 (N_20636,N_16158,N_14951);
or U20637 (N_20637,N_15381,N_13770);
or U20638 (N_20638,N_17960,N_18284);
and U20639 (N_20639,N_18053,N_11140);
and U20640 (N_20640,N_19074,N_19372);
nand U20641 (N_20641,N_17717,N_10008);
nand U20642 (N_20642,N_19674,N_11461);
and U20643 (N_20643,N_15270,N_18772);
nand U20644 (N_20644,N_14272,N_15017);
nand U20645 (N_20645,N_16574,N_19821);
nor U20646 (N_20646,N_17387,N_13087);
nand U20647 (N_20647,N_11223,N_18040);
nor U20648 (N_20648,N_13098,N_18065);
and U20649 (N_20649,N_12106,N_18119);
and U20650 (N_20650,N_13181,N_17757);
or U20651 (N_20651,N_16035,N_12975);
nor U20652 (N_20652,N_10043,N_10206);
nor U20653 (N_20653,N_13204,N_13796);
or U20654 (N_20654,N_14317,N_15751);
and U20655 (N_20655,N_10517,N_17952);
nand U20656 (N_20656,N_16916,N_16256);
nand U20657 (N_20657,N_13850,N_10480);
nand U20658 (N_20658,N_18120,N_12272);
and U20659 (N_20659,N_13768,N_11356);
and U20660 (N_20660,N_15407,N_17058);
or U20661 (N_20661,N_13803,N_13830);
nand U20662 (N_20662,N_19765,N_14517);
and U20663 (N_20663,N_11791,N_17799);
or U20664 (N_20664,N_14758,N_10115);
nand U20665 (N_20665,N_13302,N_19559);
or U20666 (N_20666,N_12059,N_18117);
nand U20667 (N_20667,N_14824,N_13252);
and U20668 (N_20668,N_14487,N_12745);
nor U20669 (N_20669,N_15303,N_19052);
nand U20670 (N_20670,N_10961,N_13239);
nor U20671 (N_20671,N_12747,N_14433);
nand U20672 (N_20672,N_11664,N_17938);
nor U20673 (N_20673,N_19351,N_14222);
and U20674 (N_20674,N_12792,N_13372);
and U20675 (N_20675,N_10342,N_18332);
nand U20676 (N_20676,N_17698,N_11697);
and U20677 (N_20677,N_17711,N_16507);
or U20678 (N_20678,N_11869,N_12821);
xor U20679 (N_20679,N_16395,N_15355);
nor U20680 (N_20680,N_15421,N_17910);
nand U20681 (N_20681,N_15493,N_18128);
or U20682 (N_20682,N_14324,N_18690);
or U20683 (N_20683,N_11940,N_15088);
nand U20684 (N_20684,N_15132,N_16759);
and U20685 (N_20685,N_14257,N_11511);
or U20686 (N_20686,N_19606,N_16627);
or U20687 (N_20687,N_17065,N_14008);
nand U20688 (N_20688,N_18016,N_13219);
nor U20689 (N_20689,N_17750,N_17573);
nor U20690 (N_20690,N_11898,N_18949);
and U20691 (N_20691,N_15384,N_17534);
or U20692 (N_20692,N_13056,N_18295);
nor U20693 (N_20693,N_19947,N_18754);
or U20694 (N_20694,N_17632,N_10867);
nor U20695 (N_20695,N_17077,N_18334);
nand U20696 (N_20696,N_10927,N_10870);
or U20697 (N_20697,N_11295,N_17128);
nor U20698 (N_20698,N_10221,N_17031);
nor U20699 (N_20699,N_18132,N_19456);
or U20700 (N_20700,N_19673,N_11410);
nand U20701 (N_20701,N_15759,N_12192);
nand U20702 (N_20702,N_10053,N_11370);
or U20703 (N_20703,N_15277,N_11257);
or U20704 (N_20704,N_18234,N_10882);
nand U20705 (N_20705,N_10096,N_11840);
nand U20706 (N_20706,N_13626,N_16543);
or U20707 (N_20707,N_11386,N_19009);
nand U20708 (N_20708,N_16264,N_14288);
nand U20709 (N_20709,N_11347,N_17167);
and U20710 (N_20710,N_15111,N_17544);
nand U20711 (N_20711,N_15750,N_19486);
or U20712 (N_20712,N_19139,N_16882);
nand U20713 (N_20713,N_16889,N_19084);
and U20714 (N_20714,N_17520,N_19169);
nand U20715 (N_20715,N_15378,N_17378);
and U20716 (N_20716,N_14673,N_14486);
or U20717 (N_20717,N_12930,N_15780);
and U20718 (N_20718,N_15084,N_15488);
and U20719 (N_20719,N_12514,N_14483);
nand U20720 (N_20720,N_17778,N_12604);
xnor U20721 (N_20721,N_17304,N_15729);
nand U20722 (N_20722,N_12543,N_10763);
xor U20723 (N_20723,N_17202,N_15914);
nand U20724 (N_20724,N_18094,N_15519);
and U20725 (N_20725,N_10017,N_12890);
nor U20726 (N_20726,N_17776,N_10144);
nand U20727 (N_20727,N_10005,N_11063);
and U20728 (N_20728,N_19980,N_19356);
and U20729 (N_20729,N_10441,N_17817);
and U20730 (N_20730,N_16250,N_15185);
or U20731 (N_20731,N_15440,N_14055);
or U20732 (N_20732,N_14206,N_15775);
nor U20733 (N_20733,N_16967,N_17641);
and U20734 (N_20734,N_12395,N_19518);
nand U20735 (N_20735,N_19453,N_17740);
nor U20736 (N_20736,N_13257,N_18759);
xnor U20737 (N_20737,N_13464,N_14034);
nand U20738 (N_20738,N_17671,N_11863);
nand U20739 (N_20739,N_13046,N_17100);
and U20740 (N_20740,N_17788,N_18875);
and U20741 (N_20741,N_12538,N_11792);
nor U20742 (N_20742,N_10485,N_11949);
or U20743 (N_20743,N_15480,N_16911);
and U20744 (N_20744,N_17905,N_11036);
and U20745 (N_20745,N_18558,N_14987);
and U20746 (N_20746,N_19313,N_13583);
nor U20747 (N_20747,N_11757,N_16550);
and U20748 (N_20748,N_16748,N_19922);
nand U20749 (N_20749,N_14150,N_18515);
and U20750 (N_20750,N_18617,N_18311);
nor U20751 (N_20751,N_12789,N_12836);
or U20752 (N_20752,N_17780,N_11080);
and U20753 (N_20753,N_16196,N_13971);
and U20754 (N_20754,N_11557,N_14968);
nand U20755 (N_20755,N_18427,N_11263);
or U20756 (N_20756,N_13034,N_14809);
nor U20757 (N_20757,N_16226,N_19509);
or U20758 (N_20758,N_10698,N_11012);
nor U20759 (N_20759,N_17845,N_19973);
and U20760 (N_20760,N_16835,N_15311);
or U20761 (N_20761,N_10294,N_11614);
nand U20762 (N_20762,N_15013,N_17330);
and U20763 (N_20763,N_18839,N_14610);
or U20764 (N_20764,N_16117,N_19570);
nand U20765 (N_20765,N_18104,N_19715);
nor U20766 (N_20766,N_13077,N_15760);
or U20767 (N_20767,N_10497,N_12571);
and U20768 (N_20768,N_10617,N_12216);
nand U20769 (N_20769,N_19862,N_15520);
nor U20770 (N_20770,N_11700,N_11536);
nor U20771 (N_20771,N_14226,N_15848);
nand U20772 (N_20772,N_16908,N_19007);
or U20773 (N_20773,N_19112,N_14726);
and U20774 (N_20774,N_13949,N_17441);
or U20775 (N_20775,N_17319,N_11450);
nand U20776 (N_20776,N_15572,N_19466);
nor U20777 (N_20777,N_11630,N_12215);
and U20778 (N_20778,N_11158,N_11927);
and U20779 (N_20779,N_16462,N_16791);
or U20780 (N_20780,N_18404,N_12997);
nor U20781 (N_20781,N_11175,N_15218);
nand U20782 (N_20782,N_16706,N_13863);
or U20783 (N_20783,N_16358,N_14106);
nor U20784 (N_20784,N_11581,N_18599);
or U20785 (N_20785,N_10407,N_14703);
nand U20786 (N_20786,N_13658,N_16660);
nand U20787 (N_20787,N_18896,N_16869);
nor U20788 (N_20788,N_16532,N_10495);
nand U20789 (N_20789,N_17341,N_13477);
nor U20790 (N_20790,N_12230,N_15892);
or U20791 (N_20791,N_10752,N_19083);
or U20792 (N_20792,N_14542,N_11605);
and U20793 (N_20793,N_19324,N_15858);
nor U20794 (N_20794,N_17113,N_12325);
and U20795 (N_20795,N_18327,N_11770);
and U20796 (N_20796,N_19708,N_13980);
and U20797 (N_20797,N_15465,N_17111);
nor U20798 (N_20798,N_16966,N_18038);
or U20799 (N_20799,N_14544,N_15955);
nor U20800 (N_20800,N_11787,N_10493);
nor U20801 (N_20801,N_17045,N_19266);
and U20802 (N_20802,N_16650,N_19550);
and U20803 (N_20803,N_15807,N_13593);
nor U20804 (N_20804,N_14037,N_14068);
nor U20805 (N_20805,N_16279,N_11518);
nand U20806 (N_20806,N_12917,N_10697);
and U20807 (N_20807,N_14686,N_19668);
and U20808 (N_20808,N_12040,N_11321);
nand U20809 (N_20809,N_17871,N_11038);
and U20810 (N_20810,N_16075,N_17352);
nand U20811 (N_20811,N_16821,N_15649);
or U20812 (N_20812,N_10920,N_15057);
or U20813 (N_20813,N_12495,N_18747);
or U20814 (N_20814,N_17609,N_16749);
or U20815 (N_20815,N_18694,N_18312);
nor U20816 (N_20816,N_17357,N_11789);
and U20817 (N_20817,N_15859,N_12783);
and U20818 (N_20818,N_12115,N_16560);
nor U20819 (N_20819,N_16657,N_17085);
or U20820 (N_20820,N_19966,N_13447);
or U20821 (N_20821,N_11242,N_14070);
nor U20822 (N_20822,N_11422,N_16531);
nor U20823 (N_20823,N_11112,N_10197);
and U20824 (N_20824,N_15148,N_11301);
nand U20825 (N_20825,N_18265,N_14519);
nor U20826 (N_20826,N_16741,N_15693);
or U20827 (N_20827,N_12489,N_13881);
and U20828 (N_20828,N_13685,N_12270);
and U20829 (N_20829,N_17396,N_18627);
nand U20830 (N_20830,N_16511,N_11086);
nor U20831 (N_20831,N_17311,N_18824);
or U20832 (N_20832,N_14762,N_12385);
nand U20833 (N_20833,N_12654,N_19212);
or U20834 (N_20834,N_15906,N_11701);
nor U20835 (N_20835,N_14119,N_17576);
xor U20836 (N_20836,N_19205,N_12036);
and U20837 (N_20837,N_17140,N_16015);
and U20838 (N_20838,N_12797,N_11615);
nor U20839 (N_20839,N_13605,N_16926);
or U20840 (N_20840,N_13198,N_13051);
nor U20841 (N_20841,N_17909,N_17177);
or U20842 (N_20842,N_16830,N_14332);
nand U20843 (N_20843,N_16797,N_11320);
nor U20844 (N_20844,N_12692,N_16658);
nor U20845 (N_20845,N_19533,N_19195);
or U20846 (N_20846,N_19721,N_12818);
and U20847 (N_20847,N_14269,N_16166);
or U20848 (N_20848,N_12334,N_19824);
xnor U20849 (N_20849,N_18274,N_16649);
or U20850 (N_20850,N_11823,N_17294);
nand U20851 (N_20851,N_11941,N_13828);
nor U20852 (N_20852,N_14970,N_14477);
nand U20853 (N_20853,N_15194,N_12522);
nor U20854 (N_20854,N_19813,N_15882);
and U20855 (N_20855,N_14854,N_15886);
nor U20856 (N_20856,N_13878,N_16739);
or U20857 (N_20857,N_18381,N_16994);
and U20858 (N_20858,N_19423,N_11040);
nand U20859 (N_20859,N_13912,N_15650);
nor U20860 (N_20860,N_13481,N_11119);
or U20861 (N_20861,N_14293,N_11204);
or U20862 (N_20862,N_16564,N_18975);
nor U20863 (N_20863,N_10700,N_19763);
or U20864 (N_20864,N_10660,N_10102);
or U20865 (N_20865,N_12062,N_12308);
and U20866 (N_20866,N_12596,N_17769);
nand U20867 (N_20867,N_17297,N_10193);
and U20868 (N_20868,N_17189,N_10048);
nand U20869 (N_20869,N_18748,N_10605);
nor U20870 (N_20870,N_15536,N_10087);
and U20871 (N_20871,N_12328,N_12029);
nand U20872 (N_20872,N_17894,N_12980);
nor U20873 (N_20873,N_13292,N_17714);
and U20874 (N_20874,N_15325,N_10349);
or U20875 (N_20875,N_14735,N_11942);
or U20876 (N_20876,N_17701,N_11081);
and U20877 (N_20877,N_17642,N_15905);
nand U20878 (N_20878,N_15902,N_16494);
and U20879 (N_20879,N_18616,N_11681);
nor U20880 (N_20880,N_14255,N_16527);
or U20881 (N_20881,N_17945,N_12830);
nor U20882 (N_20882,N_12496,N_15121);
and U20883 (N_20883,N_14821,N_10453);
nand U20884 (N_20884,N_14214,N_17585);
nand U20885 (N_20885,N_12015,N_18278);
or U20886 (N_20886,N_12033,N_11448);
and U20887 (N_20887,N_16052,N_19920);
nor U20888 (N_20888,N_13263,N_19956);
and U20889 (N_20889,N_17133,N_11053);
or U20890 (N_20890,N_14036,N_15067);
and U20891 (N_20891,N_14934,N_13755);
nor U20892 (N_20892,N_19389,N_15140);
and U20893 (N_20893,N_12738,N_14731);
and U20894 (N_20894,N_18082,N_16536);
and U20895 (N_20895,N_18355,N_16775);
or U20896 (N_20896,N_13948,N_10735);
nor U20897 (N_20897,N_10822,N_18471);
nor U20898 (N_20898,N_12741,N_19190);
or U20899 (N_20899,N_12766,N_18318);
nor U20900 (N_20900,N_13522,N_15940);
or U20901 (N_20901,N_15204,N_11028);
and U20902 (N_20902,N_19350,N_12314);
and U20903 (N_20903,N_14005,N_11883);
nand U20904 (N_20904,N_11746,N_10267);
and U20905 (N_20905,N_13780,N_16383);
nor U20906 (N_20906,N_11774,N_11417);
and U20907 (N_20907,N_19616,N_10898);
or U20908 (N_20908,N_19346,N_16430);
xor U20909 (N_20909,N_12197,N_10355);
nand U20910 (N_20910,N_16157,N_12623);
nor U20911 (N_20911,N_11131,N_12427);
and U20912 (N_20912,N_18800,N_14149);
or U20913 (N_20913,N_12761,N_13959);
and U20914 (N_20914,N_14465,N_12503);
or U20915 (N_20915,N_15769,N_10645);
nand U20916 (N_20916,N_11219,N_16562);
nor U20917 (N_20917,N_16876,N_15216);
or U20918 (N_20918,N_16281,N_14235);
or U20919 (N_20919,N_19230,N_14729);
nor U20920 (N_20920,N_12873,N_17195);
and U20921 (N_20921,N_16252,N_13639);
nand U20922 (N_20922,N_12921,N_17006);
or U20923 (N_20923,N_17853,N_10942);
nand U20924 (N_20924,N_17546,N_15147);
or U20925 (N_20925,N_14667,N_18813);
or U20926 (N_20926,N_18408,N_11547);
and U20927 (N_20927,N_19957,N_12191);
nand U20928 (N_20928,N_14344,N_17374);
nor U20929 (N_20929,N_15475,N_15644);
nor U20930 (N_20930,N_18071,N_13509);
nor U20931 (N_20931,N_10070,N_12257);
and U20932 (N_20932,N_18526,N_12527);
nor U20933 (N_20933,N_14932,N_18745);
or U20934 (N_20934,N_17075,N_11676);
nor U20935 (N_20935,N_18464,N_15264);
nor U20936 (N_20936,N_15628,N_10518);
and U20937 (N_20937,N_19814,N_12784);
nor U20938 (N_20938,N_18508,N_17875);
nand U20939 (N_20939,N_10940,N_14308);
nor U20940 (N_20940,N_17432,N_15158);
nand U20941 (N_20941,N_17379,N_10015);
nor U20942 (N_20942,N_12005,N_13393);
or U20943 (N_20943,N_11146,N_13769);
nand U20944 (N_20944,N_12486,N_11425);
nand U20945 (N_20945,N_17439,N_19832);
or U20946 (N_20946,N_11198,N_18609);
or U20947 (N_20947,N_12610,N_19946);
nor U20948 (N_20948,N_17619,N_15598);
nand U20949 (N_20949,N_10584,N_11185);
nand U20950 (N_20950,N_15420,N_10959);
nor U20951 (N_20951,N_10028,N_17071);
nor U20952 (N_20952,N_11749,N_16675);
and U20953 (N_20953,N_18924,N_10852);
nand U20954 (N_20954,N_15734,N_11708);
or U20955 (N_20955,N_12653,N_11913);
and U20956 (N_20956,N_11718,N_16500);
or U20957 (N_20957,N_19749,N_14368);
nand U20958 (N_20958,N_15703,N_19369);
nor U20959 (N_20959,N_16026,N_12335);
nand U20960 (N_20960,N_10526,N_13965);
and U20961 (N_20961,N_17486,N_11526);
nor U20962 (N_20962,N_12322,N_19907);
or U20963 (N_20963,N_17484,N_15458);
or U20964 (N_20964,N_13695,N_10163);
and U20965 (N_20965,N_15677,N_14535);
and U20966 (N_20966,N_17438,N_14405);
and U20967 (N_20967,N_15872,N_12774);
nor U20968 (N_20968,N_19005,N_14229);
nor U20969 (N_20969,N_19037,N_13904);
nand U20970 (N_20970,N_13288,N_13216);
nor U20971 (N_20971,N_11366,N_14779);
or U20972 (N_20972,N_17175,N_11932);
nand U20973 (N_20973,N_17815,N_10601);
and U20974 (N_20974,N_10039,N_15073);
or U20975 (N_20975,N_13451,N_12867);
nand U20976 (N_20976,N_11946,N_16444);
nor U20977 (N_20977,N_18506,N_19905);
and U20978 (N_20978,N_14007,N_12249);
nand U20979 (N_20979,N_16487,N_10192);
or U20980 (N_20980,N_13926,N_18160);
or U20981 (N_20981,N_12943,N_18316);
or U20982 (N_20982,N_17917,N_14636);
and U20983 (N_20983,N_18945,N_12602);
nor U20984 (N_20984,N_16356,N_19060);
nor U20985 (N_20985,N_11688,N_16793);
nand U20986 (N_20986,N_16718,N_11510);
or U20987 (N_20987,N_17327,N_12252);
nand U20988 (N_20988,N_10340,N_14387);
and U20989 (N_20989,N_12086,N_11598);
nand U20990 (N_20990,N_11077,N_16360);
or U20991 (N_20991,N_16558,N_19484);
or U20992 (N_20992,N_19704,N_10156);
nand U20993 (N_20993,N_14989,N_13299);
nand U20994 (N_20994,N_13108,N_18227);
and U20995 (N_20995,N_14000,N_18648);
or U20996 (N_20996,N_19468,N_11992);
and U20997 (N_20997,N_19496,N_10658);
or U20998 (N_20998,N_10498,N_19960);
or U20999 (N_20999,N_19860,N_16208);
nand U21000 (N_21000,N_11767,N_17626);
nand U21001 (N_21001,N_19648,N_10628);
or U21002 (N_21002,N_14189,N_11478);
nand U21003 (N_21003,N_16457,N_15308);
nand U21004 (N_21004,N_13931,N_12946);
nor U21005 (N_21005,N_14675,N_19379);
and U21006 (N_21006,N_14144,N_13029);
nand U21007 (N_21007,N_19852,N_11981);
nor U21008 (N_21008,N_13625,N_19121);
nor U21009 (N_21009,N_11758,N_13194);
nand U21010 (N_21010,N_16887,N_15314);
nor U21011 (N_21011,N_12177,N_14159);
and U21012 (N_21012,N_17742,N_13564);
and U21013 (N_21013,N_13157,N_16450);
nor U21014 (N_21014,N_12819,N_11973);
and U21015 (N_21015,N_15938,N_18095);
nor U21016 (N_21016,N_11302,N_11843);
or U21017 (N_21017,N_14723,N_15953);
nor U21018 (N_21018,N_17644,N_19868);
nand U21019 (N_21019,N_13371,N_17762);
nor U21020 (N_21020,N_15100,N_17809);
nor U21021 (N_21021,N_19662,N_14549);
and U21022 (N_21022,N_12346,N_19815);
nand U21023 (N_21023,N_11723,N_18687);
nor U21024 (N_21024,N_14307,N_18453);
and U21025 (N_21025,N_16103,N_10009);
or U21026 (N_21026,N_10458,N_10683);
or U21027 (N_21027,N_10426,N_10590);
nor U21028 (N_21028,N_10329,N_19487);
and U21029 (N_21029,N_11747,N_13446);
and U21030 (N_21030,N_16690,N_10860);
nor U21031 (N_21031,N_17147,N_16101);
and U21032 (N_21032,N_11374,N_17826);
nor U21033 (N_21033,N_15999,N_18671);
or U21034 (N_21034,N_11048,N_18530);
nand U21035 (N_21035,N_14228,N_19692);
and U21036 (N_21036,N_18787,N_15595);
or U21037 (N_21037,N_11603,N_17744);
nand U21038 (N_21038,N_15704,N_17257);
nand U21039 (N_21039,N_16673,N_16262);
nor U21040 (N_21040,N_18409,N_12994);
nor U21041 (N_21041,N_19792,N_14700);
and U21042 (N_21042,N_11437,N_17343);
or U21043 (N_21043,N_11069,N_14309);
nor U21044 (N_21044,N_12534,N_18091);
nor U21045 (N_21045,N_10552,N_13763);
nor U21046 (N_21046,N_15857,N_13632);
nand U21047 (N_21047,N_13405,N_18953);
or U21048 (N_21048,N_17333,N_13696);
nand U21049 (N_21049,N_17976,N_12472);
and U21050 (N_21050,N_15642,N_19568);
nand U21051 (N_21051,N_10831,N_18280);
and U21052 (N_21052,N_11962,N_19775);
and U21053 (N_21053,N_11194,N_14321);
nand U21054 (N_21054,N_19424,N_16633);
nand U21055 (N_21055,N_19760,N_11035);
and U21056 (N_21056,N_12565,N_12925);
nand U21057 (N_21057,N_17563,N_10421);
xor U21058 (N_21058,N_16400,N_13120);
and U21059 (N_21059,N_11684,N_19107);
nand U21060 (N_21060,N_10301,N_13387);
nor U21061 (N_21061,N_14021,N_11443);
and U21062 (N_21062,N_16175,N_19078);
and U21063 (N_21063,N_10513,N_14102);
and U21064 (N_21064,N_17630,N_16091);
or U21065 (N_21065,N_19969,N_19215);
and U21066 (N_21066,N_12112,N_13615);
nor U21067 (N_21067,N_13047,N_14628);
and U21068 (N_21068,N_12586,N_18400);
nand U21069 (N_21069,N_14199,N_14792);
or U21070 (N_21070,N_13319,N_12474);
nand U21071 (N_21071,N_15952,N_17268);
nand U21072 (N_21072,N_13384,N_17281);
or U21073 (N_21073,N_12154,N_13113);
nor U21074 (N_21074,N_12451,N_19899);
nor U21075 (N_21075,N_15604,N_13729);
or U21076 (N_21076,N_16595,N_13021);
nor U21077 (N_21077,N_15957,N_11202);
nor U21078 (N_21078,N_14715,N_17461);
nor U21079 (N_21079,N_15449,N_13065);
nand U21080 (N_21080,N_11027,N_14471);
and U21081 (N_21081,N_13140,N_16085);
or U21082 (N_21082,N_15560,N_13304);
or U21083 (N_21083,N_11296,N_13307);
and U21084 (N_21084,N_15773,N_17283);
or U21085 (N_21085,N_18908,N_10712);
nand U21086 (N_21086,N_15786,N_19699);
nand U21087 (N_21087,N_16847,N_17413);
and U21088 (N_21088,N_16417,N_16098);
nand U21089 (N_21089,N_18414,N_18715);
nand U21090 (N_21090,N_14900,N_10751);
nand U21091 (N_21091,N_11910,N_10641);
or U21092 (N_21092,N_14547,N_15060);
and U21093 (N_21093,N_11641,N_18493);
or U21094 (N_21094,N_18835,N_15798);
nor U21095 (N_21095,N_10859,N_15685);
nand U21096 (N_21096,N_10376,N_12399);
and U21097 (N_21097,N_18330,N_15897);
nor U21098 (N_21098,N_16611,N_10569);
nor U21099 (N_21099,N_11447,N_13958);
nor U21100 (N_21100,N_18476,N_11472);
or U21101 (N_21101,N_12699,N_14997);
or U21102 (N_21102,N_12315,N_12152);
nor U21103 (N_21103,N_13565,N_19122);
nand U21104 (N_21104,N_10823,N_12972);
and U21105 (N_21105,N_15756,N_19607);
or U21106 (N_21106,N_15030,N_15558);
or U21107 (N_21107,N_15806,N_18391);
nand U21108 (N_21108,N_11466,N_10981);
and U21109 (N_21109,N_12105,N_19103);
nor U21110 (N_21110,N_16186,N_14192);
and U21111 (N_21111,N_13715,N_14178);
nor U21112 (N_21112,N_13280,N_14281);
and U21113 (N_21113,N_10209,N_15899);
nand U21114 (N_21114,N_15095,N_18989);
nor U21115 (N_21115,N_10408,N_14764);
nor U21116 (N_21116,N_19733,N_17842);
nand U21117 (N_21117,N_19878,N_17376);
and U21118 (N_21118,N_11224,N_11595);
or U21119 (N_21119,N_12241,N_18046);
nor U21120 (N_21120,N_17138,N_12352);
nand U21121 (N_21121,N_17032,N_10071);
and U21122 (N_21122,N_18556,N_13502);
nand U21123 (N_21123,N_19194,N_11822);
or U21124 (N_21124,N_10116,N_15714);
and U21125 (N_21125,N_11604,N_17161);
or U21126 (N_21126,N_15856,N_11602);
and U21127 (N_21127,N_19264,N_16331);
and U21128 (N_21128,N_17855,N_18782);
nor U21129 (N_21129,N_18885,N_15680);
nor U21130 (N_21130,N_15610,N_13621);
and U21131 (N_21131,N_16270,N_15128);
or U21132 (N_21132,N_16044,N_15586);
or U21133 (N_21133,N_11678,N_14902);
or U21134 (N_21134,N_11929,N_12273);
and U21135 (N_21135,N_13153,N_18608);
or U21136 (N_21136,N_10253,N_18751);
or U21137 (N_21137,N_14136,N_13914);
nor U21138 (N_21138,N_19040,N_14502);
nand U21139 (N_21139,N_11921,N_18272);
nor U21140 (N_21140,N_16388,N_10135);
nor U21141 (N_21141,N_19534,N_13109);
and U21142 (N_21142,N_12616,N_13468);
and U21143 (N_21143,N_13409,N_17287);
or U21144 (N_21144,N_19996,N_17785);
and U21145 (N_21145,N_15051,N_13826);
and U21146 (N_21146,N_11553,N_15031);
nor U21147 (N_21147,N_14647,N_18780);
nor U21148 (N_21148,N_13620,N_18317);
and U21149 (N_21149,N_10359,N_16377);
nor U21150 (N_21150,N_15994,N_18305);
and U21151 (N_21151,N_18974,N_19903);
nand U21152 (N_21152,N_13661,N_15253);
nand U21153 (N_21153,N_11300,N_14920);
and U21154 (N_21154,N_17937,N_19884);
or U21155 (N_21155,N_11365,N_10512);
nand U21156 (N_21156,N_18329,N_14898);
and U21157 (N_21157,N_15293,N_13591);
and U21158 (N_21158,N_17519,N_11124);
or U21159 (N_21159,N_11031,N_12553);
and U21160 (N_21160,N_14551,N_16980);
nor U21161 (N_21161,N_15180,N_12089);
and U21162 (N_21162,N_11055,N_12881);
and U21163 (N_21163,N_10782,N_19510);
xor U21164 (N_21164,N_11556,N_14131);
or U21165 (N_21165,N_18049,N_10347);
or U21166 (N_21166,N_14707,N_15514);
nor U21167 (N_21167,N_18064,N_10774);
and U21168 (N_21168,N_17192,N_18216);
nand U21169 (N_21169,N_12122,N_16901);
nand U21170 (N_21170,N_18643,N_17918);
nor U21171 (N_21171,N_12828,N_17532);
or U21172 (N_21172,N_12061,N_19840);
or U21173 (N_21173,N_13019,N_19297);
nand U21174 (N_21174,N_17810,N_16483);
and U21175 (N_21175,N_17827,N_19398);
nand U21176 (N_21176,N_13441,N_16486);
and U21177 (N_21177,N_19555,N_15269);
or U21178 (N_21178,N_17572,N_15653);
nand U21179 (N_21179,N_17716,N_11982);
and U21180 (N_21180,N_18682,N_11200);
or U21181 (N_21181,N_17713,N_15544);
nor U21182 (N_21182,N_11902,N_14826);
nor U21183 (N_21183,N_11005,N_10381);
or U21184 (N_21184,N_12069,N_13266);
xor U21185 (N_21185,N_11148,N_19085);
nor U21186 (N_21186,N_14232,N_14407);
nor U21187 (N_21187,N_18358,N_16467);
and U21188 (N_21188,N_16033,N_10159);
nor U21189 (N_21189,N_17335,N_12286);
nand U21190 (N_21190,N_19856,N_13277);
or U21191 (N_21191,N_17101,N_16549);
and U21192 (N_21192,N_14734,N_19728);
and U21193 (N_21193,N_10561,N_11613);
or U21194 (N_21194,N_15722,N_13519);
and U21195 (N_21195,N_12817,N_19569);
nand U21196 (N_21196,N_11188,N_17249);
and U21197 (N_21197,N_16850,N_15850);
or U21198 (N_21198,N_11010,N_19245);
or U21199 (N_21199,N_12428,N_10766);
nor U21200 (N_21200,N_10716,N_14666);
or U21201 (N_21201,N_11421,N_19483);
and U21202 (N_21202,N_11108,N_16665);
nor U21203 (N_21203,N_13874,N_11164);
or U21204 (N_21204,N_10386,N_19641);
nor U21205 (N_21205,N_16839,N_13152);
or U21206 (N_21206,N_18276,N_14972);
nand U21207 (N_21207,N_15700,N_14093);
nand U21208 (N_21208,N_14819,N_11832);
nor U21209 (N_21209,N_10618,N_17092);
or U21210 (N_21210,N_14894,N_15021);
nand U21211 (N_21211,N_16230,N_13316);
and U21212 (N_21212,N_18761,N_10328);
or U21213 (N_21213,N_11689,N_19713);
and U21214 (N_21214,N_11323,N_18727);
nor U21215 (N_21215,N_10973,N_15291);
or U21216 (N_21216,N_18698,N_11247);
nor U21217 (N_21217,N_14839,N_13312);
nand U21218 (N_21218,N_14424,N_11157);
nand U21219 (N_21219,N_12344,N_13294);
nor U21220 (N_21220,N_19827,N_10422);
nand U21221 (N_21221,N_10452,N_19115);
nor U21222 (N_21222,N_16943,N_13355);
or U21223 (N_21223,N_18535,N_10974);
nand U21224 (N_21224,N_15496,N_15551);
or U21225 (N_21225,N_14345,N_16153);
nor U21226 (N_21226,N_10175,N_14743);
nand U21227 (N_21227,N_16603,N_10504);
and U21228 (N_21228,N_12362,N_19291);
or U21229 (N_21229,N_13964,N_17877);
and U21230 (N_21230,N_14223,N_11548);
and U21231 (N_21231,N_15117,N_19006);
or U21232 (N_21232,N_15761,N_19612);
nand U21233 (N_21233,N_10343,N_11282);
nor U21234 (N_21234,N_13689,N_19013);
and U21235 (N_21235,N_19433,N_19970);
nor U21236 (N_21236,N_13381,N_18383);
and U21237 (N_21237,N_13733,N_10311);
nand U21238 (N_21238,N_11473,N_12714);
nor U21239 (N_21239,N_19177,N_15438);
nor U21240 (N_21240,N_14914,N_17131);
and U21241 (N_21241,N_12998,N_16592);
and U21242 (N_21242,N_11919,N_18823);
nor U21243 (N_21243,N_18313,N_16368);
nor U21244 (N_21244,N_10727,N_19426);
nand U21245 (N_21245,N_19854,N_10184);
and U21246 (N_21246,N_11703,N_15425);
nand U21247 (N_21247,N_12351,N_16651);
and U21248 (N_21248,N_19978,N_17254);
nor U21249 (N_21249,N_19571,N_15340);
nor U21250 (N_21250,N_10798,N_15887);
nor U21251 (N_21251,N_10353,N_13414);
nor U21252 (N_21252,N_17427,N_12573);
nand U21253 (N_21253,N_15326,N_14861);
nand U21254 (N_21254,N_14123,N_19590);
nor U21255 (N_21255,N_15377,N_16449);
and U21256 (N_21256,N_19777,N_14377);
or U21257 (N_21257,N_15790,N_10657);
and U21258 (N_21258,N_12088,N_17073);
and U21259 (N_21259,N_11818,N_13852);
or U21260 (N_21260,N_17224,N_14054);
and U21261 (N_21261,N_14162,N_12608);
nor U21262 (N_21262,N_12008,N_14399);
or U21263 (N_21263,N_12967,N_10045);
nand U21264 (N_21264,N_17347,N_16622);
and U21265 (N_21265,N_19964,N_15470);
nor U21266 (N_21266,N_12645,N_19087);
and U21267 (N_21267,N_18789,N_14524);
or U21268 (N_21268,N_16404,N_14640);
or U21269 (N_21269,N_19865,N_10089);
or U21270 (N_21270,N_19019,N_16465);
nor U21271 (N_21271,N_10032,N_18518);
or U21272 (N_21272,N_16664,N_12476);
or U21273 (N_21273,N_15737,N_18876);
and U21274 (N_21274,N_18029,N_18459);
and U21275 (N_21275,N_18081,N_16064);
and U21276 (N_21276,N_14795,N_14057);
nand U21277 (N_21277,N_18002,N_19176);
nand U21278 (N_21278,N_14955,N_16171);
or U21279 (N_21279,N_13691,N_11879);
and U21280 (N_21280,N_10276,N_17260);
or U21281 (N_21281,N_16106,N_10153);
nor U21282 (N_21282,N_17210,N_19823);
nor U21283 (N_21283,N_14728,N_10263);
nor U21284 (N_21284,N_17245,N_19300);
and U21285 (N_21285,N_14168,N_14305);
and U21286 (N_21286,N_14639,N_15056);
nand U21287 (N_21287,N_19929,N_18319);
nor U21288 (N_21288,N_10026,N_17340);
and U21289 (N_21289,N_13742,N_14670);
nor U21290 (N_21290,N_11238,N_19252);
or U21291 (N_21291,N_14600,N_17209);
and U21292 (N_21292,N_15328,N_19588);
nand U21293 (N_21293,N_16273,N_11897);
nand U21294 (N_21294,N_10171,N_14566);
nand U21295 (N_21295,N_10037,N_10801);
or U21296 (N_21296,N_18335,N_13431);
and U21297 (N_21297,N_17392,N_10982);
or U21298 (N_21298,N_18478,N_13323);
or U21299 (N_21299,N_10725,N_17962);
nor U21300 (N_21300,N_11135,N_18981);
xnor U21301 (N_21301,N_15730,N_17156);
nand U21302 (N_21302,N_15439,N_12023);
and U21303 (N_21303,N_17931,N_13512);
or U21304 (N_21304,N_10431,N_15323);
and U21305 (N_21305,N_16469,N_18129);
or U21306 (N_21306,N_13127,N_17469);
nand U21307 (N_21307,N_15636,N_16348);
nor U21308 (N_21308,N_16553,N_19882);
and U21309 (N_21309,N_18510,N_13313);
nand U21310 (N_21310,N_14665,N_16827);
nand U21311 (N_21311,N_19254,N_13727);
nor U21312 (N_21312,N_11167,N_14693);
or U21313 (N_21313,N_16598,N_15265);
nor U21314 (N_21314,N_18337,N_16357);
or U21315 (N_21315,N_12938,N_14496);
or U21316 (N_21316,N_16302,N_10921);
nor U21317 (N_21317,N_15089,N_19624);
nand U21318 (N_21318,N_14155,N_15462);
nor U21319 (N_21319,N_12291,N_16470);
or U21320 (N_21320,N_16258,N_13840);
or U21321 (N_21321,N_12544,N_11706);
or U21322 (N_21322,N_15478,N_18922);
or U21323 (N_21323,N_19425,N_19493);
and U21324 (N_21324,N_10824,N_16411);
nand U21325 (N_21325,N_17001,N_12979);
nor U21326 (N_21326,N_19613,N_19056);
and U21327 (N_21327,N_14532,N_12795);
and U21328 (N_21328,N_14924,N_14221);
nor U21329 (N_21329,N_14323,N_17253);
nand U21330 (N_21330,N_11468,N_18399);
or U21331 (N_21331,N_14545,N_14512);
and U21332 (N_21332,N_13364,N_13030);
nor U21333 (N_21333,N_19686,N_10886);
or U21334 (N_21334,N_19363,N_14182);
nor U21335 (N_21335,N_19816,N_10316);
and U21336 (N_21336,N_12358,N_13456);
and U21337 (N_21337,N_14490,N_10644);
nand U21338 (N_21338,N_10255,N_10729);
or U21339 (N_21339,N_18815,N_13932);
and U21340 (N_21340,N_17044,N_16554);
and U21341 (N_21341,N_14491,N_15419);
nand U21342 (N_21342,N_18540,N_18848);
and U21343 (N_21343,N_16801,N_12952);
nor U21344 (N_21344,N_12394,N_19023);
nor U21345 (N_21345,N_17783,N_18786);
or U21346 (N_21346,N_13599,N_13154);
nand U21347 (N_21347,N_11878,N_12071);
nor U21348 (N_21348,N_17662,N_18704);
nor U21349 (N_21349,N_18910,N_11303);
nand U21350 (N_21350,N_16485,N_10460);
and U21351 (N_21351,N_10896,N_13894);
nor U21352 (N_21352,N_19967,N_11060);
nor U21353 (N_21353,N_13986,N_11326);
or U21354 (N_21354,N_16642,N_12756);
nor U21355 (N_21355,N_16986,N_13099);
or U21356 (N_21356,N_19825,N_12021);
or U21357 (N_21357,N_11663,N_18846);
or U21358 (N_21358,N_14859,N_13787);
nand U21359 (N_21359,N_11888,N_12401);
nor U21360 (N_21360,N_19203,N_12625);
nand U21361 (N_21361,N_16736,N_17220);
or U21362 (N_21362,N_16872,N_11454);
nor U21363 (N_21363,N_10250,N_12691);
nand U21364 (N_21364,N_18345,N_16920);
or U21365 (N_21365,N_17243,N_14284);
nand U21366 (N_21366,N_17155,N_19638);
and U21367 (N_21367,N_14418,N_14946);
nand U21368 (N_21368,N_14851,N_14336);
nand U21369 (N_21369,N_17269,N_18739);
and U21370 (N_21370,N_17943,N_16572);
nand U21371 (N_21371,N_19011,N_13470);
nand U21372 (N_21372,N_10772,N_15487);
or U21373 (N_21373,N_15825,N_13513);
nor U21374 (N_21374,N_13673,N_11667);
nor U21375 (N_21375,N_10198,N_18495);
nor U21376 (N_21376,N_13269,N_17391);
nand U21377 (N_21377,N_19049,N_16582);
or U21378 (N_21378,N_15457,N_17097);
nand U21379 (N_21379,N_16180,N_17538);
and U21380 (N_21380,N_16890,N_12306);
nor U21381 (N_21381,N_10999,N_11462);
nand U21382 (N_21382,N_11159,N_17425);
or U21383 (N_21383,N_10050,N_13495);
or U21384 (N_21384,N_15623,N_14403);
or U21385 (N_21385,N_12803,N_13892);
or U21386 (N_21386,N_15504,N_11796);
or U21387 (N_21387,N_10055,N_18651);
or U21388 (N_21388,N_10025,N_15004);
xor U21389 (N_21389,N_10560,N_17405);
nand U21390 (N_21390,N_19782,N_14419);
and U21391 (N_21391,N_11844,N_12816);
and U21392 (N_21392,N_13124,N_18597);
nand U21393 (N_21393,N_17759,N_15178);
nand U21394 (N_21394,N_15945,N_10370);
nand U21395 (N_21395,N_13062,N_10265);
nor U21396 (N_21396,N_19138,N_10293);
or U21397 (N_21397,N_19747,N_12657);
or U21398 (N_21398,N_13135,N_18259);
or U21399 (N_21399,N_17412,N_15571);
and U21400 (N_21400,N_12367,N_12927);
nand U21401 (N_21401,N_18181,N_16496);
nor U21402 (N_21402,N_15622,N_10811);
and U21403 (N_21403,N_17975,N_19332);
nor U21404 (N_21404,N_14776,N_17234);
and U21405 (N_21405,N_17027,N_11064);
or U21406 (N_21406,N_18141,N_16345);
and U21407 (N_21407,N_18640,N_15179);
xnor U21408 (N_21408,N_13846,N_17591);
and U21409 (N_21409,N_16447,N_14543);
and U21410 (N_21410,N_18321,N_12049);
nor U21411 (N_21411,N_13880,N_11128);
nor U21412 (N_21412,N_14739,N_13331);
and U21413 (N_21413,N_14588,N_12207);
nand U21414 (N_21414,N_17775,N_16151);
and U21415 (N_21415,N_18479,N_18422);
xor U21416 (N_21416,N_12510,N_13784);
and U21417 (N_21417,N_11162,N_15345);
and U21418 (N_21418,N_11037,N_16076);
and U21419 (N_21419,N_17465,N_16414);
nor U21420 (N_21420,N_11197,N_13068);
and U21421 (N_21421,N_16546,N_16597);
or U21422 (N_21422,N_10390,N_13547);
and U21423 (N_21423,N_17649,N_16849);
nand U21424 (N_21424,N_13498,N_11520);
or U21425 (N_21425,N_19061,N_15684);
or U21426 (N_21426,N_19268,N_18764);
or U21427 (N_21427,N_15980,N_11880);
or U21428 (N_21428,N_13574,N_13645);
and U21429 (N_21429,N_12077,N_13609);
and U21430 (N_21430,N_16022,N_11882);
nand U21431 (N_21431,N_15634,N_18301);
nand U21432 (N_21432,N_16614,N_18564);
nor U21433 (N_21433,N_18802,N_14455);
and U21434 (N_21434,N_17103,N_19505);
nand U21435 (N_21435,N_18057,N_14431);
or U21436 (N_21436,N_16109,N_12924);
nor U21437 (N_21437,N_10875,N_15154);
and U21438 (N_21438,N_11456,N_10332);
nand U21439 (N_21439,N_18586,N_17942);
or U21440 (N_21440,N_11939,N_10979);
nand U21441 (N_21441,N_13774,N_17672);
and U21442 (N_21442,N_12603,N_15175);
nand U21443 (N_21443,N_13270,N_11743);
or U21444 (N_21444,N_15909,N_18971);
nand U21445 (N_21445,N_12019,N_15150);
or U21446 (N_21446,N_10462,N_12274);
nor U21447 (N_21447,N_14618,N_18455);
and U21448 (N_21448,N_10190,N_15927);
nor U21449 (N_21449,N_11419,N_15996);
nor U21450 (N_21450,N_19497,N_16918);
and U21451 (N_21451,N_11964,N_13792);
nand U21452 (N_21452,N_18622,N_18629);
nor U21453 (N_21453,N_16110,N_14197);
nand U21454 (N_21454,N_10357,N_15924);
nor U21455 (N_21455,N_14857,N_10680);
or U21456 (N_21456,N_13112,N_10685);
and U21457 (N_21457,N_13167,N_17473);
and U21458 (N_21458,N_18468,N_12390);
nand U21459 (N_21459,N_10708,N_10520);
xnor U21460 (N_21460,N_13855,N_19063);
nor U21461 (N_21461,N_19998,N_19726);
and U21462 (N_21462,N_10871,N_19150);
or U21463 (N_21463,N_17301,N_15666);
or U21464 (N_21464,N_13262,N_18729);
or U21465 (N_21465,N_18350,N_10640);
or U21466 (N_21466,N_19417,N_11229);
nor U21467 (N_21467,N_17207,N_17881);
and U21468 (N_21468,N_14270,N_13668);
nor U21469 (N_21469,N_17735,N_19409);
nor U21470 (N_21470,N_10863,N_18781);
or U21471 (N_21471,N_11006,N_11430);
and U21472 (N_21472,N_19738,N_17807);
nand U21473 (N_21473,N_12148,N_10162);
or U21474 (N_21474,N_10743,N_19689);
nand U21475 (N_21475,N_14806,N_18380);
or U21476 (N_21476,N_16819,N_16587);
nor U21477 (N_21477,N_14367,N_13119);
and U21478 (N_21478,N_13942,N_19573);
nand U21479 (N_21479,N_14173,N_18904);
nand U21480 (N_21480,N_12278,N_13941);
and U21481 (N_21481,N_19393,N_15974);
nand U21482 (N_21482,N_12222,N_14264);
and U21483 (N_21483,N_15366,N_11671);
nor U21484 (N_21484,N_15129,N_17684);
and U21485 (N_21485,N_19410,N_10167);
nand U21486 (N_21486,N_10274,N_16248);
or U21487 (N_21487,N_17115,N_15163);
nand U21488 (N_21488,N_15453,N_17252);
and U21489 (N_21489,N_16866,N_12304);
and U21490 (N_21490,N_12170,N_17979);
and U21491 (N_21491,N_18933,N_12311);
or U21492 (N_21492,N_17499,N_15990);
or U21493 (N_21493,N_15742,N_16762);
and U21494 (N_21494,N_19436,N_13631);
and U21495 (N_21495,N_19100,N_17037);
nand U21496 (N_21496,N_15492,N_10219);
nand U21497 (N_21497,N_17939,N_19694);
nor U21498 (N_21498,N_18618,N_13078);
nand U21499 (N_21499,N_18454,N_16977);
nor U21500 (N_21500,N_17372,N_12895);
nand U21501 (N_21501,N_14373,N_12804);
nor U21502 (N_21502,N_17540,N_19239);
nand U21503 (N_21503,N_19362,N_15526);
nor U21504 (N_21504,N_16201,N_16393);
and U21505 (N_21505,N_13663,N_13766);
nand U21506 (N_21506,N_16445,N_15764);
and U21507 (N_21507,N_15145,N_15611);
or U21508 (N_21508,N_16350,N_19774);
or U21509 (N_21509,N_17650,N_18534);
or U21510 (N_21510,N_17236,N_12575);
nor U21511 (N_21511,N_14979,N_13536);
nor U21512 (N_21512,N_14994,N_19828);
nor U21513 (N_21513,N_17021,N_12377);
and U21514 (N_21514,N_15811,N_16482);
nand U21515 (N_21515,N_19469,N_17504);
nand U21516 (N_21516,N_19522,N_14977);
and U21517 (N_21517,N_13994,N_12212);
nor U21518 (N_21518,N_18201,N_10861);
nand U21519 (N_21519,N_11686,N_13423);
and U21520 (N_21520,N_14637,N_11727);
and U21521 (N_21521,N_12001,N_10636);
nor U21522 (N_21522,N_15074,N_15336);
or U21523 (N_21523,N_12512,N_14777);
nor U21524 (N_21524,N_14638,N_11660);
nor U21525 (N_21525,N_15284,N_13643);
nor U21526 (N_21526,N_13988,N_19474);
and U21527 (N_21527,N_11587,N_12871);
and U21528 (N_21528,N_12743,N_13096);
or U21529 (N_21529,N_19965,N_11390);
nor U21530 (N_21530,N_16515,N_11333);
or U21531 (N_21531,N_14505,N_16353);
or U21532 (N_21532,N_16930,N_16856);
xor U21533 (N_21533,N_17011,N_15437);
nor U21534 (N_21534,N_10031,N_13907);
nor U21535 (N_21535,N_13543,N_11655);
nand U21536 (N_21536,N_12079,N_18183);
or U21537 (N_21537,N_16343,N_15161);
and U21538 (N_21538,N_13735,N_12569);
nand U21539 (N_21539,N_12228,N_13374);
or U21540 (N_21540,N_17739,N_18821);
or U21541 (N_21541,N_17652,N_17689);
nor U21542 (N_21542,N_15671,N_16316);
nand U21543 (N_21543,N_14064,N_17516);
xor U21544 (N_21544,N_18134,N_17836);
or U21545 (N_21545,N_12173,N_10016);
or U21546 (N_21546,N_11549,N_13440);
nor U21547 (N_21547,N_16027,N_11936);
nor U21548 (N_21548,N_13683,N_10842);
nand U21549 (N_21549,N_11072,N_17966);
nand U21550 (N_21550,N_12285,N_16375);
or U21551 (N_21551,N_19506,N_18108);
nand U21552 (N_21552,N_17230,N_14711);
nor U21553 (N_21553,N_18577,N_17164);
nand U21554 (N_21554,N_10041,N_18356);
nand U21555 (N_21555,N_15191,N_11228);
nand U21556 (N_21556,N_15259,N_13707);
and U21557 (N_21557,N_15958,N_13879);
and U21558 (N_21558,N_17049,N_15400);
or U21559 (N_21559,N_19577,N_11870);
or U21560 (N_21560,N_14392,N_12083);
nor U21561 (N_21561,N_18112,N_12028);
and U21562 (N_21562,N_11754,N_13017);
nand U21563 (N_21563,N_11647,N_11380);
nand U21564 (N_21564,N_14488,N_11142);
or U21565 (N_21565,N_12916,N_17346);
or U21566 (N_21566,N_17009,N_19621);
nor U21567 (N_21567,N_18143,N_10674);
and U21568 (N_21568,N_13206,N_10365);
and U21569 (N_21569,N_14873,N_19219);
and U21570 (N_21570,N_17510,N_16234);
nand U21571 (N_21571,N_17906,N_11464);
nand U21572 (N_21572,N_19068,N_11955);
and U21573 (N_21573,N_13767,N_10655);
or U21574 (N_21574,N_10706,N_15533);
nand U21575 (N_21575,N_18543,N_18229);
and U21576 (N_21576,N_16072,N_12366);
nor U21577 (N_21577,N_16586,N_11795);
or U21578 (N_21578,N_11368,N_18520);
or U21579 (N_21579,N_17959,N_10180);
or U21580 (N_21580,N_12973,N_13570);
and U21581 (N_21581,N_19843,N_19033);
nand U21582 (N_21582,N_18010,N_10218);
or U21583 (N_21583,N_12659,N_19189);
and U21584 (N_21584,N_14752,N_10269);
xnor U21585 (N_21585,N_15249,N_13436);
nand U21586 (N_21586,N_14536,N_13086);
xnor U21587 (N_21587,N_12519,N_17683);
and U21588 (N_21588,N_12876,N_18533);
nor U21589 (N_21589,N_14312,N_10011);
or U21590 (N_21590,N_14903,N_17593);
nor U21591 (N_21591,N_14886,N_12389);
or U21592 (N_21592,N_13079,N_16956);
nand U21593 (N_21593,N_14065,N_17114);
and U21594 (N_21594,N_18998,N_13596);
and U21595 (N_21595,N_17796,N_17091);
and U21596 (N_21596,N_13282,N_17456);
nor U21597 (N_21597,N_18900,N_18268);
and U21598 (N_21598,N_15796,N_15411);
nor U21599 (N_21599,N_17797,N_15431);
nand U21600 (N_21600,N_17197,N_10140);
and U21601 (N_21601,N_12165,N_17908);
nor U21602 (N_21602,N_18709,N_17476);
or U21603 (N_21603,N_11925,N_14230);
nor U21604 (N_21604,N_11173,N_10412);
and U21605 (N_21605,N_15599,N_10220);
and U21606 (N_21606,N_15559,N_15565);
nand U21607 (N_21607,N_19271,N_13106);
nand U21608 (N_21608,N_12347,N_19382);
or U21609 (N_21609,N_14635,N_12153);
and U21610 (N_21610,N_11730,N_16418);
and U21611 (N_21611,N_17248,N_10595);
or U21612 (N_21612,N_10849,N_17270);
and U21613 (N_21613,N_11306,N_18228);
or U21614 (N_21614,N_17599,N_15646);
nand U21615 (N_21615,N_13145,N_15956);
nand U21616 (N_21616,N_17417,N_14443);
nand U21617 (N_21617,N_17096,N_18254);
and U21618 (N_21618,N_19891,N_10051);
xor U21619 (N_21619,N_16195,N_19997);
nand U21620 (N_21620,N_19598,N_16335);
and U21621 (N_21621,N_11433,N_18489);
and U21622 (N_21622,N_11408,N_18589);
and U21623 (N_21623,N_10599,N_13902);
nor U21624 (N_21624,N_10139,N_16362);
and U21625 (N_21625,N_11193,N_11947);
nor U21626 (N_21626,N_16129,N_11311);
nor U21627 (N_21627,N_11958,N_14732);
or U21628 (N_21628,N_19632,N_18054);
and U21629 (N_21629,N_10014,N_12357);
nand U21630 (N_21630,N_18401,N_18466);
nor U21631 (N_21631,N_11088,N_14437);
and U21632 (N_21632,N_15301,N_19517);
nor U21633 (N_21633,N_11763,N_14917);
nand U21634 (N_21634,N_13847,N_19260);
and U21635 (N_21635,N_18689,N_19201);
nand U21636 (N_21636,N_16401,N_11156);
or U21637 (N_21637,N_17012,N_12965);
and U21638 (N_21638,N_14382,N_16808);
and U21639 (N_21639,N_18090,N_18784);
nor U21640 (N_21640,N_16361,N_12843);
and U21641 (N_21641,N_17054,N_19408);
and U21642 (N_21642,N_17530,N_12327);
nand U21643 (N_21643,N_19651,N_17638);
and U21644 (N_21644,N_15934,N_12696);
and U21645 (N_21645,N_13842,N_16655);
and U21646 (N_21646,N_10440,N_18646);
or U21647 (N_21647,N_14613,N_19388);
nor U21648 (N_21648,N_12324,N_14672);
and U21649 (N_21649,N_12644,N_19341);
and U21650 (N_21650,N_15134,N_14379);
nor U21651 (N_21651,N_13180,N_16304);
and U21652 (N_21652,N_11995,N_13937);
nand U21653 (N_21653,N_17595,N_17231);
or U21654 (N_21654,N_17828,N_10608);
or U21655 (N_21655,N_16429,N_18827);
nand U21656 (N_21656,N_19937,N_11141);
nor U21657 (N_21657,N_13133,N_18561);
nor U21658 (N_21658,N_15402,N_15135);
or U21659 (N_21659,N_10568,N_10319);
nand U21660 (N_21660,N_13438,N_19327);
or U21661 (N_21661,N_14325,N_19223);
and U21662 (N_21662,N_11244,N_19317);
nand U21663 (N_21663,N_10519,N_13720);
nand U21664 (N_21664,N_13434,N_18857);
or U21665 (N_21665,N_13883,N_14183);
nand U21666 (N_21666,N_10802,N_19459);
and U21667 (N_21667,N_17812,N_16105);
and U21668 (N_21668,N_13217,N_18096);
nand U21669 (N_21669,N_13242,N_13341);
or U21670 (N_21670,N_19072,N_15304);
or U21671 (N_21671,N_14528,N_13786);
nor U21672 (N_21672,N_17887,N_15114);
xor U21673 (N_21673,N_18283,N_12178);
and U21674 (N_21674,N_15339,N_16124);
or U21675 (N_21675,N_18398,N_18982);
and U21676 (N_21676,N_19753,N_12850);
or U21677 (N_21677,N_11212,N_12827);
and U21678 (N_21678,N_15359,N_13637);
nand U21679 (N_21679,N_16581,N_14785);
nand U21680 (N_21680,N_13598,N_11318);
and U21681 (N_21681,N_14579,N_18950);
nor U21682 (N_21682,N_10086,N_14930);
nor U21683 (N_21683,N_17371,N_19880);
or U21684 (N_21684,N_14511,N_18390);
or U21685 (N_21685,N_15615,N_19055);
and U21686 (N_21686,N_15635,N_11865);
or U21687 (N_21687,N_17565,N_19707);
xnor U21688 (N_21688,N_12719,N_11354);
nor U21689 (N_21689,N_17420,N_11262);
nor U21690 (N_21690,N_15706,N_14770);
and U21691 (N_21691,N_15812,N_18418);
or U21692 (N_21692,N_18490,N_13011);
nor U21693 (N_21693,N_14615,N_10227);
nor U21694 (N_21694,N_18450,N_14180);
and U21695 (N_21695,N_19293,N_12572);
nor U21696 (N_21696,N_18962,N_15290);
or U21697 (N_21697,N_15871,N_13197);
or U21698 (N_21698,N_11809,N_16484);
xor U21699 (N_21699,N_13256,N_13503);
and U21700 (N_21700,N_11106,N_17968);
nor U21701 (N_21701,N_11423,N_19225);
nor U21702 (N_21702,N_16701,N_10297);
nand U21703 (N_21703,N_13745,N_18325);
and U21704 (N_21704,N_16461,N_15556);
nand U21705 (N_21705,N_11074,N_17002);
or U21706 (N_21706,N_18523,N_14048);
nor U21707 (N_21707,N_11911,N_19818);
or U21708 (N_21708,N_17601,N_11093);
and U21709 (N_21709,N_15699,N_15659);
nand U21710 (N_21710,N_13104,N_10758);
nand U21711 (N_21711,N_15554,N_16770);
and U21712 (N_21712,N_15441,N_13946);
or U21713 (N_21713,N_11748,N_19690);
nor U21714 (N_21714,N_18200,N_19375);
or U21715 (N_21715,N_14164,N_13708);
nor U21716 (N_21716,N_14259,N_12832);
nor U21717 (N_21717,N_11505,N_11486);
or U21718 (N_21718,N_13141,N_10878);
and U21719 (N_21719,N_18632,N_12710);
or U21720 (N_21720,N_16000,N_10245);
and U21721 (N_21721,N_13022,N_10834);
and U21722 (N_21722,N_19735,N_16215);
or U21723 (N_21723,N_13101,N_10088);
and U21724 (N_21724,N_19640,N_10228);
xnor U21725 (N_21725,N_16993,N_14061);
nor U21726 (N_21726,N_12091,N_13489);
and U21727 (N_21727,N_17664,N_13484);
nor U21728 (N_21728,N_10231,N_13701);
nor U21729 (N_21729,N_17529,N_19428);
or U21730 (N_21730,N_17201,N_16846);
or U21731 (N_21731,N_14427,N_14509);
and U21732 (N_21732,N_11075,N_10582);
or U21733 (N_21733,N_11030,N_19119);
or U21734 (N_21734,N_11760,N_14705);
and U21735 (N_21735,N_14371,N_14599);
or U21736 (N_21736,N_13858,N_13311);
nand U21737 (N_21737,N_18711,N_10322);
nor U21738 (N_21738,N_10846,N_12101);
and U21739 (N_21739,N_16059,N_17079);
and U21740 (N_21740,N_14204,N_17719);
or U21741 (N_21741,N_13537,N_17514);
and U21742 (N_21742,N_12048,N_15950);
or U21743 (N_21743,N_17503,N_11575);
or U21744 (N_21744,N_11230,N_10409);
or U21745 (N_21745,N_19578,N_17560);
and U21746 (N_21746,N_13032,N_18806);
nand U21747 (N_21747,N_11481,N_17761);
nor U21748 (N_21748,N_12044,N_17211);
or U21749 (N_21749,N_19799,N_13718);
nand U21750 (N_21750,N_14661,N_13771);
or U21751 (N_21751,N_19396,N_16325);
nor U21752 (N_21752,N_13175,N_19660);
nand U21753 (N_21753,N_19941,N_18718);
and U21754 (N_21754,N_12985,N_11579);
nor U21755 (N_21755,N_17721,N_14546);
or U21756 (N_21756,N_15597,N_12780);
or U21757 (N_21757,N_11110,N_10237);
nor U21758 (N_21758,N_12250,N_15363);
nand U21759 (N_21759,N_17535,N_14448);
nand U21760 (N_21760,N_17925,N_14076);
and U21761 (N_21761,N_10764,N_10847);
nand U21762 (N_21762,N_15461,N_12664);
or U21763 (N_21763,N_10173,N_18338);
and U21764 (N_21764,N_14200,N_11653);
and U21765 (N_21765,N_18963,N_10536);
and U21766 (N_21766,N_18395,N_13368);
nor U21767 (N_21767,N_18566,N_18724);
and U21768 (N_21768,N_15664,N_10223);
xor U21769 (N_21769,N_16829,N_12209);
or U21770 (N_21770,N_13943,N_18041);
nand U21771 (N_21771,N_13339,N_11820);
and U21772 (N_21772,N_13657,N_18849);
and U21773 (N_21773,N_11966,N_13024);
and U21774 (N_21774,N_19269,N_13606);
and U21775 (N_21775,N_17375,N_11360);
nand U21776 (N_21776,N_14540,N_12157);
or U21777 (N_21777,N_16987,N_16011);
nor U21778 (N_21778,N_11658,N_19627);
and U21779 (N_21779,N_17153,N_10844);
nor U21780 (N_21780,N_11874,N_10624);
nand U21781 (N_21781,N_15570,N_10178);
or U21782 (N_21782,N_14847,N_14499);
nor U21783 (N_21783,N_17036,N_11248);
nand U21784 (N_21784,N_12198,N_12411);
nand U21785 (N_21785,N_13717,N_15891);
nor U21786 (N_21786,N_11611,N_11574);
and U21787 (N_21787,N_13237,N_17863);
nor U21788 (N_21788,N_18863,N_10024);
nand U21789 (N_21789,N_11117,N_16905);
nand U21790 (N_21790,N_11276,N_12098);
or U21791 (N_21791,N_15767,N_12406);
nand U21792 (N_21792,N_17951,N_14254);
and U21793 (N_21793,N_12114,N_18903);
or U21794 (N_21794,N_10838,N_19438);
nor U21795 (N_21795,N_15240,N_12236);
nor U21796 (N_21796,N_13318,N_16773);
or U21797 (N_21797,N_17258,N_11288);
or U21798 (N_21798,N_14213,N_19482);
and U21799 (N_21799,N_16838,N_12991);
nand U21800 (N_21800,N_11532,N_11011);
nor U21801 (N_21801,N_14107,N_10770);
nand U21802 (N_21802,N_11286,N_19240);
nand U21803 (N_21803,N_15619,N_15482);
and U21804 (N_21804,N_19282,N_10869);
nor U21805 (N_21805,N_17697,N_17141);
nand U21806 (N_21806,N_12947,N_17168);
or U21807 (N_21807,N_14163,N_11491);
nand U21808 (N_21808,N_15071,N_17935);
and U21809 (N_21809,N_16004,N_18832);
nand U21810 (N_21810,N_17734,N_18098);
or U21811 (N_21811,N_12158,N_11371);
and U21812 (N_21812,N_15788,N_16936);
nor U21813 (N_21813,N_16426,N_14146);
nand U21814 (N_21814,N_14702,N_19370);
nor U21815 (N_21815,N_12387,N_18354);
and U21816 (N_21816,N_11528,N_12171);
or U21817 (N_21817,N_19623,N_17646);
or U21818 (N_21818,N_10969,N_17452);
and U21819 (N_21819,N_13420,N_12957);
nor U21820 (N_21820,N_16699,N_18252);
nor U21821 (N_21821,N_15045,N_17605);
or U21822 (N_21822,N_11659,N_16787);
and U21823 (N_21823,N_13977,N_11259);
nor U21824 (N_21824,N_13354,N_17095);
and U21825 (N_21825,N_17726,N_10444);
nand U21826 (N_21826,N_16925,N_17145);
nand U21827 (N_21827,N_11355,N_15110);
nand U21828 (N_21828,N_19357,N_10819);
nor U21829 (N_21829,N_16503,N_14033);
nor U21830 (N_21830,N_18107,N_10922);
nor U21831 (N_21831,N_16096,N_19419);
nand U21832 (N_21832,N_10583,N_13160);
nand U21833 (N_21833,N_18067,N_10881);
or U21834 (N_21834,N_18084,N_13807);
or U21835 (N_21835,N_11588,N_16924);
nor U21836 (N_21836,N_13365,N_16042);
or U21837 (N_21837,N_15362,N_19106);
or U21838 (N_21838,N_12889,N_14755);
or U21839 (N_21839,N_18760,N_17615);
and U21840 (N_21840,N_11834,N_19645);
nand U21841 (N_21841,N_15606,N_11291);
or U21842 (N_21842,N_12459,N_15525);
nor U21843 (N_21843,N_19310,N_14582);
and U21844 (N_21844,N_13508,N_16666);
nand U21845 (N_21845,N_17206,N_16257);
or U21846 (N_21846,N_14030,N_18505);
nand U21847 (N_21847,N_12545,N_11451);
nor U21848 (N_21848,N_15946,N_16676);
nand U21849 (N_21849,N_10378,N_17927);
nor U21850 (N_21850,N_16834,N_17973);
nand U21851 (N_21851,N_11350,N_16616);
and U21852 (N_21852,N_14504,N_11225);
or U21853 (N_21853,N_10653,N_13379);
nor U21854 (N_21854,N_16288,N_14273);
nor U21855 (N_21855,N_10461,N_16396);
nand U21856 (N_21856,N_10413,N_13479);
nor U21857 (N_21857,N_14569,N_16238);
nor U21858 (N_21858,N_14923,N_14763);
nor U21859 (N_21859,N_17481,N_10445);
nor U21860 (N_21860,N_10054,N_11061);
or U21861 (N_21861,N_10499,N_13212);
and U21862 (N_21862,N_13584,N_11214);
nor U21863 (N_21863,N_16156,N_16421);
nand U21864 (N_21864,N_15485,N_16760);
nand U21865 (N_21865,N_10474,N_13839);
nor U21866 (N_21866,N_19368,N_12463);
nand U21867 (N_21867,N_19652,N_15686);
nor U21868 (N_21868,N_14811,N_19961);
nand U21869 (N_21869,N_18844,N_19349);
nor U21870 (N_21870,N_12375,N_15166);
nor U21871 (N_21871,N_19073,N_10243);
nor U21872 (N_21872,N_18916,N_18897);
or U21873 (N_21873,N_16097,N_16419);
nand U21874 (N_21874,N_11772,N_17262);
nor U21875 (N_21875,N_16895,N_19807);
nor U21876 (N_21876,N_16056,N_15229);
xnor U21877 (N_21877,N_16541,N_16314);
or U21878 (N_21878,N_13190,N_11352);
and U21879 (N_21879,N_10079,N_18753);
and U21880 (N_21880,N_15048,N_18929);
and U21881 (N_21881,N_11813,N_19767);
nor U21882 (N_21882,N_15921,N_15404);
nand U21883 (N_21883,N_10128,N_12168);
and U21884 (N_21884,N_17303,N_19525);
and U21885 (N_21885,N_15091,N_17517);
or U21886 (N_21886,N_17434,N_17835);
nor U21887 (N_21887,N_16533,N_14571);
and U21888 (N_21888,N_18058,N_12723);
and U21889 (N_21889,N_15317,N_13186);
and U21890 (N_21890,N_14268,N_16771);
and U21891 (N_21891,N_17240,N_19377);
nor U21892 (N_21892,N_19908,N_17990);
and U21893 (N_21893,N_17545,N_19512);
nor U21894 (N_21894,N_17801,N_19270);
and U21895 (N_21895,N_18262,N_18662);
and U21896 (N_21896,N_12958,N_14507);
or U21897 (N_21897,N_10667,N_12749);
nor U21898 (N_21898,N_12478,N_16422);
or U21899 (N_21899,N_10036,N_12176);
or U21900 (N_21900,N_14420,N_10510);
and U21901 (N_21901,N_17814,N_10174);
nor U21902 (N_21902,N_16534,N_13264);
nor U21903 (N_21903,N_17695,N_19342);
nand U21904 (N_21904,N_16412,N_10433);
and U21905 (N_21905,N_10417,N_12940);
nor U21906 (N_21906,N_13700,N_15594);
and U21907 (N_21907,N_12711,N_15094);
nor U21908 (N_21908,N_18239,N_13213);
nand U21909 (N_21909,N_10176,N_11362);
nor U21910 (N_21910,N_11210,N_17401);
or U21911 (N_21911,N_13698,N_17838);
and U21912 (N_21912,N_12677,N_12840);
and U21913 (N_21913,N_17286,N_11722);
nand U21914 (N_21914,N_19415,N_17526);
or U21915 (N_21915,N_10626,N_17399);
nor U21916 (N_21916,N_17284,N_13814);
nor U21917 (N_21917,N_16732,N_19622);
nand U21918 (N_21918,N_15739,N_14591);
nor U21919 (N_21919,N_18893,N_12452);
and U21920 (N_21920,N_19229,N_13825);
and U21921 (N_21921,N_12027,N_10841);
or U21922 (N_21922,N_12473,N_18569);
nor U21923 (N_21923,N_10383,N_17700);
and U21924 (N_21924,N_11237,N_15155);
nand U21925 (N_21925,N_16219,N_10367);
nand U21926 (N_21926,N_10757,N_19940);
nand U21927 (N_21927,N_17654,N_15310);
or U21928 (N_21928,N_10515,N_18649);
nor U21929 (N_21929,N_12446,N_17292);
nand U21930 (N_21930,N_18368,N_18818);
nor U21931 (N_21931,N_17729,N_16161);
and U21932 (N_21932,N_10570,N_15196);
or U21933 (N_21933,N_18796,N_14357);
nand U21934 (N_21934,N_19259,N_17035);
nand U21935 (N_21935,N_17026,N_18644);
or U21936 (N_21936,N_17659,N_16596);
nand U21937 (N_21937,N_17265,N_12552);
and U21938 (N_21938,N_17844,N_12404);
nand U21939 (N_21939,N_13835,N_19529);
and U21940 (N_21940,N_16081,N_14594);
nor U21941 (N_21941,N_12342,N_16624);
nand U21942 (N_21942,N_14883,N_16251);
and U21943 (N_21943,N_14003,N_14769);
nand U21944 (N_21944,N_19875,N_15169);
nor U21945 (N_21945,N_12116,N_18549);
and U21946 (N_21946,N_14962,N_15118);
nand U21947 (N_21947,N_19999,N_18822);
nor U21948 (N_21948,N_10808,N_13553);
and U21949 (N_21949,N_14927,N_10887);
nand U21950 (N_21950,N_10603,N_14023);
nand U21951 (N_21951,N_18918,N_17186);
and U21952 (N_21952,N_10400,N_19944);
or U21953 (N_21953,N_11766,N_16189);
and U21954 (N_21954,N_15152,N_11418);
or U21955 (N_21955,N_15200,N_12856);
nand U21956 (N_21956,N_15915,N_15012);
nand U21957 (N_21957,N_17680,N_17191);
or U21958 (N_21958,N_14024,N_17431);
nand U21959 (N_21959,N_19418,N_10194);
nand U21960 (N_21960,N_17699,N_11687);
nor U21961 (N_21961,N_17367,N_15397);
nand U21962 (N_21962,N_13515,N_10980);
and U21963 (N_21963,N_10188,N_14812);
nor U21964 (N_21964,N_18247,N_14478);
or U21965 (N_21965,N_18164,N_16857);
nor U21966 (N_21966,N_12150,N_16740);
and U21967 (N_21967,N_17833,N_12849);
nand U21968 (N_21968,N_14059,N_11645);
and U21969 (N_21969,N_18808,N_18198);
nand U21970 (N_21970,N_12360,N_17539);
nand U21971 (N_21971,N_11682,N_12589);
and U21972 (N_21972,N_15823,N_12633);
and U21973 (N_21973,N_19321,N_15413);
and U21974 (N_21974,N_18985,N_18142);
nor U21975 (N_21975,N_12689,N_17409);
or U21976 (N_21976,N_15254,N_15038);
nand U21977 (N_21977,N_10111,N_19574);
or U21978 (N_21978,N_12524,N_13891);
or U21979 (N_21979,N_13833,N_18056);
or U21980 (N_21980,N_11340,N_14585);
or U21981 (N_21981,N_14127,N_16990);
nor U21982 (N_21982,N_14166,N_11475);
nand U21983 (N_21983,N_15188,N_10935);
nor U21984 (N_21984,N_12185,N_12103);
and U21985 (N_21985,N_19987,N_12383);
or U21986 (N_21986,N_10562,N_12443);
or U21987 (N_21987,N_18623,N_16962);
nor U21988 (N_21988,N_11804,N_12568);
nor U21989 (N_21989,N_14009,N_13520);
or U21990 (N_21990,N_13042,N_16253);
or U21991 (N_21991,N_10496,N_18385);
and U21992 (N_21992,N_10216,N_18099);
or U21993 (N_21993,N_15687,N_13084);
nor U21994 (N_21994,N_14969,N_15149);
and U21995 (N_21995,N_10596,N_13466);
nand U21996 (N_21996,N_10058,N_12926);
nor U21997 (N_21997,N_12369,N_16970);
nand U21998 (N_21998,N_16800,N_18592);
or U21999 (N_21999,N_19479,N_18544);
or U22000 (N_22000,N_14249,N_17023);
nor U22001 (N_22001,N_15895,N_16437);
nand U22002 (N_22002,N_16468,N_14157);
and U22003 (N_22003,N_11477,N_15251);
or U22004 (N_22004,N_18498,N_19146);
nand U22005 (N_22005,N_13514,N_13306);
nand U22006 (N_22006,N_15701,N_16945);
nand U22007 (N_22007,N_16439,N_19226);
nor U22008 (N_22008,N_12120,N_10021);
or U22009 (N_22009,N_13603,N_14774);
nor U22010 (N_22010,N_10555,N_18934);
and U22011 (N_22011,N_16187,N_12128);
nor U22012 (N_22012,N_15582,N_11013);
nor U22013 (N_22013,N_18036,N_11704);
and U22014 (N_22014,N_15327,N_10964);
and U22015 (N_22015,N_13619,N_11089);
and U22016 (N_22016,N_16111,N_12667);
nand U22017 (N_22017,N_17505,N_11851);
nand U22018 (N_22018,N_19541,N_13957);
or U22019 (N_22019,N_11750,N_13352);
and U22020 (N_22020,N_17753,N_10170);
or U22021 (N_22021,N_18052,N_11000);
nor U22022 (N_22022,N_13188,N_16750);
and U22023 (N_22023,N_15749,N_18135);
and U22024 (N_22024,N_19881,N_12675);
or U22025 (N_22025,N_11498,N_14689);
and U22026 (N_22026,N_19075,N_11324);
or U22027 (N_22027,N_12698,N_10784);
nand U22028 (N_22028,N_12978,N_15926);
or U22029 (N_22029,N_10234,N_18744);
and U22030 (N_22030,N_17751,N_18771);
or U22031 (N_22031,N_18917,N_10673);
or U22032 (N_22032,N_17313,N_11589);
nor U22033 (N_22033,N_19768,N_14472);
or U22034 (N_22034,N_15846,N_14177);
or U22035 (N_22035,N_13562,N_19267);
or U22036 (N_22036,N_14663,N_18116);
or U22037 (N_22037,N_15835,N_11852);
nor U22038 (N_22038,N_11096,N_17361);
and U22039 (N_22039,N_18854,N_18743);
and U22040 (N_22040,N_15369,N_14253);
or U22041 (N_22041,N_11917,N_13161);
nor U22042 (N_22042,N_10872,N_14616);
nor U22043 (N_22043,N_10717,N_13070);
nand U22044 (N_22044,N_12234,N_14333);
and U22045 (N_22045,N_15563,N_11091);
nor U22046 (N_22046,N_13286,N_16877);
nor U22047 (N_22047,N_17344,N_18557);
and U22048 (N_22048,N_16127,N_15929);
nand U22049 (N_22049,N_11310,N_10754);
and U22050 (N_22050,N_13559,N_19397);
nand U22051 (N_22051,N_15679,N_15032);
nand U22052 (N_22052,N_18279,N_12652);
and U22053 (N_22053,N_16663,N_15066);
or U22054 (N_22054,N_12578,N_17903);
and U22055 (N_22055,N_14828,N_19784);
nand U22056 (N_22056,N_11432,N_13837);
or U22057 (N_22057,N_13841,N_12196);
nor U22058 (N_22058,N_14294,N_14130);
nor U22059 (N_22059,N_12760,N_12992);
or U22060 (N_22060,N_12372,N_17410);
nand U22061 (N_22061,N_19800,N_16018);
nor U22062 (N_22062,N_12694,N_11965);
nand U22063 (N_22063,N_15967,N_10317);
or U22064 (N_22064,N_16684,N_16599);
and U22065 (N_22065,N_11745,N_12834);
and U22066 (N_22066,N_16236,N_17331);
nand U22067 (N_22067,N_11594,N_12506);
and U22068 (N_22068,N_13709,N_14301);
nand U22069 (N_22069,N_10179,N_10286);
or U22070 (N_22070,N_15667,N_12757);
nor U22071 (N_22071,N_14867,N_17172);
and U22072 (N_22072,N_12755,N_10491);
nor U22073 (N_22073,N_18452,N_17588);
or U22074 (N_22074,N_11578,N_15236);
and U22075 (N_22075,N_13429,N_17923);
nand U22076 (N_22076,N_13975,N_18720);
nand U22077 (N_22077,N_17345,N_14646);
or U22078 (N_22078,N_19584,N_15454);
nor U22079 (N_22079,N_16213,N_16577);
nand U22080 (N_22080,N_14300,N_17436);
and U22081 (N_22081,N_19488,N_19567);
nor U22082 (N_22082,N_15009,N_14022);
or U22083 (N_22083,N_12650,N_11904);
nor U22084 (N_22084,N_15123,N_13557);
and U22085 (N_22085,N_19371,N_18944);
or U22086 (N_22086,N_14991,N_15389);
and U22087 (N_22087,N_15753,N_15464);
nand U22088 (N_22088,N_13326,N_15266);
nor U22089 (N_22089,N_17487,N_10785);
and U22090 (N_22090,N_16523,N_14422);
or U22091 (N_22091,N_13159,N_17957);
and U22092 (N_22092,N_13421,N_12728);
nor U22093 (N_22093,N_12075,N_12536);
nor U22094 (N_22094,N_15361,N_19401);
nand U22095 (N_22095,N_11226,N_14231);
and U22096 (N_22096,N_15689,N_13813);
or U22097 (N_22097,N_16863,N_15401);
nor U22098 (N_22098,N_11546,N_10790);
or U22099 (N_22099,N_19077,N_16060);
and U22100 (N_22100,N_11485,N_14058);
nor U22101 (N_22101,N_10534,N_10117);
or U22102 (N_22102,N_14798,N_19144);
nor U22103 (N_22103,N_12283,N_11833);
nor U22104 (N_22104,N_12790,N_19001);
nand U22105 (N_22105,N_16192,N_19237);
nor U22106 (N_22106,N_11403,N_17123);
or U22107 (N_22107,N_17971,N_13404);
and U22108 (N_22108,N_14028,N_15079);
nand U22109 (N_22109,N_11786,N_17087);
nand U22110 (N_22110,N_12662,N_14412);
and U22111 (N_22111,N_11458,N_18791);
or U22112 (N_22112,N_11821,N_19618);
and U22113 (N_22113,N_10222,N_19196);
and U22114 (N_22114,N_16584,N_19508);
or U22115 (N_22115,N_14953,N_11233);
or U22116 (N_22116,N_13577,N_12933);
and U22117 (N_22117,N_12959,N_11201);
or U22118 (N_22118,N_18113,N_11361);
nand U22119 (N_22119,N_19028,N_17451);
nand U22120 (N_22120,N_11195,N_12841);
nor U22121 (N_22121,N_19183,N_14326);
nor U22122 (N_22122,N_14966,N_16826);
and U22123 (N_22123,N_12237,N_19684);
nand U22124 (N_22124,N_13279,N_12591);
nor U22125 (N_22125,N_19090,N_15376);
or U22126 (N_22126,N_12541,N_18955);
nor U22127 (N_22127,N_12823,N_19117);
nor U22128 (N_22128,N_13320,N_18734);
and U22129 (N_22129,N_15652,N_11025);
nand U22130 (N_22130,N_14746,N_15851);
or U22131 (N_22131,N_13155,N_15052);
or U22132 (N_22132,N_14738,N_13506);
or U22133 (N_22133,N_14435,N_11893);
nor U22134 (N_22134,N_14878,N_17298);
nor U22135 (N_22135,N_13903,N_18163);
or U22136 (N_22136,N_19136,N_11489);
nand U22137 (N_22137,N_17868,N_15630);
nor U22138 (N_22138,N_17466,N_14185);
and U22139 (N_22139,N_14280,N_17743);
and U22140 (N_22140,N_19535,N_12786);
nor U22141 (N_22141,N_17459,N_19720);
nor U22142 (N_22142,N_19785,N_12287);
nor U22143 (N_22143,N_12909,N_11534);
or U22144 (N_22144,N_10814,N_16102);
or U22145 (N_22145,N_12186,N_17897);
or U22146 (N_22146,N_19234,N_19485);
nor U22147 (N_22147,N_15992,N_10557);
and U22148 (N_22148,N_15585,N_19105);
and U22149 (N_22149,N_10356,N_12225);
nor U22150 (N_22150,N_17834,N_11264);
and U22151 (N_22151,N_18869,N_12982);
and U22152 (N_22152,N_18030,N_15358);
nor U22153 (N_22153,N_13624,N_16593);
nor U22154 (N_22154,N_14461,N_14786);
or U22155 (N_22155,N_19585,N_15840);
or U22156 (N_22156,N_16817,N_11297);
nand U22157 (N_22157,N_14045,N_14612);
nand U22158 (N_22158,N_14462,N_17617);
or U22159 (N_22159,N_18964,N_13000);
and U22160 (N_22160,N_12298,N_16521);
or U22161 (N_22161,N_11584,N_19769);
and U22162 (N_22162,N_11029,N_13580);
nor U22163 (N_22163,N_18872,N_12118);
nand U22164 (N_22164,N_11413,N_12010);
nand U22165 (N_22165,N_14145,N_19411);
or U22166 (N_22166,N_10230,N_12733);
nor U22167 (N_22167,N_11867,N_11920);
and U22168 (N_22168,N_15661,N_13889);
or U22169 (N_22169,N_10687,N_16540);
nor U22170 (N_22170,N_15516,N_18996);
or U22171 (N_22171,N_17929,N_15596);
or U22172 (N_22172,N_11635,N_11442);
and U22173 (N_22173,N_12337,N_16731);
and U22174 (N_22174,N_19095,N_19445);
nor U22175 (N_22175,N_12026,N_19286);
or U22176 (N_22176,N_16185,N_10266);
nand U22177 (N_22177,N_11446,N_17733);
nand U22178 (N_22178,N_13014,N_15579);
nand U22179 (N_22179,N_12600,N_17448);
and U22180 (N_22180,N_18109,N_13638);
and U22181 (N_22181,N_18375,N_12276);
and U22182 (N_22182,N_17592,N_19093);
and U22183 (N_22183,N_17985,N_15137);
nand U22184 (N_22184,N_16958,N_19516);
nor U22185 (N_22185,N_16202,N_19309);
and U22186 (N_22186,N_19276,N_16844);
nand U22187 (N_22187,N_19809,N_13804);
or U22188 (N_22188,N_17880,N_17482);
nand U22189 (N_22189,N_10759,N_10279);
nor U22190 (N_22190,N_13690,N_12467);
nor U22191 (N_22191,N_12981,N_14960);
or U22192 (N_22192,N_10694,N_18983);
and U22193 (N_22193,N_11891,N_13363);
or U22194 (N_22194,N_12374,N_19930);
and U22195 (N_22195,N_13283,N_16460);
nand U22196 (N_22196,N_15663,N_19977);
or U22197 (N_22197,N_14203,N_18956);
or U22198 (N_22198,N_14347,N_19924);
xor U22199 (N_22199,N_15515,N_15505);
nand U22200 (N_22200,N_12500,N_11427);
nor U22201 (N_22201,N_17756,N_14990);
or U22202 (N_22202,N_18156,N_10702);
nand U22203 (N_22203,N_11755,N_13601);
nor U22204 (N_22204,N_10395,N_19540);
or U22205 (N_22205,N_11800,N_11975);
xor U22206 (N_22206,N_13220,N_11254);
and U22207 (N_22207,N_15947,N_16653);
and U22208 (N_22208,N_17478,N_19581);
nor U22209 (N_22209,N_19180,N_11907);
and U22210 (N_22210,N_16431,N_17916);
and U22211 (N_22211,N_18630,N_11187);
nand U22212 (N_22212,N_11525,N_12035);
nor U22213 (N_22213,N_11283,N_10427);
or U22214 (N_22214,N_13822,N_11068);
or U22215 (N_22215,N_10331,N_11695);
nor U22216 (N_22216,N_19855,N_18080);
and U22217 (N_22217,N_11533,N_18992);
and U22218 (N_22218,N_15969,N_17803);
nor U22219 (N_22219,N_10521,N_10715);
and U22220 (N_22220,N_16522,N_18240);
and U22221 (N_22221,N_16277,N_14067);
and U22222 (N_22222,N_12320,N_11241);
nor U22223 (N_22223,N_18699,N_16969);
nand U22224 (N_22224,N_19065,N_10337);
nor U22225 (N_22225,N_11831,N_19988);
and U22226 (N_22226,N_12960,N_18001);
nor U22227 (N_22227,N_17174,N_16885);
or U22228 (N_22228,N_18828,N_15913);
nor U22229 (N_22229,N_10938,N_13556);
and U22230 (N_22230,N_13616,N_14010);
nand U22231 (N_22231,N_10414,N_14978);
and U22232 (N_22232,N_13973,N_19628);
and U22233 (N_22233,N_17349,N_14766);
and U22234 (N_22234,N_18587,N_18717);
nand U22235 (N_22235,N_17837,N_18213);
nand U22236 (N_22236,N_14737,N_18007);
nand U22237 (N_22237,N_13369,N_13362);
nand U22238 (N_22238,N_17285,N_19990);
nand U22239 (N_22239,N_13272,N_19594);
nand U22240 (N_22240,N_12497,N_13754);
and U22241 (N_22241,N_12961,N_10271);
nor U22242 (N_22242,N_10084,N_15616);
or U22243 (N_22243,N_18702,N_18359);
and U22244 (N_22244,N_15725,N_12811);
and U22245 (N_22245,N_14449,N_10207);
nor U22246 (N_22246,N_12882,N_18594);
nand U22247 (N_22247,N_11876,N_13013);
or U22248 (N_22248,N_14609,N_14973);
nor U22249 (N_22249,N_15356,N_19343);
or U22250 (N_22250,N_15353,N_13360);
nor U22251 (N_22251,N_15436,N_14383);
or U22252 (N_22252,N_16285,N_14335);
nor U22253 (N_22253,N_10813,N_15262);
or U22254 (N_22254,N_14112,N_15500);
and U22255 (N_22255,N_18633,N_17613);
or U22256 (N_22256,N_11858,N_15838);
or U22257 (N_22257,N_16183,N_17857);
nor U22258 (N_22258,N_18410,N_10249);
nand U22259 (N_22259,N_19273,N_17169);
nand U22260 (N_22260,N_12460,N_10945);
nor U22261 (N_22261,N_10363,N_12939);
and U22262 (N_22262,N_14800,N_10915);
and U22263 (N_22263,N_16644,N_16165);
nand U22264 (N_22264,N_14218,N_17219);
nor U22265 (N_22265,N_18994,N_19680);
nor U22266 (N_22266,N_16246,N_16023);
or U22267 (N_22267,N_10586,N_15986);
nand U22268 (N_22268,N_10483,N_11900);
and U22269 (N_22269,N_19158,N_14078);
or U22270 (N_22270,N_13614,N_14396);
nand U22271 (N_22271,N_12632,N_10391);
nand U22272 (N_22272,N_18184,N_19323);
nand U22273 (N_22273,N_11668,N_18932);
or U22274 (N_22274,N_19336,N_17954);
and U22275 (N_22275,N_12038,N_15022);
or U22276 (N_22276,N_11272,N_17370);
or U22277 (N_22277,N_18968,N_10866);
or U22278 (N_22278,N_16338,N_18755);
nand U22279 (N_22279,N_10675,N_12898);
nor U22280 (N_22280,N_17216,N_14868);
nand U22281 (N_22281,N_13773,N_12599);
and U22282 (N_22282,N_19029,N_19731);
nor U22283 (N_22283,N_14744,N_18320);
and U22284 (N_22284,N_11166,N_10081);
nand U22285 (N_22285,N_11875,N_14375);
nor U22286 (N_22286,N_10795,N_11058);
nand U22287 (N_22287,N_15550,N_14128);
and U22288 (N_22288,N_19446,N_12051);
or U22289 (N_22289,N_19319,N_11149);
or U22290 (N_22290,N_18426,N_16057);
and U22291 (N_22291,N_19002,N_18340);
xor U22292 (N_22292,N_15660,N_17643);
nor U22293 (N_22293,N_18020,N_14742);
nor U22294 (N_22294,N_15748,N_18641);
nand U22295 (N_22295,N_19199,N_11951);
and U22296 (N_22296,N_16613,N_15638);
or U22297 (N_22297,N_11873,N_17718);
nor U22298 (N_22298,N_13195,N_11479);
nor U22299 (N_22299,N_19134,N_16239);
nand U22300 (N_22300,N_14831,N_16211);
and U22301 (N_22301,N_14088,N_13410);
or U22302 (N_22302,N_10165,N_19547);
xnor U22303 (N_22303,N_11482,N_11050);
and U22304 (N_22304,N_16816,N_18140);
and U22305 (N_22305,N_19284,N_11406);
nor U22306 (N_22306,N_13648,N_11661);
and U22307 (N_22307,N_18277,N_16919);
and U22308 (N_22308,N_10585,N_18467);
nand U22309 (N_22309,N_17282,N_12627);
or U22310 (N_22310,N_18516,N_12726);
or U22311 (N_22311,N_15587,N_14963);
nand U22312 (N_22312,N_15854,N_14196);
nand U22313 (N_22313,N_12437,N_14501);
nor U22314 (N_22314,N_12701,N_10615);
nor U22315 (N_22315,N_16093,N_12410);
and U22316 (N_22316,N_15861,N_14649);
or U22317 (N_22317,N_18188,N_14825);
nand U22318 (N_22318,N_18434,N_15245);
or U22319 (N_22319,N_19700,N_14139);
and U22320 (N_22320,N_16785,N_16788);
or U22321 (N_22321,N_14469,N_10738);
nand U22322 (N_22322,N_19603,N_14108);
nor U22323 (N_22323,N_11953,N_14282);
nor U22324 (N_22324,N_17050,N_18856);
and U22325 (N_22325,N_15395,N_12136);
nor U22326 (N_22326,N_10046,N_10494);
or U22327 (N_22327,N_14931,N_19047);
or U22328 (N_22328,N_16233,N_17507);
or U22329 (N_22329,N_15025,N_16240);
nor U22330 (N_22330,N_11784,N_13548);
and U22331 (N_22331,N_11646,N_14265);
or U22332 (N_22332,N_10290,N_15908);
or U22333 (N_22333,N_19091,N_11693);
or U22334 (N_22334,N_11379,N_14843);
or U22335 (N_22335,N_16654,N_19213);
and U22336 (N_22336,N_14414,N_19027);
nor U22337 (N_22337,N_12160,N_11812);
and U22338 (N_22338,N_12143,N_16142);
or U22339 (N_22339,N_12720,N_15298);
nor U22340 (N_22340,N_16755,N_18055);
or U22341 (N_22341,N_13037,N_12735);
and U22342 (N_22342,N_16312,N_14556);
nand U22343 (N_22343,N_19558,N_12671);
and U22344 (N_22344,N_12254,N_15307);
or U22345 (N_22345,N_12341,N_12742);
or U22346 (N_22346,N_19523,N_19702);
nor U22347 (N_22347,N_18150,N_15399);
nand U22348 (N_22348,N_19330,N_14389);
or U22349 (N_22349,N_18958,N_15822);
and U22350 (N_22350,N_13249,N_11621);
nor U22351 (N_22351,N_15795,N_13232);
and U22352 (N_22352,N_19819,N_19246);
and U22353 (N_22353,N_19873,N_18705);
or U22354 (N_22354,N_19015,N_19936);
and U22355 (N_22355,N_10403,N_16961);
nand U22356 (N_22356,N_17749,N_18895);
nor U22357 (N_22357,N_13043,N_15321);
or U22358 (N_22358,N_18841,N_16859);
xor U22359 (N_22359,N_18287,N_15676);
nor U22360 (N_22360,N_15302,N_16781);
nor U22361 (N_22361,N_19786,N_16938);
nand U22362 (N_22362,N_12974,N_10287);
and U22363 (N_22363,N_13010,N_10126);
nand U22364 (N_22364,N_10597,N_18710);
nor U22365 (N_22365,N_18563,N_12966);
and U22366 (N_22366,N_17611,N_16282);
xor U22367 (N_22367,N_19945,N_18525);
or U22368 (N_22368,N_12614,N_12243);
and U22369 (N_22369,N_12310,N_11719);
or U22370 (N_22370,N_15566,N_12605);
and U22371 (N_22371,N_11742,N_13697);
and U22372 (N_22372,N_18746,N_16893);
or U22373 (N_22373,N_16207,N_12309);
and U22374 (N_22374,N_14075,N_10233);
nor U22375 (N_22375,N_13569,N_14698);
nor U22376 (N_22376,N_16807,N_11903);
nor U22377 (N_22377,N_19302,N_15509);
nor U22378 (N_22378,N_13856,N_11023);
or U22379 (N_22379,N_17276,N_13261);
or U22380 (N_22380,N_12646,N_11109);
nand U22381 (N_22381,N_11334,N_17074);
or U22382 (N_22382,N_18788,N_16317);
nor U22383 (N_22383,N_10344,N_19892);
nand U22384 (N_22384,N_18574,N_16416);
or U22385 (N_22385,N_12265,N_12996);
or U22386 (N_22386,N_11597,N_13490);
nand U22387 (N_22387,N_17200,N_15037);
nand U22388 (N_22388,N_13380,N_17882);
nand U22389 (N_22389,N_19004,N_19165);
and U22390 (N_22390,N_15532,N_18322);
nor U22391 (N_22391,N_10392,N_11349);
nor U22392 (N_22392,N_15698,N_19030);
or U22393 (N_22393,N_16505,N_15476);
or U22394 (N_22394,N_10939,N_18008);
and U22395 (N_22395,N_17825,N_15131);
and U22396 (N_22396,N_13067,N_19608);
nor U22397 (N_22397,N_12725,N_13761);
nand U22398 (N_22398,N_15332,N_12621);
and U22399 (N_22399,N_18212,N_16860);
or U22400 (N_22400,N_19863,N_14862);
nand U22401 (N_22401,N_11956,N_19187);
nor U22402 (N_22402,N_15092,N_13646);
nor U22403 (N_22403,N_14531,N_14749);
nor U22404 (N_22404,N_11328,N_17232);
nand U22405 (N_22405,N_18959,N_14992);
and U22406 (N_22406,N_10778,N_18880);
or U22407 (N_22407,N_17782,N_16999);
and U22408 (N_22408,N_16833,N_16672);
nand U22409 (N_22409,N_15018,N_12562);
nand U22410 (N_22410,N_12744,N_14974);
or U22411 (N_22411,N_11937,N_13171);
or U22412 (N_22412,N_19975,N_19932);
nor U22413 (N_22413,N_13604,N_12750);
and U22414 (N_22414,N_12564,N_17321);
nand U22415 (N_22415,N_14911,N_11968);
or U22416 (N_22416,N_16551,N_14761);
nand U22417 (N_22417,N_16712,N_10902);
nor U22418 (N_22418,N_15517,N_16931);
and U22419 (N_22419,N_10120,N_12976);
and U22420 (N_22420,N_19380,N_16851);
and U22421 (N_22421,N_19258,N_15512);
or U22422 (N_22422,N_16478,N_15683);
nand U22423 (N_22423,N_12680,N_16235);
nand U22424 (N_22424,N_17386,N_16524);
or U22425 (N_22425,N_19141,N_14198);
and U22426 (N_22426,N_12668,N_11399);
or U22427 (N_22427,N_17446,N_13053);
nor U22428 (N_22428,N_17625,N_17108);
nand U22429 (N_22429,N_13023,N_10166);
or U22430 (N_22430,N_14258,N_12874);
nor U22431 (N_22431,N_15809,N_13739);
nor U22432 (N_22432,N_15228,N_14985);
nor U22433 (N_22433,N_13435,N_11996);
or U22434 (N_22434,N_11814,N_17846);
nand U22435 (N_22435,N_19942,N_10434);
nor U22436 (N_22436,N_17121,N_18957);
nand U22437 (N_22437,N_16609,N_13527);
or U22438 (N_22438,N_19447,N_10554);
nor U22439 (N_22439,N_13334,N_16490);
and U22440 (N_22440,N_12239,N_16359);
and U22441 (N_22441,N_18203,N_17213);
nand U22442 (N_22442,N_15125,N_16710);
and U22443 (N_22443,N_18907,N_16618);
or U22444 (N_22444,N_12093,N_12223);
or U22445 (N_22445,N_19345,N_13137);
nand U22446 (N_22446,N_17789,N_15494);
nor U22447 (N_22447,N_11003,N_17577);
or U22448 (N_22448,N_14397,N_13336);
or U22449 (N_22449,N_10701,N_12880);
nor U22450 (N_22450,N_13664,N_11261);
nand U22451 (N_22451,N_18257,N_13585);
or U22452 (N_22452,N_11652,N_13704);
or U22453 (N_22453,N_10540,N_12683);
and U22454 (N_22454,N_19897,N_19207);
nand U22455 (N_22455,N_14928,N_13670);
nor U22456 (N_22456,N_18100,N_13333);
nor U22457 (N_22457,N_18842,N_11121);
nand U22458 (N_22458,N_16861,N_13218);
nand U22459 (N_22459,N_18169,N_17949);
and U22460 (N_22460,N_14101,N_17557);
and U22461 (N_22461,N_19352,N_13714);
and U22462 (N_22462,N_13179,N_12941);
nor U22463 (N_22463,N_10786,N_11776);
nor U22464 (N_22464,N_13156,N_11974);
or U22465 (N_22465,N_18470,N_11062);
nand U22466 (N_22466,N_12348,N_16025);
nor U22467 (N_22467,N_14069,N_11353);
nand U22468 (N_22468,N_15855,N_15019);
nand U22469 (N_22469,N_14584,N_14884);
nor U22470 (N_22470,N_16451,N_19444);
nor U22471 (N_22471,N_16041,N_18289);
and U22472 (N_22472,N_11705,N_17528);
and U22473 (N_22473,N_13662,N_14099);
nor U22474 (N_22474,N_17600,N_13834);
nand U22475 (N_22475,N_11751,N_13617);
nor U22476 (N_22476,N_10010,N_14384);
or U22477 (N_22477,N_14514,N_13654);
or U22478 (N_22478,N_13924,N_13998);
nor U22479 (N_22479,N_10528,N_19220);
and U22480 (N_22480,N_17273,N_12702);
nand U22481 (N_22481,N_13054,N_12579);
and U22482 (N_22482,N_13586,N_14658);
nor U22483 (N_22483,N_14913,N_19766);
nand U22484 (N_22484,N_17368,N_10642);
and U22485 (N_22485,N_18899,N_13719);
and U22486 (N_22486,N_16803,N_13274);
nand U22487 (N_22487,N_14668,N_14815);
nand U22488 (N_22488,N_18367,N_14877);
nor U22489 (N_22489,N_16225,N_12529);
nor U22490 (N_22490,N_15757,N_19387);
or U22491 (N_22491,N_18138,N_14052);
nand U22492 (N_22492,N_12042,N_17978);
nand U22493 (N_22493,N_10793,N_11912);
and U22494 (N_22494,N_16274,N_12356);
and U22495 (N_22495,N_17218,N_10429);
or U22496 (N_22496,N_15322,N_11500);
or U22497 (N_22497,N_10791,N_18343);
nand U22498 (N_22498,N_19457,N_12855);
nand U22499 (N_22499,N_15351,N_17669);
nor U22500 (N_22500,N_11861,N_13290);
and U22501 (N_22501,N_19890,N_19109);
nor U22502 (N_22502,N_13549,N_18539);
nand U22503 (N_22503,N_16276,N_10364);
nor U22504 (N_22504,N_18349,N_13182);
nor U22505 (N_22505,N_18309,N_16209);
or U22506 (N_22506,N_15477,N_18264);
nor U22507 (N_22507,N_10573,N_19788);
or U22508 (N_22508,N_17428,N_11954);
nor U22509 (N_22509,N_16843,N_15078);
nand U22510 (N_22510,N_18232,N_19507);
and U22511 (N_22511,N_15834,N_11836);
or U22512 (N_22512,N_13567,N_17948);
nor U22513 (N_22513,N_16220,N_19789);
nor U22514 (N_22514,N_11057,N_13057);
nand U22515 (N_22515,N_16167,N_12679);
or U22516 (N_22516,N_11779,N_17681);
or U22517 (N_22517,N_17822,N_14109);
nand U22518 (N_22518,N_17934,N_17194);
nor U22519 (N_22519,N_12398,N_14679);
nor U22520 (N_22520,N_19972,N_10456);
and U22521 (N_22521,N_18360,N_19737);
nor U22522 (N_22522,N_13123,N_15235);
nand U22523 (N_22523,N_14717,N_12847);
nand U22524 (N_22524,N_16724,N_15102);
nand U22525 (N_22525,N_10145,N_13925);
and U22526 (N_22526,N_13273,N_10721);
or U22527 (N_22527,N_19913,N_13587);
and U22528 (N_22528,N_15954,N_17501);
and U22529 (N_22529,N_18170,N_19639);
and U22530 (N_22530,N_19429,N_12502);
or U22531 (N_22531,N_13001,N_17046);
or U22532 (N_22532,N_11067,N_19399);
or U22533 (N_22533,N_10676,N_10779);
nor U22534 (N_22534,N_11170,N_17403);
nand U22535 (N_22535,N_19620,N_11332);
or U22536 (N_22536,N_14560,N_12718);
and U22537 (N_22537,N_10099,N_14975);
nand U22538 (N_22538,N_16328,N_13291);
nand U22539 (N_22539,N_10885,N_11545);
and U22540 (N_22540,N_12397,N_19086);
and U22541 (N_22541,N_11083,N_12073);
nand U22542 (N_22542,N_15849,N_15274);
nand U22543 (N_22543,N_18601,N_15978);
nor U22544 (N_22544,N_13936,N_15448);
nor U22545 (N_22545,N_11381,N_12704);
or U22546 (N_22546,N_18521,N_14793);
nor U22547 (N_22547,N_15273,N_10063);
nor U22548 (N_22548,N_14438,N_13255);
and U22549 (N_22549,N_12526,N_13031);
or U22550 (N_22550,N_13978,N_19576);
nand U22551 (N_22551,N_19817,N_14167);
nor U22552 (N_22552,N_12030,N_13058);
or U22553 (N_22553,N_12113,N_12753);
nor U22554 (N_22554,N_18794,N_10268);
and U22555 (N_22555,N_14561,N_19779);
nand U22556 (N_22556,N_11654,N_14401);
nor U22557 (N_22557,N_13345,N_18292);
and U22558 (N_22558,N_18123,N_17568);
nand U22559 (N_22559,N_14374,N_14025);
nand U22560 (N_22560,N_17690,N_19058);
nor U22561 (N_22561,N_12521,N_18442);
and U22562 (N_22562,N_13114,N_16454);
and U22563 (N_22563,N_18588,N_13538);
or U22564 (N_22564,N_18158,N_19295);
nand U22565 (N_22565,N_14858,N_10443);
and U22566 (N_22566,N_11778,N_19764);
or U22567 (N_22567,N_17157,N_15151);
or U22568 (N_22568,N_17854,N_16615);
and U22569 (N_22569,N_16583,N_10923);
and U22570 (N_22570,N_14629,N_15146);
nand U22571 (N_22571,N_18189,N_10127);
nand U22572 (N_22572,N_17687,N_11078);
and U22573 (N_22573,N_18736,N_17512);
nor U22574 (N_22574,N_12261,N_15718);
or U22575 (N_22575,N_14756,N_13652);
or U22576 (N_22576,N_17596,N_14937);
nand U22577 (N_22577,N_13809,N_13602);
nor U22578 (N_22578,N_13300,N_10916);
and U22579 (N_22579,N_19894,N_19322);
or U22580 (N_22580,N_19948,N_15451);
and U22581 (N_22581,N_15640,N_10327);
and U22582 (N_22582,N_16504,N_18481);
or U22583 (N_22583,N_18267,N_17038);
nor U22584 (N_22584,N_12202,N_12928);
nand U22585 (N_22585,N_13445,N_11848);
or U22586 (N_22586,N_13228,N_15029);
nor U22587 (N_22587,N_13711,N_16638);
nand U22588 (N_22588,N_18865,N_10537);
and U22589 (N_22589,N_18656,N_14121);
and U22590 (N_22590,N_12433,N_10183);
and U22591 (N_22591,N_16600,N_16456);
nand U22592 (N_22592,N_18859,N_18448);
and U22593 (N_22593,N_14580,N_15460);
or U22594 (N_22594,N_16698,N_12100);
and U22595 (N_22595,N_18571,N_15600);
nand U22596 (N_22596,N_13823,N_10730);
or U22597 (N_22597,N_11741,N_10957);
or U22598 (N_22598,N_14047,N_17723);
nor U22599 (N_22599,N_11207,N_15740);
nand U22600 (N_22600,N_11409,N_16245);
nor U22601 (N_22601,N_12831,N_14350);
nor U22602 (N_22602,N_11986,N_17813);
nor U22603 (N_22603,N_17819,N_18999);
and U22604 (N_22604,N_10753,N_12937);
or U22605 (N_22605,N_19495,N_13920);
or U22606 (N_22606,N_19554,N_12131);
nand U22607 (N_22607,N_15885,N_14497);
nand U22608 (N_22608,N_11183,N_10611);
and U22609 (N_22609,N_14380,N_16443);
nor U22610 (N_22610,N_17859,N_16464);
or U22611 (N_22611,N_19893,N_16867);
and U22612 (N_22612,N_10619,N_17033);
and U22613 (N_22613,N_16020,N_14789);
nor U22614 (N_22614,N_14090,N_12490);
nor U22615 (N_22615,N_17154,N_16384);
or U22616 (N_22616,N_18386,N_16875);
or U22617 (N_22617,N_14901,N_15398);
nand U22618 (N_22618,N_15613,N_10314);
nor U22619 (N_22619,N_19440,N_12963);
and U22620 (N_22620,N_18529,N_16491);
nor U22621 (N_22621,N_17536,N_19951);
nor U22622 (N_22622,N_12861,N_19385);
and U22623 (N_22623,N_12200,N_11513);
nand U22624 (N_22624,N_19838,N_18628);
and U22625 (N_22625,N_17777,N_17955);
nand U22626 (N_22626,N_18732,N_10884);
nand U22627 (N_22627,N_11338,N_19441);
and U22628 (N_22628,N_15853,N_13693);
nor U22629 (N_22629,N_11402,N_10629);
nor U22630 (N_22630,N_13815,N_10783);
and U22631 (N_22631,N_10262,N_14378);
or U22632 (N_22632,N_17354,N_10744);
nor U22633 (N_22633,N_12531,N_19392);
or U22634 (N_22634,N_13760,N_15736);
or U22635 (N_22635,N_16008,N_18492);
and U22636 (N_22636,N_10681,N_19292);
or U22637 (N_22637,N_17589,N_13985);
or U22638 (N_22638,N_18887,N_16671);
and U22639 (N_22639,N_17278,N_16392);
and U22640 (N_22640,N_19935,N_19355);
nand U22641 (N_22641,N_18439,N_17255);
and U22642 (N_22642,N_19889,N_11651);
or U22643 (N_22643,N_11133,N_11503);
nand U22644 (N_22644,N_17977,N_12634);
nor U22645 (N_22645,N_14631,N_14339);
nand U22646 (N_22646,N_15982,N_18419);
or U22647 (N_22647,N_15719,N_10625);
or U22648 (N_22648,N_14823,N_11391);
and U22649 (N_22649,N_10066,N_18144);
and U22650 (N_22650,N_15713,N_18299);
or U22651 (N_22651,N_14586,N_16617);
nor U22652 (N_22652,N_10346,N_16610);
or U22653 (N_22653,N_15192,N_16473);
nor U22654 (N_22654,N_16526,N_10985);
nand U22655 (N_22655,N_11775,N_18852);
and U22656 (N_22656,N_16029,N_19463);
or U22657 (N_22657,N_16006,N_15837);
nand U22658 (N_22658,N_17148,N_15285);
nand U22659 (N_22659,N_18740,N_15034);
xor U22660 (N_22660,N_13590,N_11002);
or U22661 (N_22661,N_16337,N_18892);
or U22662 (N_22662,N_13541,N_16912);
nor U22663 (N_22663,N_15984,N_14202);
and U22664 (N_22664,N_13947,N_10503);
or U22665 (N_22665,N_15869,N_14840);
and U22666 (N_22666,N_15624,N_19549);
nand U22667 (N_22667,N_17467,N_12778);
nor U22668 (N_22668,N_11020,N_19669);
and U22669 (N_22669,N_17856,N_19217);
nor U22670 (N_22670,N_18315,N_16804);
nor U22671 (N_22671,N_14238,N_10141);
or U22672 (N_22672,N_13284,N_13329);
or U22673 (N_22673,N_19614,N_14866);
nand U22674 (N_22674,N_13854,N_17125);
nand U22675 (N_22675,N_12911,N_10666);
nand U22676 (N_22676,N_10374,N_15334);
and U22677 (N_22677,N_17914,N_11971);
nand U22678 (N_22678,N_17779,N_10821);
or U22679 (N_22679,N_19909,N_10734);
nor U22680 (N_22680,N_18328,N_13651);
and U22681 (N_22681,N_18673,N_19857);
nor U22682 (N_22682,N_19776,N_16031);
nor U22683 (N_22683,N_16518,N_15691);
nor U22684 (N_22684,N_13066,N_11540);
and U22685 (N_22685,N_10550,N_16563);
and U22686 (N_22686,N_14250,N_14644);
and U22687 (N_22687,N_12056,N_18654);
nor U22688 (N_22688,N_16570,N_17598);
nor U22689 (N_22689,N_19580,N_17886);
nand U22690 (N_22690,N_14848,N_18003);
nand U22691 (N_22691,N_11065,N_14938);
nor U22692 (N_22692,N_12217,N_17730);
xor U22693 (N_22693,N_12525,N_10069);
nand U22694 (N_22694,N_15501,N_13105);
nand U22695 (N_22695,N_18826,N_17670);
nor U22696 (N_22696,N_17398,N_14340);
nand U22697 (N_22697,N_18022,N_14778);
or U22698 (N_22698,N_18491,N_15306);
or U22699 (N_22699,N_10182,N_14912);
nor U22700 (N_22700,N_19184,N_16896);
nor U22701 (N_22701,N_19298,N_17508);
or U22702 (N_22702,N_18101,N_12773);
xnor U22703 (N_22703,N_11837,N_14888);
or U22704 (N_22704,N_17360,N_17369);
and U22705 (N_22705,N_10654,N_14964);
and U22706 (N_22706,N_19188,N_16406);
or U22707 (N_22707,N_11790,N_13471);
nand U22708 (N_22708,N_14498,N_19575);
nor U22709 (N_22709,N_17048,N_12282);
nor U22710 (N_22710,N_10558,N_17865);
nand U22711 (N_22711,N_15113,N_10448);
or U22712 (N_22712,N_13093,N_14337);
nor U22713 (N_22713,N_15209,N_13425);
and U22714 (N_22714,N_12447,N_19963);
or U22715 (N_22715,N_13192,N_10545);
and U22716 (N_22716,N_15053,N_14916);
or U22717 (N_22717,N_10960,N_14573);
or U22718 (N_22718,N_17890,N_12323);
nand U22719 (N_22719,N_11771,N_19602);
nor U22720 (N_22720,N_13049,N_10027);
and U22721 (N_22721,N_11304,N_19232);
and U22722 (N_22722,N_14314,N_10976);
or U22723 (N_22723,N_15422,N_11810);
nand U22724 (N_22724,N_19250,N_15620);
nor U22725 (N_22725,N_18965,N_11265);
nand U22726 (N_22726,N_14895,N_14961);
or U22727 (N_22727,N_10298,N_14304);
nand U22728 (N_22728,N_19841,N_18877);
and U22729 (N_22729,N_15061,N_16727);
nand U22730 (N_22730,N_15511,N_13215);
nor U22731 (N_22731,N_10098,N_12693);
nor U22732 (N_22732,N_12908,N_11607);
nand U22733 (N_22733,N_10236,N_13117);
nor U22734 (N_22734,N_15580,N_15674);
nand U22735 (N_22735,N_11032,N_18941);
nand U22736 (N_22736,N_11440,N_19354);
nand U22737 (N_22737,N_13592,N_12142);
and U22738 (N_22738,N_14650,N_14385);
or U22739 (N_22739,N_14027,N_10052);
and U22740 (N_22740,N_15727,N_17542);
or U22741 (N_22741,N_14186,N_12343);
nand U22742 (N_22742,N_14287,N_17648);
or U22743 (N_22743,N_16413,N_11782);
nand U22744 (N_22744,N_11275,N_15618);
or U22745 (N_22745,N_17165,N_12533);
nand U22746 (N_22746,N_12076,N_16766);
and U22747 (N_22747,N_13505,N_16068);
nor U22748 (N_22748,N_16707,N_18244);
and U22749 (N_22749,N_13955,N_12969);
or U22750 (N_22750,N_15054,N_16681);
or U22751 (N_22751,N_15876,N_11571);
and U22752 (N_22752,N_11015,N_14049);
or U22753 (N_22753,N_13419,N_18548);
nor U22754 (N_22754,N_11066,N_13785);
and U22755 (N_22755,N_15543,N_13015);
and U22756 (N_22756,N_19758,N_10926);
nand U22757 (N_22757,N_10239,N_14559);
and U22758 (N_22758,N_15879,N_14084);
and U22759 (N_22759,N_16249,N_12092);
and U22760 (N_22760,N_14896,N_16083);
and U22761 (N_22761,N_19403,N_16805);
nand U22762 (N_22762,N_19931,N_12597);
and U22763 (N_22763,N_11008,N_13686);
and U22764 (N_22764,N_12144,N_13656);
nand U22765 (N_22765,N_17068,N_13597);
and U22766 (N_22766,N_19877,N_15591);
nand U22767 (N_22767,N_12211,N_10459);
nand U22768 (N_22768,N_14662,N_18445);
nor U22769 (N_22769,N_19224,N_15943);
and U22770 (N_22770,N_19734,N_14454);
nand U22771 (N_22771,N_11392,N_14376);
nand U22772 (N_22772,N_15894,N_13430);
nor U22773 (N_22773,N_10323,N_18829);
nand U22774 (N_22774,N_19954,N_18256);
nor U22775 (N_22775,N_16498,N_18294);
nor U22776 (N_22776,N_19572,N_15617);
or U22777 (N_22777,N_11044,N_11573);
and U22778 (N_22778,N_17963,N_12869);
or U22779 (N_22779,N_18997,N_18513);
and U22780 (N_22780,N_18282,N_16387);
or U22781 (N_22781,N_18559,N_18795);
or U22782 (N_22782,N_18298,N_14515);
nand U22783 (N_22783,N_14999,N_14550);
nand U22784 (N_22784,N_16099,N_16631);
nor U22785 (N_22785,N_17579,N_10133);
or U22786 (N_22786,N_15167,N_14696);
or U22787 (N_22787,N_13103,N_17639);
nor U22788 (N_22788,N_13530,N_10125);
nor U22789 (N_22789,N_12163,N_11999);
or U22790 (N_22790,N_11009,N_11216);
and U22791 (N_22791,N_17429,N_10901);
or U22792 (N_22792,N_12203,N_11424);
nand U22793 (N_22793,N_14727,N_16620);
nor U22794 (N_22794,N_13758,N_12271);
or U22795 (N_22795,N_10247,N_18300);
nand U22796 (N_22796,N_16294,N_11452);
and U22797 (N_22797,N_12012,N_11090);
nand U22798 (N_22798,N_12736,N_13935);
and U22799 (N_22799,N_15479,N_18713);
and U22800 (N_22800,N_17702,N_17013);
or U22801 (N_22801,N_14351,N_13437);
nor U22802 (N_22802,N_17196,N_19831);
or U22803 (N_22803,N_12127,N_16480);
or U22804 (N_22804,N_18218,N_11269);
or U22805 (N_22805,N_13121,N_15486);
and U22806 (N_22806,N_12897,N_19544);
or U22807 (N_22807,N_13130,N_16630);
nor U22808 (N_22808,N_13731,N_11100);
nor U22809 (N_22809,N_14558,N_17794);
nand U22810 (N_22810,N_10061,N_14805);
or U22811 (N_22811,N_18830,N_16332);
nand U22812 (N_22812,N_11805,N_16275);
and U22813 (N_22813,N_13487,N_18995);
nand U22814 (N_22814,N_14032,N_16728);
and U22815 (N_22815,N_10748,N_18810);
or U22816 (N_22816,N_16899,N_13350);
nand U22817 (N_22817,N_17607,N_13246);
nand U22818 (N_22818,N_14441,N_15637);
or U22819 (N_22819,N_13861,N_19600);
and U22820 (N_22820,N_14741,N_19231);
nand U22821 (N_22821,N_18834,N_13783);
nand U22822 (N_22822,N_17440,N_13516);
and U22823 (N_22823,N_11116,N_15112);
nor U22824 (N_22824,N_11961,N_17590);
and U22825 (N_22825,N_12638,N_11985);
nand U22826 (N_22826,N_12550,N_12950);
or U22827 (N_22827,N_14098,N_11506);
nor U22828 (N_22828,N_11669,N_10324);
or U22829 (N_22829,N_10270,N_13342);
nor U22830 (N_22830,N_11892,N_14290);
nor U22831 (N_22831,N_14853,N_16154);
or U22832 (N_22832,N_10455,N_13401);
nand U22833 (N_22833,N_10739,N_16892);
nand U22834 (N_22834,N_16715,N_16053);
nor U22835 (N_22835,N_15841,N_10777);
or U22836 (N_22836,N_15276,N_15944);
or U22837 (N_22837,N_18211,N_14091);
nand U22838 (N_22838,N_16566,N_11945);
and U22839 (N_22839,N_18804,N_15539);
nor U22840 (N_22840,N_13636,N_15911);
nor U22841 (N_22841,N_12380,N_17843);
or U22842 (N_22842,N_17158,N_18352);
nand U22843 (N_22843,N_12609,N_14480);
nand U22844 (N_22844,N_16366,N_19353);
nand U22845 (N_22845,N_17594,N_11950);
and U22846 (N_22846,N_17627,N_11043);
and U22847 (N_22847,N_15741,N_17030);
nor U22848 (N_22848,N_13716,N_17395);
nor U22849 (N_22849,N_12554,N_19591);
nor U22850 (N_22850,N_11211,N_10085);
nand U22851 (N_22851,N_19845,N_18407);
nor U22852 (N_22852,N_19994,N_16799);
and U22853 (N_22853,N_10439,N_18249);
and U22854 (N_22854,N_12954,N_14348);
or U22855 (N_22855,N_14459,N_19914);
nor U22856 (N_22856,N_15824,N_10986);
nand U22857 (N_22857,N_12758,N_15385);
nor U22858 (N_22858,N_15917,N_15173);
nand U22859 (N_22859,N_10765,N_11854);
nand U22860 (N_22860,N_17660,N_10348);
and U22861 (N_22861,N_11103,N_14195);
nor U22862 (N_22862,N_19045,N_14525);
nor U22863 (N_22863,N_12037,N_18087);
nand U22864 (N_22864,N_16806,N_17610);
and U22865 (N_22865,N_18378,N_15867);
or U22866 (N_22866,N_17798,N_18182);
nor U22867 (N_22867,N_17551,N_10944);
nand U22868 (N_22868,N_12665,N_19214);
or U22869 (N_22869,N_13588,N_11056);
nor U22870 (N_22870,N_15625,N_12822);
nand U22871 (N_22871,N_11764,N_19649);
or U22872 (N_22872,N_17351,N_15380);
and U22873 (N_22873,N_12074,N_18447);
nor U22874 (N_22874,N_14467,N_17678);
nor U22875 (N_22875,N_12159,N_11762);
or U22876 (N_22876,N_17816,N_11414);
or U22877 (N_22877,N_15222,N_15452);
nor U22878 (N_22878,N_12201,N_11101);
or U22879 (N_22879,N_11376,N_12767);
and U22880 (N_22880,N_12530,N_17913);
or U22881 (N_22881,N_18700,N_14426);
nor U22882 (N_22882,N_16525,N_15287);
nand U22883 (N_22883,N_18579,N_16499);
nand U22884 (N_22884,N_11174,N_16198);
nand U22885 (N_22885,N_18901,N_13982);
or U22886 (N_22886,N_16995,N_17706);
or U22887 (N_22887,N_10825,N_15463);
and U22888 (N_22888,N_18093,N_16845);
nor U22889 (N_22889,N_14239,N_10312);
or U22890 (N_22890,N_19465,N_13129);
nand U22891 (N_22891,N_16181,N_19082);
and U22892 (N_22892,N_17067,N_11484);
nand U22893 (N_22893,N_12303,N_12635);
nor U22894 (N_22894,N_16370,N_13896);
and U22895 (N_22895,N_17062,N_11938);
or U22896 (N_22896,N_18653,N_10256);
nand U22897 (N_22897,N_15865,N_13552);
or U22898 (N_22898,N_15206,N_13571);
and U22899 (N_22899,N_13390,N_18106);
nor U22900 (N_22900,N_14276,N_18031);
nand U22901 (N_22901,N_18546,N_19985);
nor U22902 (N_22902,N_14706,N_13377);
nor U22903 (N_22903,N_18293,N_16694);
and U22904 (N_22904,N_14652,N_11740);
or U22905 (N_22905,N_13073,N_14621);
nor U22906 (N_22906,N_17081,N_18602);
nor U22907 (N_22907,N_14154,N_12280);
or U22908 (N_22908,N_14242,N_13398);
nor U22909 (N_22909,N_13026,N_12220);
and U22910 (N_22910,N_13148,N_19102);
nor U22911 (N_22911,N_19163,N_14751);
xnor U22912 (N_22912,N_14432,N_19993);
or U22913 (N_22913,N_11115,N_18915);
nand U22914 (N_22914,N_15866,N_16159);
and U22915 (N_22915,N_14388,N_10958);
nand U22916 (N_22916,N_10211,N_17109);
and U22917 (N_22917,N_11665,N_18797);
and U22918 (N_22918,N_15442,N_18517);
nor U22919 (N_22919,N_17891,N_14802);
nand U22920 (N_22920,N_18424,N_11877);
nand U22921 (N_22921,N_14194,N_19933);
or U22922 (N_22922,N_12703,N_10661);
nor U22923 (N_22923,N_18685,N_17382);
and U22924 (N_22924,N_15658,N_16182);
or U22925 (N_22925,N_12914,N_14338);
nor U22926 (N_22926,N_10598,N_17818);
and U22927 (N_22927,N_13366,N_17724);
or U22928 (N_22928,N_16692,N_11221);
nor U22929 (N_22929,N_14522,N_13641);
or U22930 (N_22930,N_16028,N_10695);
and U22931 (N_22931,N_18136,N_14681);
and U22932 (N_22932,N_12802,N_18749);
nor U22933 (N_22933,N_19953,N_15675);
or U22934 (N_22934,N_15374,N_16623);
nor U22935 (N_22935,N_11739,N_12643);
or U22936 (N_22936,N_18637,N_19477);
nor U22937 (N_22937,N_18688,N_11281);
and U22938 (N_22938,N_12386,N_16528);
nand U22939 (N_22939,N_14816,N_17936);
nand U22940 (N_22940,N_18914,N_16559);
or U22941 (N_22941,N_13394,N_12864);
or U22942 (N_22942,N_17365,N_11502);
and U22943 (N_22943,N_12584,N_19599);
or U22944 (N_22944,N_18668,N_19663);
nor U22945 (N_22945,N_10607,N_19148);
or U22946 (N_22946,N_18770,N_14404);
or U22947 (N_22947,N_10936,N_18463);
nor U22948 (N_22948,N_16364,N_18884);
or U22949 (N_22949,N_10151,N_10929);
or U22950 (N_22950,N_14208,N_14002);
or U22951 (N_22951,N_14087,N_15608);
or U22952 (N_22952,N_13871,N_15827);
nor U22953 (N_22953,N_12853,N_19869);
or U22954 (N_22954,N_10214,N_13916);
and U22955 (N_22955,N_14444,N_13126);
nor U22956 (N_22956,N_15928,N_13868);
nor U22957 (N_22957,N_11623,N_11690);
nor U22958 (N_22958,N_15621,N_19358);
nand U22959 (N_22959,N_13517,N_13151);
nand U22960 (N_22960,N_19783,N_19081);
nand U22961 (N_22961,N_12923,N_13173);
nand U22962 (N_22962,N_14804,N_12697);
or U22963 (N_22963,N_12259,N_16293);
nand U22964 (N_22964,N_16376,N_15900);
nand U22965 (N_22965,N_14311,N_16259);
or U22966 (N_22966,N_16998,N_15329);
and U22967 (N_22967,N_14587,N_11542);
and U22968 (N_22968,N_10195,N_15315);
or U22969 (N_22969,N_16601,N_17322);
nor U22970 (N_22970,N_13660,N_11330);
nor U22971 (N_22971,N_17099,N_12242);
and U22972 (N_22972,N_19676,N_11004);
nor U22973 (N_22973,N_12307,N_19197);
or U22974 (N_22974,N_18341,N_14835);
nand U22975 (N_22975,N_12054,N_16148);
or U22976 (N_22976,N_18037,N_17561);
and U22977 (N_22977,N_12499,N_19902);
nor U22978 (N_22978,N_15105,N_18044);
nand U22979 (N_22979,N_17604,N_10890);
nand U22980 (N_22980,N_14563,N_12104);
nand U22981 (N_22981,N_17570,N_18051);
nor U22982 (N_22982,N_19830,N_13347);
nor U22983 (N_22983,N_16751,N_13953);
nand U22984 (N_22984,N_11137,N_13712);
nand U22985 (N_22985,N_19422,N_15207);
nand U22986 (N_22986,N_13480,N_11944);
and U22987 (N_22987,N_16786,N_12631);
or U22988 (N_22988,N_13003,N_11899);
and U22989 (N_22989,N_10468,N_12297);
or U22990 (N_22990,N_18921,N_15087);
and U22991 (N_22991,N_10507,N_18658);
or U22992 (N_22992,N_17728,N_15168);
nor U22993 (N_22993,N_10937,N_14085);
or U22994 (N_22994,N_15789,N_11592);
and U22995 (N_22995,N_12031,N_17676);
and U22996 (N_22996,N_19706,N_16287);
nand U22997 (N_22997,N_19125,N_13991);
or U22998 (N_22998,N_12006,N_12866);
nand U22999 (N_22999,N_10121,N_18074);
or U23000 (N_23000,N_17359,N_11435);
xor U23001 (N_23001,N_18420,N_13573);
or U23002 (N_23002,N_15023,N_13373);
nor U23003 (N_23003,N_17039,N_18376);
nand U23004 (N_23004,N_17086,N_16475);
or U23005 (N_23005,N_19044,N_10868);
nand U23006 (N_23006,N_16047,N_16408);
nor U23007 (N_23007,N_19887,N_15272);
or U23008 (N_23008,N_19536,N_12319);
nor U23009 (N_23009,N_16172,N_19762);
or U23010 (N_23010,N_15472,N_17640);
and U23011 (N_23011,N_13499,N_17858);
and U23012 (N_23012,N_15852,N_13672);
or U23013 (N_23013,N_18634,N_10112);
and U23014 (N_23014,N_17166,N_19367);
nand U23015 (N_23015,N_12686,N_11637);
and U23016 (N_23016,N_16955,N_15130);
nand U23017 (N_23017,N_13110,N_16626);
or U23018 (N_23018,N_13243,N_15282);
or U23019 (N_23019,N_16904,N_11492);
and U23020 (N_23020,N_10398,N_14237);
and U23021 (N_23021,N_14807,N_19670);
and U23022 (N_23022,N_15584,N_11179);
nor U23023 (N_23023,N_17288,N_15768);
and U23024 (N_23024,N_15320,N_11930);
nor U23025 (N_23025,N_17422,N_13271);
nor U23026 (N_23026,N_17204,N_19142);
and U23027 (N_23027,N_17418,N_18836);
and U23028 (N_23028,N_16017,N_18550);
and U23029 (N_23029,N_19307,N_11841);
and U23030 (N_23030,N_13507,N_14641);
and U23031 (N_23031,N_12462,N_13930);
nand U23032 (N_23032,N_19116,N_14188);
and U23033 (N_23033,N_14611,N_13063);
nor U23034 (N_23034,N_15567,N_14175);
nand U23035 (N_23035,N_14220,N_12842);
and U23036 (N_23036,N_12682,N_14012);
and U23037 (N_23037,N_12064,N_19548);
or U23038 (N_23038,N_12312,N_16336);
nand U23039 (N_23039,N_15468,N_13492);
or U23040 (N_23040,N_19564,N_11924);
nand U23041 (N_23041,N_17527,N_15581);
nand U23042 (N_23042,N_19218,N_13642);
nor U23043 (N_23043,N_13576,N_17381);
and U23044 (N_23044,N_17679,N_17821);
nor U23045 (N_23045,N_13005,N_12045);
nor U23046 (N_23046,N_19858,N_19311);
or U23047 (N_23047,N_17363,N_16326);
nand U23048 (N_23048,N_10396,N_13009);
nand U23049 (N_23049,N_16268,N_13359);
and U23050 (N_23050,N_16049,N_16100);
nand U23051 (N_23051,N_11322,N_15360);
or U23052 (N_23052,N_17904,N_18114);
or U23053 (N_23053,N_13082,N_12868);
and U23054 (N_23054,N_14939,N_14042);
and U23055 (N_23055,N_18242,N_17214);
nor U23056 (N_23056,N_18092,N_11098);
and U23057 (N_23057,N_19542,N_17063);
nor U23058 (N_23058,N_15044,N_11359);
nor U23059 (N_23059,N_13849,N_18088);
nor U23060 (N_23060,N_14004,N_10952);
nor U23061 (N_23061,N_17228,N_15498);
nor U23062 (N_23062,N_11314,N_13260);
or U23063 (N_23063,N_19846,N_16680);
or U23064 (N_23064,N_19740,N_16218);
and U23065 (N_23065,N_12396,N_18946);
or U23066 (N_23066,N_13199,N_15669);
and U23067 (N_23067,N_16292,N_11756);
and U23068 (N_23068,N_12034,N_10371);
or U23069 (N_23069,N_15305,N_19414);
and U23070 (N_23070,N_15971,N_10354);
nor U23071 (N_23071,N_19149,N_13753);
nor U23072 (N_23072,N_17543,N_11488);
or U23073 (N_23073,N_11906,N_19228);
or U23074 (N_23074,N_15068,N_16190);
and U23075 (N_23075,N_18033,N_14074);
or U23076 (N_23076,N_16795,N_15096);
nand U23077 (N_23077,N_18960,N_12598);
or U23078 (N_23078,N_17019,N_19556);
or U23079 (N_23079,N_11169,N_12630);
and U23080 (N_23080,N_10907,N_13721);
nor U23081 (N_23081,N_11650,N_16865);
or U23082 (N_23082,N_15408,N_19303);
nand U23083 (N_23083,N_18015,N_17150);
and U23084 (N_23084,N_15589,N_16458);
nand U23085 (N_23085,N_19805,N_14554);
nor U23086 (N_23086,N_12438,N_16389);
nand U23087 (N_23087,N_15036,N_15490);
nor U23088 (N_23088,N_16340,N_11561);
and U23089 (N_23089,N_14716,N_19532);
or U23090 (N_23090,N_16569,N_16688);
nor U23091 (N_23091,N_15965,N_14386);
nor U23092 (N_23092,N_11984,N_19308);
or U23093 (N_23093,N_10013,N_14513);
nor U23094 (N_23094,N_16402,N_11319);
or U23095 (N_23095,N_15781,N_19565);
or U23096 (N_23096,N_12557,N_19871);
or U23097 (N_23097,N_17663,N_13111);
nor U23098 (N_23098,N_15238,N_17233);
nor U23099 (N_23099,N_10289,N_17029);
nand U23100 (N_23100,N_10812,N_14608);
xnor U23101 (N_23101,N_13433,N_15733);
nor U23102 (N_23102,N_11445,N_19826);
or U23103 (N_23103,N_15535,N_19129);
or U23104 (N_23104,N_19917,N_19864);
or U23105 (N_23105,N_12145,N_15588);
and U23106 (N_23106,N_17685,N_17443);
and U23107 (N_23107,N_11970,N_10464);
nor U23108 (N_23108,N_12915,N_15473);
nor U23109 (N_23109,N_18661,N_15919);
and U23110 (N_23110,N_19563,N_18703);
and U23111 (N_23111,N_10578,N_13016);
nand U23112 (N_23112,N_13076,N_18461);
nor U23113 (N_23113,N_11236,N_10001);
nand U23114 (N_23114,N_10587,N_11868);
nand U23115 (N_23115,N_11429,N_14837);
or U23116 (N_23116,N_19161,N_16137);
nor U23117 (N_23117,N_15198,N_19952);
or U23118 (N_23118,N_11099,N_14458);
nor U23119 (N_23119,N_15058,N_12805);
nor U23120 (N_23120,N_15747,N_19473);
and U23121 (N_23121,N_19743,N_17618);
nand U23122 (N_23122,N_12296,N_13298);
or U23123 (N_23123,N_17080,N_10191);
or U23124 (N_23124,N_10352,N_12402);
or U23125 (N_23125,N_17328,N_15101);
or U23126 (N_23126,N_13666,N_12640);
or U23127 (N_23127,N_17061,N_10296);
or U23128 (N_23128,N_18444,N_18831);
or U23129 (N_23129,N_17151,N_16119);
nand U23130 (N_23130,N_10888,N_19280);
nand U23131 (N_23131,N_15787,N_10482);
or U23132 (N_23132,N_17547,N_14445);
and U23133 (N_23133,N_14747,N_14850);
nand U23134 (N_23134,N_10731,N_13128);
nor U23135 (N_23135,N_10994,N_15190);
and U23136 (N_23136,N_19586,N_16939);
nand U23137 (N_23137,N_12509,N_15989);
and U23138 (N_23138,N_19478,N_18178);
or U23139 (N_23139,N_18245,N_10002);
and U23140 (N_23140,N_13954,N_18882);
nand U23141 (N_23141,N_15975,N_16311);
nand U23142 (N_23142,N_12580,N_10064);
nor U23143 (N_23143,N_15313,N_16453);
and U23144 (N_23144,N_19643,N_15063);
and U23145 (N_23145,N_19400,N_11172);
and U23146 (N_23146,N_19167,N_19140);
and U23147 (N_23147,N_11196,N_19406);
nand U23148 (N_23148,N_15797,N_10472);
or U23149 (N_23149,N_10131,N_16122);
nand U23150 (N_23150,N_11385,N_15893);
and U23151 (N_23151,N_14879,N_11348);
nand U23152 (N_23152,N_18779,N_11819);
nand U23153 (N_23153,N_17329,N_12641);
nor U23154 (N_23154,N_14017,N_19653);
and U23155 (N_23155,N_17760,N_10278);
and U23156 (N_23156,N_15868,N_14125);
nand U23157 (N_23157,N_18364,N_18638);
nand U23158 (N_23158,N_14097,N_18167);
nor U23159 (N_23159,N_11539,N_10007);
nand U23160 (N_23160,N_17057,N_14306);
and U23161 (N_23161,N_19076,N_15344);
nor U23162 (N_23162,N_14736,N_12672);
or U23163 (N_23163,N_15961,N_12626);
and U23164 (N_23164,N_10199,N_17709);
or U23165 (N_23165,N_17988,N_19804);
and U23166 (N_23166,N_13353,N_11838);
nand U23167 (N_23167,N_12561,N_17450);
nor U23168 (N_23168,N_13893,N_16764);
nand U23169 (N_23169,N_14642,N_14832);
or U23170 (N_23170,N_13676,N_12595);
and U23171 (N_23171,N_17199,N_14733);
nor U23172 (N_23172,N_14124,N_12361);
nor U23173 (N_23173,N_18202,N_14355);
and U23174 (N_23174,N_13884,N_10204);
and U23175 (N_23175,N_12011,N_11076);
or U23176 (N_23176,N_12466,N_16662);
and U23177 (N_23177,N_13184,N_15416);
nor U23178 (N_23178,N_16138,N_15880);
nor U23179 (N_23179,N_10742,N_19071);
nand U23180 (N_23180,N_12080,N_11886);
or U23181 (N_23181,N_18676,N_16116);
nor U23182 (N_23182,N_18235,N_18765);
nand U23183 (N_23183,N_13843,N_11580);
and U23184 (N_23184,N_14945,N_17435);
and U23185 (N_23185,N_14904,N_10899);
and U23186 (N_23186,N_13531,N_10839);
or U23187 (N_23187,N_19579,N_10580);
and U23188 (N_23188,N_14527,N_13483);
and U23189 (N_23189,N_13448,N_15081);
or U23190 (N_23190,N_16820,N_12906);
and U23191 (N_23191,N_18927,N_16030);
nor U23192 (N_23192,N_15632,N_12155);
nor U23193 (N_23193,N_10637,N_17860);
or U23194 (N_23194,N_12999,N_12384);
and U23195 (N_23195,N_18168,N_17310);
nor U23196 (N_23196,N_18537,N_13832);
nand U23197 (N_23197,N_10930,N_16114);
nor U23198 (N_23198,N_16510,N_16232);
nand U23199 (N_23199,N_13040,N_14083);
and U23200 (N_23200,N_16810,N_10484);
and U23201 (N_23201,N_15354,N_19174);
or U23202 (N_23202,N_14267,N_12860);
nand U23203 (N_23203,N_13497,N_15647);
nor U23204 (N_23204,N_12886,N_17995);
nor U23205 (N_23205,N_10692,N_19859);
nor U23206 (N_23206,N_10240,N_18619);
nor U23207 (N_23207,N_11092,N_18115);
nand U23208 (N_23208,N_12857,N_11871);
and U23209 (N_23209,N_17110,N_11342);
or U23210 (N_23210,N_12560,N_18310);
or U23211 (N_23211,N_11590,N_19288);
or U23212 (N_23212,N_10146,N_19886);
and U23213 (N_23213,N_18253,N_15724);
or U23214 (N_23214,N_12739,N_16915);
nor U23215 (N_23215,N_19080,N_18585);
nor U23216 (N_23216,N_18125,N_14518);
or U23217 (N_23217,N_17293,N_16113);
nand U23218 (N_23218,N_12859,N_16798);
and U23219 (N_23219,N_11617,N_19432);
nor U23220 (N_23220,N_18017,N_10851);
and U23221 (N_23221,N_14687,N_18288);
nor U23222 (N_23222,N_13781,N_10094);
or U23223 (N_23223,N_18776,N_11797);
or U23224 (N_23224,N_15836,N_15888);
and U23225 (N_23225,N_12416,N_18421);
and U23226 (N_23226,N_14342,N_10393);
nor U23227 (N_23227,N_18103,N_13055);
or U23228 (N_23228,N_10690,N_12845);
or U23229 (N_23229,N_15072,N_14520);
nor U23230 (N_23230,N_15316,N_12434);
or U23231 (N_23231,N_13176,N_19521);
nor U23232 (N_23232,N_12458,N_17225);
xor U23233 (N_23233,N_14086,N_12948);
nand U23234 (N_23234,N_18208,N_13554);
and U23235 (N_23235,N_13388,N_12408);
nand U23236 (N_23236,N_11928,N_15491);
or U23237 (N_23237,N_17987,N_12081);
nand U23238 (N_23238,N_13488,N_16738);
and U23239 (N_23239,N_17383,N_17180);
or U23240 (N_23240,N_11372,N_15433);
or U23241 (N_23241,N_11351,N_11373);
nor U23242 (N_23242,N_19659,N_17184);
nand U23243 (N_23243,N_17564,N_11363);
and U23244 (N_23244,N_14105,N_15935);
or U23245 (N_23245,N_10745,N_15268);
and U23246 (N_23246,N_16355,N_16374);
or U23247 (N_23247,N_14750,N_15901);
and U23248 (N_23248,N_16051,N_17802);
or U23249 (N_23249,N_15059,N_15506);
nor U23250 (N_23250,N_17237,N_12267);
or U23251 (N_23251,N_18737,N_10471);
nor U23252 (N_23252,N_18499,N_16822);
and U23253 (N_23253,N_13952,N_12391);
nor U23254 (N_23254,N_13857,N_13187);
nand U23255 (N_23255,N_13888,N_17558);
and U23256 (N_23256,N_17178,N_16693);
or U23257 (N_23257,N_17419,N_14688);
or U23258 (N_23258,N_15005,N_10130);
nor U23259 (N_23259,N_18889,N_10213);
xnor U23260 (N_23260,N_13147,N_10900);
nand U23261 (N_23261,N_17586,N_10097);
nand U23262 (N_23262,N_10362,N_11327);
or U23263 (N_23263,N_12058,N_14724);
nor U23264 (N_23264,N_13475,N_10473);
or U23265 (N_23265,N_17864,N_10656);
nor U23266 (N_23266,N_13454,N_18937);
or U23267 (N_23267,N_16001,N_14784);
xor U23268 (N_23268,N_12681,N_17014);
nor U23269 (N_23269,N_14880,N_17051);
or U23270 (N_23270,N_11721,N_10442);
nor U23271 (N_23271,N_16054,N_11270);
and U23272 (N_23272,N_19480,N_12724);
or U23273 (N_23273,N_10895,N_15372);
nor U23274 (N_23274,N_17119,N_11463);
nand U23275 (N_23275,N_16131,N_19242);
and U23276 (N_23276,N_13200,N_12321);
or U23277 (N_23277,N_19126,N_19339);
or U23278 (N_23278,N_17076,N_11147);
and U23279 (N_23279,N_17426,N_10313);
or U23280 (N_23280,N_18133,N_13322);
nand U23281 (N_23281,N_14581,N_17571);
and U23282 (N_23282,N_13812,N_12359);
nand U23283 (N_23283,N_12229,N_13848);
nor U23284 (N_23284,N_12636,N_15962);
nor U23285 (N_23285,N_19455,N_14564);
nor U23286 (N_23286,N_16152,N_16765);
nand U23287 (N_23287,N_15645,N_10368);
and U23288 (N_23288,N_13558,N_18032);
and U23289 (N_23289,N_15177,N_14720);
or U23290 (N_23290,N_10572,N_17261);
nor U23291 (N_23291,N_12879,N_12123);
and U23292 (N_23292,N_14645,N_11189);
nor U23293 (N_23293,N_16753,N_17229);
and U23294 (N_23294,N_15903,N_12642);
nor U23295 (N_23295,N_18270,N_15627);
and U23296 (N_23296,N_11828,N_17584);
and U23297 (N_23297,N_12740,N_16385);
or U23298 (N_23298,N_11933,N_16769);
or U23299 (N_23299,N_15172,N_12825);
nand U23300 (N_23300,N_13146,N_18496);
or U23301 (N_23301,N_16488,N_15164);
and U23302 (N_23302,N_16922,N_12376);
or U23303 (N_23303,N_16173,N_12214);
or U23304 (N_23304,N_16090,N_10854);
or U23305 (N_23305,N_19048,N_15949);
or U23306 (N_23306,N_14833,N_17239);
nor U23307 (N_23307,N_11120,N_18066);
nor U23308 (N_23308,N_16971,N_19746);
nor U23309 (N_23309,N_10769,N_12440);
nand U23310 (N_23310,N_12414,N_14479);
or U23311 (N_23311,N_17947,N_13623);
nand U23312 (N_23312,N_12260,N_17666);
and U23313 (N_23313,N_17502,N_15097);
or U23314 (N_23314,N_18457,N_10242);
nand U23315 (N_23315,N_15076,N_10149);
or U23316 (N_23316,N_14172,N_17453);
or U23317 (N_23317,N_14354,N_19798);
or U23318 (N_23318,N_16545,N_19551);
nor U23319 (N_23319,N_13025,N_15870);
nand U23320 (N_23320,N_18692,N_15715);
or U23321 (N_23321,N_15931,N_18231);
nand U23322 (N_23322,N_11182,N_18045);
and U23323 (N_23323,N_15697,N_11459);
and U23324 (N_23324,N_17991,N_16988);
and U23325 (N_23325,N_16442,N_12009);
nand U23326 (N_23326,N_14754,N_18224);
or U23327 (N_23327,N_10208,N_18060);
nand U23328 (N_23328,N_17130,N_15220);
and U23329 (N_23329,N_13335,N_12097);
nand U23330 (N_23330,N_19593,N_17708);
or U23331 (N_23331,N_18261,N_13831);
or U23332 (N_23332,N_13305,N_17056);
nor U23333 (N_23333,N_14982,N_10280);
or U23334 (N_23334,N_14066,N_18572);
nor U23335 (N_23335,N_13327,N_11150);
and U23336 (N_23336,N_19861,N_15564);
or U23337 (N_23337,N_12117,N_16214);
and U23338 (N_23338,N_15070,N_11769);
nor U23339 (N_23339,N_13244,N_17758);
and U23340 (N_23340,N_17430,N_17562);
or U23341 (N_23341,N_14589,N_16009);
nor U23342 (N_23342,N_19277,N_15732);
and U23343 (N_23343,N_16776,N_18790);
nor U23344 (N_23344,N_11780,N_11441);
and U23345 (N_23345,N_18861,N_19021);
nor U23346 (N_23346,N_12067,N_16542);
and U23347 (N_23347,N_18233,N_14111);
nand U23348 (N_23348,N_19008,N_11559);
nor U23349 (N_23349,N_16315,N_11345);
or U23350 (N_23350,N_11474,N_13085);
or U23351 (N_23351,N_15370,N_13012);
nor U23352 (N_23352,N_11543,N_11591);
or U23353 (N_23353,N_14191,N_18675);
nor U23354 (N_23354,N_12810,N_19476);
and U23355 (N_23355,N_14598,N_19515);
nand U23356 (N_23356,N_13222,N_11192);
nand U23357 (N_23357,N_15257,N_16074);
or U23358 (N_23358,N_19168,N_10684);
nor U23359 (N_23359,N_18681,N_17449);
and U23360 (N_23360,N_16589,N_17059);
and U23361 (N_23361,N_16697,N_15964);
or U23362 (N_23362,N_16299,N_19490);
or U23363 (N_23363,N_16588,N_13122);
nand U23364 (N_23364,N_16879,N_17090);
nand U23365 (N_23365,N_13532,N_12910);
and U23366 (N_23366,N_11616,N_16607);
and U23367 (N_23367,N_16568,N_12505);
nor U23368 (N_23368,N_11284,N_19094);
and U23369 (N_23369,N_13818,N_16034);
nor U23370 (N_23370,N_15942,N_14808);
or U23371 (N_23371,N_11783,N_19099);
and U23372 (N_23372,N_10100,N_10577);
nand U23373 (N_23373,N_10579,N_11691);
or U23374 (N_23374,N_14944,N_16714);
or U23375 (N_23375,N_13240,N_19808);
nand U23376 (N_23376,N_15673,N_17205);
nor U23377 (N_23377,N_16132,N_10103);
nand U23378 (N_23378,N_13208,N_12674);
nor U23379 (N_23379,N_15717,N_13250);
nor U23380 (N_23380,N_12108,N_17624);
nand U23381 (N_23381,N_13174,N_10616);
nand U23382 (N_23382,N_17553,N_13253);
or U23383 (N_23383,N_12727,N_17767);
or U23384 (N_23384,N_16378,N_19610);
nor U23385 (N_23385,N_18488,N_12620);
nor U23386 (N_23386,N_17388,N_18221);
or U23387 (N_23387,N_19644,N_14794);
and U23388 (N_23388,N_19822,N_11290);
nor U23389 (N_23389,N_18297,N_17022);
nand U23390 (N_23390,N_15230,N_15080);
and U23391 (N_23391,N_10506,N_12903);
or U23392 (N_23392,N_18484,N_14948);
and U23393 (N_23393,N_19489,N_18304);
or U23394 (N_23394,N_13330,N_19794);
nor U23395 (N_23395,N_17289,N_17964);
or U23396 (N_23396,N_12090,N_19925);
nand U23397 (N_23397,N_15923,N_18862);
nor U23398 (N_23398,N_13951,N_17623);
or U23399 (N_23399,N_16050,N_15510);
nand U23400 (N_23400,N_13684,N_12799);
xor U23401 (N_23401,N_14193,N_13356);
nand U23402 (N_23402,N_11576,N_19278);
and U23403 (N_23403,N_11431,N_10523);
nand U23404 (N_23404,N_12673,N_19470);
nand U23405 (N_23405,N_18429,N_12381);
nor U23406 (N_23406,N_17302,N_18394);
nand U23407 (N_23407,N_15654,N_18553);
and U23408 (N_23408,N_13737,N_16077);
nand U23409 (N_23409,N_15000,N_10714);
and U23410 (N_23410,N_14864,N_13671);
nand U23411 (N_23411,N_10451,N_10792);
nand U23412 (N_23412,N_19926,N_16177);
nand U23413 (N_23413,N_11469,N_18258);
or U23414 (N_23414,N_19714,N_18223);
nand U23415 (N_23415,N_14271,N_14745);
and U23416 (N_23416,N_17280,N_10627);
or U23417 (N_23417,N_14006,N_16441);
and U23418 (N_23418,N_18636,N_11393);
and U23419 (N_23419,N_17053,N_11329);
nor U23420 (N_23420,N_19853,N_18369);
or U23421 (N_23421,N_18723,N_14593);
nand U23422 (N_23422,N_12313,N_18596);
nor U23423 (N_23423,N_15141,N_10350);
or U23424 (N_23424,N_18192,N_19986);
or U23425 (N_23425,N_19524,N_16434);
or U23426 (N_23426,N_17861,N_18285);
nand U23427 (N_23427,N_17521,N_11165);
or U23428 (N_23428,N_12339,N_15878);
nand U23429 (N_23429,N_16539,N_14690);
and U23430 (N_23430,N_10065,N_11178);
or U23431 (N_23431,N_14283,N_10592);
and U23432 (N_23432,N_15607,N_14625);
nand U23433 (N_23433,N_17772,N_10563);
and U23434 (N_23434,N_11926,N_12422);
nor U23435 (N_23435,N_15874,N_17587);
and U23436 (N_23436,N_15612,N_17120);
or U23437 (N_23437,N_14041,N_16205);
nand U23438 (N_23438,N_18624,N_19687);
nand U23439 (N_23439,N_11190,N_10741);
nor U23440 (N_23440,N_18845,N_12629);
nand U23441 (N_23441,N_10479,N_19079);
nand U23442 (N_23442,N_17793,N_13824);
nor U23443 (N_23443,N_18642,N_10967);
or U23444 (N_23444,N_17308,N_14890);
or U23445 (N_23445,N_11827,N_14411);
nand U23446 (N_23446,N_13045,N_14801);
nand U23447 (N_23447,N_11387,N_11794);
nor U23448 (N_23448,N_10341,N_18353);
and U23449 (N_23449,N_19750,N_14205);
and U23450 (N_23450,N_18625,N_10914);
or U23451 (N_23451,N_10203,N_12284);
or U23452 (N_23452,N_15075,N_17970);
or U23453 (N_23453,N_13064,N_19464);
nor U23454 (N_23454,N_16244,N_12363);
nand U23455 (N_23455,N_16349,N_10123);
nor U23456 (N_23456,N_12066,N_13917);
or U23457 (N_23457,N_10889,N_18206);
or U23458 (N_23458,N_17878,N_16204);
or U23459 (N_23459,N_14133,N_19751);
nand U23460 (N_23460,N_15225,N_16585);
or U23461 (N_23461,N_10843,N_16629);
and U23462 (N_23462,N_17028,N_14684);
or U23463 (N_23463,N_19305,N_11720);
and U23464 (N_23464,N_12305,N_12894);
nor U23465 (N_23465,N_11104,N_13877);
nor U23466 (N_23466,N_16237,N_12378);
nor U23467 (N_23467,N_10143,N_10076);
nor U23468 (N_23468,N_17000,N_15239);
nor U23469 (N_23469,N_19675,N_16637);
nand U23470 (N_23470,N_13324,N_12990);
or U23471 (N_23471,N_17122,N_10845);
and U23472 (N_23472,N_16351,N_18159);
and U23473 (N_23473,N_12017,N_14018);
and U23474 (N_23474,N_12461,N_14118);
nand U23475 (N_23475,N_15138,N_14620);
nor U23476 (N_23476,N_11287,N_15765);
nand U23477 (N_23477,N_15711,N_15352);
and U23478 (N_23478,N_10547,N_18803);
or U23479 (N_23479,N_10318,N_14860);
nand U23480 (N_23480,N_13940,N_16723);
nor U23481 (N_23481,N_17102,N_10983);
or U23482 (N_23482,N_17791,N_10273);
and U23483 (N_23483,N_13417,N_12746);
or U23484 (N_23484,N_15983,N_11631);
nand U23485 (N_23485,N_18180,N_12412);
nor U23486 (N_23486,N_15810,N_13416);
nand U23487 (N_23487,N_16917,N_16960);
or U23488 (N_23488,N_18286,N_19018);
or U23489 (N_23489,N_17173,N_18593);
and U23490 (N_23490,N_14014,N_12338);
or U23491 (N_23491,N_19546,N_17915);
nand U23492 (N_23492,N_12548,N_12226);
or U23493 (N_23493,N_15197,N_11205);
nor U23494 (N_23494,N_10740,N_12125);
or U23495 (N_23495,N_15762,N_16367);
nand U23496 (N_23496,N_15782,N_14395);
or U23497 (N_23497,N_12413,N_12350);
or U23498 (N_23498,N_13150,N_14659);
and U23499 (N_23499,N_16420,N_11018);
or U23500 (N_23500,N_17999,N_11729);
nand U23501 (N_23501,N_19820,N_10235);
nand U23502 (N_23502,N_10018,N_18149);
nor U23503 (N_23503,N_13370,N_16552);
and U23504 (N_23504,N_11922,N_14721);
or U23505 (N_23505,N_10931,N_18451);
nand U23506 (N_23506,N_14818,N_12000);
nor U23507 (N_23507,N_18598,N_18154);
or U23508 (N_23508,N_18825,N_16298);
and U23509 (N_23509,N_14243,N_17661);
and U23510 (N_23510,N_10670,N_19626);
and U23511 (N_23511,N_16746,N_18175);
and U23512 (N_23512,N_13911,N_18626);
nor U23513 (N_23513,N_10975,N_19285);
nand U23514 (N_23514,N_19123,N_15208);
nand U23515 (N_23515,N_11017,N_18187);
nand U23516 (N_23516,N_17295,N_13864);
nand U23517 (N_23517,N_10023,N_14349);
or U23518 (N_23518,N_18483,N_18938);
or U23519 (N_23519,N_14334,N_19172);
nand U23520 (N_23520,N_18006,N_14094);
and U23521 (N_23521,N_13806,N_17720);
or U23522 (N_23522,N_18415,N_10602);
nor U23523 (N_23523,N_11231,N_19193);
or U23524 (N_23524,N_10877,N_12813);
and U23525 (N_23525,N_15260,N_16352);
and U23526 (N_23526,N_13866,N_14568);
nor U23527 (N_23527,N_19637,N_13395);
or U23528 (N_23528,N_14137,N_12007);
or U23529 (N_23529,N_13044,N_13462);
and U23530 (N_23530,N_15418,N_18580);
nor U23531 (N_23531,N_12887,N_16324);
and U23532 (N_23532,N_19566,N_19204);
or U23533 (N_23533,N_10699,N_14788);
or U23534 (N_23534,N_11977,N_16269);
or U23535 (N_23535,N_15233,N_18926);
or U23536 (N_23536,N_19918,N_15119);
or U23537 (N_23537,N_16197,N_14285);
nor U23538 (N_23538,N_15392,N_14360);
nand U23539 (N_23539,N_14633,N_14062);
nor U23540 (N_23540,N_17524,N_14072);
and U23541 (N_23541,N_18840,N_16107);
and U23542 (N_23542,N_15417,N_16286);
and U23543 (N_23543,N_10750,N_11550);
and U23544 (N_23544,N_12213,N_12826);
or U23545 (N_23545,N_16576,N_16391);
nand U23546 (N_23546,N_17475,N_10924);
and U23547 (N_23547,N_17445,N_12732);
and U23548 (N_23548,N_17338,N_18614);
nor U23549 (N_23549,N_10177,N_11847);
nand U23550 (N_23550,N_11713,N_17137);
nand U23551 (N_23551,N_11218,N_10998);
nand U23552 (N_23552,N_16066,N_13795);
or U23553 (N_23553,N_17636,N_15153);
and U23554 (N_23554,N_17290,N_13172);
or U23555 (N_23555,N_15324,N_10285);
and U23556 (N_23556,N_18973,N_11983);
nand U23557 (N_23557,N_14872,N_15939);
nor U23558 (N_23558,N_10397,N_13071);
nor U23559 (N_23559,N_12844,N_18621);
or U23560 (N_23560,N_19386,N_11289);
nor U23561 (N_23561,N_16479,N_19325);
nor U23562 (N_23562,N_19101,N_17870);
or U23563 (N_23563,N_10385,N_12060);
and U23564 (N_23564,N_12588,N_15545);
or U23565 (N_23565,N_16289,N_19155);
nand U23566 (N_23566,N_15232,N_16932);
and U23567 (N_23567,N_15605,N_10150);
and U23568 (N_23568,N_16767,N_18339);
or U23569 (N_23569,N_10669,N_13050);
or U23570 (N_23570,N_12523,N_11639);
nor U23571 (N_23571,N_10475,N_12731);
nor U23572 (N_23572,N_13033,N_10737);
nor U23573 (N_23573,N_10864,N_16900);
nand U23574 (N_23574,N_14983,N_16472);
nand U23575 (N_23575,N_16079,N_16868);
nand U23576 (N_23576,N_17996,N_17020);
nand U23577 (N_23577,N_10997,N_12199);
or U23578 (N_23578,N_12355,N_13296);
or U23579 (N_23579,N_10722,N_16372);
xor U23580 (N_23580,N_11662,N_13992);
nor U23581 (N_23581,N_14740,N_17575);
or U23582 (N_23582,N_17873,N_13710);
and U23583 (N_23583,N_10402,N_13679);
and U23584 (N_23584,N_11777,N_19026);
nand U23585 (N_23585,N_16648,N_14538);
nor U23586 (N_23586,N_19553,N_15083);
and U23587 (N_23587,N_18145,N_12364);
or U23588 (N_23588,N_10522,N_11596);
or U23589 (N_23589,N_14849,N_12676);
and U23590 (N_23590,N_18722,N_18969);
or U23591 (N_23591,N_15583,N_15103);
and U23592 (N_23592,N_10621,N_10810);
nor U23593 (N_23593,N_16147,N_15860);
nand U23594 (N_23594,N_14656,N_17852);
nand U23595 (N_23595,N_19092,N_14709);
or U23596 (N_23596,N_19797,N_16141);
nor U23597 (N_23597,N_19261,N_12126);
or U23598 (N_23598,N_18545,N_18230);
nor U23599 (N_23599,N_15443,N_18172);
nor U23600 (N_23600,N_16702,N_14967);
nor U23601 (N_23601,N_13827,N_10571);
or U23602 (N_23602,N_15368,N_18214);
or U23603 (N_23603,N_10746,N_12477);
nand U23604 (N_23604,N_16021,N_10893);
or U23605 (N_23605,N_15593,N_12953);
or U23606 (N_23606,N_16886,N_12039);
nor U23607 (N_23607,N_18393,N_16260);
nand U23608 (N_23608,N_11266,N_13450);
or U23609 (N_23609,N_18494,N_12993);
or U23610 (N_23610,N_13939,N_14701);
and U23611 (N_23611,N_12102,N_13138);
or U23612 (N_23612,N_11398,N_13170);
or U23613 (N_23613,N_12266,N_11383);
nand U23614 (N_23614,N_15690,N_11860);
and U23615 (N_23615,N_18570,N_13072);
nor U23616 (N_23616,N_13221,N_19682);
or U23617 (N_23617,N_15424,N_17160);
and U23618 (N_23618,N_19407,N_15707);
nand U23619 (N_23619,N_10581,N_14567);
or U23620 (N_23620,N_17275,N_15844);
and U23621 (N_23621,N_15255,N_19801);
nand U23622 (N_23622,N_19885,N_15024);
nor U23623 (N_23623,N_19238,N_11544);
and U23624 (N_23624,N_14922,N_19333);
and U23625 (N_23625,N_10110,N_17912);
nor U23626 (N_23626,N_11052,N_11051);
nor U23627 (N_23627,N_13968,N_18370);
or U23628 (N_23628,N_16647,N_15108);
or U23629 (N_23629,N_11715,N_12611);
or U23630 (N_23630,N_16544,N_17364);
nand U23631 (N_23631,N_12612,N_18351);
nand U23632 (N_23632,N_12289,N_13533);
nor U23633 (N_23633,N_13682,N_16774);
or U23634 (N_23634,N_10425,N_15115);
or U23635 (N_23635,N_14771,N_16933);
and U23636 (N_23636,N_19850,N_11972);
nor U23637 (N_23637,N_11675,N_11568);
nor U23638 (N_23638,N_14279,N_11407);
and U23639 (N_23639,N_15694,N_10358);
or U23640 (N_23640,N_10264,N_18672);
and U23641 (N_23641,N_12581,N_10186);
nand U23642 (N_23642,N_15830,N_12302);
and U23643 (N_23643,N_12235,N_12190);
nor U23644 (N_23644,N_11389,N_16972);
or U23645 (N_23645,N_11470,N_17179);
nand U23646 (N_23646,N_13885,N_19050);
and U23647 (N_23647,N_13999,N_14980);
or U23648 (N_23648,N_11309,N_18948);
nor U23649 (N_23649,N_15275,N_12877);
nand U23650 (N_23650,N_14718,N_12785);
nand U23651 (N_23651,N_15382,N_11712);
or U23652 (N_23652,N_18843,N_17355);
nand U23653 (N_23653,N_13525,N_13996);
and U23654 (N_23654,N_14452,N_19611);
and U23655 (N_23655,N_18430,N_11803);
and U23656 (N_23656,N_19722,N_19338);
nand U23657 (N_23657,N_16870,N_18547);
and U23658 (N_23658,N_11384,N_16704);
nor U23659 (N_23659,N_18173,N_18811);
or U23660 (N_23660,N_11785,N_10210);
and U23661 (N_23661,N_12585,N_19421);
nor U23662 (N_23662,N_11862,N_18441);
or U23663 (N_23663,N_13563,N_18465);
and U23664 (N_23664,N_10118,N_14215);
nand U23665 (N_23665,N_12796,N_13929);
or U23666 (N_23666,N_15281,N_11294);
and U23667 (N_23667,N_17787,N_19329);
xor U23668 (N_23668,N_15350,N_10906);
or U23669 (N_23669,N_19334,N_14623);
or U23670 (N_23670,N_13338,N_12983);
and U23671 (N_23671,N_12016,N_19504);
or U23672 (N_23672,N_14450,N_15481);
nand U23673 (N_23673,N_18425,N_19454);
and U23674 (N_23674,N_11168,N_19384);
nand U23675 (N_23675,N_14179,N_17831);
or U23676 (N_23676,N_10404,N_17658);
or U23677 (N_23677,N_15279,N_16493);
and U23678 (N_23678,N_19010,N_12658);
or U23679 (N_23679,N_17692,N_13798);
nor U23680 (N_23680,N_11453,N_16777);
nor U23681 (N_23681,N_16729,N_10040);
or U23682 (N_23682,N_15142,N_14060);
or U23683 (N_23683,N_14869,N_15712);
nand U23684 (N_23684,N_10029,N_17893);
nor U23685 (N_23685,N_19472,N_15162);
or U23686 (N_23686,N_14541,N_10736);
nor U23687 (N_23687,N_17034,N_13004);
or U23688 (N_23688,N_18686,N_10246);
nor U23689 (N_23689,N_15124,N_12454);
and U23690 (N_23690,N_17402,N_12063);
nand U23691 (N_23691,N_12295,N_11896);
nand U23692 (N_23692,N_19347,N_10138);
or U23693 (N_23693,N_10612,N_11041);
xnor U23694 (N_23694,N_14557,N_13075);
nand U23695 (N_23695,N_14413,N_11565);
nand U23696 (N_23696,N_16446,N_16217);
or U23697 (N_23697,N_17134,N_13008);
nor U23698 (N_23698,N_11987,N_16319);
or U23699 (N_23699,N_18565,N_11989);
or U23700 (N_23700,N_15819,N_11134);
or U23701 (N_23701,N_16455,N_13231);
or U23702 (N_23702,N_13789,N_14575);
nand U23703 (N_23703,N_13214,N_16155);
or U23704 (N_23704,N_16703,N_15227);
nor U23705 (N_23705,N_19137,N_17415);
nor U23706 (N_23706,N_11829,N_14871);
nor U23707 (N_23707,N_12556,N_16509);
and U23708 (N_23708,N_18819,N_18432);
nand U23709 (N_23709,N_10951,N_10768);
nor U23710 (N_23710,N_16538,N_14671);
nor U23711 (N_23711,N_14328,N_12070);
and U23712 (N_23712,N_17667,N_17920);
and U23713 (N_23713,N_15816,N_14915);
or U23714 (N_23714,N_11555,N_19066);
nand U23715 (N_23715,N_18062,N_19315);
and U23716 (N_23716,N_13987,N_17358);
and U23717 (N_23717,N_11227,N_14475);
or U23718 (N_23718,N_13741,N_12508);
nand U23719 (N_23719,N_10664,N_12498);
and U23720 (N_23720,N_10950,N_11600);
and U23721 (N_23721,N_16685,N_13035);
nor U23722 (N_23722,N_15423,N_11026);
xor U23723 (N_23723,N_16974,N_13485);
and U23724 (N_23724,N_18972,N_14570);
nand U23725 (N_23725,N_12423,N_10012);
or U23726 (N_23726,N_14925,N_10394);
and U23727 (N_23727,N_10299,N_10990);
nor U23728 (N_23728,N_10432,N_10004);
nor U23729 (N_23729,N_10375,N_18721);
or U23730 (N_23730,N_12340,N_17188);
or U23731 (N_23731,N_19120,N_19202);
and U23732 (N_23732,N_18905,N_14050);
nand U23733 (N_23733,N_12169,N_18647);
nor U23734 (N_23734,N_13376,N_19661);
nand U23735 (N_23735,N_15549,N_18275);
nor U23736 (N_23736,N_10067,N_16216);
or U23737 (N_23737,N_15042,N_13385);
nand U23738 (N_23738,N_13317,N_10836);
or U23739 (N_23739,N_11773,N_10129);
nor U23740 (N_23740,N_15391,N_16858);
or U23741 (N_23741,N_12002,N_19128);
nor U23742 (N_23742,N_11735,N_14372);
nor U23743 (N_23743,N_15531,N_17162);
nor U23744 (N_23744,N_14783,N_17537);
nor U23745 (N_23745,N_14423,N_18043);
and U23746 (N_23746,N_10651,N_19124);
nand U23747 (N_23747,N_12316,N_16813);
and U23748 (N_23748,N_14865,N_18942);
or U23749 (N_23749,N_18225,N_13579);
nand U23750 (N_23750,N_12195,N_15256);
and U23751 (N_23751,N_15800,N_16884);
or U23752 (N_23752,N_16754,N_17665);
or U23753 (N_23753,N_13667,N_19538);
and U23754 (N_23754,N_18665,N_10003);
and U23755 (N_23755,N_18379,N_11558);
or U23756 (N_23756,N_13782,N_10282);
nand U23757 (N_23757,N_14533,N_19562);
nand U23758 (N_23758,N_11260,N_10963);
and U23759 (N_23759,N_11634,N_18118);
or U23760 (N_23760,N_15547,N_17673);
nand U23761 (N_23761,N_18615,N_10487);
and U23762 (N_23762,N_16968,N_11308);
or U23763 (N_23763,N_19810,N_12166);
and U23764 (N_23764,N_10478,N_14634);
and U23765 (N_23765,N_11535,N_16897);
xor U23766 (N_23766,N_10304,N_10201);
nor U23767 (N_23767,N_17105,N_11416);
and U23768 (N_23768,N_19629,N_19736);
or U23769 (N_23769,N_13418,N_11948);
or U23770 (N_23770,N_12808,N_17841);
or U23771 (N_23771,N_17674,N_17458);
or U23772 (N_23772,N_10377,N_11788);
or U23773 (N_23773,N_10077,N_19127);
and U23774 (N_23774,N_18273,N_16669);
and U23775 (N_23775,N_15242,N_16862);
nor U23776 (N_23776,N_19923,N_11095);
nor U23777 (N_23777,N_15001,N_12292);
and U23778 (N_23778,N_17738,N_18102);
or U23779 (N_23779,N_17279,N_12240);
or U23780 (N_23780,N_14710,N_18076);
nor U23781 (N_23781,N_10874,N_12468);
nor U23782 (N_23782,N_19537,N_12469);
or U23783 (N_23783,N_12507,N_16725);
nand U23784 (N_23784,N_17336,N_14116);
and U23785 (N_23785,N_16466,N_18296);
or U23786 (N_23786,N_12119,N_12542);
and U23787 (N_23787,N_14791,N_10481);
and U23788 (N_23788,N_14329,N_10724);
and U23789 (N_23789,N_11305,N_13439);
and U23790 (N_23790,N_15792,N_17997);
or U23791 (N_23791,N_11467,N_10388);
nor U23792 (N_23792,N_11280,N_18864);
nand U23793 (N_23793,N_19391,N_19709);
or U23794 (N_23794,N_14929,N_18460);
nand U23795 (N_23795,N_14627,N_13740);
or U23796 (N_23796,N_17773,N_19427);
nand U23797 (N_23797,N_15176,N_13100);
nand U23798 (N_23798,N_11683,N_11636);
nor U23799 (N_23799,N_13589,N_17444);
nor U23800 (N_23800,N_16149,N_14870);
and U23801 (N_23801,N_14494,N_16772);
nor U23802 (N_23802,N_10879,N_14918);
nand U23803 (N_23803,N_10865,N_10389);
or U23804 (N_23804,N_13310,N_14719);
nor U23805 (N_23805,N_17956,N_12516);
nor U23806 (N_23806,N_15629,N_19130);
nand U23807 (N_23807,N_11943,N_11694);
nor U23808 (N_23808,N_10564,N_11890);
nand U23809 (N_23809,N_16398,N_10366);
nand U23810 (N_23810,N_15445,N_15985);
and U23811 (N_23811,N_14876,N_16716);
nand U23812 (N_23812,N_10970,N_19475);
nand U23813 (N_23813,N_17993,N_12419);
nand U23814 (N_23814,N_18475,N_12149);
nand U23815 (N_23815,N_14247,N_12902);
nor U23816 (N_23816,N_18347,N_12944);
nor U23817 (N_23817,N_11046,N_13545);
nor U23818 (N_23818,N_16742,N_10142);
and U23819 (N_23819,N_11564,N_10613);
nand U23820 (N_23820,N_13268,N_11824);
and U23821 (N_23821,N_15174,N_14122);
nor U23822 (N_23822,N_12558,N_18089);
nor U23823 (N_23823,N_18507,N_12400);
nand U23824 (N_23824,N_11094,N_18416);
nor U23825 (N_23825,N_18667,N_16913);
xnor U23826 (N_23826,N_18603,N_17320);
nor U23827 (N_23827,N_11499,N_17317);
nor U23828 (N_23828,N_15049,N_12464);
nor U23829 (N_23829,N_13622,N_17911);
nand U23830 (N_23830,N_19032,N_18913);
and U23831 (N_23831,N_17221,N_18756);
or U23832 (N_23832,N_19178,N_10000);
or U23833 (N_23833,N_15523,N_18344);
or U23834 (N_23834,N_10610,N_15456);
nand U23835 (N_23835,N_18176,N_17385);
nand U23836 (N_23836,N_12888,N_14942);
and U23837 (N_23837,N_19025,N_11521);
nor U23838 (N_23838,N_18954,N_11420);
nand U23839 (N_23839,N_12403,N_15972);
nand U23840 (N_23840,N_10336,N_16594);
nand U23841 (N_23841,N_11915,N_11122);
nor U23842 (N_23842,N_13974,N_17830);
nand U23843 (N_23843,N_16143,N_16296);
nand U23844 (N_23844,N_10080,N_17454);
or U23845 (N_23845,N_19732,N_19038);
or U23846 (N_23846,N_18204,N_10093);
nand U23847 (N_23847,N_15278,N_16903);
nor U23848 (N_23848,N_13289,N_17480);
or U23849 (N_23849,N_19635,N_14548);
and U23850 (N_23850,N_19003,N_14829);
nand U23851 (N_23851,N_19992,N_11405);
nand U23852 (N_23852,N_16223,N_10682);
nand U23853 (N_23853,N_15201,N_16278);
nor U23854 (N_23854,N_18021,N_10947);
or U23855 (N_23855,N_19039,N_12371);
nor U23856 (N_23856,N_16104,N_11569);
or U23857 (N_23857,N_19135,N_13713);
or U23858 (N_23858,N_12904,N_18260);
nor U23859 (N_23859,N_18707,N_17745);
or U23860 (N_23860,N_16435,N_14572);
or U23861 (N_23861,N_15814,N_18742);
or U23862 (N_23862,N_12809,N_14262);
nand U23863 (N_23863,N_19159,N_12984);
and U23864 (N_23864,N_14327,N_19131);
and U23865 (N_23865,N_11524,N_15815);
nor U23866 (N_23866,N_11161,N_10804);
nor U23867 (N_23867,N_19378,N_11341);
or U23868 (N_23868,N_19316,N_16265);
nor U23869 (N_23869,N_10101,N_10155);
or U23870 (N_23870,N_14343,N_16636);
nand U23871 (N_23871,N_19395,N_15047);
nand U23872 (N_23872,N_11490,N_16635);
or U23873 (N_23873,N_15937,N_11087);
and U23874 (N_23874,N_18792,N_10857);
nor U23875 (N_23875,N_19716,N_16184);
xnor U23876 (N_23876,N_17688,N_11377);
nand U23877 (N_23877,N_13136,N_12420);
nor U23878 (N_23878,N_17182,N_16709);
or U23879 (N_23879,N_17989,N_19949);
or U23880 (N_23880,N_14863,N_15365);
and U23881 (N_23881,N_19359,N_11388);
nand U23882 (N_23882,N_17362,N_12829);
nand U23883 (N_23883,N_18977,N_17094);
nand U23884 (N_23884,N_16696,N_18500);
nand U23885 (N_23885,N_17574,N_15602);
and U23886 (N_23886,N_17907,N_14473);
nand U23887 (N_23887,N_17318,N_19110);
nor U23888 (N_23888,N_16333,N_10909);
or U23889 (N_23889,N_16088,N_11537);
nand U23890 (N_23890,N_18858,N_17763);
nand U23891 (N_23891,N_13860,N_11054);
or U23892 (N_23892,N_11531,N_12511);
xnor U23893 (N_23893,N_14319,N_11752);
nor U23894 (N_23894,N_11672,N_14440);
or U23895 (N_23895,N_10773,N_12801);
and U23896 (N_23896,N_15065,N_10991);
and U23897 (N_23897,N_15820,N_11487);
or U23898 (N_23898,N_15337,N_11240);
and U23899 (N_23899,N_19910,N_15979);
nor U23900 (N_23900,N_18485,N_12762);
nor U23901 (N_23901,N_11160,N_11802);
nand U23902 (N_23902,N_12318,N_15746);
nor U23903 (N_23903,N_14617,N_12899);
nor U23904 (N_23904,N_10514,N_14212);
or U23905 (N_23905,N_12052,N_15633);
nor U23906 (N_23906,N_11274,N_10307);
nand U23907 (N_23907,N_17850,N_16329);
nor U23908 (N_23908,N_18783,N_18131);
and U23909 (N_23909,N_17969,N_15548);
nor U23910 (N_23910,N_11918,N_13039);
nor U23911 (N_23911,N_16067,N_19394);
nor U23912 (N_23912,N_10787,N_11118);
nand U23913 (N_23913,N_17703,N_14539);
nand U23914 (N_23914,N_15446,N_15847);
or U23915 (N_23915,N_15246,N_11127);
or U23916 (N_23916,N_17715,N_13578);
and U23917 (N_23917,N_19835,N_11507);
or U23918 (N_23918,N_11967,N_15104);
and U23919 (N_23919,N_19275,N_18610);
nand U23920 (N_23920,N_15672,N_10035);
nand U23921 (N_23921,N_10771,N_17212);
nor U23922 (N_23922,N_10154,N_17490);
nand U23923 (N_23923,N_12301,N_17411);
or U23924 (N_23924,N_13791,N_10283);
nor U23925 (N_23925,N_14217,N_11501);
nand U23926 (N_23926,N_15818,N_12865);
or U23927 (N_23927,N_18663,N_11567);
nand U23928 (N_23928,N_17581,N_17495);
and U23929 (N_23929,N_10196,N_19088);
nor U23930 (N_23930,N_16743,N_15294);
nor U23931 (N_23931,N_19443,N_15987);
nand U23932 (N_23932,N_15771,N_12751);
or U23933 (N_23933,N_17578,N_12354);
nand U23934 (N_23934,N_14722,N_13910);
nor U23935 (N_23935,N_12326,N_18930);
nand U23936 (N_23936,N_12279,N_19062);
nor U23937 (N_23937,N_16530,N_18449);
nor U23938 (N_23938,N_10075,N_11724);
nor U23939 (N_23939,N_18324,N_17394);
or U23940 (N_23940,N_13177,N_12435);
or U23941 (N_23941,N_15692,N_15527);
nor U23942 (N_23942,N_15447,N_16848);
nand U23943 (N_23943,N_16921,N_19143);
nand U23944 (N_23944,N_13460,N_15831);
and U23945 (N_23945,N_14246,N_13938);
and U23946 (N_23946,N_17986,N_17400);
and U23947 (N_23947,N_11572,N_10631);
nor U23948 (N_23948,N_14674,N_15050);
and U23949 (N_23949,N_15347,N_19513);
nand U23950 (N_23950,N_14889,N_14596);
nor U23951 (N_23951,N_15383,N_15064);
and U23952 (N_23952,N_17820,N_14834);
or U23953 (N_23953,N_12082,N_18677);
or U23954 (N_23954,N_17296,N_14954);
and U23955 (N_23955,N_18939,N_16947);
nor U23956 (N_23956,N_15991,N_12513);
or U23957 (N_23957,N_12453,N_16573);
and U23958 (N_23958,N_19904,N_14135);
and U23959 (N_23959,N_13432,N_19790);
nand U23960 (N_23960,N_17876,N_19778);
nor U23961 (N_23961,N_15182,N_18413);
and U23962 (N_23962,N_14781,N_11107);
nor U23963 (N_23963,N_12574,N_11299);
and U23964 (N_23964,N_16888,N_14370);
nor U23965 (N_23965,N_17479,N_18943);
or U23966 (N_23966,N_18669,N_12047);
nor U23967 (N_23967,N_13131,N_19181);
nor U23968 (N_23968,N_14120,N_10943);
and U23969 (N_23969,N_19460,N_11105);
nand U23970 (N_23970,N_17946,N_18210);
nor U23971 (N_23971,N_14984,N_17804);
and U23972 (N_23972,N_18059,N_12929);
nand U23973 (N_23973,N_18323,N_13259);
or U23974 (N_23974,N_19247,N_18382);
nand U23975 (N_23975,N_19328,N_15643);
or U23976 (N_23976,N_12624,N_12883);
or U23977 (N_23977,N_15346,N_17901);
nor U23978 (N_23978,N_11279,N_14773);
nand U23979 (N_23979,N_18855,N_16752);
nor U23980 (N_23980,N_14768,N_11988);
nand U23981 (N_23981,N_10147,N_11976);
nor U23982 (N_23982,N_15912,N_10059);
nor U23983 (N_23983,N_16678,N_17597);
nand U23984 (N_23984,N_12594,N_18680);
and U23985 (N_23985,N_17433,N_15720);
and U23986 (N_23986,N_19502,N_12480);
and U23987 (N_23987,N_14320,N_14708);
nand U23988 (N_23988,N_14952,N_12737);
nor U23989 (N_23989,N_16590,N_11551);
nand U23990 (N_23990,N_13655,N_11312);
nor U23991 (N_23991,N_12986,N_15062);
nor U23992 (N_23992,N_14114,N_15373);
or U23993 (N_23993,N_14772,N_11358);
or U23994 (N_23994,N_13728,N_14019);
or U23995 (N_23995,N_17142,N_11343);
and U23996 (N_23996,N_10113,N_18763);
nand U23997 (N_23997,N_17104,N_11768);
nor U23998 (N_23998,N_14038,N_18436);
nor U23999 (N_23999,N_14132,N_11071);
nor U24000 (N_24000,N_10691,N_14410);
or U24001 (N_24001,N_15406,N_17129);
nor U24002 (N_24002,N_17447,N_15466);
and U24003 (N_24003,N_14908,N_13224);
nor U24004 (N_24004,N_10955,N_16003);
nor U24005 (N_24005,N_10912,N_10488);
nor U24006 (N_24006,N_16632,N_13402);
and U24007 (N_24007,N_16628,N_15728);
nand U24008 (N_24008,N_18631,N_13223);
nand U24009 (N_24009,N_11457,N_14356);
or U24010 (N_24010,N_16228,N_15817);
or U24011 (N_24011,N_14562,N_16950);
or U24012 (N_24012,N_15367,N_19405);
and U24013 (N_24013,N_15941,N_16365);
and U24014 (N_24014,N_12224,N_10648);
and U24015 (N_24015,N_19519,N_10137);
nor U24016 (N_24016,N_18019,N_18731);
and U24017 (N_24017,N_12262,N_10406);
nor U24018 (N_24018,N_15540,N_10082);
nor U24019 (N_24019,N_11643,N_12838);
nand U24020 (N_24020,N_15099,N_14643);
nand U24021 (N_24021,N_16118,N_14081);
or U24022 (N_24022,N_17580,N_13699);
or U24023 (N_24023,N_13928,N_13898);
or U24024 (N_24024,N_19283,N_11963);
and U24025 (N_24025,N_19272,N_14361);
and U24026 (N_24026,N_18034,N_10829);
nand U24027 (N_24027,N_14578,N_13983);
nand U24028 (N_24028,N_15997,N_19494);
and U24029 (N_24029,N_12798,N_11816);
and U24030 (N_24030,N_18814,N_16506);
nor U24031 (N_24031,N_19420,N_16070);
nor U24032 (N_24032,N_18480,N_17414);
nand U24033 (N_24033,N_11085,N_19539);
nand U24034 (N_24034,N_16295,N_16997);
or U24035 (N_24035,N_16063,N_18388);
and U24036 (N_24036,N_18947,N_11625);
nor U24037 (N_24037,N_12134,N_15966);
nor U24038 (N_24038,N_12707,N_15709);
or U24039 (N_24039,N_18805,N_13607);
and U24040 (N_24040,N_11737,N_18979);
and U24041 (N_24041,N_19035,N_15793);
or U24042 (N_24042,N_14891,N_16502);
and U24043 (N_24043,N_18373,N_12570);
or U24044 (N_24044,N_10254,N_19211);
and U24045 (N_24045,N_19152,N_12050);
xor U24046 (N_24046,N_12072,N_10856);
xnor U24047 (N_24047,N_13805,N_13905);
nand U24048 (N_24048,N_12288,N_16914);
or U24049 (N_24049,N_19617,N_10284);
nor U24050 (N_24050,N_16086,N_19742);
nor U24051 (N_24051,N_18238,N_13706);
nand U24052 (N_24052,N_14400,N_10062);
and U24053 (N_24053,N_10606,N_14943);
nand U24054 (N_24054,N_17334,N_19051);
nor U24055 (N_24055,N_12540,N_12839);
and U24056 (N_24056,N_14224,N_18291);
nand U24057 (N_24057,N_16341,N_13463);
nor U24058 (N_24058,N_18816,N_12576);
nand U24059 (N_24059,N_17795,N_16386);
nor U24060 (N_24060,N_17500,N_14691);
or U24061 (N_24061,N_10707,N_15805);
xnor U24062 (N_24062,N_19844,N_18269);
and U24063 (N_24063,N_16737,N_12639);
nor U24064 (N_24064,N_10508,N_11633);
nand U24065 (N_24065,N_10380,N_14495);
or U24066 (N_24066,N_18195,N_10988);
nand U24067 (N_24067,N_19912,N_12405);
nand U24068 (N_24068,N_15503,N_10410);
and U24069 (N_24069,N_16557,N_19812);
or U24070 (N_24070,N_15090,N_11426);
nand U24071 (N_24071,N_17862,N_17024);
and U24072 (N_24072,N_12666,N_15873);
nor U24073 (N_24073,N_10351,N_12763);
nor U24074 (N_24074,N_10723,N_12781);
nand U24075 (N_24075,N_13960,N_10405);
xor U24076 (N_24076,N_14236,N_11438);
and U24077 (N_24077,N_19118,N_17025);
xnor U24078 (N_24078,N_17159,N_16902);
nor U24079 (N_24079,N_10226,N_11895);
nor U24080 (N_24080,N_17933,N_18993);
or U24081 (N_24081,N_13634,N_16330);
and U24082 (N_24082,N_14181,N_13945);
xor U24083 (N_24083,N_18402,N_16229);
nor U24084 (N_24084,N_16934,N_10789);
nand U24085 (N_24085,N_17393,N_17583);
and U24086 (N_24086,N_15267,N_11586);
nand U24087 (N_24087,N_16061,N_10306);
nor U24088 (N_24088,N_18012,N_12934);
and U24089 (N_24089,N_15126,N_16040);
nand U24090 (N_24090,N_13235,N_13424);
or U24091 (N_24091,N_16713,N_10622);
nand U24092 (N_24092,N_19114,N_18978);
nand U24093 (N_24093,N_19235,N_19695);
nor U24094 (N_24094,N_16146,N_19503);
and U24095 (N_24095,N_13426,N_19757);
nand U24096 (N_24096,N_19374,N_17631);
and U24097 (N_24097,N_18708,N_19360);
nand U24098 (N_24098,N_17634,N_14170);
or U24099 (N_24099,N_17107,N_16403);
and U24100 (N_24100,N_18684,N_17043);
nand U24101 (N_24101,N_15286,N_11523);
and U24102 (N_24102,N_18660,N_14207);
or U24103 (N_24103,N_13542,N_13205);
nor U24104 (N_24104,N_14619,N_15093);
nand U24105 (N_24105,N_19511,N_12532);
and U24106 (N_24106,N_19655,N_17637);
and U24107 (N_24107,N_18606,N_17921);
and U24108 (N_24108,N_19849,N_10325);
and U24109 (N_24109,N_12483,N_18387);
nand U24110 (N_24110,N_15414,N_10466);
nor U24111 (N_24111,N_12722,N_19160);
and U24112 (N_24112,N_14080,N_18542);
and U24113 (N_24113,N_16959,N_10060);
nand U24114 (N_24114,N_12365,N_17112);
nor U24115 (N_24115,N_18248,N_17016);
or U24116 (N_24116,N_17582,N_18177);
and U24117 (N_24117,N_14161,N_14353);
nor U24118 (N_24118,N_18874,N_17606);
nor U24119 (N_24119,N_17732,N_12479);
nand U24120 (N_24120,N_16271,N_14079);
nand U24121 (N_24121,N_12151,N_19934);
and U24122 (N_24122,N_11620,N_18538);
and U24123 (N_24123,N_11935,N_16019);
nor U24124 (N_24124,N_12835,N_19896);
or U24125 (N_24125,N_12875,N_12248);
and U24126 (N_24126,N_16957,N_15829);
or U24127 (N_24127,N_17093,N_15098);
nor U24128 (N_24128,N_13092,N_18486);
and U24129 (N_24129,N_19729,N_14555);
nor U24130 (N_24130,N_15839,N_10543);
nand U24131 (N_24131,N_16300,N_15755);
xnor U24132 (N_24132,N_14363,N_19745);
nor U24133 (N_24133,N_10463,N_12293);
nand U24134 (N_24134,N_18807,N_10905);
nand U24135 (N_24135,N_17271,N_14063);
or U24136 (N_24136,N_17222,N_10733);
and U24137 (N_24137,N_14695,N_11884);
or U24138 (N_24138,N_19024,N_19067);
nand U24139 (N_24139,N_19796,N_14460);
or U24140 (N_24140,N_17309,N_11401);
nand U24141 (N_24141,N_15499,N_12807);
and U24142 (N_24142,N_15552,N_18501);
and U24143 (N_24143,N_15731,N_12592);
nor U24144 (N_24144,N_13094,N_13776);
nor U24145 (N_24145,N_19314,N_14790);
or U24146 (N_24146,N_19451,N_12648);
or U24147 (N_24147,N_13278,N_18511);
nor U24148 (N_24148,N_13899,N_15002);
nand U24149 (N_24149,N_17132,N_16188);
nand U24150 (N_24150,N_17088,N_10501);
and U24151 (N_24151,N_18725,N_16305);
and U24152 (N_24152,N_12146,N_16212);
or U24153 (N_24153,N_12615,N_16221);
nor U24154 (N_24154,N_14492,N_16508);
nor U24155 (N_24155,N_10038,N_12373);
and U24156 (N_24156,N_11808,N_16133);
nor U24157 (N_24157,N_17900,N_10749);
nor U24158 (N_24158,N_19928,N_15655);
nand U24159 (N_24159,N_12734,N_16112);
nor U24160 (N_24160,N_13901,N_15601);
nor U24161 (N_24161,N_15444,N_15244);
nor U24162 (N_24162,N_13116,N_11278);
and U24163 (N_24163,N_13984,N_11034);
and U24164 (N_24164,N_13007,N_14529);
and U24165 (N_24165,N_19318,N_16125);
or U24166 (N_24166,N_14712,N_13844);
and U24167 (N_24167,N_11887,N_18987);
nor U24168 (N_24168,N_12244,N_16318);
or U24169 (N_24169,N_14838,N_12931);
xnor U24170 (N_24170,N_10259,N_18693);
or U24171 (N_24171,N_13166,N_16836);
nor U24172 (N_24172,N_17533,N_13236);
nand U24173 (N_24173,N_11998,N_19373);
and U24174 (N_24174,N_13752,N_15184);
or U24175 (N_24175,N_14261,N_17737);
nor U24176 (N_24176,N_12870,N_18417);
and U24177 (N_24177,N_10546,N_16578);
nor U24178 (N_24178,N_19552,N_18562);
or U24179 (N_24179,N_18853,N_17084);
and U24180 (N_24180,N_19802,N_12417);
and U24181 (N_24181,N_19257,N_12563);
and U24182 (N_24182,N_16555,N_11901);
or U24183 (N_24183,N_10776,N_13203);
or U24184 (N_24184,N_13267,N_12945);
nand U24185 (N_24185,N_17008,N_16840);
nand U24186 (N_24186,N_18902,N_18363);
and U24187 (N_24187,N_16982,N_13613);
nand U24188 (N_24188,N_17306,N_12263);
or U24189 (N_24189,N_19210,N_11991);
nor U24190 (N_24190,N_16163,N_10796);
or U24191 (N_24191,N_10835,N_13276);
or U24192 (N_24192,N_17506,N_19192);
nand U24193 (N_24193,N_18697,N_11642);
and U24194 (N_24194,N_11251,N_11317);
or U24195 (N_24195,N_13118,N_19156);
and U24196 (N_24196,N_14653,N_17694);
nand U24197 (N_24197,N_15471,N_15705);
nand U24198 (N_24198,N_16953,N_12637);
or U24199 (N_24199,N_19289,N_18502);
and U24200 (N_24200,N_17722,N_17824);
nand U24201 (N_24201,N_13995,N_17126);
nor U24202 (N_24202,N_17754,N_11734);
nor U24203 (N_24203,N_14409,N_14216);
or U24204 (N_24204,N_17407,N_17620);
nand U24205 (N_24205,N_12264,N_11698);
nor U24206 (N_24206,N_18255,N_13069);
or U24207 (N_24207,N_17198,N_16024);
and U24208 (N_24208,N_12111,N_19133);
nand U24209 (N_24209,N_12065,N_17511);
nand U24210 (N_24210,N_13125,N_18591);
nor U24211 (N_24211,N_19811,N_14767);
nand U24212 (N_24212,N_13872,N_14485);
or U24213 (N_24213,N_13600,N_11344);
or U24214 (N_24214,N_12800,N_11674);
or U24215 (N_24215,N_15484,N_18179);
nor U24216 (N_24216,N_13343,N_15507);
or U24217 (N_24217,N_13472,N_13060);
or U24218 (N_24218,N_15428,N_11155);
nor U24219 (N_24219,N_10411,N_10719);
nor U24220 (N_24220,N_12025,N_12180);
nor U24221 (N_24221,N_16290,N_12705);
nand U24222 (N_24222,N_18085,N_10232);
nor U24223 (N_24223,N_15390,N_14406);
and U24224 (N_24224,N_10435,N_10450);
nand U24225 (N_24225,N_19761,N_11759);
and U24226 (N_24226,N_13927,N_15122);
and U24227 (N_24227,N_10251,N_11632);
and U24228 (N_24228,N_15165,N_13819);
nand U24229 (N_24229,N_15040,N_19171);
or U24230 (N_24230,N_16756,N_16825);
nor U24231 (N_24231,N_15435,N_14291);
nor U24232 (N_24232,N_17924,N_16038);
and U24233 (N_24233,N_18241,N_12294);
nor U24234 (N_24234,N_10588,N_14260);
or U24235 (N_24235,N_16824,N_16679);
or U24236 (N_24236,N_19147,N_19683);
and U24237 (N_24237,N_17651,N_10335);
nor U24238 (N_24238,N_19587,N_17404);
nand U24239 (N_24239,N_13853,N_18527);
or U24240 (N_24240,N_17098,N_19335);
nand U24241 (N_24241,N_10428,N_11570);
nor U24242 (N_24242,N_13346,N_15614);
nor U24243 (N_24243,N_11114,N_15271);
nand U24244 (N_24244,N_10780,N_18042);
or U24245 (N_24245,N_15813,N_10662);
and U24246 (N_24246,N_18870,N_16942);
or U24247 (N_24247,N_16301,N_16145);
or U24248 (N_24248,N_11673,N_19365);
and U24249 (N_24249,N_13301,N_17867);
or U24250 (N_24250,N_18568,N_10932);
nor U24251 (N_24251,N_12690,N_10169);
or U24252 (N_24252,N_11411,N_14753);
or U24253 (N_24253,N_11258,N_19020);
or U24254 (N_24254,N_16039,N_11496);
nand U24255 (N_24255,N_12708,N_12430);
nand U24256 (N_24256,N_12547,N_17653);
and U24257 (N_24257,N_10261,N_15171);
and U24258 (N_24258,N_14510,N_16951);
and U24259 (N_24259,N_12771,N_15668);
and U24260 (N_24260,N_14630,N_19671);
or U24261 (N_24261,N_10711,N_13102);
nor U24262 (N_24262,N_11577,N_19064);
nor U24263 (N_24263,N_11622,N_16092);
or U24264 (N_24264,N_14313,N_18083);
nor U24265 (N_24265,N_15574,N_17848);
or U24266 (N_24266,N_18251,N_13328);
nand U24267 (N_24267,N_15086,N_16621);
nor U24268 (N_24268,N_10873,N_18555);
nand U24269 (N_24269,N_14330,N_16344);
xnor U24270 (N_24270,N_11716,N_13551);
nand U24271 (N_24271,N_12622,N_14160);
and U24272 (N_24272,N_13725,N_13997);
nor U24273 (N_24273,N_19381,N_19097);
nand U24274 (N_24274,N_11232,N_13178);
nor U24275 (N_24275,N_11923,N_13738);
nor U24276 (N_24276,N_16043,N_14757);
or U24277 (N_24277,N_13906,N_11990);
nor U24278 (N_24278,N_12655,N_13539);
and U24279 (N_24279,N_13444,N_16652);
nand U24280 (N_24280,N_10217,N_17350);
nand U24281 (N_24281,N_15394,N_13132);
nand U24282 (N_24282,N_14082,N_10291);
or U24283 (N_24283,N_10639,N_16089);
nor U24284 (N_24284,N_19173,N_15904);
nand U24285 (N_24285,N_19326,N_13281);
nand U24286 (N_24286,N_11465,N_15432);
nor U24287 (N_24287,N_12164,N_13332);
xnor U24288 (N_24288,N_19057,N_13397);
nand U24289 (N_24289,N_10820,N_17682);
nor U24290 (N_24290,N_12450,N_14676);
and U24291 (N_24291,N_10321,N_13873);
and U24292 (N_24292,N_13059,N_10848);
and U24293 (N_24293,N_17710,N_12218);
and U24294 (N_24294,N_10574,N_16492);
and U24295 (N_24295,N_18552,N_17004);
and U24296 (N_24296,N_13765,N_18153);
nor U24297 (N_24297,N_18898,N_18207);
and U24298 (N_24298,N_16761,N_14020);
and U24299 (N_24299,N_17005,N_10530);
nand U24300 (N_24300,N_16321,N_10292);
or U24301 (N_24301,N_15875,N_12812);
and U24302 (N_24302,N_19901,N_19348);
nor U24303 (N_24303,N_10775,N_17982);
or U24304 (N_24304,N_15170,N_18438);
or U24305 (N_24305,N_14001,N_18757);
nor U24306 (N_24306,N_14655,N_18620);
and U24307 (N_24307,N_13209,N_19255);
nor U24308 (N_24308,N_14153,N_12078);
and U24309 (N_24309,N_17567,N_13640);
or U24310 (N_24310,N_11582,N_15778);
nor U24311 (N_24311,N_12455,N_11395);
nand U24312 (N_24312,N_17655,N_18411);
and U24313 (N_24313,N_17277,N_19430);
or U24314 (N_24314,N_15335,N_12457);
nor U24315 (N_24315,N_19911,N_14907);
nor U24316 (N_24316,N_10505,N_18714);
or U24317 (N_24317,N_13534,N_14476);
or U24318 (N_24318,N_12901,N_12546);
xor U24319 (N_24319,N_18151,N_11846);
nand U24320 (N_24320,N_10057,N_12779);
or U24321 (N_24321,N_11480,N_13981);
or U24322 (N_24322,N_16203,N_16891);
and U24323 (N_24323,N_17851,N_14051);
nand U24324 (N_24324,N_13908,N_14941);
nand U24325 (N_24325,N_17771,N_12441);
or U24326 (N_24326,N_10369,N_15592);
nor U24327 (N_24327,N_14470,N_19955);
and U24328 (N_24328,N_12837,N_15770);
nor U24329 (N_24329,N_11583,N_16513);
and U24330 (N_24330,N_11250,N_10106);
or U24331 (N_24331,N_19491,N_12833);
and U24332 (N_24332,N_17238,N_17463);
or U24333 (N_24333,N_13653,N_11806);
and U24334 (N_24334,N_19837,N_17635);
and U24335 (N_24335,N_19492,N_16946);
and U24336 (N_24336,N_12493,N_11145);
and U24337 (N_24337,N_14390,N_15375);
nor U24338 (N_24338,N_19759,N_13297);
nand U24339 (N_24339,N_18762,N_19874);
nand U24340 (N_24340,N_16078,N_10164);
nor U24341 (N_24341,N_19437,N_18878);
and U24342 (N_24342,N_15963,N_19748);
nor U24343 (N_24343,N_18696,N_18078);
or U24344 (N_24344,N_19895,N_16342);
and U24345 (N_24345,N_13572,N_10531);
nor U24346 (N_24346,N_19132,N_10034);
nand U24347 (N_24347,N_18121,N_18678);
or U24348 (N_24348,N_16136,N_14697);
or U24349 (N_24349,N_10832,N_18512);
nand U24350 (N_24350,N_14169,N_19705);
or U24351 (N_24351,N_11045,N_19744);
or U24352 (N_24352,N_12084,N_19679);
and U24353 (N_24353,N_10728,N_14956);
nor U24354 (N_24354,N_12174,N_16757);
nor U24355 (N_24355,N_18991,N_19191);
or U24356 (N_24356,N_13677,N_19631);
and U24357 (N_24357,N_13802,N_17267);
or U24358 (N_24358,N_14394,N_10941);
or U24359 (N_24359,N_12444,N_16140);
nor U24360 (N_24360,N_17889,N_10148);
nor U24361 (N_24361,N_16178,N_14949);
nor U24362 (N_24362,N_16983,N_13315);
nand U24363 (N_24363,N_13389,N_13510);
and U24364 (N_24364,N_14986,N_19089);
nand U24365 (N_24365,N_18077,N_12179);
and U24366 (N_24366,N_19262,N_19022);
or U24367 (N_24367,N_19989,N_11014);
and U24368 (N_24368,N_17015,N_17786);
nand U24369 (N_24369,N_18073,N_17770);
nor U24370 (N_24370,N_19458,N_10078);
nand U24371 (N_24371,N_19696,N_11130);
nor U24372 (N_24372,N_18237,N_17227);
or U24373 (N_24373,N_11249,N_14429);
and U24374 (N_24374,N_15785,N_14810);
and U24375 (N_24375,N_10277,N_11619);
nor U24376 (N_24376,N_11811,N_11519);
and U24377 (N_24377,N_14096,N_11522);
or U24378 (N_24378,N_11807,N_14240);
or U24379 (N_24379,N_13459,N_12484);
nor U24380 (N_24380,N_15429,N_11113);
or U24381 (N_24381,N_16432,N_14322);
nor U24382 (N_24382,N_14016,N_10614);
nand U24383 (N_24383,N_14415,N_13627);
or U24384 (N_24384,N_12618,N_18560);
and U24385 (N_24385,N_17811,N_16379);
or U24386 (N_24386,N_19331,N_19054);
nor U24387 (N_24387,N_14583,N_18127);
nand U24388 (N_24388,N_10334,N_14906);
nand U24389 (N_24389,N_18469,N_10092);
or U24390 (N_24390,N_19795,N_14252);
nand U24391 (N_24391,N_10384,N_19979);
and U24392 (N_24392,N_12593,N_18768);
and U24393 (N_24393,N_13486,N_15434);
or U24394 (N_24394,N_10989,N_19274);
nand U24395 (N_24395,N_19983,N_10638);
and U24396 (N_24396,N_19279,N_12617);
nor U24397 (N_24397,N_18474,N_19560);
and U24398 (N_24398,N_17136,N_13474);
or U24399 (N_24399,N_12188,N_13337);
xnor U24400 (N_24400,N_16604,N_12210);
nand U24401 (N_24401,N_11171,N_15289);
nor U24402 (N_24402,N_14044,N_16399);
nor U24403 (N_24403,N_11154,N_10747);
nand U24404 (N_24404,N_13207,N_16778);
or U24405 (N_24405,N_16210,N_13838);
nor U24406 (N_24406,N_17069,N_16514);
nand U24407 (N_24407,N_18456,N_15578);
nand U24408 (N_24408,N_12907,N_16423);
and U24409 (N_24409,N_11243,N_10107);
nor U24410 (N_24410,N_16476,N_13036);
nor U24411 (N_24411,N_10689,N_11905);
nand U24412 (N_24412,N_18812,N_14602);
nor U24413 (N_24413,N_14958,N_14521);
and U24414 (N_24414,N_13168,N_17437);
or U24415 (N_24415,N_11914,N_17241);
and U24416 (N_24416,N_10212,N_12099);
or U24417 (N_24417,N_11969,N_11530);
or U24418 (N_24418,N_15569,N_14393);
nor U24419 (N_24419,N_11022,N_16864);
and U24420 (N_24420,N_17171,N_15889);
or U24421 (N_24421,N_16045,N_17883);
and U24422 (N_24422,N_15553,N_18980);
nor U24423 (N_24423,N_16410,N_12329);
or U24424 (N_24424,N_10248,N_19938);
nor U24425 (N_24425,N_14151,N_17965);
and U24426 (N_24426,N_12392,N_14457);
nor U24427 (N_24427,N_14817,N_13788);
and U24428 (N_24428,N_13169,N_15410);
nand U24429 (N_24429,N_13457,N_10486);
and U24430 (N_24430,N_16160,N_16082);
or U24431 (N_24431,N_13561,N_16909);
nand U24432 (N_24432,N_10806,N_13523);
nor U24433 (N_24433,N_18639,N_11677);
or U24434 (N_24434,N_16247,N_16780);
nand U24435 (N_24435,N_17727,N_14481);
or U24436 (N_24436,N_12770,N_14820);
or U24437 (N_24437,N_12754,N_18497);
and U24438 (N_24438,N_11021,N_11710);
or U24439 (N_24439,N_16992,N_14316);
nand U24440 (N_24440,N_17902,N_15020);
or U24441 (N_24441,N_13491,N_14245);
nand U24442 (N_24442,N_16730,N_17898);
nand U24443 (N_24443,N_10006,N_11186);
nand U24444 (N_24444,N_19340,N_13211);
and U24445 (N_24445,N_12439,N_18266);
nand U24446 (N_24446,N_15877,N_13808);
or U24447 (N_24447,N_10566,N_16409);
nand U24448 (N_24448,N_10136,N_16065);
nor U24449 (N_24449,N_15495,N_19741);
and U24450 (N_24450,N_13196,N_19672);
or U24451 (N_24451,N_12730,N_15970);
nor U24452 (N_24452,N_17515,N_14576);
or U24453 (N_24453,N_12806,N_10168);
nand U24454 (N_24454,N_16069,N_11136);
and U24455 (N_24455,N_15133,N_13473);
or U24456 (N_24456,N_10732,N_17462);
or U24457 (N_24457,N_12619,N_17118);
and U24458 (N_24458,N_13191,N_10643);
nand U24459 (N_24459,N_18886,N_13540);
and U24460 (N_24460,N_15542,N_12456);
nor U24461 (N_24461,N_14315,N_19833);
or U24462 (N_24462,N_17072,N_13183);
nor U24463 (N_24463,N_13900,N_14950);
and U24464 (N_24464,N_16571,N_13134);
nor U24465 (N_24465,N_18219,N_12331);
nand U24466 (N_24466,N_10686,N_15388);
and U24467 (N_24467,N_15405,N_16965);
nor U24468 (N_24468,N_16164,N_17497);
or U24469 (N_24469,N_12935,N_19848);
or U24470 (N_24470,N_12764,N_13287);
and U24471 (N_24471,N_13678,N_10995);
nor U24472 (N_24472,N_14366,N_18984);
or U24473 (N_24473,N_18928,N_15783);
or U24474 (N_24474,N_12332,N_13308);
nand U24475 (N_24475,N_16390,N_18923);
or U24476 (N_24476,N_13482,N_18473);
nand U24477 (N_24477,N_11111,N_10345);
nor U24478 (N_24478,N_16842,N_12684);
nor U24479 (N_24479,N_12504,N_18952);
nand U24480 (N_24480,N_16979,N_10987);
nor U24481 (N_24481,N_14565,N_16489);
and U24482 (N_24482,N_17185,N_16512);
nor U24483 (N_24483,N_17614,N_10593);
nor U24484 (N_24484,N_19376,N_14362);
nand U24485 (N_24485,N_17494,N_18906);
or U24486 (N_24486,N_11799,N_10326);
nand U24487 (N_24487,N_17483,N_16363);
and U24488 (N_24488,N_19145,N_17117);
or U24489 (N_24489,N_17847,N_17250);
and U24490 (N_24490,N_14553,N_15754);
and U24491 (N_24491,N_13772,N_19253);
nor U24492 (N_24492,N_14603,N_19725);
and U24493 (N_24493,N_17083,N_18967);
nor U24494 (N_24494,N_13455,N_12492);
nor U24495 (N_24495,N_12251,N_10533);
nand U24496 (N_24496,N_15576,N_16721);
or U24497 (N_24497,N_16717,N_15247);
and U24498 (N_24498,N_12759,N_17748);
or U24499 (N_24499,N_11277,N_14998);
nand U24500 (N_24500,N_18883,N_14919);
nand U24501 (N_24501,N_10609,N_10993);
nand U24502 (N_24502,N_10200,N_15136);
nand U24503 (N_24503,N_16952,N_11714);
nor U24504 (N_24504,N_17808,N_13702);
and U24505 (N_24505,N_14013,N_10794);
nor U24506 (N_24506,N_18014,N_17832);
nand U24507 (N_24507,N_16477,N_19531);
and U24508 (N_24508,N_10436,N_17849);
nor U24509 (N_24509,N_15726,N_12606);
nor U24510 (N_24510,N_15035,N_14446);
nand U24511 (N_24511,N_18925,N_11346);
nand U24512 (N_24512,N_11460,N_14077);
nor U24513 (N_24513,N_12094,N_13265);
nand U24514 (N_24514,N_16224,N_13674);
or U24515 (N_24515,N_16369,N_15430);
or U24516 (N_24516,N_12687,N_14574);
nand U24517 (N_24517,N_16397,N_18331);
and U24518 (N_24518,N_13724,N_19773);
xnor U24519 (N_24519,N_18405,N_12055);
nand U24520 (N_24520,N_12872,N_11826);
nor U24521 (N_24521,N_19876,N_11215);
xor U24522 (N_24522,N_10446,N_10122);
nand U24523 (N_24523,N_15312,N_19781);
nor U24524 (N_24524,N_15537,N_12256);
and U24525 (N_24525,N_17705,N_10949);
or U24526 (N_24526,N_16309,N_14844);
or U24527 (N_24527,N_19604,N_11707);
nand U24528 (N_24528,N_10134,N_13478);
and U24529 (N_24529,N_14682,N_17555);
or U24530 (N_24530,N_17455,N_10418);
nand U24531 (N_24531,N_12715,N_10073);
or U24532 (N_24532,N_18199,N_13870);
nand U24533 (N_24533,N_16784,N_19681);
nand U24534 (N_24534,N_11042,N_19248);
and U24535 (N_24535,N_16481,N_15028);
or U24536 (N_24536,N_19249,N_14095);
or U24537 (N_24537,N_17552,N_18028);
nor U24538 (N_24538,N_18583,N_10858);
or U24539 (N_24539,N_11733,N_19597);
or U24540 (N_24540,N_16852,N_12139);
nor U24541 (N_24541,N_16048,N_19301);
and U24542 (N_24542,N_17548,N_14402);
or U24543 (N_24543,N_14241,N_11375);
or U24544 (N_24544,N_12794,N_16266);
and U24545 (N_24545,N_15280,N_15120);
and U24546 (N_24546,N_19787,N_13321);
nor U24547 (N_24547,N_11271,N_11601);
nand U24548 (N_24548,N_15263,N_13396);
nand U24549 (N_24549,N_14803,N_11781);
nor U24550 (N_24550,N_15497,N_15412);
and U24551 (N_24551,N_14782,N_13962);
and U24552 (N_24552,N_12129,N_15930);
or U24553 (N_24553,N_17928,N_17550);
or U24554 (N_24554,N_13412,N_17747);
or U24555 (N_24555,N_16708,N_15735);
nand U24556 (N_24556,N_16645,N_10809);
or U24557 (N_24557,N_10416,N_11208);
nand U24558 (N_24558,N_16547,N_14201);
or U24559 (N_24559,N_18194,N_15745);
and U24560 (N_24560,N_17888,N_14100);
nor U24561 (N_24561,N_14624,N_14234);
nor U24562 (N_24562,N_12820,N_19017);
nor U24563 (N_24563,N_11628,N_10668);
xor U24564 (N_24564,N_17442,N_19227);
and U24565 (N_24565,N_15541,N_16973);
nand U24566 (N_24566,N_12878,N_10913);
nor U24567 (N_24567,N_15010,N_14748);
nand U24568 (N_24568,N_11960,N_14142);
nor U24569 (N_24569,N_10828,N_19113);
nor U24570 (N_24570,N_14993,N_11163);
xnor U24571 (N_24571,N_12245,N_18970);
and U24572 (N_24572,N_12549,N_13821);
or U24573 (N_24573,N_16139,N_10549);
nor U24574 (N_24574,N_10189,N_18026);
or U24575 (N_24575,N_18217,N_14503);
and U24576 (N_24576,N_15833,N_18048);
and U24577 (N_24577,N_17974,N_12628);
or U24578 (N_24578,N_18196,N_13201);
and U24579 (N_24579,N_14822,N_10575);
nor U24580 (N_24580,N_15015,N_14474);
and U24581 (N_24581,N_19306,N_11908);
xnor U24582 (N_24582,N_13800,N_14391);
nor U24583 (N_24583,N_17244,N_10850);
or U24584 (N_24584,N_14278,N_10161);
nor U24585 (N_24585,N_16474,N_15189);
and U24586 (N_24586,N_10713,N_12768);
or U24587 (N_24587,N_12854,N_10511);
or U24588 (N_24588,N_18482,N_12227);
and U24589 (N_24589,N_18290,N_11872);
or U24590 (N_24590,N_12587,N_19803);
nand U24591 (N_24591,N_16991,N_17342);
nor U24592 (N_24592,N_14836,N_19870);
and U24593 (N_24593,N_19467,N_13097);
or U24594 (N_24594,N_11612,N_14523);
nand U24595 (N_24595,N_16659,N_16497);
and U24596 (N_24596,N_19625,N_16677);
or U24597 (N_24597,N_11931,N_11129);
nor U24598 (N_24598,N_14365,N_13351);
and U24599 (N_24599,N_13158,N_11449);
or U24600 (N_24600,N_16162,N_18226);
and U24601 (N_24601,N_19528,N_15007);
or U24602 (N_24602,N_19041,N_10880);
nand U24603 (N_24603,N_16241,N_10548);
or U24604 (N_24604,N_16745,N_17781);
and U24605 (N_24605,N_10158,N_11765);
or U24606 (N_24606,N_14508,N_17879);
nand U24607 (N_24607,N_19939,N_11554);
or U24608 (N_24608,N_16121,N_16855);
and U24609 (N_24609,N_18205,N_18397);
and U24610 (N_24610,N_17622,N_12884);
or U24611 (N_24611,N_15217,N_10894);
nor U24612 (N_24612,N_18712,N_10181);
nor U24613 (N_24613,N_12660,N_18576);
nand U24614 (N_24614,N_13020,N_15993);
or U24615 (N_24615,N_19976,N_12345);
nor U24616 (N_24616,N_15665,N_17149);
or U24617 (N_24617,N_17647,N_12862);
and U24618 (N_24618,N_13325,N_14303);
nand U24619 (N_24619,N_12491,N_15521);
and U24620 (N_24620,N_13705,N_14148);
nor U24621 (N_24621,N_13722,N_14143);
or U24622 (N_24622,N_18271,N_10401);
and U24623 (N_24623,N_15881,N_12087);
nand U24624 (N_24624,N_12814,N_10623);
or U24625 (N_24625,N_14482,N_14796);
nand U24626 (N_24626,N_13406,N_11509);
or U24627 (N_24627,N_11618,N_11397);
or U24628 (N_24628,N_17082,N_11267);
nand U24629 (N_24629,N_18072,N_13966);
and U24630 (N_24630,N_19501,N_17992);
or U24631 (N_24631,N_16606,N_17208);
or U24632 (N_24632,N_13990,N_18551);
nand U24633 (N_24633,N_16308,N_12172);
and U24634 (N_24634,N_16135,N_11316);
or U24635 (N_24635,N_18148,N_18976);
or U24636 (N_24636,N_14537,N_18838);
or U24637 (N_24637,N_11177,N_19866);
and U24638 (N_24638,N_16046,N_17339);
nor U24639 (N_24639,N_17272,N_12905);
nand U24640 (N_24640,N_10338,N_10984);
nor U24641 (N_24641,N_10781,N_15211);
nand U24642 (N_24642,N_17124,N_18645);
and U24643 (N_24643,N_16174,N_19364);
and U24644 (N_24644,N_11515,N_16927);
nand U24645 (N_24645,N_12515,N_10556);
nor U24646 (N_24646,N_14657,N_16115);
nand U24647 (N_24647,N_17522,N_16758);
nor U24648 (N_24648,N_15842,N_12649);
and U24649 (N_24649,N_14219,N_17397);
nand U24650 (N_24650,N_19281,N_13694);
nor U24651 (N_24651,N_14506,N_14297);
nand U24652 (N_24652,N_15046,N_16823);
nand U24653 (N_24653,N_12046,N_18000);
or U24654 (N_24654,N_14648,N_10815);
nor U24655 (N_24655,N_12333,N_14905);
and U24656 (N_24656,N_17423,N_17668);
and U24657 (N_24657,N_18061,N_17457);
nor U24658 (N_24658,N_15241,N_17146);
nor U24659 (N_24659,N_14439,N_15292);
nor U24660 (N_24660,N_18738,N_16719);
or U24661 (N_24661,N_12776,N_10309);
nand U24662 (N_24662,N_19950,N_15393);
and U24663 (N_24663,N_17736,N_19439);
nor U24664 (N_24664,N_19958,N_14606);
nor U24665 (N_24665,N_12182,N_10807);
nand U24666 (N_24666,N_18047,N_16689);
nor U24667 (N_24667,N_17135,N_16619);
or U24668 (N_24668,N_18365,N_17675);
or U24669 (N_24669,N_10762,N_10476);
or U24670 (N_24670,N_10330,N_16734);
and U24671 (N_24671,N_10152,N_13449);
nor U24672 (N_24672,N_15221,N_10817);
or U24673 (N_24673,N_10799,N_11881);
nor U24674 (N_24674,N_19299,N_15681);
nand U24675 (N_24675,N_18215,N_10525);
nor U24676 (N_24676,N_18931,N_17603);
and U24677 (N_24677,N_11132,N_14725);
or U24678 (N_24678,N_11516,N_10310);
nor U24679 (N_24679,N_15529,N_10837);
and U24680 (N_24680,N_14552,N_13759);
and U24681 (N_24681,N_16199,N_11024);
or U24682 (N_24682,N_19157,N_17491);
and U24683 (N_24683,N_17408,N_14408);
or U24684 (N_24684,N_10091,N_15688);
nand U24685 (N_24685,N_17312,N_12482);
nand U24686 (N_24686,N_19791,N_12987);
nor U24687 (N_24687,N_13524,N_10591);
nand U24688 (N_24688,N_18752,N_13107);
and U24689 (N_24689,N_13358,N_13829);
or U24690 (N_24690,N_17384,N_11857);
and U24691 (N_24691,N_13820,N_15116);
or U24692 (N_24692,N_10538,N_18139);
or U24693 (N_24693,N_16415,N_14015);
or U24694 (N_24694,N_17307,N_10962);
nand U24695 (N_24695,N_15379,N_13340);
nor U24696 (N_24696,N_18920,N_14210);
nor U24697 (N_24697,N_16346,N_10399);
and U24698 (N_24698,N_17556,N_10465);
and U24699 (N_24699,N_11627,N_17170);
or U24700 (N_24700,N_17764,N_13193);
nand U24701 (N_24701,N_11894,N_14026);
or U24702 (N_24702,N_18412,N_14893);
and U24703 (N_24703,N_10275,N_16193);
nand U24704 (N_24704,N_18988,N_16646);
nand U24705 (N_24705,N_13692,N_18798);
nand U24706 (N_24706,N_16733,N_18174);
nor U24707 (N_24707,N_11563,N_17314);
nand U24708 (N_24708,N_14965,N_18820);
nor U24709 (N_24709,N_11849,N_18531);
nor U24710 (N_24710,N_16537,N_13669);
and U24711 (N_24711,N_11039,N_16254);
and U24712 (N_24712,N_16424,N_13777);
nor U24713 (N_24713,N_11753,N_19883);
nor U24714 (N_24714,N_13811,N_19633);
or U24715 (N_24715,N_13687,N_10419);
nand U24716 (N_24716,N_16425,N_15237);
or U24717 (N_24717,N_19337,N_16126);
nand U24718 (N_24718,N_10238,N_16267);
nand U24719 (N_24719,N_11728,N_12567);
or U24720 (N_24720,N_14447,N_10229);
or U24721 (N_24721,N_18766,N_15562);
nand U24722 (N_24722,N_16894,N_13869);
and U24723 (N_24723,N_11560,N_11656);
and U24724 (N_24724,N_19693,N_16880);
nand U24725 (N_24725,N_17712,N_11246);
or U24726 (N_24726,N_16440,N_15702);
and U24727 (N_24727,N_13189,N_16012);
or U24728 (N_24728,N_12161,N_18392);
nor U24729 (N_24729,N_13115,N_13566);
nand U24730 (N_24730,N_11798,N_19723);
and U24731 (N_24731,N_12891,N_15802);
and U24732 (N_24732,N_15186,N_17984);
nor U24733 (N_24733,N_12194,N_15648);
nor U24734 (N_24734,N_18443,N_12551);
nor U24735 (N_24735,N_17332,N_13895);
nand U24736 (N_24736,N_10030,N_15784);
nor U24737 (N_24737,N_12791,N_17940);
and U24738 (N_24738,N_19111,N_15215);
nor U24739 (N_24739,N_10971,N_17470);
nor U24740 (N_24740,N_15603,N_17040);
nand U24741 (N_24741,N_14295,N_14364);
nand U24742 (N_24742,N_16929,N_13230);
or U24743 (N_24743,N_12140,N_10756);
or U24744 (N_24744,N_13139,N_10816);
or U24745 (N_24745,N_15331,N_15300);
or U24746 (N_24746,N_16438,N_18578);
or U24747 (N_24747,N_19448,N_16005);
nand U24748 (N_24748,N_19200,N_10020);
nand U24749 (N_24749,N_11842,N_13386);
nand U24750 (N_24750,N_14211,N_14607);
nand U24751 (N_24751,N_17356,N_14765);
or U24752 (N_24752,N_11298,N_11471);
and U24753 (N_24753,N_16529,N_19404);
and U24754 (N_24754,N_14971,N_15016);
and U24755 (N_24755,N_18023,N_16747);
or U24756 (N_24756,N_16002,N_10529);
and U24757 (N_24757,N_11610,N_12353);
or U24758 (N_24758,N_18069,N_18130);
or U24759 (N_24759,N_13344,N_16055);
nor U24760 (N_24760,N_14289,N_15863);
and U24761 (N_24761,N_19596,N_14981);
nand U24762 (N_24762,N_16310,N_14660);
nand U24763 (N_24763,N_14352,N_15193);
and U24764 (N_24764,N_16427,N_15862);
and U24765 (N_24765,N_10449,N_15538);
nand U24766 (N_24766,N_15213,N_15297);
or U24767 (N_24767,N_15252,N_11541);
nor U24768 (N_24768,N_15738,N_19772);
or U24769 (N_24769,N_10604,N_18314);
nor U24770 (N_24770,N_13967,N_15338);
xnor U24771 (N_24771,N_16036,N_12537);
and U24772 (N_24772,N_14126,N_13247);
nand U24773 (N_24773,N_17731,N_17566);
nor U24774 (N_24774,N_12729,N_17958);
or U24775 (N_24775,N_10853,N_17930);
nor U24776 (N_24776,N_16016,N_11815);
and U24777 (N_24777,N_18659,N_14073);
or U24778 (N_24778,N_11711,N_13309);
nor U24779 (N_24779,N_11696,N_10956);
and U24780 (N_24780,N_17264,N_18124);
or U24781 (N_24781,N_10415,N_13649);
nand U24782 (N_24782,N_15959,N_10225);
or U24783 (N_24783,N_16394,N_13091);
and U24784 (N_24784,N_14592,N_14035);
nor U24785 (N_24785,N_19834,N_11666);
or U24786 (N_24786,N_14921,N_19582);
or U24787 (N_24787,N_16735,N_10671);
or U24788 (N_24788,N_12918,N_12555);
nor U24789 (N_24789,N_10469,N_13383);
xnor U24790 (N_24790,N_10966,N_10072);
nor U24791 (N_24791,N_12661,N_15590);
and U24792 (N_24792,N_18147,N_17139);
or U24793 (N_24793,N_17645,N_18573);
or U24794 (N_24794,N_12706,N_19619);
nand U24795 (N_24795,N_10933,N_11126);
nand U24796 (N_24796,N_17950,N_15981);
and U24797 (N_24797,N_12535,N_16954);
nor U24798 (N_24798,N_16428,N_10387);
nand U24799 (N_24799,N_18302,N_19233);
nor U24800 (N_24800,N_18503,N_10033);
or U24801 (N_24801,N_15843,N_17677);
and U24802 (N_24802,N_18303,N_10620);
and U24803 (N_24803,N_11199,N_15055);
nand U24804 (N_24804,N_12713,N_16691);
or U24805 (N_24805,N_16941,N_13427);
nor U24806 (N_24806,N_16433,N_19657);
nand U24807 (N_24807,N_19164,N_14190);
or U24808 (N_24808,N_13675,N_10019);
nor U24809 (N_24809,N_15626,N_16720);
nand U24810 (N_24810,N_15483,N_12656);
nor U24811 (N_24811,N_11640,N_16120);
and U24812 (N_24812,N_17866,N_12709);
or U24813 (N_24813,N_17389,N_12968);
or U24814 (N_24814,N_16280,N_19724);
and U24815 (N_24815,N_10559,N_12130);
or U24816 (N_24816,N_16327,N_13867);
nand U24817 (N_24817,N_16200,N_19900);
nor U24818 (N_24818,N_10524,N_14614);
nand U24819 (N_24819,N_18171,N_13560);
nand U24820 (N_24820,N_11830,N_11234);
or U24821 (N_24821,N_14814,N_17353);
nor U24822 (N_24822,N_18990,N_15522);
nor U24823 (N_24823,N_13876,N_18068);
and U24824 (N_24824,N_14651,N_13550);
nand U24825 (N_24825,N_15014,N_16873);
nor U24826 (N_24826,N_17163,N_17421);
and U24827 (N_24827,N_19754,N_15766);
nand U24828 (N_24828,N_15199,N_12181);
and U24829 (N_24829,N_16179,N_16722);
and U24830 (N_24830,N_15933,N_16695);
nor U24831 (N_24831,N_12995,N_10509);
nand U24832 (N_24832,N_11293,N_17235);
or U24833 (N_24833,N_13922,N_17932);
nand U24834 (N_24834,N_16579,N_13367);
nor U24835 (N_24835,N_11151,N_11702);
or U24836 (N_24836,N_12349,N_12772);
nand U24837 (N_24837,N_10876,N_19609);
nand U24838 (N_24838,N_16459,N_14165);
nor U24839 (N_24839,N_13164,N_18567);
nor U24840 (N_24840,N_19847,N_15467);
nand U24841 (N_24841,N_17047,N_10918);
nor U24842 (N_24842,N_19175,N_16996);
or U24843 (N_24843,N_16818,N_15427);
and U24844 (N_24844,N_12299,N_11497);
nand U24845 (N_24845,N_10704,N_12246);
or U24846 (N_24846,N_12388,N_15723);
nand U24847 (N_24847,N_18774,N_18361);
and U24848 (N_24848,N_16284,N_13535);
and U24849 (N_24849,N_17223,N_12053);
nor U24850 (N_24850,N_15033,N_11864);
or U24851 (N_24851,N_10688,N_14780);
nor U24852 (N_24852,N_15976,N_10305);
or U24853 (N_24853,N_11508,N_15555);
or U24854 (N_24854,N_15250,N_14141);
nor U24855 (N_24855,N_17569,N_11566);
nor U24856 (N_24856,N_14910,N_16535);
or U24857 (N_24857,N_11717,N_11853);
nand U24858 (N_24858,N_12138,N_11335);
nor U24859 (N_24859,N_12208,N_10659);
nor U24860 (N_24860,N_11206,N_16381);
nor U24861 (N_24861,N_19361,N_16548);
and U24862 (N_24862,N_18584,N_18778);
nor U24863 (N_24863,N_19995,N_17872);
or U24864 (N_24864,N_11382,N_14359);
and U24865 (N_24865,N_17806,N_16058);
and U24866 (N_24866,N_10042,N_13162);
or U24867 (N_24867,N_19514,N_13413);
and U24868 (N_24868,N_17691,N_13993);
nand U24869 (N_24869,N_16556,N_13610);
xor U24870 (N_24870,N_17116,N_18611);
nor U24871 (N_24871,N_15609,N_18657);
xnor U24872 (N_24872,N_13052,N_15936);
or U24873 (N_24873,N_12717,N_13961);
and U24874 (N_24874,N_13750,N_18371);
nor U24875 (N_24875,N_19462,N_15139);
nor U24876 (N_24876,N_12189,N_18706);
nand U24877 (N_24877,N_11059,N_17266);
or U24878 (N_24878,N_15995,N_17316);
and U24879 (N_24879,N_11909,N_18166);
nor U24880 (N_24880,N_15502,N_19520);
and U24881 (N_24881,N_13411,N_16874);
nand U24882 (N_24882,N_17300,N_19981);
or U24883 (N_24883,N_10205,N_16898);
or U24884 (N_24884,N_11699,N_16975);
nor U24885 (N_24885,N_11439,N_14926);
nor U24886 (N_24886,N_19589,N_12520);
and U24887 (N_24887,N_15143,N_13897);
nor U24888 (N_24888,N_11047,N_12848);
nand U24889 (N_24889,N_14147,N_18122);
nand U24890 (N_24890,N_15085,N_17498);
nor U24891 (N_24891,N_10300,N_15744);
and U24892 (N_24892,N_18879,N_19244);
and U24893 (N_24893,N_18384,N_12445);
and U24894 (N_24894,N_17215,N_13251);
nand U24895 (N_24895,N_17492,N_18472);
nor U24896 (N_24896,N_17805,N_14275);
nor U24897 (N_24897,N_15832,N_10215);
or U24898 (N_24898,N_11337,N_11292);
nand U24899 (N_24899,N_16789,N_19014);
nor U24900 (N_24900,N_19685,N_15656);
nor U24901 (N_24901,N_17961,N_18146);
nor U24902 (N_24902,N_15195,N_19646);
nand U24903 (N_24903,N_15318,N_13756);
nand U24904 (N_24904,N_19366,N_12057);
and U24905 (N_24905,N_15226,N_10862);
nand U24906 (N_24906,N_15156,N_14251);
or U24907 (N_24907,N_19561,N_14453);
nand U24908 (N_24908,N_18785,N_10600);
or U24909 (N_24909,N_11493,N_17406);
nand U24910 (N_24910,N_10904,N_19647);
nor U24911 (N_24911,N_15364,N_14669);
nor U24912 (N_24912,N_18357,N_14683);
and U24913 (N_24913,N_11624,N_12590);
and U24914 (N_24914,N_15678,N_13862);
nor U24915 (N_24915,N_12712,N_10996);
nor U24916 (N_24916,N_14526,N_18582);
or U24917 (N_24917,N_15932,N_10492);
nor U24918 (N_24918,N_12787,N_13254);
and U24919 (N_24919,N_17496,N_16448);
and U24920 (N_24920,N_13392,N_18986);
nor U24921 (N_24921,N_10840,N_11394);
nand U24922 (N_24922,N_10202,N_18590);
nand U24923 (N_24923,N_12989,N_12685);
nor U24924 (N_24924,N_16744,N_13442);
and U24925 (N_24925,N_17707,N_19636);
nand U24926 (N_24926,N_15203,N_19654);
and U24927 (N_24927,N_13285,N_12436);
or U24928 (N_24928,N_19770,N_17523);
or U24929 (N_24929,N_16878,N_14043);
and U24930 (N_24930,N_19771,N_16313);
nand U24931 (N_24931,N_17472,N_14933);
xnor U24932 (N_24932,N_12382,N_16407);
and U24933 (N_24933,N_12815,N_19198);
xnor U24934 (N_24934,N_11538,N_18406);
and U24935 (N_24935,N_13314,N_17489);
or U24936 (N_24936,N_19665,N_15127);
nand U24937 (N_24937,N_14341,N_11978);
or U24938 (N_24938,N_10438,N_13229);
nand U24939 (N_24939,N_16007,N_13185);
nand U24940 (N_24940,N_17633,N_17488);
nand U24941 (N_24941,N_15319,N_18063);
or U24942 (N_24942,N_16640,N_11455);
and U24943 (N_24943,N_18890,N_13790);
nand U24944 (N_24944,N_17656,N_19658);
and U24945 (N_24945,N_18683,N_14138);
or U24946 (N_24946,N_13149,N_19499);
or U24947 (N_24947,N_12167,N_16625);
and U24948 (N_24948,N_19170,N_16790);
nand U24949 (N_24949,N_19166,N_14995);
and U24950 (N_24950,N_19919,N_18209);
and U24951 (N_24951,N_16854,N_15008);
and U24952 (N_24952,N_16334,N_14115);
or U24953 (N_24953,N_15845,N_12896);
and U24954 (N_24954,N_18575,N_16674);
nor U24955 (N_24955,N_13234,N_15907);
nand U24956 (N_24956,N_14428,N_11213);
nand U24957 (N_24957,N_18524,N_10447);
nor U24958 (N_24958,N_10500,N_12175);
nor U24959 (N_24959,N_13629,N_16243);
nor U24960 (N_24960,N_13382,N_12032);
or U24961 (N_24961,N_12846,N_19615);
nor U24962 (N_24962,N_13915,N_14595);
nor U24963 (N_24963,N_18487,N_19921);
and U24964 (N_24964,N_13275,N_19601);
nand U24965 (N_24965,N_13703,N_18961);
or U24966 (N_24966,N_19867,N_19526);
nor U24967 (N_24967,N_10830,N_10565);
and U24968 (N_24968,N_14104,N_12669);
nor U24969 (N_24969,N_10678,N_15794);
and U24970 (N_24970,N_13083,N_13630);
xor U24971 (N_24971,N_17060,N_16928);
nand U24972 (N_24972,N_16014,N_19104);
or U24973 (N_24973,N_14730,N_15333);
nand U24974 (N_24974,N_15489,N_15396);
nand U24975 (N_24975,N_15960,N_18528);
or U24976 (N_24976,N_18679,N_17390);
nand U24977 (N_24977,N_18868,N_12132);
nand U24978 (N_24978,N_13933,N_10693);
or U24979 (N_24979,N_19312,N_16602);
nand U24980 (N_24980,N_12281,N_14841);
and U24981 (N_24981,N_11268,N_14654);
or U24982 (N_24982,N_12494,N_11606);
nor U24983 (N_24983,N_18086,N_18111);
or U24984 (N_24984,N_13890,N_18162);
and U24985 (N_24985,N_17324,N_12424);
nor U24986 (N_24986,N_19927,N_14605);
nand U24987 (N_24987,N_15695,N_11644);
and U24988 (N_24988,N_13723,N_14852);
and U24989 (N_24989,N_14604,N_17628);
nand U24990 (N_24990,N_14468,N_16565);
and U24991 (N_24991,N_15371,N_14813);
and U24992 (N_24992,N_10187,N_18758);
nand U24993 (N_24993,N_14881,N_13612);
and U24994 (N_24994,N_12475,N_19543);
or U24995 (N_24995,N_10090,N_10797);
or U24996 (N_24996,N_16516,N_15922);
nand U24997 (N_24997,N_18437,N_18635);
nand U24998 (N_24998,N_10761,N_17190);
and U24999 (N_24999,N_15524,N_18650);
nand U25000 (N_25000,N_18247,N_10562);
and U25001 (N_25001,N_11145,N_17003);
nand U25002 (N_25002,N_10570,N_19744);
and U25003 (N_25003,N_15123,N_16974);
or U25004 (N_25004,N_19433,N_18971);
or U25005 (N_25005,N_14621,N_13848);
and U25006 (N_25006,N_11647,N_13322);
and U25007 (N_25007,N_12754,N_15050);
nor U25008 (N_25008,N_16549,N_15164);
and U25009 (N_25009,N_13123,N_18424);
nand U25010 (N_25010,N_10782,N_15485);
or U25011 (N_25011,N_16960,N_18745);
and U25012 (N_25012,N_16542,N_18124);
or U25013 (N_25013,N_16448,N_17663);
nor U25014 (N_25014,N_17545,N_15058);
or U25015 (N_25015,N_10053,N_16322);
and U25016 (N_25016,N_12875,N_17712);
and U25017 (N_25017,N_14596,N_18308);
and U25018 (N_25018,N_16180,N_15980);
nand U25019 (N_25019,N_17509,N_17142);
or U25020 (N_25020,N_15011,N_14563);
and U25021 (N_25021,N_17787,N_13568);
and U25022 (N_25022,N_18409,N_15518);
nor U25023 (N_25023,N_17951,N_19807);
nand U25024 (N_25024,N_19581,N_10826);
or U25025 (N_25025,N_12393,N_18611);
nand U25026 (N_25026,N_11128,N_10484);
nor U25027 (N_25027,N_16593,N_16582);
or U25028 (N_25028,N_15468,N_16978);
or U25029 (N_25029,N_12655,N_18050);
nor U25030 (N_25030,N_17100,N_13590);
and U25031 (N_25031,N_19168,N_15761);
nor U25032 (N_25032,N_15805,N_13862);
nand U25033 (N_25033,N_10899,N_16722);
or U25034 (N_25034,N_12983,N_15451);
nand U25035 (N_25035,N_17902,N_17240);
nand U25036 (N_25036,N_16774,N_12971);
nand U25037 (N_25037,N_18155,N_12945);
and U25038 (N_25038,N_12262,N_11994);
nor U25039 (N_25039,N_16682,N_13380);
and U25040 (N_25040,N_17620,N_18534);
nor U25041 (N_25041,N_10501,N_15290);
nand U25042 (N_25042,N_16906,N_18108);
or U25043 (N_25043,N_13768,N_14564);
nor U25044 (N_25044,N_10255,N_13119);
or U25045 (N_25045,N_11985,N_14159);
and U25046 (N_25046,N_15934,N_11860);
or U25047 (N_25047,N_15086,N_14094);
and U25048 (N_25048,N_10766,N_17069);
and U25049 (N_25049,N_12812,N_10491);
nand U25050 (N_25050,N_16855,N_10957);
nor U25051 (N_25051,N_13385,N_11837);
and U25052 (N_25052,N_10940,N_16135);
nand U25053 (N_25053,N_15518,N_13142);
nor U25054 (N_25054,N_16834,N_15676);
nor U25055 (N_25055,N_17661,N_12629);
and U25056 (N_25056,N_13389,N_10967);
and U25057 (N_25057,N_14827,N_15198);
nand U25058 (N_25058,N_10207,N_17274);
nand U25059 (N_25059,N_18671,N_18144);
nand U25060 (N_25060,N_16965,N_11314);
nor U25061 (N_25061,N_12379,N_13746);
or U25062 (N_25062,N_17144,N_10799);
nor U25063 (N_25063,N_16993,N_18845);
and U25064 (N_25064,N_12497,N_13785);
or U25065 (N_25065,N_10752,N_13887);
or U25066 (N_25066,N_16228,N_13698);
nor U25067 (N_25067,N_19301,N_12853);
nand U25068 (N_25068,N_15520,N_13290);
nor U25069 (N_25069,N_15544,N_18540);
or U25070 (N_25070,N_12017,N_13380);
and U25071 (N_25071,N_18300,N_10742);
nand U25072 (N_25072,N_12306,N_17393);
xnor U25073 (N_25073,N_11981,N_14673);
nor U25074 (N_25074,N_17060,N_13363);
nand U25075 (N_25075,N_18421,N_17266);
and U25076 (N_25076,N_11622,N_11370);
and U25077 (N_25077,N_10824,N_19359);
and U25078 (N_25078,N_16836,N_17792);
nand U25079 (N_25079,N_10152,N_11280);
nor U25080 (N_25080,N_17330,N_10280);
or U25081 (N_25081,N_10990,N_18332);
or U25082 (N_25082,N_10431,N_15489);
or U25083 (N_25083,N_14336,N_18686);
nor U25084 (N_25084,N_12228,N_15137);
and U25085 (N_25085,N_10025,N_16115);
and U25086 (N_25086,N_12007,N_17879);
nand U25087 (N_25087,N_11097,N_11781);
nand U25088 (N_25088,N_18502,N_18948);
nand U25089 (N_25089,N_10889,N_15156);
or U25090 (N_25090,N_16116,N_11737);
or U25091 (N_25091,N_16985,N_12745);
or U25092 (N_25092,N_13146,N_17426);
nor U25093 (N_25093,N_14827,N_12854);
nand U25094 (N_25094,N_11336,N_19553);
nor U25095 (N_25095,N_16842,N_16568);
nand U25096 (N_25096,N_15645,N_13865);
nand U25097 (N_25097,N_12130,N_10902);
and U25098 (N_25098,N_10037,N_16583);
and U25099 (N_25099,N_14304,N_10156);
nand U25100 (N_25100,N_15737,N_17601);
or U25101 (N_25101,N_18192,N_12557);
nor U25102 (N_25102,N_12163,N_16133);
and U25103 (N_25103,N_12153,N_11672);
and U25104 (N_25104,N_13525,N_16495);
or U25105 (N_25105,N_13609,N_11938);
and U25106 (N_25106,N_17090,N_10041);
nand U25107 (N_25107,N_16150,N_11310);
nor U25108 (N_25108,N_16962,N_10813);
and U25109 (N_25109,N_17234,N_17071);
or U25110 (N_25110,N_18372,N_11260);
nor U25111 (N_25111,N_18472,N_12840);
and U25112 (N_25112,N_15093,N_17477);
nand U25113 (N_25113,N_11167,N_16380);
nand U25114 (N_25114,N_19707,N_19539);
and U25115 (N_25115,N_12608,N_14292);
and U25116 (N_25116,N_11030,N_13199);
or U25117 (N_25117,N_16268,N_15543);
or U25118 (N_25118,N_10028,N_15350);
and U25119 (N_25119,N_16021,N_14155);
nand U25120 (N_25120,N_19500,N_18548);
and U25121 (N_25121,N_14839,N_19451);
nand U25122 (N_25122,N_19101,N_16208);
or U25123 (N_25123,N_18781,N_19087);
or U25124 (N_25124,N_10046,N_14043);
and U25125 (N_25125,N_18764,N_14464);
nor U25126 (N_25126,N_11052,N_13871);
or U25127 (N_25127,N_18294,N_18569);
nor U25128 (N_25128,N_17478,N_11333);
nor U25129 (N_25129,N_18840,N_14433);
nor U25130 (N_25130,N_11375,N_12271);
nand U25131 (N_25131,N_17104,N_12089);
and U25132 (N_25132,N_15154,N_17553);
nor U25133 (N_25133,N_12926,N_15461);
nor U25134 (N_25134,N_18977,N_15682);
or U25135 (N_25135,N_19855,N_13621);
and U25136 (N_25136,N_10079,N_14458);
or U25137 (N_25137,N_17971,N_16583);
nand U25138 (N_25138,N_11716,N_19123);
nand U25139 (N_25139,N_15649,N_11108);
or U25140 (N_25140,N_12895,N_13398);
and U25141 (N_25141,N_19100,N_13929);
nor U25142 (N_25142,N_17596,N_19918);
or U25143 (N_25143,N_10255,N_14354);
nor U25144 (N_25144,N_14231,N_16782);
nor U25145 (N_25145,N_18157,N_19304);
nor U25146 (N_25146,N_19844,N_14171);
or U25147 (N_25147,N_19123,N_13046);
nand U25148 (N_25148,N_17317,N_11891);
nor U25149 (N_25149,N_10377,N_19237);
nor U25150 (N_25150,N_10525,N_17822);
or U25151 (N_25151,N_11806,N_11383);
nand U25152 (N_25152,N_12578,N_11964);
nor U25153 (N_25153,N_17914,N_12408);
nand U25154 (N_25154,N_13782,N_14945);
and U25155 (N_25155,N_15208,N_15892);
and U25156 (N_25156,N_13632,N_11149);
or U25157 (N_25157,N_11850,N_19233);
and U25158 (N_25158,N_17932,N_12654);
and U25159 (N_25159,N_13555,N_15272);
and U25160 (N_25160,N_17292,N_11819);
nor U25161 (N_25161,N_14714,N_17052);
nor U25162 (N_25162,N_12941,N_10309);
and U25163 (N_25163,N_15122,N_19062);
nand U25164 (N_25164,N_11278,N_12780);
nand U25165 (N_25165,N_10249,N_16987);
and U25166 (N_25166,N_14248,N_10851);
nor U25167 (N_25167,N_12202,N_14865);
nand U25168 (N_25168,N_16640,N_13816);
nand U25169 (N_25169,N_10028,N_18389);
nor U25170 (N_25170,N_10986,N_11697);
or U25171 (N_25171,N_18887,N_19574);
xor U25172 (N_25172,N_14655,N_10769);
and U25173 (N_25173,N_19613,N_18586);
nand U25174 (N_25174,N_16040,N_17441);
nand U25175 (N_25175,N_14462,N_13480);
nor U25176 (N_25176,N_12205,N_19332);
nor U25177 (N_25177,N_10840,N_18588);
or U25178 (N_25178,N_15775,N_14799);
or U25179 (N_25179,N_19618,N_10234);
or U25180 (N_25180,N_16220,N_12272);
nor U25181 (N_25181,N_19383,N_13786);
or U25182 (N_25182,N_16377,N_18077);
or U25183 (N_25183,N_11446,N_19507);
and U25184 (N_25184,N_12179,N_10214);
and U25185 (N_25185,N_17340,N_15901);
and U25186 (N_25186,N_15654,N_16679);
or U25187 (N_25187,N_15253,N_15498);
nand U25188 (N_25188,N_18818,N_14599);
nor U25189 (N_25189,N_10296,N_15771);
and U25190 (N_25190,N_11312,N_17440);
or U25191 (N_25191,N_10187,N_11294);
and U25192 (N_25192,N_16953,N_16633);
or U25193 (N_25193,N_18095,N_10048);
nor U25194 (N_25194,N_12867,N_18986);
and U25195 (N_25195,N_11527,N_13289);
and U25196 (N_25196,N_19046,N_14315);
nand U25197 (N_25197,N_13743,N_11057);
nor U25198 (N_25198,N_13911,N_11831);
and U25199 (N_25199,N_17192,N_12118);
nor U25200 (N_25200,N_10187,N_12037);
or U25201 (N_25201,N_16363,N_12795);
nand U25202 (N_25202,N_15746,N_13839);
or U25203 (N_25203,N_18711,N_14631);
nand U25204 (N_25204,N_11914,N_17272);
and U25205 (N_25205,N_12641,N_10485);
or U25206 (N_25206,N_13918,N_14176);
nor U25207 (N_25207,N_15395,N_13834);
or U25208 (N_25208,N_18330,N_18513);
and U25209 (N_25209,N_14384,N_10022);
or U25210 (N_25210,N_19259,N_16331);
nor U25211 (N_25211,N_13966,N_11538);
nand U25212 (N_25212,N_19690,N_10927);
or U25213 (N_25213,N_17444,N_18635);
nand U25214 (N_25214,N_19308,N_17596);
nor U25215 (N_25215,N_15765,N_16371);
and U25216 (N_25216,N_14097,N_14417);
nor U25217 (N_25217,N_18963,N_15554);
and U25218 (N_25218,N_11849,N_18640);
nand U25219 (N_25219,N_13160,N_19735);
or U25220 (N_25220,N_11012,N_12967);
and U25221 (N_25221,N_13216,N_13083);
and U25222 (N_25222,N_18389,N_16085);
or U25223 (N_25223,N_16465,N_15411);
or U25224 (N_25224,N_13583,N_12878);
nor U25225 (N_25225,N_14047,N_14958);
nand U25226 (N_25226,N_15622,N_15640);
or U25227 (N_25227,N_14630,N_14465);
and U25228 (N_25228,N_12601,N_19422);
nor U25229 (N_25229,N_13230,N_10701);
or U25230 (N_25230,N_17586,N_16671);
and U25231 (N_25231,N_18763,N_17274);
nand U25232 (N_25232,N_12221,N_12847);
and U25233 (N_25233,N_10664,N_18373);
nor U25234 (N_25234,N_18743,N_14955);
nand U25235 (N_25235,N_12658,N_17613);
and U25236 (N_25236,N_12700,N_13766);
nand U25237 (N_25237,N_18055,N_18936);
and U25238 (N_25238,N_10764,N_19487);
nand U25239 (N_25239,N_15319,N_16154);
and U25240 (N_25240,N_14240,N_19593);
nand U25241 (N_25241,N_15762,N_10253);
nand U25242 (N_25242,N_15939,N_14253);
nor U25243 (N_25243,N_15961,N_18803);
nand U25244 (N_25244,N_13905,N_10995);
and U25245 (N_25245,N_18243,N_10031);
or U25246 (N_25246,N_14791,N_15185);
or U25247 (N_25247,N_12958,N_17892);
nand U25248 (N_25248,N_12410,N_17757);
nand U25249 (N_25249,N_12502,N_16565);
nand U25250 (N_25250,N_14600,N_10712);
nor U25251 (N_25251,N_10915,N_18073);
and U25252 (N_25252,N_12568,N_13726);
or U25253 (N_25253,N_11360,N_19856);
nand U25254 (N_25254,N_19046,N_19491);
nand U25255 (N_25255,N_15166,N_13077);
nor U25256 (N_25256,N_15137,N_11531);
and U25257 (N_25257,N_17593,N_13799);
or U25258 (N_25258,N_17416,N_13913);
or U25259 (N_25259,N_15665,N_15686);
and U25260 (N_25260,N_14475,N_11973);
nor U25261 (N_25261,N_19953,N_15143);
nand U25262 (N_25262,N_15750,N_15905);
or U25263 (N_25263,N_14822,N_10105);
xor U25264 (N_25264,N_18997,N_11958);
nand U25265 (N_25265,N_14390,N_12858);
nor U25266 (N_25266,N_19224,N_17461);
and U25267 (N_25267,N_17662,N_10288);
and U25268 (N_25268,N_10165,N_10520);
and U25269 (N_25269,N_10113,N_11290);
or U25270 (N_25270,N_10931,N_16602);
or U25271 (N_25271,N_12183,N_15539);
or U25272 (N_25272,N_17896,N_15184);
nor U25273 (N_25273,N_10019,N_16517);
nor U25274 (N_25274,N_19694,N_11932);
xnor U25275 (N_25275,N_14906,N_13146);
and U25276 (N_25276,N_16295,N_11732);
or U25277 (N_25277,N_19744,N_15927);
nand U25278 (N_25278,N_17114,N_13838);
nor U25279 (N_25279,N_15401,N_10708);
nor U25280 (N_25280,N_14702,N_11880);
nor U25281 (N_25281,N_16659,N_12244);
and U25282 (N_25282,N_10601,N_10610);
and U25283 (N_25283,N_11554,N_11254);
nor U25284 (N_25284,N_13662,N_11857);
or U25285 (N_25285,N_19009,N_15099);
nor U25286 (N_25286,N_10304,N_12612);
nor U25287 (N_25287,N_10080,N_13288);
nand U25288 (N_25288,N_11154,N_13574);
and U25289 (N_25289,N_18002,N_10843);
and U25290 (N_25290,N_14260,N_18607);
nor U25291 (N_25291,N_17682,N_17540);
and U25292 (N_25292,N_12109,N_15244);
nand U25293 (N_25293,N_15902,N_15816);
or U25294 (N_25294,N_15917,N_11912);
and U25295 (N_25295,N_15570,N_13334);
or U25296 (N_25296,N_11097,N_11920);
and U25297 (N_25297,N_10759,N_18814);
nor U25298 (N_25298,N_16218,N_14776);
and U25299 (N_25299,N_10364,N_14213);
and U25300 (N_25300,N_19896,N_14421);
nand U25301 (N_25301,N_17979,N_19853);
nor U25302 (N_25302,N_13159,N_12377);
or U25303 (N_25303,N_14704,N_13767);
nand U25304 (N_25304,N_16812,N_13652);
nor U25305 (N_25305,N_17449,N_14730);
nor U25306 (N_25306,N_19735,N_11119);
and U25307 (N_25307,N_16772,N_16412);
or U25308 (N_25308,N_11112,N_11376);
and U25309 (N_25309,N_12729,N_10996);
and U25310 (N_25310,N_15149,N_12456);
or U25311 (N_25311,N_15247,N_12200);
nand U25312 (N_25312,N_14191,N_19137);
or U25313 (N_25313,N_10903,N_10776);
nand U25314 (N_25314,N_16022,N_17774);
or U25315 (N_25315,N_14350,N_10030);
and U25316 (N_25316,N_19111,N_11387);
and U25317 (N_25317,N_16697,N_18129);
nor U25318 (N_25318,N_17650,N_18580);
nor U25319 (N_25319,N_15648,N_13310);
or U25320 (N_25320,N_16952,N_12099);
nor U25321 (N_25321,N_15031,N_15806);
nand U25322 (N_25322,N_13031,N_12116);
nor U25323 (N_25323,N_19012,N_12372);
nand U25324 (N_25324,N_16242,N_10746);
nor U25325 (N_25325,N_11965,N_13660);
or U25326 (N_25326,N_18136,N_19348);
nand U25327 (N_25327,N_18924,N_12358);
nor U25328 (N_25328,N_14210,N_10846);
or U25329 (N_25329,N_16762,N_16177);
or U25330 (N_25330,N_18730,N_15282);
and U25331 (N_25331,N_14946,N_17221);
or U25332 (N_25332,N_17418,N_16717);
nor U25333 (N_25333,N_16398,N_13027);
or U25334 (N_25334,N_12174,N_11406);
nor U25335 (N_25335,N_17707,N_19904);
and U25336 (N_25336,N_14293,N_12990);
nor U25337 (N_25337,N_16562,N_18627);
nor U25338 (N_25338,N_10255,N_11974);
or U25339 (N_25339,N_10536,N_10391);
nor U25340 (N_25340,N_18648,N_18592);
nor U25341 (N_25341,N_11177,N_17957);
nor U25342 (N_25342,N_12722,N_14945);
nor U25343 (N_25343,N_16079,N_11371);
nor U25344 (N_25344,N_13336,N_17241);
or U25345 (N_25345,N_16748,N_15155);
nand U25346 (N_25346,N_19297,N_15163);
or U25347 (N_25347,N_15375,N_15034);
nor U25348 (N_25348,N_11500,N_19935);
nand U25349 (N_25349,N_16863,N_14728);
or U25350 (N_25350,N_16059,N_14234);
or U25351 (N_25351,N_14833,N_15547);
nor U25352 (N_25352,N_14832,N_16927);
nor U25353 (N_25353,N_16431,N_13880);
or U25354 (N_25354,N_11482,N_11085);
nand U25355 (N_25355,N_13500,N_17035);
and U25356 (N_25356,N_12810,N_14431);
or U25357 (N_25357,N_13089,N_10233);
nor U25358 (N_25358,N_11636,N_10768);
or U25359 (N_25359,N_15180,N_16522);
nor U25360 (N_25360,N_13465,N_18756);
nor U25361 (N_25361,N_17059,N_15297);
nand U25362 (N_25362,N_16512,N_19160);
nor U25363 (N_25363,N_11837,N_14919);
nor U25364 (N_25364,N_14306,N_10634);
nor U25365 (N_25365,N_17416,N_15294);
or U25366 (N_25366,N_16154,N_17256);
nand U25367 (N_25367,N_18312,N_10042);
nor U25368 (N_25368,N_11487,N_17597);
nand U25369 (N_25369,N_19083,N_13335);
and U25370 (N_25370,N_16430,N_19025);
and U25371 (N_25371,N_12751,N_14563);
nor U25372 (N_25372,N_15644,N_14002);
nand U25373 (N_25373,N_14224,N_16193);
and U25374 (N_25374,N_15205,N_18688);
nand U25375 (N_25375,N_14084,N_12489);
nand U25376 (N_25376,N_14004,N_17905);
or U25377 (N_25377,N_12778,N_15105);
nor U25378 (N_25378,N_14965,N_13444);
or U25379 (N_25379,N_15140,N_19869);
and U25380 (N_25380,N_18875,N_19391);
nand U25381 (N_25381,N_10844,N_14226);
or U25382 (N_25382,N_11904,N_16523);
nor U25383 (N_25383,N_12154,N_14172);
and U25384 (N_25384,N_15191,N_18851);
nand U25385 (N_25385,N_18678,N_18764);
nor U25386 (N_25386,N_14758,N_12135);
nor U25387 (N_25387,N_19740,N_19700);
nand U25388 (N_25388,N_11988,N_18223);
or U25389 (N_25389,N_11148,N_18669);
nor U25390 (N_25390,N_14065,N_12405);
nor U25391 (N_25391,N_10119,N_18850);
and U25392 (N_25392,N_12932,N_18328);
or U25393 (N_25393,N_15748,N_18919);
or U25394 (N_25394,N_13838,N_13512);
nor U25395 (N_25395,N_19695,N_14763);
nor U25396 (N_25396,N_15779,N_15031);
xnor U25397 (N_25397,N_15141,N_14415);
and U25398 (N_25398,N_12965,N_15583);
and U25399 (N_25399,N_15248,N_10354);
nor U25400 (N_25400,N_10334,N_10080);
nor U25401 (N_25401,N_14608,N_11326);
or U25402 (N_25402,N_18316,N_19859);
nor U25403 (N_25403,N_14073,N_18813);
and U25404 (N_25404,N_15578,N_11981);
nand U25405 (N_25405,N_15841,N_18512);
nand U25406 (N_25406,N_13207,N_12952);
nand U25407 (N_25407,N_13462,N_16946);
and U25408 (N_25408,N_13857,N_19042);
or U25409 (N_25409,N_18116,N_15820);
xor U25410 (N_25410,N_16812,N_11941);
nand U25411 (N_25411,N_17405,N_11918);
nor U25412 (N_25412,N_19686,N_15781);
nor U25413 (N_25413,N_12780,N_16443);
or U25414 (N_25414,N_17578,N_18641);
or U25415 (N_25415,N_17952,N_16910);
or U25416 (N_25416,N_19693,N_16954);
or U25417 (N_25417,N_11581,N_11013);
nor U25418 (N_25418,N_15224,N_13123);
nor U25419 (N_25419,N_19646,N_17020);
nand U25420 (N_25420,N_14426,N_11595);
and U25421 (N_25421,N_17743,N_12420);
nand U25422 (N_25422,N_16126,N_16664);
or U25423 (N_25423,N_15657,N_16278);
and U25424 (N_25424,N_16964,N_12247);
and U25425 (N_25425,N_14907,N_13961);
nor U25426 (N_25426,N_17599,N_17511);
and U25427 (N_25427,N_11457,N_14332);
or U25428 (N_25428,N_15394,N_18735);
nand U25429 (N_25429,N_10319,N_16099);
nor U25430 (N_25430,N_19838,N_13204);
or U25431 (N_25431,N_10801,N_15139);
nand U25432 (N_25432,N_15917,N_11590);
or U25433 (N_25433,N_14150,N_15298);
and U25434 (N_25434,N_17654,N_15028);
and U25435 (N_25435,N_13609,N_14591);
nor U25436 (N_25436,N_13658,N_19779);
nand U25437 (N_25437,N_13701,N_17881);
and U25438 (N_25438,N_10044,N_16945);
nor U25439 (N_25439,N_15064,N_11138);
or U25440 (N_25440,N_10464,N_13519);
nor U25441 (N_25441,N_18685,N_11204);
nor U25442 (N_25442,N_14589,N_18967);
and U25443 (N_25443,N_18989,N_19351);
or U25444 (N_25444,N_12699,N_13688);
and U25445 (N_25445,N_17687,N_11549);
nor U25446 (N_25446,N_19585,N_15847);
nand U25447 (N_25447,N_11655,N_13098);
or U25448 (N_25448,N_12337,N_11247);
nor U25449 (N_25449,N_19749,N_15709);
or U25450 (N_25450,N_14440,N_17098);
and U25451 (N_25451,N_15298,N_11441);
or U25452 (N_25452,N_18180,N_11621);
nand U25453 (N_25453,N_11859,N_10779);
nor U25454 (N_25454,N_15160,N_11961);
xnor U25455 (N_25455,N_18162,N_16953);
and U25456 (N_25456,N_14438,N_14607);
nand U25457 (N_25457,N_19979,N_12939);
or U25458 (N_25458,N_19066,N_18568);
nor U25459 (N_25459,N_10954,N_10890);
nand U25460 (N_25460,N_13421,N_18771);
nor U25461 (N_25461,N_17995,N_14439);
nor U25462 (N_25462,N_16480,N_17146);
nand U25463 (N_25463,N_19247,N_17429);
nor U25464 (N_25464,N_14532,N_16543);
and U25465 (N_25465,N_10738,N_14671);
nand U25466 (N_25466,N_14430,N_11300);
nor U25467 (N_25467,N_18901,N_19953);
and U25468 (N_25468,N_10183,N_14447);
or U25469 (N_25469,N_14498,N_11364);
nand U25470 (N_25470,N_14013,N_18080);
and U25471 (N_25471,N_12379,N_19286);
nand U25472 (N_25472,N_18906,N_17149);
nor U25473 (N_25473,N_17396,N_13452);
nand U25474 (N_25474,N_19512,N_15892);
nor U25475 (N_25475,N_18735,N_15350);
xor U25476 (N_25476,N_16541,N_17353);
nor U25477 (N_25477,N_13056,N_19609);
and U25478 (N_25478,N_17798,N_17761);
or U25479 (N_25479,N_11164,N_13837);
nand U25480 (N_25480,N_10351,N_16296);
nor U25481 (N_25481,N_17983,N_10173);
nor U25482 (N_25482,N_17765,N_12800);
and U25483 (N_25483,N_16124,N_13425);
and U25484 (N_25484,N_14421,N_14806);
and U25485 (N_25485,N_12635,N_13478);
and U25486 (N_25486,N_13897,N_12516);
nor U25487 (N_25487,N_13131,N_19023);
nand U25488 (N_25488,N_19071,N_11931);
or U25489 (N_25489,N_11460,N_16549);
nor U25490 (N_25490,N_14555,N_19292);
and U25491 (N_25491,N_10595,N_15909);
and U25492 (N_25492,N_10127,N_17051);
nand U25493 (N_25493,N_15950,N_11476);
and U25494 (N_25494,N_19605,N_14242);
or U25495 (N_25495,N_15307,N_11252);
and U25496 (N_25496,N_13864,N_14327);
or U25497 (N_25497,N_14034,N_13432);
nor U25498 (N_25498,N_16324,N_12892);
nor U25499 (N_25499,N_13356,N_10990);
or U25500 (N_25500,N_12522,N_18095);
nor U25501 (N_25501,N_18578,N_14077);
or U25502 (N_25502,N_11792,N_10322);
and U25503 (N_25503,N_14425,N_15917);
or U25504 (N_25504,N_18009,N_14696);
or U25505 (N_25505,N_16331,N_13999);
nor U25506 (N_25506,N_14201,N_13318);
or U25507 (N_25507,N_17635,N_11135);
nand U25508 (N_25508,N_17498,N_17002);
nor U25509 (N_25509,N_18496,N_15344);
and U25510 (N_25510,N_15349,N_12473);
nor U25511 (N_25511,N_18866,N_10397);
nand U25512 (N_25512,N_10306,N_17426);
or U25513 (N_25513,N_19154,N_10204);
or U25514 (N_25514,N_11647,N_13496);
nor U25515 (N_25515,N_11589,N_11099);
nor U25516 (N_25516,N_12821,N_18339);
and U25517 (N_25517,N_13992,N_14311);
nor U25518 (N_25518,N_18455,N_15758);
or U25519 (N_25519,N_15831,N_11888);
nor U25520 (N_25520,N_17293,N_12874);
nor U25521 (N_25521,N_15101,N_16960);
and U25522 (N_25522,N_19760,N_14212);
nor U25523 (N_25523,N_11762,N_10005);
or U25524 (N_25524,N_13541,N_14790);
nor U25525 (N_25525,N_16571,N_12327);
nor U25526 (N_25526,N_13760,N_19334);
nand U25527 (N_25527,N_13385,N_19510);
and U25528 (N_25528,N_18643,N_10017);
xnor U25529 (N_25529,N_16518,N_14706);
or U25530 (N_25530,N_10019,N_13281);
and U25531 (N_25531,N_16691,N_10110);
nand U25532 (N_25532,N_14024,N_19717);
and U25533 (N_25533,N_19766,N_11769);
and U25534 (N_25534,N_10821,N_11058);
nor U25535 (N_25535,N_17937,N_11309);
nand U25536 (N_25536,N_17910,N_14611);
nand U25537 (N_25537,N_14857,N_19465);
or U25538 (N_25538,N_14775,N_11958);
nand U25539 (N_25539,N_17975,N_16886);
nor U25540 (N_25540,N_10333,N_18236);
or U25541 (N_25541,N_19661,N_17617);
and U25542 (N_25542,N_11528,N_14180);
or U25543 (N_25543,N_11451,N_14234);
and U25544 (N_25544,N_11354,N_12667);
nand U25545 (N_25545,N_10501,N_18387);
and U25546 (N_25546,N_15392,N_17491);
nand U25547 (N_25547,N_15976,N_11235);
xnor U25548 (N_25548,N_19409,N_10218);
or U25549 (N_25549,N_11464,N_10253);
nor U25550 (N_25550,N_18416,N_13081);
and U25551 (N_25551,N_15193,N_11541);
or U25552 (N_25552,N_10720,N_15350);
nand U25553 (N_25553,N_19617,N_13487);
nor U25554 (N_25554,N_16006,N_13519);
nor U25555 (N_25555,N_17616,N_14182);
nand U25556 (N_25556,N_17913,N_18770);
nor U25557 (N_25557,N_15882,N_12430);
and U25558 (N_25558,N_11897,N_11339);
and U25559 (N_25559,N_18999,N_16292);
nor U25560 (N_25560,N_10043,N_16866);
nand U25561 (N_25561,N_14051,N_14388);
nand U25562 (N_25562,N_15813,N_11830);
or U25563 (N_25563,N_13150,N_19120);
nor U25564 (N_25564,N_14417,N_18821);
and U25565 (N_25565,N_12832,N_15402);
or U25566 (N_25566,N_18694,N_11305);
nand U25567 (N_25567,N_19303,N_15712);
nor U25568 (N_25568,N_19614,N_14544);
and U25569 (N_25569,N_16467,N_11194);
nand U25570 (N_25570,N_14822,N_18685);
or U25571 (N_25571,N_11503,N_17412);
or U25572 (N_25572,N_12016,N_17051);
nand U25573 (N_25573,N_14030,N_16784);
or U25574 (N_25574,N_14450,N_15296);
or U25575 (N_25575,N_19192,N_16758);
or U25576 (N_25576,N_12153,N_11808);
nor U25577 (N_25577,N_18545,N_19820);
or U25578 (N_25578,N_10932,N_18739);
and U25579 (N_25579,N_15794,N_14778);
or U25580 (N_25580,N_15723,N_14021);
or U25581 (N_25581,N_14025,N_17767);
or U25582 (N_25582,N_18213,N_13415);
or U25583 (N_25583,N_19923,N_13437);
nand U25584 (N_25584,N_10900,N_14122);
and U25585 (N_25585,N_17777,N_12793);
and U25586 (N_25586,N_19332,N_13183);
nor U25587 (N_25587,N_15234,N_12727);
or U25588 (N_25588,N_10225,N_11183);
nor U25589 (N_25589,N_15236,N_19502);
xnor U25590 (N_25590,N_17692,N_16253);
and U25591 (N_25591,N_16543,N_11541);
nand U25592 (N_25592,N_12556,N_15270);
nor U25593 (N_25593,N_12321,N_16727);
and U25594 (N_25594,N_13946,N_18400);
nor U25595 (N_25595,N_18085,N_12143);
or U25596 (N_25596,N_13698,N_13950);
nand U25597 (N_25597,N_10519,N_19945);
nor U25598 (N_25598,N_15616,N_11447);
xor U25599 (N_25599,N_18086,N_19024);
nor U25600 (N_25600,N_19513,N_15172);
or U25601 (N_25601,N_14279,N_15282);
and U25602 (N_25602,N_16487,N_18409);
and U25603 (N_25603,N_10903,N_14255);
nand U25604 (N_25604,N_11811,N_18352);
nand U25605 (N_25605,N_10914,N_16367);
nor U25606 (N_25606,N_15007,N_14445);
nand U25607 (N_25607,N_11645,N_16411);
or U25608 (N_25608,N_14210,N_10750);
or U25609 (N_25609,N_12190,N_13335);
nor U25610 (N_25610,N_10841,N_10995);
nor U25611 (N_25611,N_14336,N_13674);
xnor U25612 (N_25612,N_16528,N_16553);
nor U25613 (N_25613,N_18265,N_17428);
or U25614 (N_25614,N_10958,N_12990);
or U25615 (N_25615,N_16868,N_12519);
nand U25616 (N_25616,N_12054,N_14697);
or U25617 (N_25617,N_18936,N_17560);
or U25618 (N_25618,N_12560,N_14867);
or U25619 (N_25619,N_12704,N_11098);
nand U25620 (N_25620,N_12211,N_13746);
and U25621 (N_25621,N_15844,N_14183);
nand U25622 (N_25622,N_19560,N_13124);
nand U25623 (N_25623,N_19243,N_17275);
xor U25624 (N_25624,N_19021,N_18555);
nor U25625 (N_25625,N_13585,N_19078);
or U25626 (N_25626,N_13413,N_11867);
or U25627 (N_25627,N_19971,N_17183);
or U25628 (N_25628,N_19295,N_14607);
and U25629 (N_25629,N_12791,N_18350);
and U25630 (N_25630,N_14941,N_11879);
and U25631 (N_25631,N_18903,N_10843);
and U25632 (N_25632,N_18742,N_12937);
and U25633 (N_25633,N_18369,N_14443);
and U25634 (N_25634,N_13812,N_18306);
or U25635 (N_25635,N_16334,N_15190);
nand U25636 (N_25636,N_19541,N_14028);
nor U25637 (N_25637,N_10522,N_14322);
nand U25638 (N_25638,N_16575,N_18430);
and U25639 (N_25639,N_14254,N_10778);
and U25640 (N_25640,N_11699,N_13444);
nor U25641 (N_25641,N_11245,N_13242);
and U25642 (N_25642,N_10863,N_15252);
and U25643 (N_25643,N_15737,N_11183);
nand U25644 (N_25644,N_17518,N_10793);
nor U25645 (N_25645,N_14957,N_12486);
xor U25646 (N_25646,N_18400,N_19167);
nor U25647 (N_25647,N_15093,N_18566);
nand U25648 (N_25648,N_11271,N_18948);
and U25649 (N_25649,N_16620,N_19381);
xnor U25650 (N_25650,N_15672,N_19314);
nor U25651 (N_25651,N_18141,N_11888);
nor U25652 (N_25652,N_15841,N_12142);
nor U25653 (N_25653,N_12206,N_11695);
or U25654 (N_25654,N_19970,N_16826);
nor U25655 (N_25655,N_17109,N_17588);
nor U25656 (N_25656,N_15044,N_14347);
nand U25657 (N_25657,N_14401,N_13904);
and U25658 (N_25658,N_11765,N_12622);
and U25659 (N_25659,N_12703,N_15808);
nand U25660 (N_25660,N_13440,N_12141);
nor U25661 (N_25661,N_17173,N_14930);
nand U25662 (N_25662,N_11198,N_14779);
and U25663 (N_25663,N_13874,N_11936);
nand U25664 (N_25664,N_11068,N_18278);
and U25665 (N_25665,N_16294,N_16890);
or U25666 (N_25666,N_19052,N_10363);
or U25667 (N_25667,N_12289,N_15169);
or U25668 (N_25668,N_15571,N_15533);
nor U25669 (N_25669,N_13627,N_10818);
nor U25670 (N_25670,N_19157,N_10538);
nand U25671 (N_25671,N_16302,N_10328);
or U25672 (N_25672,N_16380,N_11394);
or U25673 (N_25673,N_11826,N_13724);
nand U25674 (N_25674,N_10084,N_16102);
xor U25675 (N_25675,N_12406,N_19247);
nand U25676 (N_25676,N_12134,N_16376);
or U25677 (N_25677,N_18140,N_11887);
nand U25678 (N_25678,N_14994,N_12156);
and U25679 (N_25679,N_18556,N_13895);
and U25680 (N_25680,N_19105,N_15187);
or U25681 (N_25681,N_15834,N_11986);
and U25682 (N_25682,N_11825,N_14215);
or U25683 (N_25683,N_18866,N_16164);
and U25684 (N_25684,N_10750,N_18965);
nand U25685 (N_25685,N_10634,N_13811);
nand U25686 (N_25686,N_10515,N_18968);
and U25687 (N_25687,N_10279,N_10517);
nand U25688 (N_25688,N_16347,N_18056);
nand U25689 (N_25689,N_12069,N_18742);
and U25690 (N_25690,N_16410,N_16104);
and U25691 (N_25691,N_12240,N_17278);
nor U25692 (N_25692,N_15847,N_16052);
or U25693 (N_25693,N_18357,N_14577);
nand U25694 (N_25694,N_18699,N_10591);
or U25695 (N_25695,N_19148,N_12735);
nor U25696 (N_25696,N_18810,N_18053);
and U25697 (N_25697,N_16388,N_18654);
or U25698 (N_25698,N_17953,N_17937);
nand U25699 (N_25699,N_11738,N_18786);
or U25700 (N_25700,N_13948,N_11335);
nand U25701 (N_25701,N_18147,N_11729);
and U25702 (N_25702,N_16745,N_14475);
nor U25703 (N_25703,N_14152,N_15093);
nor U25704 (N_25704,N_18769,N_17430);
nand U25705 (N_25705,N_17890,N_15032);
nor U25706 (N_25706,N_16115,N_19664);
or U25707 (N_25707,N_13542,N_18209);
and U25708 (N_25708,N_15670,N_14324);
or U25709 (N_25709,N_16278,N_11719);
or U25710 (N_25710,N_13883,N_16188);
and U25711 (N_25711,N_12637,N_12079);
nor U25712 (N_25712,N_16125,N_10909);
nor U25713 (N_25713,N_12504,N_18011);
or U25714 (N_25714,N_19667,N_16092);
or U25715 (N_25715,N_13395,N_12619);
nor U25716 (N_25716,N_19151,N_13971);
nor U25717 (N_25717,N_10949,N_18416);
nor U25718 (N_25718,N_15745,N_12492);
nor U25719 (N_25719,N_10227,N_18844);
nor U25720 (N_25720,N_16912,N_14691);
nand U25721 (N_25721,N_10605,N_13044);
nor U25722 (N_25722,N_18679,N_11188);
or U25723 (N_25723,N_19136,N_13149);
nand U25724 (N_25724,N_12317,N_16061);
and U25725 (N_25725,N_12268,N_16490);
and U25726 (N_25726,N_14645,N_10702);
nand U25727 (N_25727,N_18931,N_17958);
and U25728 (N_25728,N_14983,N_18701);
nand U25729 (N_25729,N_13786,N_16357);
nor U25730 (N_25730,N_12023,N_17448);
or U25731 (N_25731,N_17162,N_14480);
and U25732 (N_25732,N_18609,N_19997);
nor U25733 (N_25733,N_13372,N_11018);
or U25734 (N_25734,N_17214,N_11041);
nand U25735 (N_25735,N_14292,N_15660);
or U25736 (N_25736,N_16419,N_11534);
or U25737 (N_25737,N_13546,N_15829);
nand U25738 (N_25738,N_11962,N_19039);
nor U25739 (N_25739,N_14989,N_18125);
and U25740 (N_25740,N_11352,N_18421);
nor U25741 (N_25741,N_10069,N_14723);
nand U25742 (N_25742,N_15376,N_18319);
nor U25743 (N_25743,N_15211,N_15873);
nor U25744 (N_25744,N_19750,N_14666);
nand U25745 (N_25745,N_17656,N_16955);
nor U25746 (N_25746,N_16126,N_15972);
or U25747 (N_25747,N_18106,N_10805);
nand U25748 (N_25748,N_13677,N_19817);
nand U25749 (N_25749,N_15015,N_15530);
or U25750 (N_25750,N_16787,N_15050);
xnor U25751 (N_25751,N_18821,N_11826);
nor U25752 (N_25752,N_14792,N_13827);
or U25753 (N_25753,N_12334,N_19088);
nand U25754 (N_25754,N_15895,N_13257);
nor U25755 (N_25755,N_13897,N_19878);
or U25756 (N_25756,N_18526,N_16787);
nor U25757 (N_25757,N_13676,N_19049);
or U25758 (N_25758,N_18583,N_10005);
or U25759 (N_25759,N_16933,N_11001);
nor U25760 (N_25760,N_19092,N_19693);
nand U25761 (N_25761,N_16923,N_14180);
or U25762 (N_25762,N_15192,N_19683);
or U25763 (N_25763,N_19408,N_17649);
nor U25764 (N_25764,N_19239,N_11598);
or U25765 (N_25765,N_15052,N_18751);
nand U25766 (N_25766,N_19143,N_17391);
nor U25767 (N_25767,N_12520,N_15449);
xnor U25768 (N_25768,N_11959,N_19179);
xnor U25769 (N_25769,N_14729,N_13463);
and U25770 (N_25770,N_15339,N_13163);
and U25771 (N_25771,N_16966,N_14266);
or U25772 (N_25772,N_13954,N_19554);
or U25773 (N_25773,N_10372,N_10514);
or U25774 (N_25774,N_10787,N_15822);
nor U25775 (N_25775,N_16572,N_16772);
nand U25776 (N_25776,N_11335,N_10119);
or U25777 (N_25777,N_18288,N_13737);
nor U25778 (N_25778,N_15043,N_11269);
and U25779 (N_25779,N_17146,N_11885);
and U25780 (N_25780,N_14105,N_10047);
or U25781 (N_25781,N_14035,N_17865);
nor U25782 (N_25782,N_18172,N_11748);
nand U25783 (N_25783,N_10783,N_12872);
nand U25784 (N_25784,N_16751,N_18695);
nor U25785 (N_25785,N_16960,N_16509);
nor U25786 (N_25786,N_16384,N_14826);
nor U25787 (N_25787,N_14015,N_12147);
or U25788 (N_25788,N_18962,N_10598);
nor U25789 (N_25789,N_16857,N_13819);
or U25790 (N_25790,N_12044,N_17469);
nor U25791 (N_25791,N_10635,N_15942);
and U25792 (N_25792,N_10129,N_11207);
nand U25793 (N_25793,N_12974,N_14571);
and U25794 (N_25794,N_10998,N_12993);
nor U25795 (N_25795,N_13527,N_11686);
nor U25796 (N_25796,N_15535,N_11537);
nand U25797 (N_25797,N_19430,N_10630);
nor U25798 (N_25798,N_15275,N_19865);
nand U25799 (N_25799,N_13794,N_14194);
and U25800 (N_25800,N_11781,N_17698);
nor U25801 (N_25801,N_13728,N_18955);
and U25802 (N_25802,N_16812,N_12359);
and U25803 (N_25803,N_15009,N_19540);
nor U25804 (N_25804,N_19794,N_10390);
or U25805 (N_25805,N_12936,N_13124);
and U25806 (N_25806,N_13264,N_16778);
or U25807 (N_25807,N_14247,N_18152);
and U25808 (N_25808,N_19338,N_13988);
and U25809 (N_25809,N_14944,N_16818);
and U25810 (N_25810,N_15512,N_18094);
or U25811 (N_25811,N_11696,N_14773);
nor U25812 (N_25812,N_15339,N_16191);
or U25813 (N_25813,N_18876,N_12431);
and U25814 (N_25814,N_16761,N_15104);
nor U25815 (N_25815,N_12161,N_16063);
nor U25816 (N_25816,N_12227,N_18145);
and U25817 (N_25817,N_14839,N_12484);
or U25818 (N_25818,N_15734,N_18394);
or U25819 (N_25819,N_15036,N_19728);
or U25820 (N_25820,N_13334,N_17868);
or U25821 (N_25821,N_18804,N_12874);
and U25822 (N_25822,N_15407,N_18747);
or U25823 (N_25823,N_18546,N_12963);
and U25824 (N_25824,N_17145,N_12432);
or U25825 (N_25825,N_12045,N_15181);
nor U25826 (N_25826,N_10265,N_19644);
nand U25827 (N_25827,N_10379,N_14776);
nand U25828 (N_25828,N_19832,N_18029);
and U25829 (N_25829,N_17681,N_11512);
and U25830 (N_25830,N_13113,N_18179);
nor U25831 (N_25831,N_16721,N_16052);
nand U25832 (N_25832,N_14044,N_15587);
or U25833 (N_25833,N_12257,N_19561);
nand U25834 (N_25834,N_14907,N_15286);
nor U25835 (N_25835,N_16249,N_16570);
or U25836 (N_25836,N_16508,N_12695);
and U25837 (N_25837,N_11854,N_19446);
nand U25838 (N_25838,N_18766,N_14255);
nor U25839 (N_25839,N_19631,N_18626);
nor U25840 (N_25840,N_17941,N_13861);
nand U25841 (N_25841,N_10425,N_13423);
nand U25842 (N_25842,N_15313,N_14509);
nand U25843 (N_25843,N_11603,N_13548);
and U25844 (N_25844,N_14284,N_17785);
or U25845 (N_25845,N_13587,N_12828);
nand U25846 (N_25846,N_14027,N_16827);
or U25847 (N_25847,N_11977,N_19211);
nand U25848 (N_25848,N_12622,N_13272);
nor U25849 (N_25849,N_10686,N_16819);
and U25850 (N_25850,N_12202,N_17708);
or U25851 (N_25851,N_10493,N_15906);
and U25852 (N_25852,N_11731,N_16168);
and U25853 (N_25853,N_15275,N_17904);
nand U25854 (N_25854,N_12249,N_19077);
nand U25855 (N_25855,N_14931,N_15492);
and U25856 (N_25856,N_13220,N_17196);
nor U25857 (N_25857,N_14078,N_10025);
nand U25858 (N_25858,N_13271,N_15056);
and U25859 (N_25859,N_10808,N_19345);
or U25860 (N_25860,N_10164,N_17048);
or U25861 (N_25861,N_13816,N_15159);
and U25862 (N_25862,N_10569,N_11558);
and U25863 (N_25863,N_11783,N_14357);
nand U25864 (N_25864,N_17012,N_18415);
nor U25865 (N_25865,N_12894,N_18328);
or U25866 (N_25866,N_15237,N_14733);
and U25867 (N_25867,N_12016,N_11310);
or U25868 (N_25868,N_10295,N_10119);
and U25869 (N_25869,N_12794,N_15767);
nand U25870 (N_25870,N_16455,N_19675);
nand U25871 (N_25871,N_10232,N_14399);
or U25872 (N_25872,N_14632,N_14271);
and U25873 (N_25873,N_11674,N_18220);
or U25874 (N_25874,N_17531,N_11647);
nor U25875 (N_25875,N_14196,N_16332);
and U25876 (N_25876,N_13483,N_18083);
or U25877 (N_25877,N_11080,N_15008);
nor U25878 (N_25878,N_12696,N_19203);
xnor U25879 (N_25879,N_11426,N_16390);
and U25880 (N_25880,N_12566,N_18411);
or U25881 (N_25881,N_10622,N_17404);
or U25882 (N_25882,N_11397,N_13127);
nand U25883 (N_25883,N_15249,N_18380);
nor U25884 (N_25884,N_17392,N_15413);
nand U25885 (N_25885,N_10029,N_15132);
or U25886 (N_25886,N_13516,N_10075);
nand U25887 (N_25887,N_14365,N_13662);
nor U25888 (N_25888,N_13708,N_10318);
or U25889 (N_25889,N_14440,N_17373);
and U25890 (N_25890,N_15572,N_17907);
nor U25891 (N_25891,N_19129,N_17472);
nand U25892 (N_25892,N_14699,N_13587);
nand U25893 (N_25893,N_19773,N_10656);
nand U25894 (N_25894,N_17758,N_15653);
nand U25895 (N_25895,N_15689,N_10178);
and U25896 (N_25896,N_12923,N_13970);
nor U25897 (N_25897,N_19646,N_19074);
and U25898 (N_25898,N_11423,N_19244);
or U25899 (N_25899,N_14886,N_19732);
and U25900 (N_25900,N_18236,N_18534);
nand U25901 (N_25901,N_15453,N_18763);
and U25902 (N_25902,N_18220,N_19518);
nand U25903 (N_25903,N_12394,N_12180);
nor U25904 (N_25904,N_18188,N_15587);
nor U25905 (N_25905,N_14755,N_16602);
xnor U25906 (N_25906,N_11207,N_11493);
or U25907 (N_25907,N_12472,N_17346);
nand U25908 (N_25908,N_12919,N_17374);
or U25909 (N_25909,N_15700,N_19438);
and U25910 (N_25910,N_16398,N_14364);
nor U25911 (N_25911,N_11787,N_17252);
nand U25912 (N_25912,N_16848,N_11415);
or U25913 (N_25913,N_16336,N_12463);
and U25914 (N_25914,N_16364,N_10791);
and U25915 (N_25915,N_18120,N_15359);
nor U25916 (N_25916,N_11961,N_13832);
nor U25917 (N_25917,N_18873,N_13901);
and U25918 (N_25918,N_10737,N_16249);
nor U25919 (N_25919,N_17989,N_10426);
or U25920 (N_25920,N_19167,N_17512);
nor U25921 (N_25921,N_16986,N_16972);
xor U25922 (N_25922,N_16680,N_11937);
nor U25923 (N_25923,N_11492,N_11570);
and U25924 (N_25924,N_19849,N_16090);
nor U25925 (N_25925,N_18242,N_18071);
nand U25926 (N_25926,N_14859,N_11829);
or U25927 (N_25927,N_14168,N_18778);
nand U25928 (N_25928,N_10207,N_17479);
or U25929 (N_25929,N_18723,N_12734);
nand U25930 (N_25930,N_17664,N_12262);
nor U25931 (N_25931,N_19261,N_10367);
or U25932 (N_25932,N_18070,N_14268);
nor U25933 (N_25933,N_11043,N_16225);
nand U25934 (N_25934,N_16813,N_15076);
or U25935 (N_25935,N_14753,N_17859);
and U25936 (N_25936,N_12735,N_19686);
nand U25937 (N_25937,N_17961,N_16081);
xor U25938 (N_25938,N_12793,N_14541);
nor U25939 (N_25939,N_13013,N_13088);
nand U25940 (N_25940,N_13161,N_19425);
nor U25941 (N_25941,N_13615,N_18132);
and U25942 (N_25942,N_14306,N_14240);
and U25943 (N_25943,N_12856,N_13262);
and U25944 (N_25944,N_11645,N_10675);
nand U25945 (N_25945,N_19665,N_11438);
or U25946 (N_25946,N_17871,N_15923);
nor U25947 (N_25947,N_19755,N_11315);
nand U25948 (N_25948,N_10798,N_12667);
nor U25949 (N_25949,N_15869,N_16740);
and U25950 (N_25950,N_12550,N_16222);
nor U25951 (N_25951,N_12900,N_12285);
or U25952 (N_25952,N_17844,N_17959);
nand U25953 (N_25953,N_19517,N_16657);
or U25954 (N_25954,N_10720,N_13581);
or U25955 (N_25955,N_11978,N_17738);
or U25956 (N_25956,N_18792,N_18099);
and U25957 (N_25957,N_17509,N_15181);
or U25958 (N_25958,N_17945,N_11713);
or U25959 (N_25959,N_13372,N_14620);
nand U25960 (N_25960,N_14551,N_18371);
and U25961 (N_25961,N_15397,N_13029);
nand U25962 (N_25962,N_14584,N_18415);
nor U25963 (N_25963,N_10969,N_15726);
nand U25964 (N_25964,N_10040,N_18352);
or U25965 (N_25965,N_19832,N_16293);
nor U25966 (N_25966,N_14159,N_17044);
nor U25967 (N_25967,N_13020,N_11102);
nand U25968 (N_25968,N_10255,N_13768);
and U25969 (N_25969,N_10833,N_11984);
and U25970 (N_25970,N_15060,N_18009);
nor U25971 (N_25971,N_12302,N_18510);
or U25972 (N_25972,N_10260,N_15655);
or U25973 (N_25973,N_18500,N_14554);
nor U25974 (N_25974,N_12010,N_10025);
or U25975 (N_25975,N_13080,N_15016);
and U25976 (N_25976,N_19547,N_15015);
and U25977 (N_25977,N_18833,N_18759);
nand U25978 (N_25978,N_18795,N_11893);
nand U25979 (N_25979,N_11045,N_13462);
nor U25980 (N_25980,N_17931,N_12803);
and U25981 (N_25981,N_17768,N_19075);
nand U25982 (N_25982,N_13140,N_14666);
and U25983 (N_25983,N_11953,N_11569);
and U25984 (N_25984,N_11698,N_11015);
nor U25985 (N_25985,N_19826,N_18468);
nand U25986 (N_25986,N_16020,N_16985);
and U25987 (N_25987,N_13606,N_10290);
and U25988 (N_25988,N_18790,N_11358);
nand U25989 (N_25989,N_17803,N_17584);
or U25990 (N_25990,N_16264,N_12280);
and U25991 (N_25991,N_16930,N_14899);
nor U25992 (N_25992,N_17406,N_15307);
nand U25993 (N_25993,N_18859,N_15811);
or U25994 (N_25994,N_19091,N_17184);
or U25995 (N_25995,N_10721,N_13925);
and U25996 (N_25996,N_11058,N_19242);
nor U25997 (N_25997,N_15445,N_17488);
xor U25998 (N_25998,N_13396,N_14534);
and U25999 (N_25999,N_15732,N_19242);
nand U26000 (N_26000,N_18709,N_13448);
nand U26001 (N_26001,N_16226,N_14050);
nand U26002 (N_26002,N_10937,N_11538);
or U26003 (N_26003,N_19394,N_16283);
and U26004 (N_26004,N_16962,N_13756);
nor U26005 (N_26005,N_11235,N_19237);
nor U26006 (N_26006,N_14207,N_18517);
or U26007 (N_26007,N_15453,N_18815);
or U26008 (N_26008,N_19361,N_13884);
nand U26009 (N_26009,N_19064,N_18785);
or U26010 (N_26010,N_16863,N_10340);
or U26011 (N_26011,N_16886,N_19180);
nand U26012 (N_26012,N_16644,N_14576);
nor U26013 (N_26013,N_12884,N_13374);
nand U26014 (N_26014,N_14519,N_17985);
nand U26015 (N_26015,N_18111,N_11081);
nor U26016 (N_26016,N_12203,N_11098);
nor U26017 (N_26017,N_11321,N_13991);
and U26018 (N_26018,N_19546,N_13377);
nor U26019 (N_26019,N_13342,N_19652);
nor U26020 (N_26020,N_17120,N_13297);
or U26021 (N_26021,N_15193,N_10125);
and U26022 (N_26022,N_15858,N_11634);
or U26023 (N_26023,N_13716,N_14454);
or U26024 (N_26024,N_18330,N_10543);
nor U26025 (N_26025,N_16420,N_18990);
nor U26026 (N_26026,N_17945,N_17518);
and U26027 (N_26027,N_11516,N_18607);
and U26028 (N_26028,N_16418,N_19338);
nand U26029 (N_26029,N_12637,N_19233);
nor U26030 (N_26030,N_12314,N_18544);
nor U26031 (N_26031,N_10337,N_14611);
and U26032 (N_26032,N_13411,N_14357);
and U26033 (N_26033,N_17640,N_16448);
nor U26034 (N_26034,N_11893,N_19572);
nand U26035 (N_26035,N_13000,N_14439);
nor U26036 (N_26036,N_19481,N_13951);
nor U26037 (N_26037,N_12796,N_17484);
and U26038 (N_26038,N_13639,N_14502);
nand U26039 (N_26039,N_12179,N_12996);
or U26040 (N_26040,N_15618,N_12341);
nand U26041 (N_26041,N_17013,N_12463);
and U26042 (N_26042,N_15962,N_13556);
nand U26043 (N_26043,N_17593,N_18541);
nand U26044 (N_26044,N_14285,N_14115);
or U26045 (N_26045,N_16411,N_16921);
and U26046 (N_26046,N_19932,N_18121);
nand U26047 (N_26047,N_12856,N_13104);
nand U26048 (N_26048,N_11107,N_17951);
or U26049 (N_26049,N_13446,N_17187);
and U26050 (N_26050,N_13534,N_13833);
and U26051 (N_26051,N_17769,N_11841);
and U26052 (N_26052,N_17210,N_16704);
nand U26053 (N_26053,N_17196,N_10886);
nor U26054 (N_26054,N_13064,N_19042);
nor U26055 (N_26055,N_17752,N_10809);
or U26056 (N_26056,N_16978,N_10707);
nand U26057 (N_26057,N_18919,N_17459);
or U26058 (N_26058,N_19350,N_13701);
or U26059 (N_26059,N_12379,N_16216);
and U26060 (N_26060,N_14913,N_17184);
and U26061 (N_26061,N_16514,N_11602);
and U26062 (N_26062,N_17225,N_19664);
or U26063 (N_26063,N_10181,N_15150);
and U26064 (N_26064,N_16609,N_12444);
or U26065 (N_26065,N_15137,N_13715);
or U26066 (N_26066,N_15161,N_10776);
nand U26067 (N_26067,N_17865,N_19389);
nand U26068 (N_26068,N_14778,N_12425);
nand U26069 (N_26069,N_15360,N_16710);
or U26070 (N_26070,N_11140,N_10224);
or U26071 (N_26071,N_15468,N_18509);
nand U26072 (N_26072,N_18797,N_17294);
or U26073 (N_26073,N_18740,N_10955);
or U26074 (N_26074,N_15003,N_18805);
nand U26075 (N_26075,N_19158,N_10240);
nor U26076 (N_26076,N_13090,N_11871);
nor U26077 (N_26077,N_19533,N_17690);
and U26078 (N_26078,N_13330,N_14250);
nand U26079 (N_26079,N_15430,N_11423);
nand U26080 (N_26080,N_12860,N_16847);
nor U26081 (N_26081,N_12006,N_19561);
nand U26082 (N_26082,N_16492,N_15375);
and U26083 (N_26083,N_14781,N_13478);
nor U26084 (N_26084,N_13503,N_12696);
or U26085 (N_26085,N_18858,N_12652);
and U26086 (N_26086,N_16220,N_14036);
and U26087 (N_26087,N_13079,N_10354);
and U26088 (N_26088,N_15059,N_12594);
xor U26089 (N_26089,N_16023,N_17099);
nand U26090 (N_26090,N_19707,N_11296);
and U26091 (N_26091,N_17221,N_13890);
and U26092 (N_26092,N_15780,N_11276);
or U26093 (N_26093,N_14031,N_12631);
nor U26094 (N_26094,N_16357,N_12033);
and U26095 (N_26095,N_18066,N_18875);
nand U26096 (N_26096,N_11071,N_13019);
and U26097 (N_26097,N_19134,N_11428);
nor U26098 (N_26098,N_17976,N_16532);
nand U26099 (N_26099,N_11920,N_15648);
nor U26100 (N_26100,N_18599,N_19123);
nand U26101 (N_26101,N_13704,N_14412);
nor U26102 (N_26102,N_17045,N_15388);
or U26103 (N_26103,N_14619,N_15571);
and U26104 (N_26104,N_10154,N_19852);
and U26105 (N_26105,N_17401,N_16672);
nand U26106 (N_26106,N_17583,N_12894);
and U26107 (N_26107,N_19481,N_12207);
and U26108 (N_26108,N_13757,N_19509);
nor U26109 (N_26109,N_18577,N_19547);
nor U26110 (N_26110,N_12924,N_17057);
and U26111 (N_26111,N_13102,N_18674);
or U26112 (N_26112,N_13633,N_18031);
and U26113 (N_26113,N_13266,N_15818);
nor U26114 (N_26114,N_15830,N_10504);
nor U26115 (N_26115,N_18239,N_12007);
or U26116 (N_26116,N_19230,N_11677);
nor U26117 (N_26117,N_19841,N_19012);
or U26118 (N_26118,N_14184,N_14318);
and U26119 (N_26119,N_13951,N_13827);
and U26120 (N_26120,N_15900,N_12330);
nor U26121 (N_26121,N_18043,N_10981);
or U26122 (N_26122,N_11616,N_10015);
xnor U26123 (N_26123,N_16430,N_14645);
and U26124 (N_26124,N_16535,N_19806);
nand U26125 (N_26125,N_12961,N_16530);
and U26126 (N_26126,N_16678,N_11547);
nor U26127 (N_26127,N_18046,N_12195);
or U26128 (N_26128,N_15017,N_11057);
nand U26129 (N_26129,N_16762,N_12344);
or U26130 (N_26130,N_12236,N_17678);
nand U26131 (N_26131,N_12541,N_12087);
or U26132 (N_26132,N_18415,N_11644);
nor U26133 (N_26133,N_16104,N_19832);
and U26134 (N_26134,N_16403,N_12414);
or U26135 (N_26135,N_17467,N_10221);
nor U26136 (N_26136,N_17975,N_16794);
and U26137 (N_26137,N_12599,N_12201);
nor U26138 (N_26138,N_18257,N_18905);
or U26139 (N_26139,N_14685,N_12764);
nand U26140 (N_26140,N_16872,N_15948);
and U26141 (N_26141,N_17694,N_15605);
or U26142 (N_26142,N_10764,N_12398);
nand U26143 (N_26143,N_17502,N_15972);
nor U26144 (N_26144,N_19085,N_14004);
nand U26145 (N_26145,N_12349,N_10738);
nor U26146 (N_26146,N_13191,N_12432);
xor U26147 (N_26147,N_12411,N_13747);
nor U26148 (N_26148,N_19616,N_11291);
nand U26149 (N_26149,N_18874,N_17316);
nor U26150 (N_26150,N_16399,N_12115);
or U26151 (N_26151,N_18399,N_17580);
or U26152 (N_26152,N_14460,N_11179);
and U26153 (N_26153,N_18420,N_10951);
nor U26154 (N_26154,N_15476,N_13487);
nand U26155 (N_26155,N_15473,N_14955);
and U26156 (N_26156,N_14472,N_12888);
nand U26157 (N_26157,N_16980,N_13929);
or U26158 (N_26158,N_10238,N_13395);
and U26159 (N_26159,N_10321,N_12233);
nor U26160 (N_26160,N_12480,N_17981);
nor U26161 (N_26161,N_16957,N_19069);
and U26162 (N_26162,N_11888,N_16959);
nand U26163 (N_26163,N_14031,N_18688);
nor U26164 (N_26164,N_11509,N_12169);
and U26165 (N_26165,N_19147,N_16911);
or U26166 (N_26166,N_11068,N_10066);
nor U26167 (N_26167,N_16596,N_19375);
and U26168 (N_26168,N_18316,N_11534);
or U26169 (N_26169,N_10591,N_11234);
xor U26170 (N_26170,N_16473,N_10809);
nor U26171 (N_26171,N_14938,N_16033);
and U26172 (N_26172,N_19915,N_11559);
nor U26173 (N_26173,N_10376,N_19941);
nor U26174 (N_26174,N_18807,N_13284);
nand U26175 (N_26175,N_18867,N_12712);
nor U26176 (N_26176,N_15650,N_17265);
and U26177 (N_26177,N_18222,N_12347);
nor U26178 (N_26178,N_14694,N_13610);
nor U26179 (N_26179,N_18516,N_15140);
nor U26180 (N_26180,N_11826,N_18921);
or U26181 (N_26181,N_14343,N_16144);
and U26182 (N_26182,N_17108,N_15990);
nand U26183 (N_26183,N_18886,N_16617);
and U26184 (N_26184,N_14204,N_14982);
nand U26185 (N_26185,N_11251,N_15661);
nor U26186 (N_26186,N_10518,N_15026);
nor U26187 (N_26187,N_18507,N_19894);
and U26188 (N_26188,N_11751,N_19174);
or U26189 (N_26189,N_15315,N_10590);
nand U26190 (N_26190,N_11682,N_10218);
or U26191 (N_26191,N_17293,N_13460);
or U26192 (N_26192,N_11810,N_14437);
nor U26193 (N_26193,N_13835,N_15086);
and U26194 (N_26194,N_19961,N_13751);
nand U26195 (N_26195,N_18126,N_10884);
nor U26196 (N_26196,N_13553,N_15849);
or U26197 (N_26197,N_18276,N_14660);
nand U26198 (N_26198,N_16756,N_18285);
and U26199 (N_26199,N_10961,N_17908);
nor U26200 (N_26200,N_16027,N_16542);
or U26201 (N_26201,N_18387,N_18576);
or U26202 (N_26202,N_17358,N_15991);
and U26203 (N_26203,N_19928,N_19710);
nand U26204 (N_26204,N_14924,N_13348);
nand U26205 (N_26205,N_18048,N_14092);
and U26206 (N_26206,N_13592,N_10121);
and U26207 (N_26207,N_11307,N_14366);
nand U26208 (N_26208,N_10793,N_14563);
and U26209 (N_26209,N_18563,N_14174);
nand U26210 (N_26210,N_11619,N_12143);
nor U26211 (N_26211,N_12376,N_19208);
or U26212 (N_26212,N_10917,N_19054);
nor U26213 (N_26213,N_18660,N_14298);
nand U26214 (N_26214,N_10894,N_11227);
nand U26215 (N_26215,N_15483,N_17176);
nand U26216 (N_26216,N_12879,N_10173);
nand U26217 (N_26217,N_15834,N_12757);
nor U26218 (N_26218,N_15765,N_11865);
and U26219 (N_26219,N_13366,N_12914);
and U26220 (N_26220,N_11138,N_19224);
and U26221 (N_26221,N_12984,N_11208);
nor U26222 (N_26222,N_11365,N_13531);
nor U26223 (N_26223,N_16045,N_16398);
and U26224 (N_26224,N_12694,N_16691);
nor U26225 (N_26225,N_16396,N_11736);
and U26226 (N_26226,N_10151,N_18217);
and U26227 (N_26227,N_13473,N_13816);
and U26228 (N_26228,N_19089,N_12118);
nor U26229 (N_26229,N_13048,N_18560);
nor U26230 (N_26230,N_16015,N_17714);
nand U26231 (N_26231,N_16020,N_17031);
and U26232 (N_26232,N_17906,N_18997);
or U26233 (N_26233,N_11249,N_17718);
nand U26234 (N_26234,N_19086,N_18986);
nor U26235 (N_26235,N_15955,N_15517);
or U26236 (N_26236,N_11127,N_10292);
or U26237 (N_26237,N_18214,N_15328);
or U26238 (N_26238,N_12608,N_16563);
and U26239 (N_26239,N_13877,N_19934);
or U26240 (N_26240,N_10869,N_14735);
or U26241 (N_26241,N_19216,N_12912);
nor U26242 (N_26242,N_16240,N_17200);
nand U26243 (N_26243,N_11060,N_10983);
nand U26244 (N_26244,N_13276,N_15110);
nor U26245 (N_26245,N_15330,N_11524);
nor U26246 (N_26246,N_15152,N_17214);
nor U26247 (N_26247,N_10034,N_11130);
or U26248 (N_26248,N_14935,N_12827);
and U26249 (N_26249,N_14984,N_14806);
nor U26250 (N_26250,N_12722,N_15230);
nand U26251 (N_26251,N_12685,N_11403);
nand U26252 (N_26252,N_18424,N_16098);
or U26253 (N_26253,N_19710,N_13543);
nand U26254 (N_26254,N_12745,N_11084);
or U26255 (N_26255,N_16567,N_10895);
nand U26256 (N_26256,N_14859,N_15476);
nor U26257 (N_26257,N_14724,N_14498);
nand U26258 (N_26258,N_11569,N_10674);
nor U26259 (N_26259,N_10639,N_15450);
or U26260 (N_26260,N_14371,N_13099);
or U26261 (N_26261,N_17737,N_11539);
nor U26262 (N_26262,N_17262,N_17805);
nand U26263 (N_26263,N_19098,N_17902);
and U26264 (N_26264,N_11576,N_13063);
nand U26265 (N_26265,N_16683,N_13483);
nand U26266 (N_26266,N_13563,N_16332);
or U26267 (N_26267,N_18237,N_15930);
nor U26268 (N_26268,N_17684,N_10148);
nand U26269 (N_26269,N_19391,N_15810);
nor U26270 (N_26270,N_14800,N_15612);
nand U26271 (N_26271,N_16244,N_11422);
and U26272 (N_26272,N_13818,N_10807);
nand U26273 (N_26273,N_14790,N_18670);
and U26274 (N_26274,N_15904,N_11487);
nand U26275 (N_26275,N_10119,N_19096);
nor U26276 (N_26276,N_19335,N_10805);
and U26277 (N_26277,N_10861,N_16459);
and U26278 (N_26278,N_19051,N_11404);
and U26279 (N_26279,N_10305,N_18956);
or U26280 (N_26280,N_10482,N_12645);
nand U26281 (N_26281,N_13852,N_16176);
nand U26282 (N_26282,N_18680,N_11955);
nand U26283 (N_26283,N_14789,N_11798);
or U26284 (N_26284,N_13522,N_14223);
and U26285 (N_26285,N_19746,N_10454);
nor U26286 (N_26286,N_12116,N_15616);
nand U26287 (N_26287,N_17232,N_14621);
and U26288 (N_26288,N_11655,N_12980);
nand U26289 (N_26289,N_10176,N_14543);
or U26290 (N_26290,N_13982,N_19919);
nand U26291 (N_26291,N_10222,N_15652);
or U26292 (N_26292,N_10175,N_13865);
nand U26293 (N_26293,N_11895,N_11911);
nand U26294 (N_26294,N_18048,N_13615);
nand U26295 (N_26295,N_16623,N_13873);
and U26296 (N_26296,N_13306,N_13841);
nor U26297 (N_26297,N_16296,N_10747);
or U26298 (N_26298,N_11401,N_10049);
or U26299 (N_26299,N_17180,N_10934);
nor U26300 (N_26300,N_11041,N_15548);
and U26301 (N_26301,N_16718,N_10437);
and U26302 (N_26302,N_10222,N_19423);
or U26303 (N_26303,N_12824,N_14268);
and U26304 (N_26304,N_13647,N_14413);
nor U26305 (N_26305,N_15802,N_13254);
and U26306 (N_26306,N_13738,N_17168);
and U26307 (N_26307,N_16324,N_15430);
and U26308 (N_26308,N_14693,N_16770);
nand U26309 (N_26309,N_15449,N_11896);
nand U26310 (N_26310,N_16854,N_14069);
nand U26311 (N_26311,N_19341,N_18433);
or U26312 (N_26312,N_14597,N_13346);
nand U26313 (N_26313,N_19283,N_17267);
nor U26314 (N_26314,N_15068,N_18361);
and U26315 (N_26315,N_14545,N_13910);
or U26316 (N_26316,N_16740,N_14352);
and U26317 (N_26317,N_18083,N_19445);
and U26318 (N_26318,N_17767,N_15592);
nand U26319 (N_26319,N_19680,N_18825);
nand U26320 (N_26320,N_16835,N_13208);
and U26321 (N_26321,N_10531,N_12763);
and U26322 (N_26322,N_17285,N_16665);
or U26323 (N_26323,N_15134,N_10032);
or U26324 (N_26324,N_15950,N_12888);
or U26325 (N_26325,N_13648,N_10389);
or U26326 (N_26326,N_14492,N_14487);
and U26327 (N_26327,N_15199,N_17625);
nor U26328 (N_26328,N_19017,N_16719);
nor U26329 (N_26329,N_17850,N_19689);
nand U26330 (N_26330,N_13426,N_19722);
or U26331 (N_26331,N_10564,N_12410);
nor U26332 (N_26332,N_11652,N_18083);
nand U26333 (N_26333,N_12584,N_14608);
xnor U26334 (N_26334,N_16437,N_10867);
or U26335 (N_26335,N_17636,N_19181);
or U26336 (N_26336,N_13240,N_16751);
or U26337 (N_26337,N_17394,N_15876);
or U26338 (N_26338,N_18350,N_18460);
nor U26339 (N_26339,N_18103,N_13342);
or U26340 (N_26340,N_10107,N_14140);
nand U26341 (N_26341,N_19992,N_18508);
nand U26342 (N_26342,N_18147,N_14636);
and U26343 (N_26343,N_14138,N_17371);
and U26344 (N_26344,N_11344,N_14201);
and U26345 (N_26345,N_10110,N_14071);
nor U26346 (N_26346,N_15457,N_12085);
xor U26347 (N_26347,N_17804,N_12970);
and U26348 (N_26348,N_11536,N_13351);
nand U26349 (N_26349,N_10455,N_18946);
or U26350 (N_26350,N_17426,N_12944);
or U26351 (N_26351,N_13245,N_14823);
nand U26352 (N_26352,N_10098,N_16724);
nor U26353 (N_26353,N_18386,N_10428);
or U26354 (N_26354,N_16745,N_10894);
nor U26355 (N_26355,N_10692,N_12249);
nor U26356 (N_26356,N_17512,N_17682);
nand U26357 (N_26357,N_12431,N_18991);
nand U26358 (N_26358,N_18993,N_13568);
nor U26359 (N_26359,N_10871,N_13409);
nor U26360 (N_26360,N_19871,N_11465);
or U26361 (N_26361,N_15086,N_14832);
nor U26362 (N_26362,N_15216,N_17459);
nand U26363 (N_26363,N_18006,N_11781);
nand U26364 (N_26364,N_19825,N_15947);
and U26365 (N_26365,N_18056,N_19906);
or U26366 (N_26366,N_12319,N_18684);
nand U26367 (N_26367,N_18267,N_10794);
xnor U26368 (N_26368,N_14666,N_17642);
and U26369 (N_26369,N_13110,N_18781);
nand U26370 (N_26370,N_13858,N_15888);
nor U26371 (N_26371,N_18833,N_15310);
nor U26372 (N_26372,N_14166,N_16240);
or U26373 (N_26373,N_11256,N_12889);
or U26374 (N_26374,N_19825,N_11123);
or U26375 (N_26375,N_13936,N_13423);
and U26376 (N_26376,N_11997,N_14229);
and U26377 (N_26377,N_11704,N_15349);
or U26378 (N_26378,N_12935,N_17129);
nor U26379 (N_26379,N_11315,N_12271);
and U26380 (N_26380,N_12155,N_14123);
nor U26381 (N_26381,N_17445,N_19613);
and U26382 (N_26382,N_16274,N_15758);
or U26383 (N_26383,N_12707,N_10850);
and U26384 (N_26384,N_13316,N_16804);
nand U26385 (N_26385,N_13098,N_13631);
and U26386 (N_26386,N_17533,N_14777);
and U26387 (N_26387,N_14749,N_19015);
or U26388 (N_26388,N_13691,N_15166);
and U26389 (N_26389,N_13338,N_16081);
and U26390 (N_26390,N_14694,N_15127);
and U26391 (N_26391,N_19773,N_17925);
and U26392 (N_26392,N_17829,N_17405);
and U26393 (N_26393,N_14924,N_17242);
nand U26394 (N_26394,N_12842,N_11466);
nand U26395 (N_26395,N_15699,N_10260);
nor U26396 (N_26396,N_12903,N_16120);
nor U26397 (N_26397,N_13063,N_14991);
or U26398 (N_26398,N_12608,N_10991);
or U26399 (N_26399,N_13467,N_14129);
and U26400 (N_26400,N_17876,N_13467);
or U26401 (N_26401,N_10780,N_12100);
nor U26402 (N_26402,N_16274,N_19302);
and U26403 (N_26403,N_12125,N_17587);
nand U26404 (N_26404,N_10025,N_11221);
nand U26405 (N_26405,N_19273,N_15545);
or U26406 (N_26406,N_16339,N_17850);
or U26407 (N_26407,N_18292,N_18869);
and U26408 (N_26408,N_16727,N_16477);
or U26409 (N_26409,N_10931,N_13765);
or U26410 (N_26410,N_16833,N_13174);
and U26411 (N_26411,N_10948,N_17648);
nor U26412 (N_26412,N_12678,N_16497);
and U26413 (N_26413,N_17397,N_15036);
or U26414 (N_26414,N_12619,N_10752);
and U26415 (N_26415,N_17680,N_13288);
and U26416 (N_26416,N_18078,N_14279);
nand U26417 (N_26417,N_18951,N_18216);
nor U26418 (N_26418,N_14534,N_18633);
nand U26419 (N_26419,N_12904,N_12847);
nand U26420 (N_26420,N_14338,N_17150);
nor U26421 (N_26421,N_18165,N_12606);
nor U26422 (N_26422,N_13708,N_19514);
nand U26423 (N_26423,N_18937,N_11717);
and U26424 (N_26424,N_14388,N_18851);
and U26425 (N_26425,N_19802,N_16512);
nand U26426 (N_26426,N_10428,N_17398);
or U26427 (N_26427,N_18365,N_13762);
or U26428 (N_26428,N_13727,N_15030);
and U26429 (N_26429,N_14125,N_19899);
or U26430 (N_26430,N_10632,N_15172);
and U26431 (N_26431,N_10229,N_12988);
xnor U26432 (N_26432,N_14950,N_12244);
nor U26433 (N_26433,N_15861,N_11734);
and U26434 (N_26434,N_15773,N_18211);
or U26435 (N_26435,N_18767,N_13573);
or U26436 (N_26436,N_16594,N_12968);
nor U26437 (N_26437,N_13779,N_17295);
nor U26438 (N_26438,N_15217,N_17902);
nor U26439 (N_26439,N_13076,N_16519);
nor U26440 (N_26440,N_12144,N_13418);
or U26441 (N_26441,N_11339,N_16323);
and U26442 (N_26442,N_19772,N_18125);
or U26443 (N_26443,N_11132,N_15727);
nand U26444 (N_26444,N_19267,N_13806);
or U26445 (N_26445,N_16689,N_17076);
and U26446 (N_26446,N_16223,N_16231);
or U26447 (N_26447,N_10380,N_15546);
and U26448 (N_26448,N_19733,N_19904);
and U26449 (N_26449,N_17851,N_15415);
nand U26450 (N_26450,N_10061,N_12870);
and U26451 (N_26451,N_12319,N_12911);
nor U26452 (N_26452,N_18542,N_13030);
nor U26453 (N_26453,N_14913,N_19247);
or U26454 (N_26454,N_12603,N_14949);
nand U26455 (N_26455,N_17920,N_19285);
or U26456 (N_26456,N_15908,N_18667);
nor U26457 (N_26457,N_14749,N_18859);
and U26458 (N_26458,N_11525,N_18165);
nor U26459 (N_26459,N_13060,N_10981);
and U26460 (N_26460,N_14622,N_14549);
nand U26461 (N_26461,N_12483,N_12100);
xor U26462 (N_26462,N_18560,N_14757);
nor U26463 (N_26463,N_12385,N_14981);
nand U26464 (N_26464,N_11065,N_13580);
nand U26465 (N_26465,N_15909,N_16580);
nand U26466 (N_26466,N_17399,N_17737);
nor U26467 (N_26467,N_16007,N_16178);
and U26468 (N_26468,N_14639,N_11005);
nand U26469 (N_26469,N_10395,N_19213);
nand U26470 (N_26470,N_18906,N_15025);
and U26471 (N_26471,N_15574,N_19192);
nor U26472 (N_26472,N_18089,N_17724);
and U26473 (N_26473,N_10858,N_16631);
nand U26474 (N_26474,N_12837,N_16543);
or U26475 (N_26475,N_19827,N_14587);
and U26476 (N_26476,N_12813,N_16045);
nor U26477 (N_26477,N_11040,N_15628);
xor U26478 (N_26478,N_18886,N_13421);
or U26479 (N_26479,N_18595,N_14286);
and U26480 (N_26480,N_13356,N_15309);
and U26481 (N_26481,N_15392,N_10433);
or U26482 (N_26482,N_16731,N_16880);
and U26483 (N_26483,N_15530,N_16961);
or U26484 (N_26484,N_18989,N_13424);
and U26485 (N_26485,N_17524,N_17943);
nor U26486 (N_26486,N_11766,N_17477);
nor U26487 (N_26487,N_10743,N_10735);
and U26488 (N_26488,N_16174,N_11189);
and U26489 (N_26489,N_19077,N_19982);
and U26490 (N_26490,N_16337,N_19927);
and U26491 (N_26491,N_19261,N_19386);
nor U26492 (N_26492,N_15576,N_17597);
nand U26493 (N_26493,N_19721,N_17128);
nor U26494 (N_26494,N_16223,N_14249);
nor U26495 (N_26495,N_13170,N_17320);
or U26496 (N_26496,N_16385,N_17746);
nor U26497 (N_26497,N_10738,N_16466);
and U26498 (N_26498,N_18283,N_16575);
nand U26499 (N_26499,N_18207,N_17500);
or U26500 (N_26500,N_11588,N_10971);
xnor U26501 (N_26501,N_13659,N_15386);
nor U26502 (N_26502,N_10540,N_15249);
nor U26503 (N_26503,N_18312,N_10928);
nor U26504 (N_26504,N_15949,N_19032);
nand U26505 (N_26505,N_16419,N_18571);
nand U26506 (N_26506,N_10149,N_18899);
nand U26507 (N_26507,N_15111,N_16172);
and U26508 (N_26508,N_11624,N_12322);
and U26509 (N_26509,N_11817,N_12394);
and U26510 (N_26510,N_10091,N_17016);
nand U26511 (N_26511,N_15927,N_16644);
and U26512 (N_26512,N_17758,N_16459);
or U26513 (N_26513,N_15595,N_17958);
and U26514 (N_26514,N_15052,N_17865);
nor U26515 (N_26515,N_19087,N_14903);
or U26516 (N_26516,N_17508,N_17539);
and U26517 (N_26517,N_18131,N_12617);
xor U26518 (N_26518,N_12470,N_19881);
nand U26519 (N_26519,N_16395,N_18350);
or U26520 (N_26520,N_15105,N_13824);
and U26521 (N_26521,N_14114,N_17143);
nor U26522 (N_26522,N_14911,N_11244);
nor U26523 (N_26523,N_17512,N_15405);
or U26524 (N_26524,N_13019,N_12980);
nor U26525 (N_26525,N_11616,N_11878);
or U26526 (N_26526,N_10634,N_10638);
or U26527 (N_26527,N_19155,N_13949);
nand U26528 (N_26528,N_17086,N_11952);
nand U26529 (N_26529,N_10843,N_14710);
or U26530 (N_26530,N_11336,N_17405);
nor U26531 (N_26531,N_17198,N_11264);
and U26532 (N_26532,N_11909,N_13713);
or U26533 (N_26533,N_19677,N_15133);
and U26534 (N_26534,N_19059,N_12012);
nand U26535 (N_26535,N_14988,N_12198);
nand U26536 (N_26536,N_16251,N_10721);
nor U26537 (N_26537,N_19578,N_13939);
or U26538 (N_26538,N_18487,N_15525);
or U26539 (N_26539,N_13538,N_14351);
nand U26540 (N_26540,N_10026,N_16398);
or U26541 (N_26541,N_16537,N_12639);
and U26542 (N_26542,N_19265,N_15044);
nor U26543 (N_26543,N_13957,N_15646);
or U26544 (N_26544,N_19481,N_13195);
nand U26545 (N_26545,N_17963,N_18457);
and U26546 (N_26546,N_18788,N_16582);
or U26547 (N_26547,N_19702,N_17715);
nor U26548 (N_26548,N_17758,N_10202);
nand U26549 (N_26549,N_17421,N_13704);
nor U26550 (N_26550,N_17977,N_16424);
nor U26551 (N_26551,N_11330,N_15863);
nor U26552 (N_26552,N_17677,N_15009);
and U26553 (N_26553,N_10980,N_18733);
or U26554 (N_26554,N_11212,N_10869);
nand U26555 (N_26555,N_19930,N_12422);
or U26556 (N_26556,N_14779,N_19857);
nor U26557 (N_26557,N_11460,N_12948);
or U26558 (N_26558,N_14520,N_19800);
and U26559 (N_26559,N_12821,N_13052);
and U26560 (N_26560,N_10886,N_15075);
nand U26561 (N_26561,N_12490,N_12106);
or U26562 (N_26562,N_13830,N_15270);
nor U26563 (N_26563,N_14619,N_12207);
and U26564 (N_26564,N_10109,N_19358);
or U26565 (N_26565,N_14341,N_11717);
nor U26566 (N_26566,N_11179,N_15871);
nor U26567 (N_26567,N_10001,N_14962);
nor U26568 (N_26568,N_19567,N_13660);
nor U26569 (N_26569,N_11167,N_13788);
or U26570 (N_26570,N_16923,N_18454);
nor U26571 (N_26571,N_19758,N_18860);
nor U26572 (N_26572,N_12077,N_12794);
nor U26573 (N_26573,N_12390,N_17549);
and U26574 (N_26574,N_10372,N_18421);
and U26575 (N_26575,N_17043,N_18810);
and U26576 (N_26576,N_10503,N_17345);
and U26577 (N_26577,N_10450,N_13536);
nor U26578 (N_26578,N_19871,N_16185);
nand U26579 (N_26579,N_13834,N_12927);
or U26580 (N_26580,N_18698,N_14257);
nor U26581 (N_26581,N_13560,N_17906);
or U26582 (N_26582,N_17230,N_10799);
nand U26583 (N_26583,N_11058,N_18580);
nand U26584 (N_26584,N_17560,N_12458);
nor U26585 (N_26585,N_18317,N_16737);
nand U26586 (N_26586,N_18685,N_18417);
or U26587 (N_26587,N_10815,N_19020);
or U26588 (N_26588,N_17163,N_14270);
nand U26589 (N_26589,N_16406,N_18587);
and U26590 (N_26590,N_17675,N_19633);
nand U26591 (N_26591,N_14368,N_10451);
nand U26592 (N_26592,N_18329,N_14310);
or U26593 (N_26593,N_15152,N_13816);
and U26594 (N_26594,N_13585,N_18661);
nor U26595 (N_26595,N_11960,N_18695);
or U26596 (N_26596,N_10740,N_18129);
nand U26597 (N_26597,N_16792,N_14186);
nand U26598 (N_26598,N_11516,N_19636);
nand U26599 (N_26599,N_13318,N_18522);
or U26600 (N_26600,N_19288,N_19949);
nor U26601 (N_26601,N_12947,N_15451);
or U26602 (N_26602,N_18299,N_11340);
nor U26603 (N_26603,N_17900,N_18667);
nor U26604 (N_26604,N_11859,N_15381);
nand U26605 (N_26605,N_18920,N_17852);
or U26606 (N_26606,N_16351,N_11755);
nor U26607 (N_26607,N_10728,N_11571);
or U26608 (N_26608,N_13166,N_16351);
nor U26609 (N_26609,N_17277,N_16633);
or U26610 (N_26610,N_12429,N_19403);
nand U26611 (N_26611,N_16543,N_15564);
nand U26612 (N_26612,N_14684,N_14338);
and U26613 (N_26613,N_10530,N_19141);
nand U26614 (N_26614,N_16960,N_13485);
and U26615 (N_26615,N_17273,N_19188);
xnor U26616 (N_26616,N_17781,N_19177);
or U26617 (N_26617,N_11959,N_19088);
nand U26618 (N_26618,N_17459,N_13114);
nand U26619 (N_26619,N_13559,N_13173);
or U26620 (N_26620,N_10940,N_15281);
nand U26621 (N_26621,N_16219,N_17034);
nand U26622 (N_26622,N_16453,N_16510);
and U26623 (N_26623,N_12271,N_17555);
nand U26624 (N_26624,N_10691,N_17494);
nor U26625 (N_26625,N_14068,N_18495);
or U26626 (N_26626,N_12873,N_14268);
and U26627 (N_26627,N_10938,N_16229);
nor U26628 (N_26628,N_15352,N_17202);
nor U26629 (N_26629,N_13691,N_16547);
nand U26630 (N_26630,N_12997,N_15300);
or U26631 (N_26631,N_18246,N_10635);
nor U26632 (N_26632,N_10650,N_13477);
and U26633 (N_26633,N_11140,N_13012);
or U26634 (N_26634,N_14494,N_17420);
or U26635 (N_26635,N_18464,N_12446);
and U26636 (N_26636,N_17701,N_19902);
nand U26637 (N_26637,N_15762,N_15419);
or U26638 (N_26638,N_15167,N_18822);
or U26639 (N_26639,N_13777,N_18228);
nand U26640 (N_26640,N_10940,N_16031);
or U26641 (N_26641,N_17691,N_10847);
nand U26642 (N_26642,N_10143,N_10130);
and U26643 (N_26643,N_19564,N_10211);
nor U26644 (N_26644,N_15908,N_15697);
and U26645 (N_26645,N_10524,N_13652);
nand U26646 (N_26646,N_18485,N_14438);
or U26647 (N_26647,N_10563,N_13814);
and U26648 (N_26648,N_11074,N_17276);
nand U26649 (N_26649,N_12713,N_10231);
nand U26650 (N_26650,N_11948,N_19283);
and U26651 (N_26651,N_10706,N_11351);
nor U26652 (N_26652,N_16990,N_15455);
nor U26653 (N_26653,N_12059,N_15710);
nor U26654 (N_26654,N_12309,N_15437);
or U26655 (N_26655,N_18130,N_15911);
and U26656 (N_26656,N_14845,N_13243);
or U26657 (N_26657,N_13973,N_19962);
or U26658 (N_26658,N_13258,N_14801);
and U26659 (N_26659,N_10927,N_10329);
nor U26660 (N_26660,N_13845,N_18191);
nor U26661 (N_26661,N_19709,N_19296);
nand U26662 (N_26662,N_12659,N_18581);
nor U26663 (N_26663,N_12851,N_10529);
nor U26664 (N_26664,N_17436,N_15050);
nand U26665 (N_26665,N_19676,N_10825);
or U26666 (N_26666,N_13124,N_19561);
nand U26667 (N_26667,N_17059,N_16764);
or U26668 (N_26668,N_19049,N_12127);
or U26669 (N_26669,N_12057,N_13210);
or U26670 (N_26670,N_13011,N_12179);
nor U26671 (N_26671,N_13558,N_17324);
nand U26672 (N_26672,N_11596,N_19571);
nor U26673 (N_26673,N_15617,N_17922);
or U26674 (N_26674,N_11872,N_14036);
or U26675 (N_26675,N_11086,N_13066);
nand U26676 (N_26676,N_16860,N_13080);
nor U26677 (N_26677,N_16318,N_10008);
and U26678 (N_26678,N_16240,N_14418);
nand U26679 (N_26679,N_15728,N_10863);
nor U26680 (N_26680,N_15356,N_19453);
nor U26681 (N_26681,N_10646,N_13589);
and U26682 (N_26682,N_14040,N_11121);
and U26683 (N_26683,N_17126,N_17961);
or U26684 (N_26684,N_14009,N_12683);
nor U26685 (N_26685,N_15445,N_12609);
or U26686 (N_26686,N_14856,N_14650);
nor U26687 (N_26687,N_18878,N_15336);
and U26688 (N_26688,N_16565,N_14657);
or U26689 (N_26689,N_12933,N_14662);
nor U26690 (N_26690,N_18627,N_19920);
nor U26691 (N_26691,N_19016,N_14927);
nor U26692 (N_26692,N_15251,N_13106);
and U26693 (N_26693,N_11540,N_10571);
nor U26694 (N_26694,N_12436,N_18778);
and U26695 (N_26695,N_16115,N_15512);
nor U26696 (N_26696,N_14178,N_11973);
nand U26697 (N_26697,N_11828,N_18351);
and U26698 (N_26698,N_14173,N_16587);
or U26699 (N_26699,N_12431,N_17909);
or U26700 (N_26700,N_12344,N_19377);
nor U26701 (N_26701,N_19999,N_11404);
nand U26702 (N_26702,N_10605,N_16950);
and U26703 (N_26703,N_12549,N_11422);
and U26704 (N_26704,N_12174,N_13762);
and U26705 (N_26705,N_14734,N_18139);
and U26706 (N_26706,N_19801,N_12525);
and U26707 (N_26707,N_12349,N_14195);
xnor U26708 (N_26708,N_14988,N_14417);
nor U26709 (N_26709,N_11584,N_16448);
and U26710 (N_26710,N_19854,N_15647);
nand U26711 (N_26711,N_14536,N_12081);
and U26712 (N_26712,N_10295,N_17409);
nor U26713 (N_26713,N_17062,N_11256);
nor U26714 (N_26714,N_16808,N_19909);
or U26715 (N_26715,N_14986,N_14870);
or U26716 (N_26716,N_19225,N_17150);
nand U26717 (N_26717,N_14176,N_18954);
nand U26718 (N_26718,N_19966,N_11907);
or U26719 (N_26719,N_18007,N_10876);
nor U26720 (N_26720,N_10174,N_16909);
and U26721 (N_26721,N_16807,N_15653);
or U26722 (N_26722,N_12684,N_19018);
and U26723 (N_26723,N_11092,N_15812);
nand U26724 (N_26724,N_19930,N_15819);
nor U26725 (N_26725,N_12411,N_11431);
nand U26726 (N_26726,N_14058,N_16698);
nor U26727 (N_26727,N_18148,N_18363);
or U26728 (N_26728,N_10901,N_19067);
and U26729 (N_26729,N_14104,N_18059);
nor U26730 (N_26730,N_16131,N_14512);
or U26731 (N_26731,N_19933,N_12645);
or U26732 (N_26732,N_16894,N_10833);
and U26733 (N_26733,N_16945,N_13330);
nor U26734 (N_26734,N_13225,N_10180);
or U26735 (N_26735,N_15575,N_11398);
and U26736 (N_26736,N_12151,N_15158);
nand U26737 (N_26737,N_15936,N_16123);
nor U26738 (N_26738,N_14045,N_17383);
or U26739 (N_26739,N_15061,N_16942);
nand U26740 (N_26740,N_11469,N_13445);
or U26741 (N_26741,N_13881,N_16821);
nand U26742 (N_26742,N_15072,N_18031);
nor U26743 (N_26743,N_14680,N_12398);
or U26744 (N_26744,N_16839,N_17001);
and U26745 (N_26745,N_10668,N_16058);
nor U26746 (N_26746,N_17797,N_14829);
or U26747 (N_26747,N_18714,N_11791);
or U26748 (N_26748,N_17589,N_12439);
nor U26749 (N_26749,N_16652,N_15890);
or U26750 (N_26750,N_17462,N_17734);
xor U26751 (N_26751,N_18968,N_13391);
and U26752 (N_26752,N_11908,N_16678);
and U26753 (N_26753,N_16263,N_12512);
nor U26754 (N_26754,N_11700,N_18273);
and U26755 (N_26755,N_19645,N_12679);
and U26756 (N_26756,N_12550,N_17012);
and U26757 (N_26757,N_11690,N_12463);
or U26758 (N_26758,N_14253,N_16654);
nand U26759 (N_26759,N_11768,N_17795);
nor U26760 (N_26760,N_17013,N_17600);
or U26761 (N_26761,N_11530,N_16861);
nand U26762 (N_26762,N_12861,N_18456);
or U26763 (N_26763,N_10608,N_19008);
nand U26764 (N_26764,N_16650,N_16323);
or U26765 (N_26765,N_17691,N_14923);
nor U26766 (N_26766,N_15162,N_14717);
nand U26767 (N_26767,N_18299,N_16754);
nor U26768 (N_26768,N_14620,N_17408);
or U26769 (N_26769,N_15900,N_11727);
nand U26770 (N_26770,N_14359,N_16157);
nor U26771 (N_26771,N_16532,N_13416);
nor U26772 (N_26772,N_18061,N_15994);
nor U26773 (N_26773,N_13900,N_18431);
nand U26774 (N_26774,N_15122,N_13986);
nor U26775 (N_26775,N_17837,N_11867);
nor U26776 (N_26776,N_10822,N_14253);
or U26777 (N_26777,N_13811,N_12543);
and U26778 (N_26778,N_15083,N_12271);
and U26779 (N_26779,N_16557,N_15278);
nand U26780 (N_26780,N_11309,N_18062);
nor U26781 (N_26781,N_19377,N_14155);
or U26782 (N_26782,N_15121,N_11248);
nand U26783 (N_26783,N_12599,N_16427);
nand U26784 (N_26784,N_15529,N_13089);
xor U26785 (N_26785,N_16792,N_19516);
or U26786 (N_26786,N_12542,N_18081);
or U26787 (N_26787,N_15722,N_10858);
or U26788 (N_26788,N_11957,N_15937);
nand U26789 (N_26789,N_13931,N_11704);
nor U26790 (N_26790,N_18371,N_14350);
nor U26791 (N_26791,N_16350,N_13965);
and U26792 (N_26792,N_17157,N_18100);
nand U26793 (N_26793,N_10028,N_19436);
nor U26794 (N_26794,N_17462,N_14213);
or U26795 (N_26795,N_18440,N_18753);
nand U26796 (N_26796,N_11839,N_18473);
or U26797 (N_26797,N_16476,N_13298);
xor U26798 (N_26798,N_10856,N_14717);
nand U26799 (N_26799,N_18982,N_19448);
and U26800 (N_26800,N_11282,N_16061);
and U26801 (N_26801,N_14476,N_18290);
and U26802 (N_26802,N_15985,N_18293);
or U26803 (N_26803,N_15161,N_18744);
nand U26804 (N_26804,N_18114,N_15195);
nand U26805 (N_26805,N_19009,N_14298);
nor U26806 (N_26806,N_13351,N_17041);
nor U26807 (N_26807,N_12116,N_15459);
or U26808 (N_26808,N_18305,N_19563);
nand U26809 (N_26809,N_14761,N_14120);
nor U26810 (N_26810,N_13832,N_17192);
nand U26811 (N_26811,N_12851,N_15048);
nand U26812 (N_26812,N_19412,N_17204);
nor U26813 (N_26813,N_18094,N_15917);
nor U26814 (N_26814,N_10600,N_15031);
and U26815 (N_26815,N_13216,N_15825);
or U26816 (N_26816,N_10220,N_10267);
nand U26817 (N_26817,N_10501,N_13080);
nor U26818 (N_26818,N_14779,N_11584);
or U26819 (N_26819,N_10891,N_10588);
nor U26820 (N_26820,N_19211,N_12914);
nand U26821 (N_26821,N_14586,N_16333);
and U26822 (N_26822,N_12337,N_18448);
nand U26823 (N_26823,N_12489,N_19467);
and U26824 (N_26824,N_12793,N_15899);
nand U26825 (N_26825,N_14409,N_10042);
nand U26826 (N_26826,N_12631,N_11220);
nor U26827 (N_26827,N_16841,N_15422);
nor U26828 (N_26828,N_18746,N_14250);
xnor U26829 (N_26829,N_13101,N_10408);
and U26830 (N_26830,N_15552,N_19329);
or U26831 (N_26831,N_14061,N_16144);
nor U26832 (N_26832,N_19252,N_10037);
or U26833 (N_26833,N_15548,N_19070);
nor U26834 (N_26834,N_11121,N_18383);
nand U26835 (N_26835,N_12546,N_11521);
nand U26836 (N_26836,N_19194,N_14060);
and U26837 (N_26837,N_12485,N_15423);
or U26838 (N_26838,N_15717,N_10327);
and U26839 (N_26839,N_14403,N_10495);
or U26840 (N_26840,N_15876,N_13688);
or U26841 (N_26841,N_15651,N_10516);
or U26842 (N_26842,N_15559,N_12383);
or U26843 (N_26843,N_15234,N_16689);
and U26844 (N_26844,N_16290,N_14970);
nand U26845 (N_26845,N_10474,N_14404);
or U26846 (N_26846,N_14755,N_11098);
or U26847 (N_26847,N_14708,N_17093);
nand U26848 (N_26848,N_16651,N_11153);
and U26849 (N_26849,N_13774,N_18624);
nand U26850 (N_26850,N_16944,N_15029);
and U26851 (N_26851,N_18543,N_16641);
and U26852 (N_26852,N_17593,N_16741);
and U26853 (N_26853,N_17728,N_18743);
and U26854 (N_26854,N_10650,N_13991);
and U26855 (N_26855,N_11435,N_16785);
and U26856 (N_26856,N_19404,N_12819);
or U26857 (N_26857,N_16419,N_18092);
and U26858 (N_26858,N_16901,N_17632);
nand U26859 (N_26859,N_11285,N_18192);
nor U26860 (N_26860,N_15522,N_17487);
or U26861 (N_26861,N_19600,N_15069);
and U26862 (N_26862,N_10033,N_13184);
nand U26863 (N_26863,N_18199,N_16178);
nor U26864 (N_26864,N_17904,N_13571);
nand U26865 (N_26865,N_10214,N_13773);
nand U26866 (N_26866,N_12347,N_17996);
nand U26867 (N_26867,N_13800,N_15832);
and U26868 (N_26868,N_16425,N_12605);
or U26869 (N_26869,N_14117,N_15968);
nand U26870 (N_26870,N_16866,N_11317);
or U26871 (N_26871,N_16279,N_13914);
nor U26872 (N_26872,N_17520,N_17072);
and U26873 (N_26873,N_14335,N_14834);
nor U26874 (N_26874,N_11616,N_11463);
or U26875 (N_26875,N_17869,N_11794);
nand U26876 (N_26876,N_12896,N_15532);
and U26877 (N_26877,N_13194,N_18783);
or U26878 (N_26878,N_10034,N_18259);
nand U26879 (N_26879,N_17395,N_10643);
or U26880 (N_26880,N_14544,N_16196);
and U26881 (N_26881,N_16461,N_14223);
nor U26882 (N_26882,N_10096,N_16254);
or U26883 (N_26883,N_16444,N_16119);
nand U26884 (N_26884,N_15124,N_18461);
nand U26885 (N_26885,N_13687,N_11544);
and U26886 (N_26886,N_18962,N_17365);
and U26887 (N_26887,N_13970,N_17695);
nor U26888 (N_26888,N_11439,N_13328);
nor U26889 (N_26889,N_19748,N_19681);
and U26890 (N_26890,N_17267,N_10850);
nor U26891 (N_26891,N_15842,N_14300);
nor U26892 (N_26892,N_12105,N_19161);
nor U26893 (N_26893,N_17591,N_10449);
and U26894 (N_26894,N_14971,N_19959);
or U26895 (N_26895,N_10014,N_19402);
and U26896 (N_26896,N_14199,N_15861);
and U26897 (N_26897,N_15436,N_13951);
and U26898 (N_26898,N_11009,N_16551);
or U26899 (N_26899,N_10873,N_10142);
or U26900 (N_26900,N_10075,N_15173);
nand U26901 (N_26901,N_11725,N_14829);
or U26902 (N_26902,N_11881,N_11080);
or U26903 (N_26903,N_18371,N_16194);
nand U26904 (N_26904,N_16546,N_12816);
nor U26905 (N_26905,N_12193,N_12970);
nor U26906 (N_26906,N_14409,N_12976);
nand U26907 (N_26907,N_18492,N_13151);
nand U26908 (N_26908,N_14217,N_14403);
or U26909 (N_26909,N_13166,N_12231);
nand U26910 (N_26910,N_11819,N_11737);
nand U26911 (N_26911,N_18526,N_17258);
nand U26912 (N_26912,N_14624,N_10568);
nor U26913 (N_26913,N_13675,N_10716);
and U26914 (N_26914,N_17318,N_13923);
nor U26915 (N_26915,N_12079,N_16689);
or U26916 (N_26916,N_18758,N_10212);
nand U26917 (N_26917,N_12450,N_12320);
nand U26918 (N_26918,N_11909,N_10500);
nand U26919 (N_26919,N_13126,N_17346);
and U26920 (N_26920,N_16307,N_16261);
or U26921 (N_26921,N_13002,N_18389);
and U26922 (N_26922,N_18602,N_19104);
and U26923 (N_26923,N_13025,N_16948);
nor U26924 (N_26924,N_11810,N_13956);
nor U26925 (N_26925,N_13535,N_19310);
nor U26926 (N_26926,N_15593,N_13531);
and U26927 (N_26927,N_17114,N_10729);
nor U26928 (N_26928,N_17528,N_10845);
or U26929 (N_26929,N_19037,N_15248);
nor U26930 (N_26930,N_10756,N_16469);
and U26931 (N_26931,N_13785,N_12139);
nor U26932 (N_26932,N_17731,N_13667);
nand U26933 (N_26933,N_19017,N_18164);
and U26934 (N_26934,N_13900,N_12640);
and U26935 (N_26935,N_17284,N_12177);
and U26936 (N_26936,N_19571,N_13304);
nor U26937 (N_26937,N_13648,N_11250);
or U26938 (N_26938,N_14417,N_14025);
or U26939 (N_26939,N_19060,N_15464);
and U26940 (N_26940,N_19444,N_16149);
or U26941 (N_26941,N_10108,N_11971);
nor U26942 (N_26942,N_11681,N_18271);
or U26943 (N_26943,N_19758,N_15573);
nand U26944 (N_26944,N_13564,N_11622);
nor U26945 (N_26945,N_19194,N_16980);
or U26946 (N_26946,N_11329,N_12399);
and U26947 (N_26947,N_15756,N_14668);
nand U26948 (N_26948,N_12559,N_19602);
and U26949 (N_26949,N_11588,N_13246);
nor U26950 (N_26950,N_12032,N_19359);
nor U26951 (N_26951,N_12274,N_19908);
or U26952 (N_26952,N_18438,N_10764);
nand U26953 (N_26953,N_18625,N_11618);
nand U26954 (N_26954,N_15765,N_11081);
nor U26955 (N_26955,N_19109,N_16106);
and U26956 (N_26956,N_12109,N_17616);
nand U26957 (N_26957,N_12152,N_19813);
and U26958 (N_26958,N_16787,N_14766);
nor U26959 (N_26959,N_13402,N_17529);
nand U26960 (N_26960,N_11755,N_16763);
or U26961 (N_26961,N_18322,N_18046);
nor U26962 (N_26962,N_10020,N_15188);
or U26963 (N_26963,N_12346,N_14932);
nand U26964 (N_26964,N_17185,N_18716);
nor U26965 (N_26965,N_12083,N_19756);
and U26966 (N_26966,N_12701,N_12611);
nor U26967 (N_26967,N_19245,N_12275);
nand U26968 (N_26968,N_15650,N_11280);
or U26969 (N_26969,N_10464,N_16261);
and U26970 (N_26970,N_14415,N_11641);
or U26971 (N_26971,N_19157,N_18594);
and U26972 (N_26972,N_10589,N_18959);
nand U26973 (N_26973,N_10684,N_13129);
nor U26974 (N_26974,N_19934,N_12515);
or U26975 (N_26975,N_13537,N_14304);
nor U26976 (N_26976,N_18296,N_17558);
or U26977 (N_26977,N_10267,N_10609);
nand U26978 (N_26978,N_15615,N_15419);
nand U26979 (N_26979,N_17826,N_13469);
xor U26980 (N_26980,N_13096,N_17070);
nor U26981 (N_26981,N_15320,N_12241);
nand U26982 (N_26982,N_14706,N_19746);
nor U26983 (N_26983,N_12175,N_16890);
and U26984 (N_26984,N_11431,N_13258);
or U26985 (N_26985,N_17689,N_16089);
nand U26986 (N_26986,N_17136,N_13680);
nand U26987 (N_26987,N_16927,N_12225);
and U26988 (N_26988,N_19697,N_12353);
and U26989 (N_26989,N_12665,N_16932);
nor U26990 (N_26990,N_17450,N_12328);
and U26991 (N_26991,N_14355,N_17506);
and U26992 (N_26992,N_10077,N_14499);
nand U26993 (N_26993,N_16317,N_18680);
nand U26994 (N_26994,N_10102,N_17999);
nand U26995 (N_26995,N_11399,N_17540);
or U26996 (N_26996,N_17649,N_10765);
and U26997 (N_26997,N_15008,N_19344);
and U26998 (N_26998,N_10425,N_11839);
and U26999 (N_26999,N_15965,N_12514);
nor U27000 (N_27000,N_12591,N_16377);
and U27001 (N_27001,N_16665,N_10494);
nand U27002 (N_27002,N_18268,N_11760);
and U27003 (N_27003,N_15244,N_14313);
and U27004 (N_27004,N_15187,N_14625);
nor U27005 (N_27005,N_15934,N_16952);
or U27006 (N_27006,N_13480,N_11617);
nor U27007 (N_27007,N_15499,N_10940);
or U27008 (N_27008,N_18697,N_17179);
and U27009 (N_27009,N_13148,N_10327);
nor U27010 (N_27010,N_17053,N_19070);
or U27011 (N_27011,N_10739,N_16818);
nor U27012 (N_27012,N_14566,N_15520);
and U27013 (N_27013,N_18943,N_18364);
nor U27014 (N_27014,N_19350,N_18986);
or U27015 (N_27015,N_14450,N_18746);
or U27016 (N_27016,N_10102,N_17415);
nor U27017 (N_27017,N_15156,N_16716);
nand U27018 (N_27018,N_12180,N_14980);
and U27019 (N_27019,N_17307,N_11774);
or U27020 (N_27020,N_12014,N_11362);
nand U27021 (N_27021,N_17987,N_14791);
and U27022 (N_27022,N_13396,N_15267);
nor U27023 (N_27023,N_16005,N_16489);
nor U27024 (N_27024,N_10878,N_14396);
and U27025 (N_27025,N_11775,N_13230);
and U27026 (N_27026,N_11610,N_17863);
and U27027 (N_27027,N_14478,N_15657);
or U27028 (N_27028,N_18165,N_13320);
and U27029 (N_27029,N_19882,N_12154);
nor U27030 (N_27030,N_14758,N_19018);
nor U27031 (N_27031,N_17221,N_12224);
nor U27032 (N_27032,N_11774,N_11986);
and U27033 (N_27033,N_12584,N_19328);
nor U27034 (N_27034,N_12491,N_12268);
or U27035 (N_27035,N_10285,N_14762);
and U27036 (N_27036,N_17996,N_13210);
and U27037 (N_27037,N_12152,N_17491);
nand U27038 (N_27038,N_16221,N_11340);
or U27039 (N_27039,N_11432,N_13310);
nor U27040 (N_27040,N_14758,N_18102);
nor U27041 (N_27041,N_19629,N_13767);
and U27042 (N_27042,N_13613,N_15698);
or U27043 (N_27043,N_11453,N_11279);
or U27044 (N_27044,N_12594,N_11739);
nor U27045 (N_27045,N_13901,N_13123);
nor U27046 (N_27046,N_19811,N_11696);
nor U27047 (N_27047,N_12198,N_15249);
nand U27048 (N_27048,N_16577,N_10919);
or U27049 (N_27049,N_15855,N_13072);
or U27050 (N_27050,N_16160,N_19135);
and U27051 (N_27051,N_18178,N_11815);
and U27052 (N_27052,N_14059,N_13789);
nand U27053 (N_27053,N_10172,N_19163);
or U27054 (N_27054,N_15319,N_18557);
nor U27055 (N_27055,N_14394,N_14631);
nor U27056 (N_27056,N_17027,N_15559);
nand U27057 (N_27057,N_19441,N_18156);
or U27058 (N_27058,N_11166,N_18091);
nor U27059 (N_27059,N_11868,N_17459);
or U27060 (N_27060,N_15074,N_11401);
and U27061 (N_27061,N_19213,N_19022);
nand U27062 (N_27062,N_12276,N_13399);
nand U27063 (N_27063,N_19510,N_11220);
nor U27064 (N_27064,N_15576,N_13081);
or U27065 (N_27065,N_11587,N_13369);
nor U27066 (N_27066,N_19062,N_11255);
and U27067 (N_27067,N_10681,N_15075);
nor U27068 (N_27068,N_16314,N_16231);
nor U27069 (N_27069,N_11971,N_13771);
or U27070 (N_27070,N_17101,N_19679);
and U27071 (N_27071,N_13607,N_17220);
nand U27072 (N_27072,N_18928,N_12840);
or U27073 (N_27073,N_13115,N_17284);
and U27074 (N_27074,N_12746,N_17034);
nor U27075 (N_27075,N_19431,N_10160);
or U27076 (N_27076,N_18341,N_16299);
or U27077 (N_27077,N_18170,N_18560);
and U27078 (N_27078,N_19770,N_11365);
nand U27079 (N_27079,N_14015,N_16807);
nor U27080 (N_27080,N_16373,N_12484);
nand U27081 (N_27081,N_12494,N_13745);
nand U27082 (N_27082,N_14658,N_17942);
nand U27083 (N_27083,N_18838,N_17352);
or U27084 (N_27084,N_10256,N_15885);
and U27085 (N_27085,N_14156,N_12234);
nor U27086 (N_27086,N_14851,N_10084);
nor U27087 (N_27087,N_10831,N_18172);
and U27088 (N_27088,N_14593,N_19953);
and U27089 (N_27089,N_17036,N_11161);
nand U27090 (N_27090,N_17525,N_17149);
and U27091 (N_27091,N_13170,N_12350);
and U27092 (N_27092,N_15180,N_11159);
and U27093 (N_27093,N_18809,N_10475);
and U27094 (N_27094,N_11709,N_16004);
and U27095 (N_27095,N_17225,N_12856);
nand U27096 (N_27096,N_10663,N_18876);
or U27097 (N_27097,N_13453,N_10661);
nand U27098 (N_27098,N_10641,N_19766);
or U27099 (N_27099,N_13151,N_13222);
nand U27100 (N_27100,N_16199,N_18248);
nor U27101 (N_27101,N_13669,N_11560);
and U27102 (N_27102,N_17932,N_19508);
nor U27103 (N_27103,N_12086,N_19875);
or U27104 (N_27104,N_18922,N_17172);
nand U27105 (N_27105,N_11970,N_11476);
nand U27106 (N_27106,N_10573,N_15616);
nor U27107 (N_27107,N_17863,N_13292);
and U27108 (N_27108,N_10400,N_13253);
or U27109 (N_27109,N_14187,N_10693);
nor U27110 (N_27110,N_10763,N_13084);
nor U27111 (N_27111,N_11617,N_17672);
and U27112 (N_27112,N_13074,N_18796);
xnor U27113 (N_27113,N_16564,N_10843);
or U27114 (N_27114,N_18684,N_15439);
nand U27115 (N_27115,N_11671,N_19101);
or U27116 (N_27116,N_15530,N_12393);
nor U27117 (N_27117,N_14140,N_17230);
or U27118 (N_27118,N_18338,N_16227);
nor U27119 (N_27119,N_17661,N_14726);
nand U27120 (N_27120,N_14788,N_14400);
or U27121 (N_27121,N_16817,N_14697);
nor U27122 (N_27122,N_19219,N_10628);
or U27123 (N_27123,N_18380,N_16684);
nand U27124 (N_27124,N_16208,N_10690);
and U27125 (N_27125,N_16355,N_12788);
or U27126 (N_27126,N_12749,N_14686);
nor U27127 (N_27127,N_13054,N_19609);
nor U27128 (N_27128,N_19564,N_13400);
nand U27129 (N_27129,N_19050,N_17985);
nand U27130 (N_27130,N_15475,N_18094);
nor U27131 (N_27131,N_18419,N_11060);
nand U27132 (N_27132,N_15220,N_12615);
nor U27133 (N_27133,N_15580,N_12510);
and U27134 (N_27134,N_18994,N_17305);
and U27135 (N_27135,N_10949,N_17761);
nand U27136 (N_27136,N_10401,N_15949);
nor U27137 (N_27137,N_15889,N_18678);
nand U27138 (N_27138,N_11107,N_12921);
nor U27139 (N_27139,N_15498,N_17721);
and U27140 (N_27140,N_17583,N_13243);
and U27141 (N_27141,N_18634,N_18046);
and U27142 (N_27142,N_16836,N_12418);
nor U27143 (N_27143,N_19567,N_17456);
and U27144 (N_27144,N_18586,N_12097);
nand U27145 (N_27145,N_18216,N_14849);
and U27146 (N_27146,N_11823,N_14740);
and U27147 (N_27147,N_18730,N_19600);
or U27148 (N_27148,N_19776,N_16820);
or U27149 (N_27149,N_12772,N_10665);
nand U27150 (N_27150,N_19181,N_10652);
nor U27151 (N_27151,N_12919,N_16834);
nor U27152 (N_27152,N_17823,N_10019);
or U27153 (N_27153,N_14925,N_10010);
nor U27154 (N_27154,N_14980,N_16905);
nor U27155 (N_27155,N_11511,N_13153);
nand U27156 (N_27156,N_18328,N_16409);
and U27157 (N_27157,N_18182,N_19889);
nor U27158 (N_27158,N_11672,N_18005);
or U27159 (N_27159,N_18328,N_17197);
or U27160 (N_27160,N_16379,N_10851);
nand U27161 (N_27161,N_17685,N_13840);
and U27162 (N_27162,N_10526,N_18601);
nand U27163 (N_27163,N_14930,N_19032);
nand U27164 (N_27164,N_18912,N_14822);
nor U27165 (N_27165,N_19535,N_12934);
nand U27166 (N_27166,N_18861,N_14551);
and U27167 (N_27167,N_18565,N_14986);
nand U27168 (N_27168,N_14660,N_10475);
and U27169 (N_27169,N_19838,N_18140);
nor U27170 (N_27170,N_18322,N_12323);
nor U27171 (N_27171,N_19013,N_15939);
nor U27172 (N_27172,N_13684,N_17362);
nand U27173 (N_27173,N_11048,N_19498);
nand U27174 (N_27174,N_17843,N_15568);
nand U27175 (N_27175,N_12205,N_10925);
and U27176 (N_27176,N_10778,N_10211);
nor U27177 (N_27177,N_11173,N_13660);
xor U27178 (N_27178,N_11175,N_15359);
or U27179 (N_27179,N_15610,N_13005);
and U27180 (N_27180,N_14112,N_11792);
nand U27181 (N_27181,N_17465,N_15191);
or U27182 (N_27182,N_18609,N_11422);
and U27183 (N_27183,N_10232,N_11598);
nand U27184 (N_27184,N_16345,N_11934);
and U27185 (N_27185,N_15886,N_18717);
nor U27186 (N_27186,N_12379,N_16281);
nand U27187 (N_27187,N_15853,N_10590);
nor U27188 (N_27188,N_14634,N_11514);
and U27189 (N_27189,N_11237,N_18392);
nor U27190 (N_27190,N_15446,N_19580);
and U27191 (N_27191,N_19643,N_17688);
or U27192 (N_27192,N_12421,N_12850);
nor U27193 (N_27193,N_14936,N_10489);
and U27194 (N_27194,N_10275,N_16963);
or U27195 (N_27195,N_13863,N_11742);
or U27196 (N_27196,N_11699,N_19145);
and U27197 (N_27197,N_13516,N_19344);
nand U27198 (N_27198,N_15903,N_13448);
and U27199 (N_27199,N_11954,N_12955);
or U27200 (N_27200,N_16199,N_17638);
nand U27201 (N_27201,N_18177,N_12855);
nor U27202 (N_27202,N_19121,N_18132);
nor U27203 (N_27203,N_13575,N_19964);
nor U27204 (N_27204,N_11852,N_19088);
and U27205 (N_27205,N_18670,N_11426);
nor U27206 (N_27206,N_11037,N_17206);
and U27207 (N_27207,N_12163,N_17174);
nand U27208 (N_27208,N_19045,N_17670);
nand U27209 (N_27209,N_14755,N_19492);
nand U27210 (N_27210,N_12629,N_15084);
nand U27211 (N_27211,N_14417,N_14765);
and U27212 (N_27212,N_11184,N_15512);
and U27213 (N_27213,N_13729,N_19341);
nand U27214 (N_27214,N_15751,N_18256);
or U27215 (N_27215,N_11868,N_18254);
and U27216 (N_27216,N_18173,N_16130);
and U27217 (N_27217,N_14647,N_11841);
nand U27218 (N_27218,N_18513,N_18089);
xor U27219 (N_27219,N_18858,N_14526);
or U27220 (N_27220,N_17000,N_19705);
nand U27221 (N_27221,N_16632,N_18986);
nor U27222 (N_27222,N_13405,N_17102);
nor U27223 (N_27223,N_17075,N_12026);
or U27224 (N_27224,N_18790,N_17936);
nor U27225 (N_27225,N_14846,N_12589);
or U27226 (N_27226,N_17555,N_11956);
nor U27227 (N_27227,N_14307,N_15385);
nand U27228 (N_27228,N_12685,N_11134);
nand U27229 (N_27229,N_14263,N_19778);
or U27230 (N_27230,N_12925,N_11275);
or U27231 (N_27231,N_18509,N_15233);
or U27232 (N_27232,N_17032,N_11874);
and U27233 (N_27233,N_16065,N_13639);
nand U27234 (N_27234,N_15533,N_13616);
nor U27235 (N_27235,N_14458,N_15979);
nor U27236 (N_27236,N_14908,N_12965);
nor U27237 (N_27237,N_19726,N_19363);
nand U27238 (N_27238,N_19374,N_14178);
nor U27239 (N_27239,N_19079,N_12482);
and U27240 (N_27240,N_19368,N_17123);
or U27241 (N_27241,N_15322,N_13794);
and U27242 (N_27242,N_17008,N_15048);
nand U27243 (N_27243,N_10845,N_11774);
or U27244 (N_27244,N_10935,N_11646);
and U27245 (N_27245,N_12093,N_16917);
nand U27246 (N_27246,N_13107,N_13741);
nor U27247 (N_27247,N_17413,N_12440);
nand U27248 (N_27248,N_17977,N_11083);
nor U27249 (N_27249,N_19410,N_19568);
nor U27250 (N_27250,N_12989,N_13545);
nor U27251 (N_27251,N_19298,N_10449);
nor U27252 (N_27252,N_12989,N_12250);
nand U27253 (N_27253,N_16701,N_11824);
nand U27254 (N_27254,N_19172,N_16792);
nor U27255 (N_27255,N_14585,N_12552);
nor U27256 (N_27256,N_18828,N_14343);
nor U27257 (N_27257,N_17953,N_15903);
or U27258 (N_27258,N_18738,N_18772);
and U27259 (N_27259,N_12341,N_14073);
nand U27260 (N_27260,N_15598,N_10933);
or U27261 (N_27261,N_18503,N_16223);
or U27262 (N_27262,N_10150,N_19742);
or U27263 (N_27263,N_11204,N_10727);
nand U27264 (N_27264,N_19745,N_10330);
and U27265 (N_27265,N_18125,N_10576);
nor U27266 (N_27266,N_12421,N_12217);
nand U27267 (N_27267,N_16260,N_12495);
nor U27268 (N_27268,N_16962,N_18514);
nand U27269 (N_27269,N_11276,N_12659);
nand U27270 (N_27270,N_19981,N_14134);
nor U27271 (N_27271,N_14246,N_16884);
or U27272 (N_27272,N_11550,N_17098);
and U27273 (N_27273,N_14955,N_10503);
nand U27274 (N_27274,N_11991,N_10024);
and U27275 (N_27275,N_17406,N_17223);
nor U27276 (N_27276,N_15494,N_11760);
xnor U27277 (N_27277,N_16842,N_12883);
and U27278 (N_27278,N_13521,N_11027);
or U27279 (N_27279,N_16393,N_16942);
xor U27280 (N_27280,N_14855,N_15825);
xor U27281 (N_27281,N_11229,N_13289);
nor U27282 (N_27282,N_10459,N_11921);
nor U27283 (N_27283,N_10814,N_10690);
or U27284 (N_27284,N_13738,N_10996);
nand U27285 (N_27285,N_12847,N_14910);
and U27286 (N_27286,N_18402,N_18610);
nand U27287 (N_27287,N_18369,N_10627);
or U27288 (N_27288,N_15862,N_11044);
and U27289 (N_27289,N_14732,N_15898);
nand U27290 (N_27290,N_14551,N_14599);
or U27291 (N_27291,N_14351,N_19487);
or U27292 (N_27292,N_18232,N_19627);
nand U27293 (N_27293,N_16263,N_10786);
nor U27294 (N_27294,N_16886,N_10642);
or U27295 (N_27295,N_19561,N_18712);
and U27296 (N_27296,N_13770,N_11939);
and U27297 (N_27297,N_18811,N_17264);
and U27298 (N_27298,N_14844,N_11188);
nor U27299 (N_27299,N_11010,N_15755);
or U27300 (N_27300,N_11388,N_18744);
nor U27301 (N_27301,N_13738,N_17651);
and U27302 (N_27302,N_12574,N_12451);
nand U27303 (N_27303,N_15865,N_12048);
or U27304 (N_27304,N_17181,N_14677);
nand U27305 (N_27305,N_17217,N_18708);
or U27306 (N_27306,N_15625,N_12103);
nor U27307 (N_27307,N_14918,N_13172);
or U27308 (N_27308,N_17462,N_13317);
and U27309 (N_27309,N_12024,N_16143);
or U27310 (N_27310,N_14404,N_14397);
and U27311 (N_27311,N_17394,N_14776);
and U27312 (N_27312,N_10121,N_14109);
and U27313 (N_27313,N_12588,N_13539);
and U27314 (N_27314,N_15434,N_17035);
nor U27315 (N_27315,N_16837,N_14201);
nand U27316 (N_27316,N_12856,N_11516);
nor U27317 (N_27317,N_14972,N_19912);
nand U27318 (N_27318,N_10392,N_14915);
or U27319 (N_27319,N_16173,N_15688);
or U27320 (N_27320,N_13839,N_15905);
nor U27321 (N_27321,N_18473,N_16931);
nor U27322 (N_27322,N_13902,N_14137);
nand U27323 (N_27323,N_10552,N_17537);
nand U27324 (N_27324,N_15727,N_18011);
and U27325 (N_27325,N_17800,N_14280);
or U27326 (N_27326,N_15076,N_19104);
and U27327 (N_27327,N_10309,N_13982);
or U27328 (N_27328,N_11899,N_15643);
nor U27329 (N_27329,N_16701,N_18504);
nand U27330 (N_27330,N_10994,N_11789);
and U27331 (N_27331,N_18573,N_13830);
or U27332 (N_27332,N_16237,N_18621);
nor U27333 (N_27333,N_10582,N_10090);
and U27334 (N_27334,N_13618,N_18264);
or U27335 (N_27335,N_12832,N_19277);
or U27336 (N_27336,N_18929,N_18886);
nor U27337 (N_27337,N_16852,N_10805);
nor U27338 (N_27338,N_11198,N_10255);
nor U27339 (N_27339,N_17464,N_14403);
nor U27340 (N_27340,N_19998,N_17294);
or U27341 (N_27341,N_18783,N_17214);
nor U27342 (N_27342,N_10623,N_18771);
xnor U27343 (N_27343,N_19427,N_14904);
and U27344 (N_27344,N_16094,N_14539);
or U27345 (N_27345,N_17521,N_10471);
and U27346 (N_27346,N_11098,N_15416);
and U27347 (N_27347,N_16429,N_12717);
and U27348 (N_27348,N_11992,N_19110);
nor U27349 (N_27349,N_10557,N_16625);
and U27350 (N_27350,N_13338,N_16061);
nand U27351 (N_27351,N_18281,N_14160);
or U27352 (N_27352,N_15944,N_15246);
or U27353 (N_27353,N_15126,N_17276);
nor U27354 (N_27354,N_15766,N_18781);
and U27355 (N_27355,N_19662,N_15601);
and U27356 (N_27356,N_19742,N_12304);
nand U27357 (N_27357,N_13922,N_19901);
nor U27358 (N_27358,N_16836,N_17531);
nand U27359 (N_27359,N_15101,N_11710);
or U27360 (N_27360,N_18773,N_17833);
or U27361 (N_27361,N_14834,N_13779);
and U27362 (N_27362,N_10415,N_10353);
and U27363 (N_27363,N_10166,N_19117);
nor U27364 (N_27364,N_18666,N_18270);
and U27365 (N_27365,N_16282,N_10709);
or U27366 (N_27366,N_15845,N_11728);
or U27367 (N_27367,N_16610,N_19742);
or U27368 (N_27368,N_19618,N_16265);
and U27369 (N_27369,N_12340,N_14888);
or U27370 (N_27370,N_15527,N_13552);
and U27371 (N_27371,N_10390,N_14093);
or U27372 (N_27372,N_10727,N_18331);
nand U27373 (N_27373,N_16386,N_10606);
or U27374 (N_27374,N_12332,N_18126);
or U27375 (N_27375,N_18267,N_18942);
nand U27376 (N_27376,N_13216,N_17558);
nor U27377 (N_27377,N_14842,N_14250);
nor U27378 (N_27378,N_11741,N_17271);
and U27379 (N_27379,N_10709,N_18574);
nand U27380 (N_27380,N_16251,N_14722);
nand U27381 (N_27381,N_13142,N_13894);
nor U27382 (N_27382,N_17533,N_14332);
nor U27383 (N_27383,N_12001,N_16807);
or U27384 (N_27384,N_18962,N_10680);
nor U27385 (N_27385,N_11248,N_13076);
nand U27386 (N_27386,N_10405,N_18218);
or U27387 (N_27387,N_11711,N_11986);
nand U27388 (N_27388,N_11798,N_14377);
nand U27389 (N_27389,N_15507,N_16049);
or U27390 (N_27390,N_11622,N_16132);
nand U27391 (N_27391,N_10641,N_17947);
or U27392 (N_27392,N_17693,N_10882);
and U27393 (N_27393,N_14938,N_11969);
or U27394 (N_27394,N_16498,N_18307);
or U27395 (N_27395,N_17689,N_11189);
or U27396 (N_27396,N_18933,N_10966);
and U27397 (N_27397,N_14066,N_11992);
and U27398 (N_27398,N_15818,N_19049);
or U27399 (N_27399,N_19248,N_19095);
or U27400 (N_27400,N_19281,N_14629);
and U27401 (N_27401,N_12003,N_17797);
or U27402 (N_27402,N_14579,N_19244);
and U27403 (N_27403,N_13990,N_14017);
nand U27404 (N_27404,N_13018,N_18312);
nand U27405 (N_27405,N_14877,N_13050);
or U27406 (N_27406,N_15459,N_10572);
nand U27407 (N_27407,N_13816,N_19281);
or U27408 (N_27408,N_16439,N_17831);
nand U27409 (N_27409,N_18587,N_15626);
nand U27410 (N_27410,N_14526,N_11118);
or U27411 (N_27411,N_15172,N_18722);
and U27412 (N_27412,N_12491,N_10117);
and U27413 (N_27413,N_16219,N_18333);
nor U27414 (N_27414,N_18220,N_12481);
nor U27415 (N_27415,N_18291,N_12818);
nand U27416 (N_27416,N_17649,N_11539);
nor U27417 (N_27417,N_16067,N_18669);
xor U27418 (N_27418,N_15503,N_12114);
xnor U27419 (N_27419,N_14274,N_15376);
nor U27420 (N_27420,N_19141,N_19097);
nand U27421 (N_27421,N_10621,N_16595);
nand U27422 (N_27422,N_19700,N_11211);
or U27423 (N_27423,N_17588,N_11419);
nand U27424 (N_27424,N_13879,N_13667);
and U27425 (N_27425,N_19255,N_18030);
or U27426 (N_27426,N_15839,N_11644);
or U27427 (N_27427,N_17193,N_14639);
and U27428 (N_27428,N_14625,N_11409);
nand U27429 (N_27429,N_13758,N_12299);
or U27430 (N_27430,N_16804,N_13694);
nand U27431 (N_27431,N_17196,N_10444);
nor U27432 (N_27432,N_18687,N_14634);
nor U27433 (N_27433,N_13336,N_19999);
nand U27434 (N_27434,N_15418,N_12477);
nand U27435 (N_27435,N_16729,N_17054);
nor U27436 (N_27436,N_19047,N_11408);
nand U27437 (N_27437,N_10128,N_13543);
nor U27438 (N_27438,N_14131,N_17890);
nand U27439 (N_27439,N_16465,N_18239);
nor U27440 (N_27440,N_10185,N_18774);
and U27441 (N_27441,N_18003,N_16997);
and U27442 (N_27442,N_10942,N_10046);
or U27443 (N_27443,N_10894,N_17536);
and U27444 (N_27444,N_15791,N_15072);
nand U27445 (N_27445,N_13391,N_14461);
nand U27446 (N_27446,N_15831,N_13241);
nand U27447 (N_27447,N_15912,N_12422);
or U27448 (N_27448,N_14616,N_12393);
nand U27449 (N_27449,N_19825,N_19284);
or U27450 (N_27450,N_14986,N_12383);
nor U27451 (N_27451,N_14179,N_14946);
nor U27452 (N_27452,N_11135,N_10333);
or U27453 (N_27453,N_10083,N_16921);
or U27454 (N_27454,N_15130,N_17103);
or U27455 (N_27455,N_11188,N_19221);
nor U27456 (N_27456,N_11357,N_19679);
nor U27457 (N_27457,N_10635,N_14587);
nor U27458 (N_27458,N_12351,N_10569);
nor U27459 (N_27459,N_12562,N_13587);
and U27460 (N_27460,N_10773,N_19062);
and U27461 (N_27461,N_10437,N_19581);
or U27462 (N_27462,N_12590,N_14126);
nor U27463 (N_27463,N_16197,N_19986);
nand U27464 (N_27464,N_19632,N_11946);
nand U27465 (N_27465,N_12089,N_19245);
or U27466 (N_27466,N_13680,N_12765);
or U27467 (N_27467,N_14628,N_11669);
xor U27468 (N_27468,N_12250,N_18673);
nand U27469 (N_27469,N_15905,N_12725);
and U27470 (N_27470,N_11642,N_13985);
or U27471 (N_27471,N_17508,N_16933);
or U27472 (N_27472,N_10250,N_15528);
nand U27473 (N_27473,N_14624,N_17822);
nand U27474 (N_27474,N_13048,N_18989);
nor U27475 (N_27475,N_18914,N_11388);
or U27476 (N_27476,N_10258,N_14689);
and U27477 (N_27477,N_11837,N_11527);
or U27478 (N_27478,N_15989,N_19307);
nor U27479 (N_27479,N_10964,N_19466);
nand U27480 (N_27480,N_18496,N_13344);
or U27481 (N_27481,N_16530,N_12669);
nand U27482 (N_27482,N_16725,N_10585);
nand U27483 (N_27483,N_19056,N_10308);
and U27484 (N_27484,N_11613,N_18955);
nand U27485 (N_27485,N_12125,N_13185);
or U27486 (N_27486,N_13728,N_15979);
nor U27487 (N_27487,N_19111,N_15683);
and U27488 (N_27488,N_12183,N_10142);
or U27489 (N_27489,N_18882,N_13561);
and U27490 (N_27490,N_11680,N_16820);
and U27491 (N_27491,N_11000,N_15853);
and U27492 (N_27492,N_13883,N_12558);
nor U27493 (N_27493,N_13266,N_15909);
nor U27494 (N_27494,N_16824,N_14105);
or U27495 (N_27495,N_16853,N_17400);
nor U27496 (N_27496,N_19921,N_10277);
nand U27497 (N_27497,N_14839,N_16998);
nand U27498 (N_27498,N_13319,N_14286);
nand U27499 (N_27499,N_12267,N_17627);
or U27500 (N_27500,N_18411,N_16058);
nor U27501 (N_27501,N_14317,N_12329);
nor U27502 (N_27502,N_19251,N_18619);
nor U27503 (N_27503,N_14055,N_18451);
nand U27504 (N_27504,N_10955,N_12762);
or U27505 (N_27505,N_13321,N_16583);
or U27506 (N_27506,N_18994,N_19260);
nand U27507 (N_27507,N_16158,N_19542);
and U27508 (N_27508,N_19961,N_14602);
and U27509 (N_27509,N_12334,N_15257);
or U27510 (N_27510,N_17750,N_14259);
nor U27511 (N_27511,N_13952,N_10682);
and U27512 (N_27512,N_16928,N_13546);
nor U27513 (N_27513,N_17972,N_19308);
nor U27514 (N_27514,N_11044,N_19192);
nor U27515 (N_27515,N_17391,N_10073);
or U27516 (N_27516,N_14748,N_19439);
nor U27517 (N_27517,N_16544,N_11681);
and U27518 (N_27518,N_17597,N_10936);
or U27519 (N_27519,N_13949,N_18375);
and U27520 (N_27520,N_18231,N_13616);
and U27521 (N_27521,N_15686,N_18605);
or U27522 (N_27522,N_15403,N_16467);
nand U27523 (N_27523,N_14181,N_11228);
nor U27524 (N_27524,N_13934,N_19969);
nand U27525 (N_27525,N_14121,N_12218);
or U27526 (N_27526,N_17110,N_16154);
nor U27527 (N_27527,N_17941,N_17113);
nand U27528 (N_27528,N_11361,N_19176);
nor U27529 (N_27529,N_10975,N_13701);
nor U27530 (N_27530,N_10856,N_10459);
nor U27531 (N_27531,N_12216,N_10999);
and U27532 (N_27532,N_10734,N_17205);
nand U27533 (N_27533,N_19585,N_14267);
nand U27534 (N_27534,N_11595,N_18209);
and U27535 (N_27535,N_13822,N_15358);
or U27536 (N_27536,N_10110,N_13664);
nor U27537 (N_27537,N_10470,N_13732);
or U27538 (N_27538,N_14280,N_14867);
and U27539 (N_27539,N_16939,N_14253);
and U27540 (N_27540,N_16019,N_16338);
nor U27541 (N_27541,N_17863,N_15836);
nor U27542 (N_27542,N_13849,N_13012);
nand U27543 (N_27543,N_19305,N_16347);
nor U27544 (N_27544,N_12524,N_11122);
nand U27545 (N_27545,N_10757,N_14697);
xor U27546 (N_27546,N_12909,N_15891);
or U27547 (N_27547,N_14145,N_15168);
or U27548 (N_27548,N_11198,N_18603);
nand U27549 (N_27549,N_14020,N_18676);
or U27550 (N_27550,N_18572,N_12404);
or U27551 (N_27551,N_10464,N_11432);
or U27552 (N_27552,N_14599,N_12460);
and U27553 (N_27553,N_10277,N_14078);
or U27554 (N_27554,N_17730,N_11110);
nor U27555 (N_27555,N_12777,N_13077);
or U27556 (N_27556,N_10721,N_16797);
nor U27557 (N_27557,N_14283,N_10122);
nand U27558 (N_27558,N_16568,N_12215);
nand U27559 (N_27559,N_17775,N_19227);
or U27560 (N_27560,N_11178,N_10510);
and U27561 (N_27561,N_17638,N_15056);
and U27562 (N_27562,N_17728,N_13514);
nand U27563 (N_27563,N_18692,N_19968);
nand U27564 (N_27564,N_12687,N_17292);
nand U27565 (N_27565,N_12268,N_14722);
nor U27566 (N_27566,N_12225,N_13702);
and U27567 (N_27567,N_15581,N_18597);
and U27568 (N_27568,N_18188,N_16192);
or U27569 (N_27569,N_10875,N_13260);
and U27570 (N_27570,N_11287,N_16857);
and U27571 (N_27571,N_18475,N_11575);
nand U27572 (N_27572,N_13169,N_15658);
or U27573 (N_27573,N_13656,N_12303);
or U27574 (N_27574,N_12505,N_17919);
nand U27575 (N_27575,N_16160,N_17552);
or U27576 (N_27576,N_14152,N_16981);
nor U27577 (N_27577,N_14549,N_13384);
nand U27578 (N_27578,N_12845,N_11220);
nor U27579 (N_27579,N_12467,N_13585);
or U27580 (N_27580,N_12904,N_14425);
or U27581 (N_27581,N_19620,N_15454);
nand U27582 (N_27582,N_13242,N_19692);
or U27583 (N_27583,N_19703,N_19415);
or U27584 (N_27584,N_13407,N_15167);
nand U27585 (N_27585,N_13626,N_13386);
or U27586 (N_27586,N_13269,N_12242);
or U27587 (N_27587,N_15614,N_11569);
nor U27588 (N_27588,N_12542,N_15283);
nand U27589 (N_27589,N_17405,N_10083);
nor U27590 (N_27590,N_10813,N_13335);
or U27591 (N_27591,N_10689,N_12995);
and U27592 (N_27592,N_17222,N_19382);
nand U27593 (N_27593,N_12905,N_17728);
and U27594 (N_27594,N_16063,N_15324);
and U27595 (N_27595,N_14199,N_19063);
or U27596 (N_27596,N_10487,N_15493);
nand U27597 (N_27597,N_11806,N_13773);
and U27598 (N_27598,N_18041,N_15413);
nand U27599 (N_27599,N_18325,N_11930);
and U27600 (N_27600,N_13524,N_18964);
nor U27601 (N_27601,N_18922,N_13298);
or U27602 (N_27602,N_18731,N_12896);
nand U27603 (N_27603,N_16181,N_17547);
or U27604 (N_27604,N_17707,N_17428);
nand U27605 (N_27605,N_14550,N_12847);
and U27606 (N_27606,N_11267,N_15796);
nand U27607 (N_27607,N_14474,N_11143);
nand U27608 (N_27608,N_16936,N_18143);
and U27609 (N_27609,N_18220,N_13900);
and U27610 (N_27610,N_10213,N_18762);
or U27611 (N_27611,N_19523,N_15226);
nor U27612 (N_27612,N_10631,N_18421);
nand U27613 (N_27613,N_11372,N_14311);
nor U27614 (N_27614,N_12373,N_17260);
and U27615 (N_27615,N_16155,N_10263);
and U27616 (N_27616,N_11096,N_14306);
and U27617 (N_27617,N_10325,N_10946);
nand U27618 (N_27618,N_10419,N_17985);
or U27619 (N_27619,N_18687,N_11390);
nand U27620 (N_27620,N_18355,N_17003);
and U27621 (N_27621,N_11702,N_17021);
nor U27622 (N_27622,N_15289,N_15326);
nor U27623 (N_27623,N_17298,N_12663);
or U27624 (N_27624,N_17825,N_11389);
nor U27625 (N_27625,N_18918,N_14848);
nand U27626 (N_27626,N_14380,N_16611);
and U27627 (N_27627,N_11875,N_19222);
and U27628 (N_27628,N_11346,N_15819);
and U27629 (N_27629,N_13251,N_14763);
nand U27630 (N_27630,N_19146,N_10451);
nor U27631 (N_27631,N_17306,N_12724);
and U27632 (N_27632,N_14064,N_11178);
nand U27633 (N_27633,N_13092,N_11682);
or U27634 (N_27634,N_19135,N_13236);
or U27635 (N_27635,N_15180,N_16713);
nor U27636 (N_27636,N_17679,N_17307);
or U27637 (N_27637,N_19156,N_17098);
and U27638 (N_27638,N_11085,N_18714);
and U27639 (N_27639,N_11824,N_19072);
nand U27640 (N_27640,N_11457,N_11712);
nor U27641 (N_27641,N_16061,N_11095);
xor U27642 (N_27642,N_14513,N_19516);
and U27643 (N_27643,N_18586,N_19329);
and U27644 (N_27644,N_15571,N_11367);
nand U27645 (N_27645,N_14157,N_11276);
and U27646 (N_27646,N_15456,N_18739);
and U27647 (N_27647,N_13461,N_18550);
nand U27648 (N_27648,N_18599,N_13513);
or U27649 (N_27649,N_10746,N_13181);
and U27650 (N_27650,N_10004,N_15960);
or U27651 (N_27651,N_15049,N_13541);
nand U27652 (N_27652,N_19801,N_12626);
or U27653 (N_27653,N_11455,N_14000);
nand U27654 (N_27654,N_19981,N_12873);
nor U27655 (N_27655,N_17379,N_10507);
nand U27656 (N_27656,N_16284,N_14251);
and U27657 (N_27657,N_12936,N_13058);
nor U27658 (N_27658,N_19871,N_12955);
or U27659 (N_27659,N_15086,N_17600);
and U27660 (N_27660,N_18104,N_17163);
nand U27661 (N_27661,N_16553,N_16086);
and U27662 (N_27662,N_13006,N_15530);
nand U27663 (N_27663,N_12407,N_13680);
nor U27664 (N_27664,N_13502,N_18776);
nor U27665 (N_27665,N_16138,N_17787);
and U27666 (N_27666,N_16965,N_11805);
or U27667 (N_27667,N_12605,N_15300);
or U27668 (N_27668,N_11274,N_19969);
nor U27669 (N_27669,N_18180,N_19639);
or U27670 (N_27670,N_14277,N_12394);
or U27671 (N_27671,N_13120,N_13820);
and U27672 (N_27672,N_15855,N_12237);
or U27673 (N_27673,N_15115,N_18352);
or U27674 (N_27674,N_10147,N_12544);
nor U27675 (N_27675,N_14489,N_11361);
xor U27676 (N_27676,N_10956,N_10148);
and U27677 (N_27677,N_17556,N_14882);
nor U27678 (N_27678,N_19790,N_15736);
or U27679 (N_27679,N_18729,N_18886);
nand U27680 (N_27680,N_17932,N_19740);
or U27681 (N_27681,N_11108,N_10153);
and U27682 (N_27682,N_11832,N_12807);
and U27683 (N_27683,N_17878,N_19204);
or U27684 (N_27684,N_16326,N_18290);
and U27685 (N_27685,N_12134,N_10799);
nor U27686 (N_27686,N_16686,N_11518);
or U27687 (N_27687,N_14748,N_19009);
nor U27688 (N_27688,N_11417,N_17238);
and U27689 (N_27689,N_15718,N_13112);
nand U27690 (N_27690,N_17234,N_19282);
or U27691 (N_27691,N_19532,N_16521);
nand U27692 (N_27692,N_17921,N_14569);
and U27693 (N_27693,N_13237,N_12531);
nand U27694 (N_27694,N_12752,N_17443);
or U27695 (N_27695,N_15471,N_18860);
and U27696 (N_27696,N_18053,N_17827);
and U27697 (N_27697,N_19411,N_12233);
nand U27698 (N_27698,N_14502,N_14106);
nand U27699 (N_27699,N_11735,N_15777);
nand U27700 (N_27700,N_17464,N_15517);
and U27701 (N_27701,N_12675,N_14314);
or U27702 (N_27702,N_15517,N_12065);
or U27703 (N_27703,N_18015,N_11095);
and U27704 (N_27704,N_15841,N_12198);
or U27705 (N_27705,N_12624,N_10800);
nand U27706 (N_27706,N_15803,N_12990);
nand U27707 (N_27707,N_14165,N_15480);
and U27708 (N_27708,N_10785,N_17798);
xor U27709 (N_27709,N_17825,N_19415);
or U27710 (N_27710,N_13698,N_12889);
or U27711 (N_27711,N_15831,N_19388);
nand U27712 (N_27712,N_13745,N_18527);
nand U27713 (N_27713,N_17725,N_15592);
nor U27714 (N_27714,N_18437,N_15082);
nand U27715 (N_27715,N_19992,N_18668);
nor U27716 (N_27716,N_11574,N_14756);
and U27717 (N_27717,N_14156,N_10620);
nor U27718 (N_27718,N_16851,N_13765);
or U27719 (N_27719,N_18006,N_17178);
and U27720 (N_27720,N_10792,N_19281);
or U27721 (N_27721,N_18388,N_16470);
nor U27722 (N_27722,N_14510,N_10376);
nor U27723 (N_27723,N_12089,N_18184);
nand U27724 (N_27724,N_16809,N_11190);
or U27725 (N_27725,N_19105,N_17168);
nand U27726 (N_27726,N_19020,N_10646);
and U27727 (N_27727,N_16980,N_10373);
nor U27728 (N_27728,N_18083,N_19624);
nand U27729 (N_27729,N_18934,N_19040);
or U27730 (N_27730,N_15419,N_17058);
or U27731 (N_27731,N_17498,N_11282);
and U27732 (N_27732,N_11387,N_13905);
xor U27733 (N_27733,N_17715,N_15789);
nor U27734 (N_27734,N_19828,N_18098);
and U27735 (N_27735,N_15881,N_14002);
nand U27736 (N_27736,N_10830,N_14933);
nor U27737 (N_27737,N_11224,N_16174);
or U27738 (N_27738,N_10310,N_14691);
or U27739 (N_27739,N_14582,N_13667);
or U27740 (N_27740,N_13582,N_12818);
nor U27741 (N_27741,N_10421,N_19930);
and U27742 (N_27742,N_12807,N_11342);
xor U27743 (N_27743,N_10624,N_17892);
nand U27744 (N_27744,N_18590,N_17227);
nor U27745 (N_27745,N_15587,N_19815);
nand U27746 (N_27746,N_18621,N_17629);
nand U27747 (N_27747,N_11493,N_10870);
and U27748 (N_27748,N_18785,N_12660);
nor U27749 (N_27749,N_19968,N_10309);
or U27750 (N_27750,N_11263,N_17774);
nand U27751 (N_27751,N_19501,N_10322);
nand U27752 (N_27752,N_15344,N_11082);
or U27753 (N_27753,N_13523,N_16268);
and U27754 (N_27754,N_13631,N_19428);
xnor U27755 (N_27755,N_19378,N_13612);
nand U27756 (N_27756,N_12869,N_19808);
nand U27757 (N_27757,N_15537,N_11030);
or U27758 (N_27758,N_11214,N_16548);
nor U27759 (N_27759,N_15593,N_15421);
or U27760 (N_27760,N_19338,N_13527);
or U27761 (N_27761,N_14659,N_14664);
nor U27762 (N_27762,N_16497,N_16644);
and U27763 (N_27763,N_16047,N_14006);
or U27764 (N_27764,N_15001,N_11757);
or U27765 (N_27765,N_13815,N_17602);
or U27766 (N_27766,N_11102,N_12755);
nor U27767 (N_27767,N_16022,N_12951);
nor U27768 (N_27768,N_16842,N_17122);
and U27769 (N_27769,N_12567,N_19536);
or U27770 (N_27770,N_14730,N_16557);
nor U27771 (N_27771,N_15978,N_16982);
nand U27772 (N_27772,N_10850,N_13772);
nor U27773 (N_27773,N_17499,N_10187);
nand U27774 (N_27774,N_15804,N_13537);
and U27775 (N_27775,N_11115,N_18934);
or U27776 (N_27776,N_11856,N_19507);
or U27777 (N_27777,N_10652,N_13427);
nor U27778 (N_27778,N_12538,N_10215);
or U27779 (N_27779,N_11614,N_15531);
nand U27780 (N_27780,N_15290,N_10686);
nor U27781 (N_27781,N_12674,N_19323);
xnor U27782 (N_27782,N_17931,N_13144);
and U27783 (N_27783,N_12219,N_10371);
or U27784 (N_27784,N_17311,N_12048);
or U27785 (N_27785,N_10689,N_19690);
nor U27786 (N_27786,N_14604,N_12264);
and U27787 (N_27787,N_11500,N_16805);
nor U27788 (N_27788,N_14384,N_11236);
nand U27789 (N_27789,N_10432,N_13051);
or U27790 (N_27790,N_14244,N_12114);
and U27791 (N_27791,N_17563,N_16448);
nor U27792 (N_27792,N_10125,N_13847);
nor U27793 (N_27793,N_10347,N_19873);
nand U27794 (N_27794,N_15339,N_17599);
or U27795 (N_27795,N_16029,N_12846);
nor U27796 (N_27796,N_11763,N_10500);
or U27797 (N_27797,N_14377,N_13589);
or U27798 (N_27798,N_16778,N_15390);
and U27799 (N_27799,N_17204,N_16693);
and U27800 (N_27800,N_16854,N_19266);
and U27801 (N_27801,N_17327,N_19216);
nand U27802 (N_27802,N_12549,N_10608);
and U27803 (N_27803,N_11368,N_15317);
nand U27804 (N_27804,N_11685,N_10016);
or U27805 (N_27805,N_13732,N_19808);
nor U27806 (N_27806,N_11859,N_18255);
nor U27807 (N_27807,N_11292,N_19340);
and U27808 (N_27808,N_16902,N_18740);
nor U27809 (N_27809,N_11345,N_16176);
nor U27810 (N_27810,N_13050,N_11105);
nor U27811 (N_27811,N_11308,N_19305);
nand U27812 (N_27812,N_10759,N_19341);
xor U27813 (N_27813,N_15459,N_12466);
or U27814 (N_27814,N_12425,N_16853);
nand U27815 (N_27815,N_19836,N_18913);
or U27816 (N_27816,N_14778,N_11214);
nor U27817 (N_27817,N_17007,N_12213);
and U27818 (N_27818,N_14542,N_14266);
nor U27819 (N_27819,N_12762,N_19880);
and U27820 (N_27820,N_17150,N_10502);
nand U27821 (N_27821,N_17247,N_10375);
nor U27822 (N_27822,N_17388,N_12482);
nand U27823 (N_27823,N_15669,N_19840);
nand U27824 (N_27824,N_15031,N_13714);
and U27825 (N_27825,N_16260,N_12208);
or U27826 (N_27826,N_16534,N_15291);
or U27827 (N_27827,N_10871,N_14350);
nand U27828 (N_27828,N_16204,N_10922);
or U27829 (N_27829,N_18656,N_17267);
or U27830 (N_27830,N_16267,N_13835);
or U27831 (N_27831,N_12378,N_12462);
or U27832 (N_27832,N_13199,N_19926);
nand U27833 (N_27833,N_16092,N_10556);
nor U27834 (N_27834,N_14176,N_16276);
nor U27835 (N_27835,N_12603,N_12377);
nand U27836 (N_27836,N_10088,N_14154);
and U27837 (N_27837,N_12078,N_19076);
nand U27838 (N_27838,N_19508,N_14043);
xor U27839 (N_27839,N_19260,N_13081);
and U27840 (N_27840,N_11035,N_10883);
nand U27841 (N_27841,N_14367,N_15171);
nor U27842 (N_27842,N_19901,N_18124);
and U27843 (N_27843,N_19158,N_18646);
nor U27844 (N_27844,N_16694,N_12487);
nand U27845 (N_27845,N_17258,N_13166);
or U27846 (N_27846,N_10116,N_14545);
and U27847 (N_27847,N_13284,N_14174);
nor U27848 (N_27848,N_16432,N_17388);
or U27849 (N_27849,N_18033,N_16893);
nand U27850 (N_27850,N_13651,N_18207);
or U27851 (N_27851,N_17485,N_13722);
or U27852 (N_27852,N_18373,N_13851);
nor U27853 (N_27853,N_16094,N_15412);
or U27854 (N_27854,N_18166,N_16266);
or U27855 (N_27855,N_15028,N_14771);
and U27856 (N_27856,N_10109,N_14334);
or U27857 (N_27857,N_18960,N_14278);
nand U27858 (N_27858,N_18396,N_12282);
xor U27859 (N_27859,N_11555,N_16843);
nor U27860 (N_27860,N_13136,N_17205);
or U27861 (N_27861,N_13282,N_10753);
and U27862 (N_27862,N_13036,N_11256);
nor U27863 (N_27863,N_16568,N_19425);
and U27864 (N_27864,N_10591,N_19481);
nor U27865 (N_27865,N_10854,N_12354);
nor U27866 (N_27866,N_16097,N_15477);
and U27867 (N_27867,N_19422,N_18770);
and U27868 (N_27868,N_11135,N_16707);
and U27869 (N_27869,N_17667,N_18077);
nor U27870 (N_27870,N_18048,N_17625);
nand U27871 (N_27871,N_12878,N_18465);
or U27872 (N_27872,N_18815,N_12640);
nand U27873 (N_27873,N_17926,N_13473);
and U27874 (N_27874,N_16587,N_11742);
nor U27875 (N_27875,N_18712,N_14946);
nand U27876 (N_27876,N_16867,N_13304);
or U27877 (N_27877,N_13765,N_16527);
or U27878 (N_27878,N_19439,N_18529);
nor U27879 (N_27879,N_17006,N_16504);
or U27880 (N_27880,N_10768,N_14137);
or U27881 (N_27881,N_16421,N_11683);
or U27882 (N_27882,N_19724,N_16749);
or U27883 (N_27883,N_12724,N_19377);
nor U27884 (N_27884,N_12053,N_12098);
nor U27885 (N_27885,N_11298,N_19905);
nand U27886 (N_27886,N_16316,N_13041);
or U27887 (N_27887,N_13360,N_19508);
and U27888 (N_27888,N_10716,N_19292);
nor U27889 (N_27889,N_14995,N_18401);
nand U27890 (N_27890,N_15849,N_17558);
and U27891 (N_27891,N_14200,N_12527);
nor U27892 (N_27892,N_10514,N_12175);
and U27893 (N_27893,N_16229,N_11475);
and U27894 (N_27894,N_19015,N_19523);
or U27895 (N_27895,N_15776,N_13043);
nand U27896 (N_27896,N_17745,N_17761);
or U27897 (N_27897,N_15896,N_17607);
and U27898 (N_27898,N_16074,N_15899);
and U27899 (N_27899,N_14288,N_12836);
or U27900 (N_27900,N_16496,N_18458);
or U27901 (N_27901,N_10399,N_10873);
nor U27902 (N_27902,N_10387,N_14760);
nor U27903 (N_27903,N_13654,N_12880);
nand U27904 (N_27904,N_17617,N_16941);
nand U27905 (N_27905,N_18591,N_11177);
nor U27906 (N_27906,N_15071,N_13389);
or U27907 (N_27907,N_15429,N_10720);
nand U27908 (N_27908,N_17991,N_14821);
xor U27909 (N_27909,N_12355,N_10775);
nand U27910 (N_27910,N_19981,N_11827);
and U27911 (N_27911,N_11199,N_11734);
nor U27912 (N_27912,N_13119,N_17077);
nor U27913 (N_27913,N_11392,N_11135);
or U27914 (N_27914,N_17986,N_14509);
nor U27915 (N_27915,N_19408,N_14304);
xnor U27916 (N_27916,N_13536,N_19475);
nor U27917 (N_27917,N_12834,N_19969);
or U27918 (N_27918,N_10462,N_15500);
nand U27919 (N_27919,N_15544,N_14297);
and U27920 (N_27920,N_12093,N_17763);
nor U27921 (N_27921,N_18657,N_14462);
or U27922 (N_27922,N_18446,N_19205);
nand U27923 (N_27923,N_18042,N_14870);
and U27924 (N_27924,N_15726,N_15576);
or U27925 (N_27925,N_19505,N_18150);
nor U27926 (N_27926,N_17803,N_17867);
nor U27927 (N_27927,N_19337,N_11977);
and U27928 (N_27928,N_19956,N_14483);
or U27929 (N_27929,N_19257,N_18537);
and U27930 (N_27930,N_11377,N_18581);
nor U27931 (N_27931,N_19049,N_12880);
or U27932 (N_27932,N_19584,N_13098);
nor U27933 (N_27933,N_17931,N_13094);
and U27934 (N_27934,N_13694,N_19034);
nor U27935 (N_27935,N_10023,N_10047);
or U27936 (N_27936,N_15904,N_16103);
and U27937 (N_27937,N_10438,N_10092);
nand U27938 (N_27938,N_17428,N_10794);
and U27939 (N_27939,N_14409,N_10706);
or U27940 (N_27940,N_16173,N_15395);
and U27941 (N_27941,N_15643,N_11626);
nor U27942 (N_27942,N_11852,N_17456);
nand U27943 (N_27943,N_18271,N_11406);
or U27944 (N_27944,N_17219,N_17753);
and U27945 (N_27945,N_16983,N_11167);
nand U27946 (N_27946,N_18085,N_14838);
nand U27947 (N_27947,N_11104,N_12187);
nand U27948 (N_27948,N_11143,N_19520);
or U27949 (N_27949,N_13033,N_16845);
nand U27950 (N_27950,N_15850,N_18515);
or U27951 (N_27951,N_19530,N_13352);
and U27952 (N_27952,N_14452,N_16154);
nor U27953 (N_27953,N_19938,N_14532);
nor U27954 (N_27954,N_19349,N_17148);
and U27955 (N_27955,N_17906,N_15619);
nor U27956 (N_27956,N_12514,N_18181);
nand U27957 (N_27957,N_15799,N_12550);
nor U27958 (N_27958,N_12819,N_13078);
nor U27959 (N_27959,N_19772,N_17771);
nand U27960 (N_27960,N_14331,N_10257);
or U27961 (N_27961,N_16528,N_12048);
and U27962 (N_27962,N_11922,N_17437);
nor U27963 (N_27963,N_13062,N_18196);
nand U27964 (N_27964,N_17586,N_19983);
nand U27965 (N_27965,N_15496,N_16349);
and U27966 (N_27966,N_17496,N_16357);
or U27967 (N_27967,N_10529,N_17130);
or U27968 (N_27968,N_17796,N_11618);
or U27969 (N_27969,N_14268,N_17699);
nor U27970 (N_27970,N_17253,N_19983);
and U27971 (N_27971,N_10153,N_17117);
nor U27972 (N_27972,N_13779,N_17942);
and U27973 (N_27973,N_15855,N_14275);
nor U27974 (N_27974,N_18228,N_11168);
and U27975 (N_27975,N_18105,N_18160);
and U27976 (N_27976,N_18522,N_12625);
nor U27977 (N_27977,N_11392,N_18355);
nor U27978 (N_27978,N_10092,N_15593);
xor U27979 (N_27979,N_14214,N_19917);
nor U27980 (N_27980,N_12597,N_10242);
nand U27981 (N_27981,N_12364,N_14461);
nor U27982 (N_27982,N_18993,N_17918);
nor U27983 (N_27983,N_17506,N_19155);
nor U27984 (N_27984,N_14231,N_13180);
or U27985 (N_27985,N_19896,N_18189);
or U27986 (N_27986,N_16487,N_14425);
and U27987 (N_27987,N_10389,N_12350);
nor U27988 (N_27988,N_16275,N_12315);
nor U27989 (N_27989,N_18484,N_10473);
and U27990 (N_27990,N_17102,N_10370);
and U27991 (N_27991,N_15336,N_12759);
and U27992 (N_27992,N_10184,N_16079);
or U27993 (N_27993,N_12846,N_17054);
nor U27994 (N_27994,N_11267,N_16049);
or U27995 (N_27995,N_11473,N_17472);
and U27996 (N_27996,N_19802,N_10776);
nand U27997 (N_27997,N_10636,N_19729);
nor U27998 (N_27998,N_10646,N_16654);
xnor U27999 (N_27999,N_19913,N_14896);
nand U28000 (N_28000,N_14622,N_13820);
or U28001 (N_28001,N_10118,N_18429);
nand U28002 (N_28002,N_19391,N_10550);
or U28003 (N_28003,N_11343,N_12087);
and U28004 (N_28004,N_13107,N_18992);
and U28005 (N_28005,N_15932,N_19971);
and U28006 (N_28006,N_12150,N_15865);
or U28007 (N_28007,N_12068,N_14047);
and U28008 (N_28008,N_13529,N_19990);
or U28009 (N_28009,N_18312,N_10109);
or U28010 (N_28010,N_14940,N_14606);
nand U28011 (N_28011,N_10606,N_16040);
and U28012 (N_28012,N_18480,N_13988);
or U28013 (N_28013,N_18841,N_14891);
nand U28014 (N_28014,N_17407,N_16485);
or U28015 (N_28015,N_13063,N_14223);
or U28016 (N_28016,N_17757,N_16122);
nand U28017 (N_28017,N_12426,N_15369);
or U28018 (N_28018,N_15267,N_18748);
and U28019 (N_28019,N_17563,N_12509);
nor U28020 (N_28020,N_15512,N_15981);
nor U28021 (N_28021,N_12226,N_15757);
nand U28022 (N_28022,N_14264,N_17871);
or U28023 (N_28023,N_13606,N_19476);
xnor U28024 (N_28024,N_17267,N_16570);
nor U28025 (N_28025,N_15597,N_11169);
nor U28026 (N_28026,N_18947,N_13453);
and U28027 (N_28027,N_12184,N_11498);
and U28028 (N_28028,N_13486,N_15113);
nand U28029 (N_28029,N_13923,N_16180);
nand U28030 (N_28030,N_10993,N_14573);
or U28031 (N_28031,N_12733,N_18703);
nand U28032 (N_28032,N_13835,N_14921);
nand U28033 (N_28033,N_14484,N_15749);
nor U28034 (N_28034,N_16755,N_13355);
nor U28035 (N_28035,N_14372,N_13512);
nand U28036 (N_28036,N_18945,N_12687);
and U28037 (N_28037,N_13236,N_14659);
nand U28038 (N_28038,N_18756,N_19038);
nor U28039 (N_28039,N_14817,N_17546);
nand U28040 (N_28040,N_13970,N_12096);
nand U28041 (N_28041,N_16767,N_12326);
or U28042 (N_28042,N_19666,N_17848);
nand U28043 (N_28043,N_12728,N_17887);
nand U28044 (N_28044,N_16813,N_11737);
nor U28045 (N_28045,N_16300,N_13242);
and U28046 (N_28046,N_11426,N_15760);
and U28047 (N_28047,N_12482,N_19663);
and U28048 (N_28048,N_14127,N_13270);
nand U28049 (N_28049,N_13091,N_12183);
or U28050 (N_28050,N_11594,N_15332);
nand U28051 (N_28051,N_14777,N_10357);
nand U28052 (N_28052,N_14393,N_17406);
or U28053 (N_28053,N_19125,N_15233);
nor U28054 (N_28054,N_13247,N_11807);
nand U28055 (N_28055,N_13983,N_12491);
nand U28056 (N_28056,N_15560,N_10180);
nand U28057 (N_28057,N_13412,N_12701);
and U28058 (N_28058,N_18028,N_16246);
nor U28059 (N_28059,N_16027,N_12099);
nor U28060 (N_28060,N_14052,N_11466);
nand U28061 (N_28061,N_14312,N_12493);
and U28062 (N_28062,N_13895,N_16115);
and U28063 (N_28063,N_12740,N_10434);
or U28064 (N_28064,N_13676,N_16074);
nand U28065 (N_28065,N_18454,N_15639);
nand U28066 (N_28066,N_12870,N_11038);
or U28067 (N_28067,N_14494,N_10423);
nand U28068 (N_28068,N_18025,N_14800);
or U28069 (N_28069,N_11391,N_18412);
or U28070 (N_28070,N_13311,N_15066);
and U28071 (N_28071,N_17376,N_10546);
nor U28072 (N_28072,N_14645,N_13756);
nor U28073 (N_28073,N_19682,N_13461);
nor U28074 (N_28074,N_18743,N_19694);
or U28075 (N_28075,N_18953,N_18133);
or U28076 (N_28076,N_18456,N_13215);
nand U28077 (N_28077,N_19200,N_13216);
or U28078 (N_28078,N_11649,N_16383);
nor U28079 (N_28079,N_11761,N_14614);
nand U28080 (N_28080,N_13652,N_14932);
and U28081 (N_28081,N_11898,N_12129);
nor U28082 (N_28082,N_19773,N_17965);
nor U28083 (N_28083,N_11740,N_16328);
nand U28084 (N_28084,N_18625,N_11553);
and U28085 (N_28085,N_12758,N_17797);
or U28086 (N_28086,N_10340,N_19707);
or U28087 (N_28087,N_12432,N_11818);
or U28088 (N_28088,N_16761,N_15355);
nor U28089 (N_28089,N_17170,N_18403);
nor U28090 (N_28090,N_19287,N_12724);
nor U28091 (N_28091,N_13282,N_10244);
nand U28092 (N_28092,N_19333,N_16677);
or U28093 (N_28093,N_12913,N_15332);
nand U28094 (N_28094,N_19022,N_10151);
and U28095 (N_28095,N_16232,N_10614);
nor U28096 (N_28096,N_18038,N_12455);
nor U28097 (N_28097,N_15792,N_14755);
nor U28098 (N_28098,N_14365,N_18901);
nand U28099 (N_28099,N_10371,N_12874);
and U28100 (N_28100,N_12358,N_12255);
nand U28101 (N_28101,N_17035,N_17418);
and U28102 (N_28102,N_18109,N_17468);
and U28103 (N_28103,N_12350,N_13653);
nor U28104 (N_28104,N_16754,N_18755);
nor U28105 (N_28105,N_10012,N_14722);
nand U28106 (N_28106,N_13427,N_14570);
nor U28107 (N_28107,N_13230,N_12007);
nand U28108 (N_28108,N_13760,N_17506);
nor U28109 (N_28109,N_17838,N_10752);
nand U28110 (N_28110,N_12374,N_16022);
or U28111 (N_28111,N_19398,N_18832);
and U28112 (N_28112,N_13845,N_11869);
nor U28113 (N_28113,N_10028,N_12950);
nand U28114 (N_28114,N_16052,N_13920);
or U28115 (N_28115,N_13975,N_19495);
nand U28116 (N_28116,N_10637,N_12031);
or U28117 (N_28117,N_15169,N_16200);
or U28118 (N_28118,N_15474,N_10364);
nand U28119 (N_28119,N_17182,N_11206);
and U28120 (N_28120,N_12278,N_18429);
nor U28121 (N_28121,N_18238,N_13548);
or U28122 (N_28122,N_14736,N_14761);
nand U28123 (N_28123,N_14695,N_11905);
nor U28124 (N_28124,N_11818,N_12060);
nor U28125 (N_28125,N_18501,N_11878);
nor U28126 (N_28126,N_17967,N_14792);
nand U28127 (N_28127,N_18716,N_14888);
nand U28128 (N_28128,N_18002,N_10379);
nor U28129 (N_28129,N_19115,N_14621);
and U28130 (N_28130,N_10023,N_12948);
nor U28131 (N_28131,N_12630,N_18154);
nor U28132 (N_28132,N_16373,N_18346);
nand U28133 (N_28133,N_17020,N_16647);
nand U28134 (N_28134,N_11840,N_17605);
or U28135 (N_28135,N_14062,N_15371);
or U28136 (N_28136,N_17118,N_19722);
nor U28137 (N_28137,N_12875,N_18636);
or U28138 (N_28138,N_13325,N_12165);
nand U28139 (N_28139,N_11125,N_19040);
xnor U28140 (N_28140,N_10638,N_17470);
nor U28141 (N_28141,N_16580,N_18960);
nand U28142 (N_28142,N_17801,N_11095);
and U28143 (N_28143,N_18464,N_15122);
or U28144 (N_28144,N_17348,N_11123);
nor U28145 (N_28145,N_11215,N_19528);
or U28146 (N_28146,N_17146,N_10650);
or U28147 (N_28147,N_15973,N_11917);
or U28148 (N_28148,N_11158,N_14153);
or U28149 (N_28149,N_16186,N_13632);
and U28150 (N_28150,N_11846,N_15442);
nor U28151 (N_28151,N_19514,N_18459);
or U28152 (N_28152,N_11120,N_11725);
or U28153 (N_28153,N_18735,N_19952);
and U28154 (N_28154,N_17474,N_19678);
nor U28155 (N_28155,N_14981,N_18508);
or U28156 (N_28156,N_18119,N_14202);
and U28157 (N_28157,N_16330,N_16051);
nand U28158 (N_28158,N_13387,N_18233);
and U28159 (N_28159,N_11193,N_11458);
or U28160 (N_28160,N_16850,N_19923);
and U28161 (N_28161,N_19008,N_19853);
or U28162 (N_28162,N_17256,N_19285);
nand U28163 (N_28163,N_18828,N_18927);
nor U28164 (N_28164,N_18490,N_14573);
or U28165 (N_28165,N_16468,N_16449);
or U28166 (N_28166,N_19239,N_15945);
or U28167 (N_28167,N_10200,N_18892);
or U28168 (N_28168,N_12715,N_16529);
nand U28169 (N_28169,N_12648,N_14133);
nor U28170 (N_28170,N_13784,N_13738);
nor U28171 (N_28171,N_12747,N_13732);
and U28172 (N_28172,N_17578,N_16389);
or U28173 (N_28173,N_11690,N_14635);
nor U28174 (N_28174,N_18987,N_15864);
nor U28175 (N_28175,N_13177,N_15553);
nand U28176 (N_28176,N_12452,N_15594);
nor U28177 (N_28177,N_18822,N_16819);
and U28178 (N_28178,N_12940,N_11556);
or U28179 (N_28179,N_14124,N_11184);
and U28180 (N_28180,N_16841,N_17220);
or U28181 (N_28181,N_16328,N_16495);
nor U28182 (N_28182,N_13478,N_19833);
nand U28183 (N_28183,N_16059,N_11001);
or U28184 (N_28184,N_19500,N_16358);
nand U28185 (N_28185,N_12515,N_19977);
nand U28186 (N_28186,N_18352,N_13525);
or U28187 (N_28187,N_19205,N_16483);
nor U28188 (N_28188,N_19105,N_15856);
nor U28189 (N_28189,N_16486,N_19708);
or U28190 (N_28190,N_11604,N_13293);
and U28191 (N_28191,N_13591,N_17473);
and U28192 (N_28192,N_16187,N_12330);
and U28193 (N_28193,N_17587,N_16334);
nand U28194 (N_28194,N_18204,N_14042);
or U28195 (N_28195,N_15017,N_15339);
and U28196 (N_28196,N_10788,N_13182);
xnor U28197 (N_28197,N_13571,N_13227);
or U28198 (N_28198,N_19984,N_12989);
nor U28199 (N_28199,N_10456,N_19673);
or U28200 (N_28200,N_19316,N_17827);
nand U28201 (N_28201,N_11724,N_14289);
nor U28202 (N_28202,N_10660,N_19579);
or U28203 (N_28203,N_14820,N_10231);
nor U28204 (N_28204,N_12580,N_13567);
nor U28205 (N_28205,N_12743,N_16321);
nor U28206 (N_28206,N_15241,N_11451);
or U28207 (N_28207,N_15267,N_10174);
nor U28208 (N_28208,N_19338,N_14495);
nor U28209 (N_28209,N_11839,N_14699);
or U28210 (N_28210,N_10079,N_18300);
nor U28211 (N_28211,N_19560,N_18276);
nand U28212 (N_28212,N_18328,N_13215);
or U28213 (N_28213,N_18311,N_13957);
or U28214 (N_28214,N_13222,N_11670);
and U28215 (N_28215,N_15568,N_17888);
nor U28216 (N_28216,N_19864,N_16395);
or U28217 (N_28217,N_18861,N_13245);
and U28218 (N_28218,N_10694,N_18954);
or U28219 (N_28219,N_10440,N_13978);
nor U28220 (N_28220,N_14689,N_17274);
nand U28221 (N_28221,N_10471,N_11488);
nor U28222 (N_28222,N_11833,N_13167);
or U28223 (N_28223,N_14372,N_10280);
and U28224 (N_28224,N_19827,N_11422);
nor U28225 (N_28225,N_19598,N_15938);
or U28226 (N_28226,N_11177,N_15231);
xor U28227 (N_28227,N_13857,N_10472);
nand U28228 (N_28228,N_18686,N_11296);
and U28229 (N_28229,N_13738,N_18849);
or U28230 (N_28230,N_14396,N_15342);
or U28231 (N_28231,N_10028,N_12106);
nand U28232 (N_28232,N_17865,N_18155);
nand U28233 (N_28233,N_16570,N_11199);
nand U28234 (N_28234,N_14312,N_11156);
and U28235 (N_28235,N_19218,N_12772);
nor U28236 (N_28236,N_13983,N_14304);
or U28237 (N_28237,N_17085,N_10237);
nor U28238 (N_28238,N_12467,N_15303);
or U28239 (N_28239,N_12307,N_13832);
nand U28240 (N_28240,N_17212,N_15230);
and U28241 (N_28241,N_15311,N_10033);
nor U28242 (N_28242,N_17510,N_18339);
nor U28243 (N_28243,N_12402,N_14556);
and U28244 (N_28244,N_16702,N_17238);
nand U28245 (N_28245,N_12622,N_17026);
nand U28246 (N_28246,N_13115,N_14165);
nor U28247 (N_28247,N_19046,N_19913);
and U28248 (N_28248,N_12198,N_10586);
or U28249 (N_28249,N_18033,N_11003);
nand U28250 (N_28250,N_13013,N_17094);
nand U28251 (N_28251,N_10200,N_15564);
nand U28252 (N_28252,N_19602,N_15038);
nor U28253 (N_28253,N_17747,N_16722);
nand U28254 (N_28254,N_17188,N_18835);
and U28255 (N_28255,N_17949,N_10960);
or U28256 (N_28256,N_18473,N_13719);
nand U28257 (N_28257,N_18355,N_19710);
nand U28258 (N_28258,N_11486,N_12057);
and U28259 (N_28259,N_15790,N_16129);
nand U28260 (N_28260,N_12557,N_18481);
nand U28261 (N_28261,N_13804,N_17035);
nor U28262 (N_28262,N_17184,N_11467);
nand U28263 (N_28263,N_14777,N_16702);
nand U28264 (N_28264,N_14304,N_13864);
or U28265 (N_28265,N_17384,N_14477);
nand U28266 (N_28266,N_10438,N_15612);
nand U28267 (N_28267,N_13967,N_16067);
nor U28268 (N_28268,N_18755,N_18576);
and U28269 (N_28269,N_18210,N_11721);
nor U28270 (N_28270,N_11437,N_17304);
or U28271 (N_28271,N_11589,N_19104);
nor U28272 (N_28272,N_11116,N_11476);
nand U28273 (N_28273,N_15461,N_17517);
or U28274 (N_28274,N_16136,N_12567);
and U28275 (N_28275,N_10318,N_16162);
nand U28276 (N_28276,N_17034,N_18394);
and U28277 (N_28277,N_11724,N_16908);
nor U28278 (N_28278,N_19038,N_12824);
or U28279 (N_28279,N_10811,N_10915);
nor U28280 (N_28280,N_18841,N_14037);
or U28281 (N_28281,N_10768,N_14465);
nor U28282 (N_28282,N_11365,N_18558);
nor U28283 (N_28283,N_19981,N_12811);
or U28284 (N_28284,N_19438,N_15544);
nor U28285 (N_28285,N_14650,N_14399);
nand U28286 (N_28286,N_11225,N_17531);
nand U28287 (N_28287,N_17525,N_12679);
nand U28288 (N_28288,N_17671,N_13533);
xnor U28289 (N_28289,N_15760,N_18964);
nor U28290 (N_28290,N_11944,N_14231);
nor U28291 (N_28291,N_15121,N_12300);
nor U28292 (N_28292,N_15953,N_15411);
nand U28293 (N_28293,N_17891,N_18040);
or U28294 (N_28294,N_11994,N_18725);
nor U28295 (N_28295,N_15218,N_13253);
and U28296 (N_28296,N_14532,N_15399);
nand U28297 (N_28297,N_11626,N_12412);
or U28298 (N_28298,N_18512,N_19935);
and U28299 (N_28299,N_19749,N_12033);
or U28300 (N_28300,N_11176,N_18585);
or U28301 (N_28301,N_14101,N_12517);
nand U28302 (N_28302,N_18675,N_11960);
nand U28303 (N_28303,N_13566,N_18132);
nor U28304 (N_28304,N_18892,N_12859);
or U28305 (N_28305,N_11645,N_14504);
nor U28306 (N_28306,N_11996,N_10786);
and U28307 (N_28307,N_10702,N_12310);
or U28308 (N_28308,N_10988,N_13792);
or U28309 (N_28309,N_15733,N_12592);
or U28310 (N_28310,N_14158,N_15482);
nand U28311 (N_28311,N_16040,N_13821);
and U28312 (N_28312,N_18209,N_16534);
nor U28313 (N_28313,N_14827,N_17899);
nand U28314 (N_28314,N_16869,N_11504);
or U28315 (N_28315,N_17822,N_11687);
nand U28316 (N_28316,N_14270,N_11531);
nor U28317 (N_28317,N_15182,N_18604);
nand U28318 (N_28318,N_14295,N_16869);
and U28319 (N_28319,N_18596,N_18455);
or U28320 (N_28320,N_14403,N_10314);
nand U28321 (N_28321,N_18845,N_17252);
and U28322 (N_28322,N_12425,N_16180);
nor U28323 (N_28323,N_19441,N_18305);
nand U28324 (N_28324,N_16525,N_15054);
or U28325 (N_28325,N_13669,N_12269);
or U28326 (N_28326,N_11339,N_12968);
and U28327 (N_28327,N_19016,N_13769);
nor U28328 (N_28328,N_13857,N_14218);
nand U28329 (N_28329,N_17521,N_11556);
nand U28330 (N_28330,N_15239,N_19417);
or U28331 (N_28331,N_12600,N_16721);
nor U28332 (N_28332,N_14758,N_11795);
or U28333 (N_28333,N_17790,N_17114);
and U28334 (N_28334,N_12191,N_14300);
or U28335 (N_28335,N_11559,N_16430);
nand U28336 (N_28336,N_18554,N_19172);
and U28337 (N_28337,N_15586,N_14007);
nor U28338 (N_28338,N_17139,N_18760);
nand U28339 (N_28339,N_14945,N_18342);
or U28340 (N_28340,N_16590,N_11851);
and U28341 (N_28341,N_15394,N_12037);
nand U28342 (N_28342,N_19147,N_14664);
or U28343 (N_28343,N_12164,N_16193);
or U28344 (N_28344,N_14959,N_14616);
or U28345 (N_28345,N_15900,N_18599);
nor U28346 (N_28346,N_13981,N_10939);
nand U28347 (N_28347,N_13447,N_18504);
nor U28348 (N_28348,N_17406,N_15238);
nor U28349 (N_28349,N_14138,N_13074);
nor U28350 (N_28350,N_17033,N_10134);
or U28351 (N_28351,N_15881,N_15269);
and U28352 (N_28352,N_14942,N_17233);
nor U28353 (N_28353,N_12695,N_12288);
nor U28354 (N_28354,N_13365,N_12329);
or U28355 (N_28355,N_13876,N_19972);
nor U28356 (N_28356,N_10713,N_10287);
or U28357 (N_28357,N_10865,N_13328);
and U28358 (N_28358,N_10179,N_18042);
or U28359 (N_28359,N_12795,N_12454);
nor U28360 (N_28360,N_19533,N_18847);
or U28361 (N_28361,N_18316,N_18090);
nor U28362 (N_28362,N_17518,N_17992);
nand U28363 (N_28363,N_10270,N_11509);
nand U28364 (N_28364,N_14591,N_17945);
nor U28365 (N_28365,N_12342,N_19583);
or U28366 (N_28366,N_11935,N_16401);
nand U28367 (N_28367,N_14308,N_18758);
or U28368 (N_28368,N_17270,N_11536);
nand U28369 (N_28369,N_15636,N_17374);
nor U28370 (N_28370,N_18263,N_13510);
and U28371 (N_28371,N_14627,N_19800);
nor U28372 (N_28372,N_16714,N_13596);
and U28373 (N_28373,N_18300,N_17469);
or U28374 (N_28374,N_12099,N_13268);
nand U28375 (N_28375,N_11496,N_13524);
nor U28376 (N_28376,N_15022,N_14911);
and U28377 (N_28377,N_18335,N_13151);
or U28378 (N_28378,N_19002,N_13093);
nand U28379 (N_28379,N_11040,N_15216);
and U28380 (N_28380,N_17786,N_15438);
or U28381 (N_28381,N_10979,N_15835);
nor U28382 (N_28382,N_11356,N_15272);
nand U28383 (N_28383,N_19294,N_17098);
nor U28384 (N_28384,N_11888,N_19683);
nor U28385 (N_28385,N_12927,N_14348);
and U28386 (N_28386,N_11546,N_15037);
or U28387 (N_28387,N_10183,N_16708);
or U28388 (N_28388,N_10906,N_12458);
and U28389 (N_28389,N_19456,N_15941);
nand U28390 (N_28390,N_11370,N_14896);
or U28391 (N_28391,N_19590,N_11260);
nand U28392 (N_28392,N_12091,N_11322);
nor U28393 (N_28393,N_13045,N_14773);
or U28394 (N_28394,N_13501,N_19366);
or U28395 (N_28395,N_17681,N_12370);
nor U28396 (N_28396,N_11690,N_18697);
and U28397 (N_28397,N_19011,N_10075);
nand U28398 (N_28398,N_15477,N_14486);
and U28399 (N_28399,N_10305,N_19376);
or U28400 (N_28400,N_11833,N_11938);
nand U28401 (N_28401,N_13452,N_14199);
or U28402 (N_28402,N_16534,N_10706);
and U28403 (N_28403,N_18314,N_11056);
and U28404 (N_28404,N_15425,N_12846);
or U28405 (N_28405,N_12503,N_15443);
or U28406 (N_28406,N_16385,N_18003);
and U28407 (N_28407,N_11953,N_16189);
and U28408 (N_28408,N_16724,N_11545);
and U28409 (N_28409,N_19835,N_11120);
and U28410 (N_28410,N_13463,N_10632);
nand U28411 (N_28411,N_16845,N_19809);
nor U28412 (N_28412,N_17528,N_13462);
and U28413 (N_28413,N_18280,N_16777);
nand U28414 (N_28414,N_15609,N_13084);
or U28415 (N_28415,N_10942,N_13261);
nor U28416 (N_28416,N_16887,N_17650);
nand U28417 (N_28417,N_17226,N_11363);
nand U28418 (N_28418,N_18551,N_11773);
or U28419 (N_28419,N_16488,N_15545);
nor U28420 (N_28420,N_11054,N_10576);
and U28421 (N_28421,N_14383,N_12755);
or U28422 (N_28422,N_18197,N_18526);
nor U28423 (N_28423,N_16846,N_17480);
or U28424 (N_28424,N_10112,N_16293);
or U28425 (N_28425,N_19297,N_14233);
nand U28426 (N_28426,N_12378,N_18949);
nor U28427 (N_28427,N_12384,N_10890);
or U28428 (N_28428,N_17233,N_11888);
nor U28429 (N_28429,N_12904,N_11752);
nor U28430 (N_28430,N_10087,N_11281);
nand U28431 (N_28431,N_11977,N_16081);
or U28432 (N_28432,N_17458,N_12864);
nor U28433 (N_28433,N_17633,N_15268);
nor U28434 (N_28434,N_12545,N_17809);
and U28435 (N_28435,N_19624,N_12281);
nand U28436 (N_28436,N_16981,N_18366);
and U28437 (N_28437,N_17218,N_19118);
nand U28438 (N_28438,N_10312,N_10562);
and U28439 (N_28439,N_19549,N_16948);
and U28440 (N_28440,N_11047,N_10211);
and U28441 (N_28441,N_10304,N_13658);
or U28442 (N_28442,N_14744,N_16624);
and U28443 (N_28443,N_18246,N_12489);
nand U28444 (N_28444,N_19702,N_17023);
nor U28445 (N_28445,N_15702,N_10345);
nor U28446 (N_28446,N_18281,N_10618);
nand U28447 (N_28447,N_16276,N_15611);
and U28448 (N_28448,N_14259,N_11757);
or U28449 (N_28449,N_14089,N_19250);
and U28450 (N_28450,N_15060,N_16888);
and U28451 (N_28451,N_10835,N_14624);
and U28452 (N_28452,N_11587,N_15697);
or U28453 (N_28453,N_13218,N_12691);
nand U28454 (N_28454,N_10701,N_12677);
or U28455 (N_28455,N_11033,N_11929);
or U28456 (N_28456,N_19319,N_16101);
nand U28457 (N_28457,N_12111,N_16231);
nor U28458 (N_28458,N_15414,N_18223);
nand U28459 (N_28459,N_18946,N_12809);
nand U28460 (N_28460,N_16145,N_19838);
or U28461 (N_28461,N_12636,N_10341);
and U28462 (N_28462,N_15037,N_15571);
or U28463 (N_28463,N_14118,N_18330);
and U28464 (N_28464,N_19704,N_16922);
and U28465 (N_28465,N_16991,N_10104);
nor U28466 (N_28466,N_18804,N_15983);
nor U28467 (N_28467,N_10501,N_10070);
nor U28468 (N_28468,N_12633,N_15675);
nor U28469 (N_28469,N_13217,N_15694);
and U28470 (N_28470,N_13250,N_12866);
or U28471 (N_28471,N_18805,N_16664);
nand U28472 (N_28472,N_15604,N_13525);
and U28473 (N_28473,N_16872,N_11068);
nand U28474 (N_28474,N_11015,N_19016);
nand U28475 (N_28475,N_14365,N_13081);
or U28476 (N_28476,N_19702,N_11740);
nand U28477 (N_28477,N_17320,N_16167);
nor U28478 (N_28478,N_14042,N_10128);
or U28479 (N_28479,N_10920,N_15832);
nor U28480 (N_28480,N_13826,N_13172);
nand U28481 (N_28481,N_10178,N_14990);
nor U28482 (N_28482,N_12752,N_18986);
nand U28483 (N_28483,N_13550,N_17411);
or U28484 (N_28484,N_10913,N_18286);
nand U28485 (N_28485,N_19673,N_14434);
nand U28486 (N_28486,N_15458,N_10723);
nand U28487 (N_28487,N_11639,N_14459);
nand U28488 (N_28488,N_12715,N_19867);
nand U28489 (N_28489,N_15848,N_17078);
and U28490 (N_28490,N_18285,N_10725);
nand U28491 (N_28491,N_17226,N_19998);
nand U28492 (N_28492,N_17877,N_19058);
or U28493 (N_28493,N_16797,N_10605);
or U28494 (N_28494,N_10144,N_15802);
nand U28495 (N_28495,N_10502,N_14144);
or U28496 (N_28496,N_15065,N_19934);
nand U28497 (N_28497,N_16525,N_16646);
nand U28498 (N_28498,N_18679,N_14352);
and U28499 (N_28499,N_15935,N_12453);
or U28500 (N_28500,N_12829,N_11757);
nand U28501 (N_28501,N_18246,N_11939);
and U28502 (N_28502,N_19421,N_19761);
nor U28503 (N_28503,N_17089,N_15844);
and U28504 (N_28504,N_11516,N_15432);
or U28505 (N_28505,N_13149,N_16357);
and U28506 (N_28506,N_16122,N_10556);
nor U28507 (N_28507,N_19130,N_19636);
and U28508 (N_28508,N_18265,N_14861);
nor U28509 (N_28509,N_13329,N_19070);
xnor U28510 (N_28510,N_19766,N_14328);
and U28511 (N_28511,N_11429,N_15170);
or U28512 (N_28512,N_14102,N_12770);
or U28513 (N_28513,N_16851,N_10222);
or U28514 (N_28514,N_12972,N_17903);
or U28515 (N_28515,N_17590,N_10031);
nand U28516 (N_28516,N_16424,N_15673);
nor U28517 (N_28517,N_15299,N_19181);
and U28518 (N_28518,N_10005,N_19821);
or U28519 (N_28519,N_15006,N_18679);
xor U28520 (N_28520,N_10856,N_17523);
and U28521 (N_28521,N_15537,N_14741);
and U28522 (N_28522,N_15116,N_17026);
and U28523 (N_28523,N_12684,N_17989);
and U28524 (N_28524,N_12806,N_10550);
nand U28525 (N_28525,N_15082,N_14378);
nand U28526 (N_28526,N_18302,N_18740);
and U28527 (N_28527,N_19165,N_10730);
or U28528 (N_28528,N_13708,N_11501);
or U28529 (N_28529,N_19548,N_19977);
or U28530 (N_28530,N_11939,N_12660);
nor U28531 (N_28531,N_13512,N_19715);
or U28532 (N_28532,N_12981,N_18349);
or U28533 (N_28533,N_19235,N_10135);
nand U28534 (N_28534,N_17428,N_12506);
or U28535 (N_28535,N_11014,N_14023);
and U28536 (N_28536,N_19875,N_17196);
nand U28537 (N_28537,N_14387,N_18561);
or U28538 (N_28538,N_19665,N_14376);
nand U28539 (N_28539,N_17327,N_11341);
nand U28540 (N_28540,N_17666,N_15692);
or U28541 (N_28541,N_10741,N_18709);
or U28542 (N_28542,N_17679,N_18568);
nor U28543 (N_28543,N_16226,N_18845);
nand U28544 (N_28544,N_17758,N_14271);
nor U28545 (N_28545,N_10145,N_11947);
nand U28546 (N_28546,N_15783,N_13133);
nor U28547 (N_28547,N_15433,N_14490);
nand U28548 (N_28548,N_11762,N_11216);
nor U28549 (N_28549,N_10691,N_18297);
and U28550 (N_28550,N_10897,N_13981);
nand U28551 (N_28551,N_14254,N_10245);
nor U28552 (N_28552,N_11008,N_12895);
xnor U28553 (N_28553,N_12402,N_19154);
nand U28554 (N_28554,N_13708,N_18368);
and U28555 (N_28555,N_12494,N_13396);
or U28556 (N_28556,N_17113,N_10076);
nand U28557 (N_28557,N_13782,N_19858);
nand U28558 (N_28558,N_17522,N_19768);
and U28559 (N_28559,N_13716,N_12650);
and U28560 (N_28560,N_17421,N_16363);
or U28561 (N_28561,N_15499,N_10809);
or U28562 (N_28562,N_10134,N_16248);
and U28563 (N_28563,N_19391,N_16046);
nand U28564 (N_28564,N_11327,N_13395);
and U28565 (N_28565,N_13618,N_12444);
nor U28566 (N_28566,N_17184,N_19044);
nor U28567 (N_28567,N_13770,N_13186);
nor U28568 (N_28568,N_10729,N_18311);
or U28569 (N_28569,N_14041,N_10682);
and U28570 (N_28570,N_10179,N_10975);
and U28571 (N_28571,N_11636,N_17372);
nor U28572 (N_28572,N_17323,N_18507);
or U28573 (N_28573,N_11410,N_15621);
and U28574 (N_28574,N_19128,N_17713);
or U28575 (N_28575,N_15771,N_12111);
nand U28576 (N_28576,N_16398,N_11413);
nand U28577 (N_28577,N_16753,N_15070);
or U28578 (N_28578,N_10218,N_19450);
nor U28579 (N_28579,N_13533,N_17717);
or U28580 (N_28580,N_17897,N_11363);
and U28581 (N_28581,N_13230,N_18787);
nor U28582 (N_28582,N_10218,N_17697);
and U28583 (N_28583,N_15358,N_18106);
or U28584 (N_28584,N_11952,N_13833);
nor U28585 (N_28585,N_13155,N_17135);
and U28586 (N_28586,N_12617,N_11051);
nand U28587 (N_28587,N_17376,N_12533);
nand U28588 (N_28588,N_16865,N_13130);
nand U28589 (N_28589,N_17750,N_13262);
nor U28590 (N_28590,N_14977,N_14831);
or U28591 (N_28591,N_13727,N_12254);
nor U28592 (N_28592,N_19708,N_16159);
and U28593 (N_28593,N_17964,N_18383);
nor U28594 (N_28594,N_18448,N_16556);
or U28595 (N_28595,N_19946,N_14381);
and U28596 (N_28596,N_14691,N_14310);
nand U28597 (N_28597,N_14884,N_12218);
and U28598 (N_28598,N_16960,N_10694);
or U28599 (N_28599,N_11481,N_15341);
or U28600 (N_28600,N_11765,N_19648);
nand U28601 (N_28601,N_13652,N_14407);
nand U28602 (N_28602,N_14003,N_13295);
nor U28603 (N_28603,N_19944,N_16642);
nand U28604 (N_28604,N_14656,N_19391);
nor U28605 (N_28605,N_13591,N_15727);
or U28606 (N_28606,N_10718,N_18908);
nor U28607 (N_28607,N_16981,N_12632);
nor U28608 (N_28608,N_10351,N_19117);
nor U28609 (N_28609,N_12329,N_16239);
nor U28610 (N_28610,N_18933,N_13250);
nor U28611 (N_28611,N_17357,N_11525);
nand U28612 (N_28612,N_13527,N_14358);
or U28613 (N_28613,N_18108,N_18686);
or U28614 (N_28614,N_11641,N_16779);
xnor U28615 (N_28615,N_19065,N_14063);
or U28616 (N_28616,N_15047,N_16653);
nand U28617 (N_28617,N_14597,N_18429);
nand U28618 (N_28618,N_13529,N_12393);
nand U28619 (N_28619,N_11301,N_18906);
or U28620 (N_28620,N_16870,N_12944);
nand U28621 (N_28621,N_16951,N_13765);
nand U28622 (N_28622,N_12924,N_19423);
and U28623 (N_28623,N_11680,N_18279);
and U28624 (N_28624,N_14969,N_11210);
nand U28625 (N_28625,N_11462,N_12870);
nand U28626 (N_28626,N_11130,N_10824);
or U28627 (N_28627,N_12136,N_19224);
or U28628 (N_28628,N_12601,N_13400);
nand U28629 (N_28629,N_15117,N_10704);
and U28630 (N_28630,N_17397,N_12540);
nor U28631 (N_28631,N_19057,N_18938);
and U28632 (N_28632,N_14723,N_10185);
nor U28633 (N_28633,N_18212,N_11870);
and U28634 (N_28634,N_17747,N_10645);
or U28635 (N_28635,N_14657,N_10527);
nor U28636 (N_28636,N_11919,N_14399);
nor U28637 (N_28637,N_15898,N_10409);
or U28638 (N_28638,N_14242,N_16435);
or U28639 (N_28639,N_15743,N_16221);
nor U28640 (N_28640,N_16731,N_16758);
xor U28641 (N_28641,N_15383,N_11380);
or U28642 (N_28642,N_19408,N_19370);
nand U28643 (N_28643,N_12952,N_13176);
or U28644 (N_28644,N_10483,N_17930);
and U28645 (N_28645,N_16332,N_15405);
nand U28646 (N_28646,N_15402,N_18340);
or U28647 (N_28647,N_12617,N_16892);
nor U28648 (N_28648,N_14017,N_18050);
and U28649 (N_28649,N_19306,N_16212);
and U28650 (N_28650,N_14781,N_14266);
nor U28651 (N_28651,N_18048,N_13891);
nand U28652 (N_28652,N_14041,N_12808);
nor U28653 (N_28653,N_19964,N_12772);
or U28654 (N_28654,N_17598,N_15645);
and U28655 (N_28655,N_17502,N_18498);
nand U28656 (N_28656,N_19761,N_15852);
nor U28657 (N_28657,N_16506,N_15393);
and U28658 (N_28658,N_16604,N_18982);
or U28659 (N_28659,N_13628,N_17806);
nor U28660 (N_28660,N_17673,N_11322);
and U28661 (N_28661,N_12684,N_14066);
or U28662 (N_28662,N_13762,N_17857);
nor U28663 (N_28663,N_17754,N_10817);
or U28664 (N_28664,N_12655,N_14623);
or U28665 (N_28665,N_18969,N_18088);
and U28666 (N_28666,N_11299,N_16492);
nor U28667 (N_28667,N_16232,N_16844);
and U28668 (N_28668,N_10081,N_17341);
nor U28669 (N_28669,N_19918,N_11114);
nor U28670 (N_28670,N_19790,N_13406);
and U28671 (N_28671,N_13258,N_11853);
and U28672 (N_28672,N_17946,N_10287);
nor U28673 (N_28673,N_19584,N_16039);
or U28674 (N_28674,N_16784,N_16561);
nand U28675 (N_28675,N_17027,N_10225);
xnor U28676 (N_28676,N_16752,N_14496);
nor U28677 (N_28677,N_13125,N_13010);
or U28678 (N_28678,N_18923,N_16650);
nand U28679 (N_28679,N_14230,N_16932);
or U28680 (N_28680,N_19258,N_13310);
or U28681 (N_28681,N_12875,N_10397);
or U28682 (N_28682,N_12918,N_10640);
nor U28683 (N_28683,N_15695,N_19827);
and U28684 (N_28684,N_16431,N_16836);
or U28685 (N_28685,N_10805,N_10505);
nand U28686 (N_28686,N_12607,N_14853);
nor U28687 (N_28687,N_11496,N_16036);
nor U28688 (N_28688,N_13872,N_17275);
nand U28689 (N_28689,N_15870,N_15873);
and U28690 (N_28690,N_10047,N_11932);
nor U28691 (N_28691,N_18374,N_18129);
nor U28692 (N_28692,N_11035,N_15817);
nand U28693 (N_28693,N_12607,N_11165);
or U28694 (N_28694,N_16920,N_16982);
or U28695 (N_28695,N_16290,N_12210);
and U28696 (N_28696,N_11193,N_13634);
and U28697 (N_28697,N_12210,N_11840);
or U28698 (N_28698,N_12928,N_15340);
or U28699 (N_28699,N_17039,N_16093);
or U28700 (N_28700,N_19357,N_13377);
nor U28701 (N_28701,N_10037,N_11570);
nand U28702 (N_28702,N_15943,N_18462);
nand U28703 (N_28703,N_10121,N_17057);
or U28704 (N_28704,N_12353,N_18889);
or U28705 (N_28705,N_16308,N_10238);
nor U28706 (N_28706,N_12280,N_15789);
nor U28707 (N_28707,N_12611,N_19832);
and U28708 (N_28708,N_18008,N_18208);
or U28709 (N_28709,N_11357,N_11810);
or U28710 (N_28710,N_19466,N_18250);
nor U28711 (N_28711,N_18261,N_13412);
nand U28712 (N_28712,N_11976,N_12515);
nand U28713 (N_28713,N_13334,N_11917);
and U28714 (N_28714,N_11008,N_18172);
and U28715 (N_28715,N_13560,N_10383);
nand U28716 (N_28716,N_10213,N_15413);
nand U28717 (N_28717,N_14588,N_10021);
and U28718 (N_28718,N_19276,N_18732);
nand U28719 (N_28719,N_16765,N_17792);
nor U28720 (N_28720,N_17184,N_10660);
nor U28721 (N_28721,N_16403,N_13798);
and U28722 (N_28722,N_10514,N_16854);
nand U28723 (N_28723,N_14126,N_18507);
nor U28724 (N_28724,N_10705,N_17318);
or U28725 (N_28725,N_16749,N_13823);
nor U28726 (N_28726,N_12851,N_17229);
and U28727 (N_28727,N_10155,N_16486);
nor U28728 (N_28728,N_16720,N_16423);
nor U28729 (N_28729,N_12091,N_19687);
or U28730 (N_28730,N_19201,N_12897);
or U28731 (N_28731,N_19435,N_10619);
nand U28732 (N_28732,N_15795,N_14958);
and U28733 (N_28733,N_11766,N_18298);
nor U28734 (N_28734,N_12991,N_13114);
nand U28735 (N_28735,N_11527,N_12619);
nand U28736 (N_28736,N_19754,N_14576);
and U28737 (N_28737,N_12816,N_10080);
xnor U28738 (N_28738,N_14436,N_11909);
and U28739 (N_28739,N_11333,N_12788);
xor U28740 (N_28740,N_12545,N_14779);
nand U28741 (N_28741,N_13336,N_15194);
and U28742 (N_28742,N_17585,N_19530);
or U28743 (N_28743,N_17899,N_14457);
or U28744 (N_28744,N_19970,N_16936);
nand U28745 (N_28745,N_19699,N_10634);
or U28746 (N_28746,N_10327,N_16761);
or U28747 (N_28747,N_11589,N_12919);
nand U28748 (N_28748,N_10161,N_11829);
nand U28749 (N_28749,N_12862,N_19674);
nor U28750 (N_28750,N_14733,N_18536);
nand U28751 (N_28751,N_12452,N_16101);
or U28752 (N_28752,N_18770,N_14256);
nor U28753 (N_28753,N_18845,N_13227);
nor U28754 (N_28754,N_18471,N_16723);
or U28755 (N_28755,N_17052,N_16717);
nand U28756 (N_28756,N_12937,N_17160);
or U28757 (N_28757,N_16130,N_18947);
and U28758 (N_28758,N_15208,N_16647);
nand U28759 (N_28759,N_11623,N_13924);
nand U28760 (N_28760,N_10948,N_10784);
or U28761 (N_28761,N_15322,N_13421);
nor U28762 (N_28762,N_18634,N_11840);
nor U28763 (N_28763,N_10714,N_17962);
xor U28764 (N_28764,N_16393,N_18417);
or U28765 (N_28765,N_19822,N_11587);
and U28766 (N_28766,N_14567,N_16501);
and U28767 (N_28767,N_15900,N_16616);
or U28768 (N_28768,N_15535,N_13486);
nor U28769 (N_28769,N_18464,N_10959);
nor U28770 (N_28770,N_19991,N_11772);
nand U28771 (N_28771,N_12680,N_16613);
nand U28772 (N_28772,N_19973,N_13764);
and U28773 (N_28773,N_13343,N_19336);
or U28774 (N_28774,N_15774,N_15359);
and U28775 (N_28775,N_18591,N_19085);
nor U28776 (N_28776,N_18335,N_16990);
nand U28777 (N_28777,N_11877,N_11737);
nor U28778 (N_28778,N_17403,N_18628);
and U28779 (N_28779,N_13531,N_12211);
nand U28780 (N_28780,N_17796,N_15339);
and U28781 (N_28781,N_10200,N_13111);
nand U28782 (N_28782,N_13262,N_10956);
and U28783 (N_28783,N_12662,N_14913);
nor U28784 (N_28784,N_13948,N_12117);
nor U28785 (N_28785,N_14368,N_19756);
nor U28786 (N_28786,N_14299,N_13432);
nand U28787 (N_28787,N_15260,N_13168);
and U28788 (N_28788,N_11436,N_10101);
or U28789 (N_28789,N_14827,N_16444);
and U28790 (N_28790,N_14352,N_17609);
nor U28791 (N_28791,N_13359,N_16372);
or U28792 (N_28792,N_12463,N_11636);
and U28793 (N_28793,N_19474,N_11188);
or U28794 (N_28794,N_10078,N_17830);
and U28795 (N_28795,N_18353,N_12216);
and U28796 (N_28796,N_10797,N_16144);
nor U28797 (N_28797,N_18430,N_18104);
xor U28798 (N_28798,N_13172,N_17104);
and U28799 (N_28799,N_17657,N_12800);
nand U28800 (N_28800,N_18097,N_19738);
or U28801 (N_28801,N_14167,N_16610);
nand U28802 (N_28802,N_18670,N_15568);
or U28803 (N_28803,N_13769,N_17142);
nand U28804 (N_28804,N_15452,N_16803);
nor U28805 (N_28805,N_10561,N_15571);
or U28806 (N_28806,N_19424,N_10828);
nor U28807 (N_28807,N_14671,N_13414);
and U28808 (N_28808,N_12223,N_10576);
and U28809 (N_28809,N_18157,N_18116);
xor U28810 (N_28810,N_10259,N_11412);
or U28811 (N_28811,N_14568,N_19691);
nand U28812 (N_28812,N_16301,N_19961);
nor U28813 (N_28813,N_10912,N_13773);
nor U28814 (N_28814,N_11775,N_12836);
or U28815 (N_28815,N_12967,N_19145);
nand U28816 (N_28816,N_14151,N_13788);
or U28817 (N_28817,N_15804,N_16880);
nand U28818 (N_28818,N_14795,N_14401);
nor U28819 (N_28819,N_17430,N_18111);
nor U28820 (N_28820,N_10240,N_16394);
nor U28821 (N_28821,N_16438,N_12076);
or U28822 (N_28822,N_16040,N_11347);
nand U28823 (N_28823,N_16353,N_16157);
nor U28824 (N_28824,N_19318,N_18983);
nor U28825 (N_28825,N_11419,N_15634);
or U28826 (N_28826,N_14768,N_17547);
nor U28827 (N_28827,N_12621,N_17747);
nor U28828 (N_28828,N_13817,N_12053);
nand U28829 (N_28829,N_13690,N_19456);
nor U28830 (N_28830,N_12286,N_17158);
nor U28831 (N_28831,N_19807,N_17505);
nor U28832 (N_28832,N_11414,N_19899);
and U28833 (N_28833,N_12958,N_15321);
or U28834 (N_28834,N_14917,N_16571);
or U28835 (N_28835,N_16378,N_14230);
nor U28836 (N_28836,N_10608,N_19030);
and U28837 (N_28837,N_16873,N_10502);
or U28838 (N_28838,N_10349,N_12560);
nand U28839 (N_28839,N_12586,N_15675);
and U28840 (N_28840,N_17640,N_17333);
nand U28841 (N_28841,N_14041,N_13621);
nor U28842 (N_28842,N_13293,N_13455);
nor U28843 (N_28843,N_12563,N_17301);
xnor U28844 (N_28844,N_11535,N_17616);
or U28845 (N_28845,N_13166,N_14867);
xor U28846 (N_28846,N_14784,N_15655);
nor U28847 (N_28847,N_11008,N_11287);
nand U28848 (N_28848,N_18348,N_14921);
nor U28849 (N_28849,N_16919,N_16159);
and U28850 (N_28850,N_11582,N_16621);
or U28851 (N_28851,N_17904,N_11980);
and U28852 (N_28852,N_17647,N_11992);
and U28853 (N_28853,N_15570,N_12692);
xnor U28854 (N_28854,N_14638,N_12464);
nor U28855 (N_28855,N_13446,N_11127);
nand U28856 (N_28856,N_19630,N_17145);
nand U28857 (N_28857,N_13766,N_11920);
nand U28858 (N_28858,N_11037,N_19229);
nand U28859 (N_28859,N_11008,N_15767);
nand U28860 (N_28860,N_12255,N_14044);
or U28861 (N_28861,N_12048,N_17229);
or U28862 (N_28862,N_15949,N_12274);
nor U28863 (N_28863,N_14624,N_17655);
nand U28864 (N_28864,N_16492,N_11103);
nand U28865 (N_28865,N_17093,N_12746);
nand U28866 (N_28866,N_16013,N_17869);
and U28867 (N_28867,N_12635,N_13072);
or U28868 (N_28868,N_14979,N_12665);
nor U28869 (N_28869,N_11176,N_12332);
or U28870 (N_28870,N_17350,N_18251);
or U28871 (N_28871,N_15995,N_16291);
nor U28872 (N_28872,N_14766,N_13416);
nor U28873 (N_28873,N_17172,N_14553);
or U28874 (N_28874,N_19318,N_14160);
or U28875 (N_28875,N_15238,N_12195);
nor U28876 (N_28876,N_13818,N_10417);
nand U28877 (N_28877,N_19022,N_15095);
nor U28878 (N_28878,N_19808,N_10328);
nand U28879 (N_28879,N_17039,N_17678);
or U28880 (N_28880,N_16674,N_19337);
nand U28881 (N_28881,N_13818,N_15310);
nand U28882 (N_28882,N_10818,N_11264);
nor U28883 (N_28883,N_10215,N_12017);
nand U28884 (N_28884,N_16475,N_16080);
nand U28885 (N_28885,N_11840,N_15214);
nand U28886 (N_28886,N_12414,N_11193);
nand U28887 (N_28887,N_11166,N_18970);
and U28888 (N_28888,N_11936,N_13576);
nor U28889 (N_28889,N_18489,N_11722);
or U28890 (N_28890,N_14645,N_10991);
nor U28891 (N_28891,N_18588,N_13629);
or U28892 (N_28892,N_15035,N_12651);
or U28893 (N_28893,N_18112,N_11738);
nand U28894 (N_28894,N_15789,N_19857);
or U28895 (N_28895,N_11689,N_17571);
nor U28896 (N_28896,N_14814,N_13552);
and U28897 (N_28897,N_13519,N_17360);
and U28898 (N_28898,N_18391,N_12136);
nor U28899 (N_28899,N_13692,N_19713);
nor U28900 (N_28900,N_19223,N_18578);
and U28901 (N_28901,N_17282,N_12153);
and U28902 (N_28902,N_13650,N_12455);
xnor U28903 (N_28903,N_10859,N_11136);
nor U28904 (N_28904,N_13513,N_16843);
or U28905 (N_28905,N_10039,N_14710);
nand U28906 (N_28906,N_13316,N_14844);
nand U28907 (N_28907,N_14804,N_14644);
nor U28908 (N_28908,N_15582,N_14945);
nand U28909 (N_28909,N_19849,N_13493);
and U28910 (N_28910,N_14389,N_18962);
nand U28911 (N_28911,N_11731,N_16674);
and U28912 (N_28912,N_12418,N_10412);
or U28913 (N_28913,N_17914,N_15488);
nor U28914 (N_28914,N_16420,N_13014);
nor U28915 (N_28915,N_14781,N_17901);
or U28916 (N_28916,N_11475,N_11413);
or U28917 (N_28917,N_15808,N_15138);
nor U28918 (N_28918,N_13249,N_15123);
and U28919 (N_28919,N_17120,N_13976);
and U28920 (N_28920,N_17849,N_18605);
nor U28921 (N_28921,N_10118,N_15939);
or U28922 (N_28922,N_15947,N_15458);
and U28923 (N_28923,N_10516,N_10104);
or U28924 (N_28924,N_19865,N_16443);
nor U28925 (N_28925,N_16417,N_18626);
and U28926 (N_28926,N_18159,N_16358);
nand U28927 (N_28927,N_15903,N_18887);
or U28928 (N_28928,N_16547,N_17192);
nand U28929 (N_28929,N_12421,N_14259);
nand U28930 (N_28930,N_16638,N_10537);
nor U28931 (N_28931,N_17781,N_19231);
and U28932 (N_28932,N_16432,N_10032);
nand U28933 (N_28933,N_15624,N_15015);
nand U28934 (N_28934,N_16683,N_14506);
nand U28935 (N_28935,N_15651,N_12987);
and U28936 (N_28936,N_15008,N_19907);
nand U28937 (N_28937,N_14372,N_19559);
or U28938 (N_28938,N_13057,N_19911);
and U28939 (N_28939,N_12032,N_13204);
or U28940 (N_28940,N_11241,N_19127);
nor U28941 (N_28941,N_14402,N_17918);
nor U28942 (N_28942,N_12025,N_16337);
and U28943 (N_28943,N_16130,N_12095);
or U28944 (N_28944,N_16551,N_11979);
or U28945 (N_28945,N_19525,N_11312);
or U28946 (N_28946,N_19750,N_11070);
nor U28947 (N_28947,N_15201,N_11255);
or U28948 (N_28948,N_19810,N_14439);
or U28949 (N_28949,N_12787,N_16254);
nor U28950 (N_28950,N_17978,N_17499);
and U28951 (N_28951,N_17542,N_17527);
nand U28952 (N_28952,N_16317,N_15581);
nor U28953 (N_28953,N_19063,N_15031);
and U28954 (N_28954,N_13387,N_16522);
nor U28955 (N_28955,N_11580,N_14824);
nor U28956 (N_28956,N_11820,N_15771);
nand U28957 (N_28957,N_14041,N_16735);
or U28958 (N_28958,N_12876,N_17395);
xor U28959 (N_28959,N_15197,N_15136);
or U28960 (N_28960,N_11618,N_18628);
nor U28961 (N_28961,N_11588,N_12521);
nand U28962 (N_28962,N_15781,N_12125);
nor U28963 (N_28963,N_18090,N_10778);
nand U28964 (N_28964,N_13850,N_15253);
nor U28965 (N_28965,N_17408,N_16208);
and U28966 (N_28966,N_12579,N_14848);
nor U28967 (N_28967,N_16308,N_10720);
and U28968 (N_28968,N_12918,N_13197);
nor U28969 (N_28969,N_15138,N_16445);
and U28970 (N_28970,N_18895,N_17736);
nor U28971 (N_28971,N_16843,N_18934);
nand U28972 (N_28972,N_12861,N_17250);
and U28973 (N_28973,N_16650,N_10721);
or U28974 (N_28974,N_14231,N_14684);
nand U28975 (N_28975,N_18544,N_15100);
nand U28976 (N_28976,N_11492,N_16860);
nand U28977 (N_28977,N_16941,N_11959);
and U28978 (N_28978,N_11040,N_17787);
nor U28979 (N_28979,N_15508,N_16697);
and U28980 (N_28980,N_14636,N_10630);
nor U28981 (N_28981,N_19795,N_14006);
or U28982 (N_28982,N_12182,N_19421);
nand U28983 (N_28983,N_12944,N_19321);
and U28984 (N_28984,N_14937,N_19264);
or U28985 (N_28985,N_18339,N_12450);
xnor U28986 (N_28986,N_12480,N_17534);
and U28987 (N_28987,N_13392,N_12057);
nor U28988 (N_28988,N_12362,N_19108);
nand U28989 (N_28989,N_13509,N_10127);
nor U28990 (N_28990,N_14442,N_12154);
nor U28991 (N_28991,N_11566,N_11386);
nand U28992 (N_28992,N_10661,N_13644);
or U28993 (N_28993,N_10666,N_15825);
and U28994 (N_28994,N_13850,N_14061);
and U28995 (N_28995,N_12119,N_12932);
and U28996 (N_28996,N_14464,N_16474);
or U28997 (N_28997,N_17250,N_14724);
nor U28998 (N_28998,N_19053,N_12714);
nor U28999 (N_28999,N_18211,N_19374);
nor U29000 (N_29000,N_13252,N_14911);
nor U29001 (N_29001,N_13394,N_13717);
nor U29002 (N_29002,N_10521,N_17337);
and U29003 (N_29003,N_11295,N_16794);
nand U29004 (N_29004,N_15986,N_13475);
or U29005 (N_29005,N_10553,N_19787);
and U29006 (N_29006,N_19139,N_10315);
nor U29007 (N_29007,N_17013,N_14792);
or U29008 (N_29008,N_10904,N_13267);
nand U29009 (N_29009,N_10525,N_19579);
or U29010 (N_29010,N_16450,N_14362);
and U29011 (N_29011,N_13730,N_13403);
nor U29012 (N_29012,N_10730,N_14869);
nand U29013 (N_29013,N_11929,N_16330);
nand U29014 (N_29014,N_19153,N_17717);
nand U29015 (N_29015,N_12400,N_19408);
nor U29016 (N_29016,N_10131,N_11754);
nand U29017 (N_29017,N_19673,N_18535);
or U29018 (N_29018,N_16353,N_12168);
nand U29019 (N_29019,N_19195,N_16699);
or U29020 (N_29020,N_18968,N_11651);
nand U29021 (N_29021,N_10997,N_10555);
and U29022 (N_29022,N_19891,N_14863);
nand U29023 (N_29023,N_15105,N_19580);
or U29024 (N_29024,N_14557,N_19419);
or U29025 (N_29025,N_18032,N_17956);
nand U29026 (N_29026,N_17502,N_11305);
and U29027 (N_29027,N_19256,N_11361);
nor U29028 (N_29028,N_11866,N_15393);
and U29029 (N_29029,N_12847,N_18851);
nand U29030 (N_29030,N_19395,N_17333);
nand U29031 (N_29031,N_10613,N_19718);
nand U29032 (N_29032,N_11678,N_18382);
or U29033 (N_29033,N_19264,N_14690);
and U29034 (N_29034,N_15046,N_14977);
nand U29035 (N_29035,N_15644,N_11749);
nor U29036 (N_29036,N_18967,N_13988);
or U29037 (N_29037,N_15528,N_16055);
nand U29038 (N_29038,N_15522,N_17865);
nand U29039 (N_29039,N_11371,N_16370);
nor U29040 (N_29040,N_11430,N_11914);
nand U29041 (N_29041,N_13876,N_14416);
and U29042 (N_29042,N_16104,N_12345);
nor U29043 (N_29043,N_19751,N_12317);
nand U29044 (N_29044,N_11686,N_13694);
or U29045 (N_29045,N_15051,N_16693);
nor U29046 (N_29046,N_18163,N_16975);
nor U29047 (N_29047,N_13537,N_12724);
or U29048 (N_29048,N_10785,N_13344);
and U29049 (N_29049,N_12294,N_11274);
nand U29050 (N_29050,N_10579,N_15329);
and U29051 (N_29051,N_16720,N_17797);
or U29052 (N_29052,N_14922,N_16934);
and U29053 (N_29053,N_15014,N_18909);
nand U29054 (N_29054,N_19695,N_11952);
or U29055 (N_29055,N_16052,N_18164);
nand U29056 (N_29056,N_17973,N_15106);
nand U29057 (N_29057,N_17943,N_15702);
nand U29058 (N_29058,N_12857,N_13621);
nand U29059 (N_29059,N_13047,N_12692);
nand U29060 (N_29060,N_18577,N_12424);
or U29061 (N_29061,N_12097,N_13888);
and U29062 (N_29062,N_16299,N_17588);
and U29063 (N_29063,N_13436,N_11493);
or U29064 (N_29064,N_10121,N_12587);
nor U29065 (N_29065,N_14947,N_14297);
or U29066 (N_29066,N_10757,N_17987);
nor U29067 (N_29067,N_17423,N_11503);
and U29068 (N_29068,N_15171,N_16964);
nor U29069 (N_29069,N_18627,N_14911);
or U29070 (N_29070,N_10762,N_18141);
nand U29071 (N_29071,N_17445,N_12113);
or U29072 (N_29072,N_13488,N_15081);
nor U29073 (N_29073,N_13569,N_13616);
and U29074 (N_29074,N_18300,N_13158);
nor U29075 (N_29075,N_12764,N_15128);
xnor U29076 (N_29076,N_19305,N_13944);
nor U29077 (N_29077,N_18593,N_17638);
nor U29078 (N_29078,N_19435,N_15633);
and U29079 (N_29079,N_15937,N_12627);
and U29080 (N_29080,N_14910,N_16678);
or U29081 (N_29081,N_11550,N_14317);
nor U29082 (N_29082,N_15933,N_14266);
or U29083 (N_29083,N_13942,N_12958);
nand U29084 (N_29084,N_10376,N_13099);
and U29085 (N_29085,N_18670,N_16829);
or U29086 (N_29086,N_14014,N_17616);
or U29087 (N_29087,N_16151,N_10594);
nand U29088 (N_29088,N_16236,N_11115);
nand U29089 (N_29089,N_16476,N_19690);
or U29090 (N_29090,N_12969,N_14733);
nor U29091 (N_29091,N_18077,N_19693);
or U29092 (N_29092,N_18052,N_14500);
nand U29093 (N_29093,N_10285,N_14126);
or U29094 (N_29094,N_16271,N_15842);
or U29095 (N_29095,N_13461,N_17348);
nor U29096 (N_29096,N_15791,N_12845);
or U29097 (N_29097,N_10400,N_15182);
nand U29098 (N_29098,N_16862,N_19725);
nor U29099 (N_29099,N_10772,N_14584);
or U29100 (N_29100,N_18714,N_11843);
or U29101 (N_29101,N_15435,N_13013);
nor U29102 (N_29102,N_13716,N_15651);
xor U29103 (N_29103,N_13667,N_12696);
nand U29104 (N_29104,N_14121,N_19456);
or U29105 (N_29105,N_14704,N_17762);
and U29106 (N_29106,N_12033,N_11618);
and U29107 (N_29107,N_18816,N_18865);
nor U29108 (N_29108,N_18220,N_10808);
nand U29109 (N_29109,N_19300,N_15929);
nor U29110 (N_29110,N_16676,N_13961);
nand U29111 (N_29111,N_16489,N_15432);
nand U29112 (N_29112,N_11175,N_16845);
and U29113 (N_29113,N_12600,N_12331);
and U29114 (N_29114,N_11997,N_16739);
and U29115 (N_29115,N_14262,N_16073);
nor U29116 (N_29116,N_12650,N_19467);
nand U29117 (N_29117,N_12599,N_10666);
nor U29118 (N_29118,N_17598,N_14381);
nor U29119 (N_29119,N_18431,N_17833);
nand U29120 (N_29120,N_14678,N_18188);
and U29121 (N_29121,N_15262,N_13621);
nand U29122 (N_29122,N_18081,N_14343);
or U29123 (N_29123,N_11180,N_15411);
or U29124 (N_29124,N_12903,N_11970);
nor U29125 (N_29125,N_17984,N_14542);
or U29126 (N_29126,N_12843,N_19969);
or U29127 (N_29127,N_17639,N_16922);
or U29128 (N_29128,N_17114,N_18760);
nor U29129 (N_29129,N_14755,N_10724);
nor U29130 (N_29130,N_15728,N_12136);
nand U29131 (N_29131,N_15681,N_18066);
or U29132 (N_29132,N_14248,N_11352);
and U29133 (N_29133,N_17466,N_13688);
nor U29134 (N_29134,N_16703,N_11673);
nand U29135 (N_29135,N_16929,N_10705);
nand U29136 (N_29136,N_16215,N_14711);
nor U29137 (N_29137,N_19138,N_16138);
and U29138 (N_29138,N_17106,N_18757);
nor U29139 (N_29139,N_17272,N_16389);
nor U29140 (N_29140,N_18764,N_11252);
nand U29141 (N_29141,N_11266,N_18141);
and U29142 (N_29142,N_17424,N_16595);
and U29143 (N_29143,N_16323,N_18811);
or U29144 (N_29144,N_17570,N_17846);
nand U29145 (N_29145,N_16882,N_17423);
or U29146 (N_29146,N_14939,N_13301);
nor U29147 (N_29147,N_16846,N_10483);
and U29148 (N_29148,N_18015,N_17258);
or U29149 (N_29149,N_17126,N_15996);
nor U29150 (N_29150,N_17089,N_13344);
or U29151 (N_29151,N_18289,N_14673);
nand U29152 (N_29152,N_18443,N_12028);
and U29153 (N_29153,N_12970,N_14752);
nand U29154 (N_29154,N_15900,N_19707);
or U29155 (N_29155,N_10397,N_11184);
xor U29156 (N_29156,N_15347,N_10258);
nor U29157 (N_29157,N_10412,N_10727);
nand U29158 (N_29158,N_12464,N_16106);
nor U29159 (N_29159,N_16326,N_10712);
nand U29160 (N_29160,N_14858,N_10039);
and U29161 (N_29161,N_10681,N_12154);
nand U29162 (N_29162,N_12014,N_17270);
or U29163 (N_29163,N_17113,N_13666);
nand U29164 (N_29164,N_19153,N_16923);
or U29165 (N_29165,N_14540,N_16635);
nor U29166 (N_29166,N_13624,N_11309);
and U29167 (N_29167,N_17703,N_17170);
nor U29168 (N_29168,N_18459,N_17409);
nand U29169 (N_29169,N_11143,N_10929);
or U29170 (N_29170,N_18957,N_14135);
nor U29171 (N_29171,N_11685,N_19233);
nand U29172 (N_29172,N_14836,N_13340);
nor U29173 (N_29173,N_10337,N_15516);
xor U29174 (N_29174,N_10988,N_16855);
nor U29175 (N_29175,N_14464,N_10276);
or U29176 (N_29176,N_14028,N_12697);
nand U29177 (N_29177,N_12374,N_11182);
and U29178 (N_29178,N_18286,N_17276);
and U29179 (N_29179,N_14418,N_11563);
nor U29180 (N_29180,N_14734,N_12979);
and U29181 (N_29181,N_16460,N_19481);
or U29182 (N_29182,N_17825,N_15230);
and U29183 (N_29183,N_17265,N_16144);
or U29184 (N_29184,N_18710,N_13373);
nand U29185 (N_29185,N_13805,N_14687);
nor U29186 (N_29186,N_11565,N_11178);
nor U29187 (N_29187,N_13692,N_10754);
or U29188 (N_29188,N_16030,N_11267);
nor U29189 (N_29189,N_12982,N_14550);
nor U29190 (N_29190,N_13594,N_18123);
nor U29191 (N_29191,N_11318,N_17029);
or U29192 (N_29192,N_13080,N_10112);
or U29193 (N_29193,N_16678,N_14382);
or U29194 (N_29194,N_17772,N_13332);
or U29195 (N_29195,N_10496,N_18570);
and U29196 (N_29196,N_14039,N_10263);
and U29197 (N_29197,N_16107,N_16140);
nand U29198 (N_29198,N_16814,N_13981);
nand U29199 (N_29199,N_11277,N_11341);
or U29200 (N_29200,N_17419,N_19306);
nor U29201 (N_29201,N_15876,N_14778);
nor U29202 (N_29202,N_14583,N_11265);
xnor U29203 (N_29203,N_14601,N_17801);
nor U29204 (N_29204,N_10258,N_14269);
and U29205 (N_29205,N_19091,N_19111);
nand U29206 (N_29206,N_19130,N_13121);
nand U29207 (N_29207,N_18964,N_13701);
and U29208 (N_29208,N_17412,N_12308);
and U29209 (N_29209,N_12802,N_15079);
or U29210 (N_29210,N_14932,N_18946);
nor U29211 (N_29211,N_12766,N_10390);
nand U29212 (N_29212,N_13862,N_19176);
and U29213 (N_29213,N_11131,N_18896);
nor U29214 (N_29214,N_13226,N_16070);
or U29215 (N_29215,N_10592,N_10888);
nand U29216 (N_29216,N_15319,N_16027);
nand U29217 (N_29217,N_17823,N_17551);
or U29218 (N_29218,N_16979,N_17642);
nor U29219 (N_29219,N_19789,N_13727);
nand U29220 (N_29220,N_18988,N_17169);
and U29221 (N_29221,N_16662,N_18025);
and U29222 (N_29222,N_16214,N_18571);
nand U29223 (N_29223,N_10987,N_15365);
or U29224 (N_29224,N_10210,N_14033);
nor U29225 (N_29225,N_12328,N_16075);
nor U29226 (N_29226,N_10708,N_10315);
nand U29227 (N_29227,N_16860,N_16990);
or U29228 (N_29228,N_19300,N_10374);
nand U29229 (N_29229,N_17515,N_10844);
nor U29230 (N_29230,N_16958,N_17985);
or U29231 (N_29231,N_12499,N_13916);
and U29232 (N_29232,N_15175,N_17852);
nand U29233 (N_29233,N_14140,N_15263);
or U29234 (N_29234,N_15934,N_19948);
and U29235 (N_29235,N_16935,N_19867);
nor U29236 (N_29236,N_10492,N_10271);
and U29237 (N_29237,N_14889,N_16063);
nor U29238 (N_29238,N_17875,N_14078);
nor U29239 (N_29239,N_13571,N_19104);
nand U29240 (N_29240,N_19433,N_13302);
or U29241 (N_29241,N_19363,N_15223);
and U29242 (N_29242,N_16112,N_14100);
nor U29243 (N_29243,N_18688,N_15686);
or U29244 (N_29244,N_15795,N_15978);
xnor U29245 (N_29245,N_18272,N_13160);
and U29246 (N_29246,N_18768,N_14446);
nor U29247 (N_29247,N_18343,N_11702);
or U29248 (N_29248,N_19617,N_15271);
nor U29249 (N_29249,N_12042,N_15166);
nor U29250 (N_29250,N_12157,N_19908);
and U29251 (N_29251,N_19360,N_17997);
xnor U29252 (N_29252,N_17554,N_18020);
nand U29253 (N_29253,N_13515,N_17619);
nor U29254 (N_29254,N_18377,N_12255);
nor U29255 (N_29255,N_16680,N_12803);
or U29256 (N_29256,N_11982,N_12864);
or U29257 (N_29257,N_16276,N_16504);
nand U29258 (N_29258,N_13534,N_18014);
or U29259 (N_29259,N_13715,N_17226);
or U29260 (N_29260,N_12074,N_11413);
nand U29261 (N_29261,N_12928,N_13005);
xor U29262 (N_29262,N_19335,N_11846);
or U29263 (N_29263,N_15101,N_15074);
nor U29264 (N_29264,N_12827,N_19310);
nand U29265 (N_29265,N_13485,N_12030);
nor U29266 (N_29266,N_14951,N_10549);
or U29267 (N_29267,N_18291,N_19901);
nor U29268 (N_29268,N_19611,N_16767);
nor U29269 (N_29269,N_15620,N_18477);
nand U29270 (N_29270,N_12555,N_19869);
and U29271 (N_29271,N_12514,N_18938);
or U29272 (N_29272,N_13345,N_11265);
nand U29273 (N_29273,N_10620,N_15491);
and U29274 (N_29274,N_12429,N_10754);
and U29275 (N_29275,N_18734,N_14807);
nand U29276 (N_29276,N_16146,N_11137);
or U29277 (N_29277,N_18354,N_14000);
or U29278 (N_29278,N_19280,N_10405);
nand U29279 (N_29279,N_15394,N_17698);
nor U29280 (N_29280,N_10488,N_12088);
or U29281 (N_29281,N_13578,N_15896);
nor U29282 (N_29282,N_14541,N_16165);
nor U29283 (N_29283,N_15769,N_16224);
nand U29284 (N_29284,N_18930,N_11559);
nor U29285 (N_29285,N_15001,N_17075);
or U29286 (N_29286,N_12189,N_15736);
nand U29287 (N_29287,N_14094,N_16437);
and U29288 (N_29288,N_10332,N_12492);
nand U29289 (N_29289,N_12893,N_19202);
and U29290 (N_29290,N_15792,N_13133);
nor U29291 (N_29291,N_16530,N_10725);
and U29292 (N_29292,N_13444,N_11504);
nor U29293 (N_29293,N_10221,N_18328);
or U29294 (N_29294,N_15239,N_10844);
nand U29295 (N_29295,N_19434,N_17463);
or U29296 (N_29296,N_18138,N_13230);
nand U29297 (N_29297,N_10788,N_10930);
or U29298 (N_29298,N_14844,N_14508);
nand U29299 (N_29299,N_13733,N_12818);
nand U29300 (N_29300,N_16265,N_17932);
nor U29301 (N_29301,N_17596,N_18238);
nand U29302 (N_29302,N_18268,N_14825);
nor U29303 (N_29303,N_11525,N_14250);
or U29304 (N_29304,N_12072,N_13921);
nand U29305 (N_29305,N_19937,N_18678);
and U29306 (N_29306,N_19428,N_19436);
and U29307 (N_29307,N_16824,N_13897);
or U29308 (N_29308,N_18030,N_13353);
or U29309 (N_29309,N_15641,N_11931);
nor U29310 (N_29310,N_10931,N_17597);
nor U29311 (N_29311,N_11472,N_19320);
nand U29312 (N_29312,N_12848,N_16216);
nand U29313 (N_29313,N_18782,N_13837);
nor U29314 (N_29314,N_13332,N_12226);
or U29315 (N_29315,N_15339,N_16582);
or U29316 (N_29316,N_10710,N_14595);
nor U29317 (N_29317,N_13843,N_14704);
or U29318 (N_29318,N_18808,N_13158);
xor U29319 (N_29319,N_15507,N_13198);
or U29320 (N_29320,N_11216,N_13462);
nand U29321 (N_29321,N_14133,N_16663);
nand U29322 (N_29322,N_12993,N_13575);
nor U29323 (N_29323,N_15294,N_13337);
or U29324 (N_29324,N_11860,N_16264);
nand U29325 (N_29325,N_16862,N_19294);
nand U29326 (N_29326,N_16173,N_12678);
nor U29327 (N_29327,N_18595,N_14775);
and U29328 (N_29328,N_16679,N_17051);
and U29329 (N_29329,N_11086,N_16262);
and U29330 (N_29330,N_12734,N_19803);
nor U29331 (N_29331,N_14512,N_19387);
and U29332 (N_29332,N_13698,N_15739);
nor U29333 (N_29333,N_19262,N_15909);
or U29334 (N_29334,N_10759,N_18781);
nor U29335 (N_29335,N_10043,N_15661);
nor U29336 (N_29336,N_17095,N_15954);
and U29337 (N_29337,N_12535,N_13360);
nand U29338 (N_29338,N_19118,N_13530);
or U29339 (N_29339,N_13647,N_19155);
and U29340 (N_29340,N_16732,N_17973);
or U29341 (N_29341,N_10437,N_12015);
nor U29342 (N_29342,N_18672,N_14843);
and U29343 (N_29343,N_17390,N_11622);
or U29344 (N_29344,N_17271,N_14781);
nand U29345 (N_29345,N_13337,N_10723);
nor U29346 (N_29346,N_12953,N_18866);
nand U29347 (N_29347,N_11293,N_19389);
nand U29348 (N_29348,N_17220,N_14616);
nor U29349 (N_29349,N_12648,N_11840);
nor U29350 (N_29350,N_13442,N_15768);
nand U29351 (N_29351,N_19694,N_10533);
nor U29352 (N_29352,N_17991,N_11854);
nand U29353 (N_29353,N_13915,N_14248);
nand U29354 (N_29354,N_12408,N_14470);
nand U29355 (N_29355,N_19788,N_15208);
and U29356 (N_29356,N_19881,N_10637);
or U29357 (N_29357,N_10369,N_10263);
or U29358 (N_29358,N_16757,N_19340);
nor U29359 (N_29359,N_11368,N_14957);
and U29360 (N_29360,N_14965,N_19194);
nor U29361 (N_29361,N_16191,N_10134);
or U29362 (N_29362,N_10876,N_16783);
and U29363 (N_29363,N_13476,N_10341);
and U29364 (N_29364,N_14542,N_16695);
or U29365 (N_29365,N_12301,N_19855);
or U29366 (N_29366,N_10558,N_19297);
nor U29367 (N_29367,N_18650,N_10067);
nor U29368 (N_29368,N_15462,N_15819);
or U29369 (N_29369,N_14282,N_17523);
nor U29370 (N_29370,N_19891,N_13534);
nor U29371 (N_29371,N_11354,N_18156);
nor U29372 (N_29372,N_11604,N_10286);
and U29373 (N_29373,N_13774,N_10173);
nor U29374 (N_29374,N_14479,N_13079);
nand U29375 (N_29375,N_14582,N_19660);
or U29376 (N_29376,N_14446,N_14048);
and U29377 (N_29377,N_14722,N_14472);
nor U29378 (N_29378,N_18011,N_11430);
and U29379 (N_29379,N_15875,N_11517);
nor U29380 (N_29380,N_12746,N_19390);
or U29381 (N_29381,N_17481,N_15809);
and U29382 (N_29382,N_12594,N_11412);
nand U29383 (N_29383,N_13103,N_10899);
nor U29384 (N_29384,N_18797,N_17763);
xor U29385 (N_29385,N_16957,N_17779);
or U29386 (N_29386,N_17526,N_14643);
and U29387 (N_29387,N_10117,N_18635);
nand U29388 (N_29388,N_16600,N_12899);
nor U29389 (N_29389,N_17165,N_17785);
xor U29390 (N_29390,N_15585,N_12958);
or U29391 (N_29391,N_13370,N_16020);
and U29392 (N_29392,N_13003,N_13067);
and U29393 (N_29393,N_10138,N_10899);
nor U29394 (N_29394,N_19527,N_17611);
nand U29395 (N_29395,N_15318,N_19644);
nor U29396 (N_29396,N_11300,N_11699);
nand U29397 (N_29397,N_17566,N_19691);
or U29398 (N_29398,N_19778,N_17133);
nor U29399 (N_29399,N_10689,N_13608);
nand U29400 (N_29400,N_18696,N_16943);
nand U29401 (N_29401,N_16331,N_11671);
nor U29402 (N_29402,N_15816,N_12304);
or U29403 (N_29403,N_12375,N_19350);
nand U29404 (N_29404,N_15250,N_16515);
nor U29405 (N_29405,N_19508,N_11423);
and U29406 (N_29406,N_14226,N_15413);
or U29407 (N_29407,N_17216,N_13010);
and U29408 (N_29408,N_19193,N_10294);
nand U29409 (N_29409,N_18948,N_11363);
nand U29410 (N_29410,N_17593,N_16716);
nor U29411 (N_29411,N_14735,N_13793);
nor U29412 (N_29412,N_14708,N_11131);
nor U29413 (N_29413,N_12064,N_16510);
nand U29414 (N_29414,N_11533,N_13452);
and U29415 (N_29415,N_14610,N_19298);
or U29416 (N_29416,N_15413,N_13565);
or U29417 (N_29417,N_14298,N_12231);
or U29418 (N_29418,N_16842,N_18937);
nor U29419 (N_29419,N_13800,N_17477);
and U29420 (N_29420,N_13012,N_10877);
or U29421 (N_29421,N_12638,N_15829);
nand U29422 (N_29422,N_18200,N_18457);
nor U29423 (N_29423,N_16508,N_14441);
nor U29424 (N_29424,N_10022,N_19028);
nor U29425 (N_29425,N_17099,N_16179);
nand U29426 (N_29426,N_12507,N_18189);
nand U29427 (N_29427,N_13593,N_19491);
and U29428 (N_29428,N_18496,N_12507);
and U29429 (N_29429,N_12556,N_12889);
nor U29430 (N_29430,N_12822,N_15536);
nor U29431 (N_29431,N_12651,N_11565);
nand U29432 (N_29432,N_18657,N_10749);
nand U29433 (N_29433,N_11299,N_11932);
nand U29434 (N_29434,N_19440,N_18060);
nand U29435 (N_29435,N_15995,N_14481);
or U29436 (N_29436,N_11509,N_19969);
and U29437 (N_29437,N_13222,N_17509);
and U29438 (N_29438,N_17305,N_12699);
and U29439 (N_29439,N_10044,N_15463);
and U29440 (N_29440,N_10350,N_11255);
nor U29441 (N_29441,N_14772,N_16269);
nor U29442 (N_29442,N_19864,N_19623);
nand U29443 (N_29443,N_14373,N_16899);
or U29444 (N_29444,N_19366,N_17252);
nor U29445 (N_29445,N_16125,N_14596);
and U29446 (N_29446,N_11011,N_10708);
nand U29447 (N_29447,N_18757,N_17063);
nor U29448 (N_29448,N_15043,N_12700);
nand U29449 (N_29449,N_14302,N_10091);
or U29450 (N_29450,N_17470,N_13270);
xnor U29451 (N_29451,N_10068,N_11369);
nor U29452 (N_29452,N_17148,N_13310);
nand U29453 (N_29453,N_14123,N_13339);
nor U29454 (N_29454,N_18305,N_14688);
nor U29455 (N_29455,N_10433,N_13436);
nor U29456 (N_29456,N_14473,N_15247);
and U29457 (N_29457,N_15660,N_17285);
or U29458 (N_29458,N_11807,N_12245);
nor U29459 (N_29459,N_16230,N_11383);
and U29460 (N_29460,N_18223,N_12109);
and U29461 (N_29461,N_17507,N_19436);
and U29462 (N_29462,N_11890,N_19886);
nand U29463 (N_29463,N_16413,N_17236);
and U29464 (N_29464,N_14511,N_12522);
nor U29465 (N_29465,N_11683,N_16605);
or U29466 (N_29466,N_10129,N_16837);
and U29467 (N_29467,N_16149,N_16216);
and U29468 (N_29468,N_19185,N_14890);
and U29469 (N_29469,N_16560,N_14480);
or U29470 (N_29470,N_10649,N_14785);
nand U29471 (N_29471,N_14051,N_15377);
xnor U29472 (N_29472,N_14891,N_12460);
nor U29473 (N_29473,N_18710,N_15151);
nor U29474 (N_29474,N_14152,N_16363);
nand U29475 (N_29475,N_14035,N_18940);
nand U29476 (N_29476,N_15152,N_19529);
nand U29477 (N_29477,N_15935,N_10030);
and U29478 (N_29478,N_15020,N_17872);
and U29479 (N_29479,N_17220,N_14849);
nor U29480 (N_29480,N_10350,N_19493);
and U29481 (N_29481,N_16322,N_16467);
nand U29482 (N_29482,N_17037,N_18526);
or U29483 (N_29483,N_18479,N_10358);
or U29484 (N_29484,N_13136,N_15792);
nor U29485 (N_29485,N_15884,N_13094);
xnor U29486 (N_29486,N_14290,N_10701);
and U29487 (N_29487,N_13606,N_18355);
and U29488 (N_29488,N_11993,N_11674);
nor U29489 (N_29489,N_10694,N_17107);
nor U29490 (N_29490,N_16046,N_10471);
nor U29491 (N_29491,N_18366,N_19540);
and U29492 (N_29492,N_12990,N_10906);
and U29493 (N_29493,N_16120,N_19947);
nand U29494 (N_29494,N_16476,N_16708);
and U29495 (N_29495,N_18988,N_14590);
nand U29496 (N_29496,N_10128,N_15978);
nor U29497 (N_29497,N_18076,N_13224);
and U29498 (N_29498,N_17196,N_11641);
or U29499 (N_29499,N_10166,N_17194);
nand U29500 (N_29500,N_14054,N_13800);
nor U29501 (N_29501,N_11270,N_13902);
nor U29502 (N_29502,N_12878,N_13437);
nor U29503 (N_29503,N_14071,N_18420);
and U29504 (N_29504,N_10886,N_13856);
nor U29505 (N_29505,N_14614,N_19392);
and U29506 (N_29506,N_16317,N_18999);
or U29507 (N_29507,N_18268,N_13949);
and U29508 (N_29508,N_17185,N_14850);
nand U29509 (N_29509,N_15424,N_10654);
or U29510 (N_29510,N_13428,N_16775);
nand U29511 (N_29511,N_14342,N_17941);
or U29512 (N_29512,N_16409,N_17666);
or U29513 (N_29513,N_16343,N_15641);
or U29514 (N_29514,N_15212,N_12205);
or U29515 (N_29515,N_18503,N_11619);
nor U29516 (N_29516,N_12621,N_10609);
nor U29517 (N_29517,N_12286,N_12994);
nand U29518 (N_29518,N_19029,N_18143);
and U29519 (N_29519,N_18170,N_18502);
or U29520 (N_29520,N_19602,N_14576);
nand U29521 (N_29521,N_14905,N_14948);
and U29522 (N_29522,N_17222,N_15033);
nor U29523 (N_29523,N_15733,N_16690);
nand U29524 (N_29524,N_16981,N_11238);
nor U29525 (N_29525,N_17982,N_10068);
nor U29526 (N_29526,N_12836,N_15936);
and U29527 (N_29527,N_13790,N_12161);
nor U29528 (N_29528,N_14962,N_11712);
and U29529 (N_29529,N_14792,N_17221);
nor U29530 (N_29530,N_19225,N_11023);
nand U29531 (N_29531,N_12606,N_10216);
or U29532 (N_29532,N_13448,N_19627);
nor U29533 (N_29533,N_10430,N_11888);
nor U29534 (N_29534,N_19511,N_11790);
nor U29535 (N_29535,N_14785,N_11515);
nand U29536 (N_29536,N_17347,N_10083);
nand U29537 (N_29537,N_12782,N_10668);
nor U29538 (N_29538,N_11330,N_15422);
and U29539 (N_29539,N_11158,N_12531);
and U29540 (N_29540,N_16431,N_11483);
nand U29541 (N_29541,N_11865,N_16228);
nand U29542 (N_29542,N_13449,N_17932);
or U29543 (N_29543,N_18122,N_12688);
and U29544 (N_29544,N_19644,N_10672);
and U29545 (N_29545,N_16585,N_16740);
or U29546 (N_29546,N_15073,N_18663);
nor U29547 (N_29547,N_14547,N_16015);
nand U29548 (N_29548,N_12700,N_14707);
nand U29549 (N_29549,N_18549,N_17366);
or U29550 (N_29550,N_10759,N_10098);
nand U29551 (N_29551,N_16299,N_17617);
nor U29552 (N_29552,N_19157,N_12286);
nor U29553 (N_29553,N_17963,N_12614);
nand U29554 (N_29554,N_10857,N_12025);
nor U29555 (N_29555,N_16072,N_16764);
nor U29556 (N_29556,N_10013,N_14009);
and U29557 (N_29557,N_15485,N_19124);
nor U29558 (N_29558,N_11876,N_12083);
or U29559 (N_29559,N_14815,N_13188);
nand U29560 (N_29560,N_15876,N_12476);
nand U29561 (N_29561,N_14815,N_15785);
nand U29562 (N_29562,N_11125,N_16948);
nand U29563 (N_29563,N_18468,N_11220);
and U29564 (N_29564,N_11130,N_10014);
or U29565 (N_29565,N_14139,N_11364);
nand U29566 (N_29566,N_10579,N_18791);
nor U29567 (N_29567,N_14248,N_13434);
nand U29568 (N_29568,N_12344,N_15853);
or U29569 (N_29569,N_14100,N_19764);
and U29570 (N_29570,N_10547,N_16215);
and U29571 (N_29571,N_10092,N_15729);
nor U29572 (N_29572,N_16385,N_11239);
and U29573 (N_29573,N_13818,N_19137);
and U29574 (N_29574,N_16047,N_12172);
or U29575 (N_29575,N_14200,N_12632);
and U29576 (N_29576,N_10663,N_10789);
and U29577 (N_29577,N_13415,N_15049);
or U29578 (N_29578,N_16833,N_17686);
nand U29579 (N_29579,N_11320,N_13243);
or U29580 (N_29580,N_17554,N_15043);
or U29581 (N_29581,N_11704,N_19782);
or U29582 (N_29582,N_14839,N_17329);
or U29583 (N_29583,N_11103,N_12194);
and U29584 (N_29584,N_17607,N_17019);
and U29585 (N_29585,N_12896,N_15568);
nor U29586 (N_29586,N_16504,N_10954);
nand U29587 (N_29587,N_14422,N_18570);
nand U29588 (N_29588,N_13030,N_18255);
nor U29589 (N_29589,N_14060,N_15977);
nand U29590 (N_29590,N_18061,N_14264);
and U29591 (N_29591,N_13582,N_17820);
nor U29592 (N_29592,N_12216,N_18258);
or U29593 (N_29593,N_15887,N_14480);
nand U29594 (N_29594,N_18641,N_14868);
or U29595 (N_29595,N_12602,N_11501);
nand U29596 (N_29596,N_11965,N_16816);
nand U29597 (N_29597,N_16575,N_14530);
nand U29598 (N_29598,N_11087,N_11492);
xor U29599 (N_29599,N_13111,N_11835);
and U29600 (N_29600,N_18118,N_14429);
nand U29601 (N_29601,N_18259,N_14649);
nor U29602 (N_29602,N_15492,N_15849);
or U29603 (N_29603,N_11734,N_14249);
and U29604 (N_29604,N_14341,N_19586);
or U29605 (N_29605,N_19378,N_10717);
nor U29606 (N_29606,N_18388,N_17581);
or U29607 (N_29607,N_12196,N_10870);
nand U29608 (N_29608,N_16826,N_12792);
xnor U29609 (N_29609,N_16436,N_10755);
and U29610 (N_29610,N_18970,N_19403);
and U29611 (N_29611,N_11771,N_19889);
or U29612 (N_29612,N_16177,N_13858);
nand U29613 (N_29613,N_10030,N_15945);
and U29614 (N_29614,N_13163,N_16231);
and U29615 (N_29615,N_13181,N_14128);
nor U29616 (N_29616,N_16054,N_18082);
and U29617 (N_29617,N_19256,N_18969);
nor U29618 (N_29618,N_16663,N_17128);
and U29619 (N_29619,N_11256,N_18716);
nand U29620 (N_29620,N_18184,N_10913);
nor U29621 (N_29621,N_12396,N_10620);
and U29622 (N_29622,N_15524,N_14108);
nor U29623 (N_29623,N_10549,N_11940);
nor U29624 (N_29624,N_15307,N_17629);
or U29625 (N_29625,N_19113,N_10445);
and U29626 (N_29626,N_17236,N_12507);
nand U29627 (N_29627,N_16884,N_14502);
or U29628 (N_29628,N_11435,N_16679);
nor U29629 (N_29629,N_16838,N_18302);
nor U29630 (N_29630,N_17560,N_16267);
nand U29631 (N_29631,N_13997,N_14548);
and U29632 (N_29632,N_10967,N_15154);
nor U29633 (N_29633,N_12651,N_10938);
and U29634 (N_29634,N_12314,N_18853);
nor U29635 (N_29635,N_18196,N_18303);
xnor U29636 (N_29636,N_13923,N_16922);
or U29637 (N_29637,N_18175,N_19021);
nand U29638 (N_29638,N_13760,N_12155);
or U29639 (N_29639,N_15422,N_11904);
and U29640 (N_29640,N_14400,N_13489);
nor U29641 (N_29641,N_18379,N_17187);
or U29642 (N_29642,N_16956,N_16954);
or U29643 (N_29643,N_15768,N_12237);
and U29644 (N_29644,N_10354,N_12328);
or U29645 (N_29645,N_13371,N_15799);
nand U29646 (N_29646,N_13849,N_18000);
and U29647 (N_29647,N_12930,N_12439);
nor U29648 (N_29648,N_17991,N_17447);
nand U29649 (N_29649,N_17588,N_15628);
nor U29650 (N_29650,N_16520,N_10217);
or U29651 (N_29651,N_12962,N_17908);
nand U29652 (N_29652,N_13744,N_17438);
and U29653 (N_29653,N_15704,N_13272);
nor U29654 (N_29654,N_18390,N_15919);
and U29655 (N_29655,N_18708,N_18015);
nor U29656 (N_29656,N_11001,N_16103);
nand U29657 (N_29657,N_13663,N_19867);
nor U29658 (N_29658,N_18418,N_14845);
and U29659 (N_29659,N_16063,N_13326);
and U29660 (N_29660,N_16122,N_17618);
nor U29661 (N_29661,N_13279,N_15739);
nor U29662 (N_29662,N_15629,N_12279);
or U29663 (N_29663,N_19221,N_11823);
nand U29664 (N_29664,N_13158,N_16981);
nand U29665 (N_29665,N_11700,N_12120);
or U29666 (N_29666,N_16529,N_17103);
nor U29667 (N_29667,N_17981,N_15483);
and U29668 (N_29668,N_16674,N_18760);
or U29669 (N_29669,N_12438,N_15909);
nor U29670 (N_29670,N_18215,N_15827);
nand U29671 (N_29671,N_15964,N_15493);
nand U29672 (N_29672,N_18224,N_18014);
and U29673 (N_29673,N_14744,N_12041);
or U29674 (N_29674,N_12494,N_15958);
or U29675 (N_29675,N_19543,N_11086);
nand U29676 (N_29676,N_15022,N_10330);
nor U29677 (N_29677,N_12358,N_16550);
nand U29678 (N_29678,N_14822,N_13579);
or U29679 (N_29679,N_13302,N_19682);
nor U29680 (N_29680,N_19827,N_17544);
nand U29681 (N_29681,N_17008,N_13189);
nor U29682 (N_29682,N_15446,N_11492);
nor U29683 (N_29683,N_16364,N_14330);
or U29684 (N_29684,N_12899,N_10107);
and U29685 (N_29685,N_17173,N_10817);
nor U29686 (N_29686,N_15737,N_14781);
nor U29687 (N_29687,N_15378,N_13592);
nor U29688 (N_29688,N_18190,N_11403);
nand U29689 (N_29689,N_15352,N_12325);
or U29690 (N_29690,N_12967,N_19057);
nand U29691 (N_29691,N_10159,N_15145);
nor U29692 (N_29692,N_16808,N_11310);
and U29693 (N_29693,N_14339,N_16224);
nor U29694 (N_29694,N_14330,N_12427);
nor U29695 (N_29695,N_17452,N_11741);
or U29696 (N_29696,N_14747,N_13058);
and U29697 (N_29697,N_15287,N_11204);
nand U29698 (N_29698,N_13984,N_15081);
nor U29699 (N_29699,N_19782,N_17660);
nor U29700 (N_29700,N_19649,N_18616);
or U29701 (N_29701,N_19762,N_16853);
nand U29702 (N_29702,N_17011,N_19584);
and U29703 (N_29703,N_15735,N_13308);
nand U29704 (N_29704,N_10441,N_15782);
nand U29705 (N_29705,N_16071,N_15253);
and U29706 (N_29706,N_13873,N_14102);
and U29707 (N_29707,N_15428,N_10229);
or U29708 (N_29708,N_13558,N_17620);
and U29709 (N_29709,N_17967,N_14578);
or U29710 (N_29710,N_10431,N_19931);
and U29711 (N_29711,N_16803,N_10349);
nand U29712 (N_29712,N_17957,N_12835);
or U29713 (N_29713,N_13767,N_10889);
nor U29714 (N_29714,N_16542,N_18376);
and U29715 (N_29715,N_19731,N_17358);
nor U29716 (N_29716,N_16775,N_19831);
nor U29717 (N_29717,N_11305,N_10758);
and U29718 (N_29718,N_13451,N_12018);
and U29719 (N_29719,N_10178,N_15899);
or U29720 (N_29720,N_14077,N_16462);
nor U29721 (N_29721,N_14460,N_19931);
xor U29722 (N_29722,N_11024,N_16884);
nand U29723 (N_29723,N_10768,N_13938);
nand U29724 (N_29724,N_15824,N_11311);
and U29725 (N_29725,N_17406,N_17739);
nor U29726 (N_29726,N_11929,N_15676);
and U29727 (N_29727,N_12892,N_13167);
or U29728 (N_29728,N_13008,N_12356);
nand U29729 (N_29729,N_18665,N_19417);
or U29730 (N_29730,N_16886,N_16758);
nor U29731 (N_29731,N_15580,N_16771);
or U29732 (N_29732,N_16026,N_15458);
xnor U29733 (N_29733,N_13840,N_11485);
nand U29734 (N_29734,N_18794,N_13349);
and U29735 (N_29735,N_19116,N_13706);
nand U29736 (N_29736,N_11732,N_15499);
or U29737 (N_29737,N_12469,N_19581);
or U29738 (N_29738,N_13409,N_10574);
nand U29739 (N_29739,N_10738,N_16537);
nand U29740 (N_29740,N_14523,N_12504);
nand U29741 (N_29741,N_13224,N_10588);
and U29742 (N_29742,N_14733,N_19438);
nor U29743 (N_29743,N_11555,N_13838);
and U29744 (N_29744,N_11236,N_17634);
nor U29745 (N_29745,N_11099,N_19084);
nor U29746 (N_29746,N_16555,N_15122);
or U29747 (N_29747,N_15924,N_12353);
xor U29748 (N_29748,N_13034,N_19667);
and U29749 (N_29749,N_17888,N_11196);
xor U29750 (N_29750,N_18866,N_19715);
and U29751 (N_29751,N_17223,N_19595);
and U29752 (N_29752,N_14421,N_13201);
and U29753 (N_29753,N_13962,N_11842);
nor U29754 (N_29754,N_11728,N_16547);
or U29755 (N_29755,N_18494,N_11975);
nor U29756 (N_29756,N_18698,N_15580);
or U29757 (N_29757,N_14198,N_13999);
nand U29758 (N_29758,N_19769,N_17422);
nor U29759 (N_29759,N_15757,N_18460);
or U29760 (N_29760,N_18493,N_13947);
and U29761 (N_29761,N_19733,N_16302);
or U29762 (N_29762,N_15257,N_14315);
xor U29763 (N_29763,N_12351,N_19407);
or U29764 (N_29764,N_14519,N_12658);
nor U29765 (N_29765,N_10192,N_12460);
nor U29766 (N_29766,N_15617,N_10330);
nand U29767 (N_29767,N_12967,N_13870);
or U29768 (N_29768,N_16900,N_15223);
or U29769 (N_29769,N_13293,N_18495);
nor U29770 (N_29770,N_19745,N_10943);
or U29771 (N_29771,N_16391,N_16325);
nor U29772 (N_29772,N_12470,N_19808);
nor U29773 (N_29773,N_16098,N_18836);
nand U29774 (N_29774,N_11226,N_11460);
or U29775 (N_29775,N_11956,N_11529);
and U29776 (N_29776,N_14125,N_18230);
nand U29777 (N_29777,N_15739,N_12703);
or U29778 (N_29778,N_12268,N_10061);
nor U29779 (N_29779,N_15088,N_11531);
nand U29780 (N_29780,N_12221,N_10004);
nand U29781 (N_29781,N_17153,N_17107);
and U29782 (N_29782,N_11542,N_19832);
or U29783 (N_29783,N_16374,N_12184);
and U29784 (N_29784,N_12946,N_14199);
nand U29785 (N_29785,N_15282,N_11408);
or U29786 (N_29786,N_13317,N_14157);
and U29787 (N_29787,N_12437,N_11340);
and U29788 (N_29788,N_14857,N_15563);
nand U29789 (N_29789,N_16010,N_14328);
or U29790 (N_29790,N_15826,N_14683);
and U29791 (N_29791,N_18122,N_10559);
nor U29792 (N_29792,N_19487,N_13559);
nor U29793 (N_29793,N_19712,N_13354);
and U29794 (N_29794,N_18135,N_14684);
nor U29795 (N_29795,N_10264,N_10848);
and U29796 (N_29796,N_14040,N_17844);
and U29797 (N_29797,N_11809,N_12698);
nor U29798 (N_29798,N_12884,N_11279);
and U29799 (N_29799,N_17425,N_11999);
nor U29800 (N_29800,N_18124,N_12604);
nor U29801 (N_29801,N_19171,N_17483);
or U29802 (N_29802,N_12191,N_15663);
and U29803 (N_29803,N_14765,N_13626);
nand U29804 (N_29804,N_18371,N_16946);
nor U29805 (N_29805,N_18267,N_13036);
nand U29806 (N_29806,N_17974,N_12436);
nand U29807 (N_29807,N_13122,N_12511);
nor U29808 (N_29808,N_10722,N_14835);
nand U29809 (N_29809,N_16411,N_16752);
nor U29810 (N_29810,N_11770,N_14573);
or U29811 (N_29811,N_19060,N_13550);
nor U29812 (N_29812,N_19443,N_10920);
nand U29813 (N_29813,N_10487,N_16374);
nand U29814 (N_29814,N_18254,N_10143);
or U29815 (N_29815,N_19129,N_14180);
and U29816 (N_29816,N_12273,N_11319);
nand U29817 (N_29817,N_18543,N_19067);
and U29818 (N_29818,N_18973,N_10738);
nor U29819 (N_29819,N_14386,N_19893);
or U29820 (N_29820,N_15855,N_16571);
nor U29821 (N_29821,N_11527,N_15423);
xnor U29822 (N_29822,N_11653,N_19633);
nand U29823 (N_29823,N_17847,N_19468);
nor U29824 (N_29824,N_19487,N_11965);
nor U29825 (N_29825,N_11895,N_13100);
nand U29826 (N_29826,N_15126,N_10358);
nand U29827 (N_29827,N_10082,N_18668);
nor U29828 (N_29828,N_11712,N_15269);
nor U29829 (N_29829,N_10269,N_19884);
nor U29830 (N_29830,N_16289,N_12195);
nor U29831 (N_29831,N_12090,N_16710);
and U29832 (N_29832,N_10988,N_12009);
nor U29833 (N_29833,N_10425,N_18558);
or U29834 (N_29834,N_10683,N_16508);
nand U29835 (N_29835,N_12871,N_11497);
nor U29836 (N_29836,N_18551,N_14773);
nand U29837 (N_29837,N_19738,N_16148);
or U29838 (N_29838,N_19055,N_18894);
or U29839 (N_29839,N_18894,N_16511);
or U29840 (N_29840,N_19458,N_15336);
nor U29841 (N_29841,N_15974,N_15398);
and U29842 (N_29842,N_11576,N_14930);
and U29843 (N_29843,N_19047,N_13244);
and U29844 (N_29844,N_16925,N_15211);
nor U29845 (N_29845,N_18053,N_14198);
nand U29846 (N_29846,N_16415,N_12765);
and U29847 (N_29847,N_11262,N_17733);
nor U29848 (N_29848,N_14903,N_19159);
and U29849 (N_29849,N_10809,N_17060);
and U29850 (N_29850,N_15087,N_19950);
nor U29851 (N_29851,N_15855,N_19698);
nor U29852 (N_29852,N_18590,N_17482);
nor U29853 (N_29853,N_15534,N_15588);
and U29854 (N_29854,N_14577,N_12277);
nor U29855 (N_29855,N_17621,N_12223);
and U29856 (N_29856,N_14206,N_10805);
nand U29857 (N_29857,N_12016,N_11903);
and U29858 (N_29858,N_19232,N_10375);
nor U29859 (N_29859,N_18079,N_17891);
nor U29860 (N_29860,N_17382,N_13327);
and U29861 (N_29861,N_14018,N_18757);
and U29862 (N_29862,N_11322,N_13028);
or U29863 (N_29863,N_12462,N_11756);
nand U29864 (N_29864,N_12487,N_19618);
and U29865 (N_29865,N_16228,N_11763);
or U29866 (N_29866,N_16096,N_15216);
nor U29867 (N_29867,N_17808,N_17172);
nand U29868 (N_29868,N_12519,N_17111);
and U29869 (N_29869,N_13652,N_10500);
nand U29870 (N_29870,N_15878,N_13023);
nor U29871 (N_29871,N_10898,N_19609);
and U29872 (N_29872,N_16868,N_15081);
and U29873 (N_29873,N_19871,N_12861);
nor U29874 (N_29874,N_11061,N_17545);
and U29875 (N_29875,N_19731,N_13313);
or U29876 (N_29876,N_10265,N_12247);
nand U29877 (N_29877,N_10021,N_12428);
or U29878 (N_29878,N_15889,N_10237);
nand U29879 (N_29879,N_12396,N_11892);
nand U29880 (N_29880,N_14090,N_16784);
nor U29881 (N_29881,N_18670,N_18680);
nand U29882 (N_29882,N_14233,N_18846);
or U29883 (N_29883,N_10063,N_16962);
nand U29884 (N_29884,N_11026,N_15079);
and U29885 (N_29885,N_10067,N_13689);
nand U29886 (N_29886,N_11089,N_19159);
nor U29887 (N_29887,N_18688,N_18172);
and U29888 (N_29888,N_11977,N_14122);
nand U29889 (N_29889,N_10083,N_18954);
and U29890 (N_29890,N_12970,N_19844);
and U29891 (N_29891,N_13221,N_15659);
or U29892 (N_29892,N_16026,N_14976);
or U29893 (N_29893,N_10674,N_12810);
nand U29894 (N_29894,N_17648,N_12649);
and U29895 (N_29895,N_10651,N_14040);
xnor U29896 (N_29896,N_19685,N_19528);
nor U29897 (N_29897,N_15491,N_17968);
or U29898 (N_29898,N_15185,N_13583);
and U29899 (N_29899,N_15852,N_10664);
nand U29900 (N_29900,N_19850,N_13680);
nand U29901 (N_29901,N_10316,N_14828);
and U29902 (N_29902,N_16570,N_18597);
or U29903 (N_29903,N_10563,N_17456);
nand U29904 (N_29904,N_17995,N_17263);
or U29905 (N_29905,N_15301,N_15601);
nor U29906 (N_29906,N_11608,N_10683);
nor U29907 (N_29907,N_16000,N_15707);
nand U29908 (N_29908,N_12136,N_11729);
nand U29909 (N_29909,N_13179,N_16144);
nand U29910 (N_29910,N_19091,N_12859);
and U29911 (N_29911,N_11087,N_13505);
nand U29912 (N_29912,N_12697,N_11816);
or U29913 (N_29913,N_14512,N_16570);
or U29914 (N_29914,N_16677,N_17202);
nand U29915 (N_29915,N_13881,N_16440);
and U29916 (N_29916,N_14163,N_10222);
and U29917 (N_29917,N_11786,N_13951);
and U29918 (N_29918,N_19587,N_13720);
and U29919 (N_29919,N_10575,N_11184);
nor U29920 (N_29920,N_16148,N_14358);
nor U29921 (N_29921,N_10773,N_11276);
or U29922 (N_29922,N_16250,N_15292);
nor U29923 (N_29923,N_16636,N_19459);
and U29924 (N_29924,N_19285,N_13358);
nand U29925 (N_29925,N_13149,N_14581);
nand U29926 (N_29926,N_14887,N_16819);
nor U29927 (N_29927,N_15314,N_13083);
nor U29928 (N_29928,N_15019,N_12243);
nand U29929 (N_29929,N_19812,N_14132);
nor U29930 (N_29930,N_13788,N_16055);
nor U29931 (N_29931,N_15250,N_14122);
nor U29932 (N_29932,N_16437,N_18196);
nand U29933 (N_29933,N_11588,N_18514);
and U29934 (N_29934,N_13688,N_15332);
and U29935 (N_29935,N_15751,N_18780);
nand U29936 (N_29936,N_18078,N_13113);
nand U29937 (N_29937,N_12346,N_13791);
or U29938 (N_29938,N_18738,N_15538);
nand U29939 (N_29939,N_19806,N_11266);
or U29940 (N_29940,N_10000,N_14724);
or U29941 (N_29941,N_17260,N_18277);
xnor U29942 (N_29942,N_16138,N_19230);
nor U29943 (N_29943,N_19700,N_13277);
or U29944 (N_29944,N_13237,N_13966);
nand U29945 (N_29945,N_10726,N_15255);
nand U29946 (N_29946,N_10459,N_19229);
xnor U29947 (N_29947,N_10763,N_17923);
and U29948 (N_29948,N_16290,N_18683);
or U29949 (N_29949,N_19664,N_19502);
nand U29950 (N_29950,N_17902,N_18746);
nor U29951 (N_29951,N_15048,N_12031);
or U29952 (N_29952,N_11167,N_16709);
nor U29953 (N_29953,N_15956,N_18526);
nand U29954 (N_29954,N_16115,N_13424);
nand U29955 (N_29955,N_18948,N_13298);
nand U29956 (N_29956,N_19210,N_17557);
nor U29957 (N_29957,N_11229,N_17138);
and U29958 (N_29958,N_18602,N_12186);
nor U29959 (N_29959,N_10208,N_12162);
nand U29960 (N_29960,N_19741,N_18246);
nor U29961 (N_29961,N_18736,N_14149);
and U29962 (N_29962,N_12190,N_17451);
or U29963 (N_29963,N_11642,N_15566);
and U29964 (N_29964,N_10489,N_15704);
or U29965 (N_29965,N_19563,N_14268);
or U29966 (N_29966,N_14142,N_15499);
or U29967 (N_29967,N_17651,N_17660);
nand U29968 (N_29968,N_14140,N_17162);
and U29969 (N_29969,N_10340,N_11638);
and U29970 (N_29970,N_11177,N_11807);
and U29971 (N_29971,N_10637,N_18854);
nor U29972 (N_29972,N_14736,N_15636);
nand U29973 (N_29973,N_13468,N_15112);
and U29974 (N_29974,N_19717,N_15818);
xor U29975 (N_29975,N_19260,N_17397);
and U29976 (N_29976,N_15946,N_10516);
nor U29977 (N_29977,N_18812,N_16426);
or U29978 (N_29978,N_11194,N_12653);
and U29979 (N_29979,N_11532,N_11341);
nand U29980 (N_29980,N_16478,N_15668);
nand U29981 (N_29981,N_17048,N_17201);
nor U29982 (N_29982,N_18365,N_15725);
nand U29983 (N_29983,N_16964,N_12143);
nand U29984 (N_29984,N_10514,N_10219);
or U29985 (N_29985,N_14172,N_18972);
or U29986 (N_29986,N_10156,N_15339);
xor U29987 (N_29987,N_17718,N_10213);
or U29988 (N_29988,N_12392,N_15860);
nand U29989 (N_29989,N_19493,N_19397);
or U29990 (N_29990,N_10136,N_17672);
and U29991 (N_29991,N_11181,N_18933);
and U29992 (N_29992,N_10937,N_14040);
or U29993 (N_29993,N_14570,N_14207);
nand U29994 (N_29994,N_10753,N_14409);
nand U29995 (N_29995,N_15948,N_11410);
nor U29996 (N_29996,N_10402,N_18905);
nor U29997 (N_29997,N_15937,N_10948);
and U29998 (N_29998,N_18271,N_10199);
nand U29999 (N_29999,N_17700,N_18890);
or UO_0 (O_0,N_23550,N_24209);
and UO_1 (O_1,N_29612,N_27208);
nand UO_2 (O_2,N_26906,N_24771);
and UO_3 (O_3,N_23044,N_22577);
nor UO_4 (O_4,N_25804,N_21294);
and UO_5 (O_5,N_26668,N_29720);
nand UO_6 (O_6,N_28555,N_29064);
and UO_7 (O_7,N_20318,N_22703);
or UO_8 (O_8,N_25377,N_26714);
and UO_9 (O_9,N_23470,N_21240);
nand UO_10 (O_10,N_23201,N_27196);
nor UO_11 (O_11,N_29051,N_25882);
or UO_12 (O_12,N_23880,N_28556);
nor UO_13 (O_13,N_24075,N_22866);
nand UO_14 (O_14,N_22569,N_27479);
nor UO_15 (O_15,N_28274,N_22877);
or UO_16 (O_16,N_27298,N_24205);
and UO_17 (O_17,N_28641,N_24244);
or UO_18 (O_18,N_29717,N_28020);
xnor UO_19 (O_19,N_22677,N_25610);
or UO_20 (O_20,N_29413,N_25317);
nand UO_21 (O_21,N_23850,N_27581);
nand UO_22 (O_22,N_29588,N_27958);
or UO_23 (O_23,N_22054,N_25982);
and UO_24 (O_24,N_24939,N_20631);
and UO_25 (O_25,N_25360,N_25479);
nor UO_26 (O_26,N_24651,N_28771);
nand UO_27 (O_27,N_21079,N_20798);
nand UO_28 (O_28,N_23456,N_24758);
nor UO_29 (O_29,N_21332,N_20744);
nand UO_30 (O_30,N_20804,N_29796);
or UO_31 (O_31,N_25945,N_24826);
and UO_32 (O_32,N_27407,N_23326);
or UO_33 (O_33,N_21333,N_20557);
nor UO_34 (O_34,N_21329,N_28270);
or UO_35 (O_35,N_20877,N_24439);
nand UO_36 (O_36,N_25128,N_26918);
and UO_37 (O_37,N_24585,N_25907);
nor UO_38 (O_38,N_28924,N_21437);
or UO_39 (O_39,N_28891,N_22587);
or UO_40 (O_40,N_20600,N_26180);
or UO_41 (O_41,N_21824,N_25954);
and UO_42 (O_42,N_26027,N_23962);
and UO_43 (O_43,N_29647,N_23764);
and UO_44 (O_44,N_28315,N_25287);
or UO_45 (O_45,N_25567,N_22558);
or UO_46 (O_46,N_20442,N_28597);
or UO_47 (O_47,N_29113,N_22408);
nor UO_48 (O_48,N_27367,N_25406);
nand UO_49 (O_49,N_27275,N_28467);
nor UO_50 (O_50,N_24370,N_22377);
nor UO_51 (O_51,N_21120,N_29462);
and UO_52 (O_52,N_21905,N_24516);
and UO_53 (O_53,N_20917,N_28674);
and UO_54 (O_54,N_24317,N_20421);
nor UO_55 (O_55,N_20361,N_24621);
or UO_56 (O_56,N_21110,N_28265);
and UO_57 (O_57,N_20757,N_23282);
nand UO_58 (O_58,N_23695,N_28455);
and UO_59 (O_59,N_26012,N_28650);
or UO_60 (O_60,N_27541,N_28694);
or UO_61 (O_61,N_23637,N_23689);
and UO_62 (O_62,N_28195,N_23337);
nor UO_63 (O_63,N_27030,N_29599);
nand UO_64 (O_64,N_27097,N_20383);
nor UO_65 (O_65,N_24490,N_22177);
nand UO_66 (O_66,N_27144,N_25266);
nor UO_67 (O_67,N_25591,N_20552);
and UO_68 (O_68,N_21596,N_21526);
and UO_69 (O_69,N_25526,N_25796);
nand UO_70 (O_70,N_27133,N_23501);
or UO_71 (O_71,N_26069,N_27856);
and UO_72 (O_72,N_23538,N_21452);
nor UO_73 (O_73,N_21516,N_27558);
and UO_74 (O_74,N_23994,N_23085);
nor UO_75 (O_75,N_23448,N_28025);
or UO_76 (O_76,N_20182,N_21132);
and UO_77 (O_77,N_28197,N_22501);
nor UO_78 (O_78,N_29334,N_23471);
nor UO_79 (O_79,N_28140,N_21392);
or UO_80 (O_80,N_22679,N_27207);
nor UO_81 (O_81,N_21037,N_24068);
and UO_82 (O_82,N_22393,N_25151);
or UO_83 (O_83,N_26962,N_27811);
nand UO_84 (O_84,N_28392,N_22331);
nor UO_85 (O_85,N_26643,N_24387);
nand UO_86 (O_86,N_22832,N_22634);
nor UO_87 (O_87,N_20080,N_22388);
nand UO_88 (O_88,N_22034,N_28456);
and UO_89 (O_89,N_25502,N_27072);
nand UO_90 (O_90,N_24334,N_26353);
or UO_91 (O_91,N_29663,N_25017);
and UO_92 (O_92,N_26449,N_22508);
nor UO_93 (O_93,N_28581,N_22528);
nor UO_94 (O_94,N_24899,N_29811);
and UO_95 (O_95,N_24905,N_23883);
nor UO_96 (O_96,N_24375,N_21029);
nand UO_97 (O_97,N_26859,N_23600);
or UO_98 (O_98,N_24301,N_25076);
nor UO_99 (O_99,N_27778,N_29311);
nor UO_100 (O_100,N_23826,N_27664);
nor UO_101 (O_101,N_25941,N_28171);
nor UO_102 (O_102,N_21365,N_25776);
nand UO_103 (O_103,N_23528,N_29161);
and UO_104 (O_104,N_29314,N_27396);
or UO_105 (O_105,N_25095,N_20833);
or UO_106 (O_106,N_20957,N_26589);
nand UO_107 (O_107,N_20579,N_24887);
nor UO_108 (O_108,N_23278,N_27068);
nor UO_109 (O_109,N_22067,N_26140);
nand UO_110 (O_110,N_21755,N_24818);
nand UO_111 (O_111,N_21920,N_24610);
nor UO_112 (O_112,N_26342,N_29346);
nor UO_113 (O_113,N_24389,N_29887);
and UO_114 (O_114,N_20312,N_25346);
nor UO_115 (O_115,N_22580,N_21344);
nand UO_116 (O_116,N_26766,N_25981);
nor UO_117 (O_117,N_25558,N_22227);
and UO_118 (O_118,N_29215,N_23646);
and UO_119 (O_119,N_25938,N_25555);
nand UO_120 (O_120,N_25738,N_29292);
and UO_121 (O_121,N_22430,N_20072);
nand UO_122 (O_122,N_27901,N_29250);
nor UO_123 (O_123,N_28476,N_22032);
nor UO_124 (O_124,N_21853,N_20984);
nand UO_125 (O_125,N_22573,N_21008);
or UO_126 (O_126,N_22390,N_29231);
nor UO_127 (O_127,N_24745,N_27004);
and UO_128 (O_128,N_26059,N_28783);
and UO_129 (O_129,N_26779,N_24757);
nand UO_130 (O_130,N_28369,N_29828);
nor UO_131 (O_131,N_29926,N_24854);
and UO_132 (O_132,N_25278,N_26147);
nor UO_133 (O_133,N_21814,N_22785);
nor UO_134 (O_134,N_27355,N_21434);
or UO_135 (O_135,N_20228,N_23878);
or UO_136 (O_136,N_26210,N_25177);
and UO_137 (O_137,N_24865,N_26983);
and UO_138 (O_138,N_28287,N_26098);
nor UO_139 (O_139,N_28178,N_20776);
nor UO_140 (O_140,N_21337,N_24279);
and UO_141 (O_141,N_21607,N_24481);
or UO_142 (O_142,N_25989,N_24442);
nand UO_143 (O_143,N_24984,N_23908);
or UO_144 (O_144,N_22555,N_22953);
or UO_145 (O_145,N_23595,N_23210);
and UO_146 (O_146,N_24568,N_25734);
nand UO_147 (O_147,N_26767,N_22814);
and UO_148 (O_148,N_21559,N_22346);
nand UO_149 (O_149,N_26396,N_27807);
or UO_150 (O_150,N_23645,N_21749);
nand UO_151 (O_151,N_27404,N_25331);
and UO_152 (O_152,N_25966,N_26054);
nand UO_153 (O_153,N_22925,N_22014);
nor UO_154 (O_154,N_24801,N_20812);
nand UO_155 (O_155,N_23332,N_27334);
nand UO_156 (O_156,N_23353,N_23788);
and UO_157 (O_157,N_24584,N_29744);
nand UO_158 (O_158,N_23340,N_23674);
and UO_159 (O_159,N_22912,N_23609);
nor UO_160 (O_160,N_28857,N_21797);
or UO_161 (O_161,N_22869,N_22052);
nor UO_162 (O_162,N_26421,N_23774);
nand UO_163 (O_163,N_28010,N_23145);
nand UO_164 (O_164,N_24234,N_23296);
and UO_165 (O_165,N_25054,N_23925);
and UO_166 (O_166,N_29546,N_26478);
nor UO_167 (O_167,N_27098,N_25984);
or UO_168 (O_168,N_28344,N_20909);
or UO_169 (O_169,N_23696,N_23924);
or UO_170 (O_170,N_21599,N_23205);
or UO_171 (O_171,N_24581,N_28930);
nand UO_172 (O_172,N_28434,N_28914);
and UO_173 (O_173,N_21992,N_20771);
or UO_174 (O_174,N_26521,N_25566);
or UO_175 (O_175,N_22300,N_29089);
nand UO_176 (O_176,N_20304,N_25288);
nor UO_177 (O_177,N_26924,N_20920);
nor UO_178 (O_178,N_20605,N_23023);
and UO_179 (O_179,N_22094,N_25474);
and UO_180 (O_180,N_28114,N_29187);
or UO_181 (O_181,N_29875,N_24534);
or UO_182 (O_182,N_27863,N_21861);
or UO_183 (O_183,N_29147,N_26765);
nand UO_184 (O_184,N_28882,N_20211);
xnor UO_185 (O_185,N_27126,N_25090);
or UO_186 (O_186,N_27488,N_27322);
or UO_187 (O_187,N_24619,N_26952);
or UO_188 (O_188,N_24989,N_21153);
and UO_189 (O_189,N_27136,N_23395);
or UO_190 (O_190,N_24125,N_28093);
or UO_191 (O_191,N_26335,N_21665);
and UO_192 (O_192,N_27038,N_21378);
or UO_193 (O_193,N_29635,N_27255);
and UO_194 (O_194,N_22842,N_29754);
and UO_195 (O_195,N_28569,N_26124);
or UO_196 (O_196,N_26846,N_23983);
or UO_197 (O_197,N_21976,N_22383);
nand UO_198 (O_198,N_24257,N_26037);
and UO_199 (O_199,N_26754,N_25258);
nand UO_200 (O_200,N_24819,N_27105);
nor UO_201 (O_201,N_29065,N_22374);
xor UO_202 (O_202,N_26686,N_24299);
nand UO_203 (O_203,N_26062,N_29235);
or UO_204 (O_204,N_24091,N_21324);
nor UO_205 (O_205,N_23539,N_29383);
nor UO_206 (O_206,N_24102,N_21948);
or UO_207 (O_207,N_24893,N_26169);
nand UO_208 (O_208,N_24582,N_25390);
nand UO_209 (O_209,N_25767,N_27673);
and UO_210 (O_210,N_26129,N_24248);
or UO_211 (O_211,N_27061,N_26712);
or UO_212 (O_212,N_25753,N_25049);
and UO_213 (O_213,N_26826,N_23874);
nor UO_214 (O_214,N_28090,N_27041);
or UO_215 (O_215,N_29143,N_29670);
nor UO_216 (O_216,N_27882,N_28451);
nor UO_217 (O_217,N_28550,N_25862);
and UO_218 (O_218,N_21027,N_20689);
and UO_219 (O_219,N_27333,N_22329);
or UO_220 (O_220,N_22541,N_28798);
or UO_221 (O_221,N_26785,N_23492);
nor UO_222 (O_222,N_20396,N_27709);
nand UO_223 (O_223,N_22285,N_29050);
nor UO_224 (O_224,N_27537,N_29764);
nand UO_225 (O_225,N_28637,N_29418);
nand UO_226 (O_226,N_27375,N_26897);
and UO_227 (O_227,N_24167,N_20963);
or UO_228 (O_228,N_20912,N_29700);
nand UO_229 (O_229,N_29211,N_21161);
nor UO_230 (O_230,N_28929,N_26901);
nor UO_231 (O_231,N_28916,N_24054);
or UO_232 (O_232,N_28207,N_25570);
or UO_233 (O_233,N_26743,N_20189);
and UO_234 (O_234,N_27576,N_21021);
or UO_235 (O_235,N_29535,N_24788);
nor UO_236 (O_236,N_22975,N_22263);
and UO_237 (O_237,N_28164,N_25645);
nand UO_238 (O_238,N_29169,N_22579);
nor UO_239 (O_239,N_24652,N_23493);
and UO_240 (O_240,N_23691,N_24286);
nand UO_241 (O_241,N_28756,N_25276);
and UO_242 (O_242,N_20246,N_21511);
nand UO_243 (O_243,N_27477,N_23946);
nand UO_244 (O_244,N_24747,N_29073);
nor UO_245 (O_245,N_23710,N_22209);
and UO_246 (O_246,N_21733,N_21321);
and UO_247 (O_247,N_24936,N_26536);
nor UO_248 (O_248,N_27777,N_24417);
and UO_249 (O_249,N_21191,N_25808);
nand UO_250 (O_250,N_29677,N_21226);
nor UO_251 (O_251,N_29731,N_23923);
nor UO_252 (O_252,N_26261,N_29648);
or UO_253 (O_253,N_29365,N_21560);
and UO_254 (O_254,N_24855,N_26959);
and UO_255 (O_255,N_27867,N_28268);
nand UO_256 (O_256,N_26373,N_20352);
nand UO_257 (O_257,N_21388,N_26013);
or UO_258 (O_258,N_22255,N_22906);
and UO_259 (O_259,N_26091,N_26305);
nor UO_260 (O_260,N_24391,N_23428);
nand UO_261 (O_261,N_27115,N_29316);
and UO_262 (O_262,N_29208,N_24972);
or UO_263 (O_263,N_25120,N_26240);
and UO_264 (O_264,N_24265,N_27326);
and UO_265 (O_265,N_23629,N_28810);
and UO_266 (O_266,N_27570,N_29990);
nor UO_267 (O_267,N_24253,N_28781);
nor UO_268 (O_268,N_22556,N_20648);
and UO_269 (O_269,N_22559,N_29276);
nand UO_270 (O_270,N_20043,N_29358);
nor UO_271 (O_271,N_26250,N_24919);
nand UO_272 (O_272,N_29234,N_25313);
and UO_273 (O_273,N_23562,N_23972);
or UO_274 (O_274,N_24933,N_25033);
or UO_275 (O_275,N_25368,N_21631);
or UO_276 (O_276,N_28393,N_22804);
and UO_277 (O_277,N_25300,N_26651);
and UO_278 (O_278,N_28230,N_25219);
or UO_279 (O_279,N_24674,N_23254);
and UO_280 (O_280,N_21835,N_21427);
nor UO_281 (O_281,N_27923,N_23522);
or UO_282 (O_282,N_25135,N_23363);
nand UO_283 (O_283,N_20588,N_23662);
nor UO_284 (O_284,N_26400,N_28868);
nand UO_285 (O_285,N_21468,N_28016);
and UO_286 (O_286,N_26707,N_24115);
and UO_287 (O_287,N_24675,N_28349);
nor UO_288 (O_288,N_27135,N_24243);
nor UO_289 (O_289,N_24073,N_21401);
and UO_290 (O_290,N_20104,N_26768);
and UO_291 (O_291,N_24533,N_26220);
nand UO_292 (O_292,N_29149,N_27700);
or UO_293 (O_293,N_25028,N_23921);
or UO_294 (O_294,N_21315,N_21421);
and UO_295 (O_295,N_27185,N_22334);
and UO_296 (O_296,N_20423,N_24093);
or UO_297 (O_297,N_29706,N_23716);
nand UO_298 (O_298,N_26822,N_25792);
or UO_299 (O_299,N_23270,N_21993);
nand UO_300 (O_300,N_28473,N_26885);
nand UO_301 (O_301,N_25861,N_22619);
nor UO_302 (O_302,N_24394,N_23938);
or UO_303 (O_303,N_22483,N_24660);
nand UO_304 (O_304,N_23967,N_25158);
and UO_305 (O_305,N_25361,N_27270);
nand UO_306 (O_306,N_24733,N_21305);
nand UO_307 (O_307,N_25963,N_28224);
or UO_308 (O_308,N_23833,N_24839);
or UO_309 (O_309,N_21154,N_28128);
or UO_310 (O_310,N_20767,N_29692);
or UO_311 (O_311,N_22515,N_28867);
nor UO_312 (O_312,N_21269,N_20432);
and UO_313 (O_313,N_21568,N_22042);
nor UO_314 (O_314,N_27090,N_25829);
and UO_315 (O_315,N_21685,N_27391);
and UO_316 (O_316,N_26105,N_21571);
and UO_317 (O_317,N_23916,N_23074);
and UO_318 (O_318,N_20092,N_21639);
or UO_319 (O_319,N_25928,N_23066);
and UO_320 (O_320,N_22931,N_23312);
and UO_321 (O_321,N_26231,N_20366);
nand UO_322 (O_322,N_23378,N_29180);
nand UO_323 (O_323,N_23840,N_21082);
nand UO_324 (O_324,N_25762,N_29725);
and UO_325 (O_325,N_29908,N_24006);
nand UO_326 (O_326,N_26269,N_28541);
and UO_327 (O_327,N_22010,N_25670);
or UO_328 (O_328,N_20796,N_24732);
or UO_329 (O_329,N_20167,N_26288);
nor UO_330 (O_330,N_25402,N_29968);
nand UO_331 (O_331,N_20285,N_24037);
nor UO_332 (O_332,N_26595,N_29103);
or UO_333 (O_333,N_26040,N_23435);
or UO_334 (O_334,N_29502,N_25209);
or UO_335 (O_335,N_23888,N_29326);
nand UO_336 (O_336,N_26836,N_28013);
nor UO_337 (O_337,N_29296,N_23990);
and UO_338 (O_338,N_21695,N_24668);
or UO_339 (O_339,N_28352,N_28296);
or UO_340 (O_340,N_23286,N_21032);
nand UO_341 (O_341,N_22516,N_20682);
xor UO_342 (O_342,N_28193,N_23982);
nor UO_343 (O_343,N_22917,N_23365);
nor UO_344 (O_344,N_26513,N_23364);
and UO_345 (O_345,N_21455,N_29989);
nand UO_346 (O_346,N_26283,N_23277);
nor UO_347 (O_347,N_26183,N_26404);
and UO_348 (O_348,N_22936,N_23310);
or UO_349 (O_349,N_23051,N_28559);
nand UO_350 (O_350,N_23614,N_28062);
or UO_351 (O_351,N_24261,N_21762);
and UO_352 (O_352,N_25409,N_29821);
or UO_353 (O_353,N_29364,N_28667);
nand UO_354 (O_354,N_24691,N_24474);
and UO_355 (O_355,N_20184,N_29529);
nor UO_356 (O_356,N_20407,N_27306);
nor UO_357 (O_357,N_23249,N_28614);
nand UO_358 (O_358,N_25060,N_29660);
and UO_359 (O_359,N_20082,N_27337);
nor UO_360 (O_360,N_23742,N_22305);
nand UO_361 (O_361,N_27940,N_29911);
nor UO_362 (O_362,N_25512,N_27473);
or UO_363 (O_363,N_20333,N_21717);
or UO_364 (O_364,N_20234,N_21508);
nor UO_365 (O_365,N_26115,N_21999);
or UO_366 (O_366,N_24482,N_27766);
and UO_367 (O_367,N_21464,N_24774);
nand UO_368 (O_368,N_29129,N_28416);
and UO_369 (O_369,N_22186,N_27691);
or UO_370 (O_370,N_25321,N_22018);
and UO_371 (O_371,N_23441,N_25475);
and UO_372 (O_372,N_29685,N_26299);
nand UO_373 (O_373,N_21147,N_26413);
or UO_374 (O_374,N_22947,N_23451);
nand UO_375 (O_375,N_25681,N_25501);
nor UO_376 (O_376,N_28079,N_29701);
or UO_377 (O_377,N_24531,N_27455);
nor UO_378 (O_378,N_23827,N_23536);
and UO_379 (O_379,N_22586,N_29808);
and UO_380 (O_380,N_22273,N_28158);
nor UO_381 (O_381,N_28505,N_22357);
nor UO_382 (O_382,N_23811,N_20438);
nand UO_383 (O_383,N_20156,N_20779);
nor UO_384 (O_384,N_26516,N_23179);
or UO_385 (O_385,N_27545,N_20295);
or UO_386 (O_386,N_24084,N_21831);
nand UO_387 (O_387,N_28673,N_28886);
or UO_388 (O_388,N_28169,N_27836);
nand UO_389 (O_389,N_27213,N_24931);
nor UO_390 (O_390,N_22288,N_22985);
or UO_391 (O_391,N_22222,N_26296);
and UO_392 (O_392,N_20976,N_23639);
nand UO_393 (O_393,N_21961,N_27893);
nor UO_394 (O_394,N_29912,N_28028);
or UO_395 (O_395,N_25318,N_22883);
or UO_396 (O_396,N_29179,N_24492);
nand UO_397 (O_397,N_21909,N_27212);
nor UO_398 (O_398,N_22544,N_21164);
nand UO_399 (O_399,N_20549,N_21100);
or UO_400 (O_400,N_28679,N_21293);
nor UO_401 (O_401,N_25369,N_23948);
or UO_402 (O_402,N_24971,N_20847);
nand UO_403 (O_403,N_25186,N_27127);
nand UO_404 (O_404,N_22782,N_21043);
xnor UO_405 (O_405,N_27342,N_27027);
nand UO_406 (O_406,N_28704,N_20244);
or UO_407 (O_407,N_28995,N_28979);
nand UO_408 (O_408,N_25545,N_25880);
or UO_409 (O_409,N_26555,N_23260);
and UO_410 (O_410,N_22728,N_27518);
or UO_411 (O_411,N_25348,N_23701);
nand UO_412 (O_412,N_20801,N_28484);
nand UO_413 (O_413,N_23911,N_25611);
and UO_414 (O_414,N_26411,N_24105);
or UO_415 (O_415,N_28594,N_21202);
nor UO_416 (O_416,N_28452,N_23869);
nor UO_417 (O_417,N_21986,N_28466);
nor UO_418 (O_418,N_23980,N_27640);
nand UO_419 (O_419,N_23841,N_20155);
and UO_420 (O_420,N_21977,N_28173);
nand UO_421 (O_421,N_23581,N_29784);
or UO_422 (O_422,N_29841,N_24728);
or UO_423 (O_423,N_29831,N_20654);
or UO_424 (O_424,N_26533,N_27336);
nand UO_425 (O_425,N_27183,N_27625);
nand UO_426 (O_426,N_26356,N_26370);
nor UO_427 (O_427,N_21471,N_24550);
nor UO_428 (O_428,N_27344,N_21972);
nor UO_429 (O_429,N_21348,N_25916);
and UO_430 (O_430,N_22495,N_28699);
or UO_431 (O_431,N_20921,N_28335);
nor UO_432 (O_432,N_20529,N_24805);
or UO_433 (O_433,N_25314,N_23437);
nand UO_434 (O_434,N_20011,N_27107);
and UO_435 (O_435,N_21442,N_20695);
and UO_436 (O_436,N_29843,N_23516);
and UO_437 (O_437,N_20843,N_29712);
and UO_438 (O_438,N_21381,N_27075);
nand UO_439 (O_439,N_27617,N_28426);
nand UO_440 (O_440,N_24990,N_23618);
or UO_441 (O_441,N_21418,N_28774);
nand UO_442 (O_442,N_26033,N_20158);
nor UO_443 (O_443,N_29146,N_25865);
nand UO_444 (O_444,N_22540,N_23951);
and UO_445 (O_445,N_21433,N_29625);
or UO_446 (O_446,N_24049,N_26730);
or UO_447 (O_447,N_23915,N_26491);
or UO_448 (O_448,N_21912,N_20255);
and UO_449 (O_449,N_22595,N_26178);
or UO_450 (O_450,N_22174,N_28490);
or UO_451 (O_451,N_22621,N_26499);
and UO_452 (O_452,N_24074,N_20797);
and UO_453 (O_453,N_25002,N_29572);
and UO_454 (O_454,N_27109,N_21641);
nand UO_455 (O_455,N_28913,N_26688);
or UO_456 (O_456,N_20057,N_26067);
and UO_457 (O_457,N_25023,N_20586);
nand UO_458 (O_458,N_27274,N_25517);
nor UO_459 (O_459,N_25615,N_24506);
nand UO_460 (O_460,N_22570,N_23008);
nand UO_461 (O_461,N_24880,N_20886);
and UO_462 (O_462,N_23237,N_20416);
nor UO_463 (O_463,N_20967,N_23605);
or UO_464 (O_464,N_21454,N_24731);
and UO_465 (O_465,N_23117,N_27876);
nand UO_466 (O_466,N_22281,N_22125);
nand UO_467 (O_467,N_25602,N_28424);
or UO_468 (O_468,N_26236,N_28241);
or UO_469 (O_469,N_25943,N_29438);
or UO_470 (O_470,N_25616,N_25749);
nand UO_471 (O_471,N_25366,N_27154);
nand UO_472 (O_472,N_20379,N_22387);
nand UO_473 (O_473,N_24557,N_25304);
or UO_474 (O_474,N_23047,N_27990);
or UO_475 (O_475,N_29405,N_29549);
nand UO_476 (O_476,N_22128,N_24415);
or UO_477 (O_477,N_27378,N_24583);
nor UO_478 (O_478,N_20271,N_20709);
nor UO_479 (O_479,N_27529,N_20788);
or UO_480 (O_480,N_25710,N_29927);
or UO_481 (O_481,N_25550,N_29212);
nand UO_482 (O_482,N_26644,N_29636);
nand UO_483 (O_483,N_24716,N_20959);
and UO_484 (O_484,N_28759,N_27401);
or UO_485 (O_485,N_26815,N_20764);
nor UO_486 (O_486,N_21251,N_25872);
nor UO_487 (O_487,N_27774,N_23615);
and UO_488 (O_488,N_27040,N_28259);
nand UO_489 (O_489,N_21795,N_25335);
nor UO_490 (O_490,N_25625,N_26034);
and UO_491 (O_491,N_21543,N_21866);
nor UO_492 (O_492,N_23945,N_28498);
nand UO_493 (O_493,N_28561,N_26927);
nand UO_494 (O_494,N_20275,N_20229);
nand UO_495 (O_495,N_21754,N_24395);
or UO_496 (O_496,N_27989,N_22690);
or UO_497 (O_497,N_27631,N_20212);
nand UO_498 (O_498,N_29415,N_28937);
nand UO_499 (O_499,N_28821,N_29807);
or UO_500 (O_500,N_20621,N_26453);
or UO_501 (O_501,N_24618,N_27066);
and UO_502 (O_502,N_20934,N_29246);
nand UO_503 (O_503,N_25063,N_24240);
nor UO_504 (O_504,N_23090,N_22192);
or UO_505 (O_505,N_25196,N_29302);
nor UO_506 (O_506,N_20486,N_23466);
and UO_507 (O_507,N_23391,N_24194);
or UO_508 (O_508,N_29822,N_26979);
nand UO_509 (O_509,N_29964,N_27172);
nor UO_510 (O_510,N_25283,N_25432);
and UO_511 (O_511,N_22686,N_27044);
and UO_512 (O_512,N_26192,N_22797);
or UO_513 (O_513,N_25900,N_23534);
nand UO_514 (O_514,N_26384,N_23617);
nor UO_515 (O_515,N_25606,N_27690);
nand UO_516 (O_516,N_24891,N_26136);
or UO_517 (O_517,N_24714,N_20944);
nor UO_518 (O_518,N_29870,N_21969);
or UO_519 (O_519,N_24849,N_23527);
nand UO_520 (O_520,N_24942,N_27289);
or UO_521 (O_521,N_27972,N_29188);
nand UO_522 (O_522,N_22873,N_20310);
nand UO_523 (O_523,N_24178,N_23533);
or UO_524 (O_524,N_28727,N_22860);
or UO_525 (O_525,N_25815,N_22824);
nor UO_526 (O_526,N_24567,N_29689);
nor UO_527 (O_527,N_22594,N_28333);
nor UO_528 (O_528,N_21914,N_28531);
and UO_529 (O_529,N_25724,N_27840);
nand UO_530 (O_530,N_28862,N_24457);
nor UO_531 (O_531,N_26827,N_21005);
or UO_532 (O_532,N_28383,N_20242);
nor UO_533 (O_533,N_25967,N_26986);
and UO_534 (O_534,N_23986,N_23648);
and UO_535 (O_535,N_23784,N_21857);
or UO_536 (O_536,N_29671,N_21081);
and UO_537 (O_537,N_23120,N_21751);
nor UO_538 (O_538,N_20405,N_21156);
and UO_539 (O_539,N_25215,N_23045);
nand UO_540 (O_540,N_21459,N_24296);
and UO_541 (O_541,N_22927,N_24131);
xnor UO_542 (O_542,N_23239,N_28181);
nor UO_543 (O_543,N_25089,N_27902);
nor UO_544 (O_544,N_24454,N_23014);
or UO_545 (O_545,N_26509,N_23535);
and UO_546 (O_546,N_24410,N_26185);
nor UO_547 (O_547,N_20273,N_23782);
nand UO_548 (O_548,N_28277,N_27308);
nand UO_549 (O_549,N_26944,N_24070);
or UO_550 (O_550,N_26806,N_25843);
and UO_551 (O_551,N_23439,N_27663);
nor UO_552 (O_552,N_22773,N_27903);
nor UO_553 (O_553,N_26658,N_22812);
and UO_554 (O_554,N_26319,N_29315);
and UO_555 (O_555,N_24883,N_22693);
or UO_556 (O_556,N_25812,N_25789);
and UO_557 (O_557,N_23974,N_26244);
and UO_558 (O_558,N_22928,N_29580);
nor UO_559 (O_559,N_21128,N_26079);
or UO_560 (O_560,N_28825,N_27359);
or UO_561 (O_561,N_26753,N_24413);
and UO_562 (O_562,N_27079,N_26560);
nor UO_563 (O_563,N_24349,N_23634);
nor UO_564 (O_564,N_22744,N_21386);
or UO_565 (O_565,N_26426,N_21359);
or UO_566 (O_566,N_29124,N_26969);
and UO_567 (O_567,N_23622,N_22930);
nor UO_568 (O_568,N_26976,N_20100);
nand UO_569 (O_569,N_29293,N_23461);
nor UO_570 (O_570,N_26122,N_25344);
nor UO_571 (O_571,N_23495,N_21771);
nand UO_572 (O_572,N_22132,N_27737);
nor UO_573 (O_573,N_25417,N_28992);
and UO_574 (O_574,N_28293,N_28219);
nand UO_575 (O_575,N_28457,N_24340);
or UO_576 (O_576,N_20629,N_25066);
nor UO_577 (O_577,N_25251,N_29907);
nor UO_578 (O_578,N_26649,N_24544);
or UO_579 (O_579,N_20443,N_25687);
and UO_580 (O_580,N_27280,N_22981);
or UO_581 (O_581,N_26923,N_23769);
or UO_582 (O_582,N_25523,N_29794);
nand UO_583 (O_583,N_20402,N_29597);
nand UO_584 (O_584,N_27197,N_21941);
or UO_585 (O_585,N_26341,N_27469);
nor UO_586 (O_586,N_25078,N_27028);
or UO_587 (O_587,N_22959,N_24983);
and UO_588 (O_588,N_29531,N_22131);
and UO_589 (O_589,N_29854,N_25021);
and UO_590 (O_590,N_25944,N_20400);
nand UO_591 (O_591,N_23154,N_23889);
nor UO_592 (O_592,N_25297,N_25922);
or UO_593 (O_593,N_22863,N_21463);
and UO_594 (O_594,N_29034,N_22142);
or UO_595 (O_595,N_27203,N_25412);
nor UO_596 (O_596,N_21657,N_20759);
nor UO_597 (O_597,N_29335,N_29144);
and UO_598 (O_598,N_22440,N_22164);
or UO_599 (O_599,N_25786,N_26566);
and UO_600 (O_600,N_25323,N_25118);
or UO_601 (O_601,N_22002,N_27732);
nand UO_602 (O_602,N_29915,N_29463);
and UO_603 (O_603,N_28278,N_21565);
nand UO_604 (O_604,N_25571,N_28624);
nand UO_605 (O_605,N_29820,N_25870);
or UO_606 (O_606,N_25464,N_20842);
and UO_607 (O_607,N_29221,N_28680);
nand UO_608 (O_608,N_25978,N_29936);
nor UO_609 (O_609,N_22520,N_23262);
nor UO_610 (O_610,N_20907,N_20925);
or UO_611 (O_611,N_29929,N_28520);
or UO_612 (O_612,N_21242,N_24650);
or UO_613 (O_613,N_23699,N_20568);
and UO_614 (O_614,N_27065,N_23800);
nor UO_615 (O_615,N_22598,N_29946);
nor UO_616 (O_616,N_20997,N_29424);
nor UO_617 (O_617,N_22037,N_26622);
nor UO_618 (O_618,N_20683,N_27948);
and UO_619 (O_619,N_28718,N_28787);
nand UO_620 (O_620,N_21819,N_23656);
nand UO_621 (O_621,N_28184,N_26100);
nor UO_622 (O_622,N_29168,N_28856);
and UO_623 (O_623,N_25587,N_25126);
and UO_624 (O_624,N_22348,N_24672);
nor UO_625 (O_625,N_20497,N_21549);
nor UO_626 (O_626,N_26285,N_29425);
nor UO_627 (O_627,N_27281,N_21767);
or UO_628 (O_628,N_28433,N_21684);
nand UO_629 (O_629,N_22058,N_24719);
or UO_630 (O_630,N_24499,N_24269);
or UO_631 (O_631,N_22013,N_22428);
nor UO_632 (O_632,N_20918,N_25399);
and UO_633 (O_633,N_29253,N_28340);
or UO_634 (O_634,N_21638,N_24232);
nand UO_635 (O_635,N_22810,N_28799);
nor UO_636 (O_636,N_24762,N_24712);
nand UO_637 (O_637,N_26857,N_20686);
or UO_638 (O_638,N_22371,N_25492);
and UO_639 (O_639,N_23714,N_24468);
or UO_640 (O_640,N_28552,N_26325);
and UO_641 (O_641,N_20950,N_20954);
or UO_642 (O_642,N_29000,N_26063);
nor UO_643 (O_643,N_28938,N_23294);
nor UO_644 (O_644,N_26810,N_22498);
nor UO_645 (O_645,N_20985,N_20994);
and UO_646 (O_646,N_25431,N_22886);
nor UO_647 (O_647,N_22768,N_29856);
nand UO_648 (O_648,N_22818,N_29381);
or UO_649 (O_649,N_24536,N_25778);
nand UO_650 (O_650,N_29570,N_27215);
and UO_651 (O_651,N_22775,N_29963);
or UO_652 (O_652,N_22675,N_26866);
nand UO_653 (O_653,N_29166,N_29097);
nand UO_654 (O_654,N_27348,N_23610);
or UO_655 (O_655,N_27679,N_24042);
nand UO_656 (O_656,N_27629,N_24593);
or UO_657 (O_657,N_29458,N_22519);
nand UO_658 (O_658,N_28724,N_21786);
and UO_659 (O_659,N_26484,N_26280);
or UO_660 (O_660,N_26700,N_23557);
nor UO_661 (O_661,N_26398,N_28754);
or UO_662 (O_662,N_22948,N_20844);
nor UO_663 (O_663,N_23412,N_23193);
or UO_664 (O_664,N_27834,N_20520);
nor UO_665 (O_665,N_25677,N_20663);
nor UO_666 (O_666,N_25709,N_28469);
or UO_667 (O_667,N_27390,N_26594);
and UO_668 (O_668,N_24804,N_28870);
nor UO_669 (O_669,N_28308,N_29819);
nand UO_670 (O_670,N_27163,N_21501);
nand UO_671 (O_671,N_25743,N_26139);
nor UO_672 (O_672,N_28058,N_22176);
nor UO_673 (O_673,N_27908,N_20591);
or UO_674 (O_674,N_28738,N_21832);
or UO_675 (O_675,N_27123,N_21945);
nand UO_676 (O_676,N_29115,N_28437);
nand UO_677 (O_677,N_21577,N_22730);
nor UO_678 (O_678,N_28530,N_29779);
nor UO_679 (O_679,N_24441,N_26792);
or UO_680 (O_680,N_24840,N_22893);
nor UO_681 (O_681,N_25458,N_25232);
nand UO_682 (O_682,N_26562,N_23407);
nand UO_683 (O_683,N_21947,N_25557);
or UO_684 (O_684,N_25379,N_25388);
nand UO_685 (O_685,N_25716,N_25588);
nand UO_686 (O_686,N_26251,N_27233);
or UO_687 (O_687,N_23231,N_22436);
or UO_688 (O_688,N_24153,N_20544);
and UO_689 (O_689,N_20388,N_27287);
nand UO_690 (O_690,N_20585,N_29969);
nor UO_691 (O_691,N_25720,N_21227);
and UO_692 (O_692,N_29337,N_28925);
or UO_693 (O_693,N_27933,N_22859);
and UO_694 (O_694,N_27254,N_22189);
nor UO_695 (O_695,N_22332,N_27301);
nand UO_696 (O_696,N_21165,N_20538);
nor UO_697 (O_697,N_28073,N_26956);
or UO_698 (O_698,N_24142,N_29351);
nor UO_699 (O_699,N_22885,N_27965);
nand UO_700 (O_700,N_20566,N_27116);
nor UO_701 (O_701,N_22505,N_21297);
or UO_702 (O_702,N_21879,N_21782);
or UO_703 (O_703,N_23242,N_27253);
nor UO_704 (O_704,N_27555,N_20230);
nand UO_705 (O_705,N_25026,N_28005);
nand UO_706 (O_706,N_25350,N_28047);
and UO_707 (O_707,N_23899,N_22003);
nand UO_708 (O_708,N_28503,N_24467);
nand UO_709 (O_709,N_21439,N_27528);
and UO_710 (O_710,N_20928,N_24722);
nand UO_711 (O_711,N_20484,N_20728);
or UO_712 (O_712,N_28499,N_21644);
nand UO_713 (O_713,N_24109,N_26783);
nor UO_714 (O_714,N_29319,N_25110);
nor UO_715 (O_715,N_27548,N_28350);
or UO_716 (O_716,N_28880,N_27733);
or UO_717 (O_717,N_26995,N_29578);
nor UO_718 (O_718,N_28872,N_20163);
nor UO_719 (O_719,N_29940,N_22938);
nand UO_720 (O_720,N_25330,N_29813);
nor UO_721 (O_721,N_26585,N_27450);
nor UO_722 (O_722,N_26227,N_28752);
nand UO_723 (O_723,N_21445,N_26834);
nand UO_724 (O_724,N_26424,N_28851);
and UO_725 (O_725,N_26133,N_21591);
or UO_726 (O_726,N_27857,N_27500);
and UO_727 (O_727,N_23898,N_28255);
nand UO_728 (O_728,N_22992,N_20306);
nand UO_729 (O_729,N_27810,N_20483);
nand UO_730 (O_730,N_26257,N_22637);
or UO_731 (O_731,N_28736,N_27891);
or UO_732 (O_732,N_21523,N_26856);
nor UO_733 (O_733,N_29591,N_22397);
nand UO_734 (O_734,N_20809,N_21045);
or UO_735 (O_735,N_25263,N_27580);
nor UO_736 (O_736,N_25842,N_20009);
nand UO_737 (O_737,N_28210,N_22200);
or UO_738 (O_738,N_25204,N_24385);
xor UO_739 (O_739,N_25354,N_23027);
nand UO_740 (O_740,N_25542,N_26544);
nand UO_741 (O_741,N_25154,N_26399);
nor UO_742 (O_742,N_27100,N_25096);
or UO_743 (O_743,N_26855,N_25525);
nor UO_744 (O_744,N_25702,N_23304);
or UO_745 (O_745,N_24564,N_21680);
nand UO_746 (O_746,N_26719,N_29932);
and UO_747 (O_747,N_22705,N_23553);
and UO_748 (O_748,N_25279,N_23371);
nor UO_749 (O_749,N_25370,N_23421);
or UO_750 (O_750,N_23626,N_28567);
or UO_751 (O_751,N_23602,N_26690);
or UO_752 (O_752,N_22752,N_20935);
or UO_753 (O_753,N_21287,N_25576);
and UO_754 (O_754,N_27918,N_29356);
nor UO_755 (O_755,N_20725,N_23488);
and UO_756 (O_756,N_24678,N_24460);
or UO_757 (O_757,N_24790,N_28180);
nand UO_758 (O_758,N_22320,N_22135);
nor UO_759 (O_759,N_23103,N_28805);
and UO_760 (O_760,N_24563,N_26689);
nor UO_761 (O_761,N_20619,N_28261);
and UO_762 (O_762,N_24225,N_23158);
or UO_763 (O_763,N_23511,N_25841);
nor UO_764 (O_764,N_22517,N_28312);
or UO_765 (O_765,N_28779,N_21281);
and UO_766 (O_766,N_29773,N_26189);
and UO_767 (O_767,N_23564,N_25381);
and UO_768 (O_768,N_27033,N_26219);
and UO_769 (O_769,N_23866,N_27300);
or UO_770 (O_770,N_21563,N_21424);
nand UO_771 (O_771,N_21770,N_21811);
nor UO_772 (O_772,N_22016,N_25244);
and UO_773 (O_773,N_27104,N_28281);
or UO_774 (O_774,N_21175,N_27712);
and UO_775 (O_775,N_22477,N_28076);
nor UO_776 (O_776,N_23715,N_23099);
or UO_777 (O_777,N_23088,N_23787);
and UO_778 (O_778,N_22610,N_29299);
or UO_779 (O_779,N_25756,N_20617);
or UO_780 (O_780,N_25324,N_29522);
nor UO_781 (O_781,N_28646,N_28811);
nand UO_782 (O_782,N_28864,N_22438);
or UO_783 (O_783,N_23598,N_25062);
nand UO_784 (O_784,N_24017,N_27738);
or UO_785 (O_785,N_22386,N_28419);
or UO_786 (O_786,N_26692,N_29375);
nor UO_787 (O_787,N_23943,N_28208);
nor UO_788 (O_788,N_26415,N_21584);
or UO_789 (O_789,N_27719,N_23408);
nor UO_790 (O_790,N_27219,N_27941);
or UO_791 (O_791,N_25240,N_23829);
nand UO_792 (O_792,N_20408,N_26150);
nand UO_793 (O_793,N_24496,N_26438);
nor UO_794 (O_794,N_21031,N_22742);
or UO_795 (O_795,N_29001,N_21690);
nand UO_796 (O_796,N_22398,N_26429);
nor UO_797 (O_797,N_25238,N_25534);
nand UO_798 (O_798,N_25748,N_21148);
and UO_799 (O_799,N_29617,N_26583);
nand UO_800 (O_800,N_21431,N_24355);
nand UO_801 (O_801,N_20596,N_21958);
nor UO_802 (O_802,N_26604,N_21186);
or UO_803 (O_803,N_20702,N_20413);
or UO_804 (O_804,N_20110,N_24715);
and UO_805 (O_805,N_20819,N_22994);
nand UO_806 (O_806,N_28804,N_21592);
or UO_807 (O_807,N_21342,N_22568);
and UO_808 (O_808,N_20099,N_25983);
nor UO_809 (O_809,N_25635,N_26420);
or UO_810 (O_810,N_25535,N_24426);
nand UO_811 (O_811,N_27465,N_26940);
nor UO_812 (O_812,N_20206,N_25751);
nor UO_813 (O_813,N_29961,N_29489);
and UO_814 (O_814,N_20649,N_29571);
nor UO_815 (O_815,N_21285,N_28529);
or UO_816 (O_816,N_21859,N_26943);
or UO_817 (O_817,N_22311,N_27904);
and UO_818 (O_818,N_26871,N_29429);
and UO_819 (O_819,N_27535,N_27108);
nand UO_820 (O_820,N_23199,N_25294);
xnor UO_821 (O_821,N_25580,N_25707);
nand UO_822 (O_822,N_29366,N_23424);
and UO_823 (O_823,N_24684,N_21983);
nor UO_824 (O_824,N_28953,N_24844);
nor UO_825 (O_825,N_21363,N_20676);
nand UO_826 (O_826,N_23700,N_29446);
or UO_827 (O_827,N_23954,N_20204);
and UO_828 (O_828,N_28339,N_20718);
and UO_829 (O_829,N_23941,N_21055);
and UO_830 (O_830,N_21776,N_20034);
or UO_831 (O_831,N_24447,N_24004);
or UO_832 (O_832,N_25071,N_23436);
nand UO_833 (O_833,N_24053,N_28026);
or UO_834 (O_834,N_29735,N_22817);
and UO_835 (O_835,N_26021,N_24537);
nor UO_836 (O_836,N_23082,N_23490);
and UO_837 (O_837,N_26654,N_22097);
nand UO_838 (O_838,N_23257,N_22803);
and UO_839 (O_839,N_27470,N_20441);
nor UO_840 (O_840,N_21298,N_25662);
and UO_841 (O_841,N_26624,N_27037);
and UO_842 (O_842,N_20320,N_28571);
nor UO_843 (O_843,N_22811,N_22074);
and UO_844 (O_844,N_27858,N_21473);
nor UO_845 (O_845,N_20632,N_27981);
or UO_846 (O_846,N_23265,N_26161);
nand UO_847 (O_847,N_25895,N_20001);
nor UO_848 (O_848,N_26423,N_26964);
xnor UO_849 (O_849,N_24384,N_29576);
and UO_850 (O_850,N_22965,N_26186);
nand UO_851 (O_851,N_22103,N_29698);
or UO_852 (O_852,N_24493,N_29600);
nor UO_853 (O_853,N_20166,N_27997);
or UO_854 (O_854,N_22702,N_26552);
and UO_855 (O_855,N_20485,N_29655);
and UO_856 (O_856,N_28570,N_28375);
nand UO_857 (O_857,N_22169,N_24230);
and UO_858 (O_858,N_26331,N_23478);
or UO_859 (O_859,N_23518,N_27020);
and UO_860 (O_860,N_29896,N_26717);
and UO_861 (O_861,N_24792,N_27364);
nor UO_862 (O_862,N_20889,N_21694);
and UO_863 (O_863,N_20274,N_25579);
nor UO_864 (O_864,N_20560,N_25105);
nor UO_865 (O_865,N_21065,N_24015);
nor UO_866 (O_866,N_20299,N_22747);
or UO_867 (O_867,N_22392,N_23574);
nor UO_868 (O_868,N_20594,N_27427);
nor UO_869 (O_869,N_21453,N_20461);
or UO_870 (O_870,N_25382,N_22492);
nor UO_871 (O_871,N_22457,N_26672);
nand UO_872 (O_872,N_20698,N_21522);
and UO_873 (O_873,N_22878,N_28399);
nor UO_874 (O_874,N_21668,N_21606);
and UO_875 (O_875,N_20716,N_20023);
and UO_876 (O_876,N_20283,N_28446);
nand UO_877 (O_877,N_23857,N_22093);
nor UO_878 (O_878,N_20574,N_26289);
nand UO_879 (O_879,N_28796,N_27912);
nand UO_880 (O_880,N_27088,N_28634);
and UO_881 (O_881,N_27751,N_25583);
and UO_882 (O_882,N_25285,N_25654);
nand UO_883 (O_883,N_28066,N_26875);
and UO_884 (O_884,N_20260,N_20572);
nand UO_885 (O_885,N_24596,N_27539);
nor UO_886 (O_886,N_23531,N_29877);
nor UO_887 (O_887,N_22908,N_25665);
nand UO_888 (O_888,N_20143,N_24687);
nor UO_889 (O_889,N_23150,N_29954);
or UO_890 (O_890,N_27160,N_22354);
and UO_891 (O_891,N_26517,N_25022);
or UO_892 (O_892,N_29214,N_27311);
and UO_893 (O_893,N_28970,N_22746);
and UO_894 (O_894,N_25245,N_20027);
or UO_895 (O_895,N_20730,N_24176);
nor UO_896 (O_896,N_20208,N_23006);
or UO_897 (O_897,N_28662,N_20807);
and UO_898 (O_898,N_27329,N_23161);
nor UO_899 (O_899,N_29520,N_21432);
and UO_900 (O_900,N_20147,N_25153);
nand UO_901 (O_901,N_21371,N_27666);
and UO_902 (O_902,N_28094,N_24779);
or UO_903 (O_903,N_27187,N_21066);
nand UO_904 (O_904,N_24020,N_26458);
and UO_905 (O_905,N_21813,N_25619);
and UO_906 (O_906,N_27414,N_29400);
or UO_907 (O_907,N_27684,N_27608);
nor UO_908 (O_908,N_28497,N_27728);
and UO_909 (O_909,N_22453,N_25438);
nor UO_910 (O_910,N_27138,N_27383);
and UO_911 (O_911,N_29345,N_28949);
nand UO_912 (O_912,N_23187,N_23176);
nor UO_913 (O_913,N_25260,N_28454);
or UO_914 (O_914,N_28665,N_23392);
nand UO_915 (O_915,N_23309,N_25165);
nand UO_916 (O_916,N_21897,N_23397);
and UO_917 (O_917,N_27050,N_24270);
nor UO_918 (O_918,N_20107,N_29384);
nand UO_919 (O_919,N_25935,N_22545);
nor UO_920 (O_920,N_21934,N_26044);
nor UO_921 (O_921,N_24853,N_26097);
nor UO_922 (O_922,N_26727,N_22723);
nand UO_923 (O_923,N_23048,N_26246);
xor UO_924 (O_924,N_24975,N_22181);
nand UO_925 (O_925,N_27582,N_23050);
nor UO_926 (O_926,N_23055,N_26999);
and UO_927 (O_927,N_28196,N_23559);
or UO_928 (O_928,N_22736,N_20180);
or UO_929 (O_929,N_24767,N_24092);
nand UO_930 (O_930,N_22217,N_23390);
nor UO_931 (O_931,N_29360,N_24654);
and UO_932 (O_932,N_26745,N_28623);
nand UO_933 (O_933,N_24800,N_29046);
nor UO_934 (O_934,N_24433,N_21894);
and UO_935 (O_935,N_21647,N_20265);
nor UO_936 (O_936,N_22361,N_24289);
or UO_937 (O_937,N_25961,N_20021);
and UO_938 (O_938,N_24960,N_27380);
nor UO_939 (O_939,N_23025,N_22602);
nor UO_940 (O_940,N_20924,N_22950);
and UO_941 (O_941,N_20056,N_20878);
or UO_942 (O_942,N_20881,N_27706);
nand UO_943 (O_943,N_26374,N_23721);
and UO_944 (O_944,N_27055,N_21112);
or UO_945 (O_945,N_25793,N_29680);
nand UO_946 (O_946,N_27628,N_20546);
nand UO_947 (O_947,N_24953,N_27146);
nand UO_948 (O_948,N_24002,N_29730);
or UO_949 (O_949,N_22592,N_26575);
and UO_950 (O_950,N_26071,N_23584);
nand UO_951 (O_951,N_22609,N_23041);
nand UO_952 (O_952,N_20045,N_26726);
nand UO_953 (O_953,N_21266,N_24513);
or UO_954 (O_954,N_24987,N_21200);
or UO_955 (O_955,N_25189,N_24764);
nor UO_956 (O_956,N_20502,N_25881);
or UO_957 (O_957,N_29761,N_28788);
or UO_958 (O_958,N_20377,N_21688);
and UO_959 (O_959,N_21910,N_22664);
or UO_960 (O_960,N_28947,N_28943);
nor UO_961 (O_961,N_23491,N_21480);
nand UO_962 (O_962,N_26145,N_24233);
or UO_963 (O_963,N_28895,N_29953);
nor UO_964 (O_964,N_26549,N_29622);
nand UO_965 (O_965,N_29068,N_25851);
nand UO_966 (O_966,N_26377,N_23404);
nand UO_967 (O_967,N_24462,N_29281);
nor UO_968 (O_968,N_21497,N_24573);
nor UO_969 (O_969,N_24530,N_26151);
xnor UO_970 (O_970,N_23886,N_21962);
and UO_971 (O_971,N_21286,N_26003);
nor UO_972 (O_972,N_28166,N_24276);
nand UO_973 (O_973,N_20512,N_21290);
nor UO_974 (O_974,N_27349,N_23914);
nand UO_975 (O_975,N_28554,N_20448);
and UO_976 (O_976,N_25029,N_21375);
nand UO_977 (O_977,N_26828,N_21878);
or UO_978 (O_978,N_22645,N_25505);
nand UO_979 (O_979,N_22036,N_28092);
nand UO_980 (O_980,N_24165,N_28794);
and UO_981 (O_981,N_26209,N_28271);
or UO_982 (O_982,N_27371,N_20371);
and UO_983 (O_983,N_25162,N_25012);
or UO_984 (O_984,N_20220,N_29222);
or UO_985 (O_985,N_25732,N_29548);
and UO_986 (O_986,N_28923,N_27639);
nor UO_987 (O_987,N_22095,N_20261);
or UO_988 (O_988,N_23842,N_24908);
nand UO_989 (O_989,N_27387,N_28753);
nand UO_990 (O_990,N_21955,N_20849);
or UO_991 (O_991,N_20052,N_24669);
nand UO_992 (O_992,N_23328,N_24098);
nand UO_993 (O_993,N_22787,N_27637);
nor UO_994 (O_994,N_29736,N_27171);
or UO_995 (O_995,N_26710,N_22916);
and UO_996 (O_996,N_24734,N_29710);
and UO_997 (O_997,N_27353,N_20604);
nand UO_998 (O_998,N_24603,N_20991);
and UO_999 (O_999,N_28644,N_20339);
and UO_1000 (O_1000,N_27919,N_29978);
nand UO_1001 (O_1001,N_23612,N_29646);
and UO_1002 (O_1002,N_29209,N_29788);
nor UO_1003 (O_1003,N_28112,N_23059);
nand UO_1004 (O_1004,N_29871,N_24063);
nor UO_1005 (O_1005,N_26650,N_24686);
nor UO_1006 (O_1006,N_25471,N_24473);
or UO_1007 (O_1007,N_24282,N_20108);
or UO_1008 (O_1008,N_27218,N_29048);
nor UO_1009 (O_1009,N_28689,N_26046);
nor UO_1010 (O_1010,N_28069,N_25184);
nand UO_1011 (O_1011,N_28956,N_20162);
nor UO_1012 (O_1012,N_26390,N_22652);
or UO_1013 (O_1013,N_24377,N_28792);
or UO_1014 (O_1014,N_29696,N_26799);
nand UO_1015 (O_1015,N_29837,N_29661);
or UO_1016 (O_1016,N_24926,N_23524);
nand UO_1017 (O_1017,N_21249,N_22065);
and UO_1018 (O_1018,N_20022,N_20359);
nand UO_1019 (O_1019,N_22051,N_21042);
nor UO_1020 (O_1020,N_25385,N_20160);
or UO_1021 (O_1021,N_20091,N_27282);
nand UO_1022 (O_1022,N_23673,N_25416);
nor UO_1023 (O_1023,N_26567,N_23504);
nand UO_1024 (O_1024,N_27446,N_24700);
or UO_1025 (O_1025,N_29666,N_25307);
nand UO_1026 (O_1026,N_20965,N_29573);
or UO_1027 (O_1027,N_24896,N_25019);
nor UO_1028 (O_1028,N_20481,N_26996);
nand UO_1029 (O_1029,N_27204,N_22800);
or UO_1030 (O_1030,N_23760,N_26226);
or UO_1031 (O_1031,N_26784,N_20657);
nand UO_1032 (O_1032,N_27991,N_27372);
or UO_1033 (O_1033,N_26338,N_29174);
and UO_1034 (O_1034,N_27888,N_28876);
and UO_1035 (O_1035,N_24843,N_20929);
nand UO_1036 (O_1036,N_24171,N_21109);
nand UO_1037 (O_1037,N_27430,N_28672);
nor UO_1038 (O_1038,N_21784,N_26092);
nand UO_1039 (O_1039,N_29672,N_29045);
and UO_1040 (O_1040,N_25801,N_25633);
nand UO_1041 (O_1041,N_21049,N_20691);
nor UO_1042 (O_1042,N_22692,N_26312);
nor UO_1043 (O_1043,N_28038,N_22663);
and UO_1044 (O_1044,N_24929,N_22949);
nor UO_1045 (O_1045,N_23684,N_21697);
nand UO_1046 (O_1046,N_23680,N_20608);
and UO_1047 (O_1047,N_25311,N_28888);
and UO_1048 (O_1048,N_24156,N_25689);
nand UO_1049 (O_1049,N_28785,N_21207);
and UO_1050 (O_1050,N_21194,N_27864);
or UO_1051 (O_1051,N_26401,N_20222);
nor UO_1052 (O_1052,N_22435,N_20577);
nand UO_1053 (O_1053,N_26170,N_23011);
nand UO_1054 (O_1054,N_26895,N_29639);
nor UO_1055 (O_1055,N_22228,N_20810);
nand UO_1056 (O_1056,N_28463,N_24047);
and UO_1057 (O_1057,N_21341,N_25404);
and UO_1058 (O_1058,N_21916,N_26323);
or UO_1059 (O_1059,N_26586,N_23790);
or UO_1060 (O_1060,N_21944,N_28878);
nor UO_1061 (O_1061,N_23856,N_20226);
xor UO_1062 (O_1062,N_28808,N_20144);
nand UO_1063 (O_1063,N_21316,N_24013);
or UO_1064 (O_1064,N_24741,N_22655);
nor UO_1065 (O_1065,N_25970,N_20607);
or UO_1066 (O_1066,N_23063,N_27084);
nand UO_1067 (O_1067,N_26221,N_24260);
nor UO_1068 (O_1068,N_28945,N_26703);
nand UO_1069 (O_1069,N_29156,N_24959);
nor UO_1070 (O_1070,N_21413,N_21214);
and UO_1071 (O_1071,N_27975,N_23333);
or UO_1072 (O_1072,N_29226,N_22046);
or UO_1073 (O_1073,N_20490,N_23217);
or UO_1074 (O_1074,N_22789,N_24521);
or UO_1075 (O_1075,N_27701,N_20172);
and UO_1076 (O_1076,N_20303,N_25099);
nor UO_1077 (O_1077,N_25024,N_29162);
or UO_1078 (O_1078,N_21443,N_22352);
and UO_1079 (O_1079,N_27952,N_22004);
or UO_1080 (O_1080,N_27966,N_27512);
nor UO_1081 (O_1081,N_20947,N_26367);
nor UO_1082 (O_1082,N_22871,N_23977);
or UO_1083 (O_1083,N_22781,N_25800);
and UO_1084 (O_1084,N_23416,N_29444);
nor UO_1085 (O_1085,N_23409,N_22790);
nand UO_1086 (O_1086,N_28616,N_24995);
or UO_1087 (O_1087,N_20248,N_23512);
and UO_1088 (O_1088,N_27921,N_28858);
nor UO_1089 (O_1089,N_29739,N_25182);
and UO_1090 (O_1090,N_26684,N_22960);
nand UO_1091 (O_1091,N_24458,N_22027);
and UO_1092 (O_1092,N_22373,N_26682);
and UO_1093 (O_1093,N_23329,N_27507);
and UO_1094 (O_1094,N_28033,N_27566);
nor UO_1095 (O_1095,N_25513,N_20992);
or UO_1096 (O_1096,N_25172,N_20866);
nor UO_1097 (O_1097,N_24968,N_20774);
nand UO_1098 (O_1098,N_27720,N_20989);
and UO_1099 (O_1099,N_22445,N_21622);
or UO_1100 (O_1100,N_28203,N_22779);
or UO_1101 (O_1101,N_26776,N_24756);
nor UO_1102 (O_1102,N_23688,N_21610);
nor UO_1103 (O_1103,N_26593,N_20263);
nor UO_1104 (O_1104,N_24145,N_27223);
nand UO_1105 (O_1105,N_24403,N_26357);
nand UO_1106 (O_1106,N_22101,N_23155);
nand UO_1107 (O_1107,N_29136,N_28922);
nand UO_1108 (O_1108,N_24608,N_21072);
or UO_1109 (O_1109,N_25960,N_27636);
or UO_1110 (O_1110,N_29976,N_22945);
and UO_1111 (O_1111,N_25389,N_27297);
or UO_1112 (O_1112,N_26823,N_24859);
nor UO_1113 (O_1113,N_22265,N_24842);
nor UO_1114 (O_1114,N_26457,N_22884);
nand UO_1115 (O_1115,N_20298,N_23825);
or UO_1116 (O_1116,N_20839,N_26812);
or UO_1117 (O_1117,N_27134,N_27593);
and UO_1118 (O_1118,N_24580,N_23311);
and UO_1119 (O_1119,N_22382,N_22770);
and UO_1120 (O_1120,N_23274,N_26360);
nand UO_1121 (O_1121,N_26883,N_20395);
or UO_1122 (O_1122,N_21105,N_25061);
or UO_1123 (O_1123,N_24881,N_22849);
or UO_1124 (O_1124,N_21810,N_25408);
or UO_1125 (O_1125,N_27094,N_21618);
or UO_1126 (O_1126,N_22000,N_20846);
and UO_1127 (O_1127,N_23130,N_22823);
and UO_1128 (O_1128,N_26933,N_21580);
nand UO_1129 (O_1129,N_22301,N_23053);
nand UO_1130 (O_1130,N_29729,N_21904);
nand UO_1131 (O_1131,N_23032,N_25669);
nand UO_1132 (O_1132,N_29088,N_29853);
nand UO_1133 (O_1133,N_23372,N_22584);
and UO_1134 (O_1134,N_28122,N_29934);
and UO_1135 (O_1135,N_28521,N_29713);
and UO_1136 (O_1136,N_20908,N_29257);
nor UO_1137 (O_1137,N_26262,N_28019);
or UO_1138 (O_1138,N_27492,N_25065);
or UO_1139 (O_1139,N_22850,N_23174);
or UO_1140 (O_1140,N_23459,N_20157);
or UO_1141 (O_1141,N_25968,N_24698);
nor UO_1142 (O_1142,N_21199,N_27366);
or UO_1143 (O_1143,N_27756,N_24188);
nand UO_1144 (O_1144,N_27540,N_24451);
nor UO_1145 (O_1145,N_27243,N_20505);
nand UO_1146 (O_1146,N_25532,N_23561);
and UO_1147 (O_1147,N_22138,N_29775);
and UO_1148 (O_1148,N_22940,N_25467);
nand UO_1149 (O_1149,N_22614,N_28029);
nor UO_1150 (O_1150,N_25642,N_23606);
and UO_1151 (O_1151,N_26912,N_26673);
and UO_1152 (O_1152,N_25485,N_22389);
nand UO_1153 (O_1153,N_28977,N_27716);
nor UO_1154 (O_1154,N_21436,N_25630);
and UO_1155 (O_1155,N_22829,N_26084);
nor UO_1156 (O_1156,N_20123,N_22659);
and UO_1157 (O_1157,N_22029,N_22843);
and UO_1158 (O_1158,N_26619,N_23748);
nand UO_1159 (O_1159,N_25325,N_28084);
nand UO_1160 (O_1160,N_21046,N_23810);
nor UO_1161 (O_1161,N_28131,N_28948);
and UO_1162 (O_1162,N_21732,N_22582);
nand UO_1163 (O_1163,N_28500,N_20134);
nand UO_1164 (O_1164,N_26922,N_29176);
nand UO_1165 (O_1165,N_22345,N_28780);
and UO_1166 (O_1166,N_20637,N_24944);
nor UO_1167 (O_1167,N_23603,N_20369);
nand UO_1168 (O_1168,N_24694,N_28225);
and UO_1169 (O_1169,N_23136,N_23399);
nor UO_1170 (O_1170,N_20459,N_20346);
and UO_1171 (O_1171,N_23351,N_23919);
and UO_1172 (O_1172,N_29303,N_21699);
or UO_1173 (O_1173,N_20679,N_26194);
and UO_1174 (O_1174,N_26966,N_21553);
nand UO_1175 (O_1175,N_23144,N_28654);
and UO_1176 (O_1176,N_25839,N_26801);
and UO_1177 (O_1177,N_20873,N_27269);
xnor UO_1178 (O_1178,N_23381,N_29251);
nand UO_1179 (O_1179,N_21069,N_23965);
or UO_1180 (O_1180,N_28404,N_26410);
nand UO_1181 (O_1181,N_27224,N_22491);
or UO_1182 (O_1182,N_21358,N_22678);
nor UO_1183 (O_1183,N_27074,N_27429);
nor UO_1184 (O_1184,N_28690,N_29118);
nand UO_1185 (O_1185,N_29589,N_26452);
nand UO_1186 (O_1186,N_24828,N_23266);
nor UO_1187 (O_1187,N_20711,N_28213);
nor UO_1188 (O_1188,N_20901,N_24322);
nand UO_1189 (O_1189,N_29714,N_20006);
xor UO_1190 (O_1190,N_29852,N_23373);
and UO_1191 (O_1191,N_23717,N_21636);
and UO_1192 (O_1192,N_29803,N_20114);
and UO_1193 (O_1193,N_20444,N_26497);
nand UO_1194 (O_1194,N_21283,N_26328);
or UO_1195 (O_1195,N_28600,N_29923);
nand UO_1196 (O_1196,N_27235,N_29032);
and UO_1197 (O_1197,N_20046,N_28324);
nand UO_1198 (O_1198,N_23835,N_27626);
nor UO_1199 (O_1199,N_26017,N_24072);
nand UO_1200 (O_1200,N_27439,N_21990);
and UO_1201 (O_1201,N_23273,N_23541);
nand UO_1202 (O_1202,N_20399,N_29055);
and UO_1203 (O_1203,N_22295,N_22616);
nor UO_1204 (O_1204,N_21152,N_27161);
nand UO_1205 (O_1205,N_23792,N_20237);
nand UO_1206 (O_1206,N_23226,N_25221);
or UO_1207 (O_1207,N_23252,N_25303);
and UO_1208 (O_1208,N_23793,N_23215);
or UO_1209 (O_1209,N_20340,N_27623);
nor UO_1210 (O_1210,N_24331,N_27394);
or UO_1211 (O_1211,N_26235,N_22446);
nor UO_1212 (O_1212,N_25788,N_28458);
or UO_1213 (O_1213,N_23900,N_26663);
and UO_1214 (O_1214,N_24122,N_23664);
or UO_1215 (O_1215,N_22070,N_28893);
or UO_1216 (O_1216,N_25259,N_22466);
or UO_1217 (O_1217,N_26320,N_28243);
or UO_1218 (O_1218,N_24237,N_23068);
nor UO_1219 (O_1219,N_27262,N_22651);
nand UO_1220 (O_1220,N_23872,N_25840);
nand UO_1221 (O_1221,N_24342,N_28185);
nor UO_1222 (O_1222,N_25014,N_24586);
or UO_1223 (O_1223,N_27475,N_29318);
nor UO_1224 (O_1224,N_25846,N_26881);
nand UO_1225 (O_1225,N_21368,N_21734);
nor UO_1226 (O_1226,N_24562,N_22049);
nand UO_1227 (O_1227,N_22425,N_28258);
and UO_1228 (O_1228,N_21380,N_24673);
or UO_1229 (O_1229,N_21465,N_23824);
and UO_1230 (O_1230,N_28915,N_25484);
nor UO_1231 (O_1231,N_28279,N_25489);
or UO_1232 (O_1232,N_23807,N_25083);
nor UO_1233 (O_1233,N_24527,N_25133);
nor UO_1234 (O_1234,N_21490,N_22242);
nor UO_1235 (O_1235,N_23142,N_22646);
or UO_1236 (O_1236,N_28606,N_27800);
or UO_1237 (O_1237,N_25850,N_26788);
or UO_1238 (O_1238,N_25371,N_21748);
and UO_1239 (O_1239,N_25009,N_23418);
or UO_1240 (O_1240,N_21880,N_23839);
nor UO_1241 (O_1241,N_27827,N_22026);
nor UO_1242 (O_1242,N_26143,N_29793);
nand UO_1243 (O_1243,N_23220,N_20098);
and UO_1244 (O_1244,N_25696,N_22951);
nor UO_1245 (O_1245,N_27201,N_28999);
nor UO_1246 (O_1246,N_29511,N_29711);
or UO_1247 (O_1247,N_20062,N_22119);
nor UO_1248 (O_1248,N_25536,N_21485);
and UO_1249 (O_1249,N_23385,N_28642);
xnor UO_1250 (O_1250,N_24405,N_27808);
nand UO_1251 (O_1251,N_27851,N_29430);
or UO_1252 (O_1252,N_26154,N_26547);
nor UO_1253 (O_1253,N_23660,N_25909);
and UO_1254 (O_1254,N_25581,N_25043);
or UO_1255 (O_1255,N_22341,N_27707);
nand UO_1256 (O_1256,N_28917,N_29827);
nand UO_1257 (O_1257,N_23077,N_22901);
nand UO_1258 (O_1258,N_27753,N_27508);
nor UO_1259 (O_1259,N_21272,N_25391);
nand UO_1260 (O_1260,N_27806,N_24094);
nand UO_1261 (O_1261,N_24320,N_24048);
or UO_1262 (O_1262,N_21991,N_21367);
or UO_1263 (O_1263,N_27317,N_21068);
nor UO_1264 (O_1264,N_25256,N_29153);
nand UO_1265 (O_1265,N_29649,N_22084);
and UO_1266 (O_1266,N_29604,N_29995);
nand UO_1267 (O_1267,N_26035,N_24898);
and UO_1268 (O_1268,N_22079,N_20694);
nor UO_1269 (O_1269,N_21572,N_22836);
nand UO_1270 (O_1270,N_22193,N_27176);
or UO_1271 (O_1271,N_20602,N_24784);
or UO_1272 (O_1272,N_24749,N_24352);
nand UO_1273 (O_1273,N_26082,N_22639);
nand UO_1274 (O_1274,N_29258,N_20646);
and UO_1275 (O_1275,N_21750,N_28586);
or UO_1276 (O_1276,N_27790,N_27982);
nor UO_1277 (O_1277,N_22275,N_20386);
or UO_1278 (O_1278,N_25291,N_20964);
nand UO_1279 (O_1279,N_28847,N_21258);
or UO_1280 (O_1280,N_24794,N_29771);
nor UO_1281 (O_1281,N_27907,N_28153);
and UO_1282 (O_1282,N_27869,N_22197);
or UO_1283 (O_1283,N_25622,N_20355);
nand UO_1284 (O_1284,N_26368,N_27892);
and UO_1285 (O_1285,N_29644,N_20119);
and UO_1286 (O_1286,N_29945,N_26080);
or UO_1287 (O_1287,N_24466,N_22904);
and UO_1288 (O_1288,N_20982,N_27162);
nor UO_1289 (O_1289,N_20202,N_25441);
or UO_1290 (O_1290,N_26265,N_24934);
or UO_1291 (O_1291,N_24519,N_22221);
nor UO_1292 (O_1292,N_25679,N_24112);
or UO_1293 (O_1293,N_24295,N_24378);
nand UO_1294 (O_1294,N_26523,N_28088);
xnor UO_1295 (O_1295,N_22085,N_27604);
and UO_1296 (O_1296,N_22396,N_29797);
and UO_1297 (O_1297,N_29495,N_28205);
and UO_1298 (O_1298,N_20191,N_24297);
nand UO_1299 (O_1299,N_28841,N_28871);
nand UO_1300 (O_1300,N_24025,N_28583);
and UO_1301 (O_1301,N_27780,N_20720);
and UO_1302 (O_1302,N_22801,N_23956);
or UO_1303 (O_1303,N_27762,N_26825);
nor UO_1304 (O_1304,N_25695,N_22343);
and UO_1305 (O_1305,N_24871,N_25914);
or UO_1306 (O_1306,N_21311,N_28717);
and UO_1307 (O_1307,N_28068,N_25875);
or UO_1308 (O_1308,N_21406,N_29391);
or UO_1309 (O_1309,N_27818,N_26378);
and UO_1310 (O_1310,N_21050,N_25592);
nor UO_1311 (O_1311,N_24412,N_21924);
or UO_1312 (O_1312,N_26546,N_26042);
nand UO_1313 (O_1313,N_25745,N_29988);
and UO_1314 (O_1314,N_26364,N_20161);
and UO_1315 (O_1315,N_27894,N_26387);
or UO_1316 (O_1316,N_20131,N_29012);
or UO_1317 (O_1317,N_28056,N_24152);
and UO_1318 (O_1318,N_29419,N_23185);
nand UO_1319 (O_1319,N_25537,N_20420);
nor UO_1320 (O_1320,N_22604,N_23871);
or UO_1321 (O_1321,N_27562,N_20931);
nand UO_1322 (O_1322,N_20389,N_28234);
or UO_1323 (O_1323,N_29756,N_26466);
and UO_1324 (O_1324,N_26520,N_27140);
nor UO_1325 (O_1325,N_20071,N_26463);
nand UO_1326 (O_1326,N_22473,N_22890);
or UO_1327 (O_1327,N_21080,N_29781);
or UO_1328 (O_1328,N_22183,N_21142);
or UO_1329 (O_1329,N_24628,N_20864);
and UO_1330 (O_1330,N_29527,N_26498);
and UO_1331 (O_1331,N_29902,N_28389);
nor UO_1332 (O_1332,N_29681,N_27641);
and UO_1333 (O_1333,N_28143,N_25298);
nor UO_1334 (O_1334,N_28901,N_23801);
or UO_1335 (O_1335,N_26232,N_22648);
nand UO_1336 (O_1336,N_26655,N_29328);
nand UO_1337 (O_1337,N_20465,N_20514);
nand UO_1338 (O_1338,N_23181,N_21255);
nand UO_1339 (O_1339,N_23628,N_28260);
and UO_1340 (O_1340,N_26928,N_28332);
and UO_1341 (O_1341,N_29550,N_25777);
nor UO_1342 (O_1342,N_28012,N_25769);
or UO_1343 (O_1343,N_29037,N_27482);
or UO_1344 (O_1344,N_27960,N_29474);
and UO_1345 (O_1345,N_24664,N_25674);
and UO_1346 (O_1346,N_28604,N_21034);
and UO_1347 (O_1347,N_28712,N_22443);
nand UO_1348 (O_1348,N_27746,N_22411);
nor UO_1349 (O_1349,N_27821,N_25733);
or UO_1350 (O_1350,N_22739,N_24044);
nand UO_1351 (O_1351,N_22891,N_27645);
nor UO_1352 (O_1352,N_24941,N_22485);
and UO_1353 (O_1353,N_20516,N_23927);
or UO_1354 (O_1354,N_22588,N_23873);
nor UO_1355 (O_1355,N_22761,N_24390);
and UO_1356 (O_1356,N_28734,N_20545);
nor UO_1357 (O_1357,N_24814,N_26083);
or UO_1358 (O_1358,N_20210,N_25010);
and UO_1359 (O_1359,N_28952,N_23129);
nand UO_1360 (O_1360,N_22157,N_20615);
or UO_1361 (O_1361,N_29363,N_22165);
and UO_1362 (O_1362,N_27523,N_21956);
nor UO_1363 (O_1363,N_24776,N_23765);
nand UO_1364 (O_1364,N_23985,N_28292);
nor UO_1365 (O_1365,N_26709,N_21481);
nor UO_1366 (O_1366,N_25414,N_25904);
nor UO_1367 (O_1367,N_22421,N_25401);
and UO_1368 (O_1368,N_25211,N_26904);
or UO_1369 (O_1369,N_23879,N_23087);
nand UO_1370 (O_1370,N_26179,N_23987);
or UO_1371 (O_1371,N_25956,N_27186);
or UO_1372 (O_1372,N_28141,N_26379);
and UO_1373 (O_1373,N_22798,N_28543);
and UO_1374 (O_1374,N_28211,N_29203);
nor UO_1375 (O_1375,N_29081,N_22680);
nand UO_1376 (O_1376,N_27319,N_22786);
or UO_1377 (O_1377,N_22830,N_25296);
nor UO_1378 (O_1378,N_20522,N_23149);
or UO_1379 (O_1379,N_25356,N_25072);
nor UO_1380 (O_1380,N_25527,N_26127);
nor UO_1381 (O_1381,N_21660,N_24275);
or UO_1382 (O_1382,N_27231,N_22820);
nand UO_1383 (O_1383,N_21349,N_26832);
nor UO_1384 (O_1384,N_20825,N_28837);
nor UO_1385 (O_1385,N_22110,N_29667);
and UO_1386 (O_1386,N_25653,N_24470);
nand UO_1387 (O_1387,N_26948,N_29817);
or UO_1388 (O_1388,N_23583,N_26569);
nor UO_1389 (O_1389,N_27158,N_28696);
nand UO_1390 (O_1390,N_21504,N_29967);
nor UO_1391 (O_1391,N_21988,N_22141);
and UO_1392 (O_1392,N_25046,N_27880);
nand UO_1393 (O_1393,N_27889,N_24763);
nor UO_1394 (O_1394,N_22844,N_29507);
nand UO_1395 (O_1395,N_22336,N_21792);
and UO_1396 (O_1396,N_28625,N_26635);
nor UO_1397 (O_1397,N_21595,N_26270);
or UO_1398 (O_1398,N_20268,N_24489);
or UO_1399 (O_1399,N_24630,N_26910);
nand UO_1400 (O_1400,N_29067,N_27787);
nand UO_1401 (O_1401,N_20942,N_29709);
nand UO_1402 (O_1402,N_24241,N_26427);
or UO_1403 (O_1403,N_22865,N_27781);
nor UO_1404 (O_1404,N_28806,N_28371);
or UO_1405 (O_1405,N_25347,N_22493);
nor UO_1406 (O_1406,N_23314,N_29343);
and UO_1407 (O_1407,N_21252,N_23638);
and UO_1408 (O_1408,N_22854,N_26306);
or UO_1409 (O_1409,N_20611,N_24633);
nand UO_1410 (O_1410,N_29376,N_29121);
nand UO_1411 (O_1411,N_25871,N_27943);
nand UO_1412 (O_1412,N_20738,N_27436);
and UO_1413 (O_1413,N_20140,N_28544);
nand UO_1414 (O_1414,N_21166,N_24796);
nor UO_1415 (O_1415,N_28961,N_28933);
nand UO_1416 (O_1416,N_23042,N_25779);
and UO_1417 (O_1417,N_24028,N_28251);
nor UO_1418 (O_1418,N_26201,N_23075);
xnor UO_1419 (O_1419,N_28510,N_24857);
and UO_1420 (O_1420,N_28765,N_25857);
and UO_1421 (O_1421,N_29467,N_21720);
and UO_1422 (O_1422,N_20447,N_28540);
nand UO_1423 (O_1423,N_22982,N_28162);
nor UO_1424 (O_1424,N_29634,N_24076);
and UO_1425 (O_1425,N_28428,N_23548);
or UO_1426 (O_1426,N_24594,N_26291);
nand UO_1427 (O_1427,N_27817,N_29207);
nand UO_1428 (O_1428,N_23912,N_26073);
nand UO_1429 (O_1429,N_23630,N_25450);
or UO_1430 (O_1430,N_27624,N_21345);
and UO_1431 (O_1431,N_27310,N_28285);
and UO_1432 (O_1432,N_29024,N_26542);
and UO_1433 (O_1433,N_22944,N_26475);
nand UO_1434 (O_1434,N_23747,N_25903);
and UO_1435 (O_1435,N_24169,N_23196);
nor UO_1436 (O_1436,N_23611,N_24372);
nand UO_1437 (O_1437,N_24775,N_29966);
or UO_1438 (O_1438,N_26565,N_20897);
or UO_1439 (O_1439,N_24082,N_27421);
xor UO_1440 (O_1440,N_23207,N_20063);
nor UO_1441 (O_1441,N_27957,N_24434);
nand UO_1442 (O_1442,N_28776,N_24830);
nor UO_1443 (O_1443,N_29232,N_29728);
and UO_1444 (O_1444,N_27979,N_23566);
nand UO_1445 (O_1445,N_20456,N_28218);
and UO_1446 (O_1446,N_29043,N_20314);
or UO_1447 (O_1447,N_21848,N_27598);
nand UO_1448 (O_1448,N_25715,N_21044);
nand UO_1449 (O_1449,N_21456,N_22405);
and UO_1450 (O_1450,N_27612,N_27316);
nand UO_1451 (O_1451,N_21048,N_22538);
nand UO_1452 (O_1452,N_29984,N_28957);
and UO_1453 (O_1453,N_29295,N_21451);
nor UO_1454 (O_1454,N_27530,N_20177);
or UO_1455 (O_1455,N_26851,N_29937);
nor UO_1456 (O_1456,N_25495,N_22763);
nand UO_1457 (O_1457,N_28627,N_23109);
and UO_1458 (O_1458,N_26026,N_25770);
nand UO_1459 (O_1459,N_27816,N_21295);
nand UO_1460 (O_1460,N_27360,N_24089);
nand UO_1461 (O_1461,N_24475,N_28240);
nand UO_1462 (O_1462,N_28422,N_24374);
and UO_1463 (O_1463,N_25280,N_22615);
nor UO_1464 (O_1464,N_29755,N_20121);
or UO_1465 (O_1465,N_27463,N_27257);
nand UO_1466 (O_1466,N_27859,N_20979);
or UO_1467 (O_1467,N_24215,N_21675);
or UO_1468 (O_1468,N_22724,N_27522);
or UO_1469 (O_1469,N_25831,N_26057);
nand UO_1470 (O_1470,N_28574,N_29029);
or UO_1471 (O_1471,N_26667,N_29950);
or UO_1472 (O_1472,N_20030,N_25130);
and UO_1473 (O_1473,N_23033,N_29021);
and UO_1474 (O_1474,N_20672,N_24738);
nand UO_1475 (O_1475,N_27148,N_20300);
nor UO_1476 (O_1476,N_28687,N_23143);
nand UO_1477 (O_1477,N_29734,N_22793);
and UO_1478 (O_1478,N_26824,N_29547);
and UO_1479 (O_1479,N_25986,N_22432);
and UO_1480 (O_1480,N_24005,N_22923);
and UO_1481 (O_1481,N_21086,N_26627);
or UO_1482 (O_1482,N_24873,N_22459);
nor UO_1483 (O_1483,N_25934,N_22324);
or UO_1484 (O_1484,N_20687,N_27346);
nor UO_1485 (O_1485,N_21728,N_20037);
or UO_1486 (O_1486,N_25969,N_28709);
or UO_1487 (O_1487,N_28148,N_27491);
or UO_1488 (O_1488,N_25998,N_22199);
or UO_1489 (O_1489,N_29341,N_21652);
or UO_1490 (O_1490,N_21726,N_26732);
or UO_1491 (O_1491,N_20370,N_25050);
and UO_1492 (O_1492,N_28411,N_23949);
and UO_1493 (O_1493,N_25603,N_22628);
nor UO_1494 (O_1494,N_26195,N_28814);
and UO_1495 (O_1495,N_21160,N_27409);
nor UO_1496 (O_1496,N_23758,N_23198);
nand UO_1497 (O_1497,N_27681,N_26476);
and UO_1498 (O_1498,N_25873,N_28097);
nor UO_1499 (O_1499,N_25584,N_29086);
nand UO_1500 (O_1500,N_26366,N_20893);
nor UO_1501 (O_1501,N_22898,N_25772);
or UO_1502 (O_1502,N_21430,N_29669);
or UO_1503 (O_1503,N_23334,N_27939);
or UO_1504 (O_1504,N_21446,N_26011);
nor UO_1505 (O_1505,N_25856,N_25787);
and UO_1506 (O_1506,N_24358,N_28828);
or UO_1507 (O_1507,N_29385,N_20313);
nand UO_1508 (O_1508,N_20693,N_29746);
and UO_1509 (O_1509,N_29451,N_23652);
and UO_1510 (O_1510,N_20827,N_27307);
and UO_1511 (O_1511,N_27823,N_27510);
and UO_1512 (O_1512,N_22532,N_27328);
nor UO_1513 (O_1513,N_21678,N_25549);
nor UO_1514 (O_1514,N_25210,N_27783);
nor UO_1515 (O_1515,N_21889,N_23413);
or UO_1516 (O_1516,N_21054,N_29245);
nor UO_1517 (O_1517,N_26482,N_22121);
or UO_1518 (O_1518,N_23100,N_22076);
nor UO_1519 (O_1519,N_24491,N_25915);
or UO_1520 (O_1520,N_22460,N_27141);
or UO_1521 (O_1521,N_20922,N_22246);
and UO_1522 (O_1522,N_29224,N_22855);
or UO_1523 (O_1523,N_26985,N_28496);
and UO_1524 (O_1524,N_29504,N_21854);
or UO_1525 (O_1525,N_21807,N_22876);
and UO_1526 (O_1526,N_20500,N_21229);
nand UO_1527 (O_1527,N_21254,N_27327);
and UO_1528 (O_1528,N_24882,N_27875);
nand UO_1529 (O_1529,N_26601,N_24635);
nor UO_1530 (O_1530,N_23620,N_21738);
nand UO_1531 (O_1531,N_23599,N_21448);
and UO_1532 (O_1532,N_21387,N_24254);
nand UO_1533 (O_1533,N_27056,N_23361);
nand UO_1534 (O_1534,N_27498,N_27180);
nand UO_1535 (O_1535,N_27029,N_22123);
and UO_1536 (O_1536,N_23821,N_29403);
nor UO_1537 (O_1537,N_25397,N_21808);
xnor UO_1538 (O_1538,N_24688,N_24343);
nor UO_1539 (O_1539,N_28585,N_24350);
nand UO_1540 (O_1540,N_22983,N_21470);
nor UO_1541 (O_1541,N_23393,N_21628);
or UO_1542 (O_1542,N_25657,N_20542);
nand UO_1543 (O_1543,N_24327,N_26681);
and UO_1544 (O_1544,N_29272,N_29722);
nand UO_1545 (O_1545,N_27195,N_29261);
and UO_1546 (O_1546,N_28008,N_23909);
or UO_1547 (O_1547,N_29313,N_28447);
or UO_1548 (O_1548,N_22458,N_25655);
nor UO_1549 (O_1549,N_21541,N_20872);
or UO_1550 (O_1550,N_23362,N_24354);
or UO_1551 (O_1551,N_29325,N_29816);
and UO_1552 (O_1552,N_20489,N_22155);
nor UO_1553 (O_1553,N_28413,N_22206);
or UO_1554 (O_1554,N_29880,N_20419);
and UO_1555 (O_1555,N_25333,N_26821);
and UO_1556 (O_1556,N_27589,N_29028);
nand UO_1557 (O_1557,N_22260,N_22060);
or UO_1558 (O_1558,N_24179,N_26531);
nor UO_1559 (O_1559,N_23658,N_20640);
nand UO_1560 (O_1560,N_26171,N_21773);
or UO_1561 (O_1561,N_23167,N_28353);
nand UO_1562 (O_1562,N_20181,N_24065);
or UO_1563 (O_1563,N_21816,N_28532);
xor UO_1564 (O_1564,N_27771,N_24235);
nand UO_1565 (O_1565,N_29353,N_20256);
or UO_1566 (O_1566,N_24329,N_22212);
nor UO_1567 (O_1567,N_29185,N_21589);
and UO_1568 (O_1568,N_26314,N_26431);
or UO_1569 (O_1569,N_22062,N_25452);
or UO_1570 (O_1570,N_27620,N_21385);
or UO_1571 (O_1571,N_24910,N_29568);
nor UO_1572 (O_1572,N_23429,N_29610);
and UO_1573 (O_1573,N_21461,N_27899);
nor UO_1574 (O_1574,N_26987,N_25025);
nand UO_1575 (O_1575,N_28784,N_20526);
nand UO_1576 (O_1576,N_20078,N_24532);
nand UO_1577 (O_1577,N_23152,N_22821);
and UO_1578 (O_1578,N_28072,N_23192);
nand UO_1579 (O_1579,N_23751,N_23405);
nor UO_1580 (O_1580,N_23526,N_26344);
nand UO_1581 (O_1581,N_29790,N_26758);
nand UO_1582 (O_1582,N_26858,N_26137);
and UO_1583 (O_1583,N_26005,N_27544);
or UO_1584 (O_1584,N_23131,N_26428);
nand UO_1585 (O_1585,N_22147,N_23021);
or UO_1586 (O_1586,N_22753,N_26184);
nand UO_1587 (O_1587,N_22699,N_25282);
or UO_1588 (O_1588,N_23338,N_24143);
or UO_1589 (O_1589,N_25003,N_24088);
and UO_1590 (O_1590,N_27849,N_26442);
xnor UO_1591 (O_1591,N_29855,N_25731);
and UO_1592 (O_1592,N_29594,N_26762);
nand UO_1593 (O_1593,N_23247,N_26336);
nor UO_1594 (O_1594,N_21936,N_23236);
and UO_1595 (O_1595,N_26271,N_22194);
and UO_1596 (O_1596,N_28418,N_20765);
xor UO_1597 (O_1597,N_26206,N_21469);
and UO_1598 (O_1598,N_28789,N_20329);
and UO_1599 (O_1599,N_27936,N_20622);
nand UO_1600 (O_1600,N_25242,N_22562);
or UO_1601 (O_1601,N_22640,N_25597);
or UO_1602 (O_1602,N_21028,N_25312);
nand UO_1603 (O_1603,N_25106,N_27193);
nand UO_1604 (O_1604,N_25933,N_26863);
nor UO_1605 (O_1605,N_20292,N_21360);
nor UO_1606 (O_1606,N_29509,N_29723);
nand UO_1607 (O_1607,N_20076,N_24425);
or UO_1608 (O_1608,N_29432,N_22979);
nor UO_1609 (O_1609,N_21232,N_29849);
and UO_1610 (O_1610,N_25059,N_29038);
nor UO_1611 (O_1611,N_28605,N_24797);
and UO_1612 (O_1612,N_21764,N_21113);
nor UO_1613 (O_1613,N_21978,N_29515);
or UO_1614 (O_1614,N_27113,N_21971);
nor UO_1615 (O_1615,N_22750,N_28971);
nor UO_1616 (O_1616,N_22932,N_29514);
or UO_1617 (O_1617,N_21601,N_23320);
nand UO_1618 (O_1618,N_26304,N_22417);
or UO_1619 (O_1619,N_22480,N_27659);
nand UO_1620 (O_1620,N_27206,N_21970);
nor UO_1621 (O_1621,N_29996,N_29534);
or UO_1622 (O_1622,N_26492,N_28085);
nand UO_1623 (O_1623,N_21015,N_23071);
or UO_1624 (O_1624,N_27927,N_26576);
and UO_1625 (O_1625,N_28367,N_21129);
nor UO_1626 (O_1626,N_28345,N_26502);
nand UO_1627 (O_1627,N_25947,N_22478);
nor UO_1628 (O_1628,N_26088,N_23148);
and UO_1629 (O_1629,N_26625,N_23587);
nor UO_1630 (O_1630,N_24214,N_28280);
and UO_1631 (O_1631,N_27739,N_21098);
and UO_1632 (O_1632,N_28890,N_25763);
or UO_1633 (O_1633,N_24974,N_28172);
nand UO_1634 (O_1634,N_26049,N_28903);
nand UO_1635 (O_1635,N_20638,N_20269);
and UO_1636 (O_1636,N_25813,N_25380);
nor UO_1637 (O_1637,N_26070,N_29897);
nor UO_1638 (O_1638,N_25449,N_27886);
nor UO_1639 (O_1639,N_26965,N_26462);
xor UO_1640 (O_1640,N_29247,N_25860);
nand UO_1641 (O_1641,N_24808,N_23922);
or UO_1642 (O_1642,N_28748,N_25104);
nand UO_1643 (O_1643,N_29806,N_21313);
nor UO_1644 (O_1644,N_28777,N_27609);
nand UO_1645 (O_1645,N_24315,N_23744);
or UO_1646 (O_1646,N_29439,N_21267);
nor UO_1647 (O_1647,N_27862,N_21475);
nor UO_1648 (O_1648,N_29359,N_22529);
nor UO_1649 (O_1649,N_25476,N_22826);
nor UO_1650 (O_1650,N_28410,N_28007);
nor UO_1651 (O_1651,N_28844,N_22278);
or UO_1652 (O_1652,N_22822,N_22512);
nand UO_1653 (O_1653,N_20105,N_28048);
and UO_1654 (O_1654,N_23410,N_27680);
nor UO_1655 (O_1655,N_28981,N_29642);
or UO_1656 (O_1656,N_25912,N_26878);
nand UO_1657 (O_1657,N_24388,N_20949);
nand UO_1658 (O_1658,N_28666,N_27920);
and UO_1659 (O_1659,N_20249,N_29101);
or UO_1660 (O_1660,N_20293,N_25073);
or UO_1661 (O_1661,N_28481,N_24236);
and UO_1662 (O_1662,N_22694,N_21626);
and UO_1663 (O_1663,N_28584,N_25568);
nor UO_1664 (O_1664,N_27873,N_26793);
or UO_1665 (O_1665,N_21890,N_28655);
nand UO_1666 (O_1666,N_23049,N_29955);
nor UO_1667 (O_1667,N_27399,N_27689);
and UO_1668 (O_1668,N_21805,N_22688);
or UO_1669 (O_1669,N_26443,N_27188);
and UO_1670 (O_1670,N_23138,N_25068);
and UO_1671 (O_1671,N_26295,N_27611);
and UO_1672 (O_1672,N_24050,N_23319);
nand UO_1673 (O_1673,N_20291,N_23632);
nand UO_1674 (O_1674,N_29195,N_27916);
nor UO_1675 (O_1675,N_27538,N_20136);
or UO_1676 (O_1676,N_27909,N_22802);
or UO_1677 (O_1677,N_25690,N_28095);
or UO_1678 (O_1678,N_23520,N_28608);
and UO_1679 (O_1679,N_26233,N_25007);
or UO_1680 (O_1680,N_27881,N_26763);
nor UO_1681 (O_1681,N_20540,N_23400);
nor UO_1682 (O_1682,N_20296,N_25041);
or UO_1683 (O_1683,N_21793,N_21369);
nor UO_1684 (O_1684,N_25144,N_25919);
or UO_1685 (O_1685,N_28245,N_28237);
or UO_1686 (O_1686,N_23350,N_24095);
or UO_1687 (O_1687,N_24502,N_25834);
xor UO_1688 (O_1688,N_23718,N_20704);
nand UO_1689 (O_1689,N_24079,N_23517);
nor UO_1690 (O_1690,N_23671,N_28244);
or UO_1691 (O_1691,N_22033,N_21064);
or UO_1692 (O_1692,N_29865,N_29096);
nor UO_1693 (O_1693,N_29047,N_26775);
nand UO_1694 (O_1694,N_23579,N_28098);
or UO_1695 (O_1695,N_23292,N_21996);
or UO_1696 (O_1696,N_28381,N_21121);
nor UO_1697 (O_1697,N_26405,N_23183);
nor UO_1698 (O_1698,N_21384,N_22150);
nor UO_1699 (O_1699,N_20378,N_28622);
nand UO_1700 (O_1700,N_23367,N_27082);
nand UO_1701 (O_1701,N_28439,N_25398);
nor UO_1702 (O_1702,N_27630,N_22475);
nor UO_1703 (O_1703,N_24485,N_24665);
nand UO_1704 (O_1704,N_25496,N_29609);
nand UO_1705 (O_1705,N_23554,N_21712);
nand UO_1706 (O_1706,N_21201,N_24284);
nand UO_1707 (O_1707,N_21603,N_20446);
and UO_1708 (O_1708,N_21838,N_26656);
nand UO_1709 (O_1709,N_23509,N_24777);
nor UO_1710 (O_1710,N_25465,N_20800);
nand UO_1711 (O_1711,N_23415,N_21447);
nor UO_1712 (O_1712,N_29804,N_27343);
or UO_1713 (O_1713,N_20016,N_21901);
or UO_1714 (O_1714,N_23736,N_26081);
or UO_1715 (O_1715,N_20858,N_21763);
and UO_1716 (O_1716,N_20803,N_27596);
nand UO_1717 (O_1717,N_28911,N_22462);
or UO_1718 (O_1718,N_22031,N_22126);
and UO_1719 (O_1719,N_21741,N_23592);
nand UO_1720 (O_1720,N_26909,N_24951);
nand UO_1721 (O_1721,N_28125,N_21495);
nor UO_1722 (O_1722,N_29914,N_26131);
nor UO_1723 (O_1723,N_22856,N_21739);
or UO_1724 (O_1724,N_27200,N_29491);
nand UO_1725 (O_1725,N_23781,N_26742);
xnor UO_1726 (O_1726,N_27142,N_26636);
or UO_1727 (O_1727,N_27393,N_23438);
and UO_1728 (O_1728,N_26869,N_26382);
nor UO_1729 (O_1729,N_21204,N_23219);
nand UO_1730 (O_1730,N_24903,N_22591);
and UO_1731 (O_1731,N_23343,N_25299);
nor UO_1732 (O_1732,N_29777,N_25227);
nand UO_1733 (O_1733,N_25601,N_23594);
nand UO_1734 (O_1734,N_20933,N_28391);
or UO_1735 (O_1735,N_24141,N_25305);
and UO_1736 (O_1736,N_26669,N_20713);
and UO_1737 (O_1737,N_23867,N_24750);
and UO_1738 (O_1738,N_23697,N_28289);
nor UO_1739 (O_1739,N_27742,N_20633);
nor UO_1740 (O_1740,N_21654,N_27441);
and UO_1741 (O_1741,N_27035,N_27847);
xnor UO_1742 (O_1742,N_25888,N_23346);
nand UO_1743 (O_1743,N_23147,N_24511);
nand UO_1744 (O_1744,N_25514,N_23324);
or UO_1745 (O_1745,N_26735,N_23665);
and UO_1746 (O_1746,N_29239,N_24129);
nor UO_1747 (O_1747,N_21486,N_23678);
or UO_1748 (O_1748,N_20409,N_25187);
and UO_1749 (O_1749,N_23111,N_29198);
and UO_1750 (O_1750,N_22247,N_25185);
and UO_1751 (O_1751,N_25341,N_23661);
nor UO_1752 (O_1752,N_25006,N_21018);
or UO_1753 (O_1753,N_21624,N_25328);
or UO_1754 (O_1754,N_27525,N_27682);
and UO_1755 (O_1755,N_29145,N_26880);
nor UO_1756 (O_1756,N_27793,N_23156);
nand UO_1757 (O_1757,N_21140,N_22323);
nand UO_1758 (O_1758,N_29017,N_21217);
nor UO_1759 (O_1759,N_20028,N_29270);
nor UO_1760 (O_1760,N_25427,N_21974);
nor UO_1761 (O_1761,N_22020,N_25457);
nor UO_1762 (O_1762,N_27568,N_29518);
nor UO_1763 (O_1763,N_29085,N_25518);
nand UO_1764 (O_1764,N_21886,N_27386);
and UO_1765 (O_1765,N_29637,N_20699);
nor UO_1766 (O_1766,N_22607,N_27302);
nand UO_1767 (O_1767,N_29562,N_29486);
nor UO_1768 (O_1768,N_28157,N_20794);
or UO_1769 (O_1769,N_27260,N_22717);
nand UO_1770 (O_1770,N_26278,N_20666);
nand UO_1771 (O_1771,N_22941,N_24967);
and UO_1772 (O_1772,N_27770,N_24617);
and UO_1773 (O_1773,N_20769,N_27476);
nand UO_1774 (O_1774,N_26490,N_25456);
or UO_1775 (O_1775,N_27435,N_22424);
nor UO_1776 (O_1776,N_22636,N_25596);
nand UO_1777 (O_1777,N_20041,N_28749);
nor UO_1778 (O_1778,N_24364,N_23325);
nor UO_1779 (O_1779,N_22092,N_25500);
nor UO_1780 (O_1780,N_27168,N_25586);
or UO_1781 (O_1781,N_25905,N_22249);
nor UO_1782 (O_1782,N_24793,N_24813);
and UO_1783 (O_1783,N_28493,N_22962);
nor UO_1784 (O_1784,N_22638,N_25506);
xor UO_1785 (O_1785,N_23018,N_23168);
nor UO_1786 (O_1786,N_21220,N_25364);
nand UO_1787 (O_1787,N_22738,N_21885);
and UO_1788 (O_1788,N_24802,N_22107);
nand UO_1789 (O_1789,N_23354,N_27865);
nand UO_1790 (O_1790,N_24885,N_22205);
or UO_1791 (O_1791,N_26728,N_20958);
nand UO_1792 (O_1792,N_22395,N_24151);
or UO_1793 (O_1793,N_22791,N_25585);
nand UO_1794 (O_1794,N_26494,N_29957);
or UO_1795 (O_1795,N_27178,N_22299);
nand UO_1796 (O_1796,N_25530,N_25629);
nand UO_1797 (O_1797,N_25864,N_21000);
or UO_1798 (O_1798,N_27021,N_26128);
or UO_1799 (O_1799,N_28189,N_28610);
or UO_1800 (O_1800,N_27445,N_24162);
or UO_1801 (O_1801,N_21564,N_29965);
and UO_1802 (O_1802,N_24463,N_26581);
nor UO_1803 (O_1803,N_24161,N_23589);
or UO_1804 (O_1804,N_22550,N_24782);
nor UO_1805 (O_1805,N_20926,N_21274);
nand UO_1806 (O_1806,N_21177,N_29879);
and UO_1807 (O_1807,N_22748,N_20266);
nor UO_1808 (O_1808,N_29826,N_29607);
nand UO_1809 (O_1809,N_27091,N_26653);
nor UO_1810 (O_1810,N_29727,N_27076);
nor UO_1811 (O_1811,N_21307,N_20721);
and UO_1812 (O_1812,N_21052,N_27053);
or UO_1813 (O_1813,N_28640,N_27618);
nor UO_1814 (O_1814,N_27093,N_27573);
or UO_1815 (O_1815,N_23164,N_26311);
and UO_1816 (O_1816,N_28850,N_20826);
or UO_1817 (O_1817,N_24723,N_22056);
nand UO_1818 (O_1818,N_26153,N_28506);
nand UO_1819 (O_1819,N_28117,N_27656);
nand UO_1820 (O_1820,N_20324,N_21980);
and UO_1821 (O_1821,N_20149,N_26603);
nand UO_1822 (O_1822,N_27651,N_22572);
and UO_1823 (O_1823,N_29544,N_22910);
and UO_1824 (O_1824,N_20492,N_22970);
or UO_1825 (O_1825,N_23065,N_23083);
nor UO_1826 (O_1826,N_26167,N_24917);
or UO_1827 (O_1827,N_22482,N_27961);
nand UO_1828 (O_1828,N_24955,N_22086);
or UO_1829 (O_1829,N_29676,N_28987);
or UO_1830 (O_1830,N_26203,N_20593);
or UO_1831 (O_1831,N_29387,N_22657);
or UO_1832 (O_1832,N_23285,N_22567);
or UO_1833 (O_1833,N_26135,N_24753);
or UO_1834 (O_1834,N_26716,N_21796);
and UO_1835 (O_1835,N_23750,N_25664);
and UO_1836 (O_1836,N_25754,N_21775);
nand UO_1837 (O_1837,N_21278,N_24344);
or UO_1838 (O_1838,N_29382,N_25798);
or UO_1839 (O_1839,N_23903,N_24707);
nand UO_1840 (O_1840,N_26563,N_21399);
nor UO_1841 (O_1841,N_20351,N_20382);
or UO_1842 (O_1842,N_25375,N_24740);
and UO_1843 (O_1843,N_26109,N_24016);
nor UO_1844 (O_1844,N_20288,N_26738);
nor UO_1845 (O_1845,N_29090,N_24689);
nand UO_1846 (O_1846,N_22735,N_21398);
nor UO_1847 (O_1847,N_21729,N_26501);
or UO_1848 (O_1848,N_25363,N_22403);
nor UO_1849 (O_1849,N_23711,N_25037);
nor UO_1850 (O_1850,N_25821,N_21546);
or UO_1851 (O_1851,N_25573,N_26598);
xor UO_1852 (O_1852,N_22672,N_27551);
or UO_1853 (O_1853,N_27887,N_21921);
or UO_1854 (O_1854,N_28082,N_27969);
nand UO_1855 (O_1855,N_20816,N_26697);
or UO_1856 (O_1856,N_27603,N_25020);
nand UO_1857 (O_1857,N_27913,N_23028);
and UO_1858 (O_1858,N_23003,N_24034);
nand UO_1859 (O_1859,N_26284,N_23814);
or UO_1860 (O_1860,N_20888,N_27365);
nand UO_1861 (O_1861,N_26266,N_24010);
or UO_1862 (O_1862,N_26060,N_22838);
nand UO_1863 (O_1863,N_28589,N_22252);
nand UO_1864 (O_1864,N_26564,N_25102);
nor UO_1865 (O_1865,N_29747,N_27938);
xor UO_1866 (O_1866,N_21820,N_25833);
nand UO_1867 (O_1867,N_24022,N_21457);
and UO_1868 (O_1868,N_21933,N_25481);
or UO_1869 (O_1869,N_28677,N_25955);
nand UO_1870 (O_1870,N_22057,N_21515);
or UO_1871 (O_1871,N_28479,N_24629);
or UO_1872 (O_1872,N_25218,N_21460);
nand UO_1873 (O_1873,N_22913,N_28355);
and UO_1874 (O_1874,N_23893,N_22943);
or UO_1875 (O_1875,N_25284,N_28390);
nor UO_1876 (O_1876,N_27761,N_28106);
or UO_1877 (O_1877,N_22496,N_23578);
and UO_1878 (O_1878,N_26642,N_20364);
or UO_1879 (O_1879,N_24666,N_22630);
nor UO_1880 (O_1880,N_22437,N_20125);
nor UO_1881 (O_1881,N_28905,N_26292);
nand UO_1882 (O_1882,N_29135,N_23694);
and UO_1883 (O_1883,N_22661,N_24221);
and UO_1884 (O_1884,N_26571,N_29983);
nor UO_1885 (O_1885,N_25543,N_26982);
nand UO_1886 (O_1886,N_28057,N_29960);
nor UO_1887 (O_1887,N_26381,N_27987);
or UO_1888 (O_1888,N_28670,N_29244);
or UO_1889 (O_1889,N_29555,N_29883);
nand UO_1890 (O_1890,N_25174,N_22514);
nand UO_1891 (O_1891,N_22330,N_23306);
nor UO_1892 (O_1892,N_21642,N_26086);
and UO_1893 (O_1893,N_26078,N_25226);
nand UO_1894 (O_1894,N_25309,N_27057);
and UO_1895 (O_1895,N_29767,N_23272);
xor UO_1896 (O_1896,N_20102,N_23849);
nand UO_1897 (O_1897,N_26229,N_24999);
nand UO_1898 (O_1898,N_25483,N_24683);
or UO_1899 (O_1899,N_25809,N_24743);
or UO_1900 (O_1900,N_27559,N_24867);
xnor UO_1901 (O_1901,N_29193,N_27635);
and UO_1902 (O_1902,N_27879,N_26597);
and UO_1903 (O_1903,N_29564,N_22219);
or UO_1904 (O_1904,N_24318,N_25927);
nor UO_1905 (O_1905,N_28730,N_25486);
nand UO_1906 (O_1906,N_28006,N_28032);
and UO_1907 (O_1907,N_29596,N_28376);
or UO_1908 (O_1908,N_28710,N_29726);
nand UO_1909 (O_1909,N_28839,N_27542);
and UO_1910 (O_1910,N_20635,N_23128);
nor UO_1911 (O_1911,N_29683,N_28773);
or UO_1912 (O_1912,N_25991,N_21753);
or UO_1913 (O_1913,N_25250,N_21157);
or UO_1914 (O_1914,N_29738,N_27354);
nand UO_1915 (O_1915,N_24515,N_26761);
and UO_1916 (O_1916,N_24631,N_28725);
or UO_1917 (O_1917,N_26023,N_21827);
and UO_1918 (O_1918,N_25487,N_29157);
nand UO_1919 (O_1919,N_28620,N_25708);
nor UO_1920 (O_1920,N_21127,N_20565);
or UO_1921 (O_1921,N_27101,N_25828);
nor UO_1922 (O_1922,N_22957,N_29407);
nand UO_1923 (O_1923,N_21355,N_25848);
and UO_1924 (O_1924,N_20085,N_20095);
and UO_1925 (O_1925,N_26588,N_25994);
nor UO_1926 (O_1926,N_26422,N_27721);
nor UO_1927 (O_1927,N_20403,N_24754);
nand UO_1928 (O_1928,N_29092,N_21676);
nor UO_1929 (O_1929,N_20279,N_29780);
nor UO_1930 (O_1930,N_20731,N_27124);
and UO_1931 (O_1931,N_20127,N_20307);
or UO_1932 (O_1932,N_24765,N_25949);
or UO_1933 (O_1933,N_28091,N_26958);
nand UO_1934 (O_1934,N_20554,N_28959);
nand UO_1935 (O_1935,N_27963,N_25342);
or UO_1936 (O_1936,N_29367,N_25936);
nor UO_1937 (O_1937,N_20253,N_26355);
or UO_1938 (O_1938,N_20430,N_28965);
nand UO_1939 (O_1939,N_29074,N_29694);
nor UO_1940 (O_1940,N_29867,N_29255);
nor UO_1941 (O_1941,N_27501,N_24273);
and UO_1942 (O_1942,N_24645,N_27285);
xnor UO_1943 (O_1943,N_20330,N_25823);
and UO_1944 (O_1944,N_22499,N_24556);
and UO_1945 (O_1945,N_21714,N_26281);
nor UO_1946 (O_1946,N_27579,N_20618);
and UO_1947 (O_1947,N_26955,N_27946);
nand UO_1948 (O_1948,N_29070,N_24039);
nor UO_1949 (O_1949,N_22660,N_21670);
nand UO_1950 (O_1950,N_26637,N_28229);
nor UO_1951 (O_1951,N_22606,N_23460);
nand UO_1952 (O_1952,N_29172,N_24008);
nor UO_1953 (O_1953,N_27331,N_23091);
or UO_1954 (O_1954,N_26334,N_20017);
xor UO_1955 (O_1955,N_24498,N_27363);
or UO_1956 (O_1956,N_25116,N_21171);
nand UO_1957 (O_1957,N_29151,N_28336);
nor UO_1958 (O_1958,N_22839,N_27590);
and UO_1959 (O_1959,N_26606,N_28898);
and UO_1960 (O_1960,N_28049,N_29881);
nand UO_1961 (O_1961,N_27106,N_22268);
nor UO_1962 (O_1962,N_29308,N_25626);
nor UO_1963 (O_1963,N_20854,N_21472);
nand UO_1964 (O_1964,N_29986,N_29150);
nand UO_1965 (O_1965,N_22816,N_22226);
nand UO_1966 (O_1966,N_21602,N_28840);
nand UO_1967 (O_1967,N_27086,N_28920);
or UO_1968 (O_1968,N_20690,N_21173);
and UO_1969 (O_1969,N_24812,N_26207);
xor UO_1970 (O_1970,N_25000,N_28415);
nand UO_1971 (O_1971,N_26715,N_20259);
nor UO_1972 (O_1972,N_22809,N_23123);
nor UO_1973 (O_1973,N_28778,N_24328);
nor UO_1974 (O_1974,N_24373,N_23180);
nor UO_1975 (O_1975,N_21615,N_21524);
nand UO_1976 (O_1976,N_25243,N_24116);
and UO_1977 (O_1977,N_23636,N_28760);
or UO_1978 (O_1978,N_28420,N_24551);
or UO_1979 (O_1979,N_23799,N_24313);
or UO_1980 (O_1980,N_27791,N_27532);
nor UO_1981 (O_1981,N_23121,N_23383);
nand UO_1982 (O_1982,N_22989,N_21674);
nand UO_1983 (O_1983,N_20737,N_23819);
nand UO_1984 (O_1984,N_21851,N_24571);
nand UO_1985 (O_1985,N_29242,N_27653);
or UO_1986 (O_1986,N_26874,N_26695);
nor UO_1987 (O_1987,N_24888,N_24658);
or UO_1988 (O_1988,N_25472,N_21247);
xor UO_1989 (O_1989,N_21263,N_20668);
and UO_1990 (O_1990,N_22914,N_25436);
and UO_1991 (O_1991,N_26674,N_23204);
nand UO_1992 (O_1992,N_23355,N_24212);
and UO_1993 (O_1993,N_20550,N_22090);
nor UO_1994 (O_1994,N_26800,N_29941);
nor UO_1995 (O_1995,N_29809,N_20422);
nand UO_1996 (O_1996,N_21004,N_26890);
nor UO_1997 (O_1997,N_22963,N_20548);
or UO_1998 (O_1998,N_24272,N_20882);
nand UO_1999 (O_1999,N_28231,N_26132);
and UO_2000 (O_2000,N_20113,N_24046);
or UO_2001 (O_2001,N_28194,N_26770);
or UO_2002 (O_2002,N_28160,N_20193);
nor UO_2003 (O_2003,N_27755,N_20267);
nor UO_2004 (O_2004,N_24333,N_25340);
and UO_2005 (O_2005,N_28450,N_29959);
xor UO_2006 (O_2006,N_21010,N_28577);
nor UO_2007 (O_2007,N_25092,N_26634);
or UO_2008 (O_2008,N_25039,N_29066);
nor UO_2009 (O_2009,N_21292,N_28249);
and UO_2010 (O_2010,N_24182,N_25405);
nor UO_2011 (O_2011,N_27935,N_20286);
nor UO_2012 (O_2012,N_26001,N_22035);
nor UO_2013 (O_2013,N_22402,N_29869);
or UO_2014 (O_2014,N_23141,N_29013);
and UO_2015 (O_2015,N_29274,N_25937);
and UO_2016 (O_2016,N_29077,N_27743);
or UO_2017 (O_2017,N_28568,N_23475);
and UO_2018 (O_2018,N_21703,N_23426);
nor UO_2019 (O_2019,N_29774,N_28191);
and UO_2020 (O_2020,N_28440,N_27670);
or UO_2021 (O_2021,N_24348,N_27480);
nor UO_2022 (O_2022,N_27248,N_26677);
nand UO_2023 (O_2023,N_20272,N_25160);
or UO_2024 (O_2024,N_22044,N_29015);
nor UO_2025 (O_2025,N_28991,N_24011);
nand UO_2026 (O_2026,N_29638,N_25455);
nand UO_2027 (O_2027,N_24325,N_29893);
nand UO_2028 (O_2028,N_28364,N_21575);
and UO_2029 (O_2029,N_27304,N_21562);
and UO_2030 (O_2030,N_23970,N_25691);
or UO_2031 (O_2031,N_25836,N_21209);
or UO_2032 (O_2032,N_24642,N_26386);
and UO_2033 (O_2033,N_20015,N_20401);
or UO_2034 (O_2034,N_21586,N_26794);
nand UO_2035 (O_2035,N_26274,N_28504);
and UO_2036 (O_2036,N_29899,N_29267);
nor UO_2037 (O_2037,N_29643,N_27425);
nor UO_2038 (O_2038,N_24357,N_24937);
nor UO_2039 (O_2039,N_24314,N_29485);
or UO_2040 (O_2040,N_26076,N_23532);
and UO_2041 (O_2041,N_27833,N_26541);
or UO_2042 (O_2042,N_25791,N_29030);
nor UO_2043 (O_2043,N_28726,N_24701);
and UO_2044 (O_2044,N_23576,N_21370);
and UO_2045 (O_2045,N_26213,N_21354);
nor UO_2046 (O_2046,N_20659,N_23999);
and UO_2047 (O_2047,N_26247,N_21391);
or UO_2048 (O_2048,N_20758,N_24612);
nand UO_2049 (O_2049,N_29217,N_22450);
nand UO_2050 (O_2050,N_27578,N_25194);
nor UO_2051 (O_2051,N_25547,N_20571);
nand UO_2052 (O_2052,N_29022,N_25032);
and UO_2053 (O_2053,N_28812,N_23523);
nand UO_2054 (O_2054,N_22328,N_28688);
and UO_2055 (O_2055,N_22895,N_28358);
nand UO_2056 (O_2056,N_25426,N_22576);
nor UO_2057 (O_2057,N_25264,N_26444);
nor UO_2058 (O_2058,N_24659,N_22757);
and UO_2059 (O_2059,N_22225,N_28889);
nand UO_2060 (O_2060,N_22296,N_24362);
and UO_2061 (O_2061,N_26461,N_22756);
and UO_2062 (O_2062,N_28368,N_20719);
nor UO_2063 (O_2063,N_20150,N_25958);
nor UO_2064 (O_2064,N_20449,N_24497);
nand UO_2065 (O_2065,N_28994,N_27032);
and UO_2066 (O_2066,N_25694,N_29060);
or UO_2067 (O_2067,N_22378,N_25469);
or UO_2068 (O_2068,N_27361,N_25149);
nor UO_2069 (O_2069,N_28462,N_29475);
nand UO_2070 (O_2070,N_20952,N_25682);
or UO_2071 (O_2071,N_27416,N_21114);
or UO_2072 (O_2072,N_29305,N_29238);
or UO_2073 (O_2073,N_26024,N_26020);
xor UO_2074 (O_2074,N_23659,N_20761);
nand UO_2075 (O_2075,N_29354,N_28104);
and UO_2076 (O_2076,N_28035,N_24341);
or UO_2077 (O_2077,N_29895,N_29542);
nor UO_2078 (O_2078,N_20519,N_27754);
and UO_2079 (O_2079,N_21107,N_20732);
or UO_2080 (O_2080,N_24040,N_23846);
and UO_2081 (O_2081,N_20460,N_21843);
and UO_2082 (O_2082,N_20278,N_23830);
and UO_2083 (O_2083,N_23542,N_24174);
or UO_2084 (O_2084,N_29177,N_20427);
and UO_2085 (O_2085,N_20620,N_26068);
nor UO_2086 (O_2086,N_28486,N_22988);
nor UO_2087 (O_2087,N_20356,N_28412);
nand UO_2088 (O_2088,N_24601,N_20517);
nand UO_2089 (O_2089,N_24591,N_29269);
nor UO_2090 (O_2090,N_26847,N_21696);
nand UO_2091 (O_2091,N_25407,N_26645);
nor UO_2092 (O_2092,N_21284,N_20083);
and UO_2093 (O_2093,N_29762,N_29009);
or UO_2094 (O_2094,N_21954,N_26004);
or UO_2095 (O_2095,N_24624,N_23481);
nor UO_2096 (O_2096,N_23115,N_26117);
or UO_2097 (O_2097,N_22870,N_22676);
nor UO_2098 (O_2098,N_29565,N_27013);
nor UO_2099 (O_2099,N_27647,N_21405);
nor UO_2100 (O_2100,N_21964,N_27563);
or UO_2101 (O_2101,N_20867,N_24139);
or UO_2102 (O_2102,N_27379,N_22266);
nand UO_2103 (O_2103,N_27122,N_28174);
or UO_2104 (O_2104,N_24940,N_27846);
and UO_2105 (O_2105,N_23038,N_27634);
and UO_2106 (O_2106,N_24014,N_28658);
or UO_2107 (O_2107,N_26902,N_24140);
and UO_2108 (O_2108,N_27227,N_21965);
and UO_2109 (O_2109,N_20133,N_25241);
nand UO_2110 (O_2110,N_22503,N_24710);
or UO_2111 (O_2111,N_24943,N_28365);
or UO_2112 (O_2112,N_29072,N_27829);
nor UO_2113 (O_2113,N_22708,N_21817);
nand UO_2114 (O_2114,N_24623,N_25246);
nand UO_2115 (O_2115,N_27112,N_26789);
nand UO_2116 (O_2116,N_21167,N_22145);
nand UO_2117 (O_2117,N_22133,N_22955);
nand UO_2118 (O_2118,N_26648,N_27974);
nand UO_2119 (O_2119,N_21498,N_23139);
nor UO_2120 (O_2120,N_29119,N_29479);
nand UO_2121 (O_2121,N_24693,N_21612);
nand UO_2122 (O_2122,N_29404,N_29277);
and UO_2123 (O_2123,N_28275,N_26773);
or UO_2124 (O_2124,N_28598,N_27418);
nand UO_2125 (O_2125,N_24469,N_21547);
nor UO_2126 (O_2126,N_24670,N_23525);
nor UO_2127 (O_2127,N_20832,N_28906);
xor UO_2128 (O_2128,N_25561,N_26352);
nor UO_2129 (O_2129,N_22596,N_22566);
or UO_2130 (O_2130,N_29362,N_23848);
nand UO_2131 (O_2131,N_24452,N_21230);
nor UO_2132 (O_2132,N_22537,N_26737);
and UO_2133 (O_2133,N_22471,N_20613);
or UO_2134 (O_2134,N_28347,N_22423);
nor UO_2135 (O_2135,N_25741,N_23172);
or UO_2136 (O_2136,N_22479,N_29275);
nand UO_2137 (O_2137,N_20811,N_29863);
nand UO_2138 (O_2138,N_23623,N_21188);
nor UO_2139 (O_2139,N_27789,N_29608);
nor UO_2140 (O_2140,N_29801,N_22231);
or UO_2141 (O_2141,N_27509,N_29525);
nand UO_2142 (O_2142,N_27103,N_29823);
and UO_2143 (O_2143,N_28633,N_21053);
nor UO_2144 (O_2144,N_23463,N_20159);
nand UO_2145 (O_2145,N_21184,N_27648);
nand UO_2146 (O_2146,N_28926,N_26974);
or UO_2147 (O_2147,N_27266,N_22507);
or UO_2148 (O_2148,N_21137,N_27502);
nor UO_2149 (O_2149,N_25663,N_27683);
nor UO_2150 (O_2150,N_27861,N_23056);
and UO_2151 (O_2151,N_20116,N_26798);
or UO_2152 (O_2152,N_25302,N_28744);
nand UO_2153 (O_2153,N_22902,N_26025);
and UO_2154 (O_2154,N_26474,N_26051);
and UO_2155 (O_2155,N_21966,N_28252);
and UO_2156 (O_2156,N_22918,N_24863);
nor UO_2157 (O_2157,N_21174,N_28573);
nand UO_2158 (O_2158,N_27351,N_23280);
nand UO_2159 (O_2159,N_28142,N_26112);
or UO_2160 (O_2160,N_21487,N_21350);
nor UO_2161 (O_2161,N_24393,N_25470);
nor UO_2162 (O_2162,N_28707,N_27607);
and UO_2163 (O_2163,N_25493,N_23836);
nand UO_2164 (O_2164,N_29569,N_21483);
nor UO_2165 (O_2165,N_25997,N_26510);
nand UO_2166 (O_2166,N_21334,N_22840);
and UO_2167 (O_2167,N_24461,N_25627);
nor UO_2168 (O_2168,N_21496,N_24680);
nor UO_2169 (O_2169,N_27669,N_23078);
and UO_2170 (O_2170,N_21035,N_22153);
nand UO_2171 (O_2171,N_25652,N_28910);
nor UO_2172 (O_2172,N_21620,N_28303);
or UO_2173 (O_2173,N_27520,N_27687);
nand UO_2174 (O_2174,N_27985,N_21785);
and UO_2175 (O_2175,N_23477,N_23996);
nor UO_2176 (O_2176,N_25939,N_27192);
nand UO_2177 (O_2177,N_25761,N_20252);
nor UO_2178 (O_2178,N_27350,N_26787);
nor UO_2179 (O_2179,N_26326,N_25890);
nor UO_2180 (O_2180,N_24695,N_24785);
nor UO_2181 (O_2181,N_22825,N_29521);
nor UO_2182 (O_2182,N_20013,N_29749);
nand UO_2183 (O_2183,N_20818,N_27151);
nand UO_2184 (O_2184,N_21094,N_26199);
and UO_2185 (O_2185,N_28286,N_28807);
and UO_2186 (O_2186,N_23958,N_23321);
nand UO_2187 (O_2187,N_20146,N_22082);
and UO_2188 (O_2188,N_26932,N_21505);
nor UO_2189 (O_2189,N_25632,N_27734);
or UO_2190 (O_2190,N_23297,N_27973);
nand UO_2191 (O_2191,N_29532,N_24292);
and UO_2192 (O_2192,N_25482,N_21118);
and UO_2193 (O_2193,N_21181,N_29125);
and UO_2194 (O_2194,N_28492,N_26951);
and UO_2195 (O_2195,N_26106,N_20697);
nor UO_2196 (O_2196,N_26385,N_26007);
nand UO_2197 (O_2197,N_20642,N_26687);
or UO_2198 (O_2198,N_21876,N_29192);
and UO_2199 (O_2199,N_22564,N_24746);
nor UO_2200 (O_2200,N_23864,N_25272);
nor UO_2201 (O_2201,N_24386,N_27513);
nand UO_2202 (O_2202,N_24250,N_29394);
or UO_2203 (O_2203,N_24366,N_23370);
and UO_2204 (O_2204,N_26022,N_29724);
and UO_2205 (O_2205,N_28996,N_27451);
or UO_2206 (O_2206,N_21383,N_22124);
nor UO_2207 (O_2207,N_22808,N_24927);
and UO_2208 (O_2208,N_24699,N_22722);
xor UO_2209 (O_2209,N_20573,N_23344);
nor UO_2210 (O_2210,N_28214,N_22431);
and UO_2211 (O_2211,N_21995,N_23720);
or UO_2212 (O_2212,N_24696,N_29633);
nand UO_2213 (O_2213,N_21338,N_27241);
and UO_2214 (O_2214,N_23243,N_20813);
or UO_2215 (O_2215,N_21036,N_29613);
nand UO_2216 (O_2216,N_26156,N_28671);
nand UO_2217 (O_2217,N_20707,N_29938);
or UO_2218 (O_2218,N_27335,N_23284);
and UO_2219 (O_2219,N_21743,N_27495);
or UO_2220 (O_2220,N_23251,N_26838);
and UO_2221 (O_2221,N_20437,N_23875);
nor UO_2222 (O_2222,N_20805,N_28149);
and UO_2223 (O_2223,N_29481,N_29304);
or UO_2224 (O_2224,N_25494,N_25461);
or UO_2225 (O_2225,N_26554,N_29536);
nand UO_2226 (O_2226,N_27494,N_29592);
or UO_2227 (O_2227,N_23483,N_29473);
nand UO_2228 (O_2228,N_21417,N_28883);
nor UO_2229 (O_2229,N_22342,N_21271);
nand UO_2230 (O_2230,N_29228,N_23766);
or UO_2231 (O_2231,N_25345,N_26347);
nor UO_2232 (O_2232,N_29344,N_22463);
nor UO_2233 (O_2233,N_20597,N_21011);
or UO_2234 (O_2234,N_29876,N_29949);
or UO_2235 (O_2235,N_23724,N_28715);
and UO_2236 (O_2236,N_22721,N_20175);
xor UO_2237 (O_2237,N_25987,N_23010);
nand UO_2238 (O_2238,N_21169,N_28869);
nor UO_2239 (O_2239,N_20453,N_20282);
nand UO_2240 (O_2240,N_21846,N_23269);
nor UO_2241 (O_2241,N_29998,N_22409);
or UO_2242 (O_2242,N_29653,N_26556);
or UO_2243 (O_2243,N_24057,N_23401);
nor UO_2244 (O_2244,N_23950,N_22418);
nor UO_2245 (O_2245,N_26819,N_20152);
or UO_2246 (O_2246,N_24833,N_28060);
xor UO_2247 (O_2247,N_25609,N_22449);
nor UO_2248 (O_2248,N_29556,N_28130);
and UO_2249 (O_2249,N_26835,N_23508);
and UO_2250 (O_2250,N_22767,N_23995);
and UO_2251 (O_2251,N_23890,N_22195);
or UO_2252 (O_2252,N_22272,N_21856);
nor UO_2253 (O_2253,N_27729,N_25594);
nand UO_2254 (O_2254,N_27531,N_27157);
nand UO_2255 (O_2255,N_20766,N_27170);
nand UO_2256 (O_2256,N_26993,N_29898);
and UO_2257 (O_2257,N_28406,N_25541);
nand UO_2258 (O_2258,N_28132,N_23035);
or UO_2259 (O_2259,N_25320,N_23685);
nand UO_2260 (O_2260,N_25141,N_23506);
nor UO_2261 (O_2261,N_21410,N_29417);
and UO_2262 (O_2262,N_23759,N_21145);
or UO_2263 (O_2263,N_29975,N_25868);
and UO_2264 (O_2264,N_23230,N_29528);
or UO_2265 (O_2265,N_24083,N_22422);
nor UO_2266 (O_2266,N_24191,N_22880);
nand UO_2267 (O_2267,N_22958,N_26957);
nor UO_2268 (O_2268,N_21144,N_25070);
nand UO_2269 (O_2269,N_21759,N_20353);
xor UO_2270 (O_2270,N_26666,N_28846);
nand UO_2271 (O_2271,N_22102,N_29434);
nor UO_2272 (O_2272,N_22546,N_24110);
and UO_2273 (O_2273,N_26580,N_26496);
nand UO_2274 (O_2274,N_28762,N_25863);
nor UO_2275 (O_2275,N_28613,N_20431);
and UO_2276 (O_2276,N_25973,N_29427);
or UO_2277 (O_2277,N_27415,N_29445);
nand UO_2278 (O_2278,N_24117,N_23563);
or UO_2279 (O_2279,N_28359,N_28731);
nor UO_2280 (O_2280,N_22224,N_21521);
and UO_2281 (O_2281,N_23920,N_29409);
nand UO_2282 (O_2282,N_29158,N_28951);
nor UO_2283 (O_2283,N_20289,N_25515);
and UO_2284 (O_2284,N_28983,N_28596);
or UO_2285 (O_2285,N_21091,N_22667);
nor UO_2286 (O_2286,N_25995,N_22366);
nor UO_2287 (O_2287,N_28660,N_29310);
nand UO_2288 (O_2288,N_21488,N_29452);
nor UO_2289 (O_2289,N_21302,N_24977);
or UO_2290 (O_2290,N_26152,N_21087);
and UO_2291 (O_2291,N_21721,N_27995);
nor UO_2292 (O_2292,N_20218,N_23212);
or UO_2293 (O_2293,N_28316,N_28830);
nor UO_2294 (O_2294,N_28721,N_21051);
or UO_2295 (O_2295,N_21687,N_20558);
nor UO_2296 (O_2296,N_29690,N_21426);
xnor UO_2297 (O_2297,N_20669,N_29628);
and UO_2298 (O_2298,N_22081,N_24906);
and UO_2299 (O_2299,N_22148,N_25352);
nand UO_2300 (O_2300,N_27081,N_23728);
or UO_2301 (O_2301,N_29484,N_28111);
or UO_2302 (O_2302,N_29487,N_26300);
xor UO_2303 (O_2303,N_23445,N_23427);
nor UO_2304 (O_2304,N_28708,N_27483);
nor UO_2305 (O_2305,N_24832,N_27121);
nand UO_2306 (O_2306,N_21794,N_25077);
nor UO_2307 (O_2307,N_24735,N_23741);
nand UO_2308 (O_2308,N_21180,N_24894);
or UO_2309 (O_2309,N_29860,N_25491);
or UO_2310 (O_2310,N_20185,N_25048);
and UO_2311 (O_2311,N_25231,N_21429);
nand UO_2312 (O_2312,N_23396,N_20905);
nand UO_2313 (O_2313,N_22269,N_27814);
nor UO_2314 (O_2314,N_25794,N_27205);
nand UO_2315 (O_2315,N_20235,N_22656);
or UO_2316 (O_2316,N_25480,N_28743);
nor UO_2317 (O_2317,N_23288,N_27292);
or UO_2318 (O_2318,N_22321,N_21538);
nand UO_2319 (O_2319,N_24662,N_23000);
nand UO_2320 (O_2320,N_27060,N_28036);
and UO_2321 (O_2321,N_29668,N_28791);
nand UO_2322 (O_2322,N_26660,N_26433);
nor UO_2323 (O_2323,N_25462,N_27166);
or UO_2324 (O_2324,N_26905,N_24321);
and UO_2325 (O_2325,N_20667,N_20319);
or UO_2326 (O_2326,N_21187,N_20628);
nand UO_2327 (O_2327,N_23126,N_21361);
or UO_2328 (O_2328,N_27045,N_29410);
and UO_2329 (O_2329,N_28373,N_24078);
and UO_2330 (O_2330,N_27099,N_23402);
nor UO_2331 (O_2331,N_21938,N_26104);
nor UO_2332 (O_2332,N_29583,N_20473);
and UO_2333 (O_2333,N_26610,N_26646);
nand UO_2334 (O_2334,N_22716,N_23780);
nand UO_2335 (O_2335,N_27034,N_28822);
and UO_2336 (O_2336,N_23627,N_28449);
or UO_2337 (O_2337,N_24932,N_24001);
or UO_2338 (O_2338,N_25599,N_28239);
and UO_2339 (O_2339,N_23052,N_22179);
nor UO_2340 (O_2340,N_28304,N_29886);
or UO_2341 (O_2341,N_24539,N_29850);
nor UO_2342 (O_2342,N_29561,N_21013);
or UO_2343 (O_2343,N_23505,N_22146);
xnor UO_2344 (O_2344,N_20595,N_25281);
nand UO_2345 (O_2345,N_20039,N_26584);
nor UO_2346 (O_2346,N_24528,N_20772);
nor UO_2347 (O_2347,N_21221,N_24446);
or UO_2348 (O_2348,N_29361,N_24952);
nand UO_2349 (O_2349,N_22590,N_25359);
nor UO_2350 (O_2350,N_24429,N_20178);
or UO_2351 (O_2351,N_25497,N_25554);
and UO_2352 (O_2352,N_26432,N_26780);
nor UO_2353 (O_2353,N_28099,N_21396);
and UO_2354 (O_2354,N_21605,N_21802);
or UO_2355 (O_2355,N_28276,N_25783);
and UO_2356 (O_2356,N_27442,N_22600);
and UO_2357 (O_2357,N_28984,N_26854);
or UO_2358 (O_2358,N_21849,N_23551);
nor UO_2359 (O_2359,N_28087,N_27211);
nand UO_2360 (O_2360,N_26313,N_20977);
nand UO_2361 (O_2361,N_26705,N_20706);
nand UO_2362 (O_2362,N_26148,N_20998);
nand UO_2363 (O_2363,N_25673,N_21588);
and UO_2364 (O_2364,N_24090,N_22691);
and UO_2365 (O_2365,N_21740,N_25685);
nand UO_2366 (O_2366,N_28899,N_25932);
nand UO_2367 (O_2367,N_22710,N_27468);
nor UO_2368 (O_2368,N_27403,N_28204);
nand UO_2369 (O_2369,N_24367,N_21218);
or UO_2370 (O_2370,N_23019,N_20141);
nor UO_2371 (O_2371,N_21683,N_26095);
nor UO_2372 (O_2372,N_25004,N_21611);
nor UO_2373 (O_2373,N_20968,N_24267);
nor UO_2374 (O_2374,N_27741,N_25684);
or UO_2375 (O_2375,N_20130,N_20834);
nor UO_2376 (O_2376,N_23567,N_22005);
and UO_2377 (O_2377,N_25052,N_21864);
nor UO_2378 (O_2378,N_24107,N_24988);
nor UO_2379 (O_2379,N_25030,N_28881);
nor UO_2380 (O_2380,N_22077,N_23795);
nor UO_2381 (O_2381,N_24973,N_22367);
nor UO_2382 (O_2382,N_20525,N_22143);
nand UO_2383 (O_2383,N_28800,N_22500);
nor UO_2384 (O_2384,N_20723,N_28636);
or UO_2385 (O_2385,N_26349,N_20609);
nor UO_2386 (O_2386,N_26679,N_26641);
nor UO_2387 (O_2387,N_24399,N_21960);
nor UO_2388 (O_2388,N_24547,N_22274);
or UO_2389 (O_2389,N_29496,N_21630);
nand UO_2390 (O_2390,N_23467,N_27890);
nor UO_2391 (O_2391,N_24806,N_22028);
nand UO_2392 (O_2392,N_27321,N_28161);
nand UO_2393 (O_2393,N_29189,N_24440);
nor UO_2394 (O_2394,N_23323,N_24136);
and UO_2395 (O_2395,N_29552,N_27031);
or UO_2396 (O_2396,N_28907,N_29752);
or UO_2397 (O_2397,N_29393,N_20084);
and UO_2398 (O_2398,N_29905,N_25199);
nor UO_2399 (O_2399,N_26769,N_23446);
or UO_2400 (O_2400,N_21403,N_28494);
and UO_2401 (O_2401,N_21891,N_26607);
or UO_2402 (O_2402,N_27583,N_28302);
and UO_2403 (O_2403,N_28820,N_24448);
nand UO_2404 (O_2404,N_28080,N_23722);
nand UO_2405 (O_2405,N_20587,N_26188);
nor UO_2406 (O_2406,N_24706,N_28168);
or UO_2407 (O_2407,N_26781,N_23607);
nor UO_2408 (O_2408,N_26141,N_21841);
or UO_2409 (O_2409,N_25533,N_20936);
nor UO_2410 (O_2410,N_29140,N_28618);
nand UO_2411 (O_2411,N_29933,N_22685);
nand UO_2412 (O_2412,N_23572,N_24288);
and UO_2413 (O_2413,N_24884,N_26613);
and UO_2414 (O_2414,N_24692,N_21168);
or UO_2415 (O_2415,N_22467,N_26075);
and UO_2416 (O_2416,N_21520,N_27585);
nand UO_2417 (O_2417,N_21126,N_21183);
and UO_2418 (O_2418,N_26868,N_25879);
and UO_2419 (O_2419,N_26657,N_22196);
and UO_2420 (O_2420,N_21366,N_28217);
nand UO_2421 (O_2421,N_27405,N_20463);
nor UO_2422 (O_2422,N_27462,N_23276);
xor UO_2423 (O_2423,N_25672,N_27130);
and UO_2424 (O_2424,N_27586,N_20914);
or UO_2425 (O_2425,N_25081,N_21449);
and UO_2426 (O_2426,N_27095,N_26372);
nor UO_2427 (O_2427,N_20365,N_26303);
or UO_2428 (O_2428,N_22903,N_28421);
nand UO_2429 (O_2429,N_23184,N_21884);
nor UO_2430 (O_2430,N_22001,N_28409);
or UO_2431 (O_2431,N_26614,N_22230);
nand UO_2432 (O_2432,N_24155,N_24504);
and UO_2433 (O_2433,N_29598,N_25593);
and UO_2434 (O_2434,N_28341,N_28998);
or UO_2435 (O_2435,N_22235,N_20701);
or UO_2436 (O_2436,N_25711,N_20871);
nor UO_2437 (O_2437,N_22163,N_21967);
and UO_2438 (O_2438,N_29584,N_29241);
nand UO_2439 (O_2439,N_26090,N_24163);
or UO_2440 (O_2440,N_28054,N_28564);
or UO_2441 (O_2441,N_24423,N_25925);
or UO_2442 (O_2442,N_24505,N_21758);
and UO_2443 (O_2443,N_24737,N_24626);
and UO_2444 (O_2444,N_27953,N_24330);
or UO_2445 (O_2445,N_21158,N_29557);
nand UO_2446 (O_2446,N_21134,N_29832);
and UO_2447 (O_2447,N_24529,N_29428);
and UO_2448 (O_2448,N_20390,N_21903);
or UO_2449 (O_2449,N_29519,N_21664);
and UO_2450 (O_2450,N_25700,N_26602);
nand UO_2451 (O_2451,N_28669,N_27988);
nand UO_2452 (O_2452,N_24258,N_24945);
or UO_2453 (O_2453,N_28170,N_22347);
or UO_2454 (O_2454,N_21888,N_24845);
nand UO_2455 (O_2455,N_28267,N_28235);
nor UO_2456 (O_2456,N_22665,N_28001);
nor UO_2457 (O_2457,N_20821,N_24029);
and UO_2458 (O_2458,N_23547,N_28273);
or UO_2459 (O_2459,N_29839,N_23666);
nand UO_2460 (O_2460,N_26525,N_20987);
and UO_2461 (O_2461,N_21093,N_29117);
and UO_2462 (O_2462,N_23331,N_29127);
xnor UO_2463 (O_2463,N_21178,N_28478);
or UO_2464 (O_2464,N_29216,N_24347);
or UO_2465 (O_2465,N_29307,N_20415);
nor UO_2466 (O_2466,N_26522,N_25327);
nand UO_2467 (O_2467,N_25267,N_23017);
or UO_2468 (O_2468,N_22114,N_24307);
nor UO_2469 (O_2469,N_23250,N_21692);
and UO_2470 (O_2470,N_25170,N_27785);
nand UO_2471 (O_2471,N_27944,N_23423);
and UO_2472 (O_2472,N_20999,N_20458);
or UO_2473 (O_2473,N_23301,N_29468);
nor UO_2474 (O_2474,N_20570,N_23608);
nor UO_2475 (O_2475,N_21002,N_28236);
nor UO_2476 (O_2476,N_20899,N_21246);
nand UO_2477 (O_2477,N_21600,N_23454);
or UO_2478 (O_2478,N_27265,N_20290);
nand UO_2479 (O_2479,N_25816,N_24809);
nand UO_2480 (O_2480,N_29884,N_25447);
and UO_2481 (O_2481,N_29864,N_28711);
and UO_2482 (O_2482,N_20717,N_29396);
nand UO_2483 (O_2483,N_24892,N_22468);
and UO_2484 (O_2484,N_28657,N_25444);
nor UO_2485 (O_2485,N_26371,N_23540);
and UO_2486 (O_2486,N_23935,N_28177);
or UO_2487 (O_2487,N_27117,N_21234);
or UO_2488 (O_2488,N_20727,N_23186);
and UO_2489 (O_2489,N_23545,N_22531);
nor UO_2490 (O_2490,N_26551,N_24807);
nor UO_2491 (O_2491,N_23794,N_24815);
and UO_2492 (O_2492,N_22795,N_26361);
or UO_2493 (O_2493,N_23076,N_22709);
nand UO_2494 (O_2494,N_24298,N_25667);
nor UO_2495 (O_2495,N_26389,N_23713);
and UO_2496 (O_2496,N_26980,N_20093);
nor UO_2497 (O_2497,N_23944,N_26234);
nor UO_2498 (O_2498,N_20830,N_28338);
nor UO_2499 (O_2499,N_27249,N_27497);
and UO_2500 (O_2500,N_20115,N_23462);
and UO_2501 (O_2501,N_29866,N_22715);
nor UO_2502 (O_2502,N_25188,N_25910);
nor UO_2503 (O_2503,N_26009,N_21001);
or UO_2504 (O_2504,N_25109,N_22298);
nand UO_2505 (O_2505,N_29558,N_27983);
or UO_2506 (O_2506,N_26376,N_22381);
and UO_2507 (O_2507,N_22727,N_26652);
nor UO_2508 (O_2508,N_27288,N_20823);
or UO_2509 (O_2509,N_26831,N_23289);
nor UO_2510 (O_2510,N_26166,N_26120);
or UO_2511 (O_2511,N_25217,N_23981);
and UO_2512 (O_2512,N_23433,N_27845);
nand UO_2513 (O_2513,N_21159,N_21574);
nor UO_2514 (O_2514,N_22075,N_24190);
nor UO_2515 (O_2515,N_22333,N_25255);
or UO_2516 (O_2516,N_22993,N_27036);
or UO_2517 (O_2517,N_26316,N_24964);
nand UO_2518 (O_2518,N_29380,N_25647);
or UO_2519 (O_2519,N_24824,N_26324);
nor UO_2520 (O_2520,N_25138,N_22362);
and UO_2521 (O_2521,N_25574,N_26860);
nor UO_2522 (O_2522,N_25413,N_26971);
nand UO_2523 (O_2523,N_24408,N_23654);
or UO_2524 (O_2524,N_28835,N_21377);
nor UO_2525 (O_2525,N_22180,N_23440);
or UO_2526 (O_2526,N_23877,N_29197);
and UO_2527 (O_2527,N_20650,N_25337);
nor UO_2528 (O_2528,N_20902,N_24264);
nor UO_2529 (O_2529,N_25257,N_20060);
or UO_2530 (O_2530,N_24164,N_28528);
nand UO_2531 (O_2531,N_23746,N_27434);
or UO_2532 (O_2532,N_20555,N_21858);
nand UO_2533 (O_2533,N_21506,N_24135);
or UO_2534 (O_2534,N_26764,N_20562);
or UO_2535 (O_2535,N_28055,N_25069);
nor UO_2536 (O_2536,N_26094,N_20086);
and UO_2537 (O_2537,N_25031,N_25722);
or UO_2538 (O_2538,N_21063,N_20393);
or UO_2539 (O_2539,N_27557,N_23352);
and UO_2540 (O_2540,N_27900,N_27325);
and UO_2541 (O_2541,N_25853,N_23341);
or UO_2542 (O_2542,N_21552,N_21450);
nor UO_2543 (O_2543,N_22489,N_29478);
nand UO_2544 (O_2544,N_26623,N_29721);
and UO_2545 (O_2545,N_26243,N_28989);
and UO_2546 (O_2546,N_28127,N_20059);
or UO_2547 (O_2547,N_24834,N_25463);
nor UO_2548 (O_2548,N_29082,N_25111);
or UO_2549 (O_2549,N_25951,N_28061);
nor UO_2550 (O_2550,N_23419,N_24965);
nor UO_2551 (O_2551,N_23955,N_26572);
or UO_2552 (O_2552,N_26670,N_21122);
and UO_2553 (O_2553,N_21902,N_20940);
nor UO_2554 (O_2554,N_23585,N_23959);
and UO_2555 (O_2555,N_27731,N_22780);
nor UO_2556 (O_2556,N_27954,N_20688);
nand UO_2557 (O_2557,N_28763,N_28768);
and UO_2558 (O_2558,N_21551,N_21101);
or UO_2559 (O_2559,N_26418,N_23847);
nor UO_2560 (O_2560,N_21867,N_26640);
or UO_2561 (O_2561,N_25275,N_21090);
nor UO_2562 (O_2562,N_23670,N_25896);
or UO_2563 (O_2563,N_25200,N_27870);
nand UO_2564 (O_2564,N_26939,N_25522);
nand UO_2565 (O_2565,N_29524,N_24890);
or UO_2566 (O_2566,N_20464,N_28823);
nand UO_2567 (O_2567,N_28716,N_20553);
or UO_2568 (O_2568,N_28017,N_23852);
nand UO_2569 (O_2569,N_29040,N_27998);
or UO_2570 (O_2570,N_29450,N_21681);
and UO_2571 (O_2571,N_29925,N_29759);
nand UO_2572 (O_2572,N_20855,N_22350);
nor UO_2573 (O_2573,N_23261,N_20715);
nand UO_2574 (O_2574,N_26864,N_29494);
nor UO_2575 (O_2575,N_20559,N_26123);
or UO_2576 (O_2576,N_22370,N_25529);
or UO_2577 (O_2577,N_27725,N_23936);
nand UO_2578 (O_2578,N_27577,N_25265);
nor UO_2579 (O_2579,N_28553,N_21474);
nor UO_2580 (O_2580,N_22650,N_22220);
nand UO_2581 (O_2581,N_26225,N_21219);
and UO_2582 (O_2582,N_28772,N_23992);
nand UO_2583 (O_2583,N_22251,N_20466);
or UO_2584 (O_2584,N_29563,N_21809);
nand UO_2585 (O_2585,N_21189,N_26898);
xnor UO_2586 (O_2586,N_29970,N_22523);
nor UO_2587 (O_2587,N_20081,N_29810);
nor UO_2588 (O_2588,N_23469,N_21320);
and UO_2589 (O_2589,N_28964,N_25656);
or UO_2590 (O_2590,N_28380,N_27675);
nor UO_2591 (O_2591,N_29693,N_28861);
nand UO_2592 (O_2592,N_26066,N_27584);
and UO_2593 (O_2593,N_27089,N_22511);
nor UO_2594 (O_2594,N_21579,N_21372);
and UO_2595 (O_2595,N_28152,N_24238);
and UO_2596 (O_2596,N_23113,N_24160);
nand UO_2597 (O_2597,N_26052,N_27775);
or UO_2598 (O_2598,N_20868,N_26830);
and UO_2599 (O_2599,N_24186,N_20176);
nor UO_2600 (O_2600,N_26582,N_22857);
nand UO_2601 (O_2601,N_29080,N_26200);
nor UO_2602 (O_2602,N_26103,N_28602);
or UO_2603 (O_2603,N_25811,N_23586);
nand UO_2604 (O_2604,N_21257,N_22976);
nand UO_2605 (O_2605,N_27730,N_23738);
nand UO_2606 (O_2606,N_25429,N_28647);
nor UO_2607 (O_2607,N_28313,N_21264);
nand UO_2608 (O_2608,N_29107,N_29435);
nand UO_2609 (O_2609,N_28459,N_21195);
or UO_2610 (O_2610,N_29652,N_24003);
or UO_2611 (O_2611,N_28183,N_29488);
and UO_2612 (O_2612,N_28685,N_20817);
nand UO_2613 (O_2613,N_23342,N_22813);
nor UO_2614 (O_2614,N_26249,N_21241);
and UO_2615 (O_2615,N_27194,N_27838);
or UO_2616 (O_2616,N_29201,N_25646);
or UO_2617 (O_2617,N_26970,N_20111);
and UO_2618 (O_2618,N_22631,N_22469);
nor UO_2619 (O_2619,N_23315,N_23947);
or UO_2620 (O_2620,N_28297,N_20035);
or UO_2621 (O_2621,N_26263,N_20606);
and UO_2622 (O_2622,N_26175,N_21578);
nor UO_2623 (O_2623,N_25446,N_27714);
nor UO_2624 (O_2624,N_21123,N_29416);
or UO_2625 (O_2625,N_24487,N_20793);
nor UO_2626 (O_2626,N_28154,N_21346);
nor UO_2627 (O_2627,N_24632,N_24638);
nor UO_2628 (O_2628,N_26599,N_21844);
nand UO_2629 (O_2629,N_24486,N_20661);
nand UO_2630 (O_2630,N_26456,N_26471);
nor UO_2631 (O_2631,N_28884,N_20754);
nand UO_2632 (O_2632,N_24085,N_21103);
and UO_2633 (O_2633,N_20350,N_22461);
and UO_2634 (O_2634,N_23316,N_25575);
and UO_2635 (O_2635,N_24897,N_27315);
nor UO_2636 (O_2636,N_23202,N_28004);
nand UO_2637 (O_2637,N_21060,N_21291);
nand UO_2638 (O_2638,N_21507,N_28015);
and UO_2639 (O_2639,N_27917,N_25134);
nand UO_2640 (O_2640,N_28165,N_21062);
or UO_2641 (O_2641,N_27632,N_24206);
nand UO_2642 (O_2642,N_24599,N_22641);
or UO_2643 (O_2643,N_21003,N_20915);
or UO_2644 (O_2644,N_20655,N_21245);
and UO_2645 (O_2645,N_21326,N_21719);
nand UO_2646 (O_2646,N_23575,N_22578);
nand UO_2647 (O_2647,N_27765,N_22290);
or UO_2648 (O_2648,N_20763,N_27078);
or UO_2649 (O_2649,N_29441,N_24338);
nor UO_2650 (O_2650,N_25509,N_21994);
nor UO_2651 (O_2651,N_26238,N_29993);
and UO_2652 (O_2652,N_29763,N_24725);
or UO_2653 (O_2653,N_25693,N_26973);
nand UO_2654 (O_2654,N_20726,N_20528);
nand UO_2655 (O_2655,N_23588,N_23757);
nor UO_2656 (O_2656,N_24786,N_22733);
or UO_2657 (O_2657,N_29483,N_22754);
and UO_2658 (O_2658,N_28356,N_21289);
or UO_2659 (O_2659,N_27809,N_25639);
nor UO_2660 (O_2660,N_22137,N_27339);
nand UO_2661 (O_2661,N_24201,N_25058);
and UO_2662 (O_2662,N_25892,N_22966);
nor UO_2663 (O_2663,N_23271,N_22684);
or UO_2664 (O_2664,N_25124,N_25261);
nand UO_2665 (O_2665,N_23640,N_22047);
and UO_2666 (O_2666,N_22769,N_23303);
nand UO_2667 (O_2667,N_24229,N_28101);
nand UO_2668 (O_2668,N_26155,N_24588);
nor UO_2669 (O_2669,N_20643,N_27222);
nand UO_2670 (O_2670,N_25045,N_29266);
and UO_2671 (O_2671,N_26723,N_25692);
nor UO_2672 (O_2672,N_23264,N_28471);
nand UO_2673 (O_2673,N_20138,N_27214);
or UO_2674 (O_2674,N_21374,N_22351);
and UO_2675 (O_2675,N_21806,N_25985);
nand UO_2676 (O_2676,N_24921,N_29370);
and UO_2677 (O_2677,N_22470,N_20469);
or UO_2678 (O_2678,N_21304,N_29948);
nor UO_2679 (O_2679,N_26089,N_29397);
nor UO_2680 (O_2680,N_20673,N_26539);
and UO_2681 (O_2681,N_21222,N_22083);
and UO_2682 (O_2682,N_29227,N_23971);
or UO_2683 (O_2683,N_27968,N_23894);
and UO_2684 (O_2684,N_20321,N_25425);
and UO_2685 (O_2685,N_26032,N_22681);
or UO_2686 (O_2686,N_29674,N_22245);
and UO_2687 (O_2687,N_23515,N_21067);
or UO_2688 (O_2688,N_22312,N_22271);
nor UO_2689 (O_2689,N_28156,N_24542);
or UO_2690 (O_2690,N_22487,N_28931);
and UO_2691 (O_2691,N_21701,N_22698);
and UO_2692 (O_2692,N_25539,N_24663);
nor UO_2693 (O_2693,N_22394,N_29947);
nor UO_2694 (O_2694,N_29094,N_25392);
nand UO_2695 (O_2695,N_23619,N_26202);
nor UO_2696 (O_2696,N_27046,N_27155);
and UO_2697 (O_2697,N_29205,N_22455);
nand UO_2698 (O_2698,N_23281,N_21510);
or UO_2699 (O_2699,N_24994,N_22404);
nor UO_2700 (O_2700,N_21957,N_23861);
nor UO_2701 (O_2701,N_22997,N_23225);
or UO_2702 (O_2702,N_24476,N_25001);
nand UO_2703 (O_2703,N_23482,N_29306);
nor UO_2704 (O_2704,N_24589,N_28535);
or UO_2705 (O_2705,N_26294,N_28629);
or UO_2706 (O_2706,N_26790,N_23382);
nand UO_2707 (O_2707,N_22175,N_22158);
or UO_2708 (O_2708,N_20129,N_24613);
and UO_2709 (O_2709,N_20770,N_22380);
or UO_2710 (O_2710,N_28980,N_23007);
and UO_2711 (O_2711,N_22934,N_21761);
nor UO_2712 (O_2712,N_23499,N_28833);
nand UO_2713 (O_2713,N_25562,N_28775);
nor UO_2714 (O_2714,N_22896,N_25202);
nand UO_2715 (O_2715,N_26041,N_23313);
or UO_2716 (O_2716,N_26796,N_29582);
nand UO_2717 (O_2717,N_28400,N_26493);
nand UO_2718 (O_2718,N_22236,N_28448);
nor UO_2719 (O_2719,N_20342,N_22935);
or UO_2720 (O_2720,N_28290,N_28966);
nand UO_2721 (O_2721,N_23227,N_22250);
and UO_2722 (O_2722,N_22887,N_20534);
nand UO_2723 (O_2723,N_20660,N_25559);
or UO_2724 (O_2724,N_27910,N_20937);
nor UO_2725 (O_2725,N_21303,N_22198);
and UO_2726 (O_2726,N_26000,N_23195);
nor UO_2727 (O_2727,N_21224,N_22644);
nor UO_2728 (O_2728,N_21440,N_26197);
nand UO_2729 (O_2729,N_26757,N_20863);
and UO_2730 (O_2730,N_27926,N_20860);
and UO_2731 (O_2731,N_28928,N_22687);
and UO_2732 (O_2732,N_28698,N_29574);
nor UO_2733 (O_2733,N_21248,N_25807);
or UO_2734 (O_2734,N_21882,N_21376);
or UO_2735 (O_2735,N_29155,N_21722);
and UO_2736 (O_2736,N_22623,N_20455);
and UO_2737 (O_2737,N_29679,N_23275);
and UO_2738 (O_2738,N_23434,N_24365);
nor UO_2739 (O_2739,N_25544,N_28445);
nand UO_2740 (O_2740,N_29566,N_22280);
nor UO_2741 (O_2741,N_22261,N_23233);
or UO_2742 (O_2742,N_25768,N_27150);
or UO_2743 (O_2743,N_26190,N_24278);
nand UO_2744 (O_2744,N_20837,N_23590);
xor UO_2745 (O_2745,N_20472,N_25439);
or UO_2746 (O_2746,N_27605,N_22400);
nor UO_2747 (O_2747,N_21742,N_26849);
nand UO_2748 (O_2748,N_28330,N_25659);
xor UO_2749 (O_2749,N_27556,N_28246);
nor UO_2750 (O_2750,N_22549,N_24148);
or UO_2751 (O_2751,N_28682,N_23457);
and UO_2752 (O_2752,N_29059,N_22841);
nand UO_2753 (O_2753,N_29499,N_29433);
and UO_2754 (O_2754,N_25640,N_27677);
nand UO_2755 (O_2755,N_23359,N_27478);
nor UO_2756 (O_2756,N_21585,N_24478);
nand UO_2757 (O_2757,N_25980,N_27003);
nand UO_2758 (O_2758,N_29374,N_23754);
nand UO_2759 (O_2759,N_26694,N_28147);
nor UO_2760 (O_2760,N_27595,N_25917);
or UO_2761 (O_2761,N_28523,N_25952);
or UO_2762 (O_2762,N_23480,N_26118);
and UO_2763 (O_2763,N_24228,N_28144);
nand UO_2764 (O_2764,N_23307,N_29116);
nand UO_2765 (O_2765,N_24045,N_27271);
and UO_2766 (O_2766,N_22998,N_29891);
and UO_2767 (O_2767,N_20004,N_23984);
and UO_2768 (O_2768,N_25150,N_23870);
nor UO_2769 (O_2769,N_23015,N_24312);
and UO_2770 (O_2770,N_26843,N_21111);
nand UO_2771 (O_2771,N_26447,N_25974);
or UO_2772 (O_2772,N_23291,N_24879);
nor UO_2773 (O_2773,N_20014,N_22759);
nand UO_2774 (O_2774,N_23651,N_28317);
or UO_2775 (O_2775,N_23706,N_29122);
nor UO_2776 (O_2776,N_25893,N_25420);
nand UO_2777 (O_2777,N_22741,N_24484);
xnor UO_2778 (O_2778,N_29447,N_24052);
or UO_2779 (O_2779,N_23473,N_27092);
or UO_2780 (O_2780,N_28565,N_29697);
xor UO_2781 (O_2781,N_20506,N_25781);
nand UO_2782 (O_2782,N_21119,N_22415);
nor UO_2783 (O_2783,N_25171,N_24969);
and UO_2784 (O_2784,N_22140,N_29842);
nand UO_2785 (O_2785,N_29707,N_25845);
nor UO_2786 (O_2786,N_20636,N_27932);
nor UO_2787 (O_2787,N_28509,N_23157);
xor UO_2788 (O_2788,N_20696,N_21519);
nor UO_2789 (O_2789,N_24036,N_24309);
nand UO_2790 (O_2790,N_22776,N_20476);
or UO_2791 (O_2791,N_21070,N_22099);
nand UO_2792 (O_2792,N_28119,N_28438);
nand UO_2793 (O_2793,N_23682,N_26731);
nand UO_2794 (O_2794,N_20487,N_26661);
nand UO_2795 (O_2795,N_24268,N_27951);
xnor UO_2796 (O_2796,N_24465,N_25454);
nand UO_2797 (O_2797,N_29673,N_24397);
nor UO_2798 (O_2798,N_21756,N_29298);
and UO_2799 (O_2799,N_25157,N_28089);
nor UO_2800 (O_2800,N_26972,N_20066);
or UO_2801 (O_2801,N_29347,N_20938);
and UO_2802 (O_2802,N_21438,N_28832);
nand UO_2803 (O_2803,N_27238,N_20020);
nand UO_2804 (O_2804,N_28988,N_20197);
nor UO_2805 (O_2805,N_22059,N_22788);
nor UO_2806 (O_2806,N_20869,N_29872);
and UO_2807 (O_2807,N_28000,N_26248);
nor UO_2808 (O_2808,N_21185,N_22213);
nor UO_2809 (O_2809,N_26272,N_20482);
nor UO_2810 (O_2810,N_28737,N_21815);
nand UO_2811 (O_2811,N_21803,N_29919);
and UO_2812 (O_2812,N_24870,N_22551);
and UO_2813 (O_2813,N_29431,N_27357);
nand UO_2814 (O_2814,N_21198,N_27678);
nand UO_2815 (O_2815,N_24416,N_24647);
nand UO_2816 (O_2816,N_27484,N_29882);
nor UO_2817 (O_2817,N_22874,N_22624);
or UO_2818 (O_2818,N_26215,N_29031);
or UO_2819 (O_2819,N_29650,N_21671);
nand UO_2820 (O_2820,N_26981,N_20216);
nor UO_2821 (O_2821,N_27749,N_21513);
or UO_2822 (O_2822,N_20541,N_26168);
or UO_2823 (O_2823,N_27813,N_29054);
nor UO_2824 (O_2824,N_22547,N_23707);
nand UO_2825 (O_2825,N_26722,N_27942);
and UO_2826 (O_2826,N_24061,N_20215);
nand UO_2827 (O_2827,N_28423,N_28668);
or UO_2828 (O_2828,N_22642,N_25885);
and UO_2829 (O_2829,N_24231,N_28593);
or UO_2830 (O_2830,N_22968,N_28129);
nor UO_2831 (O_2831,N_24290,N_22178);
and UO_2832 (O_2832,N_28137,N_25180);
and UO_2833 (O_2833,N_28663,N_25957);
nor UO_2834 (O_2834,N_25374,N_20305);
nand UO_2835 (O_2835,N_28206,N_27726);
nor UO_2836 (O_2836,N_23104,N_28139);
nand UO_2837 (O_2837,N_26839,N_25338);
or UO_2838 (O_2838,N_22292,N_22539);
or UO_2839 (O_2839,N_22211,N_27234);
or UO_2840 (O_2840,N_20124,N_29533);
nor UO_2841 (O_2841,N_21594,N_22743);
or UO_2842 (O_2842,N_26030,N_27616);
and UO_2843 (O_2843,N_23838,N_24907);
nand UO_2844 (O_2844,N_28874,N_24526);
xor UO_2845 (O_2845,N_23976,N_22764);
or UO_2846 (O_2846,N_29792,N_28488);
nand UO_2847 (O_2847,N_29620,N_20040);
nand UO_2848 (O_2848,N_29095,N_24281);
nand UO_2849 (O_2849,N_25878,N_29824);
nor UO_2850 (O_2850,N_23822,N_22611);
nand UO_2851 (O_2851,N_21656,N_29093);
and UO_2852 (O_2852,N_20467,N_23973);
nor UO_2853 (O_2853,N_23768,N_29858);
and UO_2854 (O_2854,N_20746,N_27760);
or UO_2855 (O_2855,N_29052,N_23062);
nand UO_2856 (O_2856,N_26683,N_28483);
nand UO_2857 (O_2857,N_23859,N_20783);
and UO_2858 (O_2858,N_27841,N_22401);
or UO_2859 (O_2859,N_28819,N_28444);
or UO_2860 (O_2860,N_21330,N_26031);
nand UO_2861 (O_2861,N_26173,N_28548);
nor UO_2862 (O_2862,N_21317,N_22216);
and UO_2863 (O_2863,N_23061,N_24637);
nand UO_2864 (O_2864,N_22078,N_22653);
nor UO_2865 (O_2865,N_25156,N_23043);
nand UO_2866 (O_2866,N_25818,N_23256);
and UO_2867 (O_2867,N_29791,N_28934);
nor UO_2868 (O_2868,N_25396,N_24154);
or UO_2869 (O_2869,N_24825,N_26997);
or UO_2870 (O_2870,N_20527,N_29342);
or UO_2871 (O_2871,N_23770,N_20785);
and UO_2872 (O_2872,N_28542,N_29465);
and UO_2873 (O_2873,N_21084,N_26578);
and UO_2874 (O_2874,N_20120,N_20311);
and UO_2875 (O_2875,N_28294,N_27763);
and UO_2876 (O_2876,N_22072,N_20494);
nand UO_2877 (O_2877,N_26417,N_26615);
nor UO_2878 (O_2878,N_27654,N_20507);
nand UO_2879 (O_2879,N_22451,N_22358);
nand UO_2880 (O_2880,N_20224,N_29025);
or UO_2881 (O_2881,N_23124,N_27012);
or UO_2882 (O_2882,N_27959,N_27505);
nand UO_2883 (O_2883,N_23031,N_24219);
or UO_2884 (O_2884,N_22306,N_27128);
and UO_2885 (O_2885,N_28684,N_26840);
nor UO_2886 (O_2886,N_21725,N_22766);
and UO_2887 (O_2887,N_26921,N_24922);
nand UO_2888 (O_2888,N_22069,N_27571);
or UO_2889 (O_2889,N_25658,N_21915);
or UO_2890 (O_2890,N_27111,N_26953);
and UO_2891 (O_2891,N_20531,N_24071);
and UO_2892 (O_2892,N_26931,N_23108);
or UO_2893 (O_2893,N_28096,N_24361);
nand UO_2894 (O_2894,N_20024,N_23910);
nand UO_2895 (O_2895,N_28472,N_21117);
nand UO_2896 (O_2896,N_24836,N_25572);
nor UO_2897 (O_2897,N_21548,N_28733);
nor UO_2898 (O_2898,N_20784,N_29664);
and UO_2899 (O_2899,N_27373,N_29958);
and UO_2900 (O_2900,N_23216,N_25394);
nor UO_2901 (O_2901,N_21193,N_25634);
or UO_2902 (O_2902,N_26540,N_20524);
or UO_2903 (O_2903,N_26671,N_27650);
nand UO_2904 (O_2904,N_28328,N_28975);
nor UO_2905 (O_2905,N_25201,N_20575);
nor UO_2906 (O_2906,N_20903,N_20433);
nand UO_2907 (O_2907,N_27697,N_20474);
nand UO_2908 (O_2908,N_27947,N_22907);
nand UO_2909 (O_2909,N_22858,N_29225);
nand UO_2910 (O_2910,N_24904,N_26472);
nand UO_2911 (O_2911,N_28301,N_21528);
and UO_2912 (O_2912,N_29621,N_20358);
and UO_2913 (O_2913,N_21017,N_20753);
nand UO_2914 (O_2914,N_23884,N_23238);
nor UO_2915 (O_2915,N_28693,N_27703);
nand UO_2916 (O_2916,N_21953,N_26077);
and UO_2917 (O_2917,N_29106,N_25334);
or UO_2918 (O_2918,N_29044,N_29553);
or UO_2919 (O_2919,N_22286,N_26852);
or UO_2920 (O_2920,N_25608,N_20440);
nand UO_2921 (O_2921,N_26977,N_27209);
nor UO_2922 (O_2922,N_27702,N_28081);
and UO_2923 (O_2923,N_20337,N_20852);
xnor UO_2924 (O_2924,N_27772,N_21203);
and UO_2925 (O_2925,N_21518,N_21973);
and UO_2926 (O_2926,N_20829,N_26467);
and UO_2927 (O_2927,N_24577,N_21908);
and UO_2928 (O_2928,N_27824,N_27156);
and UO_2929 (O_2929,N_27646,N_21530);
nor UO_2930 (O_2930,N_26574,N_29057);
or UO_2931 (O_2931,N_26258,N_24574);
nor UO_2932 (O_2932,N_25976,N_23443);
nand UO_2933 (O_2933,N_23761,N_22726);
and UO_2934 (O_2934,N_23798,N_24023);
nand UO_2935 (O_2935,N_28253,N_28803);
nor UO_2936 (O_2936,N_21752,N_22024);
nor UO_2937 (O_2937,N_25192,N_20000);
nand UO_2938 (O_2938,N_27259,N_27058);
nand UO_2939 (O_2939,N_24224,N_20733);
and UO_2940 (O_2940,N_20932,N_29330);
nor UO_2941 (O_2941,N_26298,N_28588);
or UO_2942 (O_2942,N_24055,N_28713);
or UO_2943 (O_2943,N_20385,N_26611);
or UO_2944 (O_2944,N_23001,N_20900);
and UO_2945 (O_2945,N_27167,N_26596);
or UO_2946 (O_2946,N_20363,N_20205);
or UO_2947 (O_2947,N_29702,N_29332);
nand UO_2948 (O_2948,N_26867,N_22215);
or UO_2949 (O_2949,N_21138,N_27685);
nor UO_2950 (O_2950,N_25229,N_29603);
and UO_2951 (O_2951,N_24009,N_21923);
and UO_2952 (O_2952,N_22695,N_21407);
nor UO_2953 (O_2953,N_28703,N_24717);
or UO_2954 (O_2954,N_25393,N_21911);
nor UO_2955 (O_2955,N_22774,N_28337);
or UO_2956 (O_2956,N_24173,N_20975);
nand UO_2957 (O_2957,N_23885,N_29575);
or UO_2958 (O_2958,N_23058,N_21116);
or UO_2959 (O_2959,N_23189,N_23345);
nand UO_2960 (O_2960,N_21261,N_26101);
or UO_2961 (O_2961,N_21006,N_24555);
or UO_2962 (O_2962,N_20323,N_29369);
or UO_2963 (O_2963,N_20532,N_27930);
and UO_2964 (O_2964,N_20518,N_21462);
nor UO_2965 (O_2965,N_23022,N_28859);
and UO_2966 (O_2966,N_23134,N_23891);
and UO_2967 (O_2967,N_20462,N_22308);
or UO_2968 (O_2968,N_26537,N_22990);
and UO_2969 (O_2969,N_23046,N_27984);
or UO_2970 (O_2970,N_27438,N_29541);
nor UO_2971 (O_2971,N_24183,N_29705);
nor UO_2972 (O_2972,N_22282,N_23818);
nor UO_2973 (O_2973,N_29220,N_27191);
and UO_2974 (O_2974,N_23865,N_20354);
nand UO_2975 (O_2975,N_22426,N_29123);
and UO_2976 (O_2976,N_27242,N_24479);
or UO_2977 (O_2977,N_20775,N_29501);
and UO_2978 (O_2978,N_29802,N_20367);
nand UO_2979 (O_2979,N_23380,N_29830);
and UO_2980 (O_2980,N_29470,N_28747);
nor UO_2981 (O_2981,N_21865,N_29323);
nand UO_2982 (O_2982,N_20499,N_22307);
nand UO_2983 (O_2983,N_21007,N_28187);
or UO_2984 (O_2984,N_29042,N_29421);
nor UO_2985 (O_2985,N_27695,N_29175);
nand UO_2986 (O_2986,N_20067,N_22160);
and UO_2987 (O_2987,N_28223,N_21435);
and UO_2988 (O_2988,N_22674,N_28002);
nor UO_2989 (O_2989,N_24443,N_27614);
nor UO_2990 (O_2990,N_25600,N_27424);
or UO_2991 (O_2991,N_23558,N_20079);
nor UO_2992 (O_2992,N_26809,N_21318);
and UO_2993 (O_2993,N_28436,N_25064);
nor UO_2994 (O_2994,N_24760,N_21393);
or UO_2995 (O_2995,N_26164,N_28378);
nor UO_2996 (O_2996,N_29398,N_21057);
nand UO_2997 (O_2997,N_28826,N_21322);
and UO_2998 (O_2998,N_20387,N_20510);
or UO_2999 (O_2999,N_28626,N_23521);
nand UO_3000 (O_3000,N_27692,N_25644);
nor UO_3001 (O_3001,N_21089,N_23160);
and UO_3002 (O_3002,N_24602,N_26891);
nand UO_3003 (O_3003,N_23571,N_24431);
or UO_3004 (O_3004,N_26018,N_21679);
nor UO_3005 (O_3005,N_21645,N_23335);
and UO_3006 (O_3006,N_29601,N_22120);
nand UO_3007 (O_3007,N_23389,N_28403);
or UO_3008 (O_3008,N_24203,N_28750);
and UO_3009 (O_3009,N_29699,N_25224);
and UO_3010 (O_3010,N_23122,N_21213);
nand UO_3011 (O_3011,N_26804,N_28425);
and UO_3012 (O_3012,N_23034,N_24609);
and UO_3013 (O_3013,N_27226,N_25411);
nand UO_3014 (O_3014,N_23069,N_26205);
nor UO_3015 (O_3015,N_25520,N_21412);
nor UO_3016 (O_3016,N_29844,N_26579);
nor UO_3017 (O_3017,N_26362,N_27173);
nor UO_3018 (O_3018,N_21812,N_28918);
or UO_3019 (O_3019,N_21265,N_24430);
and UO_3020 (O_3020,N_28190,N_27782);
nand UO_3021 (O_3021,N_29586,N_28363);
and UO_3022 (O_3022,N_21822,N_26747);
nand UO_3023 (O_3023,N_26755,N_20087);
nor UO_3024 (O_3024,N_24150,N_25990);
xor UO_3025 (O_3025,N_28326,N_27443);
or UO_3026 (O_3026,N_21634,N_23232);
and UO_3027 (O_3027,N_20225,N_28746);
and UO_3028 (O_3028,N_21327,N_26545);
nand UO_3029 (O_3029,N_22166,N_20392);
or UO_3030 (O_3030,N_29913,N_21871);
or UO_3031 (O_3031,N_23072,N_26402);
and UO_3032 (O_3032,N_27877,N_22309);
and UO_3033 (O_3033,N_25744,N_20194);
or UO_3034 (O_3034,N_29992,N_26618);
nand UO_3035 (O_3035,N_29658,N_24895);
or UO_3036 (O_3036,N_20239,N_27660);
and UO_3037 (O_3037,N_24634,N_23621);
and UO_3038 (O_3038,N_27506,N_24283);
or UO_3039 (O_3039,N_24543,N_27015);
or UO_3040 (O_3040,N_29480,N_27278);
nand UO_3041 (O_3041,N_29526,N_27129);
nor UO_3042 (O_3042,N_29443,N_24404);
or UO_3043 (O_3043,N_28897,N_24121);
nor UO_3044 (O_3044,N_20930,N_26920);
nand UO_3045 (O_3045,N_25155,N_24798);
and UO_3046 (O_3046,N_26204,N_28288);
and UO_3047 (O_3047,N_23188,N_21667);
nand UO_3048 (O_3048,N_21277,N_28485);
nor UO_3049 (O_3049,N_24077,N_22385);
nand UO_3050 (O_3050,N_22248,N_28686);
nor UO_3051 (O_3051,N_23887,N_29098);
nor UO_3052 (O_3052,N_22356,N_20051);
nand UO_3053 (O_3053,N_22353,N_28719);
nor UO_3054 (O_3054,N_29789,N_22207);
or UO_3055 (O_3055,N_21223,N_23805);
or UO_3056 (O_3056,N_24957,N_22098);
and UO_3057 (O_3057,N_24310,N_24508);
nand UO_3058 (O_3058,N_21963,N_28843);
xor UO_3059 (O_3059,N_25637,N_25577);
nor UO_3060 (O_3060,N_27674,N_24761);
or UO_3061 (O_3061,N_25367,N_29278);
nand UO_3062 (O_3062,N_23268,N_28176);
nor UO_3063 (O_3063,N_24428,N_24175);
and UO_3064 (O_3064,N_24846,N_29402);
and UO_3065 (O_3065,N_29626,N_20074);
nor UO_3066 (O_3066,N_22063,N_20856);
nor UO_3067 (O_3067,N_24565,N_22007);
or UO_3068 (O_3068,N_26816,N_20048);
or UO_3069 (O_3069,N_25147,N_22264);
or UO_3070 (O_3070,N_21124,N_29952);
nand UO_3071 (O_3071,N_24541,N_21397);
nand UO_3072 (O_3072,N_20543,N_24189);
and UO_3073 (O_3073,N_25906,N_22603);
nor UO_3074 (O_3074,N_26746,N_20190);
nand UO_3075 (O_3075,N_27993,N_23300);
and UO_3076 (O_3076,N_25252,N_29178);
nor UO_3077 (O_3077,N_23843,N_28071);
or UO_3078 (O_3078,N_29273,N_29772);
nand UO_3079 (O_3079,N_23604,N_25830);
and UO_3080 (O_3080,N_24450,N_23988);
or UO_3081 (O_3081,N_28310,N_26850);
and UO_3082 (O_3082,N_23330,N_27294);
nand UO_3083 (O_3083,N_26529,N_20357);
or UO_3084 (O_3084,N_20752,N_21614);
or UO_3085 (O_3085,N_27395,N_21395);
nor UO_3086 (O_3086,N_28534,N_27190);
and UO_3087 (O_3087,N_27802,N_21236);
and UO_3088 (O_3088,N_29104,N_27411);
nor UO_3089 (O_3089,N_26913,N_28167);
or UO_3090 (O_3090,N_28968,N_26935);
or UO_3091 (O_3091,N_25867,N_25556);
and UO_3092 (O_3092,N_21328,N_27376);
nor UO_3093 (O_3093,N_25651,N_28611);
or UO_3094 (O_3094,N_21555,N_27247);
nor UO_3095 (O_3095,N_20171,N_22933);
and UO_3096 (O_3096,N_26894,N_21023);
and UO_3097 (O_3097,N_22926,N_28661);
or UO_3098 (O_3098,N_27449,N_20317);
nand UO_3099 (O_3099,N_24641,N_25225);
and UO_3100 (O_3100,N_22995,N_25747);
nor UO_3101 (O_3101,N_21713,N_26228);
or UO_3102 (O_3102,N_24360,N_28405);
or UO_3103 (O_3103,N_24032,N_28370);
and UO_3104 (O_3104,N_26527,N_22053);
nor UO_3105 (O_3105,N_25190,N_22601);
nor UO_3106 (O_3106,N_28327,N_27588);
and UO_3107 (O_3107,N_21083,N_22283);
and UO_3108 (O_3108,N_27352,N_20054);
nor UO_3109 (O_3109,N_26307,N_28579);
nor UO_3110 (O_3110,N_27014,N_24690);
and UO_3111 (O_3111,N_23834,N_20488);
or UO_3112 (O_3112,N_23776,N_24514);
and UO_3113 (O_3113,N_25620,N_27896);
and UO_3114 (O_3114,N_25430,N_27210);
and UO_3115 (O_3115,N_21737,N_22589);
or UO_3116 (O_3116,N_24956,N_20981);
and UO_3117 (O_3117,N_24311,N_28045);
and UO_3118 (O_3118,N_28904,N_29778);
nand UO_3119 (O_3119,N_20227,N_22011);
nor UO_3120 (O_3120,N_29186,N_25222);
or UO_3121 (O_3121,N_21039,N_23783);
nand UO_3122 (O_3122,N_29279,N_27225);
nor UO_3123 (O_3123,N_28118,N_28683);
nor UO_3124 (O_3124,N_26036,N_20336);
nand UO_3125 (O_3125,N_27063,N_21533);
nand UO_3126 (O_3126,N_20406,N_23016);
nand UO_3127 (O_3127,N_23339,N_20969);
nand UO_3128 (O_3128,N_20276,N_28470);
and UO_3129 (O_3129,N_26310,N_29760);
nand UO_3130 (O_3130,N_24464,N_25233);
nor UO_3131 (O_3131,N_23803,N_24559);
or UO_3132 (O_3132,N_23119,N_26949);
nand UO_3133 (O_3133,N_23642,N_20828);
and UO_3134 (O_3134,N_21783,N_24316);
nor UO_3135 (O_3135,N_21130,N_24727);
and UO_3136 (O_3136,N_23012,N_25269);
or UO_3137 (O_3137,N_21276,N_24841);
and UO_3138 (O_3138,N_24192,N_29268);
nor UO_3139 (O_3139,N_27272,N_26620);
and UO_3140 (O_3140,N_24247,N_27295);
nor UO_3141 (O_3141,N_24060,N_27794);
and UO_3142 (O_3142,N_27007,N_27658);
nor UO_3143 (O_3143,N_26406,N_24130);
or UO_3144 (O_3144,N_29906,N_21566);
or UO_3145 (O_3145,N_22061,N_21444);
nor UO_3146 (O_3146,N_27291,N_27062);
nor UO_3147 (O_3147,N_25119,N_28941);
or UO_3148 (O_3148,N_27077,N_22872);
or UO_3149 (O_3149,N_26626,N_23672);
nor UO_3150 (O_3150,N_27413,N_29805);
nand UO_3151 (O_3151,N_28257,N_25855);
nor UO_3152 (O_3152,N_22649,N_25948);
nand UO_3153 (O_3153,N_20879,N_29291);
or UO_3154 (O_3154,N_25315,N_20789);
nor UO_3155 (O_3155,N_27397,N_29981);
nor UO_3156 (O_3156,N_29757,N_22303);
or UO_3157 (O_3157,N_29401,N_24538);
or UO_3158 (O_3158,N_29003,N_22262);
or UO_3159 (O_3159,N_20005,N_22444);
nor UO_3160 (O_3160,N_21373,N_24126);
and UO_3161 (O_3161,N_20088,N_22862);
xor UO_3162 (O_3162,N_28108,N_22553);
or UO_3163 (O_3163,N_25125,N_26159);
or UO_3164 (O_3164,N_29703,N_24858);
or UO_3165 (O_3165,N_29159,N_20047);
and UO_3166 (O_3166,N_21845,N_22490);
or UO_3167 (O_3167,N_25047,N_22021);
nor UO_3168 (O_3168,N_28067,N_26872);
and UO_3169 (O_3169,N_24256,N_25636);
nand UO_3170 (O_3170,N_28900,N_23549);
nand UO_3171 (O_3171,N_26535,N_29294);
nand UO_3172 (O_3172,N_22571,N_28566);
or UO_3173 (O_3173,N_22805,N_22089);
nand UO_3174 (O_3174,N_28018,N_29971);
nor UO_3175 (O_3175,N_28740,N_21943);
nand UO_3176 (O_3176,N_20348,N_26701);
or UO_3177 (O_3177,N_26252,N_23546);
nand UO_3178 (O_3178,N_28086,N_28305);
and UO_3179 (O_3179,N_29016,N_29939);
nand UO_3180 (O_3180,N_27925,N_22315);
or UO_3181 (O_3181,N_24062,N_28742);
nor UO_3182 (O_3182,N_29079,N_29056);
nor UO_3183 (O_3183,N_26393,N_24512);
and UO_3184 (O_3184,N_28465,N_26470);
nand UO_3185 (O_3185,N_23953,N_29624);
and UO_3186 (O_3186,N_25759,N_24575);
and UO_3187 (O_3187,N_23107,N_25805);
or UO_3188 (O_3188,N_29437,N_27812);
or UO_3189 (O_3189,N_20154,N_20891);
nor UO_3190 (O_3190,N_26900,N_21353);
and UO_3191 (O_3191,N_20848,N_23913);
or UO_3192 (O_3192,N_25091,N_20070);
nor UO_3193 (O_3193,N_27263,N_25236);
and UO_3194 (O_3194,N_26002,N_21790);
and UO_3195 (O_3195,N_21881,N_27179);
and UO_3196 (O_3196,N_27198,N_25035);
and UO_3197 (O_3197,N_28050,N_23255);
or UO_3198 (O_3198,N_26557,N_22375);
nor UO_3199 (O_3199,N_26938,N_21262);
xnor UO_3200 (O_3200,N_27567,N_20360);
nor UO_3201 (O_3201,N_24744,N_23653);
or UO_3202 (O_3202,N_21270,N_20233);
nand UO_3203 (O_3203,N_24872,N_27047);
or UO_3204 (O_3204,N_24875,N_26512);
or UO_3205 (O_3205,N_27855,N_27644);
nor UO_3206 (O_3206,N_29619,N_20316);
xnor UO_3207 (O_3207,N_29300,N_22530);
nand UO_3208 (O_3208,N_26286,N_23676);
and UO_3209 (O_3209,N_29142,N_29006);
and UO_3210 (O_3210,N_24950,N_26343);
nor UO_3211 (O_3211,N_21423,N_25316);
nand UO_3212 (O_3212,N_21351,N_23228);
and UO_3213 (O_3213,N_28766,N_25179);
or UO_3214 (O_3214,N_22828,N_27369);
nand UO_3215 (O_3215,N_20493,N_25668);
and UO_3216 (O_3216,N_26446,N_21919);
nand UO_3217 (O_3217,N_21026,N_26678);
or UO_3218 (O_3218,N_28309,N_26108);
or UO_3219 (O_3219,N_23101,N_23096);
or UO_3220 (O_3220,N_24963,N_20624);
nor UO_3221 (O_3221,N_28714,N_26163);
nand UO_3222 (O_3222,N_21253,N_26968);
or UO_3223 (O_3223,N_25766,N_24226);
nor UO_3224 (O_3224,N_27054,N_20859);
and UO_3225 (O_3225,N_25785,N_20880);
nand UO_3226 (O_3226,N_22359,N_20641);
nor UO_3227 (O_3227,N_26600,N_25971);
nor UO_3228 (O_3228,N_22068,N_28003);
or UO_3229 (O_3229,N_28083,N_22420);
and UO_3230 (O_3230,N_27826,N_26267);
nor UO_3231 (O_3231,N_28135,N_21633);
nor UO_3232 (O_3232,N_24958,N_27024);
and UO_3233 (O_3233,N_21136,N_20294);
nor UO_3234 (O_3234,N_22294,N_27318);
nand UO_3235 (O_3235,N_25183,N_20895);
nand UO_3236 (O_3236,N_21025,N_27051);
or UO_3237 (O_3237,N_27665,N_26408);
and UO_3238 (O_3238,N_28441,N_21582);
nor UO_3239 (O_3239,N_23756,N_21597);
and UO_3240 (O_3240,N_25661,N_22518);
nor UO_3241 (O_3241,N_20745,N_20118);
or UO_3242 (O_3242,N_20627,N_24703);
nor UO_3243 (O_3243,N_25293,N_23496);
or UO_3244 (O_3244,N_22867,N_26724);
and UO_3245 (O_3245,N_29392,N_25946);
nand UO_3246 (O_3246,N_27574,N_20652);
nor UO_3247 (O_3247,N_26340,N_21441);
and UO_3248 (O_3248,N_29510,N_25386);
or UO_3249 (O_3249,N_28039,N_25825);
or UO_3250 (O_3250,N_26558,N_23613);
or UO_3251 (O_3251,N_27237,N_28192);
or UO_3252 (O_3252,N_29951,N_28695);
nor UO_3253 (O_3253,N_20503,N_25824);
or UO_3254 (O_3254,N_21139,N_20168);
nor UO_3255 (O_3255,N_28638,N_22229);
or UO_3256 (O_3256,N_26914,N_26099);
nand UO_3257 (O_3257,N_23417,N_22100);
and UO_3258 (O_3258,N_22796,N_25612);
and UO_3259 (O_3259,N_22509,N_22239);
nor UO_3260 (O_3260,N_25739,N_24640);
nor UO_3261 (O_3261,N_29329,N_26383);
nand UO_3262 (O_3262,N_27410,N_20137);
or UO_3263 (O_3263,N_22188,N_21071);
or UO_3264 (O_3264,N_21012,N_28398);
and UO_3265 (O_3265,N_23806,N_20951);
nand UO_3266 (O_3266,N_24721,N_26829);
nand UO_3267 (O_3267,N_23347,N_20781);
and UO_3268 (O_3268,N_29265,N_27773);
and UO_3269 (O_3269,N_29537,N_26616);
nor UO_3270 (O_3270,N_23229,N_25835);
and UO_3271 (O_3271,N_23384,N_21649);
nand UO_3272 (O_3272,N_29423,N_23815);
nand UO_3273 (O_3273,N_29455,N_22991);
and UO_3274 (O_3274,N_26138,N_22185);
or UO_3275 (O_3275,N_28678,N_29165);
nand UO_3276 (O_3276,N_20065,N_28461);
nor UO_3277 (O_3277,N_23702,N_27962);
or UO_3278 (O_3278,N_26309,N_21868);
nor UO_3279 (O_3279,N_25992,N_20101);
and UO_3280 (O_3280,N_24711,N_22091);
and UO_3281 (O_3281,N_25858,N_20425);
or UO_3282 (O_3282,N_28322,N_27432);
or UO_3283 (O_3283,N_28175,N_29078);
and UO_3284 (O_3284,N_27748,N_21576);
or UO_3285 (O_3285,N_25203,N_28159);
nor UO_3286 (O_3286,N_26862,N_20563);
or UO_3287 (O_3287,N_24263,N_22954);
nand UO_3288 (O_3288,N_28632,N_26662);
and UO_3289 (O_3289,N_21415,N_29091);
and UO_3290 (O_3290,N_21852,N_21906);
and UO_3291 (O_3291,N_22670,N_25103);
nand UO_3292 (O_3292,N_27591,N_27258);
nor UO_3293 (O_3293,N_23663,N_24305);
nand UO_3294 (O_3294,N_25213,N_23740);
or UO_3295 (O_3295,N_29223,N_26984);
and UO_3296 (O_3296,N_21356,N_28852);
or UO_3297 (O_3297,N_29688,N_24411);
and UO_3298 (O_3298,N_26369,N_28242);
nand UO_3299 (O_3299,N_27493,N_21998);
and UO_3300 (O_3300,N_25621,N_22563);
or UO_3301 (O_3301,N_25671,N_21842);
or UO_3302 (O_3302,N_29264,N_22112);
nor UO_3303 (O_3303,N_25357,N_21416);
nor UO_3304 (O_3304,N_23153,N_22474);
nor UO_3305 (O_3305,N_29373,N_29005);
nor UO_3306 (O_3306,N_22696,N_27313);
nor UO_3307 (O_3307,N_20782,N_24998);
or UO_3308 (O_3308,N_24540,N_24718);
and UO_3309 (O_3309,N_28306,N_25546);
and UO_3310 (O_3310,N_20075,N_20050);
and UO_3311 (O_3311,N_24402,N_21873);
nor UO_3312 (O_3312,N_24566,N_24653);
or UO_3313 (O_3313,N_25290,N_21874);
or UO_3314 (O_3314,N_22751,N_27011);
nand UO_3315 (O_3315,N_26409,N_28592);
and UO_3316 (O_3316,N_20454,N_23497);
nand UO_3317 (O_3317,N_26518,N_21151);
or UO_3318 (O_3318,N_27786,N_20724);
and UO_3319 (O_3319,N_28507,N_20470);
nand UO_3320 (O_3320,N_23779,N_20435);
and UO_3321 (O_3321,N_26119,N_25977);
or UO_3322 (O_3322,N_28075,N_23808);
nand UO_3323 (O_3323,N_24811,N_22161);
or UO_3324 (O_3324,N_29539,N_24445);
nand UO_3325 (O_3325,N_20412,N_28331);
nor UO_3326 (O_3326,N_25403,N_22980);
nand UO_3327 (O_3327,N_22327,N_22701);
and UO_3328 (O_3328,N_26445,N_29004);
nor UO_3329 (O_3329,N_26978,N_22254);
nand UO_3330 (O_3330,N_28824,N_20799);
nor UO_3331 (O_3331,N_28041,N_24925);
and UO_3332 (O_3332,N_25844,N_25271);
or UO_3333 (O_3333,N_27426,N_21735);
nand UO_3334 (O_3334,N_29750,N_29942);
or UO_3335 (O_3335,N_22719,N_26439);
nor UO_3336 (O_3336,N_23940,N_20480);
nor UO_3337 (O_3337,N_25799,N_24459);
nand UO_3338 (O_3338,N_20777,N_25718);
and UO_3339 (O_3339,N_27871,N_29551);
nand UO_3340 (O_3340,N_26455,N_27667);
nor UO_3341 (O_3341,N_21744,N_25351);
or UO_3342 (O_3342,N_25247,N_20835);
nand UO_3343 (O_3343,N_21092,N_29590);
nor UO_3344 (O_3344,N_27805,N_26039);
and UO_3345 (O_3345,N_27569,N_21428);
or UO_3346 (O_3346,N_26454,N_29554);
nand UO_3347 (O_3347,N_21929,N_26322);
nand UO_3348 (O_3348,N_27264,N_24661);
and UO_3349 (O_3349,N_22737,N_21791);
nand UO_3350 (O_3350,N_28990,N_25886);
nor UO_3351 (O_3351,N_28580,N_20923);
and UO_3352 (O_3352,N_29099,N_20477);
nand UO_3353 (O_3353,N_27381,N_27474);
and UO_3354 (O_3354,N_20836,N_29058);
and UO_3355 (O_3355,N_25424,N_25721);
nand UO_3356 (O_3356,N_21801,N_22136);
nand UO_3357 (O_3357,N_26749,N_27131);
and UO_3358 (O_3358,N_24480,N_23057);
nand UO_3359 (O_3359,N_29918,N_22152);
nand UO_3360 (O_3360,N_25942,N_25254);
or UO_3361 (O_3361,N_23223,N_26253);
nor UO_3362 (O_3362,N_26055,N_24249);
or UO_3363 (O_3363,N_21135,N_27073);
nand UO_3364 (O_3364,N_26915,N_20214);
or UO_3365 (O_3365,N_20345,N_27296);
or UO_3366 (O_3366,N_28226,N_26182);
and UO_3367 (O_3367,N_23178,N_28827);
nand UO_3368 (O_3368,N_23064,N_23356);
xnor UO_3369 (O_3369,N_22922,N_22203);
nand UO_3370 (O_3370,N_29787,N_28519);
or UO_3371 (O_3371,N_25433,N_22864);
and UO_3372 (O_3372,N_29459,N_28024);
nand UO_3373 (O_3373,N_21883,N_21260);
and UO_3374 (O_3374,N_27220,N_25178);
and UO_3375 (O_3375,N_28431,N_21573);
and UO_3376 (O_3376,N_25237,N_29523);
or UO_3377 (O_3377,N_29980,N_22700);
or UO_3378 (O_3378,N_20498,N_27330);
nor UO_3379 (O_3379,N_26333,N_21190);
nand UO_3380 (O_3380,N_21926,N_22319);
and UO_3381 (O_3381,N_22625,N_20515);
and UO_3382 (O_3382,N_26465,N_24000);
and UO_3383 (O_3383,N_26504,N_28728);
nor UO_3384 (O_3384,N_24923,N_27067);
nor UO_3385 (O_3385,N_27934,N_25911);
or UO_3386 (O_3386,N_21009,N_27898);
nand UO_3387 (O_3387,N_20614,N_27797);
or UO_3388 (O_3388,N_24294,N_26380);
or UO_3389 (O_3389,N_20397,N_27417);
nand UO_3390 (O_3390,N_27727,N_21765);
nand UO_3391 (O_3391,N_25094,N_22134);
nand UO_3392 (O_3392,N_25965,N_24915);
or UO_3393 (O_3393,N_27402,N_29256);
nand UO_3394 (O_3394,N_23892,N_25614);
or UO_3395 (O_3395,N_27872,N_26479);
nand UO_3396 (O_3396,N_22106,N_23960);
or UO_3397 (O_3397,N_23655,N_20714);
or UO_3398 (O_3398,N_21581,N_20747);
nor UO_3399 (O_3399,N_25056,N_23218);
and UO_3400 (O_3400,N_20513,N_23146);
nor UO_3401 (O_3401,N_29482,N_22714);
nand UO_3402 (O_3402,N_28146,N_20106);
and UO_3403 (O_3403,N_22009,N_20280);
nor UO_3404 (O_3404,N_25451,N_26437);
nor UO_3405 (O_3405,N_20281,N_20941);
nand UO_3406 (O_3406,N_25051,N_23519);
nor UO_3407 (O_3407,N_25164,N_27467);
nor UO_3408 (O_3408,N_25913,N_20599);
nand UO_3409 (O_3409,N_23112,N_27911);
nand UO_3410 (O_3410,N_22173,N_28179);
or UO_3411 (O_3411,N_23465,N_25758);
nor UO_3412 (O_3412,N_23725,N_23030);
or UO_3413 (O_3413,N_26330,N_21040);
and UO_3414 (O_3414,N_24202,N_23208);
nand UO_3415 (O_3415,N_29991,N_26837);
nand UO_3416 (O_3416,N_20670,N_28887);
nor UO_3417 (O_3417,N_22755,N_29974);
or UO_3418 (O_3418,N_29901,N_24579);
or UO_3419 (O_3419,N_29737,N_20148);
and UO_3420 (O_3420,N_29282,N_29606);
or UO_3421 (O_3421,N_24488,N_21836);
nand UO_3422 (O_3422,N_26317,N_20898);
nand UO_3423 (O_3423,N_23431,N_24087);
or UO_3424 (O_3424,N_21182,N_20375);
or UO_3425 (O_3425,N_24605,N_20896);
nor UO_3426 (O_3426,N_27268,N_24681);
and UO_3427 (O_3427,N_23635,N_28295);
nor UO_3428 (O_3428,N_28201,N_20651);
nor UO_3429 (O_3429,N_26609,N_21244);
nand UO_3430 (O_3430,N_25082,N_26487);
and UO_3431 (O_3431,N_22827,N_26329);
nand UO_3432 (O_3432,N_28150,N_20838);
nand UO_3433 (O_3433,N_22894,N_26029);
or UO_3434 (O_3434,N_27312,N_24554);
nand UO_3435 (O_3435,N_28021,N_20533);
nor UO_3436 (O_3436,N_23650,N_29753);
nand UO_3437 (O_3437,N_28802,N_24795);
nand UO_3438 (O_3438,N_25055,N_22875);
nor UO_3439 (O_3439,N_27564,N_28813);
nand UO_3440 (O_3440,N_21400,N_25100);
nand UO_3441 (O_3441,N_27842,N_23577);
or UO_3442 (O_3442,N_22712,N_23140);
nor UO_3443 (O_3443,N_24791,N_24982);
nor UO_3444 (O_3444,N_29389,N_25142);
or UO_3445 (O_3445,N_27592,N_20703);
nor UO_3446 (O_3446,N_26947,N_27010);
nor UO_3447 (O_3447,N_24622,N_23657);
nand UO_3448 (O_3448,N_23831,N_23165);
nand UO_3449 (O_3449,N_22919,N_23708);
or UO_3450 (O_3450,N_24646,N_24702);
nand UO_3451 (O_3451,N_22088,N_29331);
or UO_3452 (O_3452,N_21989,N_23582);
and UO_3453 (O_3453,N_20778,N_27852);
nand UO_3454 (O_3454,N_26543,N_23308);
nor UO_3455 (O_3455,N_24172,N_27860);
nand UO_3456 (O_3456,N_27487,N_26734);
and UO_3457 (O_3457,N_25810,N_24144);
nor UO_3458 (O_3458,N_25440,N_25503);
and UO_3459 (O_3459,N_29338,N_29075);
nor UO_3460 (O_3460,N_21711,N_29357);
nor UO_3461 (O_3461,N_26992,N_28212);
and UO_3462 (O_3462,N_26468,N_24293);
nand UO_3463 (O_3463,N_21179,N_26989);
nor UO_3464 (O_3464,N_29857,N_23596);
and UO_3465 (O_3465,N_20741,N_21235);
and UO_3466 (O_3466,N_20521,N_26480);
nor UO_3467 (O_3467,N_21296,N_20019);
nand UO_3468 (O_3468,N_27517,N_22605);
and UO_3469 (O_3469,N_25387,N_28993);
nor UO_3470 (O_3470,N_22911,N_26008);
and UO_3471 (O_3471,N_27119,N_26680);
nand UO_3472 (O_3472,N_29838,N_27217);
and UO_3473 (O_3473,N_26187,N_21702);
nor UO_3474 (O_3474,N_23357,N_28516);
nor UO_3475 (O_3475,N_27267,N_21979);
nor UO_3476 (O_3476,N_23398,N_28256);
nand UO_3477 (O_3477,N_25859,N_25736);
nor UO_3478 (O_3478,N_20284,N_28950);
nor UO_3479 (O_3479,N_22536,N_20287);
or UO_3480 (O_3480,N_25216,N_20003);
or UO_3481 (O_3481,N_20792,N_22671);
nand UO_3482 (O_3482,N_29678,N_29317);
and UO_3483 (O_3483,N_22243,N_24704);
or UO_3484 (O_3484,N_27384,N_26886);
and UO_3485 (O_3485,N_21946,N_22527);
nand UO_3486 (O_3486,N_28475,N_29848);
and UO_3487 (O_3487,N_21422,N_27883);
or UO_3488 (O_3488,N_29530,N_26460);
nand UO_3489 (O_3489,N_28954,N_26222);
nor UO_3490 (O_3490,N_25176,N_25127);
and UO_3491 (O_3491,N_21170,N_20623);
nor UO_3492 (O_3492,N_22534,N_27937);
and UO_3493 (O_3493,N_20960,N_27764);
or UO_3494 (O_3494,N_21587,N_25353);
or UO_3495 (O_3495,N_21666,N_22360);
nand UO_3496 (O_3496,N_28651,N_24437);
or UO_3497 (O_3497,N_22379,N_23823);
nand UO_3498 (O_3498,N_22159,N_23905);
nor UO_3499 (O_3499,N_20983,N_24359);
endmodule