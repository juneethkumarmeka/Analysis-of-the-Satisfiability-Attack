module basic_500_3000_500_30_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_245,In_131);
nand U1 (N_1,In_498,In_26);
or U2 (N_2,In_120,In_417);
and U3 (N_3,In_239,In_449);
or U4 (N_4,In_268,In_375);
xnor U5 (N_5,In_200,In_250);
or U6 (N_6,In_353,In_297);
and U7 (N_7,In_187,In_147);
and U8 (N_8,In_118,In_56);
nor U9 (N_9,In_448,In_179);
nand U10 (N_10,In_457,In_40);
nand U11 (N_11,In_264,In_48);
xnor U12 (N_12,In_57,In_292);
or U13 (N_13,In_153,In_441);
nand U14 (N_14,In_16,In_46);
and U15 (N_15,In_188,In_267);
and U16 (N_16,In_15,In_451);
nand U17 (N_17,In_128,In_154);
nor U18 (N_18,In_226,In_318);
nand U19 (N_19,In_143,In_204);
or U20 (N_20,In_404,In_175);
xnor U21 (N_21,In_377,In_376);
or U22 (N_22,In_446,In_371);
xor U23 (N_23,In_132,In_97);
xor U24 (N_24,In_274,In_423);
xor U25 (N_25,In_389,In_386);
or U26 (N_26,In_412,In_340);
and U27 (N_27,In_112,In_61);
nand U28 (N_28,In_430,In_462);
nor U29 (N_29,In_432,In_69);
nand U30 (N_30,In_45,In_345);
and U31 (N_31,In_18,In_477);
or U32 (N_32,In_144,In_214);
and U33 (N_33,In_124,In_436);
nand U34 (N_34,In_84,In_265);
xnor U35 (N_35,In_31,In_181);
nand U36 (N_36,In_332,In_140);
xnor U37 (N_37,In_8,In_89);
nand U38 (N_38,In_300,In_230);
xor U39 (N_39,In_242,In_355);
nor U40 (N_40,In_481,In_295);
xnor U41 (N_41,In_433,In_344);
or U42 (N_42,In_400,In_72);
xor U43 (N_43,In_485,In_74);
xor U44 (N_44,In_170,In_174);
nand U45 (N_45,In_58,In_468);
and U46 (N_46,In_201,In_497);
nand U47 (N_47,In_195,In_305);
nor U48 (N_48,In_308,In_456);
xnor U49 (N_49,In_416,In_447);
nor U50 (N_50,In_454,In_161);
nor U51 (N_51,In_299,In_329);
or U52 (N_52,In_5,In_455);
xnor U53 (N_53,In_306,In_10);
xnor U54 (N_54,In_360,In_32);
or U55 (N_55,In_358,In_190);
xnor U56 (N_56,In_166,In_491);
nand U57 (N_57,In_252,In_285);
or U58 (N_58,In_11,In_428);
xor U59 (N_59,In_328,In_396);
nor U60 (N_60,In_445,In_341);
nor U61 (N_61,In_293,In_348);
nor U62 (N_62,In_343,In_434);
nand U63 (N_63,In_439,In_381);
or U64 (N_64,In_492,In_487);
nor U65 (N_65,In_60,In_176);
xnor U66 (N_66,In_14,In_374);
or U67 (N_67,In_68,In_387);
and U68 (N_68,In_145,In_365);
xor U69 (N_69,In_474,In_425);
or U70 (N_70,In_399,In_102);
nor U71 (N_71,In_362,In_71);
xor U72 (N_72,In_431,In_415);
or U73 (N_73,In_402,In_44);
or U74 (N_74,In_108,In_167);
xor U75 (N_75,In_24,In_467);
and U76 (N_76,In_420,In_249);
xnor U77 (N_77,In_363,In_314);
xor U78 (N_78,In_159,In_38);
nor U79 (N_79,In_460,In_125);
nor U80 (N_80,In_55,In_95);
nor U81 (N_81,In_483,In_88);
or U82 (N_82,In_13,In_255);
nor U83 (N_83,In_296,In_77);
nor U84 (N_84,In_75,In_168);
or U85 (N_85,In_465,In_138);
and U86 (N_86,In_157,In_339);
xor U87 (N_87,In_127,In_391);
and U88 (N_88,In_383,In_409);
xor U89 (N_89,In_9,In_288);
nand U90 (N_90,In_189,In_107);
nand U91 (N_91,In_276,In_126);
nor U92 (N_92,In_337,In_280);
xor U93 (N_93,In_408,In_109);
nand U94 (N_94,In_466,In_461);
nor U95 (N_95,In_39,In_488);
xor U96 (N_96,In_197,In_36);
nand U97 (N_97,In_241,In_81);
xor U98 (N_98,In_104,In_272);
or U99 (N_99,In_346,In_111);
xor U100 (N_100,N_12,In_225);
nor U101 (N_101,In_327,N_32);
nor U102 (N_102,In_229,In_234);
or U103 (N_103,N_31,In_186);
or U104 (N_104,In_103,In_390);
and U105 (N_105,In_92,N_3);
nor U106 (N_106,In_22,N_67);
nor U107 (N_107,In_137,N_66);
and U108 (N_108,In_316,N_63);
or U109 (N_109,In_342,In_203);
nor U110 (N_110,In_261,In_215);
nand U111 (N_111,In_210,N_59);
nor U112 (N_112,In_76,In_495);
or U113 (N_113,In_304,In_410);
and U114 (N_114,N_86,N_38);
nand U115 (N_115,In_313,In_307);
nand U116 (N_116,In_334,In_213);
nor U117 (N_117,In_19,In_180);
or U118 (N_118,In_243,In_114);
or U119 (N_119,In_407,In_397);
xor U120 (N_120,In_294,In_217);
xor U121 (N_121,In_347,In_150);
nor U122 (N_122,In_113,In_12);
nand U123 (N_123,In_475,In_30);
xor U124 (N_124,In_62,In_379);
or U125 (N_125,In_251,In_301);
and U126 (N_126,In_248,In_489);
and U127 (N_127,In_129,In_303);
nand U128 (N_128,N_84,In_354);
and U129 (N_129,In_133,In_52);
or U130 (N_130,N_48,In_7);
or U131 (N_131,N_27,In_17);
and U132 (N_132,In_312,In_286);
nand U133 (N_133,N_90,N_14);
nor U134 (N_134,In_427,In_357);
xnor U135 (N_135,In_70,N_72);
xor U136 (N_136,N_19,In_41);
nand U137 (N_137,In_219,In_183);
or U138 (N_138,In_403,In_493);
nand U139 (N_139,N_68,In_66);
nand U140 (N_140,In_51,In_165);
nor U141 (N_141,In_260,In_254);
and U142 (N_142,N_99,In_96);
and U143 (N_143,N_40,N_0);
xnor U144 (N_144,In_42,In_473);
nand U145 (N_145,N_81,In_283);
or U146 (N_146,N_65,N_39);
xnor U147 (N_147,In_169,In_21);
nand U148 (N_148,In_78,In_149);
xor U149 (N_149,N_95,In_90);
nor U150 (N_150,In_320,N_30);
or U151 (N_151,In_115,In_437);
nand U152 (N_152,In_221,In_459);
or U153 (N_153,In_194,In_302);
xor U154 (N_154,N_53,In_392);
xor U155 (N_155,In_282,In_155);
nor U156 (N_156,In_34,N_26);
and U157 (N_157,In_336,In_240);
nand U158 (N_158,In_310,In_247);
xor U159 (N_159,N_49,In_35);
or U160 (N_160,In_435,N_78);
nor U161 (N_161,N_1,N_22);
or U162 (N_162,N_87,N_43);
nor U163 (N_163,N_15,N_23);
nor U164 (N_164,In_80,In_356);
xnor U165 (N_165,N_45,In_233);
nand U166 (N_166,N_35,In_479);
xnor U167 (N_167,N_57,In_323);
or U168 (N_168,In_232,In_289);
xor U169 (N_169,In_156,In_73);
nor U170 (N_170,In_139,N_83);
nor U171 (N_171,In_220,In_193);
and U172 (N_172,N_52,In_148);
and U173 (N_173,In_196,In_27);
and U174 (N_174,In_367,In_246);
xnor U175 (N_175,In_469,In_146);
or U176 (N_176,In_211,N_56);
xnor U177 (N_177,In_317,In_338);
xnor U178 (N_178,In_207,In_47);
or U179 (N_179,In_496,In_463);
and U180 (N_180,N_18,N_75);
or U181 (N_181,In_382,In_119);
nand U182 (N_182,In_321,In_484);
nor U183 (N_183,In_421,In_20);
xnor U184 (N_184,N_42,N_62);
nand U185 (N_185,In_1,In_351);
and U186 (N_186,In_3,In_223);
nand U187 (N_187,N_80,In_319);
xnor U188 (N_188,In_443,N_54);
or U189 (N_189,In_450,In_191);
xor U190 (N_190,N_17,N_7);
or U191 (N_191,In_476,In_65);
and U192 (N_192,In_94,In_85);
xor U193 (N_193,N_96,In_123);
and U194 (N_194,In_269,N_44);
nor U195 (N_195,In_237,In_349);
or U196 (N_196,In_398,In_257);
or U197 (N_197,In_236,In_494);
xnor U198 (N_198,In_372,N_73);
or U199 (N_199,N_41,In_152);
nand U200 (N_200,In_177,In_116);
xnor U201 (N_201,In_326,In_378);
nor U202 (N_202,In_231,N_199);
nor U203 (N_203,In_480,N_137);
and U204 (N_204,In_256,N_110);
xnor U205 (N_205,N_196,In_324);
and U206 (N_206,In_291,In_424);
nand U207 (N_207,N_120,N_155);
or U208 (N_208,N_194,N_11);
or U209 (N_209,In_82,In_262);
nor U210 (N_210,In_380,In_333);
and U211 (N_211,In_110,N_172);
or U212 (N_212,In_117,In_172);
nand U213 (N_213,In_422,In_192);
nand U214 (N_214,N_127,In_287);
nand U215 (N_215,N_161,In_298);
nor U216 (N_216,In_99,In_91);
xor U217 (N_217,In_470,In_87);
nor U218 (N_218,In_106,In_471);
and U219 (N_219,N_193,N_143);
nand U220 (N_220,In_199,In_418);
xnor U221 (N_221,In_281,N_175);
and U222 (N_222,N_107,In_164);
xor U223 (N_223,N_132,N_46);
nor U224 (N_224,In_105,N_82);
nand U225 (N_225,N_6,In_490);
nand U226 (N_226,In_212,In_100);
and U227 (N_227,In_384,N_149);
and U228 (N_228,N_163,In_361);
nand U229 (N_229,N_130,N_183);
and U230 (N_230,N_192,In_50);
and U231 (N_231,N_136,In_253);
nand U232 (N_232,In_411,N_152);
or U233 (N_233,N_154,In_184);
nand U234 (N_234,N_37,In_83);
xnor U235 (N_235,In_482,In_405);
xor U236 (N_236,In_206,In_93);
and U237 (N_237,In_130,In_228);
xnor U238 (N_238,N_47,In_185);
xor U239 (N_239,N_123,In_64);
xnor U240 (N_240,N_24,N_195);
or U241 (N_241,In_160,In_37);
xor U242 (N_242,In_53,In_98);
or U243 (N_243,In_278,In_25);
or U244 (N_244,N_61,In_369);
nand U245 (N_245,In_235,In_444);
nor U246 (N_246,In_352,N_34);
xor U247 (N_247,N_121,N_147);
or U248 (N_248,N_10,N_188);
or U249 (N_249,In_401,In_322);
nand U250 (N_250,N_180,N_118);
and U251 (N_251,In_4,N_8);
xnor U252 (N_252,In_28,N_125);
and U253 (N_253,N_106,In_359);
and U254 (N_254,N_100,N_135);
nor U255 (N_255,In_429,In_101);
nor U256 (N_256,N_60,N_20);
and U257 (N_257,N_2,N_69);
and U258 (N_258,N_146,In_419);
xnor U259 (N_259,N_28,In_216);
and U260 (N_260,N_5,N_93);
xnor U261 (N_261,N_166,N_159);
or U262 (N_262,In_393,In_438);
and U263 (N_263,N_51,In_453);
and U264 (N_264,N_101,N_109);
xor U265 (N_265,N_158,In_222);
and U266 (N_266,N_177,N_189);
nor U267 (N_267,In_136,N_187);
nor U268 (N_268,N_119,N_184);
nand U269 (N_269,In_464,N_153);
nor U270 (N_270,N_197,In_385);
nand U271 (N_271,In_330,In_173);
xnor U272 (N_272,N_79,N_145);
nor U273 (N_273,In_270,N_165);
or U274 (N_274,N_115,In_388);
and U275 (N_275,In_142,N_150);
nor U276 (N_276,In_227,N_156);
nand U277 (N_277,In_259,N_58);
xnor U278 (N_278,In_6,N_9);
or U279 (N_279,In_49,N_126);
xnor U280 (N_280,In_209,N_92);
xor U281 (N_281,In_273,N_124);
xnor U282 (N_282,N_142,N_151);
xor U283 (N_283,N_89,In_43);
nor U284 (N_284,In_266,N_174);
nand U285 (N_285,N_168,N_182);
xor U286 (N_286,In_486,In_238);
or U287 (N_287,N_162,N_102);
nor U288 (N_288,N_16,In_208);
nand U289 (N_289,N_167,N_176);
and U290 (N_290,N_134,N_122);
or U291 (N_291,In_244,In_368);
or U292 (N_292,In_311,N_181);
or U293 (N_293,N_198,In_284);
or U294 (N_294,In_413,N_33);
and U295 (N_295,N_116,In_275);
and U296 (N_296,N_94,N_160);
xnor U297 (N_297,In_134,N_148);
or U298 (N_298,In_202,In_458);
nand U299 (N_299,N_70,In_315);
nor U300 (N_300,N_104,N_242);
or U301 (N_301,In_218,N_208);
nor U302 (N_302,N_85,In_171);
nor U303 (N_303,N_50,N_276);
nand U304 (N_304,N_232,N_289);
and U305 (N_305,In_263,N_64);
nand U306 (N_306,In_29,N_253);
nand U307 (N_307,N_128,In_63);
or U308 (N_308,N_206,In_331);
and U309 (N_309,N_219,N_248);
nand U310 (N_310,In_279,N_291);
or U311 (N_311,N_265,In_426);
nor U312 (N_312,N_230,N_138);
nor U313 (N_313,N_74,N_173);
nand U314 (N_314,In_335,N_280);
and U315 (N_315,N_112,N_264);
xnor U316 (N_316,N_277,N_209);
or U317 (N_317,N_266,N_236);
nor U318 (N_318,N_296,N_249);
nand U319 (N_319,N_98,N_113);
and U320 (N_320,N_237,In_395);
nand U321 (N_321,N_213,N_212);
nor U322 (N_322,N_231,N_13);
nor U323 (N_323,N_76,N_108);
xor U324 (N_324,N_284,N_240);
and U325 (N_325,N_269,In_309);
nor U326 (N_326,N_281,N_191);
or U327 (N_327,In_325,N_260);
nor U328 (N_328,N_228,N_111);
nor U329 (N_329,N_211,N_25);
nor U330 (N_330,N_288,In_135);
and U331 (N_331,N_259,N_88);
and U332 (N_332,N_77,N_275);
or U333 (N_333,N_278,N_256);
xor U334 (N_334,N_103,N_273);
or U335 (N_335,In_158,In_163);
nand U336 (N_336,N_297,N_139);
xnor U337 (N_337,In_54,N_245);
nand U338 (N_338,N_144,N_241);
or U339 (N_339,N_250,In_366);
and U340 (N_340,In_364,N_171);
nor U341 (N_341,N_157,N_268);
xnor U342 (N_342,N_169,N_258);
nor U343 (N_343,N_190,N_207);
or U344 (N_344,N_247,N_21);
and U345 (N_345,In_478,N_200);
or U346 (N_346,In_141,In_442);
and U347 (N_347,N_252,In_79);
xor U348 (N_348,N_225,N_140);
nor U349 (N_349,N_97,N_295);
xnor U350 (N_350,N_217,In_277);
and U351 (N_351,N_224,N_234);
and U352 (N_352,N_292,N_233);
or U353 (N_353,N_55,N_229);
xor U354 (N_354,In_205,N_186);
xor U355 (N_355,N_215,N_262);
or U356 (N_356,N_294,N_287);
nand U357 (N_357,In_198,N_29);
nor U358 (N_358,In_121,N_131);
nor U359 (N_359,In_499,N_293);
and U360 (N_360,N_4,In_151);
or U361 (N_361,N_263,N_170);
or U362 (N_362,In_86,N_221);
xor U363 (N_363,N_141,N_178);
and U364 (N_364,In_67,N_210);
xor U365 (N_365,N_283,In_23);
xor U366 (N_366,In_440,N_243);
xnor U367 (N_367,N_201,In_182);
nor U368 (N_368,In_59,N_254);
and U369 (N_369,In_452,In_0);
xor U370 (N_370,In_370,N_226);
and U371 (N_371,N_279,N_261);
xnor U372 (N_372,In_290,N_71);
and U373 (N_373,N_267,N_204);
and U374 (N_374,N_272,In_2);
nor U375 (N_375,N_244,In_33);
and U376 (N_376,N_218,N_164);
nand U377 (N_377,N_105,N_282);
nor U378 (N_378,In_162,N_251);
xnor U379 (N_379,N_220,N_290);
nand U380 (N_380,In_224,In_258);
and U381 (N_381,In_271,N_117);
nand U382 (N_382,In_394,N_114);
nor U383 (N_383,N_246,N_179);
and U384 (N_384,N_238,N_133);
xor U385 (N_385,N_202,In_178);
or U386 (N_386,N_235,N_299);
and U387 (N_387,N_239,N_227);
or U388 (N_388,N_286,N_222);
nor U389 (N_389,N_205,N_257);
nor U390 (N_390,In_406,In_350);
nand U391 (N_391,N_223,N_298);
nand U392 (N_392,In_472,N_271);
nand U393 (N_393,N_255,N_36);
xnor U394 (N_394,N_203,N_91);
and U395 (N_395,N_216,N_214);
or U396 (N_396,N_129,N_270);
or U397 (N_397,N_274,In_414);
and U398 (N_398,In_122,In_373);
or U399 (N_399,N_185,N_285);
xor U400 (N_400,N_304,N_365);
nand U401 (N_401,N_333,N_393);
nand U402 (N_402,N_319,N_395);
nor U403 (N_403,N_323,N_343);
nor U404 (N_404,N_300,N_351);
or U405 (N_405,N_337,N_358);
xor U406 (N_406,N_364,N_347);
xor U407 (N_407,N_302,N_330);
and U408 (N_408,N_316,N_394);
nand U409 (N_409,N_356,N_357);
or U410 (N_410,N_391,N_369);
nor U411 (N_411,N_378,N_321);
nor U412 (N_412,N_390,N_371);
xnor U413 (N_413,N_346,N_386);
or U414 (N_414,N_373,N_320);
xnor U415 (N_415,N_329,N_375);
nand U416 (N_416,N_399,N_324);
nand U417 (N_417,N_389,N_314);
nor U418 (N_418,N_340,N_311);
and U419 (N_419,N_397,N_313);
nor U420 (N_420,N_303,N_388);
nor U421 (N_421,N_353,N_376);
nand U422 (N_422,N_381,N_398);
or U423 (N_423,N_305,N_350);
xor U424 (N_424,N_328,N_331);
or U425 (N_425,N_368,N_352);
and U426 (N_426,N_344,N_361);
or U427 (N_427,N_307,N_355);
nand U428 (N_428,N_325,N_309);
xnor U429 (N_429,N_308,N_363);
nor U430 (N_430,N_312,N_354);
or U431 (N_431,N_366,N_380);
and U432 (N_432,N_334,N_396);
nand U433 (N_433,N_318,N_349);
and U434 (N_434,N_392,N_384);
and U435 (N_435,N_315,N_326);
or U436 (N_436,N_336,N_322);
and U437 (N_437,N_377,N_306);
nand U438 (N_438,N_367,N_370);
nand U439 (N_439,N_342,N_310);
nand U440 (N_440,N_382,N_339);
nand U441 (N_441,N_317,N_383);
or U442 (N_442,N_335,N_338);
nor U443 (N_443,N_379,N_360);
nand U444 (N_444,N_387,N_348);
or U445 (N_445,N_301,N_359);
nor U446 (N_446,N_332,N_372);
or U447 (N_447,N_341,N_374);
and U448 (N_448,N_345,N_385);
and U449 (N_449,N_362,N_327);
nand U450 (N_450,N_376,N_326);
and U451 (N_451,N_310,N_304);
and U452 (N_452,N_394,N_322);
nand U453 (N_453,N_325,N_381);
xnor U454 (N_454,N_372,N_348);
nand U455 (N_455,N_306,N_360);
or U456 (N_456,N_325,N_345);
or U457 (N_457,N_324,N_325);
nand U458 (N_458,N_346,N_313);
nor U459 (N_459,N_360,N_375);
or U460 (N_460,N_373,N_359);
or U461 (N_461,N_371,N_382);
and U462 (N_462,N_398,N_370);
nand U463 (N_463,N_311,N_351);
nand U464 (N_464,N_320,N_390);
or U465 (N_465,N_335,N_325);
xor U466 (N_466,N_373,N_300);
and U467 (N_467,N_322,N_305);
nand U468 (N_468,N_322,N_350);
xnor U469 (N_469,N_303,N_340);
nor U470 (N_470,N_332,N_393);
and U471 (N_471,N_320,N_356);
nand U472 (N_472,N_324,N_309);
nor U473 (N_473,N_346,N_374);
nor U474 (N_474,N_338,N_331);
and U475 (N_475,N_316,N_365);
or U476 (N_476,N_347,N_352);
and U477 (N_477,N_317,N_385);
xor U478 (N_478,N_389,N_357);
or U479 (N_479,N_338,N_327);
nand U480 (N_480,N_308,N_340);
nor U481 (N_481,N_316,N_361);
or U482 (N_482,N_354,N_328);
or U483 (N_483,N_376,N_377);
nor U484 (N_484,N_377,N_354);
nor U485 (N_485,N_390,N_395);
or U486 (N_486,N_316,N_339);
nand U487 (N_487,N_353,N_394);
nor U488 (N_488,N_356,N_312);
or U489 (N_489,N_365,N_398);
xor U490 (N_490,N_329,N_314);
or U491 (N_491,N_360,N_324);
or U492 (N_492,N_305,N_393);
nor U493 (N_493,N_348,N_331);
or U494 (N_494,N_339,N_389);
nand U495 (N_495,N_320,N_351);
nand U496 (N_496,N_354,N_397);
xnor U497 (N_497,N_350,N_326);
xor U498 (N_498,N_336,N_348);
or U499 (N_499,N_318,N_315);
nand U500 (N_500,N_437,N_489);
nor U501 (N_501,N_463,N_406);
nand U502 (N_502,N_472,N_446);
xnor U503 (N_503,N_438,N_450);
nor U504 (N_504,N_403,N_415);
or U505 (N_505,N_467,N_453);
xor U506 (N_506,N_488,N_456);
and U507 (N_507,N_490,N_425);
or U508 (N_508,N_498,N_401);
nor U509 (N_509,N_476,N_429);
or U510 (N_510,N_451,N_436);
and U511 (N_511,N_474,N_465);
and U512 (N_512,N_428,N_458);
or U513 (N_513,N_494,N_422);
or U514 (N_514,N_411,N_452);
xnor U515 (N_515,N_445,N_486);
xnor U516 (N_516,N_447,N_431);
or U517 (N_517,N_466,N_421);
nand U518 (N_518,N_443,N_473);
and U519 (N_519,N_417,N_419);
xnor U520 (N_520,N_479,N_480);
or U521 (N_521,N_441,N_497);
nand U522 (N_522,N_424,N_496);
nand U523 (N_523,N_481,N_439);
and U524 (N_524,N_495,N_432);
xor U525 (N_525,N_423,N_409);
xnor U526 (N_526,N_483,N_444);
and U527 (N_527,N_477,N_455);
nor U528 (N_528,N_427,N_449);
nor U529 (N_529,N_430,N_454);
and U530 (N_530,N_493,N_426);
or U531 (N_531,N_460,N_404);
xor U532 (N_532,N_492,N_491);
or U533 (N_533,N_462,N_499);
nor U534 (N_534,N_457,N_416);
nand U535 (N_535,N_412,N_482);
nand U536 (N_536,N_468,N_485);
or U537 (N_537,N_408,N_418);
or U538 (N_538,N_448,N_471);
nor U539 (N_539,N_400,N_470);
nor U540 (N_540,N_413,N_475);
xor U541 (N_541,N_405,N_435);
nor U542 (N_542,N_461,N_414);
or U543 (N_543,N_402,N_410);
nand U544 (N_544,N_433,N_487);
xor U545 (N_545,N_420,N_407);
nor U546 (N_546,N_484,N_434);
xor U547 (N_547,N_478,N_469);
nor U548 (N_548,N_459,N_442);
nor U549 (N_549,N_464,N_440);
xor U550 (N_550,N_486,N_463);
or U551 (N_551,N_409,N_438);
and U552 (N_552,N_436,N_424);
or U553 (N_553,N_468,N_489);
nor U554 (N_554,N_486,N_465);
nand U555 (N_555,N_457,N_442);
nor U556 (N_556,N_408,N_412);
nor U557 (N_557,N_406,N_458);
nand U558 (N_558,N_447,N_482);
nand U559 (N_559,N_489,N_424);
xor U560 (N_560,N_439,N_463);
and U561 (N_561,N_419,N_489);
nand U562 (N_562,N_488,N_485);
nor U563 (N_563,N_497,N_430);
nand U564 (N_564,N_494,N_443);
xor U565 (N_565,N_400,N_467);
nand U566 (N_566,N_403,N_417);
xor U567 (N_567,N_422,N_492);
or U568 (N_568,N_474,N_420);
nor U569 (N_569,N_416,N_442);
nand U570 (N_570,N_489,N_467);
nor U571 (N_571,N_444,N_493);
nor U572 (N_572,N_498,N_439);
and U573 (N_573,N_484,N_481);
and U574 (N_574,N_437,N_430);
xnor U575 (N_575,N_456,N_401);
nand U576 (N_576,N_409,N_476);
and U577 (N_577,N_487,N_442);
or U578 (N_578,N_400,N_411);
and U579 (N_579,N_457,N_471);
or U580 (N_580,N_434,N_445);
xor U581 (N_581,N_499,N_470);
xnor U582 (N_582,N_451,N_490);
xor U583 (N_583,N_424,N_433);
nand U584 (N_584,N_491,N_493);
xnor U585 (N_585,N_476,N_485);
and U586 (N_586,N_468,N_497);
and U587 (N_587,N_491,N_418);
nand U588 (N_588,N_483,N_449);
or U589 (N_589,N_440,N_476);
nor U590 (N_590,N_496,N_437);
nor U591 (N_591,N_434,N_408);
and U592 (N_592,N_472,N_497);
and U593 (N_593,N_486,N_470);
and U594 (N_594,N_415,N_424);
nor U595 (N_595,N_483,N_432);
nand U596 (N_596,N_423,N_403);
nand U597 (N_597,N_438,N_435);
nand U598 (N_598,N_429,N_478);
nand U599 (N_599,N_470,N_463);
nor U600 (N_600,N_512,N_516);
and U601 (N_601,N_566,N_579);
and U602 (N_602,N_548,N_537);
xor U603 (N_603,N_506,N_505);
xnor U604 (N_604,N_561,N_597);
xor U605 (N_605,N_532,N_523);
and U606 (N_606,N_502,N_568);
or U607 (N_607,N_590,N_589);
or U608 (N_608,N_517,N_583);
xor U609 (N_609,N_539,N_529);
nand U610 (N_610,N_591,N_504);
and U611 (N_611,N_543,N_598);
xnor U612 (N_612,N_592,N_587);
nor U613 (N_613,N_530,N_554);
and U614 (N_614,N_586,N_515);
nand U615 (N_615,N_574,N_511);
and U616 (N_616,N_525,N_546);
and U617 (N_617,N_533,N_526);
xnor U618 (N_618,N_569,N_528);
nand U619 (N_619,N_536,N_552);
and U620 (N_620,N_507,N_599);
xor U621 (N_621,N_538,N_563);
nand U622 (N_622,N_581,N_585);
and U623 (N_623,N_520,N_509);
and U624 (N_624,N_524,N_514);
xor U625 (N_625,N_565,N_510);
nand U626 (N_626,N_547,N_555);
nand U627 (N_627,N_521,N_570);
and U628 (N_628,N_558,N_557);
xor U629 (N_629,N_593,N_513);
or U630 (N_630,N_508,N_544);
and U631 (N_631,N_595,N_580);
and U632 (N_632,N_562,N_594);
nor U633 (N_633,N_503,N_553);
and U634 (N_634,N_575,N_577);
xnor U635 (N_635,N_559,N_576);
nor U636 (N_636,N_542,N_501);
and U637 (N_637,N_550,N_522);
or U638 (N_638,N_564,N_540);
nor U639 (N_639,N_551,N_588);
nand U640 (N_640,N_545,N_519);
xnor U641 (N_641,N_531,N_571);
xnor U642 (N_642,N_560,N_500);
and U643 (N_643,N_527,N_556);
and U644 (N_644,N_572,N_584);
xnor U645 (N_645,N_535,N_573);
or U646 (N_646,N_534,N_596);
nand U647 (N_647,N_578,N_549);
or U648 (N_648,N_567,N_518);
nor U649 (N_649,N_541,N_582);
and U650 (N_650,N_557,N_596);
nor U651 (N_651,N_505,N_595);
nand U652 (N_652,N_537,N_547);
nand U653 (N_653,N_596,N_563);
nor U654 (N_654,N_560,N_509);
and U655 (N_655,N_581,N_524);
nor U656 (N_656,N_572,N_563);
and U657 (N_657,N_566,N_564);
and U658 (N_658,N_505,N_567);
xor U659 (N_659,N_522,N_587);
nand U660 (N_660,N_591,N_522);
or U661 (N_661,N_555,N_588);
or U662 (N_662,N_559,N_528);
or U663 (N_663,N_542,N_581);
and U664 (N_664,N_521,N_581);
and U665 (N_665,N_533,N_541);
xnor U666 (N_666,N_574,N_577);
nor U667 (N_667,N_510,N_597);
nor U668 (N_668,N_528,N_536);
nand U669 (N_669,N_577,N_595);
nand U670 (N_670,N_572,N_595);
xnor U671 (N_671,N_564,N_577);
nor U672 (N_672,N_583,N_539);
nand U673 (N_673,N_531,N_522);
or U674 (N_674,N_558,N_508);
or U675 (N_675,N_580,N_523);
nand U676 (N_676,N_594,N_517);
nor U677 (N_677,N_590,N_562);
and U678 (N_678,N_590,N_575);
nand U679 (N_679,N_570,N_539);
and U680 (N_680,N_594,N_552);
nand U681 (N_681,N_585,N_547);
xor U682 (N_682,N_585,N_590);
xnor U683 (N_683,N_539,N_589);
nor U684 (N_684,N_553,N_589);
and U685 (N_685,N_541,N_544);
nand U686 (N_686,N_509,N_599);
or U687 (N_687,N_549,N_548);
nor U688 (N_688,N_514,N_517);
xor U689 (N_689,N_522,N_589);
nand U690 (N_690,N_502,N_548);
nand U691 (N_691,N_567,N_506);
nor U692 (N_692,N_584,N_583);
or U693 (N_693,N_559,N_594);
nor U694 (N_694,N_506,N_528);
or U695 (N_695,N_586,N_556);
nor U696 (N_696,N_512,N_525);
nand U697 (N_697,N_557,N_540);
xor U698 (N_698,N_528,N_541);
nand U699 (N_699,N_577,N_529);
or U700 (N_700,N_683,N_600);
and U701 (N_701,N_654,N_686);
and U702 (N_702,N_629,N_610);
nand U703 (N_703,N_653,N_661);
xnor U704 (N_704,N_655,N_604);
and U705 (N_705,N_619,N_614);
nand U706 (N_706,N_638,N_694);
nand U707 (N_707,N_639,N_668);
xor U708 (N_708,N_692,N_627);
and U709 (N_709,N_671,N_681);
nand U710 (N_710,N_612,N_688);
nand U711 (N_711,N_689,N_673);
or U712 (N_712,N_690,N_626);
and U713 (N_713,N_669,N_618);
xor U714 (N_714,N_650,N_608);
nand U715 (N_715,N_609,N_616);
and U716 (N_716,N_660,N_684);
xnor U717 (N_717,N_602,N_634);
nand U718 (N_718,N_680,N_676);
nor U719 (N_719,N_620,N_658);
nand U720 (N_720,N_621,N_630);
xnor U721 (N_721,N_665,N_628);
nand U722 (N_722,N_622,N_656);
or U723 (N_723,N_606,N_696);
nor U724 (N_724,N_631,N_693);
nor U725 (N_725,N_674,N_699);
and U726 (N_726,N_636,N_677);
xor U727 (N_727,N_648,N_643);
nor U728 (N_728,N_659,N_695);
nor U729 (N_729,N_611,N_691);
or U730 (N_730,N_613,N_697);
and U731 (N_731,N_651,N_678);
and U732 (N_732,N_672,N_666);
nand U733 (N_733,N_641,N_652);
nor U734 (N_734,N_623,N_698);
xor U735 (N_735,N_605,N_645);
and U736 (N_736,N_603,N_682);
xnor U737 (N_737,N_635,N_687);
or U738 (N_738,N_640,N_642);
nor U739 (N_739,N_633,N_607);
nand U740 (N_740,N_625,N_667);
nor U741 (N_741,N_675,N_663);
or U742 (N_742,N_632,N_647);
nor U743 (N_743,N_646,N_670);
or U744 (N_744,N_679,N_649);
nor U745 (N_745,N_657,N_685);
nand U746 (N_746,N_644,N_617);
nor U747 (N_747,N_624,N_615);
and U748 (N_748,N_637,N_601);
xnor U749 (N_749,N_662,N_664);
or U750 (N_750,N_624,N_620);
nand U751 (N_751,N_655,N_605);
or U752 (N_752,N_641,N_610);
or U753 (N_753,N_669,N_630);
or U754 (N_754,N_660,N_672);
nor U755 (N_755,N_673,N_677);
or U756 (N_756,N_624,N_668);
or U757 (N_757,N_675,N_629);
xnor U758 (N_758,N_661,N_670);
or U759 (N_759,N_612,N_696);
nor U760 (N_760,N_621,N_646);
nand U761 (N_761,N_691,N_617);
nand U762 (N_762,N_663,N_646);
xnor U763 (N_763,N_613,N_684);
or U764 (N_764,N_639,N_622);
and U765 (N_765,N_634,N_606);
nor U766 (N_766,N_609,N_615);
xor U767 (N_767,N_687,N_653);
and U768 (N_768,N_686,N_620);
or U769 (N_769,N_645,N_626);
and U770 (N_770,N_692,N_635);
nand U771 (N_771,N_608,N_618);
nand U772 (N_772,N_698,N_614);
xnor U773 (N_773,N_627,N_686);
nand U774 (N_774,N_634,N_601);
xor U775 (N_775,N_672,N_609);
or U776 (N_776,N_676,N_692);
or U777 (N_777,N_667,N_689);
nor U778 (N_778,N_613,N_657);
or U779 (N_779,N_644,N_607);
xnor U780 (N_780,N_674,N_678);
or U781 (N_781,N_654,N_667);
and U782 (N_782,N_635,N_620);
nand U783 (N_783,N_666,N_653);
nor U784 (N_784,N_657,N_605);
or U785 (N_785,N_661,N_655);
and U786 (N_786,N_678,N_628);
nand U787 (N_787,N_634,N_687);
nor U788 (N_788,N_613,N_625);
nand U789 (N_789,N_618,N_642);
or U790 (N_790,N_671,N_664);
nor U791 (N_791,N_665,N_622);
nand U792 (N_792,N_611,N_645);
and U793 (N_793,N_631,N_678);
xor U794 (N_794,N_635,N_680);
xor U795 (N_795,N_614,N_646);
xor U796 (N_796,N_636,N_685);
xnor U797 (N_797,N_634,N_679);
or U798 (N_798,N_676,N_675);
or U799 (N_799,N_658,N_673);
nor U800 (N_800,N_703,N_757);
and U801 (N_801,N_730,N_748);
or U802 (N_802,N_790,N_783);
xnor U803 (N_803,N_701,N_763);
nor U804 (N_804,N_791,N_782);
nand U805 (N_805,N_769,N_735);
nor U806 (N_806,N_767,N_729);
and U807 (N_807,N_712,N_736);
or U808 (N_808,N_794,N_724);
or U809 (N_809,N_702,N_737);
nor U810 (N_810,N_741,N_707);
or U811 (N_811,N_708,N_739);
and U812 (N_812,N_725,N_705);
nor U813 (N_813,N_744,N_778);
or U814 (N_814,N_731,N_732);
and U815 (N_815,N_781,N_768);
xor U816 (N_816,N_770,N_713);
and U817 (N_817,N_711,N_747);
nor U818 (N_818,N_776,N_792);
xnor U819 (N_819,N_709,N_799);
or U820 (N_820,N_720,N_734);
and U821 (N_821,N_765,N_789);
or U822 (N_822,N_745,N_715);
and U823 (N_823,N_785,N_714);
nand U824 (N_824,N_700,N_780);
xor U825 (N_825,N_723,N_766);
nor U826 (N_826,N_797,N_716);
or U827 (N_827,N_743,N_722);
xor U828 (N_828,N_775,N_795);
nand U829 (N_829,N_762,N_752);
xor U830 (N_830,N_710,N_796);
and U831 (N_831,N_771,N_760);
or U832 (N_832,N_746,N_788);
xor U833 (N_833,N_784,N_777);
and U834 (N_834,N_761,N_779);
nand U835 (N_835,N_786,N_793);
or U836 (N_836,N_759,N_754);
nand U837 (N_837,N_706,N_733);
or U838 (N_838,N_738,N_717);
nand U839 (N_839,N_719,N_721);
xnor U840 (N_840,N_753,N_755);
nor U841 (N_841,N_758,N_704);
nor U842 (N_842,N_750,N_726);
nand U843 (N_843,N_756,N_749);
nand U844 (N_844,N_773,N_718);
or U845 (N_845,N_787,N_764);
nor U846 (N_846,N_740,N_798);
nand U847 (N_847,N_772,N_727);
and U848 (N_848,N_742,N_728);
xor U849 (N_849,N_774,N_751);
and U850 (N_850,N_746,N_716);
or U851 (N_851,N_744,N_748);
and U852 (N_852,N_740,N_749);
and U853 (N_853,N_753,N_735);
and U854 (N_854,N_724,N_760);
nor U855 (N_855,N_756,N_771);
xnor U856 (N_856,N_749,N_702);
nor U857 (N_857,N_775,N_717);
nor U858 (N_858,N_768,N_794);
or U859 (N_859,N_708,N_766);
nand U860 (N_860,N_797,N_764);
nand U861 (N_861,N_713,N_765);
and U862 (N_862,N_790,N_782);
and U863 (N_863,N_758,N_720);
xnor U864 (N_864,N_792,N_777);
and U865 (N_865,N_748,N_785);
nor U866 (N_866,N_752,N_749);
nor U867 (N_867,N_729,N_795);
xor U868 (N_868,N_740,N_799);
and U869 (N_869,N_702,N_762);
or U870 (N_870,N_746,N_741);
or U871 (N_871,N_772,N_710);
and U872 (N_872,N_796,N_735);
nand U873 (N_873,N_711,N_781);
xnor U874 (N_874,N_768,N_755);
nor U875 (N_875,N_758,N_733);
nand U876 (N_876,N_784,N_748);
or U877 (N_877,N_700,N_715);
and U878 (N_878,N_774,N_728);
nor U879 (N_879,N_721,N_733);
or U880 (N_880,N_756,N_760);
and U881 (N_881,N_749,N_763);
xnor U882 (N_882,N_758,N_746);
xnor U883 (N_883,N_775,N_779);
nor U884 (N_884,N_701,N_704);
nor U885 (N_885,N_744,N_739);
nor U886 (N_886,N_733,N_765);
and U887 (N_887,N_746,N_790);
xor U888 (N_888,N_764,N_765);
nand U889 (N_889,N_744,N_727);
and U890 (N_890,N_705,N_787);
nand U891 (N_891,N_756,N_736);
and U892 (N_892,N_757,N_745);
nand U893 (N_893,N_778,N_748);
or U894 (N_894,N_736,N_792);
and U895 (N_895,N_765,N_703);
or U896 (N_896,N_795,N_779);
nor U897 (N_897,N_719,N_754);
and U898 (N_898,N_715,N_716);
xnor U899 (N_899,N_746,N_773);
nor U900 (N_900,N_877,N_827);
nor U901 (N_901,N_891,N_846);
or U902 (N_902,N_868,N_876);
or U903 (N_903,N_875,N_821);
xor U904 (N_904,N_885,N_801);
or U905 (N_905,N_858,N_825);
and U906 (N_906,N_881,N_830);
nand U907 (N_907,N_835,N_855);
nor U908 (N_908,N_800,N_836);
nor U909 (N_909,N_848,N_840);
or U910 (N_910,N_823,N_857);
and U911 (N_911,N_831,N_870);
and U912 (N_912,N_871,N_834);
nor U913 (N_913,N_899,N_847);
and U914 (N_914,N_859,N_837);
and U915 (N_915,N_809,N_833);
nand U916 (N_916,N_883,N_816);
and U917 (N_917,N_882,N_851);
and U918 (N_918,N_890,N_813);
or U919 (N_919,N_892,N_802);
and U920 (N_920,N_894,N_808);
or U921 (N_921,N_895,N_874);
nor U922 (N_922,N_832,N_862);
and U923 (N_923,N_805,N_807);
xnor U924 (N_924,N_886,N_866);
nor U925 (N_925,N_878,N_863);
or U926 (N_926,N_898,N_879);
or U927 (N_927,N_828,N_869);
and U928 (N_928,N_893,N_838);
nand U929 (N_929,N_897,N_819);
and U930 (N_930,N_856,N_812);
xnor U931 (N_931,N_803,N_806);
xnor U932 (N_932,N_844,N_845);
xnor U933 (N_933,N_889,N_872);
xnor U934 (N_934,N_811,N_867);
and U935 (N_935,N_864,N_873);
nand U936 (N_936,N_829,N_841);
and U937 (N_937,N_861,N_824);
nor U938 (N_938,N_865,N_814);
nand U939 (N_939,N_804,N_896);
nor U940 (N_940,N_850,N_822);
nand U941 (N_941,N_817,N_818);
nor U942 (N_942,N_810,N_880);
xnor U943 (N_943,N_843,N_852);
or U944 (N_944,N_884,N_849);
or U945 (N_945,N_854,N_853);
and U946 (N_946,N_888,N_839);
or U947 (N_947,N_815,N_842);
or U948 (N_948,N_860,N_887);
or U949 (N_949,N_826,N_820);
nand U950 (N_950,N_854,N_803);
or U951 (N_951,N_851,N_856);
nand U952 (N_952,N_893,N_820);
nor U953 (N_953,N_808,N_825);
or U954 (N_954,N_862,N_873);
xor U955 (N_955,N_827,N_818);
xnor U956 (N_956,N_837,N_807);
nand U957 (N_957,N_817,N_884);
nor U958 (N_958,N_878,N_897);
nand U959 (N_959,N_844,N_855);
nor U960 (N_960,N_826,N_835);
xnor U961 (N_961,N_865,N_860);
nand U962 (N_962,N_810,N_854);
xor U963 (N_963,N_835,N_847);
and U964 (N_964,N_813,N_887);
nand U965 (N_965,N_875,N_804);
nand U966 (N_966,N_857,N_829);
nand U967 (N_967,N_868,N_888);
or U968 (N_968,N_841,N_855);
nand U969 (N_969,N_822,N_817);
and U970 (N_970,N_842,N_819);
and U971 (N_971,N_873,N_898);
nand U972 (N_972,N_869,N_845);
nand U973 (N_973,N_855,N_889);
xnor U974 (N_974,N_864,N_856);
nor U975 (N_975,N_887,N_806);
nand U976 (N_976,N_843,N_896);
nor U977 (N_977,N_888,N_856);
and U978 (N_978,N_849,N_871);
nor U979 (N_979,N_854,N_820);
nor U980 (N_980,N_884,N_850);
nand U981 (N_981,N_896,N_877);
nand U982 (N_982,N_867,N_864);
or U983 (N_983,N_870,N_895);
xor U984 (N_984,N_840,N_879);
xor U985 (N_985,N_884,N_856);
xnor U986 (N_986,N_872,N_829);
and U987 (N_987,N_869,N_831);
nand U988 (N_988,N_858,N_816);
and U989 (N_989,N_820,N_836);
or U990 (N_990,N_818,N_816);
and U991 (N_991,N_844,N_879);
and U992 (N_992,N_867,N_854);
nor U993 (N_993,N_880,N_825);
xor U994 (N_994,N_817,N_810);
or U995 (N_995,N_813,N_802);
or U996 (N_996,N_807,N_833);
nand U997 (N_997,N_839,N_844);
xnor U998 (N_998,N_803,N_851);
xnor U999 (N_999,N_874,N_871);
nor U1000 (N_1000,N_922,N_979);
and U1001 (N_1001,N_970,N_949);
nand U1002 (N_1002,N_912,N_928);
and U1003 (N_1003,N_985,N_929);
xnor U1004 (N_1004,N_937,N_927);
xnor U1005 (N_1005,N_989,N_926);
or U1006 (N_1006,N_908,N_911);
nor U1007 (N_1007,N_914,N_921);
or U1008 (N_1008,N_969,N_971);
nor U1009 (N_1009,N_982,N_933);
nand U1010 (N_1010,N_932,N_938);
xor U1011 (N_1011,N_915,N_995);
nand U1012 (N_1012,N_963,N_991);
nor U1013 (N_1013,N_940,N_916);
xor U1014 (N_1014,N_973,N_944);
nand U1015 (N_1015,N_947,N_900);
xnor U1016 (N_1016,N_954,N_905);
or U1017 (N_1017,N_920,N_930);
xnor U1018 (N_1018,N_980,N_955);
xor U1019 (N_1019,N_903,N_994);
or U1020 (N_1020,N_961,N_990);
or U1021 (N_1021,N_935,N_904);
and U1022 (N_1022,N_945,N_986);
and U1023 (N_1023,N_997,N_941);
or U1024 (N_1024,N_950,N_942);
nor U1025 (N_1025,N_925,N_977);
or U1026 (N_1026,N_946,N_974);
and U1027 (N_1027,N_913,N_968);
and U1028 (N_1028,N_951,N_975);
xor U1029 (N_1029,N_919,N_999);
xnor U1030 (N_1030,N_902,N_983);
nand U1031 (N_1031,N_901,N_931);
nor U1032 (N_1032,N_910,N_978);
nor U1033 (N_1033,N_998,N_967);
xnor U1034 (N_1034,N_907,N_964);
nand U1035 (N_1035,N_923,N_909);
and U1036 (N_1036,N_958,N_917);
or U1037 (N_1037,N_918,N_984);
or U1038 (N_1038,N_948,N_965);
and U1039 (N_1039,N_966,N_939);
nor U1040 (N_1040,N_996,N_943);
nor U1041 (N_1041,N_934,N_972);
nand U1042 (N_1042,N_953,N_976);
xnor U1043 (N_1043,N_960,N_959);
nor U1044 (N_1044,N_962,N_981);
or U1045 (N_1045,N_924,N_992);
and U1046 (N_1046,N_952,N_956);
or U1047 (N_1047,N_993,N_936);
nand U1048 (N_1048,N_906,N_988);
xor U1049 (N_1049,N_957,N_987);
and U1050 (N_1050,N_909,N_931);
or U1051 (N_1051,N_931,N_922);
and U1052 (N_1052,N_939,N_968);
nand U1053 (N_1053,N_920,N_965);
nand U1054 (N_1054,N_932,N_909);
or U1055 (N_1055,N_917,N_902);
or U1056 (N_1056,N_953,N_924);
xor U1057 (N_1057,N_999,N_922);
or U1058 (N_1058,N_947,N_966);
and U1059 (N_1059,N_927,N_989);
or U1060 (N_1060,N_925,N_978);
or U1061 (N_1061,N_965,N_942);
and U1062 (N_1062,N_982,N_953);
nor U1063 (N_1063,N_941,N_936);
nor U1064 (N_1064,N_993,N_972);
nor U1065 (N_1065,N_908,N_946);
and U1066 (N_1066,N_972,N_952);
and U1067 (N_1067,N_932,N_943);
xor U1068 (N_1068,N_951,N_926);
nor U1069 (N_1069,N_928,N_936);
xor U1070 (N_1070,N_936,N_988);
nand U1071 (N_1071,N_935,N_913);
nand U1072 (N_1072,N_907,N_982);
nor U1073 (N_1073,N_926,N_933);
nand U1074 (N_1074,N_997,N_910);
nor U1075 (N_1075,N_902,N_947);
xnor U1076 (N_1076,N_952,N_912);
nand U1077 (N_1077,N_974,N_934);
nand U1078 (N_1078,N_942,N_908);
and U1079 (N_1079,N_914,N_912);
nor U1080 (N_1080,N_979,N_940);
or U1081 (N_1081,N_938,N_901);
or U1082 (N_1082,N_967,N_983);
nand U1083 (N_1083,N_966,N_993);
and U1084 (N_1084,N_982,N_955);
or U1085 (N_1085,N_959,N_994);
nor U1086 (N_1086,N_975,N_948);
and U1087 (N_1087,N_992,N_909);
or U1088 (N_1088,N_946,N_929);
or U1089 (N_1089,N_919,N_979);
xnor U1090 (N_1090,N_924,N_971);
nor U1091 (N_1091,N_907,N_977);
nand U1092 (N_1092,N_985,N_968);
nand U1093 (N_1093,N_982,N_967);
xor U1094 (N_1094,N_965,N_974);
nor U1095 (N_1095,N_968,N_919);
nand U1096 (N_1096,N_941,N_978);
and U1097 (N_1097,N_929,N_915);
nor U1098 (N_1098,N_932,N_964);
nand U1099 (N_1099,N_947,N_995);
and U1100 (N_1100,N_1064,N_1035);
xnor U1101 (N_1101,N_1061,N_1022);
or U1102 (N_1102,N_1066,N_1077);
nor U1103 (N_1103,N_1088,N_1020);
and U1104 (N_1104,N_1001,N_1076);
nand U1105 (N_1105,N_1082,N_1039);
or U1106 (N_1106,N_1065,N_1055);
nand U1107 (N_1107,N_1034,N_1036);
or U1108 (N_1108,N_1002,N_1011);
or U1109 (N_1109,N_1083,N_1085);
nor U1110 (N_1110,N_1037,N_1071);
xor U1111 (N_1111,N_1046,N_1062);
or U1112 (N_1112,N_1049,N_1081);
nor U1113 (N_1113,N_1044,N_1008);
xor U1114 (N_1114,N_1097,N_1098);
or U1115 (N_1115,N_1089,N_1041);
and U1116 (N_1116,N_1025,N_1059);
or U1117 (N_1117,N_1043,N_1010);
nor U1118 (N_1118,N_1075,N_1080);
xor U1119 (N_1119,N_1005,N_1009);
or U1120 (N_1120,N_1090,N_1050);
nor U1121 (N_1121,N_1030,N_1069);
or U1122 (N_1122,N_1053,N_1006);
or U1123 (N_1123,N_1004,N_1094);
and U1124 (N_1124,N_1099,N_1054);
xor U1125 (N_1125,N_1029,N_1070);
and U1126 (N_1126,N_1087,N_1057);
xnor U1127 (N_1127,N_1026,N_1007);
or U1128 (N_1128,N_1096,N_1031);
nor U1129 (N_1129,N_1003,N_1078);
xor U1130 (N_1130,N_1072,N_1038);
nor U1131 (N_1131,N_1012,N_1074);
xor U1132 (N_1132,N_1033,N_1067);
nor U1133 (N_1133,N_1013,N_1024);
and U1134 (N_1134,N_1015,N_1040);
and U1135 (N_1135,N_1021,N_1051);
xor U1136 (N_1136,N_1068,N_1048);
or U1137 (N_1137,N_1091,N_1027);
xor U1138 (N_1138,N_1019,N_1014);
nand U1139 (N_1139,N_1092,N_1017);
xor U1140 (N_1140,N_1045,N_1095);
xnor U1141 (N_1141,N_1018,N_1042);
or U1142 (N_1142,N_1052,N_1079);
nand U1143 (N_1143,N_1047,N_1063);
nor U1144 (N_1144,N_1016,N_1000);
xor U1145 (N_1145,N_1028,N_1032);
and U1146 (N_1146,N_1084,N_1058);
xnor U1147 (N_1147,N_1073,N_1086);
xnor U1148 (N_1148,N_1093,N_1060);
xnor U1149 (N_1149,N_1023,N_1056);
and U1150 (N_1150,N_1011,N_1034);
or U1151 (N_1151,N_1076,N_1027);
or U1152 (N_1152,N_1082,N_1018);
nor U1153 (N_1153,N_1008,N_1064);
nor U1154 (N_1154,N_1089,N_1008);
nand U1155 (N_1155,N_1008,N_1002);
or U1156 (N_1156,N_1005,N_1082);
nand U1157 (N_1157,N_1015,N_1068);
nand U1158 (N_1158,N_1056,N_1030);
nor U1159 (N_1159,N_1084,N_1081);
and U1160 (N_1160,N_1052,N_1004);
nor U1161 (N_1161,N_1083,N_1067);
or U1162 (N_1162,N_1064,N_1084);
or U1163 (N_1163,N_1073,N_1047);
nand U1164 (N_1164,N_1070,N_1015);
or U1165 (N_1165,N_1069,N_1092);
or U1166 (N_1166,N_1013,N_1058);
nand U1167 (N_1167,N_1019,N_1011);
xnor U1168 (N_1168,N_1063,N_1026);
xor U1169 (N_1169,N_1079,N_1081);
nand U1170 (N_1170,N_1033,N_1074);
or U1171 (N_1171,N_1007,N_1016);
or U1172 (N_1172,N_1083,N_1088);
or U1173 (N_1173,N_1074,N_1078);
or U1174 (N_1174,N_1054,N_1073);
nand U1175 (N_1175,N_1019,N_1082);
nor U1176 (N_1176,N_1009,N_1011);
xnor U1177 (N_1177,N_1051,N_1082);
nand U1178 (N_1178,N_1064,N_1025);
and U1179 (N_1179,N_1010,N_1023);
and U1180 (N_1180,N_1003,N_1070);
or U1181 (N_1181,N_1028,N_1067);
and U1182 (N_1182,N_1074,N_1031);
nor U1183 (N_1183,N_1068,N_1097);
nand U1184 (N_1184,N_1012,N_1029);
nor U1185 (N_1185,N_1077,N_1064);
or U1186 (N_1186,N_1072,N_1021);
xnor U1187 (N_1187,N_1077,N_1020);
or U1188 (N_1188,N_1021,N_1029);
xnor U1189 (N_1189,N_1046,N_1013);
nand U1190 (N_1190,N_1092,N_1015);
nand U1191 (N_1191,N_1007,N_1069);
nor U1192 (N_1192,N_1055,N_1061);
and U1193 (N_1193,N_1065,N_1010);
or U1194 (N_1194,N_1047,N_1017);
nand U1195 (N_1195,N_1043,N_1019);
nor U1196 (N_1196,N_1043,N_1068);
and U1197 (N_1197,N_1077,N_1005);
nand U1198 (N_1198,N_1020,N_1049);
nor U1199 (N_1199,N_1007,N_1097);
nand U1200 (N_1200,N_1192,N_1160);
and U1201 (N_1201,N_1198,N_1133);
nor U1202 (N_1202,N_1171,N_1187);
and U1203 (N_1203,N_1101,N_1175);
xor U1204 (N_1204,N_1156,N_1106);
or U1205 (N_1205,N_1137,N_1132);
xnor U1206 (N_1206,N_1193,N_1141);
xor U1207 (N_1207,N_1186,N_1107);
xnor U1208 (N_1208,N_1102,N_1168);
nand U1209 (N_1209,N_1151,N_1154);
xor U1210 (N_1210,N_1169,N_1144);
nand U1211 (N_1211,N_1170,N_1134);
nand U1212 (N_1212,N_1138,N_1181);
or U1213 (N_1213,N_1123,N_1100);
nor U1214 (N_1214,N_1174,N_1108);
and U1215 (N_1215,N_1176,N_1190);
and U1216 (N_1216,N_1196,N_1185);
and U1217 (N_1217,N_1104,N_1128);
nand U1218 (N_1218,N_1164,N_1183);
nor U1219 (N_1219,N_1140,N_1112);
nor U1220 (N_1220,N_1149,N_1110);
nand U1221 (N_1221,N_1109,N_1199);
xnor U1222 (N_1222,N_1194,N_1162);
nor U1223 (N_1223,N_1166,N_1145);
or U1224 (N_1224,N_1136,N_1130);
or U1225 (N_1225,N_1191,N_1184);
or U1226 (N_1226,N_1182,N_1165);
and U1227 (N_1227,N_1167,N_1143);
and U1228 (N_1228,N_1139,N_1147);
and U1229 (N_1229,N_1142,N_1116);
nand U1230 (N_1230,N_1111,N_1157);
and U1231 (N_1231,N_1161,N_1188);
xor U1232 (N_1232,N_1163,N_1129);
or U1233 (N_1233,N_1153,N_1113);
nor U1234 (N_1234,N_1177,N_1121);
and U1235 (N_1235,N_1179,N_1173);
or U1236 (N_1236,N_1158,N_1189);
nor U1237 (N_1237,N_1105,N_1127);
nor U1238 (N_1238,N_1124,N_1114);
nand U1239 (N_1239,N_1197,N_1117);
nor U1240 (N_1240,N_1118,N_1126);
xor U1241 (N_1241,N_1146,N_1135);
or U1242 (N_1242,N_1180,N_1115);
and U1243 (N_1243,N_1122,N_1125);
and U1244 (N_1244,N_1148,N_1150);
and U1245 (N_1245,N_1120,N_1178);
or U1246 (N_1246,N_1159,N_1152);
nor U1247 (N_1247,N_1172,N_1131);
or U1248 (N_1248,N_1103,N_1155);
xnor U1249 (N_1249,N_1195,N_1119);
nand U1250 (N_1250,N_1186,N_1153);
nor U1251 (N_1251,N_1150,N_1192);
and U1252 (N_1252,N_1111,N_1191);
or U1253 (N_1253,N_1182,N_1179);
nand U1254 (N_1254,N_1185,N_1107);
and U1255 (N_1255,N_1150,N_1120);
or U1256 (N_1256,N_1151,N_1148);
nand U1257 (N_1257,N_1165,N_1124);
nand U1258 (N_1258,N_1135,N_1128);
or U1259 (N_1259,N_1112,N_1158);
xnor U1260 (N_1260,N_1154,N_1194);
nor U1261 (N_1261,N_1157,N_1125);
nor U1262 (N_1262,N_1109,N_1104);
nand U1263 (N_1263,N_1174,N_1112);
nor U1264 (N_1264,N_1123,N_1128);
xnor U1265 (N_1265,N_1109,N_1146);
nor U1266 (N_1266,N_1120,N_1164);
and U1267 (N_1267,N_1180,N_1114);
xnor U1268 (N_1268,N_1121,N_1100);
and U1269 (N_1269,N_1148,N_1152);
nor U1270 (N_1270,N_1133,N_1108);
nor U1271 (N_1271,N_1114,N_1137);
or U1272 (N_1272,N_1170,N_1115);
nand U1273 (N_1273,N_1124,N_1143);
nand U1274 (N_1274,N_1133,N_1158);
or U1275 (N_1275,N_1133,N_1113);
nor U1276 (N_1276,N_1155,N_1134);
or U1277 (N_1277,N_1141,N_1153);
or U1278 (N_1278,N_1156,N_1162);
or U1279 (N_1279,N_1147,N_1173);
xnor U1280 (N_1280,N_1138,N_1174);
xnor U1281 (N_1281,N_1105,N_1129);
and U1282 (N_1282,N_1190,N_1187);
or U1283 (N_1283,N_1116,N_1102);
or U1284 (N_1284,N_1193,N_1125);
and U1285 (N_1285,N_1112,N_1199);
xnor U1286 (N_1286,N_1171,N_1115);
and U1287 (N_1287,N_1116,N_1194);
xor U1288 (N_1288,N_1193,N_1161);
or U1289 (N_1289,N_1173,N_1171);
or U1290 (N_1290,N_1179,N_1172);
or U1291 (N_1291,N_1191,N_1170);
xnor U1292 (N_1292,N_1150,N_1100);
nor U1293 (N_1293,N_1166,N_1117);
nand U1294 (N_1294,N_1156,N_1175);
nand U1295 (N_1295,N_1113,N_1134);
nand U1296 (N_1296,N_1104,N_1148);
or U1297 (N_1297,N_1172,N_1195);
nor U1298 (N_1298,N_1142,N_1168);
nor U1299 (N_1299,N_1102,N_1126);
xor U1300 (N_1300,N_1290,N_1254);
and U1301 (N_1301,N_1240,N_1253);
nand U1302 (N_1302,N_1204,N_1270);
xnor U1303 (N_1303,N_1241,N_1209);
and U1304 (N_1304,N_1281,N_1247);
xnor U1305 (N_1305,N_1268,N_1267);
nor U1306 (N_1306,N_1231,N_1215);
and U1307 (N_1307,N_1266,N_1255);
nand U1308 (N_1308,N_1216,N_1246);
nand U1309 (N_1309,N_1202,N_1258);
or U1310 (N_1310,N_1276,N_1272);
nand U1311 (N_1311,N_1286,N_1210);
or U1312 (N_1312,N_1252,N_1248);
nand U1313 (N_1313,N_1282,N_1298);
nand U1314 (N_1314,N_1284,N_1223);
xor U1315 (N_1315,N_1283,N_1274);
xor U1316 (N_1316,N_1294,N_1278);
nand U1317 (N_1317,N_1293,N_1203);
xnor U1318 (N_1318,N_1295,N_1201);
nor U1319 (N_1319,N_1296,N_1233);
nor U1320 (N_1320,N_1229,N_1292);
or U1321 (N_1321,N_1273,N_1228);
xnor U1322 (N_1322,N_1242,N_1227);
nand U1323 (N_1323,N_1297,N_1299);
and U1324 (N_1324,N_1269,N_1262);
nor U1325 (N_1325,N_1219,N_1256);
xor U1326 (N_1326,N_1275,N_1200);
nor U1327 (N_1327,N_1237,N_1208);
nand U1328 (N_1328,N_1250,N_1260);
xor U1329 (N_1329,N_1285,N_1206);
or U1330 (N_1330,N_1279,N_1277);
and U1331 (N_1331,N_1265,N_1288);
nor U1332 (N_1332,N_1222,N_1232);
or U1333 (N_1333,N_1257,N_1205);
xor U1334 (N_1334,N_1207,N_1289);
xnor U1335 (N_1335,N_1212,N_1236);
nor U1336 (N_1336,N_1271,N_1244);
nand U1337 (N_1337,N_1243,N_1224);
xnor U1338 (N_1338,N_1211,N_1218);
xor U1339 (N_1339,N_1249,N_1226);
and U1340 (N_1340,N_1263,N_1234);
or U1341 (N_1341,N_1259,N_1239);
and U1342 (N_1342,N_1280,N_1264);
or U1343 (N_1343,N_1213,N_1221);
and U1344 (N_1344,N_1261,N_1245);
xnor U1345 (N_1345,N_1235,N_1214);
or U1346 (N_1346,N_1287,N_1291);
and U1347 (N_1347,N_1217,N_1251);
xor U1348 (N_1348,N_1238,N_1230);
and U1349 (N_1349,N_1220,N_1225);
or U1350 (N_1350,N_1210,N_1255);
nand U1351 (N_1351,N_1219,N_1289);
xor U1352 (N_1352,N_1278,N_1212);
nand U1353 (N_1353,N_1287,N_1286);
and U1354 (N_1354,N_1280,N_1226);
nand U1355 (N_1355,N_1237,N_1260);
nand U1356 (N_1356,N_1254,N_1241);
nor U1357 (N_1357,N_1205,N_1266);
and U1358 (N_1358,N_1232,N_1247);
or U1359 (N_1359,N_1253,N_1257);
or U1360 (N_1360,N_1222,N_1239);
nor U1361 (N_1361,N_1255,N_1277);
and U1362 (N_1362,N_1207,N_1238);
and U1363 (N_1363,N_1252,N_1250);
or U1364 (N_1364,N_1255,N_1228);
or U1365 (N_1365,N_1225,N_1224);
xor U1366 (N_1366,N_1294,N_1238);
nor U1367 (N_1367,N_1246,N_1234);
or U1368 (N_1368,N_1206,N_1240);
xnor U1369 (N_1369,N_1265,N_1261);
or U1370 (N_1370,N_1277,N_1228);
xnor U1371 (N_1371,N_1298,N_1283);
and U1372 (N_1372,N_1272,N_1291);
nand U1373 (N_1373,N_1223,N_1267);
and U1374 (N_1374,N_1233,N_1250);
or U1375 (N_1375,N_1210,N_1298);
and U1376 (N_1376,N_1253,N_1260);
nand U1377 (N_1377,N_1294,N_1233);
and U1378 (N_1378,N_1286,N_1202);
and U1379 (N_1379,N_1223,N_1262);
nand U1380 (N_1380,N_1202,N_1234);
or U1381 (N_1381,N_1239,N_1204);
or U1382 (N_1382,N_1284,N_1206);
or U1383 (N_1383,N_1221,N_1253);
nand U1384 (N_1384,N_1221,N_1275);
nand U1385 (N_1385,N_1288,N_1296);
nand U1386 (N_1386,N_1208,N_1249);
xnor U1387 (N_1387,N_1284,N_1296);
nor U1388 (N_1388,N_1276,N_1237);
xnor U1389 (N_1389,N_1218,N_1294);
xor U1390 (N_1390,N_1208,N_1244);
nand U1391 (N_1391,N_1208,N_1238);
or U1392 (N_1392,N_1259,N_1210);
and U1393 (N_1393,N_1253,N_1270);
xor U1394 (N_1394,N_1289,N_1299);
nor U1395 (N_1395,N_1240,N_1285);
nor U1396 (N_1396,N_1255,N_1275);
xnor U1397 (N_1397,N_1272,N_1278);
nand U1398 (N_1398,N_1270,N_1263);
or U1399 (N_1399,N_1254,N_1209);
nor U1400 (N_1400,N_1369,N_1381);
xnor U1401 (N_1401,N_1397,N_1361);
and U1402 (N_1402,N_1313,N_1391);
or U1403 (N_1403,N_1390,N_1396);
nand U1404 (N_1404,N_1387,N_1399);
or U1405 (N_1405,N_1309,N_1311);
and U1406 (N_1406,N_1373,N_1380);
xnor U1407 (N_1407,N_1314,N_1322);
nand U1408 (N_1408,N_1372,N_1333);
and U1409 (N_1409,N_1340,N_1358);
nand U1410 (N_1410,N_1303,N_1356);
or U1411 (N_1411,N_1308,N_1329);
nor U1412 (N_1412,N_1324,N_1365);
nor U1413 (N_1413,N_1343,N_1338);
xnor U1414 (N_1414,N_1346,N_1341);
and U1415 (N_1415,N_1325,N_1378);
and U1416 (N_1416,N_1382,N_1353);
xor U1417 (N_1417,N_1319,N_1334);
nor U1418 (N_1418,N_1331,N_1337);
xnor U1419 (N_1419,N_1323,N_1348);
or U1420 (N_1420,N_1398,N_1371);
nand U1421 (N_1421,N_1302,N_1394);
nor U1422 (N_1422,N_1367,N_1389);
or U1423 (N_1423,N_1363,N_1347);
nor U1424 (N_1424,N_1352,N_1386);
nor U1425 (N_1425,N_1315,N_1330);
and U1426 (N_1426,N_1335,N_1359);
nor U1427 (N_1427,N_1332,N_1326);
xor U1428 (N_1428,N_1317,N_1364);
and U1429 (N_1429,N_1357,N_1354);
xnor U1430 (N_1430,N_1306,N_1327);
xnor U1431 (N_1431,N_1384,N_1374);
nor U1432 (N_1432,N_1320,N_1392);
xnor U1433 (N_1433,N_1370,N_1349);
nor U1434 (N_1434,N_1344,N_1305);
nand U1435 (N_1435,N_1301,N_1312);
nor U1436 (N_1436,N_1388,N_1366);
and U1437 (N_1437,N_1304,N_1307);
nor U1438 (N_1438,N_1318,N_1383);
xnor U1439 (N_1439,N_1376,N_1300);
nor U1440 (N_1440,N_1379,N_1393);
or U1441 (N_1441,N_1360,N_1339);
or U1442 (N_1442,N_1336,N_1375);
and U1443 (N_1443,N_1362,N_1316);
and U1444 (N_1444,N_1351,N_1342);
nor U1445 (N_1445,N_1310,N_1321);
and U1446 (N_1446,N_1345,N_1355);
nand U1447 (N_1447,N_1377,N_1328);
or U1448 (N_1448,N_1368,N_1350);
or U1449 (N_1449,N_1385,N_1395);
xor U1450 (N_1450,N_1377,N_1346);
or U1451 (N_1451,N_1389,N_1323);
nand U1452 (N_1452,N_1366,N_1345);
or U1453 (N_1453,N_1350,N_1377);
and U1454 (N_1454,N_1390,N_1385);
or U1455 (N_1455,N_1396,N_1338);
or U1456 (N_1456,N_1318,N_1365);
nand U1457 (N_1457,N_1397,N_1309);
nor U1458 (N_1458,N_1360,N_1366);
xor U1459 (N_1459,N_1353,N_1369);
and U1460 (N_1460,N_1392,N_1351);
xor U1461 (N_1461,N_1391,N_1345);
xnor U1462 (N_1462,N_1310,N_1355);
nor U1463 (N_1463,N_1385,N_1314);
or U1464 (N_1464,N_1306,N_1339);
nand U1465 (N_1465,N_1396,N_1316);
nor U1466 (N_1466,N_1335,N_1355);
xor U1467 (N_1467,N_1333,N_1367);
nor U1468 (N_1468,N_1384,N_1332);
or U1469 (N_1469,N_1344,N_1355);
or U1470 (N_1470,N_1362,N_1340);
nor U1471 (N_1471,N_1349,N_1374);
nor U1472 (N_1472,N_1366,N_1379);
or U1473 (N_1473,N_1399,N_1352);
nor U1474 (N_1474,N_1365,N_1312);
or U1475 (N_1475,N_1307,N_1385);
nor U1476 (N_1476,N_1395,N_1352);
nor U1477 (N_1477,N_1322,N_1379);
nand U1478 (N_1478,N_1334,N_1322);
nor U1479 (N_1479,N_1383,N_1391);
and U1480 (N_1480,N_1308,N_1364);
nor U1481 (N_1481,N_1358,N_1380);
and U1482 (N_1482,N_1370,N_1396);
nor U1483 (N_1483,N_1398,N_1311);
or U1484 (N_1484,N_1381,N_1330);
nor U1485 (N_1485,N_1310,N_1368);
nand U1486 (N_1486,N_1346,N_1370);
nand U1487 (N_1487,N_1342,N_1364);
nand U1488 (N_1488,N_1333,N_1322);
nand U1489 (N_1489,N_1364,N_1379);
nor U1490 (N_1490,N_1368,N_1388);
nand U1491 (N_1491,N_1379,N_1315);
nor U1492 (N_1492,N_1379,N_1376);
nand U1493 (N_1493,N_1321,N_1373);
xnor U1494 (N_1494,N_1387,N_1372);
xor U1495 (N_1495,N_1372,N_1320);
xnor U1496 (N_1496,N_1345,N_1359);
nand U1497 (N_1497,N_1302,N_1338);
and U1498 (N_1498,N_1395,N_1327);
nor U1499 (N_1499,N_1314,N_1330);
and U1500 (N_1500,N_1406,N_1441);
or U1501 (N_1501,N_1472,N_1432);
xnor U1502 (N_1502,N_1473,N_1468);
or U1503 (N_1503,N_1435,N_1449);
xnor U1504 (N_1504,N_1481,N_1421);
or U1505 (N_1505,N_1483,N_1497);
nor U1506 (N_1506,N_1412,N_1440);
nor U1507 (N_1507,N_1451,N_1429);
and U1508 (N_1508,N_1488,N_1487);
nor U1509 (N_1509,N_1445,N_1408);
nand U1510 (N_1510,N_1477,N_1480);
nor U1511 (N_1511,N_1491,N_1409);
nor U1512 (N_1512,N_1400,N_1417);
nor U1513 (N_1513,N_1428,N_1448);
xnor U1514 (N_1514,N_1490,N_1467);
nand U1515 (N_1515,N_1456,N_1423);
nor U1516 (N_1516,N_1458,N_1434);
xnor U1517 (N_1517,N_1457,N_1413);
xnor U1518 (N_1518,N_1401,N_1460);
xnor U1519 (N_1519,N_1438,N_1419);
and U1520 (N_1520,N_1493,N_1415);
and U1521 (N_1521,N_1425,N_1465);
nor U1522 (N_1522,N_1478,N_1405);
nand U1523 (N_1523,N_1459,N_1454);
xor U1524 (N_1524,N_1424,N_1495);
nand U1525 (N_1525,N_1430,N_1422);
nor U1526 (N_1526,N_1476,N_1479);
and U1527 (N_1527,N_1410,N_1439);
and U1528 (N_1528,N_1416,N_1444);
xor U1529 (N_1529,N_1469,N_1433);
xnor U1530 (N_1530,N_1453,N_1442);
nor U1531 (N_1531,N_1466,N_1461);
and U1532 (N_1532,N_1452,N_1414);
nor U1533 (N_1533,N_1498,N_1485);
and U1534 (N_1534,N_1486,N_1492);
and U1535 (N_1535,N_1437,N_1446);
xor U1536 (N_1536,N_1420,N_1471);
or U1537 (N_1537,N_1426,N_1489);
nor U1538 (N_1538,N_1482,N_1411);
nor U1539 (N_1539,N_1418,N_1450);
nor U1540 (N_1540,N_1484,N_1431);
xnor U1541 (N_1541,N_1436,N_1403);
or U1542 (N_1542,N_1427,N_1496);
nand U1543 (N_1543,N_1455,N_1404);
nor U1544 (N_1544,N_1443,N_1464);
nand U1545 (N_1545,N_1402,N_1474);
nand U1546 (N_1546,N_1447,N_1407);
or U1547 (N_1547,N_1494,N_1499);
xor U1548 (N_1548,N_1475,N_1463);
and U1549 (N_1549,N_1470,N_1462);
nand U1550 (N_1550,N_1489,N_1402);
xor U1551 (N_1551,N_1422,N_1445);
or U1552 (N_1552,N_1419,N_1450);
nand U1553 (N_1553,N_1422,N_1478);
xnor U1554 (N_1554,N_1459,N_1410);
and U1555 (N_1555,N_1439,N_1464);
xnor U1556 (N_1556,N_1448,N_1446);
or U1557 (N_1557,N_1478,N_1414);
nor U1558 (N_1558,N_1402,N_1419);
xor U1559 (N_1559,N_1449,N_1468);
nand U1560 (N_1560,N_1411,N_1412);
and U1561 (N_1561,N_1411,N_1486);
or U1562 (N_1562,N_1416,N_1491);
or U1563 (N_1563,N_1467,N_1449);
and U1564 (N_1564,N_1485,N_1401);
nor U1565 (N_1565,N_1403,N_1437);
nand U1566 (N_1566,N_1489,N_1474);
xor U1567 (N_1567,N_1451,N_1442);
nor U1568 (N_1568,N_1498,N_1471);
xor U1569 (N_1569,N_1498,N_1423);
nand U1570 (N_1570,N_1485,N_1404);
or U1571 (N_1571,N_1476,N_1424);
nor U1572 (N_1572,N_1489,N_1419);
nand U1573 (N_1573,N_1421,N_1490);
or U1574 (N_1574,N_1434,N_1441);
and U1575 (N_1575,N_1456,N_1412);
and U1576 (N_1576,N_1400,N_1433);
nand U1577 (N_1577,N_1424,N_1400);
and U1578 (N_1578,N_1463,N_1442);
and U1579 (N_1579,N_1414,N_1407);
and U1580 (N_1580,N_1434,N_1442);
nand U1581 (N_1581,N_1465,N_1497);
and U1582 (N_1582,N_1478,N_1454);
xor U1583 (N_1583,N_1489,N_1436);
nor U1584 (N_1584,N_1434,N_1425);
xor U1585 (N_1585,N_1447,N_1490);
or U1586 (N_1586,N_1410,N_1465);
xnor U1587 (N_1587,N_1452,N_1438);
nand U1588 (N_1588,N_1430,N_1407);
xor U1589 (N_1589,N_1418,N_1457);
or U1590 (N_1590,N_1428,N_1449);
and U1591 (N_1591,N_1487,N_1484);
nand U1592 (N_1592,N_1484,N_1424);
nor U1593 (N_1593,N_1437,N_1419);
xnor U1594 (N_1594,N_1436,N_1454);
or U1595 (N_1595,N_1454,N_1483);
xor U1596 (N_1596,N_1437,N_1422);
nand U1597 (N_1597,N_1494,N_1463);
and U1598 (N_1598,N_1474,N_1433);
or U1599 (N_1599,N_1406,N_1408);
xor U1600 (N_1600,N_1578,N_1556);
or U1601 (N_1601,N_1555,N_1506);
nand U1602 (N_1602,N_1581,N_1539);
or U1603 (N_1603,N_1534,N_1508);
and U1604 (N_1604,N_1582,N_1593);
or U1605 (N_1605,N_1545,N_1527);
and U1606 (N_1606,N_1515,N_1557);
nand U1607 (N_1607,N_1513,N_1586);
nor U1608 (N_1608,N_1536,N_1559);
nor U1609 (N_1609,N_1583,N_1576);
xor U1610 (N_1610,N_1575,N_1567);
and U1611 (N_1611,N_1532,N_1503);
or U1612 (N_1612,N_1529,N_1584);
xnor U1613 (N_1613,N_1598,N_1568);
xnor U1614 (N_1614,N_1599,N_1560);
xor U1615 (N_1615,N_1591,N_1528);
xor U1616 (N_1616,N_1580,N_1590);
and U1617 (N_1617,N_1579,N_1571);
xnor U1618 (N_1618,N_1533,N_1521);
and U1619 (N_1619,N_1504,N_1572);
xor U1620 (N_1620,N_1531,N_1569);
and U1621 (N_1621,N_1552,N_1523);
nand U1622 (N_1622,N_1596,N_1562);
and U1623 (N_1623,N_1530,N_1501);
nand U1624 (N_1624,N_1519,N_1522);
or U1625 (N_1625,N_1507,N_1597);
nand U1626 (N_1626,N_1512,N_1546);
or U1627 (N_1627,N_1594,N_1505);
nor U1628 (N_1628,N_1553,N_1587);
or U1629 (N_1629,N_1585,N_1543);
and U1630 (N_1630,N_1517,N_1516);
nor U1631 (N_1631,N_1565,N_1573);
or U1632 (N_1632,N_1525,N_1514);
and U1633 (N_1633,N_1561,N_1526);
or U1634 (N_1634,N_1510,N_1563);
xnor U1635 (N_1635,N_1558,N_1588);
nor U1636 (N_1636,N_1541,N_1550);
nand U1637 (N_1637,N_1566,N_1535);
nor U1638 (N_1638,N_1511,N_1542);
xor U1639 (N_1639,N_1524,N_1574);
xnor U1640 (N_1640,N_1570,N_1548);
nand U1641 (N_1641,N_1547,N_1595);
or U1642 (N_1642,N_1500,N_1502);
xor U1643 (N_1643,N_1544,N_1554);
or U1644 (N_1644,N_1551,N_1549);
nor U1645 (N_1645,N_1564,N_1518);
nor U1646 (N_1646,N_1589,N_1509);
nand U1647 (N_1647,N_1538,N_1540);
nor U1648 (N_1648,N_1592,N_1520);
or U1649 (N_1649,N_1577,N_1537);
and U1650 (N_1650,N_1501,N_1549);
nand U1651 (N_1651,N_1527,N_1502);
xor U1652 (N_1652,N_1534,N_1530);
nor U1653 (N_1653,N_1507,N_1548);
xor U1654 (N_1654,N_1547,N_1577);
and U1655 (N_1655,N_1519,N_1568);
xnor U1656 (N_1656,N_1569,N_1519);
or U1657 (N_1657,N_1557,N_1500);
xor U1658 (N_1658,N_1529,N_1554);
or U1659 (N_1659,N_1589,N_1580);
xor U1660 (N_1660,N_1544,N_1563);
or U1661 (N_1661,N_1590,N_1505);
xor U1662 (N_1662,N_1593,N_1566);
and U1663 (N_1663,N_1533,N_1505);
xnor U1664 (N_1664,N_1575,N_1552);
nor U1665 (N_1665,N_1573,N_1599);
and U1666 (N_1666,N_1599,N_1538);
nor U1667 (N_1667,N_1538,N_1546);
and U1668 (N_1668,N_1500,N_1588);
or U1669 (N_1669,N_1549,N_1559);
xnor U1670 (N_1670,N_1593,N_1529);
nor U1671 (N_1671,N_1515,N_1550);
nor U1672 (N_1672,N_1586,N_1535);
nand U1673 (N_1673,N_1562,N_1588);
nand U1674 (N_1674,N_1544,N_1552);
xnor U1675 (N_1675,N_1592,N_1579);
xor U1676 (N_1676,N_1574,N_1552);
nor U1677 (N_1677,N_1541,N_1502);
xnor U1678 (N_1678,N_1528,N_1538);
and U1679 (N_1679,N_1572,N_1563);
nor U1680 (N_1680,N_1520,N_1593);
and U1681 (N_1681,N_1556,N_1503);
nand U1682 (N_1682,N_1519,N_1525);
nor U1683 (N_1683,N_1571,N_1525);
or U1684 (N_1684,N_1557,N_1579);
nand U1685 (N_1685,N_1590,N_1598);
or U1686 (N_1686,N_1538,N_1571);
nor U1687 (N_1687,N_1583,N_1541);
xnor U1688 (N_1688,N_1599,N_1551);
or U1689 (N_1689,N_1537,N_1542);
nor U1690 (N_1690,N_1589,N_1550);
nand U1691 (N_1691,N_1590,N_1549);
nand U1692 (N_1692,N_1566,N_1599);
xor U1693 (N_1693,N_1511,N_1557);
nand U1694 (N_1694,N_1535,N_1537);
nor U1695 (N_1695,N_1546,N_1521);
and U1696 (N_1696,N_1550,N_1503);
and U1697 (N_1697,N_1550,N_1522);
and U1698 (N_1698,N_1581,N_1576);
nand U1699 (N_1699,N_1539,N_1573);
and U1700 (N_1700,N_1683,N_1641);
nor U1701 (N_1701,N_1631,N_1689);
and U1702 (N_1702,N_1611,N_1693);
and U1703 (N_1703,N_1635,N_1640);
nand U1704 (N_1704,N_1653,N_1649);
nand U1705 (N_1705,N_1687,N_1606);
nand U1706 (N_1706,N_1696,N_1697);
nor U1707 (N_1707,N_1692,N_1691);
and U1708 (N_1708,N_1616,N_1652);
or U1709 (N_1709,N_1688,N_1698);
nand U1710 (N_1710,N_1694,N_1634);
nand U1711 (N_1711,N_1602,N_1670);
xnor U1712 (N_1712,N_1686,N_1633);
nand U1713 (N_1713,N_1672,N_1650);
nand U1714 (N_1714,N_1664,N_1646);
and U1715 (N_1715,N_1690,N_1677);
or U1716 (N_1716,N_1645,N_1699);
or U1717 (N_1717,N_1613,N_1609);
nand U1718 (N_1718,N_1623,N_1661);
xnor U1719 (N_1719,N_1695,N_1685);
and U1720 (N_1720,N_1676,N_1636);
or U1721 (N_1721,N_1674,N_1605);
or U1722 (N_1722,N_1627,N_1621);
nand U1723 (N_1723,N_1660,N_1663);
nor U1724 (N_1724,N_1600,N_1615);
xor U1725 (N_1725,N_1630,N_1607);
xnor U1726 (N_1726,N_1626,N_1603);
nor U1727 (N_1727,N_1643,N_1669);
nand U1728 (N_1728,N_1679,N_1619);
xnor U1729 (N_1729,N_1656,N_1671);
and U1730 (N_1730,N_1648,N_1637);
nand U1731 (N_1731,N_1601,N_1639);
nand U1732 (N_1732,N_1625,N_1675);
xnor U1733 (N_1733,N_1604,N_1617);
xor U1734 (N_1734,N_1651,N_1665);
nand U1735 (N_1735,N_1658,N_1644);
nand U1736 (N_1736,N_1632,N_1654);
and U1737 (N_1737,N_1682,N_1610);
and U1738 (N_1738,N_1666,N_1668);
and U1739 (N_1739,N_1673,N_1642);
and U1740 (N_1740,N_1681,N_1667);
xnor U1741 (N_1741,N_1618,N_1655);
nand U1742 (N_1742,N_1684,N_1657);
nand U1743 (N_1743,N_1612,N_1638);
xor U1744 (N_1744,N_1662,N_1622);
or U1745 (N_1745,N_1629,N_1678);
or U1746 (N_1746,N_1624,N_1680);
or U1747 (N_1747,N_1647,N_1614);
or U1748 (N_1748,N_1628,N_1620);
nand U1749 (N_1749,N_1659,N_1608);
xnor U1750 (N_1750,N_1612,N_1603);
and U1751 (N_1751,N_1649,N_1608);
and U1752 (N_1752,N_1680,N_1681);
and U1753 (N_1753,N_1678,N_1630);
nor U1754 (N_1754,N_1652,N_1637);
nand U1755 (N_1755,N_1604,N_1675);
nor U1756 (N_1756,N_1687,N_1618);
and U1757 (N_1757,N_1602,N_1682);
nand U1758 (N_1758,N_1656,N_1648);
nor U1759 (N_1759,N_1686,N_1659);
nand U1760 (N_1760,N_1624,N_1622);
and U1761 (N_1761,N_1687,N_1608);
or U1762 (N_1762,N_1650,N_1664);
nand U1763 (N_1763,N_1631,N_1672);
and U1764 (N_1764,N_1658,N_1604);
nand U1765 (N_1765,N_1637,N_1660);
nor U1766 (N_1766,N_1669,N_1636);
nor U1767 (N_1767,N_1601,N_1661);
xnor U1768 (N_1768,N_1620,N_1695);
or U1769 (N_1769,N_1671,N_1663);
or U1770 (N_1770,N_1696,N_1632);
and U1771 (N_1771,N_1642,N_1667);
nor U1772 (N_1772,N_1687,N_1631);
nor U1773 (N_1773,N_1690,N_1634);
xnor U1774 (N_1774,N_1654,N_1662);
or U1775 (N_1775,N_1627,N_1645);
and U1776 (N_1776,N_1682,N_1635);
or U1777 (N_1777,N_1655,N_1617);
and U1778 (N_1778,N_1681,N_1658);
nand U1779 (N_1779,N_1689,N_1635);
nand U1780 (N_1780,N_1636,N_1641);
and U1781 (N_1781,N_1678,N_1686);
xnor U1782 (N_1782,N_1644,N_1679);
xor U1783 (N_1783,N_1670,N_1650);
or U1784 (N_1784,N_1667,N_1621);
or U1785 (N_1785,N_1644,N_1685);
xor U1786 (N_1786,N_1619,N_1688);
xnor U1787 (N_1787,N_1684,N_1602);
or U1788 (N_1788,N_1615,N_1614);
xor U1789 (N_1789,N_1685,N_1628);
nor U1790 (N_1790,N_1691,N_1629);
nor U1791 (N_1791,N_1603,N_1695);
or U1792 (N_1792,N_1644,N_1691);
xor U1793 (N_1793,N_1665,N_1640);
xnor U1794 (N_1794,N_1616,N_1640);
and U1795 (N_1795,N_1659,N_1613);
xnor U1796 (N_1796,N_1662,N_1659);
nand U1797 (N_1797,N_1677,N_1668);
and U1798 (N_1798,N_1607,N_1624);
nand U1799 (N_1799,N_1613,N_1697);
xor U1800 (N_1800,N_1747,N_1764);
or U1801 (N_1801,N_1759,N_1741);
nor U1802 (N_1802,N_1732,N_1780);
or U1803 (N_1803,N_1726,N_1719);
or U1804 (N_1804,N_1706,N_1757);
nor U1805 (N_1805,N_1778,N_1775);
xnor U1806 (N_1806,N_1725,N_1751);
and U1807 (N_1807,N_1730,N_1761);
nand U1808 (N_1808,N_1771,N_1798);
nor U1809 (N_1809,N_1773,N_1793);
and U1810 (N_1810,N_1786,N_1738);
and U1811 (N_1811,N_1754,N_1736);
nand U1812 (N_1812,N_1745,N_1794);
and U1813 (N_1813,N_1760,N_1783);
xor U1814 (N_1814,N_1746,N_1781);
xnor U1815 (N_1815,N_1782,N_1796);
and U1816 (N_1816,N_1729,N_1717);
nand U1817 (N_1817,N_1758,N_1752);
nand U1818 (N_1818,N_1715,N_1733);
xnor U1819 (N_1819,N_1787,N_1777);
nand U1820 (N_1820,N_1756,N_1724);
xnor U1821 (N_1821,N_1767,N_1739);
or U1822 (N_1822,N_1768,N_1740);
xor U1823 (N_1823,N_1702,N_1716);
nor U1824 (N_1824,N_1711,N_1791);
or U1825 (N_1825,N_1734,N_1763);
xor U1826 (N_1826,N_1762,N_1779);
nand U1827 (N_1827,N_1755,N_1769);
xnor U1828 (N_1828,N_1721,N_1709);
xnor U1829 (N_1829,N_1765,N_1707);
and U1830 (N_1830,N_1701,N_1743);
nor U1831 (N_1831,N_1795,N_1718);
nand U1832 (N_1832,N_1723,N_1774);
xnor U1833 (N_1833,N_1735,N_1737);
or U1834 (N_1834,N_1703,N_1750);
nand U1835 (N_1835,N_1770,N_1705);
nor U1836 (N_1836,N_1784,N_1714);
or U1837 (N_1837,N_1792,N_1776);
and U1838 (N_1838,N_1722,N_1788);
xor U1839 (N_1839,N_1720,N_1797);
and U1840 (N_1840,N_1704,N_1749);
nand U1841 (N_1841,N_1766,N_1772);
or U1842 (N_1842,N_1790,N_1789);
or U1843 (N_1843,N_1744,N_1710);
and U1844 (N_1844,N_1753,N_1728);
nand U1845 (N_1845,N_1742,N_1708);
nand U1846 (N_1846,N_1712,N_1748);
or U1847 (N_1847,N_1731,N_1700);
or U1848 (N_1848,N_1785,N_1713);
or U1849 (N_1849,N_1727,N_1799);
and U1850 (N_1850,N_1728,N_1720);
or U1851 (N_1851,N_1789,N_1703);
and U1852 (N_1852,N_1766,N_1762);
and U1853 (N_1853,N_1722,N_1732);
or U1854 (N_1854,N_1703,N_1700);
nand U1855 (N_1855,N_1723,N_1752);
xor U1856 (N_1856,N_1776,N_1779);
nand U1857 (N_1857,N_1712,N_1705);
nor U1858 (N_1858,N_1707,N_1749);
and U1859 (N_1859,N_1756,N_1722);
or U1860 (N_1860,N_1770,N_1700);
xor U1861 (N_1861,N_1731,N_1776);
xor U1862 (N_1862,N_1722,N_1762);
and U1863 (N_1863,N_1763,N_1747);
xor U1864 (N_1864,N_1749,N_1736);
and U1865 (N_1865,N_1710,N_1782);
nor U1866 (N_1866,N_1735,N_1760);
nor U1867 (N_1867,N_1706,N_1762);
or U1868 (N_1868,N_1772,N_1771);
nand U1869 (N_1869,N_1707,N_1742);
nand U1870 (N_1870,N_1722,N_1780);
or U1871 (N_1871,N_1798,N_1702);
and U1872 (N_1872,N_1767,N_1792);
nand U1873 (N_1873,N_1715,N_1745);
nor U1874 (N_1874,N_1749,N_1779);
and U1875 (N_1875,N_1798,N_1787);
xnor U1876 (N_1876,N_1756,N_1787);
nor U1877 (N_1877,N_1738,N_1718);
nand U1878 (N_1878,N_1705,N_1790);
and U1879 (N_1879,N_1746,N_1757);
or U1880 (N_1880,N_1754,N_1777);
nor U1881 (N_1881,N_1722,N_1775);
nor U1882 (N_1882,N_1747,N_1767);
or U1883 (N_1883,N_1760,N_1768);
and U1884 (N_1884,N_1744,N_1785);
xor U1885 (N_1885,N_1720,N_1725);
xor U1886 (N_1886,N_1761,N_1705);
nand U1887 (N_1887,N_1776,N_1741);
xnor U1888 (N_1888,N_1776,N_1760);
nand U1889 (N_1889,N_1744,N_1789);
and U1890 (N_1890,N_1741,N_1718);
or U1891 (N_1891,N_1765,N_1764);
and U1892 (N_1892,N_1748,N_1732);
nand U1893 (N_1893,N_1782,N_1718);
xnor U1894 (N_1894,N_1787,N_1750);
or U1895 (N_1895,N_1788,N_1782);
nor U1896 (N_1896,N_1763,N_1702);
xnor U1897 (N_1897,N_1774,N_1725);
xnor U1898 (N_1898,N_1769,N_1788);
and U1899 (N_1899,N_1798,N_1790);
and U1900 (N_1900,N_1804,N_1841);
nor U1901 (N_1901,N_1879,N_1822);
nor U1902 (N_1902,N_1818,N_1894);
or U1903 (N_1903,N_1859,N_1857);
nand U1904 (N_1904,N_1816,N_1899);
nor U1905 (N_1905,N_1858,N_1836);
nand U1906 (N_1906,N_1885,N_1883);
nor U1907 (N_1907,N_1864,N_1802);
nand U1908 (N_1908,N_1846,N_1813);
and U1909 (N_1909,N_1839,N_1819);
nor U1910 (N_1910,N_1878,N_1861);
xnor U1911 (N_1911,N_1891,N_1865);
or U1912 (N_1912,N_1851,N_1853);
nor U1913 (N_1913,N_1824,N_1868);
or U1914 (N_1914,N_1863,N_1801);
nand U1915 (N_1915,N_1886,N_1848);
and U1916 (N_1916,N_1805,N_1800);
xnor U1917 (N_1917,N_1814,N_1832);
nor U1918 (N_1918,N_1809,N_1873);
nor U1919 (N_1919,N_1820,N_1874);
and U1920 (N_1920,N_1850,N_1897);
and U1921 (N_1921,N_1821,N_1896);
or U1922 (N_1922,N_1867,N_1847);
and U1923 (N_1923,N_1845,N_1881);
nor U1924 (N_1924,N_1828,N_1849);
xnor U1925 (N_1925,N_1810,N_1860);
and U1926 (N_1926,N_1869,N_1830);
nor U1927 (N_1927,N_1817,N_1815);
and U1928 (N_1928,N_1876,N_1811);
or U1929 (N_1929,N_1866,N_1843);
xnor U1930 (N_1930,N_1834,N_1871);
nand U1931 (N_1931,N_1823,N_1870);
nand U1932 (N_1932,N_1840,N_1884);
nand U1933 (N_1933,N_1888,N_1844);
and U1934 (N_1934,N_1856,N_1826);
and U1935 (N_1935,N_1835,N_1838);
xor U1936 (N_1936,N_1862,N_1837);
nand U1937 (N_1937,N_1831,N_1803);
nand U1938 (N_1938,N_1872,N_1807);
or U1939 (N_1939,N_1808,N_1898);
nor U1940 (N_1940,N_1806,N_1880);
nand U1941 (N_1941,N_1890,N_1895);
nor U1942 (N_1942,N_1833,N_1855);
xnor U1943 (N_1943,N_1892,N_1854);
nor U1944 (N_1944,N_1875,N_1877);
nand U1945 (N_1945,N_1882,N_1812);
and U1946 (N_1946,N_1889,N_1893);
nor U1947 (N_1947,N_1887,N_1825);
nor U1948 (N_1948,N_1852,N_1827);
or U1949 (N_1949,N_1842,N_1829);
nor U1950 (N_1950,N_1827,N_1828);
or U1951 (N_1951,N_1807,N_1830);
xnor U1952 (N_1952,N_1824,N_1800);
xnor U1953 (N_1953,N_1847,N_1884);
xor U1954 (N_1954,N_1864,N_1848);
or U1955 (N_1955,N_1887,N_1898);
or U1956 (N_1956,N_1852,N_1897);
xnor U1957 (N_1957,N_1812,N_1854);
and U1958 (N_1958,N_1863,N_1892);
nand U1959 (N_1959,N_1826,N_1800);
nor U1960 (N_1960,N_1863,N_1880);
or U1961 (N_1961,N_1873,N_1897);
xor U1962 (N_1962,N_1877,N_1876);
nor U1963 (N_1963,N_1820,N_1875);
and U1964 (N_1964,N_1892,N_1844);
and U1965 (N_1965,N_1801,N_1807);
nand U1966 (N_1966,N_1892,N_1845);
nor U1967 (N_1967,N_1816,N_1846);
and U1968 (N_1968,N_1841,N_1801);
nand U1969 (N_1969,N_1896,N_1878);
and U1970 (N_1970,N_1845,N_1841);
nand U1971 (N_1971,N_1861,N_1817);
nand U1972 (N_1972,N_1891,N_1876);
or U1973 (N_1973,N_1871,N_1824);
and U1974 (N_1974,N_1856,N_1839);
nand U1975 (N_1975,N_1873,N_1870);
and U1976 (N_1976,N_1838,N_1809);
and U1977 (N_1977,N_1882,N_1877);
xnor U1978 (N_1978,N_1824,N_1817);
nor U1979 (N_1979,N_1884,N_1813);
or U1980 (N_1980,N_1892,N_1873);
nor U1981 (N_1981,N_1862,N_1897);
and U1982 (N_1982,N_1848,N_1892);
or U1983 (N_1983,N_1841,N_1866);
xnor U1984 (N_1984,N_1879,N_1871);
nor U1985 (N_1985,N_1871,N_1820);
xor U1986 (N_1986,N_1891,N_1813);
nor U1987 (N_1987,N_1879,N_1870);
and U1988 (N_1988,N_1826,N_1892);
xor U1989 (N_1989,N_1818,N_1864);
xnor U1990 (N_1990,N_1876,N_1823);
or U1991 (N_1991,N_1811,N_1840);
xnor U1992 (N_1992,N_1866,N_1899);
nor U1993 (N_1993,N_1849,N_1896);
xor U1994 (N_1994,N_1862,N_1808);
and U1995 (N_1995,N_1898,N_1848);
xor U1996 (N_1996,N_1851,N_1802);
and U1997 (N_1997,N_1829,N_1801);
or U1998 (N_1998,N_1837,N_1827);
nand U1999 (N_1999,N_1837,N_1810);
nor U2000 (N_2000,N_1930,N_1921);
nand U2001 (N_2001,N_1901,N_1918);
nor U2002 (N_2002,N_1960,N_1973);
xor U2003 (N_2003,N_1925,N_1902);
nand U2004 (N_2004,N_1906,N_1942);
nor U2005 (N_2005,N_1983,N_1944);
or U2006 (N_2006,N_1933,N_1932);
and U2007 (N_2007,N_1952,N_1993);
or U2008 (N_2008,N_1994,N_1964);
nor U2009 (N_2009,N_1959,N_1957);
and U2010 (N_2010,N_1928,N_1909);
nand U2011 (N_2011,N_1910,N_1984);
or U2012 (N_2012,N_1926,N_1977);
nand U2013 (N_2013,N_1961,N_1927);
or U2014 (N_2014,N_1980,N_1978);
and U2015 (N_2015,N_1904,N_1946);
and U2016 (N_2016,N_1954,N_1951);
xnor U2017 (N_2017,N_1923,N_1945);
and U2018 (N_2018,N_1935,N_1991);
xnor U2019 (N_2019,N_1900,N_1934);
nand U2020 (N_2020,N_1986,N_1970);
and U2021 (N_2021,N_1963,N_1950);
nand U2022 (N_2022,N_1979,N_1990);
and U2023 (N_2023,N_1941,N_1943);
or U2024 (N_2024,N_1958,N_1975);
and U2025 (N_2025,N_1916,N_1968);
and U2026 (N_2026,N_1965,N_1962);
and U2027 (N_2027,N_1955,N_1936);
xnor U2028 (N_2028,N_1988,N_1924);
nand U2029 (N_2029,N_1966,N_1969);
xor U2030 (N_2030,N_1998,N_1939);
xnor U2031 (N_2031,N_1982,N_1908);
and U2032 (N_2032,N_1989,N_1919);
nor U2033 (N_2033,N_1914,N_1929);
nand U2034 (N_2034,N_1953,N_1913);
and U2035 (N_2035,N_1920,N_1985);
nor U2036 (N_2036,N_1971,N_1937);
nor U2037 (N_2037,N_1995,N_1956);
nand U2038 (N_2038,N_1940,N_1912);
nor U2039 (N_2039,N_1938,N_1997);
nand U2040 (N_2040,N_1972,N_1917);
and U2041 (N_2041,N_1903,N_1915);
or U2042 (N_2042,N_1948,N_1987);
and U2043 (N_2043,N_1976,N_1922);
and U2044 (N_2044,N_1992,N_1947);
nor U2045 (N_2045,N_1949,N_1996);
or U2046 (N_2046,N_1907,N_1905);
and U2047 (N_2047,N_1911,N_1931);
nand U2048 (N_2048,N_1981,N_1974);
or U2049 (N_2049,N_1967,N_1999);
and U2050 (N_2050,N_1927,N_1999);
or U2051 (N_2051,N_1908,N_1961);
nand U2052 (N_2052,N_1912,N_1927);
or U2053 (N_2053,N_1911,N_1983);
nand U2054 (N_2054,N_1930,N_1976);
xor U2055 (N_2055,N_1937,N_1915);
xnor U2056 (N_2056,N_1972,N_1975);
xnor U2057 (N_2057,N_1979,N_1908);
nand U2058 (N_2058,N_1964,N_1984);
nand U2059 (N_2059,N_1947,N_1995);
or U2060 (N_2060,N_1936,N_1964);
xor U2061 (N_2061,N_1983,N_1943);
nand U2062 (N_2062,N_1992,N_1995);
xor U2063 (N_2063,N_1908,N_1903);
and U2064 (N_2064,N_1928,N_1935);
nand U2065 (N_2065,N_1915,N_1967);
nor U2066 (N_2066,N_1984,N_1939);
nor U2067 (N_2067,N_1965,N_1979);
xor U2068 (N_2068,N_1960,N_1994);
and U2069 (N_2069,N_1940,N_1963);
nand U2070 (N_2070,N_1973,N_1906);
nand U2071 (N_2071,N_1989,N_1929);
nor U2072 (N_2072,N_1928,N_1963);
or U2073 (N_2073,N_1979,N_1964);
and U2074 (N_2074,N_1958,N_1994);
and U2075 (N_2075,N_1954,N_1940);
or U2076 (N_2076,N_1960,N_1977);
xnor U2077 (N_2077,N_1970,N_1925);
and U2078 (N_2078,N_1917,N_1944);
xnor U2079 (N_2079,N_1968,N_1955);
nor U2080 (N_2080,N_1931,N_1902);
nor U2081 (N_2081,N_1918,N_1943);
nand U2082 (N_2082,N_1952,N_1958);
nor U2083 (N_2083,N_1952,N_1930);
and U2084 (N_2084,N_1993,N_1909);
or U2085 (N_2085,N_1925,N_1936);
or U2086 (N_2086,N_1984,N_1905);
nand U2087 (N_2087,N_1973,N_1904);
and U2088 (N_2088,N_1973,N_1926);
or U2089 (N_2089,N_1922,N_1975);
and U2090 (N_2090,N_1920,N_1989);
nand U2091 (N_2091,N_1964,N_1970);
nor U2092 (N_2092,N_1917,N_1947);
and U2093 (N_2093,N_1932,N_1909);
xor U2094 (N_2094,N_1923,N_1908);
nor U2095 (N_2095,N_1928,N_1990);
and U2096 (N_2096,N_1975,N_1974);
nand U2097 (N_2097,N_1947,N_1931);
xor U2098 (N_2098,N_1976,N_1926);
nor U2099 (N_2099,N_1982,N_1995);
xor U2100 (N_2100,N_2011,N_2049);
nor U2101 (N_2101,N_2027,N_2046);
xnor U2102 (N_2102,N_2052,N_2085);
nor U2103 (N_2103,N_2078,N_2028);
xor U2104 (N_2104,N_2072,N_2096);
xor U2105 (N_2105,N_2013,N_2068);
nor U2106 (N_2106,N_2038,N_2000);
nor U2107 (N_2107,N_2092,N_2051);
nand U2108 (N_2108,N_2026,N_2082);
nor U2109 (N_2109,N_2083,N_2017);
xor U2110 (N_2110,N_2019,N_2097);
or U2111 (N_2111,N_2012,N_2006);
nand U2112 (N_2112,N_2075,N_2089);
or U2113 (N_2113,N_2067,N_2073);
or U2114 (N_2114,N_2070,N_2001);
and U2115 (N_2115,N_2015,N_2080);
and U2116 (N_2116,N_2009,N_2039);
nor U2117 (N_2117,N_2064,N_2054);
and U2118 (N_2118,N_2030,N_2081);
xnor U2119 (N_2119,N_2098,N_2016);
nand U2120 (N_2120,N_2093,N_2035);
nand U2121 (N_2121,N_2018,N_2084);
and U2122 (N_2122,N_2074,N_2050);
nand U2123 (N_2123,N_2020,N_2061);
and U2124 (N_2124,N_2010,N_2056);
or U2125 (N_2125,N_2058,N_2053);
or U2126 (N_2126,N_2004,N_2029);
or U2127 (N_2127,N_2099,N_2040);
or U2128 (N_2128,N_2062,N_2095);
and U2129 (N_2129,N_2032,N_2069);
xor U2130 (N_2130,N_2076,N_2021);
nor U2131 (N_2131,N_2079,N_2007);
and U2132 (N_2132,N_2065,N_2091);
nor U2133 (N_2133,N_2025,N_2086);
and U2134 (N_2134,N_2063,N_2002);
and U2135 (N_2135,N_2059,N_2005);
and U2136 (N_2136,N_2044,N_2008);
nor U2137 (N_2137,N_2077,N_2042);
xor U2138 (N_2138,N_2045,N_2090);
and U2139 (N_2139,N_2022,N_2037);
or U2140 (N_2140,N_2033,N_2094);
and U2141 (N_2141,N_2031,N_2066);
or U2142 (N_2142,N_2055,N_2088);
or U2143 (N_2143,N_2034,N_2041);
and U2144 (N_2144,N_2071,N_2014);
nor U2145 (N_2145,N_2087,N_2047);
nor U2146 (N_2146,N_2023,N_2043);
nand U2147 (N_2147,N_2057,N_2036);
and U2148 (N_2148,N_2048,N_2024);
nor U2149 (N_2149,N_2003,N_2060);
or U2150 (N_2150,N_2065,N_2017);
nand U2151 (N_2151,N_2009,N_2042);
nand U2152 (N_2152,N_2059,N_2097);
xor U2153 (N_2153,N_2060,N_2013);
or U2154 (N_2154,N_2076,N_2015);
nor U2155 (N_2155,N_2057,N_2030);
and U2156 (N_2156,N_2029,N_2022);
xnor U2157 (N_2157,N_2010,N_2009);
nor U2158 (N_2158,N_2086,N_2063);
xnor U2159 (N_2159,N_2059,N_2074);
nor U2160 (N_2160,N_2098,N_2084);
and U2161 (N_2161,N_2083,N_2062);
nor U2162 (N_2162,N_2022,N_2039);
xnor U2163 (N_2163,N_2040,N_2012);
or U2164 (N_2164,N_2037,N_2085);
and U2165 (N_2165,N_2010,N_2076);
or U2166 (N_2166,N_2048,N_2097);
nor U2167 (N_2167,N_2029,N_2030);
and U2168 (N_2168,N_2028,N_2008);
xnor U2169 (N_2169,N_2068,N_2012);
nor U2170 (N_2170,N_2057,N_2046);
nor U2171 (N_2171,N_2082,N_2081);
and U2172 (N_2172,N_2018,N_2033);
nor U2173 (N_2173,N_2000,N_2006);
nand U2174 (N_2174,N_2041,N_2059);
nand U2175 (N_2175,N_2071,N_2029);
xnor U2176 (N_2176,N_2003,N_2020);
nor U2177 (N_2177,N_2075,N_2080);
or U2178 (N_2178,N_2075,N_2098);
nor U2179 (N_2179,N_2047,N_2058);
nor U2180 (N_2180,N_2015,N_2074);
xor U2181 (N_2181,N_2067,N_2039);
or U2182 (N_2182,N_2096,N_2093);
and U2183 (N_2183,N_2069,N_2096);
xnor U2184 (N_2184,N_2047,N_2033);
and U2185 (N_2185,N_2004,N_2047);
or U2186 (N_2186,N_2053,N_2074);
nor U2187 (N_2187,N_2044,N_2002);
and U2188 (N_2188,N_2021,N_2058);
nand U2189 (N_2189,N_2024,N_2099);
nand U2190 (N_2190,N_2016,N_2086);
nor U2191 (N_2191,N_2066,N_2053);
nor U2192 (N_2192,N_2076,N_2095);
nand U2193 (N_2193,N_2018,N_2037);
or U2194 (N_2194,N_2006,N_2063);
xor U2195 (N_2195,N_2000,N_2037);
xnor U2196 (N_2196,N_2016,N_2076);
and U2197 (N_2197,N_2089,N_2046);
nor U2198 (N_2198,N_2069,N_2055);
xor U2199 (N_2199,N_2069,N_2062);
or U2200 (N_2200,N_2138,N_2173);
xnor U2201 (N_2201,N_2139,N_2132);
or U2202 (N_2202,N_2199,N_2108);
or U2203 (N_2203,N_2172,N_2113);
or U2204 (N_2204,N_2122,N_2144);
or U2205 (N_2205,N_2129,N_2106);
and U2206 (N_2206,N_2186,N_2162);
nand U2207 (N_2207,N_2116,N_2127);
or U2208 (N_2208,N_2150,N_2120);
or U2209 (N_2209,N_2149,N_2174);
nand U2210 (N_2210,N_2185,N_2187);
or U2211 (N_2211,N_2126,N_2117);
or U2212 (N_2212,N_2176,N_2131);
or U2213 (N_2213,N_2181,N_2121);
nand U2214 (N_2214,N_2133,N_2182);
nor U2215 (N_2215,N_2195,N_2103);
nor U2216 (N_2216,N_2165,N_2153);
and U2217 (N_2217,N_2169,N_2119);
nand U2218 (N_2218,N_2192,N_2175);
xor U2219 (N_2219,N_2107,N_2137);
nand U2220 (N_2220,N_2111,N_2167);
and U2221 (N_2221,N_2100,N_2171);
xor U2222 (N_2222,N_2189,N_2188);
or U2223 (N_2223,N_2164,N_2105);
xor U2224 (N_2224,N_2141,N_2142);
nand U2225 (N_2225,N_2114,N_2184);
nor U2226 (N_2226,N_2193,N_2191);
or U2227 (N_2227,N_2115,N_2148);
xnor U2228 (N_2228,N_2158,N_2123);
xnor U2229 (N_2229,N_2163,N_2170);
nand U2230 (N_2230,N_2112,N_2135);
xnor U2231 (N_2231,N_2166,N_2194);
and U2232 (N_2232,N_2140,N_2161);
nor U2233 (N_2233,N_2128,N_2190);
or U2234 (N_2234,N_2179,N_2160);
nand U2235 (N_2235,N_2147,N_2143);
and U2236 (N_2236,N_2102,N_2198);
nor U2237 (N_2237,N_2151,N_2146);
xnor U2238 (N_2238,N_2136,N_2109);
and U2239 (N_2239,N_2110,N_2197);
or U2240 (N_2240,N_2134,N_2180);
or U2241 (N_2241,N_2101,N_2196);
or U2242 (N_2242,N_2168,N_2156);
nor U2243 (N_2243,N_2125,N_2124);
and U2244 (N_2244,N_2118,N_2152);
xor U2245 (N_2245,N_2130,N_2104);
xor U2246 (N_2246,N_2159,N_2154);
and U2247 (N_2247,N_2177,N_2145);
xor U2248 (N_2248,N_2157,N_2155);
nand U2249 (N_2249,N_2178,N_2183);
xor U2250 (N_2250,N_2145,N_2138);
xnor U2251 (N_2251,N_2187,N_2177);
xnor U2252 (N_2252,N_2134,N_2141);
xnor U2253 (N_2253,N_2112,N_2199);
nor U2254 (N_2254,N_2190,N_2197);
and U2255 (N_2255,N_2194,N_2165);
or U2256 (N_2256,N_2126,N_2172);
xnor U2257 (N_2257,N_2151,N_2133);
and U2258 (N_2258,N_2136,N_2163);
or U2259 (N_2259,N_2166,N_2176);
xor U2260 (N_2260,N_2180,N_2141);
or U2261 (N_2261,N_2151,N_2125);
and U2262 (N_2262,N_2168,N_2196);
nand U2263 (N_2263,N_2133,N_2165);
and U2264 (N_2264,N_2101,N_2135);
xor U2265 (N_2265,N_2106,N_2137);
xnor U2266 (N_2266,N_2128,N_2197);
xnor U2267 (N_2267,N_2196,N_2185);
xor U2268 (N_2268,N_2175,N_2199);
nor U2269 (N_2269,N_2116,N_2146);
nand U2270 (N_2270,N_2148,N_2161);
or U2271 (N_2271,N_2186,N_2108);
nor U2272 (N_2272,N_2162,N_2155);
xor U2273 (N_2273,N_2131,N_2121);
or U2274 (N_2274,N_2151,N_2118);
xor U2275 (N_2275,N_2186,N_2128);
xor U2276 (N_2276,N_2145,N_2169);
xnor U2277 (N_2277,N_2125,N_2183);
nand U2278 (N_2278,N_2147,N_2111);
nor U2279 (N_2279,N_2117,N_2173);
nor U2280 (N_2280,N_2115,N_2130);
xnor U2281 (N_2281,N_2125,N_2133);
xnor U2282 (N_2282,N_2184,N_2197);
nor U2283 (N_2283,N_2117,N_2114);
and U2284 (N_2284,N_2165,N_2132);
nand U2285 (N_2285,N_2173,N_2172);
or U2286 (N_2286,N_2135,N_2120);
and U2287 (N_2287,N_2169,N_2171);
nand U2288 (N_2288,N_2138,N_2190);
nand U2289 (N_2289,N_2177,N_2138);
nor U2290 (N_2290,N_2138,N_2117);
nand U2291 (N_2291,N_2142,N_2183);
or U2292 (N_2292,N_2193,N_2142);
nand U2293 (N_2293,N_2103,N_2180);
and U2294 (N_2294,N_2127,N_2112);
or U2295 (N_2295,N_2151,N_2185);
nor U2296 (N_2296,N_2102,N_2143);
or U2297 (N_2297,N_2170,N_2193);
nand U2298 (N_2298,N_2159,N_2136);
xor U2299 (N_2299,N_2197,N_2121);
or U2300 (N_2300,N_2289,N_2222);
nand U2301 (N_2301,N_2291,N_2205);
nand U2302 (N_2302,N_2251,N_2252);
nor U2303 (N_2303,N_2260,N_2295);
nor U2304 (N_2304,N_2274,N_2263);
nor U2305 (N_2305,N_2265,N_2266);
and U2306 (N_2306,N_2284,N_2209);
nand U2307 (N_2307,N_2206,N_2243);
xnor U2308 (N_2308,N_2228,N_2277);
xnor U2309 (N_2309,N_2221,N_2238);
or U2310 (N_2310,N_2246,N_2210);
or U2311 (N_2311,N_2208,N_2281);
and U2312 (N_2312,N_2256,N_2283);
xnor U2313 (N_2313,N_2247,N_2226);
and U2314 (N_2314,N_2200,N_2232);
nor U2315 (N_2315,N_2239,N_2285);
or U2316 (N_2316,N_2297,N_2223);
nand U2317 (N_2317,N_2287,N_2257);
xor U2318 (N_2318,N_2264,N_2234);
nor U2319 (N_2319,N_2261,N_2279);
and U2320 (N_2320,N_2288,N_2290);
or U2321 (N_2321,N_2227,N_2278);
xor U2322 (N_2322,N_2203,N_2224);
xnor U2323 (N_2323,N_2282,N_2280);
nor U2324 (N_2324,N_2244,N_2270);
nand U2325 (N_2325,N_2214,N_2201);
nand U2326 (N_2326,N_2230,N_2253);
xnor U2327 (N_2327,N_2235,N_2215);
nor U2328 (N_2328,N_2237,N_2250);
or U2329 (N_2329,N_2218,N_2204);
nor U2330 (N_2330,N_2272,N_2236);
xnor U2331 (N_2331,N_2217,N_2271);
nor U2332 (N_2332,N_2273,N_2219);
xnor U2333 (N_2333,N_2259,N_2292);
nor U2334 (N_2334,N_2220,N_2229);
xnor U2335 (N_2335,N_2245,N_2213);
and U2336 (N_2336,N_2267,N_2225);
and U2337 (N_2337,N_2276,N_2216);
nand U2338 (N_2338,N_2298,N_2258);
nand U2339 (N_2339,N_2211,N_2286);
nor U2340 (N_2340,N_2296,N_2233);
nor U2341 (N_2341,N_2268,N_2248);
xnor U2342 (N_2342,N_2249,N_2212);
and U2343 (N_2343,N_2293,N_2275);
nand U2344 (N_2344,N_2255,N_2262);
nand U2345 (N_2345,N_2202,N_2294);
nand U2346 (N_2346,N_2269,N_2299);
and U2347 (N_2347,N_2231,N_2207);
or U2348 (N_2348,N_2242,N_2241);
xor U2349 (N_2349,N_2254,N_2240);
nor U2350 (N_2350,N_2213,N_2210);
nand U2351 (N_2351,N_2208,N_2236);
xor U2352 (N_2352,N_2237,N_2272);
or U2353 (N_2353,N_2248,N_2231);
xnor U2354 (N_2354,N_2264,N_2210);
xor U2355 (N_2355,N_2256,N_2275);
nor U2356 (N_2356,N_2280,N_2243);
xnor U2357 (N_2357,N_2243,N_2235);
nor U2358 (N_2358,N_2233,N_2287);
and U2359 (N_2359,N_2247,N_2216);
nor U2360 (N_2360,N_2220,N_2280);
and U2361 (N_2361,N_2276,N_2240);
nor U2362 (N_2362,N_2221,N_2262);
nand U2363 (N_2363,N_2224,N_2220);
or U2364 (N_2364,N_2237,N_2218);
and U2365 (N_2365,N_2202,N_2237);
nor U2366 (N_2366,N_2280,N_2277);
and U2367 (N_2367,N_2291,N_2276);
nand U2368 (N_2368,N_2248,N_2208);
or U2369 (N_2369,N_2226,N_2260);
or U2370 (N_2370,N_2207,N_2253);
xor U2371 (N_2371,N_2247,N_2218);
nand U2372 (N_2372,N_2201,N_2241);
or U2373 (N_2373,N_2250,N_2222);
and U2374 (N_2374,N_2267,N_2292);
and U2375 (N_2375,N_2221,N_2248);
xor U2376 (N_2376,N_2213,N_2254);
xnor U2377 (N_2377,N_2275,N_2224);
nor U2378 (N_2378,N_2268,N_2204);
and U2379 (N_2379,N_2205,N_2289);
and U2380 (N_2380,N_2287,N_2254);
and U2381 (N_2381,N_2218,N_2238);
xor U2382 (N_2382,N_2220,N_2201);
nor U2383 (N_2383,N_2273,N_2209);
or U2384 (N_2384,N_2230,N_2292);
or U2385 (N_2385,N_2211,N_2245);
or U2386 (N_2386,N_2282,N_2270);
xnor U2387 (N_2387,N_2254,N_2284);
and U2388 (N_2388,N_2268,N_2283);
nor U2389 (N_2389,N_2276,N_2280);
nand U2390 (N_2390,N_2281,N_2285);
or U2391 (N_2391,N_2272,N_2201);
xnor U2392 (N_2392,N_2288,N_2298);
xnor U2393 (N_2393,N_2258,N_2222);
xor U2394 (N_2394,N_2296,N_2256);
or U2395 (N_2395,N_2212,N_2224);
or U2396 (N_2396,N_2246,N_2278);
xnor U2397 (N_2397,N_2217,N_2296);
xor U2398 (N_2398,N_2242,N_2281);
nor U2399 (N_2399,N_2280,N_2269);
nand U2400 (N_2400,N_2300,N_2392);
nand U2401 (N_2401,N_2307,N_2327);
xor U2402 (N_2402,N_2365,N_2386);
nand U2403 (N_2403,N_2337,N_2324);
or U2404 (N_2404,N_2340,N_2345);
and U2405 (N_2405,N_2379,N_2305);
xnor U2406 (N_2406,N_2377,N_2397);
and U2407 (N_2407,N_2382,N_2334);
or U2408 (N_2408,N_2353,N_2389);
and U2409 (N_2409,N_2341,N_2396);
or U2410 (N_2410,N_2302,N_2380);
nor U2411 (N_2411,N_2347,N_2351);
xor U2412 (N_2412,N_2375,N_2303);
xor U2413 (N_2413,N_2306,N_2399);
nand U2414 (N_2414,N_2355,N_2391);
nand U2415 (N_2415,N_2356,N_2366);
nor U2416 (N_2416,N_2352,N_2346);
xor U2417 (N_2417,N_2398,N_2388);
nor U2418 (N_2418,N_2323,N_2372);
or U2419 (N_2419,N_2360,N_2390);
or U2420 (N_2420,N_2367,N_2363);
nand U2421 (N_2421,N_2370,N_2313);
xor U2422 (N_2422,N_2378,N_2311);
xnor U2423 (N_2423,N_2333,N_2357);
xnor U2424 (N_2424,N_2325,N_2364);
nand U2425 (N_2425,N_2374,N_2316);
nor U2426 (N_2426,N_2301,N_2385);
and U2427 (N_2427,N_2369,N_2349);
nand U2428 (N_2428,N_2381,N_2394);
or U2429 (N_2429,N_2321,N_2395);
nor U2430 (N_2430,N_2318,N_2361);
xnor U2431 (N_2431,N_2314,N_2371);
xnor U2432 (N_2432,N_2354,N_2315);
xnor U2433 (N_2433,N_2309,N_2343);
nand U2434 (N_2434,N_2308,N_2344);
xnor U2435 (N_2435,N_2383,N_2368);
xor U2436 (N_2436,N_2335,N_2319);
nand U2437 (N_2437,N_2358,N_2342);
nor U2438 (N_2438,N_2326,N_2332);
nor U2439 (N_2439,N_2330,N_2348);
or U2440 (N_2440,N_2339,N_2310);
and U2441 (N_2441,N_2384,N_2373);
nor U2442 (N_2442,N_2317,N_2387);
nand U2443 (N_2443,N_2328,N_2362);
xnor U2444 (N_2444,N_2312,N_2359);
xor U2445 (N_2445,N_2304,N_2338);
xor U2446 (N_2446,N_2393,N_2329);
nand U2447 (N_2447,N_2376,N_2331);
nand U2448 (N_2448,N_2336,N_2322);
or U2449 (N_2449,N_2320,N_2350);
xnor U2450 (N_2450,N_2334,N_2383);
xnor U2451 (N_2451,N_2369,N_2326);
nand U2452 (N_2452,N_2382,N_2355);
and U2453 (N_2453,N_2363,N_2396);
and U2454 (N_2454,N_2313,N_2331);
nand U2455 (N_2455,N_2362,N_2354);
nor U2456 (N_2456,N_2358,N_2322);
nand U2457 (N_2457,N_2326,N_2342);
nor U2458 (N_2458,N_2387,N_2321);
and U2459 (N_2459,N_2366,N_2324);
xnor U2460 (N_2460,N_2393,N_2352);
nor U2461 (N_2461,N_2335,N_2322);
nand U2462 (N_2462,N_2340,N_2374);
nand U2463 (N_2463,N_2305,N_2354);
nor U2464 (N_2464,N_2363,N_2383);
and U2465 (N_2465,N_2377,N_2384);
nand U2466 (N_2466,N_2322,N_2357);
nand U2467 (N_2467,N_2368,N_2334);
and U2468 (N_2468,N_2369,N_2307);
and U2469 (N_2469,N_2378,N_2398);
xor U2470 (N_2470,N_2367,N_2369);
and U2471 (N_2471,N_2350,N_2341);
nand U2472 (N_2472,N_2304,N_2348);
nand U2473 (N_2473,N_2369,N_2385);
xor U2474 (N_2474,N_2391,N_2328);
nand U2475 (N_2475,N_2322,N_2359);
or U2476 (N_2476,N_2360,N_2323);
xnor U2477 (N_2477,N_2342,N_2307);
nand U2478 (N_2478,N_2303,N_2314);
nand U2479 (N_2479,N_2312,N_2333);
nor U2480 (N_2480,N_2364,N_2333);
nand U2481 (N_2481,N_2345,N_2381);
nand U2482 (N_2482,N_2322,N_2303);
nand U2483 (N_2483,N_2386,N_2368);
xor U2484 (N_2484,N_2388,N_2307);
nand U2485 (N_2485,N_2379,N_2350);
or U2486 (N_2486,N_2359,N_2326);
nor U2487 (N_2487,N_2395,N_2371);
or U2488 (N_2488,N_2399,N_2303);
nor U2489 (N_2489,N_2341,N_2399);
xor U2490 (N_2490,N_2316,N_2336);
xor U2491 (N_2491,N_2399,N_2320);
xnor U2492 (N_2492,N_2392,N_2314);
or U2493 (N_2493,N_2335,N_2332);
and U2494 (N_2494,N_2338,N_2311);
xor U2495 (N_2495,N_2366,N_2375);
xnor U2496 (N_2496,N_2306,N_2377);
nor U2497 (N_2497,N_2331,N_2329);
and U2498 (N_2498,N_2377,N_2335);
nand U2499 (N_2499,N_2385,N_2395);
or U2500 (N_2500,N_2439,N_2486);
nand U2501 (N_2501,N_2432,N_2427);
nand U2502 (N_2502,N_2435,N_2431);
and U2503 (N_2503,N_2490,N_2496);
nand U2504 (N_2504,N_2423,N_2478);
xnor U2505 (N_2505,N_2416,N_2446);
nand U2506 (N_2506,N_2472,N_2499);
nor U2507 (N_2507,N_2466,N_2494);
nand U2508 (N_2508,N_2402,N_2420);
or U2509 (N_2509,N_2449,N_2400);
nand U2510 (N_2510,N_2442,N_2433);
or U2511 (N_2511,N_2497,N_2482);
nor U2512 (N_2512,N_2480,N_2414);
and U2513 (N_2513,N_2407,N_2462);
or U2514 (N_2514,N_2483,N_2463);
and U2515 (N_2515,N_2415,N_2448);
xnor U2516 (N_2516,N_2440,N_2406);
and U2517 (N_2517,N_2459,N_2451);
nand U2518 (N_2518,N_2470,N_2412);
xnor U2519 (N_2519,N_2413,N_2493);
or U2520 (N_2520,N_2488,N_2434);
nor U2521 (N_2521,N_2425,N_2473);
xor U2522 (N_2522,N_2455,N_2471);
xnor U2523 (N_2523,N_2475,N_2411);
nand U2524 (N_2524,N_2401,N_2468);
or U2525 (N_2525,N_2450,N_2487);
and U2526 (N_2526,N_2489,N_2404);
or U2527 (N_2527,N_2426,N_2476);
and U2528 (N_2528,N_2485,N_2464);
nand U2529 (N_2529,N_2460,N_2452);
xor U2530 (N_2530,N_2495,N_2403);
nor U2531 (N_2531,N_2481,N_2484);
nand U2532 (N_2532,N_2469,N_2428);
or U2533 (N_2533,N_2421,N_2458);
or U2534 (N_2534,N_2405,N_2467);
and U2535 (N_2535,N_2492,N_2479);
nand U2536 (N_2536,N_2498,N_2477);
nor U2537 (N_2537,N_2454,N_2441);
nand U2538 (N_2538,N_2418,N_2410);
or U2539 (N_2539,N_2456,N_2419);
nand U2540 (N_2540,N_2461,N_2424);
nor U2541 (N_2541,N_2408,N_2444);
or U2542 (N_2542,N_2445,N_2491);
nand U2543 (N_2543,N_2474,N_2438);
xor U2544 (N_2544,N_2409,N_2430);
nor U2545 (N_2545,N_2417,N_2443);
nor U2546 (N_2546,N_2447,N_2453);
and U2547 (N_2547,N_2429,N_2436);
xor U2548 (N_2548,N_2422,N_2437);
nor U2549 (N_2549,N_2465,N_2457);
or U2550 (N_2550,N_2461,N_2492);
nor U2551 (N_2551,N_2484,N_2406);
and U2552 (N_2552,N_2456,N_2401);
and U2553 (N_2553,N_2420,N_2478);
xor U2554 (N_2554,N_2477,N_2408);
or U2555 (N_2555,N_2453,N_2452);
xor U2556 (N_2556,N_2499,N_2449);
and U2557 (N_2557,N_2440,N_2402);
and U2558 (N_2558,N_2431,N_2414);
and U2559 (N_2559,N_2422,N_2463);
or U2560 (N_2560,N_2400,N_2406);
or U2561 (N_2561,N_2440,N_2407);
and U2562 (N_2562,N_2464,N_2486);
nor U2563 (N_2563,N_2419,N_2453);
or U2564 (N_2564,N_2414,N_2468);
xnor U2565 (N_2565,N_2440,N_2456);
nand U2566 (N_2566,N_2412,N_2478);
and U2567 (N_2567,N_2487,N_2499);
xnor U2568 (N_2568,N_2431,N_2456);
or U2569 (N_2569,N_2475,N_2423);
nand U2570 (N_2570,N_2465,N_2462);
and U2571 (N_2571,N_2464,N_2444);
and U2572 (N_2572,N_2459,N_2407);
or U2573 (N_2573,N_2476,N_2464);
or U2574 (N_2574,N_2415,N_2452);
and U2575 (N_2575,N_2406,N_2494);
nand U2576 (N_2576,N_2418,N_2470);
nand U2577 (N_2577,N_2427,N_2464);
or U2578 (N_2578,N_2492,N_2493);
nor U2579 (N_2579,N_2456,N_2402);
nor U2580 (N_2580,N_2445,N_2476);
nor U2581 (N_2581,N_2467,N_2469);
nand U2582 (N_2582,N_2451,N_2454);
nand U2583 (N_2583,N_2457,N_2479);
nand U2584 (N_2584,N_2428,N_2497);
nand U2585 (N_2585,N_2416,N_2437);
and U2586 (N_2586,N_2439,N_2450);
or U2587 (N_2587,N_2483,N_2449);
nor U2588 (N_2588,N_2452,N_2407);
and U2589 (N_2589,N_2404,N_2492);
nand U2590 (N_2590,N_2407,N_2445);
nor U2591 (N_2591,N_2401,N_2438);
xor U2592 (N_2592,N_2424,N_2415);
nor U2593 (N_2593,N_2449,N_2435);
xor U2594 (N_2594,N_2421,N_2457);
xor U2595 (N_2595,N_2453,N_2409);
nand U2596 (N_2596,N_2412,N_2459);
nor U2597 (N_2597,N_2446,N_2484);
or U2598 (N_2598,N_2420,N_2464);
xor U2599 (N_2599,N_2489,N_2471);
and U2600 (N_2600,N_2588,N_2569);
or U2601 (N_2601,N_2525,N_2590);
xnor U2602 (N_2602,N_2543,N_2512);
or U2603 (N_2603,N_2599,N_2507);
nor U2604 (N_2604,N_2538,N_2578);
nand U2605 (N_2605,N_2583,N_2530);
and U2606 (N_2606,N_2584,N_2571);
nand U2607 (N_2607,N_2515,N_2595);
and U2608 (N_2608,N_2558,N_2541);
nand U2609 (N_2609,N_2573,N_2535);
xor U2610 (N_2610,N_2516,N_2524);
nand U2611 (N_2611,N_2559,N_2597);
nor U2612 (N_2612,N_2544,N_2561);
or U2613 (N_2613,N_2593,N_2529);
and U2614 (N_2614,N_2506,N_2522);
nand U2615 (N_2615,N_2557,N_2591);
nand U2616 (N_2616,N_2501,N_2511);
or U2617 (N_2617,N_2577,N_2553);
or U2618 (N_2618,N_2539,N_2596);
nand U2619 (N_2619,N_2519,N_2545);
or U2620 (N_2620,N_2502,N_2575);
nor U2621 (N_2621,N_2518,N_2509);
nor U2622 (N_2622,N_2552,N_2548);
xnor U2623 (N_2623,N_2536,N_2562);
nor U2624 (N_2624,N_2534,N_2560);
nand U2625 (N_2625,N_2505,N_2565);
nor U2626 (N_2626,N_2526,N_2550);
or U2627 (N_2627,N_2570,N_2514);
nand U2628 (N_2628,N_2532,N_2554);
nor U2629 (N_2629,N_2576,N_2542);
or U2630 (N_2630,N_2564,N_2586);
or U2631 (N_2631,N_2563,N_2547);
and U2632 (N_2632,N_2517,N_2582);
or U2633 (N_2633,N_2580,N_2567);
and U2634 (N_2634,N_2585,N_2533);
or U2635 (N_2635,N_2598,N_2546);
or U2636 (N_2636,N_2555,N_2504);
nand U2637 (N_2637,N_2592,N_2572);
xor U2638 (N_2638,N_2589,N_2574);
or U2639 (N_2639,N_2520,N_2566);
or U2640 (N_2640,N_2503,N_2556);
nor U2641 (N_2641,N_2540,N_2513);
and U2642 (N_2642,N_2581,N_2579);
xnor U2643 (N_2643,N_2587,N_2537);
nand U2644 (N_2644,N_2594,N_2527);
or U2645 (N_2645,N_2531,N_2528);
and U2646 (N_2646,N_2500,N_2508);
xnor U2647 (N_2647,N_2521,N_2551);
and U2648 (N_2648,N_2568,N_2523);
nand U2649 (N_2649,N_2510,N_2549);
and U2650 (N_2650,N_2505,N_2543);
nand U2651 (N_2651,N_2538,N_2537);
and U2652 (N_2652,N_2508,N_2561);
and U2653 (N_2653,N_2565,N_2572);
nand U2654 (N_2654,N_2568,N_2564);
and U2655 (N_2655,N_2533,N_2517);
and U2656 (N_2656,N_2575,N_2555);
xnor U2657 (N_2657,N_2514,N_2552);
nand U2658 (N_2658,N_2598,N_2515);
and U2659 (N_2659,N_2592,N_2511);
nor U2660 (N_2660,N_2550,N_2557);
nor U2661 (N_2661,N_2540,N_2592);
or U2662 (N_2662,N_2545,N_2584);
and U2663 (N_2663,N_2578,N_2592);
xnor U2664 (N_2664,N_2511,N_2517);
xnor U2665 (N_2665,N_2554,N_2566);
nor U2666 (N_2666,N_2581,N_2595);
nand U2667 (N_2667,N_2576,N_2545);
nand U2668 (N_2668,N_2522,N_2538);
and U2669 (N_2669,N_2534,N_2516);
or U2670 (N_2670,N_2579,N_2574);
nand U2671 (N_2671,N_2500,N_2586);
nand U2672 (N_2672,N_2533,N_2540);
nand U2673 (N_2673,N_2582,N_2531);
and U2674 (N_2674,N_2508,N_2595);
xor U2675 (N_2675,N_2599,N_2508);
xnor U2676 (N_2676,N_2559,N_2516);
and U2677 (N_2677,N_2503,N_2521);
xnor U2678 (N_2678,N_2592,N_2580);
nand U2679 (N_2679,N_2515,N_2549);
xor U2680 (N_2680,N_2583,N_2549);
xnor U2681 (N_2681,N_2542,N_2547);
nor U2682 (N_2682,N_2542,N_2578);
nor U2683 (N_2683,N_2551,N_2578);
xor U2684 (N_2684,N_2577,N_2599);
xnor U2685 (N_2685,N_2546,N_2531);
nand U2686 (N_2686,N_2562,N_2527);
and U2687 (N_2687,N_2597,N_2575);
nand U2688 (N_2688,N_2541,N_2553);
or U2689 (N_2689,N_2533,N_2546);
nor U2690 (N_2690,N_2545,N_2594);
or U2691 (N_2691,N_2540,N_2507);
or U2692 (N_2692,N_2528,N_2573);
xor U2693 (N_2693,N_2523,N_2583);
xor U2694 (N_2694,N_2569,N_2533);
nand U2695 (N_2695,N_2540,N_2501);
or U2696 (N_2696,N_2504,N_2571);
xnor U2697 (N_2697,N_2599,N_2598);
nand U2698 (N_2698,N_2592,N_2542);
or U2699 (N_2699,N_2523,N_2584);
nand U2700 (N_2700,N_2678,N_2633);
or U2701 (N_2701,N_2635,N_2643);
and U2702 (N_2702,N_2691,N_2613);
and U2703 (N_2703,N_2607,N_2649);
and U2704 (N_2704,N_2627,N_2606);
nand U2705 (N_2705,N_2614,N_2619);
or U2706 (N_2706,N_2674,N_2629);
and U2707 (N_2707,N_2602,N_2654);
or U2708 (N_2708,N_2632,N_2646);
and U2709 (N_2709,N_2604,N_2653);
or U2710 (N_2710,N_2612,N_2652);
nor U2711 (N_2711,N_2623,N_2601);
xnor U2712 (N_2712,N_2666,N_2609);
xor U2713 (N_2713,N_2689,N_2656);
or U2714 (N_2714,N_2676,N_2641);
nor U2715 (N_2715,N_2667,N_2610);
or U2716 (N_2716,N_2684,N_2668);
and U2717 (N_2717,N_2673,N_2622);
xor U2718 (N_2718,N_2662,N_2686);
and U2719 (N_2719,N_2682,N_2693);
and U2720 (N_2720,N_2650,N_2648);
nor U2721 (N_2721,N_2672,N_2608);
xnor U2722 (N_2722,N_2628,N_2651);
nor U2723 (N_2723,N_2642,N_2671);
nor U2724 (N_2724,N_2620,N_2639);
and U2725 (N_2725,N_2661,N_2657);
or U2726 (N_2726,N_2624,N_2687);
nor U2727 (N_2727,N_2695,N_2655);
or U2728 (N_2728,N_2680,N_2615);
nor U2729 (N_2729,N_2605,N_2663);
nand U2730 (N_2730,N_2621,N_2677);
xor U2731 (N_2731,N_2640,N_2630);
nand U2732 (N_2732,N_2698,N_2699);
or U2733 (N_2733,N_2616,N_2626);
nor U2734 (N_2734,N_2660,N_2681);
and U2735 (N_2735,N_2685,N_2690);
nand U2736 (N_2736,N_2617,N_2631);
and U2737 (N_2737,N_2637,N_2644);
nand U2738 (N_2738,N_2603,N_2669);
nand U2739 (N_2739,N_2625,N_2696);
xnor U2740 (N_2740,N_2675,N_2670);
xor U2741 (N_2741,N_2600,N_2688);
nor U2742 (N_2742,N_2697,N_2638);
xnor U2743 (N_2743,N_2611,N_2659);
xor U2744 (N_2744,N_2694,N_2647);
or U2745 (N_2745,N_2634,N_2679);
or U2746 (N_2746,N_2658,N_2664);
nor U2747 (N_2747,N_2618,N_2692);
or U2748 (N_2748,N_2665,N_2683);
and U2749 (N_2749,N_2645,N_2636);
nand U2750 (N_2750,N_2676,N_2691);
nor U2751 (N_2751,N_2677,N_2687);
and U2752 (N_2752,N_2657,N_2608);
nand U2753 (N_2753,N_2674,N_2606);
xor U2754 (N_2754,N_2615,N_2644);
nand U2755 (N_2755,N_2684,N_2623);
nand U2756 (N_2756,N_2677,N_2652);
and U2757 (N_2757,N_2618,N_2612);
and U2758 (N_2758,N_2614,N_2648);
or U2759 (N_2759,N_2695,N_2675);
nand U2760 (N_2760,N_2614,N_2608);
xnor U2761 (N_2761,N_2651,N_2679);
nand U2762 (N_2762,N_2648,N_2668);
nor U2763 (N_2763,N_2621,N_2635);
or U2764 (N_2764,N_2618,N_2654);
xor U2765 (N_2765,N_2648,N_2695);
xor U2766 (N_2766,N_2656,N_2692);
nand U2767 (N_2767,N_2616,N_2648);
xnor U2768 (N_2768,N_2645,N_2673);
and U2769 (N_2769,N_2669,N_2629);
or U2770 (N_2770,N_2616,N_2608);
nor U2771 (N_2771,N_2683,N_2655);
nand U2772 (N_2772,N_2605,N_2691);
nand U2773 (N_2773,N_2603,N_2656);
nand U2774 (N_2774,N_2642,N_2609);
nand U2775 (N_2775,N_2619,N_2663);
and U2776 (N_2776,N_2648,N_2634);
nor U2777 (N_2777,N_2640,N_2621);
and U2778 (N_2778,N_2694,N_2685);
nor U2779 (N_2779,N_2687,N_2632);
xor U2780 (N_2780,N_2612,N_2621);
and U2781 (N_2781,N_2650,N_2632);
or U2782 (N_2782,N_2661,N_2647);
nor U2783 (N_2783,N_2620,N_2667);
or U2784 (N_2784,N_2603,N_2666);
xor U2785 (N_2785,N_2670,N_2607);
nand U2786 (N_2786,N_2621,N_2659);
and U2787 (N_2787,N_2635,N_2628);
nor U2788 (N_2788,N_2687,N_2656);
or U2789 (N_2789,N_2675,N_2604);
xnor U2790 (N_2790,N_2656,N_2617);
and U2791 (N_2791,N_2655,N_2653);
nand U2792 (N_2792,N_2664,N_2609);
and U2793 (N_2793,N_2668,N_2692);
and U2794 (N_2794,N_2616,N_2658);
and U2795 (N_2795,N_2651,N_2695);
nor U2796 (N_2796,N_2667,N_2645);
and U2797 (N_2797,N_2640,N_2641);
nand U2798 (N_2798,N_2694,N_2690);
or U2799 (N_2799,N_2697,N_2620);
xnor U2800 (N_2800,N_2735,N_2701);
nand U2801 (N_2801,N_2785,N_2746);
nor U2802 (N_2802,N_2796,N_2736);
or U2803 (N_2803,N_2780,N_2763);
or U2804 (N_2804,N_2707,N_2700);
or U2805 (N_2805,N_2748,N_2712);
and U2806 (N_2806,N_2728,N_2792);
and U2807 (N_2807,N_2711,N_2708);
and U2808 (N_2808,N_2753,N_2777);
and U2809 (N_2809,N_2782,N_2751);
nand U2810 (N_2810,N_2724,N_2754);
or U2811 (N_2811,N_2742,N_2743);
xnor U2812 (N_2812,N_2765,N_2799);
and U2813 (N_2813,N_2755,N_2718);
nand U2814 (N_2814,N_2793,N_2715);
or U2815 (N_2815,N_2769,N_2733);
or U2816 (N_2816,N_2723,N_2730);
xor U2817 (N_2817,N_2786,N_2781);
nor U2818 (N_2818,N_2713,N_2745);
xnor U2819 (N_2819,N_2714,N_2761);
and U2820 (N_2820,N_2772,N_2775);
nand U2821 (N_2821,N_2767,N_2752);
and U2822 (N_2822,N_2791,N_2727);
or U2823 (N_2823,N_2757,N_2756);
or U2824 (N_2824,N_2726,N_2705);
xor U2825 (N_2825,N_2760,N_2768);
and U2826 (N_2826,N_2778,N_2709);
and U2827 (N_2827,N_2704,N_2773);
nand U2828 (N_2828,N_2740,N_2721);
nand U2829 (N_2829,N_2747,N_2774);
nor U2830 (N_2830,N_2766,N_2749);
nand U2831 (N_2831,N_2729,N_2784);
or U2832 (N_2832,N_2798,N_2750);
nor U2833 (N_2833,N_2722,N_2732);
and U2834 (N_2834,N_2764,N_2770);
nand U2835 (N_2835,N_2737,N_2789);
nor U2836 (N_2836,N_2719,N_2716);
xnor U2837 (N_2837,N_2783,N_2725);
and U2838 (N_2838,N_2706,N_2734);
or U2839 (N_2839,N_2790,N_2771);
nand U2840 (N_2840,N_2787,N_2720);
nor U2841 (N_2841,N_2738,N_2759);
xnor U2842 (N_2842,N_2703,N_2762);
and U2843 (N_2843,N_2739,N_2797);
and U2844 (N_2844,N_2776,N_2702);
xor U2845 (N_2845,N_2744,N_2731);
xor U2846 (N_2846,N_2788,N_2710);
and U2847 (N_2847,N_2779,N_2758);
or U2848 (N_2848,N_2741,N_2795);
nand U2849 (N_2849,N_2794,N_2717);
nor U2850 (N_2850,N_2704,N_2752);
nand U2851 (N_2851,N_2711,N_2742);
and U2852 (N_2852,N_2734,N_2720);
nand U2853 (N_2853,N_2760,N_2707);
xnor U2854 (N_2854,N_2702,N_2798);
nor U2855 (N_2855,N_2718,N_2757);
and U2856 (N_2856,N_2755,N_2798);
or U2857 (N_2857,N_2703,N_2787);
or U2858 (N_2858,N_2795,N_2737);
and U2859 (N_2859,N_2779,N_2750);
and U2860 (N_2860,N_2755,N_2757);
xor U2861 (N_2861,N_2715,N_2754);
nand U2862 (N_2862,N_2739,N_2718);
and U2863 (N_2863,N_2718,N_2780);
nor U2864 (N_2864,N_2712,N_2736);
or U2865 (N_2865,N_2748,N_2781);
and U2866 (N_2866,N_2750,N_2777);
or U2867 (N_2867,N_2718,N_2772);
nor U2868 (N_2868,N_2781,N_2737);
or U2869 (N_2869,N_2791,N_2790);
nor U2870 (N_2870,N_2760,N_2765);
nand U2871 (N_2871,N_2780,N_2700);
nor U2872 (N_2872,N_2738,N_2794);
nor U2873 (N_2873,N_2767,N_2798);
nand U2874 (N_2874,N_2744,N_2738);
and U2875 (N_2875,N_2707,N_2797);
or U2876 (N_2876,N_2788,N_2724);
xor U2877 (N_2877,N_2722,N_2709);
and U2878 (N_2878,N_2718,N_2778);
and U2879 (N_2879,N_2734,N_2783);
nand U2880 (N_2880,N_2750,N_2791);
nor U2881 (N_2881,N_2759,N_2782);
nand U2882 (N_2882,N_2778,N_2748);
or U2883 (N_2883,N_2773,N_2718);
and U2884 (N_2884,N_2726,N_2760);
xnor U2885 (N_2885,N_2747,N_2729);
nand U2886 (N_2886,N_2776,N_2745);
and U2887 (N_2887,N_2731,N_2751);
nand U2888 (N_2888,N_2725,N_2737);
or U2889 (N_2889,N_2704,N_2725);
xnor U2890 (N_2890,N_2772,N_2714);
or U2891 (N_2891,N_2702,N_2708);
nor U2892 (N_2892,N_2744,N_2754);
nand U2893 (N_2893,N_2779,N_2713);
nor U2894 (N_2894,N_2769,N_2770);
xnor U2895 (N_2895,N_2726,N_2770);
and U2896 (N_2896,N_2745,N_2746);
nand U2897 (N_2897,N_2760,N_2700);
nand U2898 (N_2898,N_2726,N_2758);
nand U2899 (N_2899,N_2788,N_2723);
or U2900 (N_2900,N_2805,N_2816);
and U2901 (N_2901,N_2869,N_2871);
xnor U2902 (N_2902,N_2860,N_2810);
or U2903 (N_2903,N_2861,N_2800);
xnor U2904 (N_2904,N_2811,N_2850);
nor U2905 (N_2905,N_2887,N_2826);
nor U2906 (N_2906,N_2866,N_2827);
nand U2907 (N_2907,N_2896,N_2819);
nand U2908 (N_2908,N_2815,N_2835);
xnor U2909 (N_2909,N_2879,N_2894);
or U2910 (N_2910,N_2818,N_2849);
xnor U2911 (N_2911,N_2838,N_2868);
or U2912 (N_2912,N_2832,N_2820);
xnor U2913 (N_2913,N_2885,N_2891);
nor U2914 (N_2914,N_2863,N_2803);
nor U2915 (N_2915,N_2813,N_2830);
or U2916 (N_2916,N_2802,N_2888);
nor U2917 (N_2917,N_2876,N_2856);
or U2918 (N_2918,N_2893,N_2828);
and U2919 (N_2919,N_2872,N_2884);
nand U2920 (N_2920,N_2857,N_2847);
xnor U2921 (N_2921,N_2889,N_2874);
nand U2922 (N_2922,N_2824,N_2855);
xnor U2923 (N_2923,N_2829,N_2806);
nor U2924 (N_2924,N_2833,N_2867);
nand U2925 (N_2925,N_2823,N_2808);
nand U2926 (N_2926,N_2862,N_2831);
nor U2927 (N_2927,N_2875,N_2834);
xnor U2928 (N_2928,N_2890,N_2812);
and U2929 (N_2929,N_2865,N_2883);
nor U2930 (N_2930,N_2804,N_2845);
and U2931 (N_2931,N_2895,N_2852);
nand U2932 (N_2932,N_2878,N_2899);
nand U2933 (N_2933,N_2807,N_2892);
or U2934 (N_2934,N_2848,N_2897);
nor U2935 (N_2935,N_2843,N_2822);
or U2936 (N_2936,N_2854,N_2809);
xor U2937 (N_2937,N_2870,N_2842);
or U2938 (N_2938,N_2821,N_2841);
xnor U2939 (N_2939,N_2858,N_2844);
or U2940 (N_2940,N_2836,N_2839);
or U2941 (N_2941,N_2801,N_2881);
nor U2942 (N_2942,N_2825,N_2882);
xor U2943 (N_2943,N_2817,N_2851);
nor U2944 (N_2944,N_2873,N_2837);
or U2945 (N_2945,N_2864,N_2898);
nor U2946 (N_2946,N_2877,N_2886);
xor U2947 (N_2947,N_2853,N_2814);
nor U2948 (N_2948,N_2840,N_2880);
nor U2949 (N_2949,N_2859,N_2846);
xnor U2950 (N_2950,N_2855,N_2886);
nor U2951 (N_2951,N_2888,N_2864);
or U2952 (N_2952,N_2875,N_2891);
or U2953 (N_2953,N_2894,N_2849);
xnor U2954 (N_2954,N_2836,N_2832);
and U2955 (N_2955,N_2858,N_2849);
or U2956 (N_2956,N_2859,N_2856);
or U2957 (N_2957,N_2885,N_2873);
xor U2958 (N_2958,N_2880,N_2861);
xor U2959 (N_2959,N_2835,N_2841);
and U2960 (N_2960,N_2897,N_2885);
xnor U2961 (N_2961,N_2882,N_2851);
and U2962 (N_2962,N_2820,N_2843);
and U2963 (N_2963,N_2891,N_2811);
nand U2964 (N_2964,N_2826,N_2827);
nor U2965 (N_2965,N_2851,N_2893);
and U2966 (N_2966,N_2812,N_2899);
or U2967 (N_2967,N_2831,N_2803);
and U2968 (N_2968,N_2890,N_2804);
or U2969 (N_2969,N_2804,N_2899);
or U2970 (N_2970,N_2872,N_2839);
xor U2971 (N_2971,N_2805,N_2896);
nor U2972 (N_2972,N_2856,N_2837);
xnor U2973 (N_2973,N_2840,N_2806);
nor U2974 (N_2974,N_2873,N_2822);
nand U2975 (N_2975,N_2829,N_2815);
and U2976 (N_2976,N_2876,N_2808);
and U2977 (N_2977,N_2856,N_2852);
and U2978 (N_2978,N_2895,N_2874);
xor U2979 (N_2979,N_2831,N_2835);
nand U2980 (N_2980,N_2825,N_2803);
and U2981 (N_2981,N_2802,N_2840);
nor U2982 (N_2982,N_2882,N_2823);
nand U2983 (N_2983,N_2893,N_2873);
or U2984 (N_2984,N_2864,N_2893);
nand U2985 (N_2985,N_2855,N_2881);
xnor U2986 (N_2986,N_2826,N_2853);
nor U2987 (N_2987,N_2824,N_2861);
and U2988 (N_2988,N_2824,N_2845);
nor U2989 (N_2989,N_2899,N_2817);
nor U2990 (N_2990,N_2836,N_2895);
xnor U2991 (N_2991,N_2875,N_2850);
or U2992 (N_2992,N_2818,N_2851);
and U2993 (N_2993,N_2821,N_2881);
xor U2994 (N_2994,N_2875,N_2857);
nor U2995 (N_2995,N_2856,N_2801);
nor U2996 (N_2996,N_2840,N_2876);
nand U2997 (N_2997,N_2802,N_2853);
nand U2998 (N_2998,N_2886,N_2830);
and U2999 (N_2999,N_2802,N_2839);
xor UO_0 (O_0,N_2918,N_2967);
or UO_1 (O_1,N_2907,N_2965);
xnor UO_2 (O_2,N_2929,N_2959);
nor UO_3 (O_3,N_2989,N_2933);
xnor UO_4 (O_4,N_2909,N_2958);
nand UO_5 (O_5,N_2936,N_2985);
and UO_6 (O_6,N_2906,N_2949);
nor UO_7 (O_7,N_2923,N_2986);
nand UO_8 (O_8,N_2908,N_2943);
xnor UO_9 (O_9,N_2988,N_2999);
nand UO_10 (O_10,N_2972,N_2990);
xor UO_11 (O_11,N_2917,N_2951);
xor UO_12 (O_12,N_2993,N_2978);
and UO_13 (O_13,N_2960,N_2901);
or UO_14 (O_14,N_2922,N_2927);
xnor UO_15 (O_15,N_2997,N_2920);
nand UO_16 (O_16,N_2942,N_2973);
and UO_17 (O_17,N_2961,N_2948);
xor UO_18 (O_18,N_2925,N_2905);
nand UO_19 (O_19,N_2915,N_2977);
or UO_20 (O_20,N_2913,N_2912);
nor UO_21 (O_21,N_2966,N_2992);
nor UO_22 (O_22,N_2926,N_2979);
or UO_23 (O_23,N_2974,N_2956);
nor UO_24 (O_24,N_2968,N_2995);
xnor UO_25 (O_25,N_2940,N_2964);
xnor UO_26 (O_26,N_2928,N_2980);
nand UO_27 (O_27,N_2945,N_2935);
xnor UO_28 (O_28,N_2938,N_2996);
or UO_29 (O_29,N_2975,N_2946);
xor UO_30 (O_30,N_2934,N_2924);
or UO_31 (O_31,N_2971,N_2987);
xor UO_32 (O_32,N_2937,N_2983);
nand UO_33 (O_33,N_2939,N_2963);
nor UO_34 (O_34,N_2904,N_2984);
xor UO_35 (O_35,N_2944,N_2981);
nand UO_36 (O_36,N_2919,N_2982);
xnor UO_37 (O_37,N_2952,N_2947);
xnor UO_38 (O_38,N_2903,N_2932);
xor UO_39 (O_39,N_2976,N_2953);
xor UO_40 (O_40,N_2914,N_2921);
nor UO_41 (O_41,N_2962,N_2910);
nor UO_42 (O_42,N_2930,N_2902);
or UO_43 (O_43,N_2950,N_2994);
and UO_44 (O_44,N_2991,N_2941);
nand UO_45 (O_45,N_2900,N_2970);
xor UO_46 (O_46,N_2955,N_2916);
nand UO_47 (O_47,N_2998,N_2957);
xnor UO_48 (O_48,N_2931,N_2954);
nand UO_49 (O_49,N_2969,N_2911);
or UO_50 (O_50,N_2953,N_2902);
nor UO_51 (O_51,N_2906,N_2978);
xnor UO_52 (O_52,N_2924,N_2965);
nor UO_53 (O_53,N_2958,N_2935);
xor UO_54 (O_54,N_2941,N_2936);
xor UO_55 (O_55,N_2918,N_2997);
or UO_56 (O_56,N_2931,N_2908);
nand UO_57 (O_57,N_2995,N_2905);
and UO_58 (O_58,N_2920,N_2948);
nor UO_59 (O_59,N_2945,N_2971);
xnor UO_60 (O_60,N_2900,N_2915);
nor UO_61 (O_61,N_2994,N_2928);
and UO_62 (O_62,N_2983,N_2969);
xnor UO_63 (O_63,N_2915,N_2961);
nand UO_64 (O_64,N_2908,N_2990);
or UO_65 (O_65,N_2933,N_2901);
nand UO_66 (O_66,N_2962,N_2913);
nand UO_67 (O_67,N_2983,N_2980);
and UO_68 (O_68,N_2914,N_2950);
and UO_69 (O_69,N_2975,N_2983);
xor UO_70 (O_70,N_2963,N_2919);
or UO_71 (O_71,N_2950,N_2900);
xnor UO_72 (O_72,N_2945,N_2927);
nor UO_73 (O_73,N_2932,N_2918);
nor UO_74 (O_74,N_2908,N_2909);
and UO_75 (O_75,N_2916,N_2986);
or UO_76 (O_76,N_2905,N_2989);
and UO_77 (O_77,N_2915,N_2950);
nand UO_78 (O_78,N_2998,N_2921);
and UO_79 (O_79,N_2965,N_2951);
xor UO_80 (O_80,N_2943,N_2947);
or UO_81 (O_81,N_2929,N_2982);
xor UO_82 (O_82,N_2994,N_2990);
xor UO_83 (O_83,N_2955,N_2909);
nand UO_84 (O_84,N_2900,N_2962);
nor UO_85 (O_85,N_2920,N_2951);
and UO_86 (O_86,N_2953,N_2979);
and UO_87 (O_87,N_2917,N_2967);
xor UO_88 (O_88,N_2914,N_2923);
xor UO_89 (O_89,N_2910,N_2922);
or UO_90 (O_90,N_2978,N_2938);
and UO_91 (O_91,N_2953,N_2920);
or UO_92 (O_92,N_2950,N_2960);
and UO_93 (O_93,N_2972,N_2995);
nor UO_94 (O_94,N_2942,N_2935);
or UO_95 (O_95,N_2911,N_2991);
and UO_96 (O_96,N_2972,N_2998);
xor UO_97 (O_97,N_2995,N_2991);
and UO_98 (O_98,N_2939,N_2920);
nor UO_99 (O_99,N_2968,N_2977);
nor UO_100 (O_100,N_2989,N_2943);
and UO_101 (O_101,N_2939,N_2966);
and UO_102 (O_102,N_2907,N_2942);
nand UO_103 (O_103,N_2956,N_2900);
and UO_104 (O_104,N_2979,N_2958);
xnor UO_105 (O_105,N_2914,N_2995);
or UO_106 (O_106,N_2972,N_2981);
nor UO_107 (O_107,N_2960,N_2924);
and UO_108 (O_108,N_2912,N_2921);
nand UO_109 (O_109,N_2987,N_2916);
nor UO_110 (O_110,N_2934,N_2919);
nor UO_111 (O_111,N_2915,N_2922);
nor UO_112 (O_112,N_2976,N_2928);
xor UO_113 (O_113,N_2999,N_2917);
nor UO_114 (O_114,N_2995,N_2906);
xnor UO_115 (O_115,N_2905,N_2911);
or UO_116 (O_116,N_2973,N_2991);
nor UO_117 (O_117,N_2981,N_2919);
nor UO_118 (O_118,N_2906,N_2926);
and UO_119 (O_119,N_2915,N_2935);
nor UO_120 (O_120,N_2978,N_2930);
nor UO_121 (O_121,N_2969,N_2902);
nand UO_122 (O_122,N_2948,N_2983);
nand UO_123 (O_123,N_2974,N_2946);
nor UO_124 (O_124,N_2914,N_2951);
nor UO_125 (O_125,N_2992,N_2938);
xnor UO_126 (O_126,N_2983,N_2924);
and UO_127 (O_127,N_2930,N_2995);
and UO_128 (O_128,N_2988,N_2972);
and UO_129 (O_129,N_2987,N_2955);
nand UO_130 (O_130,N_2999,N_2933);
or UO_131 (O_131,N_2955,N_2910);
and UO_132 (O_132,N_2939,N_2937);
xor UO_133 (O_133,N_2954,N_2907);
or UO_134 (O_134,N_2908,N_2919);
xnor UO_135 (O_135,N_2900,N_2941);
nor UO_136 (O_136,N_2900,N_2933);
and UO_137 (O_137,N_2911,N_2904);
nor UO_138 (O_138,N_2941,N_2930);
nor UO_139 (O_139,N_2979,N_2955);
xor UO_140 (O_140,N_2948,N_2903);
xor UO_141 (O_141,N_2987,N_2922);
or UO_142 (O_142,N_2932,N_2908);
nor UO_143 (O_143,N_2903,N_2956);
and UO_144 (O_144,N_2935,N_2961);
or UO_145 (O_145,N_2927,N_2957);
nor UO_146 (O_146,N_2974,N_2934);
xor UO_147 (O_147,N_2997,N_2954);
and UO_148 (O_148,N_2934,N_2985);
or UO_149 (O_149,N_2916,N_2975);
or UO_150 (O_150,N_2958,N_2905);
nand UO_151 (O_151,N_2985,N_2963);
and UO_152 (O_152,N_2992,N_2999);
nand UO_153 (O_153,N_2917,N_2974);
nor UO_154 (O_154,N_2980,N_2948);
nor UO_155 (O_155,N_2955,N_2990);
nand UO_156 (O_156,N_2960,N_2905);
nand UO_157 (O_157,N_2995,N_2983);
xor UO_158 (O_158,N_2912,N_2908);
or UO_159 (O_159,N_2923,N_2975);
nand UO_160 (O_160,N_2970,N_2948);
nor UO_161 (O_161,N_2964,N_2984);
or UO_162 (O_162,N_2999,N_2990);
nor UO_163 (O_163,N_2986,N_2930);
nand UO_164 (O_164,N_2932,N_2979);
nand UO_165 (O_165,N_2960,N_2943);
and UO_166 (O_166,N_2953,N_2916);
nor UO_167 (O_167,N_2901,N_2963);
xor UO_168 (O_168,N_2931,N_2968);
and UO_169 (O_169,N_2965,N_2968);
nand UO_170 (O_170,N_2905,N_2983);
or UO_171 (O_171,N_2975,N_2985);
nand UO_172 (O_172,N_2926,N_2958);
or UO_173 (O_173,N_2988,N_2953);
and UO_174 (O_174,N_2911,N_2933);
and UO_175 (O_175,N_2938,N_2972);
xnor UO_176 (O_176,N_2928,N_2953);
nor UO_177 (O_177,N_2919,N_2931);
xor UO_178 (O_178,N_2964,N_2921);
and UO_179 (O_179,N_2920,N_2921);
nor UO_180 (O_180,N_2952,N_2907);
and UO_181 (O_181,N_2945,N_2910);
or UO_182 (O_182,N_2981,N_2922);
or UO_183 (O_183,N_2946,N_2920);
nor UO_184 (O_184,N_2961,N_2973);
and UO_185 (O_185,N_2961,N_2989);
nor UO_186 (O_186,N_2971,N_2943);
nor UO_187 (O_187,N_2958,N_2914);
xor UO_188 (O_188,N_2953,N_2993);
and UO_189 (O_189,N_2984,N_2919);
nor UO_190 (O_190,N_2982,N_2958);
nor UO_191 (O_191,N_2957,N_2951);
nor UO_192 (O_192,N_2994,N_2966);
xnor UO_193 (O_193,N_2989,N_2974);
or UO_194 (O_194,N_2945,N_2979);
nor UO_195 (O_195,N_2943,N_2940);
and UO_196 (O_196,N_2900,N_2914);
and UO_197 (O_197,N_2994,N_2925);
or UO_198 (O_198,N_2974,N_2931);
nor UO_199 (O_199,N_2901,N_2967);
and UO_200 (O_200,N_2959,N_2994);
xor UO_201 (O_201,N_2950,N_2978);
nor UO_202 (O_202,N_2989,N_2959);
nor UO_203 (O_203,N_2965,N_2901);
xnor UO_204 (O_204,N_2942,N_2959);
nor UO_205 (O_205,N_2959,N_2919);
and UO_206 (O_206,N_2974,N_2979);
nor UO_207 (O_207,N_2917,N_2915);
and UO_208 (O_208,N_2966,N_2979);
xor UO_209 (O_209,N_2969,N_2907);
xor UO_210 (O_210,N_2967,N_2927);
xnor UO_211 (O_211,N_2972,N_2964);
xnor UO_212 (O_212,N_2989,N_2921);
nor UO_213 (O_213,N_2998,N_2999);
and UO_214 (O_214,N_2915,N_2993);
nand UO_215 (O_215,N_2956,N_2957);
nor UO_216 (O_216,N_2923,N_2922);
nor UO_217 (O_217,N_2920,N_2991);
or UO_218 (O_218,N_2900,N_2988);
nor UO_219 (O_219,N_2950,N_2971);
xor UO_220 (O_220,N_2964,N_2928);
xnor UO_221 (O_221,N_2918,N_2939);
nand UO_222 (O_222,N_2936,N_2922);
nand UO_223 (O_223,N_2907,N_2997);
xor UO_224 (O_224,N_2915,N_2920);
xor UO_225 (O_225,N_2955,N_2902);
or UO_226 (O_226,N_2937,N_2911);
and UO_227 (O_227,N_2949,N_2920);
xor UO_228 (O_228,N_2939,N_2926);
or UO_229 (O_229,N_2934,N_2956);
or UO_230 (O_230,N_2907,N_2906);
or UO_231 (O_231,N_2956,N_2951);
and UO_232 (O_232,N_2962,N_2902);
nand UO_233 (O_233,N_2953,N_2910);
nor UO_234 (O_234,N_2900,N_2964);
or UO_235 (O_235,N_2975,N_2962);
xnor UO_236 (O_236,N_2972,N_2916);
and UO_237 (O_237,N_2938,N_2995);
and UO_238 (O_238,N_2999,N_2985);
nor UO_239 (O_239,N_2902,N_2981);
and UO_240 (O_240,N_2930,N_2944);
or UO_241 (O_241,N_2972,N_2915);
and UO_242 (O_242,N_2927,N_2978);
nand UO_243 (O_243,N_2923,N_2900);
xor UO_244 (O_244,N_2974,N_2900);
or UO_245 (O_245,N_2956,N_2912);
nor UO_246 (O_246,N_2997,N_2998);
or UO_247 (O_247,N_2973,N_2978);
or UO_248 (O_248,N_2909,N_2915);
xor UO_249 (O_249,N_2923,N_2950);
or UO_250 (O_250,N_2945,N_2903);
xor UO_251 (O_251,N_2998,N_2906);
xor UO_252 (O_252,N_2954,N_2959);
and UO_253 (O_253,N_2996,N_2986);
nand UO_254 (O_254,N_2924,N_2948);
xnor UO_255 (O_255,N_2915,N_2971);
or UO_256 (O_256,N_2941,N_2907);
nand UO_257 (O_257,N_2973,N_2950);
nor UO_258 (O_258,N_2977,N_2919);
nand UO_259 (O_259,N_2997,N_2966);
nand UO_260 (O_260,N_2957,N_2979);
nor UO_261 (O_261,N_2936,N_2982);
and UO_262 (O_262,N_2913,N_2995);
nand UO_263 (O_263,N_2958,N_2940);
xor UO_264 (O_264,N_2965,N_2972);
or UO_265 (O_265,N_2911,N_2915);
and UO_266 (O_266,N_2971,N_2975);
nor UO_267 (O_267,N_2902,N_2947);
or UO_268 (O_268,N_2921,N_2910);
or UO_269 (O_269,N_2981,N_2905);
nor UO_270 (O_270,N_2922,N_2973);
xnor UO_271 (O_271,N_2944,N_2909);
nand UO_272 (O_272,N_2904,N_2991);
nor UO_273 (O_273,N_2904,N_2928);
nor UO_274 (O_274,N_2989,N_2924);
nand UO_275 (O_275,N_2959,N_2983);
and UO_276 (O_276,N_2993,N_2904);
nand UO_277 (O_277,N_2901,N_2907);
xor UO_278 (O_278,N_2936,N_2951);
nor UO_279 (O_279,N_2993,N_2948);
and UO_280 (O_280,N_2971,N_2994);
or UO_281 (O_281,N_2910,N_2949);
nand UO_282 (O_282,N_2983,N_2971);
nor UO_283 (O_283,N_2952,N_2992);
xnor UO_284 (O_284,N_2950,N_2972);
and UO_285 (O_285,N_2933,N_2936);
and UO_286 (O_286,N_2956,N_2975);
and UO_287 (O_287,N_2930,N_2957);
or UO_288 (O_288,N_2991,N_2992);
nand UO_289 (O_289,N_2926,N_2965);
nand UO_290 (O_290,N_2906,N_2920);
and UO_291 (O_291,N_2983,N_2964);
nand UO_292 (O_292,N_2951,N_2935);
and UO_293 (O_293,N_2982,N_2904);
nand UO_294 (O_294,N_2988,N_2903);
xnor UO_295 (O_295,N_2942,N_2948);
or UO_296 (O_296,N_2990,N_2938);
xor UO_297 (O_297,N_2901,N_2958);
nand UO_298 (O_298,N_2920,N_2912);
nor UO_299 (O_299,N_2939,N_2955);
nand UO_300 (O_300,N_2954,N_2922);
nand UO_301 (O_301,N_2934,N_2990);
or UO_302 (O_302,N_2964,N_2957);
nand UO_303 (O_303,N_2902,N_2954);
nand UO_304 (O_304,N_2903,N_2914);
and UO_305 (O_305,N_2942,N_2965);
nand UO_306 (O_306,N_2971,N_2932);
and UO_307 (O_307,N_2927,N_2991);
or UO_308 (O_308,N_2912,N_2939);
or UO_309 (O_309,N_2986,N_2945);
nand UO_310 (O_310,N_2915,N_2998);
xor UO_311 (O_311,N_2950,N_2935);
nor UO_312 (O_312,N_2909,N_2923);
nor UO_313 (O_313,N_2902,N_2985);
nor UO_314 (O_314,N_2956,N_2930);
and UO_315 (O_315,N_2975,N_2911);
xnor UO_316 (O_316,N_2932,N_2968);
nand UO_317 (O_317,N_2959,N_2916);
xor UO_318 (O_318,N_2980,N_2951);
and UO_319 (O_319,N_2972,N_2929);
and UO_320 (O_320,N_2928,N_2939);
or UO_321 (O_321,N_2984,N_2973);
xnor UO_322 (O_322,N_2967,N_2910);
nand UO_323 (O_323,N_2930,N_2905);
xnor UO_324 (O_324,N_2919,N_2917);
nor UO_325 (O_325,N_2975,N_2954);
xnor UO_326 (O_326,N_2932,N_2913);
nor UO_327 (O_327,N_2905,N_2979);
nor UO_328 (O_328,N_2920,N_2922);
and UO_329 (O_329,N_2927,N_2907);
nand UO_330 (O_330,N_2942,N_2958);
nand UO_331 (O_331,N_2964,N_2901);
or UO_332 (O_332,N_2946,N_2999);
xnor UO_333 (O_333,N_2988,N_2964);
or UO_334 (O_334,N_2991,N_2956);
or UO_335 (O_335,N_2974,N_2910);
xnor UO_336 (O_336,N_2990,N_2996);
xor UO_337 (O_337,N_2981,N_2978);
and UO_338 (O_338,N_2984,N_2900);
xnor UO_339 (O_339,N_2961,N_2977);
nor UO_340 (O_340,N_2912,N_2969);
and UO_341 (O_341,N_2939,N_2948);
nor UO_342 (O_342,N_2920,N_2919);
and UO_343 (O_343,N_2956,N_2961);
nor UO_344 (O_344,N_2914,N_2997);
or UO_345 (O_345,N_2978,N_2921);
and UO_346 (O_346,N_2928,N_2973);
or UO_347 (O_347,N_2995,N_2920);
nand UO_348 (O_348,N_2967,N_2948);
or UO_349 (O_349,N_2978,N_2963);
xnor UO_350 (O_350,N_2921,N_2900);
xor UO_351 (O_351,N_2973,N_2983);
xor UO_352 (O_352,N_2939,N_2967);
or UO_353 (O_353,N_2937,N_2962);
nor UO_354 (O_354,N_2928,N_2998);
nand UO_355 (O_355,N_2943,N_2935);
nand UO_356 (O_356,N_2909,N_2943);
nor UO_357 (O_357,N_2972,N_2953);
xnor UO_358 (O_358,N_2919,N_2928);
nand UO_359 (O_359,N_2933,N_2913);
or UO_360 (O_360,N_2909,N_2954);
and UO_361 (O_361,N_2908,N_2958);
nand UO_362 (O_362,N_2905,N_2935);
nor UO_363 (O_363,N_2950,N_2931);
or UO_364 (O_364,N_2995,N_2928);
nor UO_365 (O_365,N_2952,N_2964);
nand UO_366 (O_366,N_2925,N_2902);
nor UO_367 (O_367,N_2906,N_2933);
nor UO_368 (O_368,N_2948,N_2916);
nand UO_369 (O_369,N_2921,N_2918);
or UO_370 (O_370,N_2989,N_2983);
and UO_371 (O_371,N_2998,N_2973);
and UO_372 (O_372,N_2985,N_2971);
and UO_373 (O_373,N_2925,N_2933);
and UO_374 (O_374,N_2912,N_2971);
nor UO_375 (O_375,N_2923,N_2995);
nand UO_376 (O_376,N_2932,N_2995);
nand UO_377 (O_377,N_2937,N_2910);
xnor UO_378 (O_378,N_2955,N_2986);
nand UO_379 (O_379,N_2982,N_2996);
and UO_380 (O_380,N_2967,N_2906);
xnor UO_381 (O_381,N_2998,N_2966);
nand UO_382 (O_382,N_2927,N_2963);
nor UO_383 (O_383,N_2943,N_2937);
or UO_384 (O_384,N_2986,N_2989);
xnor UO_385 (O_385,N_2956,N_2942);
nand UO_386 (O_386,N_2903,N_2951);
nand UO_387 (O_387,N_2965,N_2967);
nor UO_388 (O_388,N_2951,N_2938);
and UO_389 (O_389,N_2958,N_2934);
xor UO_390 (O_390,N_2905,N_2961);
or UO_391 (O_391,N_2923,N_2905);
and UO_392 (O_392,N_2948,N_2943);
and UO_393 (O_393,N_2944,N_2983);
and UO_394 (O_394,N_2917,N_2960);
nand UO_395 (O_395,N_2935,N_2955);
nor UO_396 (O_396,N_2920,N_2913);
nand UO_397 (O_397,N_2911,N_2951);
and UO_398 (O_398,N_2984,N_2972);
xnor UO_399 (O_399,N_2900,N_2954);
xor UO_400 (O_400,N_2921,N_2911);
or UO_401 (O_401,N_2929,N_2907);
xor UO_402 (O_402,N_2952,N_2982);
and UO_403 (O_403,N_2941,N_2982);
xnor UO_404 (O_404,N_2990,N_2919);
nand UO_405 (O_405,N_2956,N_2981);
or UO_406 (O_406,N_2945,N_2914);
nand UO_407 (O_407,N_2944,N_2993);
and UO_408 (O_408,N_2927,N_2988);
nor UO_409 (O_409,N_2990,N_2948);
nor UO_410 (O_410,N_2960,N_2915);
nor UO_411 (O_411,N_2939,N_2964);
nand UO_412 (O_412,N_2937,N_2970);
or UO_413 (O_413,N_2908,N_2978);
and UO_414 (O_414,N_2963,N_2970);
or UO_415 (O_415,N_2922,N_2921);
xor UO_416 (O_416,N_2979,N_2921);
or UO_417 (O_417,N_2995,N_2962);
nand UO_418 (O_418,N_2971,N_2934);
nand UO_419 (O_419,N_2973,N_2946);
nor UO_420 (O_420,N_2928,N_2971);
xnor UO_421 (O_421,N_2922,N_2911);
nor UO_422 (O_422,N_2998,N_2900);
xnor UO_423 (O_423,N_2953,N_2913);
nor UO_424 (O_424,N_2962,N_2917);
or UO_425 (O_425,N_2953,N_2986);
xnor UO_426 (O_426,N_2998,N_2916);
and UO_427 (O_427,N_2943,N_2969);
and UO_428 (O_428,N_2990,N_2947);
nor UO_429 (O_429,N_2981,N_2982);
or UO_430 (O_430,N_2926,N_2923);
xnor UO_431 (O_431,N_2964,N_2985);
and UO_432 (O_432,N_2984,N_2913);
xnor UO_433 (O_433,N_2968,N_2980);
nor UO_434 (O_434,N_2980,N_2989);
or UO_435 (O_435,N_2981,N_2941);
and UO_436 (O_436,N_2981,N_2970);
and UO_437 (O_437,N_2980,N_2939);
nand UO_438 (O_438,N_2982,N_2987);
nand UO_439 (O_439,N_2970,N_2996);
nand UO_440 (O_440,N_2955,N_2901);
nand UO_441 (O_441,N_2958,N_2951);
nor UO_442 (O_442,N_2932,N_2943);
or UO_443 (O_443,N_2950,N_2903);
xor UO_444 (O_444,N_2973,N_2974);
nor UO_445 (O_445,N_2949,N_2934);
nand UO_446 (O_446,N_2942,N_2954);
xor UO_447 (O_447,N_2985,N_2979);
xnor UO_448 (O_448,N_2904,N_2986);
or UO_449 (O_449,N_2958,N_2981);
or UO_450 (O_450,N_2966,N_2905);
or UO_451 (O_451,N_2994,N_2900);
or UO_452 (O_452,N_2990,N_2944);
and UO_453 (O_453,N_2987,N_2960);
xor UO_454 (O_454,N_2961,N_2934);
nor UO_455 (O_455,N_2974,N_2918);
xnor UO_456 (O_456,N_2966,N_2982);
and UO_457 (O_457,N_2980,N_2902);
or UO_458 (O_458,N_2919,N_2968);
nor UO_459 (O_459,N_2960,N_2906);
nor UO_460 (O_460,N_2947,N_2939);
or UO_461 (O_461,N_2918,N_2962);
xor UO_462 (O_462,N_2909,N_2910);
nor UO_463 (O_463,N_2919,N_2983);
or UO_464 (O_464,N_2913,N_2973);
nand UO_465 (O_465,N_2927,N_2955);
xnor UO_466 (O_466,N_2967,N_2914);
or UO_467 (O_467,N_2921,N_2905);
nand UO_468 (O_468,N_2976,N_2960);
and UO_469 (O_469,N_2968,N_2940);
nor UO_470 (O_470,N_2969,N_2968);
nand UO_471 (O_471,N_2963,N_2956);
nor UO_472 (O_472,N_2997,N_2904);
xnor UO_473 (O_473,N_2909,N_2978);
xnor UO_474 (O_474,N_2944,N_2912);
xnor UO_475 (O_475,N_2991,N_2917);
and UO_476 (O_476,N_2916,N_2989);
nor UO_477 (O_477,N_2920,N_2987);
nand UO_478 (O_478,N_2931,N_2947);
or UO_479 (O_479,N_2924,N_2970);
and UO_480 (O_480,N_2995,N_2970);
nand UO_481 (O_481,N_2983,N_2955);
nor UO_482 (O_482,N_2971,N_2947);
xor UO_483 (O_483,N_2989,N_2939);
nor UO_484 (O_484,N_2902,N_2900);
and UO_485 (O_485,N_2975,N_2990);
and UO_486 (O_486,N_2940,N_2996);
and UO_487 (O_487,N_2904,N_2973);
xnor UO_488 (O_488,N_2972,N_2935);
nor UO_489 (O_489,N_2916,N_2964);
and UO_490 (O_490,N_2936,N_2906);
nand UO_491 (O_491,N_2909,N_2969);
xnor UO_492 (O_492,N_2982,N_2974);
or UO_493 (O_493,N_2938,N_2994);
and UO_494 (O_494,N_2942,N_2915);
or UO_495 (O_495,N_2927,N_2948);
nor UO_496 (O_496,N_2919,N_2955);
nand UO_497 (O_497,N_2972,N_2900);
nand UO_498 (O_498,N_2963,N_2940);
nor UO_499 (O_499,N_2937,N_2975);
endmodule