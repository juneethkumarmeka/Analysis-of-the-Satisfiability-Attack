module basic_1500_15000_2000_30_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_1145,In_1344);
xor U1 (N_1,In_1102,In_1143);
and U2 (N_2,In_527,In_805);
nand U3 (N_3,In_120,In_105);
nand U4 (N_4,In_522,In_777);
xnor U5 (N_5,In_623,In_530);
nand U6 (N_6,In_406,In_679);
xnor U7 (N_7,In_664,In_1123);
nand U8 (N_8,In_1313,In_218);
and U9 (N_9,In_754,In_303);
xor U10 (N_10,In_1134,In_423);
and U11 (N_11,In_1309,In_1182);
or U12 (N_12,In_966,In_609);
or U13 (N_13,In_119,In_1129);
or U14 (N_14,In_541,In_187);
nor U15 (N_15,In_1291,In_801);
xor U16 (N_16,In_781,In_1142);
or U17 (N_17,In_1370,In_546);
xnor U18 (N_18,In_952,In_352);
or U19 (N_19,In_1114,In_419);
and U20 (N_20,In_561,In_425);
nand U21 (N_21,In_770,In_1277);
nand U22 (N_22,In_824,In_574);
or U23 (N_23,In_377,In_1491);
or U24 (N_24,In_186,In_111);
nor U25 (N_25,In_453,In_929);
xnor U26 (N_26,In_1168,In_812);
and U27 (N_27,In_1483,In_946);
nand U28 (N_28,In_1385,In_851);
or U29 (N_29,In_1167,In_697);
nand U30 (N_30,In_641,In_759);
nand U31 (N_31,In_1495,In_1332);
nand U32 (N_32,In_39,In_195);
or U33 (N_33,In_1327,In_748);
nand U34 (N_34,In_1031,In_470);
nand U35 (N_35,In_1466,In_289);
or U36 (N_36,In_294,In_213);
and U37 (N_37,In_1257,In_736);
or U38 (N_38,In_1490,In_1116);
and U39 (N_39,In_788,In_965);
nor U40 (N_40,In_655,In_771);
or U41 (N_41,In_354,In_569);
xnor U42 (N_42,In_1158,In_1341);
nand U43 (N_43,In_199,In_324);
nor U44 (N_44,In_710,In_1177);
nor U45 (N_45,In_1052,In_1380);
xnor U46 (N_46,In_415,In_5);
nor U47 (N_47,In_341,In_158);
or U48 (N_48,In_1359,In_1228);
nor U49 (N_49,In_258,In_50);
xor U50 (N_50,In_309,In_490);
and U51 (N_51,In_1269,In_862);
nand U52 (N_52,In_844,In_588);
or U53 (N_53,In_392,In_978);
nand U54 (N_54,In_480,In_1169);
nand U55 (N_55,In_662,In_1410);
nor U56 (N_56,In_845,In_765);
and U57 (N_57,In_1418,In_822);
or U58 (N_58,In_462,In_939);
nor U59 (N_59,In_133,In_1379);
xor U60 (N_60,In_672,In_854);
nand U61 (N_61,In_885,In_682);
or U62 (N_62,In_1343,In_1094);
xor U63 (N_63,In_72,In_810);
or U64 (N_64,In_432,In_927);
xor U65 (N_65,In_414,In_985);
and U66 (N_66,In_126,In_1106);
and U67 (N_67,In_300,In_1265);
nor U68 (N_68,In_257,In_1101);
nand U69 (N_69,In_1084,In_439);
and U70 (N_70,In_994,In_1172);
nand U71 (N_71,In_364,In_1024);
nand U72 (N_72,In_412,In_1246);
nor U73 (N_73,In_1464,In_458);
or U74 (N_74,In_88,In_728);
and U75 (N_75,In_1039,In_548);
or U76 (N_76,In_864,In_1331);
xor U77 (N_77,In_161,In_1258);
and U78 (N_78,In_92,In_660);
or U79 (N_79,In_367,In_15);
xnor U80 (N_80,In_476,In_832);
and U81 (N_81,In_1053,In_1063);
nor U82 (N_82,In_1465,In_1115);
xor U83 (N_83,In_659,In_694);
or U84 (N_84,In_519,In_135);
and U85 (N_85,In_1361,In_763);
or U86 (N_86,In_922,In_90);
nor U87 (N_87,In_865,In_206);
xor U88 (N_88,In_1047,In_553);
or U89 (N_89,In_245,In_311);
nand U90 (N_90,In_505,In_1077);
xnor U91 (N_91,In_350,In_1099);
nand U92 (N_92,In_1022,In_857);
nor U93 (N_93,In_1455,In_137);
or U94 (N_94,In_440,In_738);
and U95 (N_95,In_849,In_18);
nor U96 (N_96,In_1109,In_1147);
nand U97 (N_97,In_247,In_969);
or U98 (N_98,In_221,In_315);
or U99 (N_99,In_1056,In_43);
nor U100 (N_100,In_286,In_1006);
or U101 (N_101,In_614,In_704);
nor U102 (N_102,In_6,In_884);
nor U103 (N_103,In_680,In_340);
nand U104 (N_104,In_436,In_1090);
nand U105 (N_105,In_686,In_1171);
nor U106 (N_106,In_1184,In_1441);
and U107 (N_107,In_1071,In_1403);
xor U108 (N_108,In_368,In_796);
and U109 (N_109,In_1286,In_834);
nor U110 (N_110,In_671,In_915);
nor U111 (N_111,In_390,In_979);
nor U112 (N_112,In_718,In_878);
xnor U113 (N_113,In_1124,In_1021);
and U114 (N_114,In_938,In_1104);
nor U115 (N_115,In_1082,In_1268);
xor U116 (N_116,In_610,In_1356);
xor U117 (N_117,In_1007,In_1390);
and U118 (N_118,In_1191,In_262);
xor U119 (N_119,In_1315,In_1218);
and U120 (N_120,In_1243,In_651);
nand U121 (N_121,In_1453,In_427);
nand U122 (N_122,In_1272,In_1004);
nand U123 (N_123,In_215,In_358);
nand U124 (N_124,In_1451,In_403);
nand U125 (N_125,In_521,In_1381);
or U126 (N_126,In_977,In_1200);
or U127 (N_127,In_338,In_953);
nand U128 (N_128,In_1314,In_47);
nor U129 (N_129,In_1040,In_1292);
xor U130 (N_130,In_1149,In_1374);
xnor U131 (N_131,In_1264,In_850);
or U132 (N_132,In_1416,In_1035);
or U133 (N_133,In_725,In_1103);
or U134 (N_134,In_1162,In_933);
nand U135 (N_135,In_1027,In_1155);
and U136 (N_136,In_515,In_1450);
nand U137 (N_137,In_1442,In_1221);
nor U138 (N_138,In_1012,In_30);
or U139 (N_139,In_958,In_1316);
nand U140 (N_140,In_1079,In_855);
nand U141 (N_141,In_1303,In_1475);
xor U142 (N_142,In_1059,In_192);
or U143 (N_143,In_1023,In_317);
nor U144 (N_144,In_398,In_500);
or U145 (N_145,In_35,In_880);
and U146 (N_146,In_1426,In_1175);
nor U147 (N_147,In_41,In_32);
xnor U148 (N_148,In_563,In_619);
nand U149 (N_149,In_733,In_1428);
nor U150 (N_150,In_1308,In_94);
and U151 (N_151,In_1088,In_457);
xor U152 (N_152,In_1157,In_1457);
and U153 (N_153,In_1215,In_987);
nand U154 (N_154,In_591,In_255);
or U155 (N_155,In_495,In_203);
and U156 (N_156,In_1174,In_921);
xnor U157 (N_157,In_802,In_407);
or U158 (N_158,In_1140,In_113);
or U159 (N_159,In_379,In_260);
xor U160 (N_160,In_73,In_1135);
nand U161 (N_161,In_290,In_720);
nand U162 (N_162,In_983,In_210);
or U163 (N_163,In_944,In_231);
xor U164 (N_164,In_24,In_65);
xor U165 (N_165,In_321,In_346);
or U166 (N_166,In_611,In_901);
and U167 (N_167,In_755,In_523);
nand U168 (N_168,In_487,In_445);
nor U169 (N_169,In_863,In_1377);
nor U170 (N_170,In_673,In_1033);
xnor U171 (N_171,In_876,In_469);
or U172 (N_172,In_361,In_1444);
xnor U173 (N_173,In_1118,In_1041);
nand U174 (N_174,In_121,In_420);
xnor U175 (N_175,In_1132,In_70);
xnor U176 (N_176,In_1346,In_1497);
or U177 (N_177,In_993,In_26);
or U178 (N_178,In_587,In_1152);
or U179 (N_179,In_141,In_1064);
nor U180 (N_180,In_1312,In_10);
nor U181 (N_181,In_984,In_1224);
xor U182 (N_182,In_334,In_903);
xor U183 (N_183,In_417,In_230);
xnor U184 (N_184,In_1222,In_709);
and U185 (N_185,In_1065,In_1253);
nor U186 (N_186,In_1329,In_298);
nand U187 (N_187,In_526,In_1306);
nand U188 (N_188,In_349,In_20);
nand U189 (N_189,In_1443,In_394);
xor U190 (N_190,In_53,In_1122);
nor U191 (N_191,In_622,In_621);
nor U192 (N_192,In_1409,In_1494);
and U193 (N_193,In_1487,In_665);
and U194 (N_194,In_897,In_1280);
or U195 (N_195,In_595,In_846);
nand U196 (N_196,In_1354,In_1423);
and U197 (N_197,In_524,In_44);
or U198 (N_198,In_960,In_224);
xnor U199 (N_199,In_389,In_1340);
or U200 (N_200,In_163,In_740);
and U201 (N_201,In_716,In_1266);
and U202 (N_202,In_123,In_1010);
nor U203 (N_203,In_766,In_1216);
nor U204 (N_204,In_205,In_348);
xnor U205 (N_205,In_911,In_1438);
nor U206 (N_206,In_25,In_1139);
nand U207 (N_207,In_1477,In_776);
nor U208 (N_208,In_815,In_356);
nor U209 (N_209,In_607,In_745);
nand U210 (N_210,In_799,In_1435);
nor U211 (N_211,In_1239,In_148);
nand U212 (N_212,In_992,In_906);
and U213 (N_213,In_1117,In_155);
nor U214 (N_214,In_833,In_568);
nand U215 (N_215,In_613,In_792);
or U216 (N_216,In_1345,In_954);
nand U217 (N_217,In_376,In_554);
xor U218 (N_218,In_525,In_1427);
xnor U219 (N_219,In_632,In_695);
xnor U220 (N_220,In_491,In_594);
nand U221 (N_221,In_1138,In_23);
nand U222 (N_222,In_1097,In_283);
and U223 (N_223,In_624,In_475);
and U224 (N_224,In_769,In_1371);
xor U225 (N_225,In_643,In_580);
nand U226 (N_226,In_93,In_373);
nand U227 (N_227,In_516,In_1069);
nand U228 (N_228,In_1046,In_13);
and U229 (N_229,In_840,In_1034);
xor U230 (N_230,In_234,In_1202);
nand U231 (N_231,In_1323,In_971);
nor U232 (N_232,In_782,In_464);
nor U233 (N_233,In_896,In_1108);
nand U234 (N_234,In_547,In_504);
xor U235 (N_235,In_497,In_1412);
or U236 (N_236,In_1180,In_1016);
or U237 (N_237,In_335,In_78);
or U238 (N_238,In_49,In_482);
nand U239 (N_239,In_721,In_565);
nor U240 (N_240,In_1449,In_1217);
nor U241 (N_241,In_1382,In_705);
nor U242 (N_242,In_421,In_81);
nand U243 (N_243,In_450,In_1391);
or U244 (N_244,In_937,In_1296);
xor U245 (N_245,In_402,In_1244);
nor U246 (N_246,In_208,In_731);
and U247 (N_247,In_1384,In_973);
nor U248 (N_248,In_1092,In_177);
or U249 (N_249,In_1358,In_385);
xnor U250 (N_250,In_1349,In_166);
and U251 (N_251,In_919,In_575);
nor U252 (N_252,In_232,In_1375);
or U253 (N_253,In_638,In_1209);
nor U254 (N_254,In_129,In_501);
and U255 (N_255,In_484,In_685);
nor U256 (N_256,In_1458,In_396);
nand U257 (N_257,In_688,In_900);
xor U258 (N_258,In_435,In_219);
or U259 (N_259,In_512,In_917);
and U260 (N_260,In_1478,In_1001);
and U261 (N_261,In_1283,In_1201);
and U262 (N_262,In_332,In_820);
nand U263 (N_263,In_275,In_729);
nor U264 (N_264,In_183,In_1096);
and U265 (N_265,In_388,In_585);
and U266 (N_266,In_1055,In_761);
nand U267 (N_267,In_1445,In_270);
or U268 (N_268,In_925,In_606);
or U269 (N_269,In_821,In_690);
nor U270 (N_270,In_151,In_489);
nand U271 (N_271,In_399,In_1119);
or U272 (N_272,In_1018,In_276);
nor U273 (N_273,In_708,In_160);
nand U274 (N_274,In_428,In_1163);
or U275 (N_275,In_1098,In_56);
and U276 (N_276,In_1337,In_60);
nor U277 (N_277,In_456,In_254);
or U278 (N_278,In_323,In_14);
nand U279 (N_279,In_211,In_1400);
nand U280 (N_280,In_1013,In_127);
xnor U281 (N_281,In_45,In_1334);
xnor U282 (N_282,In_297,In_853);
nor U283 (N_283,In_961,In_657);
xor U284 (N_284,In_887,In_1235);
and U285 (N_285,In_413,In_401);
and U286 (N_286,In_1061,In_1166);
xnor U287 (N_287,In_1067,In_1270);
or U288 (N_288,In_583,In_787);
nor U289 (N_289,In_366,In_893);
nand U290 (N_290,In_79,In_905);
nor U291 (N_291,In_683,In_17);
nor U292 (N_292,In_443,In_764);
nand U293 (N_293,In_178,In_700);
nand U294 (N_294,In_827,In_263);
nand U295 (N_295,In_875,In_687);
nor U296 (N_296,In_916,In_1281);
nor U297 (N_297,In_89,In_1432);
or U298 (N_298,In_1000,In_804);
or U299 (N_299,In_605,In_438);
xnor U300 (N_300,In_261,In_1476);
nand U301 (N_301,In_836,In_950);
or U302 (N_302,In_68,In_835);
and U303 (N_303,In_362,In_951);
xor U304 (N_304,In_184,In_1127);
and U305 (N_305,In_1367,In_104);
or U306 (N_306,In_1363,In_816);
xnor U307 (N_307,In_779,In_1017);
nor U308 (N_308,In_517,In_191);
nand U309 (N_309,In_1299,In_238);
xor U310 (N_310,In_1369,In_1424);
nor U311 (N_311,In_593,In_1480);
nand U312 (N_312,In_1288,In_1319);
and U313 (N_313,In_1373,In_76);
and U314 (N_314,In_1398,In_1223);
and U315 (N_315,In_188,In_122);
and U316 (N_316,In_989,In_843);
or U317 (N_317,In_828,In_912);
and U318 (N_318,In_355,In_1226);
nand U319 (N_319,In_1130,In_762);
and U320 (N_320,In_3,In_856);
xor U321 (N_321,In_1318,In_964);
nor U322 (N_322,In_696,In_0);
xnor U323 (N_323,In_278,In_861);
nor U324 (N_324,In_460,In_91);
or U325 (N_325,In_1112,In_879);
xor U326 (N_326,In_1470,In_768);
or U327 (N_327,In_928,In_233);
xor U328 (N_328,In_1100,In_1275);
or U329 (N_329,In_870,In_1333);
and U330 (N_330,In_1060,In_604);
nand U331 (N_331,In_1456,In_408);
nand U332 (N_332,In_150,In_1095);
and U333 (N_333,In_790,In_1469);
or U334 (N_334,In_371,In_1324);
nor U335 (N_335,In_957,In_1290);
and U336 (N_336,In_1259,In_136);
nor U337 (N_337,In_29,In_1005);
nand U338 (N_338,In_1049,In_251);
nor U339 (N_339,In_970,In_75);
or U340 (N_340,In_1394,In_1326);
nand U341 (N_341,In_819,In_1192);
nand U342 (N_342,In_1240,In_1274);
nand U343 (N_343,In_717,In_1242);
or U344 (N_344,In_506,In_1499);
or U345 (N_345,In_532,In_806);
or U346 (N_346,In_249,In_743);
and U347 (N_347,In_99,In_847);
nor U348 (N_348,In_859,In_62);
or U349 (N_349,In_167,In_545);
nand U350 (N_350,In_502,In_59);
nor U351 (N_351,In_1225,In_981);
and U352 (N_352,In_508,In_1234);
and U353 (N_353,In_393,In_175);
xor U354 (N_354,In_132,In_883);
and U355 (N_355,In_531,In_692);
nor U356 (N_356,In_1074,In_473);
or U357 (N_357,In_809,In_567);
nor U358 (N_358,In_36,In_596);
nor U359 (N_359,In_1008,In_1219);
xnor U360 (N_360,In_1048,In_271);
nor U361 (N_361,In_1252,In_942);
and U362 (N_362,In_115,In_774);
nor U363 (N_363,In_1322,In_1485);
and U364 (N_364,In_868,In_1420);
or U365 (N_365,In_539,In_202);
or U366 (N_366,In_185,In_543);
xnor U367 (N_367,In_27,In_146);
nor U368 (N_368,In_1043,In_180);
and U369 (N_369,In_154,In_773);
or U370 (N_370,In_689,In_681);
and U371 (N_371,In_2,In_372);
xnor U372 (N_372,In_626,In_1030);
or U373 (N_373,In_772,In_182);
or U374 (N_374,In_444,In_174);
xnor U375 (N_375,In_1325,In_313);
nand U376 (N_376,In_649,In_1164);
xor U377 (N_377,In_287,In_240);
or U378 (N_378,In_194,In_1251);
nor U379 (N_379,In_1307,In_316);
xnor U380 (N_380,In_1126,In_477);
or U381 (N_381,In_320,In_107);
xnor U382 (N_382,In_314,In_248);
xnor U383 (N_383,In_1452,In_959);
xor U384 (N_384,In_503,In_1440);
nor U385 (N_385,In_38,In_882);
nor U386 (N_386,In_895,In_1111);
nand U387 (N_387,In_330,In_881);
or U388 (N_388,In_1404,In_980);
nand U389 (N_389,In_441,In_1353);
nand U390 (N_390,In_667,In_1462);
xnor U391 (N_391,In_227,In_637);
and U392 (N_392,In_1467,In_1393);
or U393 (N_393,In_923,In_1206);
nor U394 (N_394,In_706,In_1422);
or U395 (N_395,In_974,In_732);
and U396 (N_396,In_431,In_1078);
xnor U397 (N_397,In_307,In_359);
or U398 (N_398,In_829,In_1198);
and U399 (N_399,In_701,In_212);
nand U400 (N_400,In_597,In_1486);
or U401 (N_401,In_116,In_1236);
nand U402 (N_402,In_711,In_1289);
or U403 (N_403,In_351,In_1355);
and U404 (N_404,In_1014,In_246);
nand U405 (N_405,In_997,In_1137);
nand U406 (N_406,In_325,In_1399);
nand U407 (N_407,In_647,In_479);
or U408 (N_408,In_1179,In_823);
nor U409 (N_409,In_381,In_1057);
and U410 (N_410,In_1042,In_807);
xnor U411 (N_411,In_226,In_1062);
nor U412 (N_412,In_898,In_193);
nor U413 (N_413,In_308,In_21);
and U414 (N_414,In_635,In_747);
nor U415 (N_415,In_866,In_474);
nand U416 (N_416,In_319,In_1366);
nand U417 (N_417,In_726,In_889);
or U418 (N_418,In_838,In_1392);
nand U419 (N_419,In_114,In_301);
xnor U420 (N_420,In_932,In_1365);
or U421 (N_421,In_1153,In_1185);
and U422 (N_422,In_1304,In_934);
and U423 (N_423,In_1019,In_537);
or U424 (N_424,In_744,In_1181);
or U425 (N_425,In_108,In_1189);
and U426 (N_426,In_784,In_1075);
or U427 (N_427,In_1190,In_285);
and U428 (N_428,In_1335,In_165);
nand U429 (N_429,In_273,In_1386);
and U430 (N_430,In_723,In_197);
xor U431 (N_431,In_869,In_1425);
and U432 (N_432,In_1489,In_1248);
and U433 (N_433,In_1279,In_945);
and U434 (N_434,In_592,In_292);
or U435 (N_435,In_644,In_1496);
or U436 (N_436,In_1026,In_775);
nor U437 (N_437,In_280,In_256);
or U438 (N_438,In_391,In_871);
xnor U439 (N_439,In_383,In_636);
and U440 (N_440,In_57,In_466);
nor U441 (N_441,In_483,In_1032);
xnor U442 (N_442,In_693,In_363);
and U443 (N_443,In_825,In_37);
xnor U444 (N_444,In_1254,In_1473);
nand U445 (N_445,In_31,In_310);
or U446 (N_446,In_892,In_268);
or U447 (N_447,In_1342,In_702);
nand U448 (N_448,In_645,In_1232);
or U449 (N_449,In_1434,In_550);
and U450 (N_450,In_1203,In_409);
or U451 (N_451,In_1481,In_625);
nand U452 (N_452,In_749,In_1454);
nand U453 (N_453,In_424,In_198);
nand U454 (N_454,In_1054,In_877);
nand U455 (N_455,In_162,In_196);
xnor U456 (N_456,In_1003,In_1262);
and U457 (N_457,In_654,In_991);
xor U458 (N_458,In_570,In_395);
nor U459 (N_459,In_1183,In_1045);
nand U460 (N_460,In_455,In_299);
xnor U461 (N_461,In_724,In_778);
nor U462 (N_462,In_1284,In_1148);
or U463 (N_463,In_1204,In_382);
or U464 (N_464,In_318,In_1091);
nor U465 (N_465,In_481,In_968);
nor U466 (N_466,In_170,In_589);
or U467 (N_467,In_910,In_1301);
xnor U468 (N_468,In_329,In_106);
xnor U469 (N_469,In_1429,In_42);
and U470 (N_470,In_676,In_145);
nand U471 (N_471,In_164,In_343);
nor U472 (N_472,In_797,In_1421);
xor U473 (N_473,In_86,In_172);
nand U474 (N_474,In_51,In_369);
or U475 (N_475,In_976,In_85);
nor U476 (N_476,In_1472,In_698);
and U477 (N_477,In_1231,In_222);
nand U478 (N_478,In_535,In_1156);
or U479 (N_479,In_1413,In_941);
xor U480 (N_480,In_817,In_12);
xor U481 (N_481,In_757,In_328);
nor U482 (N_482,In_557,In_1213);
nand U483 (N_483,In_1468,In_511);
nand U484 (N_484,In_80,In_1247);
nand U485 (N_485,In_590,In_598);
and U486 (N_486,In_422,In_730);
nor U487 (N_487,In_1131,In_387);
and U488 (N_488,In_499,In_652);
xnor U489 (N_489,In_95,In_380);
nand U490 (N_490,In_1260,In_1241);
nand U491 (N_491,In_302,In_1237);
nand U492 (N_492,In_620,In_1348);
xnor U493 (N_493,In_1036,In_579);
or U494 (N_494,In_296,In_384);
or U495 (N_495,In_1009,In_400);
xor U496 (N_496,In_930,In_1498);
nor U497 (N_497,In_1,In_1178);
nor U498 (N_498,In_760,In_675);
nor U499 (N_499,In_117,In_128);
nand U500 (N_500,In_1160,N_185);
nor U501 (N_501,N_255,N_119);
and U502 (N_502,In_510,N_410);
nand U503 (N_503,N_115,N_128);
nor U504 (N_504,In_935,N_136);
and U505 (N_505,In_118,In_1287);
nor U506 (N_506,In_507,In_8);
or U507 (N_507,In_190,In_556);
or U508 (N_508,In_201,N_281);
nor U509 (N_509,In_831,In_176);
or U510 (N_510,N_10,N_50);
and U511 (N_511,In_584,N_144);
xor U512 (N_512,N_365,N_104);
or U513 (N_513,In_295,N_343);
xnor U514 (N_514,N_112,In_572);
or U515 (N_515,In_566,N_26);
nor U516 (N_516,N_97,In_634);
nor U517 (N_517,In_551,In_67);
xor U518 (N_518,In_1431,N_456);
xnor U519 (N_519,N_205,In_259);
and U520 (N_520,N_127,In_404);
nor U521 (N_521,N_229,In_214);
nand U522 (N_522,N_67,In_237);
nor U523 (N_523,In_55,N_325);
or U524 (N_524,N_161,In_1165);
xnor U525 (N_525,N_147,In_200);
and U526 (N_526,In_998,In_242);
or U527 (N_527,In_669,N_227);
xor U528 (N_528,In_282,In_1402);
or U529 (N_529,N_439,In_1066);
and U530 (N_530,In_179,In_872);
xor U531 (N_531,In_529,N_36);
xor U532 (N_532,In_397,In_608);
nor U533 (N_533,In_54,In_642);
nor U534 (N_534,In_66,In_9);
nor U535 (N_535,N_443,In_1113);
or U536 (N_536,In_1187,In_670);
xor U537 (N_537,In_386,In_1186);
xnor U538 (N_538,N_43,N_254);
or U539 (N_539,N_95,In_982);
nor U540 (N_540,In_1121,N_485);
nand U541 (N_541,N_352,N_186);
nand U542 (N_542,N_79,N_187);
xor U543 (N_543,In_558,N_368);
or U544 (N_544,N_350,In_808);
nand U545 (N_545,N_320,N_271);
xnor U546 (N_546,N_155,N_435);
nand U547 (N_547,N_253,N_129);
nor U548 (N_548,N_483,In_71);
and U549 (N_549,N_324,N_18);
and U550 (N_550,N_58,N_25);
nand U551 (N_551,In_209,N_384);
nor U552 (N_552,In_1089,In_988);
and U553 (N_553,In_1087,In_793);
nand U554 (N_554,N_85,In_1446);
nor U555 (N_555,In_494,N_474);
nor U556 (N_556,N_179,In_1278);
xor U557 (N_557,N_301,In_288);
and U558 (N_558,In_860,In_339);
and U559 (N_559,In_52,In_1154);
xnor U560 (N_560,N_231,N_211);
and U561 (N_561,In_616,N_134);
or U562 (N_562,N_453,In_125);
xnor U563 (N_563,In_1068,N_302);
nand U564 (N_564,N_472,In_542);
xor U565 (N_565,In_433,N_295);
and U566 (N_566,N_304,In_452);
nand U567 (N_567,N_45,N_234);
and U568 (N_568,N_489,In_1193);
xor U569 (N_569,N_65,In_873);
nor U570 (N_570,N_44,N_398);
nand U571 (N_571,N_455,In_279);
or U572 (N_572,In_442,In_1227);
or U573 (N_573,In_437,In_714);
nand U574 (N_574,N_284,In_996);
and U575 (N_575,In_972,N_82);
nand U576 (N_576,In_4,N_338);
and U577 (N_577,N_329,N_192);
and U578 (N_578,In_1263,N_375);
and U579 (N_579,N_286,N_7);
nor U580 (N_580,In_149,In_223);
or U581 (N_581,N_189,N_333);
or U582 (N_582,In_603,N_233);
nand U583 (N_583,N_174,N_240);
xor U584 (N_584,N_105,In_1170);
nand U585 (N_585,N_321,N_242);
nand U586 (N_586,N_117,In_826);
nand U587 (N_587,N_225,N_402);
or U588 (N_588,N_34,In_661);
xnor U589 (N_589,N_354,In_40);
nand U590 (N_590,In_564,N_63);
or U591 (N_591,In_1411,In_471);
nand U592 (N_592,N_389,In_253);
nor U593 (N_593,N_265,In_646);
or U594 (N_594,In_1305,N_154);
and U595 (N_595,N_118,In_780);
or U596 (N_596,In_1233,N_369);
nand U597 (N_597,In_837,In_1298);
nor U598 (N_598,In_599,In_342);
nor U599 (N_599,N_262,In_1339);
nor U600 (N_600,In_1107,N_109);
or U601 (N_601,N_54,In_272);
or U602 (N_602,N_38,N_303);
nor U603 (N_603,In_555,N_431);
xnor U604 (N_604,N_376,N_35);
and U605 (N_605,In_707,In_948);
and U606 (N_606,N_280,In_888);
nor U607 (N_607,In_767,N_392);
and U608 (N_608,In_152,N_120);
or U609 (N_609,N_148,N_313);
and U610 (N_610,In_97,N_101);
nor U611 (N_611,N_149,N_210);
nor U612 (N_612,In_265,In_360);
or U613 (N_613,In_794,In_347);
nor U614 (N_614,In_1249,In_74);
xnor U615 (N_615,N_417,In_1161);
nand U616 (N_616,N_33,In_1407);
nand U617 (N_617,N_228,N_88);
or U618 (N_618,N_94,In_269);
and U619 (N_619,In_653,N_305);
and U620 (N_620,N_257,In_947);
or U621 (N_621,N_145,In_1317);
and U622 (N_622,In_264,In_617);
nand U623 (N_623,N_459,In_1212);
xnor U624 (N_624,N_223,In_429);
xor U625 (N_625,N_486,In_1433);
or U626 (N_626,In_375,In_1229);
and U627 (N_627,In_306,N_158);
nand U628 (N_628,N_449,N_407);
nand U629 (N_629,N_465,N_66);
nand U630 (N_630,N_220,In_956);
and U631 (N_631,In_739,N_201);
nand U632 (N_632,In_1388,N_51);
nor U633 (N_633,In_1357,N_47);
nor U634 (N_634,In_1125,In_1293);
and U635 (N_635,N_414,N_328);
nor U636 (N_636,N_468,N_244);
and U637 (N_637,N_125,In_789);
or U638 (N_638,N_351,N_74);
nor U639 (N_639,N_124,N_380);
nor U640 (N_640,In_601,N_497);
and U641 (N_641,N_311,In_918);
or U642 (N_642,N_81,N_470);
or U643 (N_643,N_96,In_337);
xor U644 (N_644,In_963,In_61);
and U645 (N_645,N_230,In_405);
nand U646 (N_646,N_172,N_41);
nand U647 (N_647,N_256,N_217);
nor U648 (N_648,In_236,In_975);
nor U649 (N_649,In_345,In_674);
and U650 (N_650,In_874,In_1484);
nand U651 (N_651,In_841,In_1230);
and U652 (N_652,In_1159,N_294);
xor U653 (N_653,In_112,In_1460);
nand U654 (N_654,In_677,In_1070);
xor U655 (N_655,In_986,N_306);
or U656 (N_656,In_1085,In_684);
xor U657 (N_657,N_107,N_131);
nand U658 (N_658,N_499,In_1141);
or U659 (N_659,N_143,In_235);
or U660 (N_660,In_1430,In_353);
and U661 (N_661,N_421,In_1300);
or U662 (N_662,In_648,N_367);
and U663 (N_663,N_53,In_1482);
or U664 (N_664,N_77,N_90);
and U665 (N_665,N_12,In_1245);
xor U666 (N_666,In_274,In_454);
nor U667 (N_667,N_471,In_1133);
nor U668 (N_668,N_441,N_283);
nand U669 (N_669,N_454,N_278);
nor U670 (N_670,N_213,N_222);
or U671 (N_671,In_1011,In_962);
and U672 (N_672,N_226,N_490);
xnor U673 (N_673,In_1415,N_492);
nor U674 (N_674,In_658,In_899);
and U675 (N_675,In_538,In_1417);
and U676 (N_676,In_1020,N_184);
nand U677 (N_677,N_473,N_251);
xor U678 (N_678,N_91,N_360);
xor U679 (N_679,N_123,N_93);
and U680 (N_680,In_1086,In_411);
or U681 (N_681,In_990,In_663);
xnor U682 (N_682,In_63,N_113);
xor U683 (N_683,N_9,In_1025);
and U684 (N_684,N_14,In_82);
and U685 (N_685,In_830,N_195);
nor U686 (N_686,N_73,N_336);
nand U687 (N_687,In_281,In_147);
and U688 (N_688,N_363,In_1362);
and U689 (N_689,In_791,In_1321);
and U690 (N_690,N_23,N_122);
or U691 (N_691,N_173,In_1302);
or U692 (N_692,In_536,N_248);
nor U693 (N_693,In_138,N_175);
nor U694 (N_694,N_70,In_902);
nor U695 (N_695,N_344,In_1360);
and U696 (N_696,In_560,N_219);
or U697 (N_697,N_275,In_907);
or U698 (N_698,In_478,In_378);
or U699 (N_699,N_422,In_327);
and U700 (N_700,In_1197,In_800);
nor U701 (N_701,In_157,N_106);
and U702 (N_702,In_1205,In_576);
xnor U703 (N_703,In_168,N_37);
and U704 (N_704,In_858,In_1347);
or U705 (N_705,N_153,In_703);
and U706 (N_706,In_1448,N_214);
nand U707 (N_707,In_225,In_250);
or U708 (N_708,N_261,In_139);
xnor U709 (N_709,In_266,N_296);
or U710 (N_710,N_387,In_485);
and U711 (N_711,N_52,N_133);
xor U712 (N_712,N_42,N_335);
and U713 (N_713,N_318,N_6);
nor U714 (N_714,In_628,N_345);
or U715 (N_715,N_493,N_64);
xnor U716 (N_716,N_159,In_1120);
or U717 (N_717,In_1151,N_377);
and U718 (N_718,In_1220,In_1080);
or U719 (N_719,N_13,N_371);
nor U720 (N_720,N_146,N_243);
xor U721 (N_721,In_949,In_305);
or U722 (N_722,N_29,In_1015);
and U723 (N_723,In_217,In_640);
nand U724 (N_724,N_481,N_498);
xor U725 (N_725,In_416,N_200);
xor U726 (N_726,N_496,In_140);
xor U727 (N_727,N_452,N_362);
nor U728 (N_728,N_263,N_272);
nor U729 (N_729,N_2,In_102);
nand U730 (N_730,N_269,N_224);
and U731 (N_731,In_124,N_49);
nor U732 (N_732,In_562,N_22);
nand U733 (N_733,In_11,In_239);
xnor U734 (N_734,In_34,In_1194);
or U735 (N_735,In_924,In_451);
nor U736 (N_736,In_549,N_382);
xnor U737 (N_737,In_216,In_1207);
nor U738 (N_738,In_1461,N_89);
and U739 (N_739,N_237,N_273);
and U740 (N_740,N_98,In_229);
nand U741 (N_741,In_712,N_206);
xnor U742 (N_742,In_69,In_77);
nor U743 (N_743,N_24,N_349);
xnor U744 (N_744,N_478,N_142);
nor U745 (N_745,In_1144,N_204);
nor U746 (N_746,N_442,N_317);
nand U747 (N_747,N_406,N_78);
xnor U748 (N_748,N_432,N_258);
nand U749 (N_749,N_28,In_267);
nor U750 (N_750,In_581,N_334);
nor U751 (N_751,N_287,N_433);
nor U752 (N_752,In_612,In_46);
nand U753 (N_753,In_244,In_1419);
or U754 (N_754,N_102,N_157);
and U755 (N_755,N_193,N_183);
nor U756 (N_756,N_135,N_171);
nand U757 (N_757,N_268,In_207);
nand U758 (N_758,N_27,N_319);
nor U759 (N_759,N_277,In_908);
nor U760 (N_760,In_1479,In_1285);
and U761 (N_761,N_416,In_967);
nor U762 (N_762,In_751,In_1492);
nor U763 (N_763,In_144,N_446);
and U764 (N_764,N_482,In_573);
and U765 (N_765,N_322,N_202);
and U766 (N_766,In_131,N_130);
xor U767 (N_767,In_904,In_493);
nor U768 (N_768,N_342,N_32);
nand U769 (N_769,In_734,In_159);
or U770 (N_770,N_346,N_425);
xor U771 (N_771,In_1311,In_886);
and U772 (N_772,N_209,In_1208);
xor U773 (N_773,In_173,In_1351);
nand U774 (N_774,N_264,N_420);
or U775 (N_775,In_514,N_467);
nor U776 (N_776,N_163,In_1396);
and U777 (N_777,In_96,In_488);
nand U778 (N_778,In_153,N_21);
nor U779 (N_779,In_540,N_290);
nand U780 (N_780,N_458,N_494);
xor U781 (N_781,N_394,In_811);
or U782 (N_782,In_1401,N_68);
and U783 (N_783,N_475,N_339);
nor U784 (N_784,N_293,In_1238);
xnor U785 (N_785,In_472,In_1310);
xor U786 (N_786,N_393,In_430);
nor U787 (N_787,In_1297,In_1328);
or U788 (N_788,In_940,N_358);
nor U789 (N_789,N_450,In_64);
nand U790 (N_790,In_1173,N_20);
nand U791 (N_791,N_238,In_291);
nand U792 (N_792,In_1368,In_100);
xor U793 (N_793,N_56,N_403);
xnor U794 (N_794,In_1038,In_1378);
or U795 (N_795,In_374,In_600);
xnor U796 (N_796,N_156,N_379);
nand U797 (N_797,In_243,In_867);
xnor U798 (N_798,In_1463,N_141);
and U799 (N_799,In_633,N_137);
xnor U800 (N_800,N_86,In_842);
xnor U801 (N_801,N_167,In_1338);
xor U802 (N_802,In_467,In_1050);
nand U803 (N_803,N_419,In_1110);
nor U804 (N_804,N_162,In_204);
or U805 (N_805,N_252,In_1397);
and U806 (N_806,In_1256,N_408);
xor U807 (N_807,In_559,N_359);
xor U808 (N_808,N_182,In_84);
nand U809 (N_809,In_496,In_326);
nand U810 (N_810,N_330,N_221);
nand U811 (N_811,N_17,N_245);
and U812 (N_812,N_445,In_1072);
xor U813 (N_813,In_142,N_126);
nor U814 (N_814,In_627,In_448);
nand U815 (N_815,In_156,In_803);
or U816 (N_816,In_1352,In_520);
or U817 (N_817,N_270,N_463);
nor U818 (N_818,In_783,N_266);
or U819 (N_819,N_388,In_1146);
nor U820 (N_820,In_1037,In_1474);
or U821 (N_821,N_462,N_466);
and U822 (N_822,N_75,N_464);
and U823 (N_823,N_282,N_327);
and U824 (N_824,In_1437,N_477);
nor U825 (N_825,N_178,In_756);
xnor U826 (N_826,N_487,N_30);
nand U827 (N_827,In_463,In_58);
nand U828 (N_828,N_373,In_16);
nor U829 (N_829,In_1395,In_668);
nor U830 (N_830,N_176,N_207);
nand U831 (N_831,N_391,N_381);
nor U832 (N_832,N_397,In_336);
nor U833 (N_833,In_618,In_582);
nor U834 (N_834,N_337,In_468);
or U835 (N_835,N_423,In_995);
nand U836 (N_836,N_138,In_1447);
or U837 (N_837,N_341,N_267);
or U838 (N_838,N_434,N_438);
nor U839 (N_839,In_1294,N_332);
nor U840 (N_840,In_741,In_552);
nand U841 (N_841,In_331,N_164);
nand U842 (N_842,N_40,In_528);
nand U843 (N_843,In_1383,In_1176);
nor U844 (N_844,N_241,In_1210);
xnor U845 (N_845,In_181,In_1051);
nand U846 (N_846,In_629,In_304);
nor U847 (N_847,In_426,In_926);
nand U848 (N_848,In_818,N_461);
or U849 (N_849,N_429,In_1211);
nand U850 (N_850,In_1083,In_909);
and U851 (N_851,N_347,In_449);
xor U852 (N_852,In_143,In_852);
nand U853 (N_853,In_1044,N_5);
and U854 (N_854,In_1199,N_405);
nand U855 (N_855,N_411,N_4);
xor U856 (N_856,N_340,In_1376);
and U857 (N_857,In_735,N_298);
nand U858 (N_858,In_758,In_750);
nor U859 (N_859,N_60,N_315);
or U860 (N_860,In_1058,In_312);
nand U861 (N_861,In_914,In_446);
nand U862 (N_862,N_215,N_212);
or U863 (N_863,In_1350,N_447);
or U864 (N_864,N_395,In_498);
xor U865 (N_865,N_364,N_378);
or U866 (N_866,N_218,In_691);
and U867 (N_867,In_1282,N_259);
or U868 (N_868,In_1389,N_396);
nand U869 (N_869,In_447,N_418);
nor U870 (N_870,In_1105,N_191);
nor U871 (N_871,N_289,In_1405);
and U872 (N_872,N_170,In_220);
and U873 (N_873,N_250,N_166);
nand U874 (N_874,N_197,N_46);
nand U875 (N_875,N_401,In_252);
nor U876 (N_876,In_365,In_509);
nor U877 (N_877,N_357,In_678);
xor U878 (N_878,N_314,N_323);
or U879 (N_879,N_15,In_1195);
xnor U880 (N_880,In_656,In_890);
nand U881 (N_881,In_1459,N_100);
and U882 (N_882,In_1073,In_518);
and U883 (N_883,N_132,N_83);
xor U884 (N_884,In_486,In_1488);
and U885 (N_885,In_1271,N_372);
nand U886 (N_886,In_752,In_931);
nor U887 (N_887,N_190,In_1439);
or U888 (N_888,N_31,N_374);
xnor U889 (N_889,N_288,N_199);
or U890 (N_890,N_71,In_333);
or U891 (N_891,In_110,N_59);
or U892 (N_892,In_48,N_469);
nor U893 (N_893,In_571,In_814);
and U894 (N_894,In_715,N_415);
and U895 (N_895,N_99,In_7);
xor U896 (N_896,In_785,N_386);
or U897 (N_897,In_171,In_727);
xnor U898 (N_898,In_719,In_650);
or U899 (N_899,In_943,N_491);
xor U900 (N_900,In_999,In_894);
and U901 (N_901,N_383,N_299);
nor U902 (N_902,In_1267,In_134);
xnor U903 (N_903,In_370,In_913);
nor U904 (N_904,In_322,N_0);
or U905 (N_905,N_236,N_151);
nor U906 (N_906,N_430,N_16);
xnor U907 (N_907,N_177,In_465);
xor U908 (N_908,N_121,N_140);
nand U909 (N_909,In_1196,In_418);
nor U910 (N_910,In_631,In_1276);
nand U911 (N_911,N_181,In_544);
nor U912 (N_912,N_460,N_451);
nor U913 (N_913,N_316,In_1471);
nor U914 (N_914,N_353,N_495);
xor U915 (N_915,In_109,N_249);
xnor U916 (N_916,N_404,N_260);
or U917 (N_917,In_1128,In_19);
xor U918 (N_918,N_348,N_308);
xnor U919 (N_919,N_356,In_746);
nand U920 (N_920,N_484,In_22);
nor U921 (N_921,N_196,In_534);
nand U922 (N_922,In_737,In_1214);
and U923 (N_923,N_246,N_399);
nor U924 (N_924,In_434,N_92);
nor U925 (N_925,In_101,N_300);
or U926 (N_926,In_228,In_241);
nor U927 (N_927,N_440,In_357);
nor U928 (N_928,N_366,N_232);
nor U929 (N_929,N_285,In_891);
nor U930 (N_930,N_488,N_309);
and U931 (N_931,N_39,In_920);
and U932 (N_932,In_1436,N_480);
and U933 (N_933,In_98,N_150);
nand U934 (N_934,N_48,N_361);
nor U935 (N_935,In_1261,N_424);
nor U936 (N_936,In_410,N_198);
or U937 (N_937,In_577,In_461);
and U938 (N_938,In_1250,In_1081);
and U939 (N_939,N_412,N_326);
and U940 (N_940,In_1029,In_936);
or U941 (N_941,N_116,N_291);
nand U942 (N_942,In_742,N_69);
and U943 (N_943,In_344,In_1330);
or U944 (N_944,In_1364,N_239);
nor U945 (N_945,In_615,N_180);
nor U946 (N_946,In_277,N_169);
or U947 (N_947,In_1028,In_955);
and U948 (N_948,N_139,N_160);
nor U949 (N_949,In_578,In_169);
xnor U950 (N_950,In_513,N_80);
nand U951 (N_951,In_1076,In_1093);
or U952 (N_952,In_189,N_448);
xnor U953 (N_953,N_310,In_130);
or U954 (N_954,N_87,N_279);
and U955 (N_955,In_639,N_55);
nand U956 (N_956,In_798,N_312);
xor U957 (N_957,In_293,N_103);
nand U958 (N_958,In_630,N_409);
nand U959 (N_959,In_1150,In_28);
xnor U960 (N_960,N_57,In_87);
nor U961 (N_961,N_114,N_331);
xnor U962 (N_962,In_533,In_586);
nand U963 (N_963,In_1320,In_1188);
and U964 (N_964,N_370,N_476);
xnor U965 (N_965,In_666,In_492);
or U966 (N_966,N_292,N_62);
nand U967 (N_967,N_168,N_274);
and U968 (N_968,In_848,N_436);
xor U969 (N_969,N_1,In_459);
nand U970 (N_970,N_84,N_428);
or U971 (N_971,N_297,In_1408);
and U972 (N_972,In_795,In_1136);
nand U973 (N_973,In_786,N_8);
nand U974 (N_974,In_713,N_76);
xnor U975 (N_975,In_1273,N_208);
nor U976 (N_976,N_437,In_813);
xnor U977 (N_977,N_276,In_1336);
nor U978 (N_978,In_839,N_413);
or U979 (N_979,In_1493,N_3);
or U980 (N_980,In_1372,N_19);
or U981 (N_981,N_390,N_110);
nand U982 (N_982,In_33,N_247);
xor U983 (N_983,N_108,N_479);
xor U984 (N_984,In_284,N_165);
xnor U985 (N_985,In_1414,N_235);
nand U986 (N_986,N_426,N_11);
and U987 (N_987,N_203,N_216);
nor U988 (N_988,In_1387,N_61);
nand U989 (N_989,N_355,N_457);
or U990 (N_990,In_699,N_194);
nor U991 (N_991,N_188,N_72);
xor U992 (N_992,N_385,In_753);
xor U993 (N_993,N_111,N_444);
and U994 (N_994,N_152,N_307);
and U995 (N_995,In_602,In_722);
nor U996 (N_996,In_1406,In_1002);
nor U997 (N_997,N_400,In_1255);
and U998 (N_998,In_83,In_103);
nor U999 (N_999,N_427,In_1295);
xor U1000 (N_1000,N_820,N_534);
and U1001 (N_1001,N_964,N_619);
and U1002 (N_1002,N_547,N_985);
xor U1003 (N_1003,N_556,N_532);
nand U1004 (N_1004,N_613,N_840);
or U1005 (N_1005,N_968,N_707);
and U1006 (N_1006,N_784,N_722);
or U1007 (N_1007,N_924,N_746);
or U1008 (N_1008,N_848,N_526);
or U1009 (N_1009,N_600,N_729);
nand U1010 (N_1010,N_635,N_756);
or U1011 (N_1011,N_826,N_925);
or U1012 (N_1012,N_792,N_508);
and U1013 (N_1013,N_861,N_805);
xor U1014 (N_1014,N_793,N_958);
xnor U1015 (N_1015,N_759,N_815);
nor U1016 (N_1016,N_966,N_767);
and U1017 (N_1017,N_989,N_507);
xor U1018 (N_1018,N_592,N_512);
nand U1019 (N_1019,N_970,N_975);
nor U1020 (N_1020,N_525,N_879);
nand U1021 (N_1021,N_806,N_940);
xor U1022 (N_1022,N_655,N_789);
xor U1023 (N_1023,N_560,N_910);
nor U1024 (N_1024,N_704,N_689);
xnor U1025 (N_1025,N_607,N_736);
nor U1026 (N_1026,N_943,N_771);
nand U1027 (N_1027,N_680,N_571);
nand U1028 (N_1028,N_570,N_768);
and U1029 (N_1029,N_593,N_763);
or U1030 (N_1030,N_888,N_730);
or U1031 (N_1031,N_794,N_780);
or U1032 (N_1032,N_521,N_726);
xor U1033 (N_1033,N_732,N_823);
or U1034 (N_1034,N_828,N_865);
or U1035 (N_1035,N_682,N_870);
nor U1036 (N_1036,N_891,N_646);
nand U1037 (N_1037,N_629,N_700);
or U1038 (N_1038,N_912,N_856);
nor U1039 (N_1039,N_615,N_548);
or U1040 (N_1040,N_941,N_745);
xor U1041 (N_1041,N_765,N_712);
nand U1042 (N_1042,N_850,N_749);
nand U1043 (N_1043,N_788,N_558);
nand U1044 (N_1044,N_808,N_731);
nand U1045 (N_1045,N_775,N_995);
xnor U1046 (N_1046,N_790,N_603);
or U1047 (N_1047,N_540,N_810);
nand U1048 (N_1048,N_976,N_514);
or U1049 (N_1049,N_761,N_980);
or U1050 (N_1050,N_935,N_798);
nor U1051 (N_1051,N_868,N_596);
nor U1052 (N_1052,N_817,N_921);
and U1053 (N_1053,N_881,N_727);
nor U1054 (N_1054,N_541,N_754);
nand U1055 (N_1055,N_695,N_892);
nor U1056 (N_1056,N_679,N_711);
nor U1057 (N_1057,N_698,N_647);
xnor U1058 (N_1058,N_564,N_543);
nor U1059 (N_1059,N_779,N_716);
and U1060 (N_1060,N_758,N_533);
xnor U1061 (N_1061,N_516,N_957);
xor U1062 (N_1062,N_650,N_833);
xor U1063 (N_1063,N_709,N_530);
xor U1064 (N_1064,N_670,N_874);
nor U1065 (N_1065,N_623,N_649);
nand U1066 (N_1066,N_831,N_979);
nor U1067 (N_1067,N_760,N_883);
and U1068 (N_1068,N_747,N_671);
nor U1069 (N_1069,N_737,N_956);
and U1070 (N_1070,N_869,N_782);
and U1071 (N_1071,N_664,N_787);
or U1072 (N_1072,N_847,N_841);
xnor U1073 (N_1073,N_837,N_785);
nor U1074 (N_1074,N_813,N_836);
or U1075 (N_1075,N_901,N_987);
and U1076 (N_1076,N_626,N_706);
or U1077 (N_1077,N_984,N_648);
and U1078 (N_1078,N_988,N_884);
nand U1079 (N_1079,N_755,N_645);
nor U1080 (N_1080,N_529,N_838);
and U1081 (N_1081,N_911,N_963);
nand U1082 (N_1082,N_797,N_853);
nand U1083 (N_1083,N_715,N_520);
and U1084 (N_1084,N_550,N_799);
or U1085 (N_1085,N_574,N_518);
nand U1086 (N_1086,N_693,N_630);
and U1087 (N_1087,N_686,N_934);
nor U1088 (N_1088,N_777,N_886);
nor U1089 (N_1089,N_555,N_703);
nand U1090 (N_1090,N_948,N_708);
xnor U1091 (N_1091,N_897,N_800);
and U1092 (N_1092,N_959,N_751);
and U1093 (N_1093,N_538,N_513);
xnor U1094 (N_1094,N_617,N_567);
or U1095 (N_1095,N_927,N_791);
xnor U1096 (N_1096,N_952,N_658);
nand U1097 (N_1097,N_589,N_855);
nand U1098 (N_1098,N_922,N_599);
or U1099 (N_1099,N_931,N_638);
and U1100 (N_1100,N_981,N_580);
nand U1101 (N_1101,N_738,N_864);
and U1102 (N_1102,N_662,N_601);
nand U1103 (N_1103,N_565,N_535);
and U1104 (N_1104,N_620,N_858);
xor U1105 (N_1105,N_774,N_844);
or U1106 (N_1106,N_559,N_644);
nor U1107 (N_1107,N_549,N_812);
nor U1108 (N_1108,N_895,N_926);
or U1109 (N_1109,N_531,N_669);
xnor U1110 (N_1110,N_871,N_504);
nand U1111 (N_1111,N_552,N_832);
nand U1112 (N_1112,N_898,N_661);
xor U1113 (N_1113,N_906,N_714);
and U1114 (N_1114,N_632,N_677);
or U1115 (N_1115,N_683,N_676);
and U1116 (N_1116,N_656,N_809);
xnor U1117 (N_1117,N_743,N_503);
or U1118 (N_1118,N_945,N_867);
xor U1119 (N_1119,N_667,N_586);
xor U1120 (N_1120,N_528,N_876);
nand U1121 (N_1121,N_652,N_590);
nand U1122 (N_1122,N_843,N_933);
nor U1123 (N_1123,N_889,N_909);
nand U1124 (N_1124,N_699,N_877);
and U1125 (N_1125,N_939,N_829);
and U1126 (N_1126,N_719,N_973);
nor U1127 (N_1127,N_778,N_953);
xor U1128 (N_1128,N_986,N_852);
and U1129 (N_1129,N_748,N_666);
xor U1130 (N_1130,N_795,N_969);
xor U1131 (N_1131,N_938,N_578);
xor U1132 (N_1132,N_675,N_576);
nor U1133 (N_1133,N_903,N_611);
xor U1134 (N_1134,N_916,N_811);
xnor U1135 (N_1135,N_694,N_502);
and U1136 (N_1136,N_851,N_505);
or U1137 (N_1137,N_752,N_796);
xor U1138 (N_1138,N_998,N_557);
xor U1139 (N_1139,N_978,N_882);
xor U1140 (N_1140,N_899,N_673);
nor U1141 (N_1141,N_621,N_539);
or U1142 (N_1142,N_723,N_977);
xor U1143 (N_1143,N_907,N_517);
and U1144 (N_1144,N_818,N_955);
and U1145 (N_1145,N_622,N_616);
nand U1146 (N_1146,N_604,N_510);
and U1147 (N_1147,N_554,N_872);
or U1148 (N_1148,N_511,N_690);
nand U1149 (N_1149,N_928,N_577);
nand U1150 (N_1150,N_983,N_902);
or U1151 (N_1151,N_942,N_572);
nand U1152 (N_1152,N_993,N_522);
or U1153 (N_1153,N_643,N_608);
nor U1154 (N_1154,N_612,N_672);
xnor U1155 (N_1155,N_713,N_542);
xnor U1156 (N_1156,N_741,N_739);
nor U1157 (N_1157,N_807,N_972);
xnor U1158 (N_1158,N_725,N_653);
or U1159 (N_1159,N_637,N_609);
or U1160 (N_1160,N_750,N_606);
xnor U1161 (N_1161,N_866,N_610);
nand U1162 (N_1162,N_825,N_918);
nand U1163 (N_1163,N_618,N_814);
nand U1164 (N_1164,N_579,N_859);
and U1165 (N_1165,N_821,N_873);
and U1166 (N_1166,N_830,N_660);
or U1167 (N_1167,N_802,N_893);
nor U1168 (N_1168,N_718,N_905);
nand U1169 (N_1169,N_949,N_890);
or U1170 (N_1170,N_932,N_947);
nand U1171 (N_1171,N_994,N_584);
nand U1172 (N_1172,N_816,N_701);
nand U1173 (N_1173,N_900,N_597);
nor U1174 (N_1174,N_685,N_929);
or U1175 (N_1175,N_923,N_999);
xor U1176 (N_1176,N_733,N_634);
xnor U1177 (N_1177,N_720,N_946);
and U1178 (N_1178,N_515,N_974);
or U1179 (N_1179,N_551,N_640);
or U1180 (N_1180,N_896,N_566);
nor U1181 (N_1181,N_857,N_875);
or U1182 (N_1182,N_786,N_735);
xnor U1183 (N_1183,N_501,N_692);
nand U1184 (N_1184,N_951,N_849);
or U1185 (N_1185,N_688,N_684);
and U1186 (N_1186,N_764,N_996);
xnor U1187 (N_1187,N_598,N_509);
xnor U1188 (N_1188,N_681,N_696);
and U1189 (N_1189,N_581,N_654);
or U1190 (N_1190,N_887,N_967);
xor U1191 (N_1191,N_721,N_642);
nand U1192 (N_1192,N_631,N_545);
nor U1193 (N_1193,N_628,N_573);
nand U1194 (N_1194,N_705,N_633);
nor U1195 (N_1195,N_781,N_917);
and U1196 (N_1196,N_950,N_663);
xor U1197 (N_1197,N_659,N_668);
and U1198 (N_1198,N_863,N_553);
and U1199 (N_1199,N_568,N_527);
nand U1200 (N_1200,N_657,N_762);
or U1201 (N_1201,N_740,N_845);
or U1202 (N_1202,N_744,N_776);
nor U1203 (N_1203,N_920,N_536);
xnor U1204 (N_1204,N_561,N_724);
nor U1205 (N_1205,N_991,N_962);
xor U1206 (N_1206,N_627,N_687);
nand U1207 (N_1207,N_624,N_537);
xnor U1208 (N_1208,N_766,N_804);
or U1209 (N_1209,N_728,N_717);
nor U1210 (N_1210,N_734,N_944);
or U1211 (N_1211,N_591,N_783);
and U1212 (N_1212,N_960,N_835);
or U1213 (N_1213,N_880,N_674);
and U1214 (N_1214,N_625,N_753);
nor U1215 (N_1215,N_913,N_594);
and U1216 (N_1216,N_500,N_819);
nor U1217 (N_1217,N_954,N_636);
nand U1218 (N_1218,N_842,N_990);
and U1219 (N_1219,N_961,N_562);
and U1220 (N_1220,N_639,N_757);
nand U1221 (N_1221,N_585,N_678);
xnor U1222 (N_1222,N_506,N_575);
nor U1223 (N_1223,N_894,N_588);
or U1224 (N_1224,N_915,N_742);
nor U1225 (N_1225,N_665,N_614);
nand U1226 (N_1226,N_587,N_885);
and U1227 (N_1227,N_862,N_908);
nand U1228 (N_1228,N_803,N_914);
nand U1229 (N_1229,N_982,N_936);
xor U1230 (N_1230,N_770,N_930);
and U1231 (N_1231,N_992,N_641);
and U1232 (N_1232,N_702,N_846);
xor U1233 (N_1233,N_546,N_937);
nor U1234 (N_1234,N_772,N_519);
nor U1235 (N_1235,N_919,N_860);
or U1236 (N_1236,N_582,N_595);
xnor U1237 (N_1237,N_697,N_965);
nand U1238 (N_1238,N_822,N_710);
nor U1239 (N_1239,N_544,N_971);
nor U1240 (N_1240,N_691,N_769);
xor U1241 (N_1241,N_834,N_997);
or U1242 (N_1242,N_824,N_854);
or U1243 (N_1243,N_801,N_605);
nor U1244 (N_1244,N_524,N_523);
or U1245 (N_1245,N_904,N_827);
nor U1246 (N_1246,N_878,N_651);
xnor U1247 (N_1247,N_563,N_569);
nor U1248 (N_1248,N_583,N_839);
xnor U1249 (N_1249,N_602,N_773);
nor U1250 (N_1250,N_734,N_854);
or U1251 (N_1251,N_880,N_694);
nand U1252 (N_1252,N_909,N_546);
or U1253 (N_1253,N_704,N_634);
nand U1254 (N_1254,N_686,N_534);
and U1255 (N_1255,N_538,N_776);
nand U1256 (N_1256,N_756,N_895);
or U1257 (N_1257,N_987,N_599);
or U1258 (N_1258,N_676,N_720);
or U1259 (N_1259,N_876,N_809);
nor U1260 (N_1260,N_851,N_739);
xnor U1261 (N_1261,N_812,N_687);
xor U1262 (N_1262,N_563,N_585);
and U1263 (N_1263,N_506,N_736);
nor U1264 (N_1264,N_599,N_631);
nand U1265 (N_1265,N_827,N_533);
nor U1266 (N_1266,N_833,N_525);
and U1267 (N_1267,N_546,N_531);
nor U1268 (N_1268,N_558,N_563);
xor U1269 (N_1269,N_664,N_635);
or U1270 (N_1270,N_918,N_850);
nor U1271 (N_1271,N_884,N_729);
and U1272 (N_1272,N_527,N_593);
and U1273 (N_1273,N_743,N_849);
nor U1274 (N_1274,N_729,N_636);
nand U1275 (N_1275,N_770,N_851);
and U1276 (N_1276,N_671,N_993);
and U1277 (N_1277,N_971,N_700);
and U1278 (N_1278,N_671,N_977);
or U1279 (N_1279,N_989,N_839);
xor U1280 (N_1280,N_584,N_956);
and U1281 (N_1281,N_941,N_747);
or U1282 (N_1282,N_834,N_678);
nor U1283 (N_1283,N_698,N_894);
nor U1284 (N_1284,N_995,N_833);
nor U1285 (N_1285,N_592,N_584);
and U1286 (N_1286,N_893,N_973);
nand U1287 (N_1287,N_811,N_570);
xor U1288 (N_1288,N_801,N_823);
and U1289 (N_1289,N_596,N_933);
nand U1290 (N_1290,N_885,N_813);
and U1291 (N_1291,N_945,N_596);
or U1292 (N_1292,N_978,N_686);
xor U1293 (N_1293,N_735,N_873);
or U1294 (N_1294,N_693,N_752);
nor U1295 (N_1295,N_522,N_753);
nor U1296 (N_1296,N_856,N_709);
or U1297 (N_1297,N_738,N_765);
xor U1298 (N_1298,N_956,N_946);
and U1299 (N_1299,N_910,N_969);
or U1300 (N_1300,N_707,N_904);
xor U1301 (N_1301,N_601,N_697);
nor U1302 (N_1302,N_828,N_531);
xnor U1303 (N_1303,N_722,N_987);
xnor U1304 (N_1304,N_547,N_525);
nand U1305 (N_1305,N_660,N_769);
or U1306 (N_1306,N_602,N_571);
and U1307 (N_1307,N_610,N_577);
nand U1308 (N_1308,N_728,N_807);
nand U1309 (N_1309,N_631,N_709);
and U1310 (N_1310,N_855,N_957);
nor U1311 (N_1311,N_849,N_609);
and U1312 (N_1312,N_728,N_830);
nand U1313 (N_1313,N_764,N_798);
nor U1314 (N_1314,N_922,N_802);
nand U1315 (N_1315,N_599,N_853);
nand U1316 (N_1316,N_892,N_968);
nor U1317 (N_1317,N_839,N_523);
or U1318 (N_1318,N_884,N_822);
or U1319 (N_1319,N_612,N_860);
nand U1320 (N_1320,N_711,N_816);
nand U1321 (N_1321,N_962,N_616);
or U1322 (N_1322,N_944,N_750);
and U1323 (N_1323,N_830,N_674);
nand U1324 (N_1324,N_570,N_889);
nor U1325 (N_1325,N_736,N_873);
and U1326 (N_1326,N_646,N_708);
nor U1327 (N_1327,N_589,N_767);
xnor U1328 (N_1328,N_702,N_930);
xor U1329 (N_1329,N_831,N_503);
nand U1330 (N_1330,N_775,N_727);
xor U1331 (N_1331,N_985,N_799);
xnor U1332 (N_1332,N_657,N_731);
xor U1333 (N_1333,N_967,N_895);
and U1334 (N_1334,N_994,N_674);
and U1335 (N_1335,N_762,N_956);
xor U1336 (N_1336,N_785,N_927);
nor U1337 (N_1337,N_639,N_678);
or U1338 (N_1338,N_868,N_940);
or U1339 (N_1339,N_885,N_918);
or U1340 (N_1340,N_622,N_761);
or U1341 (N_1341,N_695,N_818);
nor U1342 (N_1342,N_562,N_993);
nor U1343 (N_1343,N_556,N_542);
and U1344 (N_1344,N_751,N_786);
xnor U1345 (N_1345,N_596,N_888);
and U1346 (N_1346,N_954,N_808);
nor U1347 (N_1347,N_541,N_750);
nor U1348 (N_1348,N_862,N_775);
xnor U1349 (N_1349,N_836,N_570);
nor U1350 (N_1350,N_649,N_731);
nand U1351 (N_1351,N_713,N_898);
xor U1352 (N_1352,N_964,N_763);
or U1353 (N_1353,N_526,N_902);
xnor U1354 (N_1354,N_945,N_756);
and U1355 (N_1355,N_623,N_944);
xor U1356 (N_1356,N_879,N_503);
nor U1357 (N_1357,N_500,N_820);
nor U1358 (N_1358,N_906,N_691);
and U1359 (N_1359,N_938,N_926);
and U1360 (N_1360,N_981,N_678);
nand U1361 (N_1361,N_974,N_697);
or U1362 (N_1362,N_665,N_547);
nand U1363 (N_1363,N_810,N_761);
and U1364 (N_1364,N_965,N_719);
nand U1365 (N_1365,N_532,N_559);
nand U1366 (N_1366,N_594,N_766);
nand U1367 (N_1367,N_737,N_770);
and U1368 (N_1368,N_763,N_709);
and U1369 (N_1369,N_982,N_528);
nor U1370 (N_1370,N_987,N_967);
nand U1371 (N_1371,N_650,N_606);
nand U1372 (N_1372,N_511,N_991);
xnor U1373 (N_1373,N_661,N_737);
nor U1374 (N_1374,N_957,N_955);
nand U1375 (N_1375,N_733,N_598);
nand U1376 (N_1376,N_714,N_655);
xor U1377 (N_1377,N_590,N_673);
nor U1378 (N_1378,N_840,N_750);
and U1379 (N_1379,N_902,N_800);
nand U1380 (N_1380,N_724,N_920);
and U1381 (N_1381,N_750,N_673);
nor U1382 (N_1382,N_605,N_809);
nor U1383 (N_1383,N_724,N_762);
or U1384 (N_1384,N_769,N_977);
nand U1385 (N_1385,N_618,N_910);
and U1386 (N_1386,N_894,N_570);
or U1387 (N_1387,N_596,N_780);
and U1388 (N_1388,N_881,N_840);
xor U1389 (N_1389,N_867,N_771);
and U1390 (N_1390,N_740,N_945);
xor U1391 (N_1391,N_523,N_956);
nor U1392 (N_1392,N_960,N_862);
xnor U1393 (N_1393,N_960,N_670);
nand U1394 (N_1394,N_771,N_878);
xor U1395 (N_1395,N_925,N_704);
or U1396 (N_1396,N_762,N_605);
nand U1397 (N_1397,N_738,N_574);
nor U1398 (N_1398,N_660,N_802);
or U1399 (N_1399,N_637,N_779);
or U1400 (N_1400,N_656,N_977);
and U1401 (N_1401,N_850,N_564);
nor U1402 (N_1402,N_959,N_641);
or U1403 (N_1403,N_717,N_520);
nor U1404 (N_1404,N_506,N_656);
and U1405 (N_1405,N_850,N_559);
and U1406 (N_1406,N_781,N_729);
xor U1407 (N_1407,N_965,N_728);
and U1408 (N_1408,N_810,N_832);
nand U1409 (N_1409,N_920,N_970);
nor U1410 (N_1410,N_621,N_661);
nand U1411 (N_1411,N_509,N_919);
or U1412 (N_1412,N_747,N_769);
nand U1413 (N_1413,N_585,N_892);
nor U1414 (N_1414,N_846,N_980);
or U1415 (N_1415,N_677,N_530);
nand U1416 (N_1416,N_953,N_577);
nand U1417 (N_1417,N_661,N_931);
or U1418 (N_1418,N_526,N_627);
or U1419 (N_1419,N_955,N_696);
xnor U1420 (N_1420,N_710,N_770);
or U1421 (N_1421,N_968,N_626);
nand U1422 (N_1422,N_702,N_851);
nand U1423 (N_1423,N_971,N_652);
and U1424 (N_1424,N_542,N_581);
or U1425 (N_1425,N_889,N_720);
or U1426 (N_1426,N_584,N_883);
xnor U1427 (N_1427,N_981,N_680);
nand U1428 (N_1428,N_896,N_644);
xnor U1429 (N_1429,N_888,N_645);
nor U1430 (N_1430,N_907,N_837);
or U1431 (N_1431,N_560,N_734);
nor U1432 (N_1432,N_973,N_853);
and U1433 (N_1433,N_840,N_993);
nor U1434 (N_1434,N_774,N_633);
or U1435 (N_1435,N_689,N_929);
nand U1436 (N_1436,N_501,N_950);
nand U1437 (N_1437,N_646,N_817);
nand U1438 (N_1438,N_949,N_551);
and U1439 (N_1439,N_519,N_564);
nand U1440 (N_1440,N_804,N_979);
nand U1441 (N_1441,N_993,N_789);
nor U1442 (N_1442,N_659,N_534);
or U1443 (N_1443,N_789,N_922);
xnor U1444 (N_1444,N_715,N_878);
and U1445 (N_1445,N_572,N_920);
or U1446 (N_1446,N_956,N_525);
nor U1447 (N_1447,N_808,N_597);
and U1448 (N_1448,N_604,N_906);
xor U1449 (N_1449,N_865,N_607);
xnor U1450 (N_1450,N_742,N_869);
nor U1451 (N_1451,N_746,N_663);
or U1452 (N_1452,N_788,N_658);
xnor U1453 (N_1453,N_720,N_584);
and U1454 (N_1454,N_735,N_844);
nor U1455 (N_1455,N_814,N_910);
or U1456 (N_1456,N_712,N_512);
or U1457 (N_1457,N_542,N_727);
and U1458 (N_1458,N_882,N_793);
nand U1459 (N_1459,N_543,N_900);
and U1460 (N_1460,N_990,N_683);
xor U1461 (N_1461,N_681,N_563);
nor U1462 (N_1462,N_700,N_679);
nor U1463 (N_1463,N_856,N_558);
nor U1464 (N_1464,N_685,N_671);
xor U1465 (N_1465,N_540,N_982);
nand U1466 (N_1466,N_790,N_956);
and U1467 (N_1467,N_958,N_893);
xnor U1468 (N_1468,N_748,N_538);
nand U1469 (N_1469,N_897,N_627);
xor U1470 (N_1470,N_555,N_816);
nand U1471 (N_1471,N_910,N_854);
or U1472 (N_1472,N_873,N_678);
xor U1473 (N_1473,N_892,N_662);
nor U1474 (N_1474,N_634,N_787);
and U1475 (N_1475,N_606,N_911);
nor U1476 (N_1476,N_729,N_594);
and U1477 (N_1477,N_757,N_577);
xnor U1478 (N_1478,N_955,N_820);
nand U1479 (N_1479,N_640,N_644);
nor U1480 (N_1480,N_995,N_611);
or U1481 (N_1481,N_586,N_724);
nand U1482 (N_1482,N_803,N_747);
xnor U1483 (N_1483,N_631,N_708);
nand U1484 (N_1484,N_569,N_595);
and U1485 (N_1485,N_616,N_734);
and U1486 (N_1486,N_942,N_695);
nand U1487 (N_1487,N_798,N_870);
nand U1488 (N_1488,N_588,N_944);
and U1489 (N_1489,N_748,N_723);
nor U1490 (N_1490,N_785,N_577);
nand U1491 (N_1491,N_671,N_799);
or U1492 (N_1492,N_576,N_570);
nand U1493 (N_1493,N_548,N_693);
nor U1494 (N_1494,N_589,N_502);
or U1495 (N_1495,N_759,N_969);
and U1496 (N_1496,N_998,N_700);
nand U1497 (N_1497,N_842,N_573);
nor U1498 (N_1498,N_583,N_539);
xnor U1499 (N_1499,N_980,N_597);
xnor U1500 (N_1500,N_1146,N_1318);
or U1501 (N_1501,N_1223,N_1492);
xor U1502 (N_1502,N_1270,N_1365);
xnor U1503 (N_1503,N_1061,N_1240);
nand U1504 (N_1504,N_1434,N_1033);
xnor U1505 (N_1505,N_1447,N_1449);
nor U1506 (N_1506,N_1302,N_1348);
and U1507 (N_1507,N_1023,N_1322);
nand U1508 (N_1508,N_1169,N_1379);
nor U1509 (N_1509,N_1339,N_1182);
xnor U1510 (N_1510,N_1350,N_1454);
xnor U1511 (N_1511,N_1151,N_1406);
xor U1512 (N_1512,N_1297,N_1370);
and U1513 (N_1513,N_1189,N_1119);
xor U1514 (N_1514,N_1135,N_1200);
nand U1515 (N_1515,N_1212,N_1368);
xnor U1516 (N_1516,N_1097,N_1430);
nor U1517 (N_1517,N_1255,N_1067);
nand U1518 (N_1518,N_1464,N_1000);
nand U1519 (N_1519,N_1310,N_1364);
xnor U1520 (N_1520,N_1329,N_1236);
nor U1521 (N_1521,N_1012,N_1170);
nand U1522 (N_1522,N_1390,N_1080);
or U1523 (N_1523,N_1109,N_1278);
nand U1524 (N_1524,N_1226,N_1056);
or U1525 (N_1525,N_1072,N_1005);
xor U1526 (N_1526,N_1399,N_1083);
and U1527 (N_1527,N_1110,N_1213);
xor U1528 (N_1528,N_1456,N_1275);
and U1529 (N_1529,N_1460,N_1301);
and U1530 (N_1530,N_1338,N_1145);
nand U1531 (N_1531,N_1076,N_1363);
and U1532 (N_1532,N_1198,N_1059);
xor U1533 (N_1533,N_1336,N_1100);
nor U1534 (N_1534,N_1139,N_1323);
and U1535 (N_1535,N_1465,N_1334);
nand U1536 (N_1536,N_1428,N_1239);
or U1537 (N_1537,N_1124,N_1105);
or U1538 (N_1538,N_1383,N_1225);
nor U1539 (N_1539,N_1332,N_1038);
nor U1540 (N_1540,N_1204,N_1260);
xor U1541 (N_1541,N_1378,N_1445);
nand U1542 (N_1542,N_1408,N_1238);
xnor U1543 (N_1543,N_1369,N_1079);
nor U1544 (N_1544,N_1263,N_1242);
and U1545 (N_1545,N_1295,N_1035);
xor U1546 (N_1546,N_1293,N_1362);
or U1547 (N_1547,N_1103,N_1398);
or U1548 (N_1548,N_1436,N_1443);
xnor U1549 (N_1549,N_1044,N_1397);
and U1550 (N_1550,N_1231,N_1307);
or U1551 (N_1551,N_1172,N_1154);
nor U1552 (N_1552,N_1114,N_1201);
and U1553 (N_1553,N_1127,N_1442);
nand U1554 (N_1554,N_1392,N_1091);
xor U1555 (N_1555,N_1459,N_1030);
or U1556 (N_1556,N_1065,N_1068);
and U1557 (N_1557,N_1308,N_1247);
or U1558 (N_1558,N_1222,N_1429);
xnor U1559 (N_1559,N_1254,N_1419);
nand U1560 (N_1560,N_1438,N_1190);
nand U1561 (N_1561,N_1498,N_1469);
xor U1562 (N_1562,N_1251,N_1249);
nor U1563 (N_1563,N_1064,N_1393);
nor U1564 (N_1564,N_1159,N_1211);
xor U1565 (N_1565,N_1279,N_1028);
nand U1566 (N_1566,N_1346,N_1437);
and U1567 (N_1567,N_1487,N_1340);
and U1568 (N_1568,N_1070,N_1253);
nor U1569 (N_1569,N_1018,N_1175);
or U1570 (N_1570,N_1243,N_1314);
nand U1571 (N_1571,N_1351,N_1384);
xnor U1572 (N_1572,N_1185,N_1401);
and U1573 (N_1573,N_1171,N_1228);
nor U1574 (N_1574,N_1244,N_1273);
nor U1575 (N_1575,N_1316,N_1111);
or U1576 (N_1576,N_1149,N_1468);
and U1577 (N_1577,N_1102,N_1446);
or U1578 (N_1578,N_1343,N_1414);
and U1579 (N_1579,N_1315,N_1161);
nor U1580 (N_1580,N_1184,N_1466);
xor U1581 (N_1581,N_1298,N_1265);
or U1582 (N_1582,N_1342,N_1326);
and U1583 (N_1583,N_1011,N_1367);
and U1584 (N_1584,N_1262,N_1413);
nor U1585 (N_1585,N_1281,N_1125);
xnor U1586 (N_1586,N_1305,N_1396);
nor U1587 (N_1587,N_1029,N_1128);
or U1588 (N_1588,N_1060,N_1163);
xor U1589 (N_1589,N_1192,N_1359);
nand U1590 (N_1590,N_1380,N_1478);
nand U1591 (N_1591,N_1054,N_1353);
xnor U1592 (N_1592,N_1021,N_1259);
xor U1593 (N_1593,N_1491,N_1188);
xor U1594 (N_1594,N_1299,N_1117);
or U1595 (N_1595,N_1294,N_1101);
nand U1596 (N_1596,N_1319,N_1328);
or U1597 (N_1597,N_1476,N_1115);
and U1598 (N_1598,N_1354,N_1164);
xnor U1599 (N_1599,N_1219,N_1327);
and U1600 (N_1600,N_1020,N_1309);
xnor U1601 (N_1601,N_1007,N_1418);
nand U1602 (N_1602,N_1410,N_1409);
nand U1603 (N_1603,N_1250,N_1395);
and U1604 (N_1604,N_1371,N_1407);
and U1605 (N_1605,N_1050,N_1321);
and U1606 (N_1606,N_1195,N_1096);
nor U1607 (N_1607,N_1349,N_1173);
xnor U1608 (N_1608,N_1152,N_1455);
and U1609 (N_1609,N_1431,N_1150);
xor U1610 (N_1610,N_1129,N_1234);
nand U1611 (N_1611,N_1156,N_1078);
xnor U1612 (N_1612,N_1218,N_1120);
or U1613 (N_1613,N_1202,N_1099);
nor U1614 (N_1614,N_1355,N_1207);
nor U1615 (N_1615,N_1009,N_1230);
or U1616 (N_1616,N_1337,N_1320);
nor U1617 (N_1617,N_1473,N_1484);
nand U1618 (N_1618,N_1043,N_1246);
nor U1619 (N_1619,N_1196,N_1074);
or U1620 (N_1620,N_1360,N_1153);
and U1621 (N_1621,N_1345,N_1062);
nor U1622 (N_1622,N_1272,N_1433);
xnor U1623 (N_1623,N_1461,N_1215);
or U1624 (N_1624,N_1095,N_1041);
and U1625 (N_1625,N_1267,N_1075);
or U1626 (N_1626,N_1168,N_1232);
nand U1627 (N_1627,N_1313,N_1143);
nand U1628 (N_1628,N_1490,N_1126);
xnor U1629 (N_1629,N_1421,N_1485);
nor U1630 (N_1630,N_1001,N_1495);
nor U1631 (N_1631,N_1214,N_1107);
nand U1632 (N_1632,N_1176,N_1049);
nand U1633 (N_1633,N_1486,N_1206);
or U1634 (N_1634,N_1417,N_1087);
or U1635 (N_1635,N_1387,N_1462);
nor U1636 (N_1636,N_1140,N_1158);
and U1637 (N_1637,N_1415,N_1084);
and U1638 (N_1638,N_1209,N_1179);
xor U1639 (N_1639,N_1098,N_1439);
or U1640 (N_1640,N_1440,N_1089);
nor U1641 (N_1641,N_1045,N_1376);
nand U1642 (N_1642,N_1463,N_1444);
nand U1643 (N_1643,N_1123,N_1481);
or U1644 (N_1644,N_1271,N_1130);
nand U1645 (N_1645,N_1121,N_1002);
and U1646 (N_1646,N_1142,N_1411);
and U1647 (N_1647,N_1488,N_1330);
nor U1648 (N_1648,N_1227,N_1136);
nand U1649 (N_1649,N_1010,N_1166);
nand U1650 (N_1650,N_1019,N_1157);
or U1651 (N_1651,N_1241,N_1248);
nor U1652 (N_1652,N_1233,N_1132);
and U1653 (N_1653,N_1147,N_1116);
nor U1654 (N_1654,N_1285,N_1208);
and U1655 (N_1655,N_1032,N_1181);
or U1656 (N_1656,N_1286,N_1258);
nand U1657 (N_1657,N_1274,N_1220);
or U1658 (N_1658,N_1288,N_1347);
or U1659 (N_1659,N_1282,N_1066);
or U1660 (N_1660,N_1221,N_1358);
nor U1661 (N_1661,N_1216,N_1494);
or U1662 (N_1662,N_1108,N_1377);
xor U1663 (N_1663,N_1134,N_1261);
xnor U1664 (N_1664,N_1489,N_1499);
xor U1665 (N_1665,N_1381,N_1324);
nor U1666 (N_1666,N_1081,N_1477);
nand U1667 (N_1667,N_1423,N_1493);
nor U1668 (N_1668,N_1372,N_1177);
xnor U1669 (N_1669,N_1194,N_1008);
and U1670 (N_1670,N_1422,N_1031);
nand U1671 (N_1671,N_1400,N_1483);
nand U1672 (N_1672,N_1266,N_1186);
and U1673 (N_1673,N_1131,N_1051);
nand U1674 (N_1674,N_1432,N_1300);
or U1675 (N_1675,N_1199,N_1069);
nor U1676 (N_1676,N_1026,N_1471);
xor U1677 (N_1677,N_1291,N_1344);
nor U1678 (N_1678,N_1312,N_1427);
nand U1679 (N_1679,N_1257,N_1224);
and U1680 (N_1680,N_1474,N_1036);
xor U1681 (N_1681,N_1458,N_1256);
or U1682 (N_1682,N_1448,N_1426);
nor U1683 (N_1683,N_1165,N_1303);
nand U1684 (N_1684,N_1388,N_1113);
nor U1685 (N_1685,N_1425,N_1148);
nor U1686 (N_1686,N_1024,N_1193);
nand U1687 (N_1687,N_1280,N_1452);
nand U1688 (N_1688,N_1073,N_1245);
and U1689 (N_1689,N_1420,N_1325);
nor U1690 (N_1690,N_1055,N_1467);
xor U1691 (N_1691,N_1450,N_1317);
or U1692 (N_1692,N_1017,N_1104);
xnor U1693 (N_1693,N_1453,N_1053);
nor U1694 (N_1694,N_1352,N_1106);
and U1695 (N_1695,N_1183,N_1482);
nor U1696 (N_1696,N_1015,N_1375);
nor U1697 (N_1697,N_1037,N_1252);
or U1698 (N_1698,N_1470,N_1394);
nand U1699 (N_1699,N_1404,N_1333);
nand U1700 (N_1700,N_1086,N_1268);
nand U1701 (N_1701,N_1144,N_1178);
nand U1702 (N_1702,N_1013,N_1237);
and U1703 (N_1703,N_1058,N_1386);
and U1704 (N_1704,N_1006,N_1361);
nor U1705 (N_1705,N_1162,N_1092);
and U1706 (N_1706,N_1269,N_1403);
or U1707 (N_1707,N_1071,N_1412);
nor U1708 (N_1708,N_1187,N_1277);
or U1709 (N_1709,N_1402,N_1122);
nor U1710 (N_1710,N_1441,N_1479);
nor U1711 (N_1711,N_1385,N_1025);
and U1712 (N_1712,N_1306,N_1382);
or U1713 (N_1713,N_1405,N_1480);
and U1714 (N_1714,N_1197,N_1210);
and U1715 (N_1715,N_1085,N_1374);
nor U1716 (N_1716,N_1203,N_1088);
nand U1717 (N_1717,N_1052,N_1496);
nor U1718 (N_1718,N_1167,N_1287);
nand U1719 (N_1719,N_1290,N_1094);
nor U1720 (N_1720,N_1497,N_1016);
and U1721 (N_1721,N_1424,N_1042);
nor U1722 (N_1722,N_1296,N_1389);
and U1723 (N_1723,N_1046,N_1451);
nand U1724 (N_1724,N_1003,N_1112);
and U1725 (N_1725,N_1160,N_1229);
or U1726 (N_1726,N_1004,N_1284);
xor U1727 (N_1727,N_1039,N_1304);
xor U1728 (N_1728,N_1435,N_1217);
nor U1729 (N_1729,N_1235,N_1174);
xor U1730 (N_1730,N_1373,N_1335);
or U1731 (N_1731,N_1048,N_1047);
nor U1732 (N_1732,N_1416,N_1063);
or U1733 (N_1733,N_1155,N_1034);
xor U1734 (N_1734,N_1093,N_1057);
or U1735 (N_1735,N_1082,N_1022);
and U1736 (N_1736,N_1118,N_1077);
nand U1737 (N_1737,N_1191,N_1331);
nor U1738 (N_1738,N_1276,N_1205);
or U1739 (N_1739,N_1311,N_1014);
and U1740 (N_1740,N_1391,N_1180);
and U1741 (N_1741,N_1138,N_1133);
nand U1742 (N_1742,N_1090,N_1357);
and U1743 (N_1743,N_1366,N_1289);
or U1744 (N_1744,N_1137,N_1264);
xnor U1745 (N_1745,N_1341,N_1292);
or U1746 (N_1746,N_1283,N_1472);
xor U1747 (N_1747,N_1141,N_1356);
and U1748 (N_1748,N_1457,N_1027);
or U1749 (N_1749,N_1040,N_1475);
nor U1750 (N_1750,N_1083,N_1061);
and U1751 (N_1751,N_1393,N_1016);
and U1752 (N_1752,N_1019,N_1290);
nand U1753 (N_1753,N_1401,N_1375);
nand U1754 (N_1754,N_1187,N_1016);
nor U1755 (N_1755,N_1368,N_1276);
nor U1756 (N_1756,N_1131,N_1299);
and U1757 (N_1757,N_1270,N_1308);
nand U1758 (N_1758,N_1458,N_1101);
nand U1759 (N_1759,N_1405,N_1469);
or U1760 (N_1760,N_1272,N_1319);
and U1761 (N_1761,N_1180,N_1331);
xor U1762 (N_1762,N_1145,N_1158);
and U1763 (N_1763,N_1363,N_1422);
xor U1764 (N_1764,N_1156,N_1424);
nand U1765 (N_1765,N_1211,N_1234);
or U1766 (N_1766,N_1207,N_1118);
and U1767 (N_1767,N_1381,N_1318);
nand U1768 (N_1768,N_1056,N_1040);
or U1769 (N_1769,N_1128,N_1099);
nand U1770 (N_1770,N_1109,N_1395);
or U1771 (N_1771,N_1395,N_1397);
nand U1772 (N_1772,N_1453,N_1454);
and U1773 (N_1773,N_1335,N_1476);
xnor U1774 (N_1774,N_1121,N_1238);
nor U1775 (N_1775,N_1270,N_1406);
nor U1776 (N_1776,N_1178,N_1085);
xor U1777 (N_1777,N_1172,N_1250);
or U1778 (N_1778,N_1087,N_1255);
or U1779 (N_1779,N_1414,N_1200);
nand U1780 (N_1780,N_1480,N_1360);
nor U1781 (N_1781,N_1424,N_1256);
nor U1782 (N_1782,N_1275,N_1214);
or U1783 (N_1783,N_1055,N_1116);
nor U1784 (N_1784,N_1436,N_1342);
and U1785 (N_1785,N_1464,N_1169);
xor U1786 (N_1786,N_1260,N_1118);
nand U1787 (N_1787,N_1093,N_1314);
or U1788 (N_1788,N_1113,N_1253);
nand U1789 (N_1789,N_1259,N_1144);
nor U1790 (N_1790,N_1440,N_1299);
xor U1791 (N_1791,N_1238,N_1347);
or U1792 (N_1792,N_1201,N_1267);
or U1793 (N_1793,N_1278,N_1448);
xor U1794 (N_1794,N_1087,N_1037);
or U1795 (N_1795,N_1258,N_1470);
xnor U1796 (N_1796,N_1125,N_1276);
xor U1797 (N_1797,N_1152,N_1420);
nor U1798 (N_1798,N_1126,N_1007);
and U1799 (N_1799,N_1385,N_1063);
and U1800 (N_1800,N_1056,N_1438);
nand U1801 (N_1801,N_1367,N_1245);
xnor U1802 (N_1802,N_1386,N_1366);
xor U1803 (N_1803,N_1028,N_1497);
xnor U1804 (N_1804,N_1260,N_1375);
nand U1805 (N_1805,N_1132,N_1172);
xnor U1806 (N_1806,N_1066,N_1083);
or U1807 (N_1807,N_1130,N_1080);
and U1808 (N_1808,N_1417,N_1487);
nor U1809 (N_1809,N_1344,N_1262);
nand U1810 (N_1810,N_1348,N_1093);
and U1811 (N_1811,N_1023,N_1421);
or U1812 (N_1812,N_1151,N_1309);
nand U1813 (N_1813,N_1061,N_1495);
nor U1814 (N_1814,N_1056,N_1433);
nand U1815 (N_1815,N_1180,N_1491);
nor U1816 (N_1816,N_1077,N_1064);
xor U1817 (N_1817,N_1165,N_1193);
or U1818 (N_1818,N_1289,N_1433);
nor U1819 (N_1819,N_1274,N_1130);
or U1820 (N_1820,N_1341,N_1040);
and U1821 (N_1821,N_1287,N_1241);
and U1822 (N_1822,N_1304,N_1025);
nor U1823 (N_1823,N_1230,N_1382);
nand U1824 (N_1824,N_1474,N_1131);
or U1825 (N_1825,N_1292,N_1484);
nor U1826 (N_1826,N_1300,N_1372);
or U1827 (N_1827,N_1037,N_1001);
or U1828 (N_1828,N_1433,N_1463);
or U1829 (N_1829,N_1011,N_1065);
or U1830 (N_1830,N_1160,N_1062);
xor U1831 (N_1831,N_1152,N_1136);
nor U1832 (N_1832,N_1498,N_1079);
xnor U1833 (N_1833,N_1159,N_1361);
nor U1834 (N_1834,N_1124,N_1238);
xor U1835 (N_1835,N_1172,N_1159);
nor U1836 (N_1836,N_1023,N_1287);
nor U1837 (N_1837,N_1308,N_1307);
nand U1838 (N_1838,N_1112,N_1021);
nand U1839 (N_1839,N_1095,N_1063);
xor U1840 (N_1840,N_1366,N_1314);
or U1841 (N_1841,N_1035,N_1280);
nand U1842 (N_1842,N_1183,N_1375);
nor U1843 (N_1843,N_1326,N_1189);
nand U1844 (N_1844,N_1307,N_1114);
and U1845 (N_1845,N_1369,N_1104);
xor U1846 (N_1846,N_1415,N_1316);
or U1847 (N_1847,N_1279,N_1445);
xnor U1848 (N_1848,N_1383,N_1389);
xnor U1849 (N_1849,N_1486,N_1414);
xor U1850 (N_1850,N_1131,N_1470);
nor U1851 (N_1851,N_1470,N_1390);
nand U1852 (N_1852,N_1077,N_1065);
nand U1853 (N_1853,N_1363,N_1003);
and U1854 (N_1854,N_1223,N_1273);
xnor U1855 (N_1855,N_1355,N_1131);
or U1856 (N_1856,N_1393,N_1102);
and U1857 (N_1857,N_1364,N_1323);
nand U1858 (N_1858,N_1496,N_1388);
or U1859 (N_1859,N_1026,N_1426);
and U1860 (N_1860,N_1061,N_1102);
or U1861 (N_1861,N_1000,N_1348);
or U1862 (N_1862,N_1344,N_1042);
nand U1863 (N_1863,N_1435,N_1461);
and U1864 (N_1864,N_1219,N_1063);
nand U1865 (N_1865,N_1494,N_1306);
nand U1866 (N_1866,N_1441,N_1235);
or U1867 (N_1867,N_1141,N_1338);
nor U1868 (N_1868,N_1184,N_1482);
or U1869 (N_1869,N_1085,N_1032);
nor U1870 (N_1870,N_1238,N_1119);
and U1871 (N_1871,N_1412,N_1472);
or U1872 (N_1872,N_1324,N_1479);
and U1873 (N_1873,N_1356,N_1437);
or U1874 (N_1874,N_1464,N_1285);
xnor U1875 (N_1875,N_1060,N_1492);
xnor U1876 (N_1876,N_1048,N_1198);
xnor U1877 (N_1877,N_1331,N_1099);
or U1878 (N_1878,N_1259,N_1148);
and U1879 (N_1879,N_1325,N_1201);
or U1880 (N_1880,N_1070,N_1322);
and U1881 (N_1881,N_1209,N_1311);
or U1882 (N_1882,N_1420,N_1051);
and U1883 (N_1883,N_1171,N_1243);
or U1884 (N_1884,N_1335,N_1166);
nand U1885 (N_1885,N_1334,N_1238);
xor U1886 (N_1886,N_1256,N_1161);
xor U1887 (N_1887,N_1468,N_1369);
nor U1888 (N_1888,N_1458,N_1492);
nand U1889 (N_1889,N_1423,N_1158);
nand U1890 (N_1890,N_1084,N_1429);
xnor U1891 (N_1891,N_1445,N_1267);
xnor U1892 (N_1892,N_1229,N_1100);
nor U1893 (N_1893,N_1477,N_1168);
xnor U1894 (N_1894,N_1454,N_1326);
nand U1895 (N_1895,N_1069,N_1433);
and U1896 (N_1896,N_1047,N_1478);
and U1897 (N_1897,N_1472,N_1333);
and U1898 (N_1898,N_1356,N_1029);
nand U1899 (N_1899,N_1070,N_1309);
or U1900 (N_1900,N_1476,N_1394);
nor U1901 (N_1901,N_1385,N_1321);
nor U1902 (N_1902,N_1366,N_1212);
and U1903 (N_1903,N_1100,N_1303);
nor U1904 (N_1904,N_1100,N_1111);
or U1905 (N_1905,N_1460,N_1386);
xor U1906 (N_1906,N_1174,N_1440);
nor U1907 (N_1907,N_1393,N_1291);
xnor U1908 (N_1908,N_1289,N_1399);
or U1909 (N_1909,N_1433,N_1246);
or U1910 (N_1910,N_1199,N_1218);
nor U1911 (N_1911,N_1190,N_1065);
nand U1912 (N_1912,N_1221,N_1160);
or U1913 (N_1913,N_1085,N_1218);
or U1914 (N_1914,N_1092,N_1307);
nand U1915 (N_1915,N_1139,N_1121);
xnor U1916 (N_1916,N_1379,N_1263);
nor U1917 (N_1917,N_1338,N_1144);
or U1918 (N_1918,N_1323,N_1051);
nor U1919 (N_1919,N_1035,N_1141);
or U1920 (N_1920,N_1164,N_1465);
nor U1921 (N_1921,N_1412,N_1320);
nand U1922 (N_1922,N_1354,N_1453);
nor U1923 (N_1923,N_1173,N_1032);
nor U1924 (N_1924,N_1049,N_1218);
nor U1925 (N_1925,N_1158,N_1029);
nor U1926 (N_1926,N_1222,N_1098);
nand U1927 (N_1927,N_1210,N_1134);
or U1928 (N_1928,N_1144,N_1475);
and U1929 (N_1929,N_1483,N_1114);
nor U1930 (N_1930,N_1058,N_1265);
or U1931 (N_1931,N_1288,N_1359);
nand U1932 (N_1932,N_1432,N_1372);
nand U1933 (N_1933,N_1227,N_1492);
nor U1934 (N_1934,N_1078,N_1084);
nand U1935 (N_1935,N_1063,N_1105);
nor U1936 (N_1936,N_1005,N_1487);
xnor U1937 (N_1937,N_1061,N_1108);
xnor U1938 (N_1938,N_1065,N_1231);
and U1939 (N_1939,N_1183,N_1472);
nand U1940 (N_1940,N_1460,N_1359);
nand U1941 (N_1941,N_1053,N_1178);
and U1942 (N_1942,N_1337,N_1089);
or U1943 (N_1943,N_1433,N_1450);
or U1944 (N_1944,N_1334,N_1004);
or U1945 (N_1945,N_1387,N_1408);
or U1946 (N_1946,N_1074,N_1235);
or U1947 (N_1947,N_1067,N_1381);
xor U1948 (N_1948,N_1120,N_1305);
or U1949 (N_1949,N_1178,N_1243);
or U1950 (N_1950,N_1462,N_1421);
or U1951 (N_1951,N_1111,N_1337);
or U1952 (N_1952,N_1435,N_1436);
xnor U1953 (N_1953,N_1007,N_1383);
nand U1954 (N_1954,N_1381,N_1422);
nor U1955 (N_1955,N_1459,N_1165);
xnor U1956 (N_1956,N_1261,N_1233);
or U1957 (N_1957,N_1189,N_1031);
xor U1958 (N_1958,N_1185,N_1177);
nand U1959 (N_1959,N_1352,N_1455);
xnor U1960 (N_1960,N_1367,N_1377);
and U1961 (N_1961,N_1468,N_1020);
nor U1962 (N_1962,N_1177,N_1349);
and U1963 (N_1963,N_1101,N_1274);
or U1964 (N_1964,N_1404,N_1366);
nor U1965 (N_1965,N_1082,N_1498);
and U1966 (N_1966,N_1449,N_1072);
and U1967 (N_1967,N_1248,N_1239);
xnor U1968 (N_1968,N_1170,N_1146);
or U1969 (N_1969,N_1436,N_1367);
nand U1970 (N_1970,N_1353,N_1119);
nand U1971 (N_1971,N_1177,N_1407);
xor U1972 (N_1972,N_1255,N_1476);
and U1973 (N_1973,N_1011,N_1329);
nor U1974 (N_1974,N_1126,N_1463);
or U1975 (N_1975,N_1492,N_1463);
nand U1976 (N_1976,N_1335,N_1079);
nand U1977 (N_1977,N_1114,N_1306);
and U1978 (N_1978,N_1298,N_1000);
nor U1979 (N_1979,N_1012,N_1162);
and U1980 (N_1980,N_1005,N_1389);
or U1981 (N_1981,N_1462,N_1145);
xor U1982 (N_1982,N_1057,N_1334);
xnor U1983 (N_1983,N_1487,N_1364);
xnor U1984 (N_1984,N_1161,N_1117);
or U1985 (N_1985,N_1382,N_1056);
nand U1986 (N_1986,N_1170,N_1108);
nand U1987 (N_1987,N_1047,N_1458);
nor U1988 (N_1988,N_1497,N_1157);
and U1989 (N_1989,N_1180,N_1313);
nor U1990 (N_1990,N_1463,N_1238);
nand U1991 (N_1991,N_1426,N_1437);
nand U1992 (N_1992,N_1209,N_1234);
or U1993 (N_1993,N_1079,N_1202);
nand U1994 (N_1994,N_1356,N_1371);
or U1995 (N_1995,N_1437,N_1130);
xor U1996 (N_1996,N_1455,N_1171);
or U1997 (N_1997,N_1257,N_1108);
or U1998 (N_1998,N_1337,N_1021);
and U1999 (N_1999,N_1412,N_1138);
nor U2000 (N_2000,N_1595,N_1887);
or U2001 (N_2001,N_1825,N_1789);
and U2002 (N_2002,N_1662,N_1728);
nor U2003 (N_2003,N_1550,N_1831);
nand U2004 (N_2004,N_1650,N_1960);
nand U2005 (N_2005,N_1577,N_1882);
nand U2006 (N_2006,N_1833,N_1516);
xnor U2007 (N_2007,N_1747,N_1954);
nand U2008 (N_2008,N_1676,N_1795);
xnor U2009 (N_2009,N_1708,N_1537);
or U2010 (N_2010,N_1930,N_1699);
nor U2011 (N_2011,N_1718,N_1838);
or U2012 (N_2012,N_1917,N_1692);
xor U2013 (N_2013,N_1848,N_1780);
xor U2014 (N_2014,N_1846,N_1619);
nand U2015 (N_2015,N_1757,N_1693);
nor U2016 (N_2016,N_1736,N_1568);
and U2017 (N_2017,N_1652,N_1905);
xnor U2018 (N_2018,N_1647,N_1709);
xor U2019 (N_2019,N_1916,N_1868);
nor U2020 (N_2020,N_1984,N_1983);
and U2021 (N_2021,N_1994,N_1678);
nand U2022 (N_2022,N_1814,N_1573);
and U2023 (N_2023,N_1951,N_1963);
xnor U2024 (N_2024,N_1752,N_1853);
or U2025 (N_2025,N_1844,N_1779);
nor U2026 (N_2026,N_1601,N_1575);
nor U2027 (N_2027,N_1944,N_1523);
or U2028 (N_2028,N_1989,N_1937);
xnor U2029 (N_2029,N_1631,N_1566);
nand U2030 (N_2030,N_1915,N_1941);
xnor U2031 (N_2031,N_1929,N_1875);
and U2032 (N_2032,N_1743,N_1547);
or U2033 (N_2033,N_1739,N_1758);
nor U2034 (N_2034,N_1856,N_1645);
xor U2035 (N_2035,N_1998,N_1629);
and U2036 (N_2036,N_1742,N_1925);
or U2037 (N_2037,N_1644,N_1809);
or U2038 (N_2038,N_1892,N_1976);
nor U2039 (N_2039,N_1625,N_1580);
and U2040 (N_2040,N_1682,N_1528);
or U2041 (N_2041,N_1689,N_1636);
nand U2042 (N_2042,N_1893,N_1648);
or U2043 (N_2043,N_1910,N_1584);
nand U2044 (N_2044,N_1734,N_1922);
or U2045 (N_2045,N_1594,N_1906);
xnor U2046 (N_2046,N_1518,N_1506);
xor U2047 (N_2047,N_1847,N_1791);
xnor U2048 (N_2048,N_1936,N_1700);
nand U2049 (N_2049,N_1766,N_1507);
nor U2050 (N_2050,N_1872,N_1551);
and U2051 (N_2051,N_1562,N_1978);
or U2052 (N_2052,N_1615,N_1639);
nor U2053 (N_2053,N_1790,N_1681);
or U2054 (N_2054,N_1590,N_1545);
or U2055 (N_2055,N_1637,N_1656);
or U2056 (N_2056,N_1874,N_1815);
and U2057 (N_2057,N_1927,N_1958);
and U2058 (N_2058,N_1920,N_1955);
xor U2059 (N_2059,N_1841,N_1623);
nand U2060 (N_2060,N_1852,N_1604);
nand U2061 (N_2061,N_1582,N_1654);
nand U2062 (N_2062,N_1785,N_1860);
or U2063 (N_2063,N_1710,N_1953);
and U2064 (N_2064,N_1737,N_1962);
nand U2065 (N_2065,N_1712,N_1756);
and U2066 (N_2066,N_1850,N_1839);
xor U2067 (N_2067,N_1898,N_1793);
nor U2068 (N_2068,N_1711,N_1957);
nand U2069 (N_2069,N_1628,N_1968);
or U2070 (N_2070,N_1558,N_1769);
or U2071 (N_2071,N_1612,N_1884);
xor U2072 (N_2072,N_1928,N_1515);
nand U2073 (N_2073,N_1913,N_1867);
or U2074 (N_2074,N_1603,N_1986);
nand U2075 (N_2075,N_1830,N_1542);
nor U2076 (N_2076,N_1688,N_1741);
xnor U2077 (N_2077,N_1776,N_1886);
nand U2078 (N_2078,N_1521,N_1883);
and U2079 (N_2079,N_1914,N_1724);
xor U2080 (N_2080,N_1630,N_1540);
nand U2081 (N_2081,N_1826,N_1849);
or U2082 (N_2082,N_1671,N_1526);
nand U2083 (N_2083,N_1613,N_1750);
nand U2084 (N_2084,N_1821,N_1802);
or U2085 (N_2085,N_1767,N_1903);
nor U2086 (N_2086,N_1858,N_1987);
xnor U2087 (N_2087,N_1836,N_1744);
xnor U2088 (N_2088,N_1806,N_1500);
nor U2089 (N_2089,N_1855,N_1900);
nor U2090 (N_2090,N_1672,N_1851);
or U2091 (N_2091,N_1857,N_1591);
and U2092 (N_2092,N_1798,N_1866);
xnor U2093 (N_2093,N_1843,N_1588);
or U2094 (N_2094,N_1907,N_1745);
xor U2095 (N_2095,N_1771,N_1760);
xnor U2096 (N_2096,N_1599,N_1570);
nor U2097 (N_2097,N_1690,N_1985);
nor U2098 (N_2098,N_1530,N_1885);
xor U2099 (N_2099,N_1977,N_1950);
and U2100 (N_2100,N_1513,N_1723);
nor U2101 (N_2101,N_1923,N_1670);
xnor U2102 (N_2102,N_1800,N_1902);
nor U2103 (N_2103,N_1572,N_1942);
xnor U2104 (N_2104,N_1979,N_1541);
nor U2105 (N_2105,N_1813,N_1600);
nor U2106 (N_2106,N_1564,N_1641);
xnor U2107 (N_2107,N_1634,N_1948);
nand U2108 (N_2108,N_1891,N_1719);
xnor U2109 (N_2109,N_1730,N_1921);
nand U2110 (N_2110,N_1546,N_1722);
nand U2111 (N_2111,N_1609,N_1655);
and U2112 (N_2112,N_1565,N_1538);
nand U2113 (N_2113,N_1919,N_1759);
xor U2114 (N_2114,N_1549,N_1614);
nor U2115 (N_2115,N_1598,N_1765);
nor U2116 (N_2116,N_1904,N_1947);
nand U2117 (N_2117,N_1535,N_1763);
or U2118 (N_2118,N_1651,N_1996);
nor U2119 (N_2119,N_1553,N_1640);
and U2120 (N_2120,N_1864,N_1532);
and U2121 (N_2121,N_1597,N_1799);
xnor U2122 (N_2122,N_1773,N_1658);
or U2123 (N_2123,N_1512,N_1509);
and U2124 (N_2124,N_1794,N_1683);
nand U2125 (N_2125,N_1596,N_1627);
and U2126 (N_2126,N_1714,N_1881);
and U2127 (N_2127,N_1684,N_1787);
nor U2128 (N_2128,N_1859,N_1797);
nor U2129 (N_2129,N_1696,N_1725);
nor U2130 (N_2130,N_1901,N_1946);
and U2131 (N_2131,N_1783,N_1805);
and U2132 (N_2132,N_1520,N_1973);
xnor U2133 (N_2133,N_1819,N_1698);
xnor U2134 (N_2134,N_1967,N_1876);
or U2135 (N_2135,N_1735,N_1931);
and U2136 (N_2136,N_1691,N_1810);
nor U2137 (N_2137,N_1685,N_1531);
xnor U2138 (N_2138,N_1638,N_1897);
and U2139 (N_2139,N_1707,N_1510);
nor U2140 (N_2140,N_1552,N_1686);
nand U2141 (N_2141,N_1772,N_1704);
and U2142 (N_2142,N_1620,N_1863);
nor U2143 (N_2143,N_1560,N_1827);
xnor U2144 (N_2144,N_1585,N_1563);
and U2145 (N_2145,N_1519,N_1932);
nand U2146 (N_2146,N_1543,N_1961);
xor U2147 (N_2147,N_1861,N_1889);
xnor U2148 (N_2148,N_1992,N_1877);
xor U2149 (N_2149,N_1970,N_1823);
xnor U2150 (N_2150,N_1605,N_1751);
or U2151 (N_2151,N_1569,N_1869);
nand U2152 (N_2152,N_1788,N_1999);
nor U2153 (N_2153,N_1695,N_1926);
nor U2154 (N_2154,N_1895,N_1908);
and U2155 (N_2155,N_1720,N_1778);
or U2156 (N_2156,N_1971,N_1626);
nand U2157 (N_2157,N_1643,N_1754);
xnor U2158 (N_2158,N_1804,N_1517);
or U2159 (N_2159,N_1924,N_1764);
or U2160 (N_2160,N_1862,N_1982);
nor U2161 (N_2161,N_1845,N_1525);
and U2162 (N_2162,N_1738,N_1579);
nor U2163 (N_2163,N_1716,N_1934);
or U2164 (N_2164,N_1508,N_1624);
or U2165 (N_2165,N_1871,N_1705);
and U2166 (N_2166,N_1988,N_1997);
nor U2167 (N_2167,N_1956,N_1571);
xor U2168 (N_2168,N_1781,N_1661);
and U2169 (N_2169,N_1608,N_1659);
or U2170 (N_2170,N_1824,N_1808);
or U2171 (N_2171,N_1803,N_1890);
and U2172 (N_2172,N_1701,N_1975);
nand U2173 (N_2173,N_1583,N_1873);
nor U2174 (N_2174,N_1727,N_1938);
xor U2175 (N_2175,N_1820,N_1837);
nor U2176 (N_2176,N_1811,N_1786);
or U2177 (N_2177,N_1993,N_1679);
nor U2178 (N_2178,N_1753,N_1567);
or U2179 (N_2179,N_1835,N_1829);
or U2180 (N_2180,N_1574,N_1592);
xnor U2181 (N_2181,N_1784,N_1677);
nand U2182 (N_2182,N_1616,N_1607);
nand U2183 (N_2183,N_1879,N_1680);
or U2184 (N_2184,N_1807,N_1702);
nand U2185 (N_2185,N_1918,N_1965);
and U2186 (N_2186,N_1694,N_1602);
nand U2187 (N_2187,N_1943,N_1717);
nand U2188 (N_2188,N_1557,N_1697);
and U2189 (N_2189,N_1854,N_1669);
nand U2190 (N_2190,N_1586,N_1980);
xor U2191 (N_2191,N_1770,N_1896);
and U2192 (N_2192,N_1834,N_1816);
and U2193 (N_2193,N_1878,N_1649);
or U2194 (N_2194,N_1664,N_1715);
nor U2195 (N_2195,N_1840,N_1865);
nand U2196 (N_2196,N_1646,N_1991);
nor U2197 (N_2197,N_1660,N_1653);
nand U2198 (N_2198,N_1524,N_1974);
xor U2199 (N_2199,N_1894,N_1606);
and U2200 (N_2200,N_1939,N_1502);
or U2201 (N_2201,N_1768,N_1534);
xor U2202 (N_2202,N_1576,N_1733);
nand U2203 (N_2203,N_1935,N_1899);
xnor U2204 (N_2204,N_1674,N_1633);
and U2205 (N_2205,N_1611,N_1663);
nor U2206 (N_2206,N_1972,N_1587);
or U2207 (N_2207,N_1703,N_1792);
xor U2208 (N_2208,N_1959,N_1777);
xnor U2209 (N_2209,N_1667,N_1561);
or U2210 (N_2210,N_1675,N_1774);
xnor U2211 (N_2211,N_1801,N_1746);
or U2212 (N_2212,N_1912,N_1589);
nand U2213 (N_2213,N_1945,N_1969);
or U2214 (N_2214,N_1556,N_1832);
xor U2215 (N_2215,N_1514,N_1617);
nor U2216 (N_2216,N_1729,N_1817);
nand U2217 (N_2217,N_1559,N_1755);
xnor U2218 (N_2218,N_1642,N_1501);
and U2219 (N_2219,N_1503,N_1544);
nor U2220 (N_2220,N_1673,N_1726);
and U2221 (N_2221,N_1554,N_1536);
or U2222 (N_2222,N_1933,N_1504);
nor U2223 (N_2223,N_1529,N_1966);
and U2224 (N_2224,N_1668,N_1995);
nor U2225 (N_2225,N_1539,N_1911);
and U2226 (N_2226,N_1610,N_1578);
nand U2227 (N_2227,N_1748,N_1749);
nand U2228 (N_2228,N_1622,N_1740);
or U2229 (N_2229,N_1687,N_1666);
nor U2230 (N_2230,N_1909,N_1761);
and U2231 (N_2231,N_1618,N_1990);
nor U2232 (N_2232,N_1796,N_1940);
or U2233 (N_2233,N_1949,N_1593);
nor U2234 (N_2234,N_1964,N_1635);
or U2235 (N_2235,N_1818,N_1822);
or U2236 (N_2236,N_1713,N_1665);
and U2237 (N_2237,N_1548,N_1828);
and U2238 (N_2238,N_1533,N_1888);
nand U2239 (N_2239,N_1657,N_1706);
nand U2240 (N_2240,N_1782,N_1812);
and U2241 (N_2241,N_1775,N_1731);
xor U2242 (N_2242,N_1505,N_1511);
xor U2243 (N_2243,N_1762,N_1555);
xnor U2244 (N_2244,N_1870,N_1981);
nand U2245 (N_2245,N_1721,N_1880);
and U2246 (N_2246,N_1842,N_1632);
nor U2247 (N_2247,N_1732,N_1621);
nor U2248 (N_2248,N_1581,N_1527);
nor U2249 (N_2249,N_1522,N_1952);
or U2250 (N_2250,N_1653,N_1993);
or U2251 (N_2251,N_1779,N_1699);
nor U2252 (N_2252,N_1713,N_1884);
nor U2253 (N_2253,N_1682,N_1985);
or U2254 (N_2254,N_1624,N_1696);
xor U2255 (N_2255,N_1599,N_1976);
and U2256 (N_2256,N_1811,N_1955);
xor U2257 (N_2257,N_1866,N_1734);
or U2258 (N_2258,N_1543,N_1835);
and U2259 (N_2259,N_1672,N_1670);
nand U2260 (N_2260,N_1506,N_1992);
or U2261 (N_2261,N_1650,N_1599);
nand U2262 (N_2262,N_1831,N_1876);
nand U2263 (N_2263,N_1813,N_1677);
xnor U2264 (N_2264,N_1916,N_1908);
and U2265 (N_2265,N_1779,N_1971);
or U2266 (N_2266,N_1576,N_1561);
xnor U2267 (N_2267,N_1697,N_1768);
nor U2268 (N_2268,N_1780,N_1806);
nor U2269 (N_2269,N_1541,N_1911);
nor U2270 (N_2270,N_1647,N_1553);
nand U2271 (N_2271,N_1537,N_1676);
or U2272 (N_2272,N_1952,N_1987);
or U2273 (N_2273,N_1758,N_1842);
and U2274 (N_2274,N_1623,N_1521);
or U2275 (N_2275,N_1953,N_1544);
nor U2276 (N_2276,N_1944,N_1909);
nor U2277 (N_2277,N_1675,N_1695);
nor U2278 (N_2278,N_1862,N_1952);
nor U2279 (N_2279,N_1850,N_1506);
nor U2280 (N_2280,N_1519,N_1891);
nand U2281 (N_2281,N_1629,N_1785);
or U2282 (N_2282,N_1906,N_1587);
nor U2283 (N_2283,N_1890,N_1513);
nand U2284 (N_2284,N_1641,N_1923);
or U2285 (N_2285,N_1800,N_1562);
nand U2286 (N_2286,N_1882,N_1744);
or U2287 (N_2287,N_1696,N_1656);
and U2288 (N_2288,N_1504,N_1809);
and U2289 (N_2289,N_1667,N_1947);
nand U2290 (N_2290,N_1806,N_1817);
and U2291 (N_2291,N_1972,N_1803);
nor U2292 (N_2292,N_1727,N_1920);
nor U2293 (N_2293,N_1515,N_1978);
or U2294 (N_2294,N_1739,N_1983);
or U2295 (N_2295,N_1998,N_1573);
or U2296 (N_2296,N_1933,N_1935);
nand U2297 (N_2297,N_1997,N_1537);
or U2298 (N_2298,N_1694,N_1991);
xnor U2299 (N_2299,N_1869,N_1913);
and U2300 (N_2300,N_1967,N_1951);
nor U2301 (N_2301,N_1645,N_1646);
xnor U2302 (N_2302,N_1997,N_1966);
nor U2303 (N_2303,N_1526,N_1550);
or U2304 (N_2304,N_1943,N_1813);
xnor U2305 (N_2305,N_1762,N_1926);
and U2306 (N_2306,N_1769,N_1672);
xnor U2307 (N_2307,N_1568,N_1795);
or U2308 (N_2308,N_1802,N_1622);
or U2309 (N_2309,N_1797,N_1959);
or U2310 (N_2310,N_1587,N_1752);
or U2311 (N_2311,N_1844,N_1958);
or U2312 (N_2312,N_1944,N_1772);
xor U2313 (N_2313,N_1855,N_1931);
nor U2314 (N_2314,N_1759,N_1570);
nand U2315 (N_2315,N_1956,N_1938);
xor U2316 (N_2316,N_1684,N_1954);
or U2317 (N_2317,N_1543,N_1827);
nand U2318 (N_2318,N_1625,N_1765);
and U2319 (N_2319,N_1932,N_1610);
and U2320 (N_2320,N_1975,N_1948);
nor U2321 (N_2321,N_1973,N_1766);
or U2322 (N_2322,N_1500,N_1870);
nand U2323 (N_2323,N_1667,N_1624);
nor U2324 (N_2324,N_1820,N_1629);
and U2325 (N_2325,N_1620,N_1802);
and U2326 (N_2326,N_1563,N_1661);
xnor U2327 (N_2327,N_1914,N_1800);
xnor U2328 (N_2328,N_1763,N_1816);
or U2329 (N_2329,N_1626,N_1897);
and U2330 (N_2330,N_1818,N_1621);
nor U2331 (N_2331,N_1510,N_1598);
nor U2332 (N_2332,N_1570,N_1832);
nor U2333 (N_2333,N_1942,N_1796);
nor U2334 (N_2334,N_1719,N_1517);
nor U2335 (N_2335,N_1704,N_1942);
nand U2336 (N_2336,N_1777,N_1559);
xnor U2337 (N_2337,N_1548,N_1573);
nand U2338 (N_2338,N_1612,N_1786);
nand U2339 (N_2339,N_1924,N_1564);
nor U2340 (N_2340,N_1952,N_1711);
or U2341 (N_2341,N_1968,N_1509);
xnor U2342 (N_2342,N_1971,N_1802);
or U2343 (N_2343,N_1664,N_1542);
and U2344 (N_2344,N_1532,N_1992);
and U2345 (N_2345,N_1757,N_1638);
or U2346 (N_2346,N_1662,N_1625);
nor U2347 (N_2347,N_1983,N_1621);
xnor U2348 (N_2348,N_1999,N_1939);
or U2349 (N_2349,N_1893,N_1779);
nand U2350 (N_2350,N_1527,N_1621);
nor U2351 (N_2351,N_1674,N_1993);
nor U2352 (N_2352,N_1790,N_1657);
or U2353 (N_2353,N_1764,N_1742);
nand U2354 (N_2354,N_1517,N_1826);
nor U2355 (N_2355,N_1866,N_1991);
xnor U2356 (N_2356,N_1847,N_1577);
and U2357 (N_2357,N_1947,N_1641);
nor U2358 (N_2358,N_1788,N_1907);
or U2359 (N_2359,N_1548,N_1836);
or U2360 (N_2360,N_1663,N_1669);
nand U2361 (N_2361,N_1893,N_1671);
nand U2362 (N_2362,N_1523,N_1850);
and U2363 (N_2363,N_1642,N_1832);
nor U2364 (N_2364,N_1559,N_1696);
nor U2365 (N_2365,N_1942,N_1843);
and U2366 (N_2366,N_1916,N_1733);
or U2367 (N_2367,N_1555,N_1564);
xnor U2368 (N_2368,N_1748,N_1889);
xnor U2369 (N_2369,N_1693,N_1852);
nor U2370 (N_2370,N_1861,N_1788);
nand U2371 (N_2371,N_1779,N_1767);
and U2372 (N_2372,N_1897,N_1919);
or U2373 (N_2373,N_1776,N_1517);
or U2374 (N_2374,N_1838,N_1557);
nor U2375 (N_2375,N_1933,N_1641);
xnor U2376 (N_2376,N_1992,N_1980);
nand U2377 (N_2377,N_1554,N_1742);
and U2378 (N_2378,N_1572,N_1654);
and U2379 (N_2379,N_1595,N_1809);
and U2380 (N_2380,N_1794,N_1785);
nand U2381 (N_2381,N_1798,N_1882);
nand U2382 (N_2382,N_1563,N_1747);
nand U2383 (N_2383,N_1892,N_1816);
nand U2384 (N_2384,N_1941,N_1897);
or U2385 (N_2385,N_1663,N_1659);
or U2386 (N_2386,N_1852,N_1979);
nand U2387 (N_2387,N_1933,N_1580);
and U2388 (N_2388,N_1966,N_1538);
nand U2389 (N_2389,N_1576,N_1535);
nor U2390 (N_2390,N_1501,N_1609);
nor U2391 (N_2391,N_1551,N_1922);
or U2392 (N_2392,N_1859,N_1769);
and U2393 (N_2393,N_1981,N_1992);
or U2394 (N_2394,N_1918,N_1805);
and U2395 (N_2395,N_1668,N_1824);
and U2396 (N_2396,N_1593,N_1578);
nand U2397 (N_2397,N_1915,N_1817);
xor U2398 (N_2398,N_1997,N_1913);
or U2399 (N_2399,N_1857,N_1850);
or U2400 (N_2400,N_1726,N_1769);
nand U2401 (N_2401,N_1829,N_1740);
or U2402 (N_2402,N_1741,N_1586);
nor U2403 (N_2403,N_1732,N_1551);
xor U2404 (N_2404,N_1700,N_1975);
and U2405 (N_2405,N_1946,N_1598);
or U2406 (N_2406,N_1805,N_1868);
or U2407 (N_2407,N_1688,N_1865);
nor U2408 (N_2408,N_1601,N_1559);
and U2409 (N_2409,N_1510,N_1718);
nor U2410 (N_2410,N_1692,N_1542);
xor U2411 (N_2411,N_1926,N_1538);
or U2412 (N_2412,N_1652,N_1805);
nand U2413 (N_2413,N_1871,N_1994);
and U2414 (N_2414,N_1603,N_1840);
and U2415 (N_2415,N_1944,N_1819);
nor U2416 (N_2416,N_1580,N_1844);
nor U2417 (N_2417,N_1773,N_1825);
or U2418 (N_2418,N_1597,N_1603);
xor U2419 (N_2419,N_1719,N_1536);
and U2420 (N_2420,N_1729,N_1866);
and U2421 (N_2421,N_1759,N_1658);
xor U2422 (N_2422,N_1514,N_1633);
and U2423 (N_2423,N_1810,N_1773);
or U2424 (N_2424,N_1553,N_1597);
and U2425 (N_2425,N_1697,N_1795);
and U2426 (N_2426,N_1515,N_1607);
nor U2427 (N_2427,N_1638,N_1818);
nand U2428 (N_2428,N_1765,N_1718);
xnor U2429 (N_2429,N_1930,N_1516);
nand U2430 (N_2430,N_1586,N_1951);
and U2431 (N_2431,N_1607,N_1728);
xor U2432 (N_2432,N_1884,N_1569);
xnor U2433 (N_2433,N_1957,N_1760);
and U2434 (N_2434,N_1858,N_1935);
nand U2435 (N_2435,N_1811,N_1736);
xnor U2436 (N_2436,N_1711,N_1599);
or U2437 (N_2437,N_1700,N_1659);
nand U2438 (N_2438,N_1724,N_1768);
or U2439 (N_2439,N_1537,N_1801);
nand U2440 (N_2440,N_1781,N_1852);
or U2441 (N_2441,N_1655,N_1856);
xnor U2442 (N_2442,N_1812,N_1821);
nor U2443 (N_2443,N_1900,N_1839);
or U2444 (N_2444,N_1761,N_1911);
and U2445 (N_2445,N_1903,N_1907);
nor U2446 (N_2446,N_1995,N_1778);
and U2447 (N_2447,N_1591,N_1929);
nand U2448 (N_2448,N_1695,N_1706);
nand U2449 (N_2449,N_1554,N_1839);
or U2450 (N_2450,N_1848,N_1978);
nor U2451 (N_2451,N_1680,N_1631);
nor U2452 (N_2452,N_1754,N_1881);
nand U2453 (N_2453,N_1561,N_1725);
and U2454 (N_2454,N_1630,N_1662);
or U2455 (N_2455,N_1688,N_1820);
or U2456 (N_2456,N_1840,N_1810);
nand U2457 (N_2457,N_1806,N_1917);
xor U2458 (N_2458,N_1568,N_1657);
nor U2459 (N_2459,N_1987,N_1726);
and U2460 (N_2460,N_1917,N_1951);
xnor U2461 (N_2461,N_1523,N_1655);
nor U2462 (N_2462,N_1618,N_1668);
or U2463 (N_2463,N_1625,N_1756);
nand U2464 (N_2464,N_1651,N_1860);
xor U2465 (N_2465,N_1843,N_1817);
or U2466 (N_2466,N_1848,N_1724);
xor U2467 (N_2467,N_1699,N_1756);
nand U2468 (N_2468,N_1978,N_1977);
or U2469 (N_2469,N_1542,N_1555);
and U2470 (N_2470,N_1709,N_1524);
nand U2471 (N_2471,N_1755,N_1642);
or U2472 (N_2472,N_1988,N_1736);
nand U2473 (N_2473,N_1797,N_1895);
and U2474 (N_2474,N_1818,N_1887);
or U2475 (N_2475,N_1853,N_1590);
and U2476 (N_2476,N_1820,N_1720);
nand U2477 (N_2477,N_1769,N_1562);
nand U2478 (N_2478,N_1768,N_1566);
nand U2479 (N_2479,N_1821,N_1720);
and U2480 (N_2480,N_1647,N_1990);
and U2481 (N_2481,N_1962,N_1614);
or U2482 (N_2482,N_1921,N_1528);
nand U2483 (N_2483,N_1701,N_1526);
xor U2484 (N_2484,N_1720,N_1762);
nor U2485 (N_2485,N_1500,N_1965);
xor U2486 (N_2486,N_1731,N_1928);
nand U2487 (N_2487,N_1765,N_1558);
nand U2488 (N_2488,N_1962,N_1917);
and U2489 (N_2489,N_1814,N_1998);
and U2490 (N_2490,N_1560,N_1646);
xnor U2491 (N_2491,N_1909,N_1510);
nor U2492 (N_2492,N_1507,N_1587);
or U2493 (N_2493,N_1587,N_1913);
nand U2494 (N_2494,N_1654,N_1964);
nand U2495 (N_2495,N_1745,N_1595);
or U2496 (N_2496,N_1746,N_1646);
or U2497 (N_2497,N_1530,N_1992);
or U2498 (N_2498,N_1959,N_1737);
or U2499 (N_2499,N_1995,N_1959);
nand U2500 (N_2500,N_2182,N_2166);
nor U2501 (N_2501,N_2013,N_2127);
and U2502 (N_2502,N_2010,N_2227);
and U2503 (N_2503,N_2172,N_2373);
nand U2504 (N_2504,N_2065,N_2395);
nand U2505 (N_2505,N_2210,N_2360);
nor U2506 (N_2506,N_2424,N_2098);
or U2507 (N_2507,N_2443,N_2019);
nor U2508 (N_2508,N_2378,N_2015);
nand U2509 (N_2509,N_2471,N_2126);
or U2510 (N_2510,N_2316,N_2004);
or U2511 (N_2511,N_2130,N_2135);
xor U2512 (N_2512,N_2413,N_2348);
or U2513 (N_2513,N_2299,N_2293);
nor U2514 (N_2514,N_2495,N_2377);
nand U2515 (N_2515,N_2344,N_2043);
xnor U2516 (N_2516,N_2338,N_2254);
nand U2517 (N_2517,N_2107,N_2426);
and U2518 (N_2518,N_2460,N_2491);
and U2519 (N_2519,N_2008,N_2416);
xnor U2520 (N_2520,N_2114,N_2129);
xor U2521 (N_2521,N_2308,N_2080);
nand U2522 (N_2522,N_2297,N_2228);
or U2523 (N_2523,N_2464,N_2234);
nor U2524 (N_2524,N_2487,N_2448);
xor U2525 (N_2525,N_2141,N_2439);
or U2526 (N_2526,N_2383,N_2396);
or U2527 (N_2527,N_2398,N_2097);
nand U2528 (N_2528,N_2068,N_2310);
and U2529 (N_2529,N_2041,N_2156);
xnor U2530 (N_2530,N_2042,N_2478);
nand U2531 (N_2531,N_2488,N_2072);
and U2532 (N_2532,N_2255,N_2260);
and U2533 (N_2533,N_2064,N_2419);
and U2534 (N_2534,N_2158,N_2021);
nor U2535 (N_2535,N_2355,N_2317);
or U2536 (N_2536,N_2112,N_2109);
nor U2537 (N_2537,N_2459,N_2270);
or U2538 (N_2538,N_2067,N_2049);
nor U2539 (N_2539,N_2380,N_2018);
nand U2540 (N_2540,N_2389,N_2334);
xnor U2541 (N_2541,N_2110,N_2306);
or U2542 (N_2542,N_2033,N_2163);
or U2543 (N_2543,N_2406,N_2083);
or U2544 (N_2544,N_2294,N_2220);
xor U2545 (N_2545,N_2428,N_2479);
nor U2546 (N_2546,N_2192,N_2390);
or U2547 (N_2547,N_2167,N_2314);
or U2548 (N_2548,N_2282,N_2438);
xor U2549 (N_2549,N_2054,N_2315);
xnor U2550 (N_2550,N_2187,N_2362);
and U2551 (N_2551,N_2272,N_2077);
xnor U2552 (N_2552,N_2468,N_2427);
nor U2553 (N_2553,N_2082,N_2052);
or U2554 (N_2554,N_2140,N_2235);
nor U2555 (N_2555,N_2216,N_2391);
and U2556 (N_2556,N_2328,N_2247);
nand U2557 (N_2557,N_2193,N_2069);
nand U2558 (N_2558,N_2145,N_2104);
and U2559 (N_2559,N_2300,N_2432);
or U2560 (N_2560,N_2000,N_2403);
or U2561 (N_2561,N_2280,N_2279);
or U2562 (N_2562,N_2274,N_2111);
or U2563 (N_2563,N_2236,N_2040);
or U2564 (N_2564,N_2132,N_2480);
xnor U2565 (N_2565,N_2195,N_2290);
nor U2566 (N_2566,N_2173,N_2092);
nor U2567 (N_2567,N_2181,N_2388);
or U2568 (N_2568,N_2006,N_2162);
and U2569 (N_2569,N_2329,N_2119);
xor U2570 (N_2570,N_2045,N_2418);
and U2571 (N_2571,N_2094,N_2327);
and U2572 (N_2572,N_2204,N_2458);
nand U2573 (N_2573,N_2277,N_2446);
nor U2574 (N_2574,N_2393,N_2245);
xor U2575 (N_2575,N_2475,N_2009);
xor U2576 (N_2576,N_2062,N_2287);
xnor U2577 (N_2577,N_2485,N_2436);
and U2578 (N_2578,N_2269,N_2024);
nor U2579 (N_2579,N_2469,N_2434);
or U2580 (N_2580,N_2307,N_2341);
and U2581 (N_2581,N_2022,N_2302);
and U2582 (N_2582,N_2183,N_2155);
xnor U2583 (N_2583,N_2169,N_2387);
nand U2584 (N_2584,N_2044,N_2440);
nand U2585 (N_2585,N_2159,N_2343);
nor U2586 (N_2586,N_2324,N_2325);
nand U2587 (N_2587,N_2447,N_2425);
xnor U2588 (N_2588,N_2311,N_2451);
and U2589 (N_2589,N_2124,N_2143);
or U2590 (N_2590,N_2101,N_2349);
or U2591 (N_2591,N_2178,N_2121);
and U2592 (N_2592,N_2492,N_2174);
xor U2593 (N_2593,N_2078,N_2081);
nand U2594 (N_2594,N_2149,N_2257);
and U2595 (N_2595,N_2401,N_2177);
nor U2596 (N_2596,N_2146,N_2090);
nor U2597 (N_2597,N_2206,N_2242);
nor U2598 (N_2598,N_2079,N_2250);
nand U2599 (N_2599,N_2455,N_2408);
and U2600 (N_2600,N_2295,N_2122);
nor U2601 (N_2601,N_2409,N_2289);
nor U2602 (N_2602,N_2266,N_2262);
nand U2603 (N_2603,N_2253,N_2025);
nand U2604 (N_2604,N_2100,N_2076);
or U2605 (N_2605,N_2211,N_2298);
or U2606 (N_2606,N_2246,N_2444);
xnor U2607 (N_2607,N_2089,N_2116);
or U2608 (N_2608,N_2356,N_2001);
nor U2609 (N_2609,N_2463,N_2496);
or U2610 (N_2610,N_2281,N_2386);
or U2611 (N_2611,N_2237,N_2256);
nand U2612 (N_2612,N_2093,N_2031);
or U2613 (N_2613,N_2481,N_2137);
and U2614 (N_2614,N_2188,N_2197);
or U2615 (N_2615,N_2131,N_2218);
nor U2616 (N_2616,N_2345,N_2472);
or U2617 (N_2617,N_2333,N_2202);
and U2618 (N_2618,N_2385,N_2309);
and U2619 (N_2619,N_2027,N_2007);
and U2620 (N_2620,N_2394,N_2452);
or U2621 (N_2621,N_2037,N_2136);
or U2622 (N_2622,N_2407,N_2264);
nand U2623 (N_2623,N_2150,N_2028);
and U2624 (N_2624,N_2346,N_2032);
and U2625 (N_2625,N_2194,N_2421);
or U2626 (N_2626,N_2005,N_2217);
nor U2627 (N_2627,N_2258,N_2200);
and U2628 (N_2628,N_2011,N_2050);
nand U2629 (N_2629,N_2352,N_2074);
or U2630 (N_2630,N_2047,N_2171);
nor U2631 (N_2631,N_2291,N_2034);
and U2632 (N_2632,N_2199,N_2108);
and U2633 (N_2633,N_2429,N_2084);
xor U2634 (N_2634,N_2382,N_2030);
nor U2635 (N_2635,N_2180,N_2445);
xnor U2636 (N_2636,N_2465,N_2118);
and U2637 (N_2637,N_2404,N_2450);
xor U2638 (N_2638,N_2437,N_2075);
xnor U2639 (N_2639,N_2326,N_2165);
nor U2640 (N_2640,N_2332,N_2186);
nand U2641 (N_2641,N_2057,N_2223);
xor U2642 (N_2642,N_2240,N_2224);
xnor U2643 (N_2643,N_2139,N_2168);
or U2644 (N_2644,N_2470,N_2369);
and U2645 (N_2645,N_2359,N_2239);
nand U2646 (N_2646,N_2157,N_2476);
nor U2647 (N_2647,N_2339,N_2190);
and U2648 (N_2648,N_2238,N_2494);
or U2649 (N_2649,N_2376,N_2196);
xnor U2650 (N_2650,N_2026,N_2128);
or U2651 (N_2651,N_2288,N_2120);
and U2652 (N_2652,N_2363,N_2219);
or U2653 (N_2653,N_2225,N_2365);
and U2654 (N_2654,N_2353,N_2248);
or U2655 (N_2655,N_2330,N_2154);
nand U2656 (N_2656,N_2466,N_2467);
nor U2657 (N_2657,N_2142,N_2420);
or U2658 (N_2658,N_2189,N_2301);
and U2659 (N_2659,N_2023,N_2207);
or U2660 (N_2660,N_2435,N_2153);
or U2661 (N_2661,N_2384,N_2482);
or U2662 (N_2662,N_2176,N_2493);
xnor U2663 (N_2663,N_2319,N_2433);
and U2664 (N_2664,N_2230,N_2441);
or U2665 (N_2665,N_2268,N_2354);
and U2666 (N_2666,N_2312,N_2321);
xnor U2667 (N_2667,N_2073,N_2414);
xnor U2668 (N_2668,N_2106,N_2051);
and U2669 (N_2669,N_2364,N_2456);
or U2670 (N_2670,N_2271,N_2374);
nor U2671 (N_2671,N_2014,N_2222);
xor U2672 (N_2672,N_2499,N_2358);
nand U2673 (N_2673,N_2400,N_2367);
xnor U2674 (N_2674,N_2267,N_2411);
or U2675 (N_2675,N_2477,N_2350);
xnor U2676 (N_2676,N_2371,N_2048);
or U2677 (N_2677,N_2088,N_2284);
and U2678 (N_2678,N_2461,N_2063);
and U2679 (N_2679,N_2261,N_2160);
xnor U2680 (N_2680,N_2086,N_2313);
and U2681 (N_2681,N_2305,N_2431);
and U2682 (N_2682,N_2351,N_2417);
xor U2683 (N_2683,N_2113,N_2203);
nand U2684 (N_2684,N_2205,N_2053);
or U2685 (N_2685,N_2347,N_2366);
nor U2686 (N_2686,N_2035,N_2296);
xor U2687 (N_2687,N_2002,N_2405);
xnor U2688 (N_2688,N_2484,N_2066);
xnor U2689 (N_2689,N_2342,N_2244);
xnor U2690 (N_2690,N_2410,N_2226);
or U2691 (N_2691,N_2125,N_2215);
nand U2692 (N_2692,N_2095,N_2148);
nor U2693 (N_2693,N_2483,N_2320);
nand U2694 (N_2694,N_2096,N_2012);
xnor U2695 (N_2695,N_2087,N_2213);
or U2696 (N_2696,N_2275,N_2060);
nand U2697 (N_2697,N_2185,N_2191);
xor U2698 (N_2698,N_2214,N_2276);
and U2699 (N_2699,N_2454,N_2133);
nand U2700 (N_2700,N_2375,N_2039);
or U2701 (N_2701,N_2415,N_2457);
and U2702 (N_2702,N_2442,N_2252);
nor U2703 (N_2703,N_2161,N_2379);
xnor U2704 (N_2704,N_2336,N_2105);
nor U2705 (N_2705,N_2020,N_2144);
and U2706 (N_2706,N_2201,N_2381);
or U2707 (N_2707,N_2249,N_2123);
xor U2708 (N_2708,N_2340,N_2091);
nand U2709 (N_2709,N_2016,N_2029);
nor U2710 (N_2710,N_2071,N_2151);
nand U2711 (N_2711,N_2292,N_2085);
nand U2712 (N_2712,N_2179,N_2208);
or U2713 (N_2713,N_2323,N_2038);
nand U2714 (N_2714,N_2059,N_2474);
xnor U2715 (N_2715,N_2241,N_2304);
nand U2716 (N_2716,N_2361,N_2498);
nand U2717 (N_2717,N_2399,N_2231);
xor U2718 (N_2718,N_2318,N_2152);
nor U2719 (N_2719,N_2453,N_2473);
and U2720 (N_2720,N_2497,N_2198);
nor U2721 (N_2721,N_2265,N_2147);
or U2722 (N_2722,N_2370,N_2285);
and U2723 (N_2723,N_2229,N_2335);
or U2724 (N_2724,N_2184,N_2058);
xor U2725 (N_2725,N_2283,N_2331);
nand U2726 (N_2726,N_2102,N_2423);
and U2727 (N_2727,N_2392,N_2322);
or U2728 (N_2728,N_2259,N_2115);
or U2729 (N_2729,N_2134,N_2056);
and U2730 (N_2730,N_2490,N_2099);
nand U2731 (N_2731,N_2422,N_2278);
nand U2732 (N_2732,N_2462,N_2209);
or U2733 (N_2733,N_2017,N_2430);
or U2734 (N_2734,N_2243,N_2221);
xor U2735 (N_2735,N_2233,N_2070);
and U2736 (N_2736,N_2337,N_2486);
nor U2737 (N_2737,N_2357,N_2303);
xnor U2738 (N_2738,N_2138,N_2212);
nor U2739 (N_2739,N_2103,N_2061);
nor U2740 (N_2740,N_2046,N_2368);
xnor U2741 (N_2741,N_2036,N_2412);
or U2742 (N_2742,N_2286,N_2251);
and U2743 (N_2743,N_2055,N_2273);
nand U2744 (N_2744,N_2175,N_2117);
nor U2745 (N_2745,N_2489,N_2003);
and U2746 (N_2746,N_2372,N_2232);
xor U2747 (N_2747,N_2402,N_2263);
xnor U2748 (N_2748,N_2397,N_2170);
nand U2749 (N_2749,N_2449,N_2164);
xnor U2750 (N_2750,N_2268,N_2290);
xor U2751 (N_2751,N_2334,N_2357);
nor U2752 (N_2752,N_2217,N_2129);
and U2753 (N_2753,N_2257,N_2313);
xnor U2754 (N_2754,N_2042,N_2289);
xnor U2755 (N_2755,N_2089,N_2041);
xnor U2756 (N_2756,N_2391,N_2054);
nor U2757 (N_2757,N_2017,N_2025);
nor U2758 (N_2758,N_2354,N_2021);
and U2759 (N_2759,N_2250,N_2425);
and U2760 (N_2760,N_2184,N_2342);
and U2761 (N_2761,N_2174,N_2083);
nor U2762 (N_2762,N_2329,N_2123);
xor U2763 (N_2763,N_2303,N_2431);
or U2764 (N_2764,N_2262,N_2322);
xor U2765 (N_2765,N_2014,N_2467);
xnor U2766 (N_2766,N_2056,N_2087);
nand U2767 (N_2767,N_2219,N_2176);
xnor U2768 (N_2768,N_2133,N_2195);
xor U2769 (N_2769,N_2104,N_2476);
and U2770 (N_2770,N_2118,N_2302);
and U2771 (N_2771,N_2003,N_2293);
xnor U2772 (N_2772,N_2395,N_2148);
or U2773 (N_2773,N_2156,N_2154);
nand U2774 (N_2774,N_2133,N_2441);
nor U2775 (N_2775,N_2346,N_2013);
xnor U2776 (N_2776,N_2324,N_2434);
xor U2777 (N_2777,N_2464,N_2201);
xor U2778 (N_2778,N_2455,N_2237);
or U2779 (N_2779,N_2443,N_2242);
nand U2780 (N_2780,N_2282,N_2028);
xor U2781 (N_2781,N_2052,N_2057);
nand U2782 (N_2782,N_2043,N_2374);
xnor U2783 (N_2783,N_2106,N_2351);
and U2784 (N_2784,N_2179,N_2063);
or U2785 (N_2785,N_2189,N_2152);
nand U2786 (N_2786,N_2450,N_2200);
xor U2787 (N_2787,N_2072,N_2196);
nand U2788 (N_2788,N_2006,N_2405);
nand U2789 (N_2789,N_2408,N_2056);
and U2790 (N_2790,N_2055,N_2255);
and U2791 (N_2791,N_2034,N_2432);
xnor U2792 (N_2792,N_2105,N_2159);
nor U2793 (N_2793,N_2275,N_2297);
xor U2794 (N_2794,N_2099,N_2473);
nor U2795 (N_2795,N_2217,N_2366);
or U2796 (N_2796,N_2317,N_2038);
nand U2797 (N_2797,N_2211,N_2133);
xor U2798 (N_2798,N_2335,N_2401);
nand U2799 (N_2799,N_2458,N_2350);
nand U2800 (N_2800,N_2100,N_2311);
xnor U2801 (N_2801,N_2052,N_2261);
and U2802 (N_2802,N_2085,N_2026);
nand U2803 (N_2803,N_2111,N_2373);
xnor U2804 (N_2804,N_2347,N_2063);
xnor U2805 (N_2805,N_2321,N_2427);
or U2806 (N_2806,N_2205,N_2313);
xor U2807 (N_2807,N_2025,N_2345);
nand U2808 (N_2808,N_2478,N_2325);
or U2809 (N_2809,N_2407,N_2008);
nand U2810 (N_2810,N_2087,N_2454);
and U2811 (N_2811,N_2338,N_2361);
nand U2812 (N_2812,N_2426,N_2126);
or U2813 (N_2813,N_2347,N_2013);
nand U2814 (N_2814,N_2212,N_2289);
xor U2815 (N_2815,N_2041,N_2317);
and U2816 (N_2816,N_2023,N_2388);
xnor U2817 (N_2817,N_2469,N_2136);
nand U2818 (N_2818,N_2239,N_2374);
or U2819 (N_2819,N_2205,N_2412);
xnor U2820 (N_2820,N_2485,N_2427);
nand U2821 (N_2821,N_2355,N_2003);
nor U2822 (N_2822,N_2065,N_2491);
nand U2823 (N_2823,N_2360,N_2119);
nand U2824 (N_2824,N_2242,N_2422);
nor U2825 (N_2825,N_2215,N_2461);
nand U2826 (N_2826,N_2328,N_2027);
xor U2827 (N_2827,N_2470,N_2313);
and U2828 (N_2828,N_2281,N_2323);
xnor U2829 (N_2829,N_2279,N_2420);
nor U2830 (N_2830,N_2203,N_2060);
xor U2831 (N_2831,N_2408,N_2180);
and U2832 (N_2832,N_2068,N_2465);
and U2833 (N_2833,N_2499,N_2498);
nand U2834 (N_2834,N_2246,N_2099);
and U2835 (N_2835,N_2065,N_2002);
xor U2836 (N_2836,N_2264,N_2050);
and U2837 (N_2837,N_2200,N_2249);
or U2838 (N_2838,N_2091,N_2174);
nand U2839 (N_2839,N_2263,N_2280);
or U2840 (N_2840,N_2237,N_2262);
nand U2841 (N_2841,N_2162,N_2263);
xnor U2842 (N_2842,N_2128,N_2425);
xor U2843 (N_2843,N_2071,N_2053);
and U2844 (N_2844,N_2226,N_2302);
nand U2845 (N_2845,N_2049,N_2456);
nor U2846 (N_2846,N_2150,N_2232);
nand U2847 (N_2847,N_2157,N_2430);
or U2848 (N_2848,N_2024,N_2140);
or U2849 (N_2849,N_2070,N_2423);
or U2850 (N_2850,N_2115,N_2472);
nand U2851 (N_2851,N_2454,N_2498);
xor U2852 (N_2852,N_2195,N_2056);
xnor U2853 (N_2853,N_2048,N_2325);
nor U2854 (N_2854,N_2066,N_2153);
nand U2855 (N_2855,N_2215,N_2389);
nor U2856 (N_2856,N_2330,N_2119);
or U2857 (N_2857,N_2431,N_2209);
nand U2858 (N_2858,N_2212,N_2076);
or U2859 (N_2859,N_2085,N_2199);
and U2860 (N_2860,N_2099,N_2401);
or U2861 (N_2861,N_2033,N_2353);
xnor U2862 (N_2862,N_2275,N_2109);
nor U2863 (N_2863,N_2310,N_2158);
xor U2864 (N_2864,N_2487,N_2412);
nand U2865 (N_2865,N_2275,N_2043);
xnor U2866 (N_2866,N_2109,N_2264);
xnor U2867 (N_2867,N_2077,N_2291);
nand U2868 (N_2868,N_2218,N_2328);
nand U2869 (N_2869,N_2102,N_2400);
nand U2870 (N_2870,N_2137,N_2444);
nor U2871 (N_2871,N_2231,N_2100);
xor U2872 (N_2872,N_2049,N_2230);
xor U2873 (N_2873,N_2324,N_2447);
and U2874 (N_2874,N_2262,N_2008);
or U2875 (N_2875,N_2232,N_2447);
or U2876 (N_2876,N_2334,N_2012);
nor U2877 (N_2877,N_2190,N_2064);
and U2878 (N_2878,N_2187,N_2139);
or U2879 (N_2879,N_2360,N_2375);
xnor U2880 (N_2880,N_2302,N_2317);
or U2881 (N_2881,N_2077,N_2413);
and U2882 (N_2882,N_2377,N_2406);
nand U2883 (N_2883,N_2004,N_2222);
or U2884 (N_2884,N_2353,N_2484);
nand U2885 (N_2885,N_2068,N_2012);
or U2886 (N_2886,N_2345,N_2282);
or U2887 (N_2887,N_2249,N_2407);
or U2888 (N_2888,N_2053,N_2315);
or U2889 (N_2889,N_2249,N_2376);
or U2890 (N_2890,N_2211,N_2461);
nor U2891 (N_2891,N_2432,N_2489);
xnor U2892 (N_2892,N_2260,N_2245);
and U2893 (N_2893,N_2419,N_2140);
nand U2894 (N_2894,N_2393,N_2306);
xnor U2895 (N_2895,N_2027,N_2170);
nor U2896 (N_2896,N_2248,N_2358);
nor U2897 (N_2897,N_2424,N_2300);
xor U2898 (N_2898,N_2221,N_2341);
or U2899 (N_2899,N_2422,N_2449);
nor U2900 (N_2900,N_2181,N_2080);
or U2901 (N_2901,N_2445,N_2426);
nand U2902 (N_2902,N_2387,N_2220);
xor U2903 (N_2903,N_2175,N_2472);
nor U2904 (N_2904,N_2145,N_2255);
xnor U2905 (N_2905,N_2257,N_2022);
xor U2906 (N_2906,N_2387,N_2175);
and U2907 (N_2907,N_2013,N_2471);
or U2908 (N_2908,N_2230,N_2208);
xnor U2909 (N_2909,N_2207,N_2416);
and U2910 (N_2910,N_2497,N_2362);
and U2911 (N_2911,N_2037,N_2156);
xnor U2912 (N_2912,N_2046,N_2084);
and U2913 (N_2913,N_2057,N_2119);
or U2914 (N_2914,N_2228,N_2261);
or U2915 (N_2915,N_2198,N_2460);
nor U2916 (N_2916,N_2190,N_2496);
xnor U2917 (N_2917,N_2460,N_2388);
xor U2918 (N_2918,N_2201,N_2062);
nand U2919 (N_2919,N_2278,N_2081);
or U2920 (N_2920,N_2463,N_2371);
and U2921 (N_2921,N_2323,N_2414);
or U2922 (N_2922,N_2481,N_2037);
nor U2923 (N_2923,N_2305,N_2434);
xnor U2924 (N_2924,N_2023,N_2084);
nand U2925 (N_2925,N_2202,N_2281);
and U2926 (N_2926,N_2070,N_2120);
and U2927 (N_2927,N_2277,N_2326);
and U2928 (N_2928,N_2084,N_2229);
nor U2929 (N_2929,N_2210,N_2434);
nor U2930 (N_2930,N_2168,N_2315);
xor U2931 (N_2931,N_2024,N_2021);
nor U2932 (N_2932,N_2368,N_2121);
and U2933 (N_2933,N_2454,N_2475);
xor U2934 (N_2934,N_2136,N_2234);
nor U2935 (N_2935,N_2451,N_2168);
or U2936 (N_2936,N_2405,N_2425);
and U2937 (N_2937,N_2045,N_2361);
nor U2938 (N_2938,N_2394,N_2011);
nor U2939 (N_2939,N_2151,N_2241);
xor U2940 (N_2940,N_2006,N_2392);
nand U2941 (N_2941,N_2222,N_2168);
xnor U2942 (N_2942,N_2093,N_2340);
or U2943 (N_2943,N_2256,N_2444);
nand U2944 (N_2944,N_2209,N_2480);
nor U2945 (N_2945,N_2227,N_2073);
and U2946 (N_2946,N_2069,N_2006);
xor U2947 (N_2947,N_2323,N_2314);
and U2948 (N_2948,N_2420,N_2275);
xor U2949 (N_2949,N_2442,N_2005);
nor U2950 (N_2950,N_2475,N_2030);
or U2951 (N_2951,N_2286,N_2408);
nand U2952 (N_2952,N_2195,N_2411);
xnor U2953 (N_2953,N_2051,N_2296);
or U2954 (N_2954,N_2493,N_2272);
nor U2955 (N_2955,N_2464,N_2150);
and U2956 (N_2956,N_2169,N_2216);
xnor U2957 (N_2957,N_2494,N_2466);
and U2958 (N_2958,N_2040,N_2232);
nor U2959 (N_2959,N_2216,N_2135);
nor U2960 (N_2960,N_2044,N_2473);
nor U2961 (N_2961,N_2027,N_2078);
nor U2962 (N_2962,N_2133,N_2064);
xnor U2963 (N_2963,N_2352,N_2327);
and U2964 (N_2964,N_2114,N_2126);
or U2965 (N_2965,N_2112,N_2472);
or U2966 (N_2966,N_2187,N_2366);
nand U2967 (N_2967,N_2333,N_2275);
and U2968 (N_2968,N_2138,N_2193);
xor U2969 (N_2969,N_2406,N_2436);
or U2970 (N_2970,N_2243,N_2076);
nor U2971 (N_2971,N_2290,N_2344);
nand U2972 (N_2972,N_2280,N_2476);
and U2973 (N_2973,N_2419,N_2300);
xor U2974 (N_2974,N_2326,N_2021);
nor U2975 (N_2975,N_2396,N_2331);
nor U2976 (N_2976,N_2010,N_2382);
xor U2977 (N_2977,N_2181,N_2336);
and U2978 (N_2978,N_2087,N_2299);
and U2979 (N_2979,N_2140,N_2070);
nand U2980 (N_2980,N_2259,N_2147);
xor U2981 (N_2981,N_2349,N_2228);
or U2982 (N_2982,N_2204,N_2077);
xnor U2983 (N_2983,N_2126,N_2306);
and U2984 (N_2984,N_2486,N_2043);
xnor U2985 (N_2985,N_2219,N_2450);
xor U2986 (N_2986,N_2381,N_2052);
nand U2987 (N_2987,N_2086,N_2360);
or U2988 (N_2988,N_2466,N_2493);
or U2989 (N_2989,N_2374,N_2049);
or U2990 (N_2990,N_2474,N_2355);
xnor U2991 (N_2991,N_2138,N_2047);
nor U2992 (N_2992,N_2234,N_2090);
nand U2993 (N_2993,N_2230,N_2460);
xnor U2994 (N_2994,N_2474,N_2293);
nand U2995 (N_2995,N_2001,N_2263);
xor U2996 (N_2996,N_2445,N_2035);
nand U2997 (N_2997,N_2242,N_2319);
xnor U2998 (N_2998,N_2364,N_2346);
or U2999 (N_2999,N_2093,N_2258);
nor U3000 (N_3000,N_2549,N_2573);
xor U3001 (N_3001,N_2669,N_2921);
nand U3002 (N_3002,N_2913,N_2515);
nand U3003 (N_3003,N_2505,N_2772);
nor U3004 (N_3004,N_2973,N_2626);
xor U3005 (N_3005,N_2998,N_2993);
nor U3006 (N_3006,N_2781,N_2634);
nor U3007 (N_3007,N_2715,N_2615);
and U3008 (N_3008,N_2743,N_2567);
nor U3009 (N_3009,N_2991,N_2992);
nor U3010 (N_3010,N_2564,N_2720);
xnor U3011 (N_3011,N_2907,N_2773);
nor U3012 (N_3012,N_2937,N_2541);
nand U3013 (N_3013,N_2905,N_2696);
nand U3014 (N_3014,N_2938,N_2956);
xor U3015 (N_3015,N_2569,N_2925);
or U3016 (N_3016,N_2857,N_2863);
nor U3017 (N_3017,N_2899,N_2860);
and U3018 (N_3018,N_2874,N_2639);
xor U3019 (N_3019,N_2592,N_2928);
and U3020 (N_3020,N_2994,N_2801);
or U3021 (N_3021,N_2616,N_2896);
nand U3022 (N_3022,N_2757,N_2789);
xnor U3023 (N_3023,N_2737,N_2710);
nand U3024 (N_3024,N_2954,N_2841);
and U3025 (N_3025,N_2837,N_2545);
xnor U3026 (N_3026,N_2783,N_2731);
nand U3027 (N_3027,N_2756,N_2680);
xor U3028 (N_3028,N_2768,N_2661);
and U3029 (N_3029,N_2791,N_2604);
nor U3030 (N_3030,N_2628,N_2562);
or U3031 (N_3031,N_2678,N_2532);
nand U3032 (N_3032,N_2817,N_2664);
nand U3033 (N_3033,N_2765,N_2693);
xnor U3034 (N_3034,N_2792,N_2811);
and U3035 (N_3035,N_2797,N_2924);
nand U3036 (N_3036,N_2514,N_2578);
and U3037 (N_3037,N_2866,N_2887);
xnor U3038 (N_3038,N_2873,N_2581);
and U3039 (N_3039,N_2605,N_2920);
or U3040 (N_3040,N_2900,N_2651);
and U3041 (N_3041,N_2527,N_2915);
or U3042 (N_3042,N_2577,N_2796);
xor U3043 (N_3043,N_2802,N_2804);
nor U3044 (N_3044,N_2936,N_2613);
xnor U3045 (N_3045,N_2629,N_2805);
and U3046 (N_3046,N_2587,N_2875);
or U3047 (N_3047,N_2555,N_2660);
nor U3048 (N_3048,N_2986,N_2823);
and U3049 (N_3049,N_2949,N_2622);
and U3050 (N_3050,N_2670,N_2542);
or U3051 (N_3051,N_2561,N_2704);
and U3052 (N_3052,N_2926,N_2812);
nor U3053 (N_3053,N_2816,N_2526);
or U3054 (N_3054,N_2788,N_2951);
xor U3055 (N_3055,N_2729,N_2927);
nand U3056 (N_3056,N_2847,N_2775);
xor U3057 (N_3057,N_2785,N_2674);
or U3058 (N_3058,N_2908,N_2895);
xor U3059 (N_3059,N_2663,N_2786);
or U3060 (N_3060,N_2962,N_2889);
xor U3061 (N_3061,N_2685,N_2643);
and U3062 (N_3062,N_2760,N_2976);
nor U3063 (N_3063,N_2929,N_2624);
xor U3064 (N_3064,N_2815,N_2647);
and U3065 (N_3065,N_2723,N_2627);
xnor U3066 (N_3066,N_2974,N_2763);
and U3067 (N_3067,N_2960,N_2984);
nor U3068 (N_3068,N_2558,N_2610);
nand U3069 (N_3069,N_2739,N_2566);
nand U3070 (N_3070,N_2885,N_2594);
or U3071 (N_3071,N_2881,N_2673);
and U3072 (N_3072,N_2912,N_2892);
xnor U3073 (N_3073,N_2935,N_2824);
nand U3074 (N_3074,N_2563,N_2808);
and U3075 (N_3075,N_2699,N_2849);
and U3076 (N_3076,N_2667,N_2834);
xnor U3077 (N_3077,N_2738,N_2518);
or U3078 (N_3078,N_2657,N_2679);
nand U3079 (N_3079,N_2883,N_2948);
xor U3080 (N_3080,N_2891,N_2982);
nor U3081 (N_3081,N_2556,N_2807);
xnor U3082 (N_3082,N_2825,N_2803);
nand U3083 (N_3083,N_2599,N_2787);
nand U3084 (N_3084,N_2658,N_2979);
nor U3085 (N_3085,N_2537,N_2560);
and U3086 (N_3086,N_2888,N_2513);
xnor U3087 (N_3087,N_2850,N_2641);
and U3088 (N_3088,N_2557,N_2827);
nand U3089 (N_3089,N_2821,N_2918);
nor U3090 (N_3090,N_2607,N_2876);
or U3091 (N_3091,N_2822,N_2902);
and U3092 (N_3092,N_2517,N_2508);
or U3093 (N_3093,N_2941,N_2602);
or U3094 (N_3094,N_2521,N_2922);
and U3095 (N_3095,N_2702,N_2632);
xnor U3096 (N_3096,N_2845,N_2846);
and U3097 (N_3097,N_2550,N_2923);
and U3098 (N_3098,N_2726,N_2844);
xor U3099 (N_3099,N_2539,N_2590);
and U3100 (N_3100,N_2869,N_2620);
and U3101 (N_3101,N_2547,N_2574);
xnor U3102 (N_3102,N_2852,N_2633);
nand U3103 (N_3103,N_2609,N_2831);
or U3104 (N_3104,N_2934,N_2770);
xor U3105 (N_3105,N_2722,N_2855);
nor U3106 (N_3106,N_2600,N_2681);
or U3107 (N_3107,N_2582,N_2886);
nor U3108 (N_3108,N_2843,N_2777);
or U3109 (N_3109,N_2799,N_2612);
nor U3110 (N_3110,N_2608,N_2870);
nand U3111 (N_3111,N_2940,N_2649);
xor U3112 (N_3112,N_2665,N_2516);
nor U3113 (N_3113,N_2961,N_2893);
xor U3114 (N_3114,N_2512,N_2753);
or U3115 (N_3115,N_2751,N_2698);
xor U3116 (N_3116,N_2551,N_2859);
xnor U3117 (N_3117,N_2759,N_2809);
and U3118 (N_3118,N_2705,N_2682);
and U3119 (N_3119,N_2636,N_2585);
and U3120 (N_3120,N_2959,N_2540);
or U3121 (N_3121,N_2964,N_2598);
and U3122 (N_3122,N_2832,N_2706);
xnor U3123 (N_3123,N_2880,N_2884);
nand U3124 (N_3124,N_2828,N_2999);
nand U3125 (N_3125,N_2712,N_2983);
xnor U3126 (N_3126,N_2583,N_2906);
nor U3127 (N_3127,N_2736,N_2637);
and U3128 (N_3128,N_2732,N_2980);
and U3129 (N_3129,N_2676,N_2793);
or U3130 (N_3130,N_2761,N_2718);
nor U3131 (N_3131,N_2656,N_2507);
and U3132 (N_3132,N_2611,N_2839);
or U3133 (N_3133,N_2575,N_2529);
nor U3134 (N_3134,N_2504,N_2691);
or U3135 (N_3135,N_2619,N_2990);
nor U3136 (N_3136,N_2543,N_2531);
and U3137 (N_3137,N_2972,N_2584);
xor U3138 (N_3138,N_2947,N_2695);
and U3139 (N_3139,N_2943,N_2588);
or U3140 (N_3140,N_2957,N_2652);
xnor U3141 (N_3141,N_2606,N_2601);
nand U3142 (N_3142,N_2591,N_2830);
xor U3143 (N_3143,N_2829,N_2953);
nand U3144 (N_3144,N_2645,N_2942);
or U3145 (N_3145,N_2501,N_2559);
or U3146 (N_3146,N_2981,N_2995);
xnor U3147 (N_3147,N_2571,N_2835);
and U3148 (N_3148,N_2523,N_2630);
and U3149 (N_3149,N_2820,N_2910);
or U3150 (N_3150,N_2528,N_2554);
xnor U3151 (N_3151,N_2795,N_2909);
and U3152 (N_3152,N_2914,N_2752);
nand U3153 (N_3153,N_2589,N_2677);
and U3154 (N_3154,N_2690,N_2684);
nand U3155 (N_3155,N_2997,N_2697);
or U3156 (N_3156,N_2689,N_2692);
or U3157 (N_3157,N_2872,N_2776);
nor U3158 (N_3158,N_2944,N_2733);
and U3159 (N_3159,N_2769,N_2520);
xnor U3160 (N_3160,N_2952,N_2919);
nand U3161 (N_3161,N_2868,N_2987);
or U3162 (N_3162,N_2700,N_2945);
or U3163 (N_3163,N_2650,N_2533);
and U3164 (N_3164,N_2764,N_2966);
nand U3165 (N_3165,N_2522,N_2848);
xnor U3166 (N_3166,N_2836,N_2818);
xor U3167 (N_3167,N_2687,N_2854);
nor U3168 (N_3168,N_2975,N_2806);
nand U3169 (N_3169,N_2683,N_2958);
xnor U3170 (N_3170,N_2666,N_2894);
nand U3171 (N_3171,N_2749,N_2734);
nor U3172 (N_3172,N_2748,N_2717);
nand U3173 (N_3173,N_2766,N_2978);
nand U3174 (N_3174,N_2780,N_2502);
nand U3175 (N_3175,N_2968,N_2813);
and U3176 (N_3176,N_2878,N_2534);
nor U3177 (N_3177,N_2969,N_2525);
or U3178 (N_3178,N_2930,N_2861);
or U3179 (N_3179,N_2635,N_2742);
nor U3180 (N_3180,N_2735,N_2595);
nor U3181 (N_3181,N_2707,N_2867);
and U3182 (N_3182,N_2955,N_2903);
or U3183 (N_3183,N_2782,N_2898);
and U3184 (N_3184,N_2916,N_2728);
and U3185 (N_3185,N_2904,N_2646);
and U3186 (N_3186,N_2901,N_2858);
nand U3187 (N_3187,N_2988,N_2890);
and U3188 (N_3188,N_2688,N_2586);
nor U3189 (N_3189,N_2826,N_2638);
and U3190 (N_3190,N_2897,N_2977);
nor U3191 (N_3191,N_2862,N_2714);
nor U3192 (N_3192,N_2882,N_2725);
and U3193 (N_3193,N_2819,N_2553);
nand U3194 (N_3194,N_2642,N_2565);
nand U3195 (N_3195,N_2967,N_2597);
or U3196 (N_3196,N_2536,N_2509);
nor U3197 (N_3197,N_2933,N_2744);
xnor U3198 (N_3198,N_2985,N_2524);
and U3199 (N_3199,N_2794,N_2570);
and U3200 (N_3200,N_2864,N_2814);
nor U3201 (N_3201,N_2740,N_2719);
or U3202 (N_3202,N_2784,N_2640);
nand U3203 (N_3203,N_2713,N_2544);
and U3204 (N_3204,N_2621,N_2576);
nor U3205 (N_3205,N_2931,N_2703);
and U3206 (N_3206,N_2970,N_2546);
xor U3207 (N_3207,N_2675,N_2686);
nor U3208 (N_3208,N_2580,N_2579);
nand U3209 (N_3209,N_2779,N_2996);
and U3210 (N_3210,N_2631,N_2668);
nor U3211 (N_3211,N_2519,N_2552);
nand U3212 (N_3212,N_2648,N_2851);
and U3213 (N_3213,N_2856,N_2654);
and U3214 (N_3214,N_2932,N_2655);
nand U3215 (N_3215,N_2755,N_2911);
and U3216 (N_3216,N_2758,N_2762);
nor U3217 (N_3217,N_2625,N_2535);
xor U3218 (N_3218,N_2939,N_2503);
nand U3219 (N_3219,N_2671,N_2871);
nor U3220 (N_3220,N_2727,N_2767);
nand U3221 (N_3221,N_2617,N_2989);
nor U3222 (N_3222,N_2614,N_2506);
nand U3223 (N_3223,N_2618,N_2708);
and U3224 (N_3224,N_2810,N_2917);
xor U3225 (N_3225,N_2842,N_2741);
or U3226 (N_3226,N_2965,N_2877);
xnor U3227 (N_3227,N_2711,N_2659);
xnor U3228 (N_3228,N_2694,N_2750);
xor U3229 (N_3229,N_2798,N_2653);
xor U3230 (N_3230,N_2745,N_2730);
nor U3231 (N_3231,N_2672,N_2701);
or U3232 (N_3232,N_2774,N_2548);
and U3233 (N_3233,N_2596,N_2724);
nand U3234 (N_3234,N_2530,N_2833);
nor U3235 (N_3235,N_2840,N_2709);
and U3236 (N_3236,N_2572,N_2747);
nor U3237 (N_3237,N_2593,N_2644);
and U3238 (N_3238,N_2510,N_2716);
or U3239 (N_3239,N_2746,N_2971);
xnor U3240 (N_3240,N_2800,N_2963);
nand U3241 (N_3241,N_2568,N_2853);
or U3242 (N_3242,N_2771,N_2603);
nor U3243 (N_3243,N_2950,N_2623);
nor U3244 (N_3244,N_2538,N_2778);
xnor U3245 (N_3245,N_2865,N_2838);
xor U3246 (N_3246,N_2721,N_2662);
nand U3247 (N_3247,N_2754,N_2946);
and U3248 (N_3248,N_2790,N_2511);
and U3249 (N_3249,N_2879,N_2500);
xor U3250 (N_3250,N_2950,N_2861);
nor U3251 (N_3251,N_2549,N_2906);
and U3252 (N_3252,N_2612,N_2763);
nor U3253 (N_3253,N_2696,N_2872);
nand U3254 (N_3254,N_2575,N_2982);
nand U3255 (N_3255,N_2778,N_2959);
nand U3256 (N_3256,N_2625,N_2791);
or U3257 (N_3257,N_2533,N_2987);
or U3258 (N_3258,N_2990,N_2905);
nand U3259 (N_3259,N_2748,N_2790);
nand U3260 (N_3260,N_2589,N_2728);
and U3261 (N_3261,N_2767,N_2918);
nand U3262 (N_3262,N_2686,N_2830);
or U3263 (N_3263,N_2745,N_2907);
nor U3264 (N_3264,N_2616,N_2731);
xor U3265 (N_3265,N_2927,N_2718);
or U3266 (N_3266,N_2934,N_2674);
xor U3267 (N_3267,N_2620,N_2582);
or U3268 (N_3268,N_2551,N_2802);
or U3269 (N_3269,N_2690,N_2595);
nand U3270 (N_3270,N_2518,N_2784);
xnor U3271 (N_3271,N_2960,N_2813);
and U3272 (N_3272,N_2508,N_2997);
xor U3273 (N_3273,N_2575,N_2662);
nand U3274 (N_3274,N_2978,N_2818);
or U3275 (N_3275,N_2711,N_2728);
xnor U3276 (N_3276,N_2885,N_2608);
and U3277 (N_3277,N_2606,N_2943);
and U3278 (N_3278,N_2781,N_2594);
and U3279 (N_3279,N_2727,N_2599);
xnor U3280 (N_3280,N_2777,N_2974);
xnor U3281 (N_3281,N_2785,N_2778);
nand U3282 (N_3282,N_2631,N_2609);
nand U3283 (N_3283,N_2768,N_2634);
nor U3284 (N_3284,N_2669,N_2764);
nand U3285 (N_3285,N_2610,N_2572);
nand U3286 (N_3286,N_2994,N_2992);
nand U3287 (N_3287,N_2977,N_2658);
nor U3288 (N_3288,N_2742,N_2808);
or U3289 (N_3289,N_2816,N_2797);
or U3290 (N_3290,N_2721,N_2701);
or U3291 (N_3291,N_2872,N_2509);
and U3292 (N_3292,N_2695,N_2980);
and U3293 (N_3293,N_2867,N_2575);
nor U3294 (N_3294,N_2850,N_2943);
nand U3295 (N_3295,N_2780,N_2772);
nand U3296 (N_3296,N_2931,N_2951);
xnor U3297 (N_3297,N_2859,N_2965);
or U3298 (N_3298,N_2670,N_2950);
or U3299 (N_3299,N_2583,N_2682);
and U3300 (N_3300,N_2881,N_2671);
nor U3301 (N_3301,N_2990,N_2951);
nor U3302 (N_3302,N_2789,N_2677);
nor U3303 (N_3303,N_2975,N_2589);
nand U3304 (N_3304,N_2550,N_2733);
xnor U3305 (N_3305,N_2765,N_2775);
nand U3306 (N_3306,N_2742,N_2910);
xor U3307 (N_3307,N_2576,N_2680);
nand U3308 (N_3308,N_2622,N_2630);
and U3309 (N_3309,N_2667,N_2739);
xnor U3310 (N_3310,N_2708,N_2905);
and U3311 (N_3311,N_2578,N_2857);
nand U3312 (N_3312,N_2917,N_2728);
nand U3313 (N_3313,N_2675,N_2595);
and U3314 (N_3314,N_2856,N_2614);
xnor U3315 (N_3315,N_2504,N_2980);
and U3316 (N_3316,N_2921,N_2556);
xor U3317 (N_3317,N_2930,N_2819);
and U3318 (N_3318,N_2613,N_2797);
and U3319 (N_3319,N_2966,N_2501);
and U3320 (N_3320,N_2546,N_2812);
or U3321 (N_3321,N_2916,N_2751);
or U3322 (N_3322,N_2856,N_2629);
nor U3323 (N_3323,N_2533,N_2740);
nand U3324 (N_3324,N_2907,N_2922);
nand U3325 (N_3325,N_2629,N_2768);
xnor U3326 (N_3326,N_2724,N_2830);
xnor U3327 (N_3327,N_2934,N_2528);
or U3328 (N_3328,N_2984,N_2547);
nand U3329 (N_3329,N_2750,N_2734);
xnor U3330 (N_3330,N_2625,N_2946);
and U3331 (N_3331,N_2607,N_2514);
xor U3332 (N_3332,N_2843,N_2573);
xnor U3333 (N_3333,N_2822,N_2733);
and U3334 (N_3334,N_2794,N_2858);
or U3335 (N_3335,N_2504,N_2897);
and U3336 (N_3336,N_2584,N_2511);
nand U3337 (N_3337,N_2802,N_2535);
nor U3338 (N_3338,N_2882,N_2674);
and U3339 (N_3339,N_2649,N_2925);
nor U3340 (N_3340,N_2785,N_2603);
nand U3341 (N_3341,N_2586,N_2810);
and U3342 (N_3342,N_2579,N_2977);
or U3343 (N_3343,N_2908,N_2962);
or U3344 (N_3344,N_2579,N_2551);
xor U3345 (N_3345,N_2825,N_2580);
nor U3346 (N_3346,N_2633,N_2664);
nand U3347 (N_3347,N_2695,N_2895);
nor U3348 (N_3348,N_2747,N_2922);
nand U3349 (N_3349,N_2700,N_2733);
nor U3350 (N_3350,N_2850,N_2778);
nand U3351 (N_3351,N_2524,N_2663);
nor U3352 (N_3352,N_2744,N_2723);
xnor U3353 (N_3353,N_2530,N_2548);
nor U3354 (N_3354,N_2708,N_2858);
nand U3355 (N_3355,N_2819,N_2613);
nand U3356 (N_3356,N_2746,N_2983);
nor U3357 (N_3357,N_2751,N_2867);
nand U3358 (N_3358,N_2709,N_2570);
or U3359 (N_3359,N_2940,N_2752);
nand U3360 (N_3360,N_2942,N_2910);
nor U3361 (N_3361,N_2794,N_2911);
nor U3362 (N_3362,N_2645,N_2921);
and U3363 (N_3363,N_2536,N_2721);
nand U3364 (N_3364,N_2695,N_2964);
xnor U3365 (N_3365,N_2746,N_2766);
nor U3366 (N_3366,N_2731,N_2535);
and U3367 (N_3367,N_2885,N_2883);
and U3368 (N_3368,N_2871,N_2827);
nand U3369 (N_3369,N_2808,N_2744);
nand U3370 (N_3370,N_2847,N_2610);
nor U3371 (N_3371,N_2908,N_2936);
or U3372 (N_3372,N_2931,N_2568);
or U3373 (N_3373,N_2518,N_2646);
nand U3374 (N_3374,N_2551,N_2717);
or U3375 (N_3375,N_2738,N_2833);
and U3376 (N_3376,N_2522,N_2811);
xnor U3377 (N_3377,N_2677,N_2519);
nand U3378 (N_3378,N_2787,N_2630);
xor U3379 (N_3379,N_2635,N_2632);
and U3380 (N_3380,N_2828,N_2756);
nand U3381 (N_3381,N_2645,N_2940);
nand U3382 (N_3382,N_2829,N_2777);
nor U3383 (N_3383,N_2644,N_2960);
nor U3384 (N_3384,N_2510,N_2694);
xnor U3385 (N_3385,N_2600,N_2874);
or U3386 (N_3386,N_2682,N_2971);
nand U3387 (N_3387,N_2559,N_2579);
or U3388 (N_3388,N_2618,N_2789);
or U3389 (N_3389,N_2903,N_2745);
or U3390 (N_3390,N_2709,N_2566);
nand U3391 (N_3391,N_2755,N_2799);
nor U3392 (N_3392,N_2725,N_2614);
xnor U3393 (N_3393,N_2610,N_2636);
or U3394 (N_3394,N_2863,N_2761);
xor U3395 (N_3395,N_2717,N_2832);
or U3396 (N_3396,N_2875,N_2829);
nand U3397 (N_3397,N_2869,N_2673);
nor U3398 (N_3398,N_2918,N_2710);
nor U3399 (N_3399,N_2520,N_2850);
nand U3400 (N_3400,N_2753,N_2920);
nor U3401 (N_3401,N_2987,N_2794);
nand U3402 (N_3402,N_2896,N_2676);
and U3403 (N_3403,N_2824,N_2963);
or U3404 (N_3404,N_2926,N_2729);
or U3405 (N_3405,N_2709,N_2563);
nand U3406 (N_3406,N_2551,N_2985);
or U3407 (N_3407,N_2790,N_2779);
nor U3408 (N_3408,N_2811,N_2521);
xnor U3409 (N_3409,N_2614,N_2638);
nor U3410 (N_3410,N_2781,N_2748);
and U3411 (N_3411,N_2510,N_2725);
xor U3412 (N_3412,N_2916,N_2541);
and U3413 (N_3413,N_2954,N_2896);
or U3414 (N_3414,N_2671,N_2667);
and U3415 (N_3415,N_2745,N_2760);
nor U3416 (N_3416,N_2962,N_2820);
nor U3417 (N_3417,N_2786,N_2714);
nor U3418 (N_3418,N_2885,N_2851);
or U3419 (N_3419,N_2809,N_2851);
and U3420 (N_3420,N_2753,N_2932);
xor U3421 (N_3421,N_2766,N_2618);
xor U3422 (N_3422,N_2685,N_2585);
nand U3423 (N_3423,N_2683,N_2508);
nor U3424 (N_3424,N_2772,N_2906);
nor U3425 (N_3425,N_2514,N_2619);
nor U3426 (N_3426,N_2776,N_2988);
nand U3427 (N_3427,N_2602,N_2710);
xnor U3428 (N_3428,N_2899,N_2741);
nand U3429 (N_3429,N_2977,N_2837);
and U3430 (N_3430,N_2906,N_2619);
or U3431 (N_3431,N_2768,N_2879);
xnor U3432 (N_3432,N_2515,N_2571);
and U3433 (N_3433,N_2863,N_2547);
and U3434 (N_3434,N_2592,N_2886);
xor U3435 (N_3435,N_2816,N_2939);
or U3436 (N_3436,N_2641,N_2981);
nor U3437 (N_3437,N_2847,N_2838);
and U3438 (N_3438,N_2559,N_2699);
or U3439 (N_3439,N_2953,N_2995);
or U3440 (N_3440,N_2888,N_2937);
or U3441 (N_3441,N_2500,N_2895);
and U3442 (N_3442,N_2848,N_2531);
or U3443 (N_3443,N_2701,N_2918);
xnor U3444 (N_3444,N_2753,N_2893);
or U3445 (N_3445,N_2870,N_2698);
or U3446 (N_3446,N_2632,N_2756);
or U3447 (N_3447,N_2849,N_2516);
nand U3448 (N_3448,N_2676,N_2538);
nand U3449 (N_3449,N_2643,N_2972);
nor U3450 (N_3450,N_2830,N_2807);
nand U3451 (N_3451,N_2766,N_2517);
xnor U3452 (N_3452,N_2970,N_2654);
nand U3453 (N_3453,N_2504,N_2776);
or U3454 (N_3454,N_2598,N_2807);
nand U3455 (N_3455,N_2796,N_2568);
nand U3456 (N_3456,N_2721,N_2521);
xor U3457 (N_3457,N_2887,N_2961);
xor U3458 (N_3458,N_2511,N_2900);
or U3459 (N_3459,N_2503,N_2768);
xor U3460 (N_3460,N_2546,N_2745);
nand U3461 (N_3461,N_2778,N_2815);
nor U3462 (N_3462,N_2715,N_2649);
and U3463 (N_3463,N_2887,N_2761);
xor U3464 (N_3464,N_2578,N_2677);
nand U3465 (N_3465,N_2903,N_2799);
and U3466 (N_3466,N_2667,N_2743);
and U3467 (N_3467,N_2947,N_2978);
xor U3468 (N_3468,N_2624,N_2963);
nor U3469 (N_3469,N_2847,N_2755);
xor U3470 (N_3470,N_2620,N_2980);
or U3471 (N_3471,N_2636,N_2888);
xnor U3472 (N_3472,N_2923,N_2532);
nor U3473 (N_3473,N_2941,N_2974);
or U3474 (N_3474,N_2835,N_2729);
nor U3475 (N_3475,N_2782,N_2952);
and U3476 (N_3476,N_2619,N_2857);
nand U3477 (N_3477,N_2662,N_2849);
nand U3478 (N_3478,N_2720,N_2546);
nor U3479 (N_3479,N_2954,N_2711);
and U3480 (N_3480,N_2587,N_2855);
or U3481 (N_3481,N_2924,N_2619);
or U3482 (N_3482,N_2641,N_2722);
nand U3483 (N_3483,N_2950,N_2771);
and U3484 (N_3484,N_2869,N_2654);
nor U3485 (N_3485,N_2630,N_2511);
xnor U3486 (N_3486,N_2730,N_2518);
xor U3487 (N_3487,N_2958,N_2630);
nand U3488 (N_3488,N_2695,N_2762);
nor U3489 (N_3489,N_2697,N_2799);
xnor U3490 (N_3490,N_2740,N_2705);
nor U3491 (N_3491,N_2702,N_2780);
xor U3492 (N_3492,N_2905,N_2743);
nand U3493 (N_3493,N_2501,N_2773);
nor U3494 (N_3494,N_2833,N_2603);
nand U3495 (N_3495,N_2886,N_2530);
and U3496 (N_3496,N_2572,N_2896);
xnor U3497 (N_3497,N_2969,N_2599);
nand U3498 (N_3498,N_2532,N_2873);
xnor U3499 (N_3499,N_2849,N_2718);
nand U3500 (N_3500,N_3335,N_3234);
nand U3501 (N_3501,N_3462,N_3048);
or U3502 (N_3502,N_3031,N_3178);
and U3503 (N_3503,N_3477,N_3490);
nand U3504 (N_3504,N_3438,N_3167);
nor U3505 (N_3505,N_3202,N_3085);
xor U3506 (N_3506,N_3053,N_3452);
xnor U3507 (N_3507,N_3212,N_3460);
nor U3508 (N_3508,N_3447,N_3141);
xor U3509 (N_3509,N_3214,N_3400);
nand U3510 (N_3510,N_3349,N_3421);
or U3511 (N_3511,N_3177,N_3489);
or U3512 (N_3512,N_3102,N_3316);
nand U3513 (N_3513,N_3379,N_3290);
or U3514 (N_3514,N_3424,N_3049);
nand U3515 (N_3515,N_3382,N_3330);
nand U3516 (N_3516,N_3044,N_3340);
xnor U3517 (N_3517,N_3001,N_3180);
nand U3518 (N_3518,N_3124,N_3226);
xor U3519 (N_3519,N_3241,N_3172);
and U3520 (N_3520,N_3188,N_3415);
nand U3521 (N_3521,N_3197,N_3487);
nor U3522 (N_3522,N_3118,N_3348);
xor U3523 (N_3523,N_3357,N_3100);
or U3524 (N_3524,N_3138,N_3484);
or U3525 (N_3525,N_3297,N_3459);
and U3526 (N_3526,N_3272,N_3485);
nand U3527 (N_3527,N_3223,N_3037);
or U3528 (N_3528,N_3018,N_3077);
nand U3529 (N_3529,N_3030,N_3215);
nor U3530 (N_3530,N_3148,N_3450);
xor U3531 (N_3531,N_3213,N_3363);
xor U3532 (N_3532,N_3155,N_3281);
xnor U3533 (N_3533,N_3029,N_3303);
and U3534 (N_3534,N_3145,N_3398);
nor U3535 (N_3535,N_3371,N_3169);
and U3536 (N_3536,N_3122,N_3367);
xor U3537 (N_3537,N_3228,N_3354);
nand U3538 (N_3538,N_3350,N_3170);
or U3539 (N_3539,N_3262,N_3404);
nand U3540 (N_3540,N_3322,N_3426);
nor U3541 (N_3541,N_3105,N_3099);
nand U3542 (N_3542,N_3005,N_3331);
nand U3543 (N_3543,N_3181,N_3098);
nor U3544 (N_3544,N_3358,N_3229);
nand U3545 (N_3545,N_3254,N_3142);
nor U3546 (N_3546,N_3417,N_3144);
and U3547 (N_3547,N_3458,N_3478);
or U3548 (N_3548,N_3461,N_3394);
nor U3549 (N_3549,N_3230,N_3004);
or U3550 (N_3550,N_3034,N_3065);
xor U3551 (N_3551,N_3020,N_3446);
or U3552 (N_3552,N_3219,N_3470);
or U3553 (N_3553,N_3119,N_3327);
xnor U3554 (N_3554,N_3043,N_3496);
or U3555 (N_3555,N_3440,N_3285);
xnor U3556 (N_3556,N_3271,N_3083);
and U3557 (N_3557,N_3027,N_3304);
and U3558 (N_3558,N_3074,N_3129);
xnor U3559 (N_3559,N_3292,N_3078);
xor U3560 (N_3560,N_3107,N_3036);
and U3561 (N_3561,N_3023,N_3052);
nor U3562 (N_3562,N_3273,N_3259);
or U3563 (N_3563,N_3301,N_3051);
nor U3564 (N_3564,N_3481,N_3407);
xnor U3565 (N_3565,N_3130,N_3439);
nor U3566 (N_3566,N_3482,N_3058);
nand U3567 (N_3567,N_3282,N_3240);
xnor U3568 (N_3568,N_3416,N_3474);
or U3569 (N_3569,N_3380,N_3066);
nor U3570 (N_3570,N_3260,N_3015);
and U3571 (N_3571,N_3498,N_3093);
nand U3572 (N_3572,N_3255,N_3256);
nand U3573 (N_3573,N_3061,N_3464);
xnor U3574 (N_3574,N_3205,N_3154);
and U3575 (N_3575,N_3243,N_3224);
or U3576 (N_3576,N_3342,N_3033);
nand U3577 (N_3577,N_3266,N_3305);
xnor U3578 (N_3578,N_3203,N_3073);
or U3579 (N_3579,N_3179,N_3465);
nand U3580 (N_3580,N_3021,N_3006);
and U3581 (N_3581,N_3242,N_3070);
nor U3582 (N_3582,N_3187,N_3325);
nor U3583 (N_3583,N_3344,N_3334);
xor U3584 (N_3584,N_3392,N_3332);
and U3585 (N_3585,N_3445,N_3200);
xnor U3586 (N_3586,N_3157,N_3261);
nand U3587 (N_3587,N_3055,N_3472);
nand U3588 (N_3588,N_3411,N_3218);
nand U3589 (N_3589,N_3391,N_3250);
xor U3590 (N_3590,N_3143,N_3289);
and U3591 (N_3591,N_3232,N_3121);
nand U3592 (N_3592,N_3311,N_3210);
and U3593 (N_3593,N_3257,N_3231);
or U3594 (N_3594,N_3026,N_3422);
and U3595 (N_3595,N_3110,N_3307);
or U3596 (N_3596,N_3333,N_3087);
and U3597 (N_3597,N_3040,N_3361);
xor U3598 (N_3598,N_3075,N_3495);
or U3599 (N_3599,N_3038,N_3296);
nor U3600 (N_3600,N_3372,N_3217);
and U3601 (N_3601,N_3024,N_3123);
nand U3602 (N_3602,N_3082,N_3265);
nor U3603 (N_3603,N_3131,N_3116);
or U3604 (N_3604,N_3427,N_3268);
nand U3605 (N_3605,N_3473,N_3329);
and U3606 (N_3606,N_3270,N_3429);
nand U3607 (N_3607,N_3430,N_3245);
xor U3608 (N_3608,N_3314,N_3192);
and U3609 (N_3609,N_3166,N_3362);
nand U3610 (N_3610,N_3396,N_3267);
nand U3611 (N_3611,N_3028,N_3189);
nor U3612 (N_3612,N_3457,N_3486);
or U3613 (N_3613,N_3084,N_3064);
nand U3614 (N_3614,N_3125,N_3211);
or U3615 (N_3615,N_3222,N_3183);
or U3616 (N_3616,N_3016,N_3184);
xor U3617 (N_3617,N_3293,N_3449);
or U3618 (N_3618,N_3012,N_3060);
and U3619 (N_3619,N_3032,N_3182);
nor U3620 (N_3620,N_3295,N_3414);
or U3621 (N_3621,N_3117,N_3199);
nor U3622 (N_3622,N_3080,N_3158);
or U3623 (N_3623,N_3162,N_3277);
and U3624 (N_3624,N_3112,N_3280);
xnor U3625 (N_3625,N_3276,N_3313);
xor U3626 (N_3626,N_3435,N_3374);
nand U3627 (N_3627,N_3089,N_3146);
or U3628 (N_3628,N_3047,N_3056);
and U3629 (N_3629,N_3017,N_3365);
nand U3630 (N_3630,N_3387,N_3364);
and U3631 (N_3631,N_3456,N_3388);
nor U3632 (N_3632,N_3386,N_3008);
and U3633 (N_3633,N_3113,N_3204);
or U3634 (N_3634,N_3244,N_3356);
nand U3635 (N_3635,N_3209,N_3366);
xor U3636 (N_3636,N_3236,N_3390);
xor U3637 (N_3637,N_3345,N_3186);
xor U3638 (N_3638,N_3299,N_3103);
nand U3639 (N_3639,N_3109,N_3191);
and U3640 (N_3640,N_3009,N_3128);
nand U3641 (N_3641,N_3347,N_3163);
or U3642 (N_3642,N_3288,N_3150);
nand U3643 (N_3643,N_3442,N_3248);
nor U3644 (N_3644,N_3448,N_3338);
or U3645 (N_3645,N_3067,N_3174);
xnor U3646 (N_3646,N_3378,N_3165);
or U3647 (N_3647,N_3010,N_3039);
or U3648 (N_3648,N_3133,N_3383);
xnor U3649 (N_3649,N_3152,N_3278);
and U3650 (N_3650,N_3171,N_3352);
nor U3651 (N_3651,N_3247,N_3463);
and U3652 (N_3652,N_3326,N_3106);
or U3653 (N_3653,N_3097,N_3403);
or U3654 (N_3654,N_3019,N_3409);
xnor U3655 (N_3655,N_3286,N_3479);
nor U3656 (N_3656,N_3441,N_3013);
and U3657 (N_3657,N_3193,N_3220);
or U3658 (N_3658,N_3007,N_3041);
or U3659 (N_3659,N_3062,N_3139);
and U3660 (N_3660,N_3090,N_3091);
nand U3661 (N_3661,N_3104,N_3094);
and U3662 (N_3662,N_3137,N_3395);
or U3663 (N_3663,N_3428,N_3443);
nand U3664 (N_3664,N_3072,N_3468);
xnor U3665 (N_3665,N_3469,N_3173);
xnor U3666 (N_3666,N_3086,N_3251);
xnor U3667 (N_3667,N_3418,N_3227);
xnor U3668 (N_3668,N_3035,N_3207);
nor U3669 (N_3669,N_3071,N_3003);
or U3670 (N_3670,N_3337,N_3323);
nor U3671 (N_3671,N_3493,N_3206);
or U3672 (N_3672,N_3042,N_3050);
nand U3673 (N_3673,N_3419,N_3114);
or U3674 (N_3674,N_3384,N_3025);
nor U3675 (N_3675,N_3059,N_3300);
and U3676 (N_3676,N_3298,N_3252);
nand U3677 (N_3677,N_3108,N_3336);
nor U3678 (N_3678,N_3111,N_3389);
nand U3679 (N_3679,N_3068,N_3431);
nand U3680 (N_3680,N_3351,N_3425);
xnor U3681 (N_3681,N_3433,N_3194);
nand U3682 (N_3682,N_3488,N_3412);
nand U3683 (N_3683,N_3263,N_3153);
xnor U3684 (N_3684,N_3476,N_3410);
nor U3685 (N_3685,N_3346,N_3014);
nand U3686 (N_3686,N_3201,N_3499);
nor U3687 (N_3687,N_3376,N_3159);
nand U3688 (N_3688,N_3161,N_3120);
nor U3689 (N_3689,N_3492,N_3360);
or U3690 (N_3690,N_3375,N_3368);
xor U3691 (N_3691,N_3399,N_3136);
xnor U3692 (N_3692,N_3216,N_3275);
nand U3693 (N_3693,N_3471,N_3381);
and U3694 (N_3694,N_3279,N_3497);
and U3695 (N_3695,N_3393,N_3175);
or U3696 (N_3696,N_3377,N_3140);
nand U3697 (N_3697,N_3246,N_3432);
or U3698 (N_3698,N_3309,N_3406);
or U3699 (N_3699,N_3317,N_3291);
nor U3700 (N_3700,N_3370,N_3324);
nor U3701 (N_3701,N_3467,N_3238);
or U3702 (N_3702,N_3233,N_3397);
and U3703 (N_3703,N_3235,N_3444);
nor U3704 (N_3704,N_3451,N_3054);
and U3705 (N_3705,N_3491,N_3373);
and U3706 (N_3706,N_3284,N_3046);
nor U3707 (N_3707,N_3002,N_3147);
and U3708 (N_3708,N_3423,N_3310);
xnor U3709 (N_3709,N_3434,N_3127);
or U3710 (N_3710,N_3359,N_3253);
xnor U3711 (N_3711,N_3302,N_3453);
and U3712 (N_3712,N_3079,N_3135);
nand U3713 (N_3713,N_3160,N_3466);
nand U3714 (N_3714,N_3000,N_3355);
nand U3715 (N_3715,N_3239,N_3405);
xnor U3716 (N_3716,N_3385,N_3195);
nor U3717 (N_3717,N_3401,N_3274);
xor U3718 (N_3718,N_3494,N_3095);
nand U3719 (N_3719,N_3308,N_3320);
and U3720 (N_3720,N_3437,N_3208);
xor U3721 (N_3721,N_3264,N_3318);
nor U3722 (N_3722,N_3101,N_3164);
or U3723 (N_3723,N_3092,N_3126);
or U3724 (N_3724,N_3294,N_3420);
and U3725 (N_3725,N_3156,N_3190);
or U3726 (N_3726,N_3088,N_3339);
and U3727 (N_3727,N_3369,N_3237);
nand U3728 (N_3728,N_3057,N_3176);
or U3729 (N_3729,N_3306,N_3096);
nand U3730 (N_3730,N_3011,N_3319);
nor U3731 (N_3731,N_3022,N_3168);
nand U3732 (N_3732,N_3198,N_3328);
or U3733 (N_3733,N_3454,N_3258);
and U3734 (N_3734,N_3076,N_3436);
or U3735 (N_3735,N_3455,N_3151);
nand U3736 (N_3736,N_3312,N_3132);
nand U3737 (N_3737,N_3081,N_3321);
or U3738 (N_3738,N_3413,N_3287);
xor U3739 (N_3739,N_3269,N_3480);
and U3740 (N_3740,N_3221,N_3341);
xnor U3741 (N_3741,N_3069,N_3283);
and U3742 (N_3742,N_3063,N_3196);
nand U3743 (N_3743,N_3353,N_3343);
nand U3744 (N_3744,N_3249,N_3185);
nor U3745 (N_3745,N_3045,N_3134);
xnor U3746 (N_3746,N_3408,N_3483);
nor U3747 (N_3747,N_3149,N_3475);
nor U3748 (N_3748,N_3315,N_3115);
or U3749 (N_3749,N_3225,N_3402);
and U3750 (N_3750,N_3199,N_3388);
or U3751 (N_3751,N_3272,N_3449);
nor U3752 (N_3752,N_3264,N_3038);
and U3753 (N_3753,N_3264,N_3337);
nand U3754 (N_3754,N_3169,N_3176);
nand U3755 (N_3755,N_3319,N_3211);
nand U3756 (N_3756,N_3120,N_3237);
xnor U3757 (N_3757,N_3022,N_3222);
or U3758 (N_3758,N_3367,N_3260);
xor U3759 (N_3759,N_3312,N_3129);
or U3760 (N_3760,N_3190,N_3191);
or U3761 (N_3761,N_3441,N_3470);
nand U3762 (N_3762,N_3220,N_3468);
nor U3763 (N_3763,N_3278,N_3249);
xnor U3764 (N_3764,N_3449,N_3151);
xor U3765 (N_3765,N_3390,N_3033);
and U3766 (N_3766,N_3081,N_3445);
nor U3767 (N_3767,N_3133,N_3163);
nor U3768 (N_3768,N_3044,N_3336);
nor U3769 (N_3769,N_3496,N_3476);
or U3770 (N_3770,N_3190,N_3276);
or U3771 (N_3771,N_3491,N_3091);
and U3772 (N_3772,N_3161,N_3060);
and U3773 (N_3773,N_3262,N_3460);
or U3774 (N_3774,N_3134,N_3175);
nor U3775 (N_3775,N_3050,N_3019);
nand U3776 (N_3776,N_3061,N_3163);
and U3777 (N_3777,N_3166,N_3210);
and U3778 (N_3778,N_3227,N_3239);
xnor U3779 (N_3779,N_3200,N_3284);
nor U3780 (N_3780,N_3116,N_3408);
nor U3781 (N_3781,N_3113,N_3232);
nand U3782 (N_3782,N_3330,N_3042);
nand U3783 (N_3783,N_3191,N_3179);
xor U3784 (N_3784,N_3066,N_3141);
or U3785 (N_3785,N_3390,N_3102);
nor U3786 (N_3786,N_3191,N_3022);
nor U3787 (N_3787,N_3293,N_3331);
and U3788 (N_3788,N_3103,N_3055);
and U3789 (N_3789,N_3013,N_3307);
nor U3790 (N_3790,N_3294,N_3457);
and U3791 (N_3791,N_3032,N_3417);
nor U3792 (N_3792,N_3407,N_3436);
nand U3793 (N_3793,N_3090,N_3118);
and U3794 (N_3794,N_3104,N_3321);
nand U3795 (N_3795,N_3325,N_3192);
or U3796 (N_3796,N_3183,N_3174);
nor U3797 (N_3797,N_3104,N_3175);
or U3798 (N_3798,N_3032,N_3058);
nand U3799 (N_3799,N_3192,N_3301);
or U3800 (N_3800,N_3049,N_3326);
or U3801 (N_3801,N_3249,N_3498);
xor U3802 (N_3802,N_3478,N_3224);
nor U3803 (N_3803,N_3008,N_3001);
nor U3804 (N_3804,N_3130,N_3418);
xor U3805 (N_3805,N_3117,N_3453);
nand U3806 (N_3806,N_3058,N_3034);
xnor U3807 (N_3807,N_3292,N_3186);
nor U3808 (N_3808,N_3352,N_3246);
nand U3809 (N_3809,N_3251,N_3345);
nand U3810 (N_3810,N_3436,N_3417);
xnor U3811 (N_3811,N_3391,N_3235);
nand U3812 (N_3812,N_3465,N_3215);
or U3813 (N_3813,N_3468,N_3050);
nand U3814 (N_3814,N_3107,N_3456);
and U3815 (N_3815,N_3263,N_3429);
or U3816 (N_3816,N_3312,N_3169);
and U3817 (N_3817,N_3473,N_3076);
xor U3818 (N_3818,N_3442,N_3193);
and U3819 (N_3819,N_3379,N_3479);
xnor U3820 (N_3820,N_3112,N_3275);
nor U3821 (N_3821,N_3005,N_3040);
xor U3822 (N_3822,N_3199,N_3395);
and U3823 (N_3823,N_3438,N_3406);
xor U3824 (N_3824,N_3188,N_3171);
xnor U3825 (N_3825,N_3004,N_3234);
and U3826 (N_3826,N_3309,N_3430);
or U3827 (N_3827,N_3099,N_3493);
or U3828 (N_3828,N_3111,N_3306);
nor U3829 (N_3829,N_3119,N_3062);
xor U3830 (N_3830,N_3357,N_3484);
and U3831 (N_3831,N_3085,N_3390);
and U3832 (N_3832,N_3132,N_3485);
nor U3833 (N_3833,N_3027,N_3150);
nand U3834 (N_3834,N_3344,N_3319);
nand U3835 (N_3835,N_3148,N_3231);
nand U3836 (N_3836,N_3045,N_3174);
and U3837 (N_3837,N_3484,N_3333);
and U3838 (N_3838,N_3268,N_3333);
and U3839 (N_3839,N_3257,N_3197);
xnor U3840 (N_3840,N_3156,N_3408);
and U3841 (N_3841,N_3197,N_3032);
or U3842 (N_3842,N_3391,N_3296);
and U3843 (N_3843,N_3139,N_3209);
nor U3844 (N_3844,N_3176,N_3336);
xor U3845 (N_3845,N_3235,N_3488);
nand U3846 (N_3846,N_3374,N_3020);
or U3847 (N_3847,N_3423,N_3184);
and U3848 (N_3848,N_3321,N_3163);
nand U3849 (N_3849,N_3274,N_3159);
nand U3850 (N_3850,N_3208,N_3337);
xor U3851 (N_3851,N_3480,N_3129);
or U3852 (N_3852,N_3375,N_3020);
or U3853 (N_3853,N_3109,N_3441);
or U3854 (N_3854,N_3356,N_3139);
and U3855 (N_3855,N_3057,N_3000);
xnor U3856 (N_3856,N_3234,N_3016);
or U3857 (N_3857,N_3149,N_3275);
xnor U3858 (N_3858,N_3004,N_3097);
xor U3859 (N_3859,N_3338,N_3489);
and U3860 (N_3860,N_3266,N_3122);
nor U3861 (N_3861,N_3234,N_3427);
xnor U3862 (N_3862,N_3112,N_3327);
or U3863 (N_3863,N_3088,N_3013);
nand U3864 (N_3864,N_3326,N_3083);
and U3865 (N_3865,N_3407,N_3187);
or U3866 (N_3866,N_3382,N_3451);
xnor U3867 (N_3867,N_3437,N_3169);
or U3868 (N_3868,N_3009,N_3013);
nand U3869 (N_3869,N_3264,N_3020);
and U3870 (N_3870,N_3322,N_3335);
and U3871 (N_3871,N_3112,N_3036);
nand U3872 (N_3872,N_3246,N_3296);
xnor U3873 (N_3873,N_3473,N_3478);
nand U3874 (N_3874,N_3197,N_3319);
xor U3875 (N_3875,N_3466,N_3390);
nor U3876 (N_3876,N_3391,N_3339);
xnor U3877 (N_3877,N_3110,N_3191);
nor U3878 (N_3878,N_3235,N_3184);
or U3879 (N_3879,N_3247,N_3455);
xor U3880 (N_3880,N_3398,N_3059);
nand U3881 (N_3881,N_3274,N_3087);
and U3882 (N_3882,N_3010,N_3122);
nor U3883 (N_3883,N_3363,N_3068);
or U3884 (N_3884,N_3401,N_3216);
nor U3885 (N_3885,N_3438,N_3131);
nor U3886 (N_3886,N_3409,N_3467);
xnor U3887 (N_3887,N_3283,N_3353);
nor U3888 (N_3888,N_3104,N_3478);
xor U3889 (N_3889,N_3050,N_3280);
nor U3890 (N_3890,N_3041,N_3100);
xor U3891 (N_3891,N_3078,N_3172);
or U3892 (N_3892,N_3153,N_3439);
nor U3893 (N_3893,N_3440,N_3025);
nor U3894 (N_3894,N_3058,N_3341);
and U3895 (N_3895,N_3341,N_3245);
xor U3896 (N_3896,N_3347,N_3081);
or U3897 (N_3897,N_3266,N_3314);
or U3898 (N_3898,N_3314,N_3337);
nor U3899 (N_3899,N_3009,N_3204);
or U3900 (N_3900,N_3383,N_3440);
or U3901 (N_3901,N_3468,N_3403);
or U3902 (N_3902,N_3469,N_3219);
nand U3903 (N_3903,N_3389,N_3461);
nor U3904 (N_3904,N_3198,N_3316);
and U3905 (N_3905,N_3498,N_3208);
or U3906 (N_3906,N_3266,N_3182);
or U3907 (N_3907,N_3113,N_3022);
nor U3908 (N_3908,N_3395,N_3129);
nor U3909 (N_3909,N_3256,N_3258);
and U3910 (N_3910,N_3027,N_3454);
xor U3911 (N_3911,N_3369,N_3061);
and U3912 (N_3912,N_3061,N_3010);
or U3913 (N_3913,N_3250,N_3386);
and U3914 (N_3914,N_3051,N_3306);
nand U3915 (N_3915,N_3422,N_3366);
xnor U3916 (N_3916,N_3403,N_3495);
nand U3917 (N_3917,N_3028,N_3351);
nor U3918 (N_3918,N_3350,N_3152);
nor U3919 (N_3919,N_3231,N_3065);
and U3920 (N_3920,N_3017,N_3234);
nor U3921 (N_3921,N_3303,N_3334);
xnor U3922 (N_3922,N_3353,N_3079);
nand U3923 (N_3923,N_3339,N_3047);
nand U3924 (N_3924,N_3151,N_3321);
nor U3925 (N_3925,N_3271,N_3395);
xnor U3926 (N_3926,N_3062,N_3291);
nand U3927 (N_3927,N_3430,N_3268);
xnor U3928 (N_3928,N_3011,N_3125);
nor U3929 (N_3929,N_3212,N_3072);
nor U3930 (N_3930,N_3036,N_3392);
or U3931 (N_3931,N_3328,N_3269);
and U3932 (N_3932,N_3195,N_3472);
nand U3933 (N_3933,N_3378,N_3035);
and U3934 (N_3934,N_3246,N_3107);
xnor U3935 (N_3935,N_3129,N_3019);
nor U3936 (N_3936,N_3035,N_3185);
nand U3937 (N_3937,N_3126,N_3498);
xor U3938 (N_3938,N_3473,N_3323);
xnor U3939 (N_3939,N_3015,N_3217);
xor U3940 (N_3940,N_3223,N_3255);
nor U3941 (N_3941,N_3459,N_3447);
nand U3942 (N_3942,N_3208,N_3281);
nor U3943 (N_3943,N_3355,N_3017);
and U3944 (N_3944,N_3160,N_3408);
or U3945 (N_3945,N_3020,N_3134);
and U3946 (N_3946,N_3060,N_3386);
xor U3947 (N_3947,N_3414,N_3087);
xnor U3948 (N_3948,N_3252,N_3214);
and U3949 (N_3949,N_3432,N_3000);
nor U3950 (N_3950,N_3440,N_3397);
nor U3951 (N_3951,N_3039,N_3357);
xor U3952 (N_3952,N_3152,N_3121);
or U3953 (N_3953,N_3288,N_3134);
nand U3954 (N_3954,N_3384,N_3026);
nand U3955 (N_3955,N_3461,N_3387);
or U3956 (N_3956,N_3068,N_3080);
and U3957 (N_3957,N_3294,N_3244);
or U3958 (N_3958,N_3416,N_3106);
nand U3959 (N_3959,N_3340,N_3176);
or U3960 (N_3960,N_3126,N_3394);
or U3961 (N_3961,N_3049,N_3145);
and U3962 (N_3962,N_3324,N_3237);
and U3963 (N_3963,N_3045,N_3453);
nor U3964 (N_3964,N_3318,N_3051);
xor U3965 (N_3965,N_3010,N_3248);
xor U3966 (N_3966,N_3017,N_3016);
or U3967 (N_3967,N_3267,N_3347);
nor U3968 (N_3968,N_3081,N_3306);
xnor U3969 (N_3969,N_3305,N_3398);
nor U3970 (N_3970,N_3158,N_3283);
nor U3971 (N_3971,N_3242,N_3010);
nand U3972 (N_3972,N_3491,N_3413);
or U3973 (N_3973,N_3113,N_3473);
nor U3974 (N_3974,N_3198,N_3265);
nor U3975 (N_3975,N_3368,N_3482);
nand U3976 (N_3976,N_3057,N_3446);
and U3977 (N_3977,N_3468,N_3316);
xnor U3978 (N_3978,N_3091,N_3108);
xnor U3979 (N_3979,N_3022,N_3104);
nand U3980 (N_3980,N_3312,N_3000);
or U3981 (N_3981,N_3197,N_3375);
nand U3982 (N_3982,N_3432,N_3361);
xor U3983 (N_3983,N_3396,N_3452);
nand U3984 (N_3984,N_3335,N_3140);
xor U3985 (N_3985,N_3016,N_3265);
xnor U3986 (N_3986,N_3444,N_3120);
nand U3987 (N_3987,N_3468,N_3216);
xnor U3988 (N_3988,N_3417,N_3203);
nand U3989 (N_3989,N_3175,N_3451);
and U3990 (N_3990,N_3481,N_3332);
xor U3991 (N_3991,N_3111,N_3073);
nor U3992 (N_3992,N_3137,N_3019);
and U3993 (N_3993,N_3472,N_3337);
or U3994 (N_3994,N_3396,N_3163);
or U3995 (N_3995,N_3327,N_3352);
xor U3996 (N_3996,N_3462,N_3210);
and U3997 (N_3997,N_3425,N_3309);
xor U3998 (N_3998,N_3052,N_3153);
nor U3999 (N_3999,N_3356,N_3430);
nand U4000 (N_4000,N_3651,N_3637);
and U4001 (N_4001,N_3760,N_3512);
and U4002 (N_4002,N_3865,N_3577);
nand U4003 (N_4003,N_3665,N_3900);
or U4004 (N_4004,N_3714,N_3984);
nand U4005 (N_4005,N_3841,N_3957);
and U4006 (N_4006,N_3664,N_3945);
and U4007 (N_4007,N_3517,N_3772);
nand U4008 (N_4008,N_3639,N_3548);
xnor U4009 (N_4009,N_3968,N_3778);
or U4010 (N_4010,N_3764,N_3542);
nand U4011 (N_4011,N_3614,N_3634);
nor U4012 (N_4012,N_3619,N_3555);
xor U4013 (N_4013,N_3518,N_3708);
xor U4014 (N_4014,N_3556,N_3944);
and U4015 (N_4015,N_3888,N_3844);
nand U4016 (N_4016,N_3591,N_3845);
and U4017 (N_4017,N_3616,N_3740);
and U4018 (N_4018,N_3713,N_3513);
or U4019 (N_4019,N_3824,N_3729);
nor U4020 (N_4020,N_3843,N_3890);
nor U4021 (N_4021,N_3802,N_3661);
nor U4022 (N_4022,N_3747,N_3910);
and U4023 (N_4023,N_3682,N_3730);
or U4024 (N_4024,N_3724,N_3981);
xor U4025 (N_4025,N_3562,N_3757);
or U4026 (N_4026,N_3761,N_3970);
or U4027 (N_4027,N_3705,N_3679);
nand U4028 (N_4028,N_3956,N_3967);
nor U4029 (N_4029,N_3774,N_3864);
nor U4030 (N_4030,N_3754,N_3991);
xnor U4031 (N_4031,N_3509,N_3744);
and U4032 (N_4032,N_3553,N_3539);
or U4033 (N_4033,N_3883,N_3769);
xor U4034 (N_4034,N_3923,N_3942);
nor U4035 (N_4035,N_3918,N_3534);
and U4036 (N_4036,N_3521,N_3540);
xor U4037 (N_4037,N_3693,N_3969);
nand U4038 (N_4038,N_3771,N_3830);
nand U4039 (N_4039,N_3554,N_3601);
nor U4040 (N_4040,N_3605,N_3751);
and U4041 (N_4041,N_3979,N_3993);
nor U4042 (N_4042,N_3711,N_3798);
nor U4043 (N_4043,N_3878,N_3580);
xor U4044 (N_4044,N_3782,N_3907);
or U4045 (N_4045,N_3533,N_3795);
nor U4046 (N_4046,N_3797,N_3777);
xnor U4047 (N_4047,N_3791,N_3612);
and U4048 (N_4048,N_3541,N_3831);
nor U4049 (N_4049,N_3884,N_3671);
xor U4050 (N_4050,N_3635,N_3698);
xnor U4051 (N_4051,N_3893,N_3881);
nor U4052 (N_4052,N_3745,N_3620);
and U4053 (N_4053,N_3852,N_3550);
and U4054 (N_4054,N_3858,N_3525);
nand U4055 (N_4055,N_3887,N_3712);
nor U4056 (N_4056,N_3787,N_3994);
nor U4057 (N_4057,N_3899,N_3790);
xnor U4058 (N_4058,N_3966,N_3765);
nor U4059 (N_4059,N_3578,N_3853);
nand U4060 (N_4060,N_3935,N_3558);
or U4061 (N_4061,N_3583,N_3503);
or U4062 (N_4062,N_3847,N_3707);
nor U4063 (N_4063,N_3709,N_3644);
nor U4064 (N_4064,N_3625,N_3850);
and U4065 (N_4065,N_3784,N_3736);
nand U4066 (N_4066,N_3986,N_3996);
nor U4067 (N_4067,N_3877,N_3546);
xnor U4068 (N_4068,N_3652,N_3813);
xnor U4069 (N_4069,N_3950,N_3727);
or U4070 (N_4070,N_3506,N_3911);
and U4071 (N_4071,N_3770,N_3628);
nor U4072 (N_4072,N_3607,N_3721);
xor U4073 (N_4073,N_3621,N_3660);
xnor U4074 (N_4074,N_3814,N_3516);
xnor U4075 (N_4075,N_3735,N_3692);
or U4076 (N_4076,N_3915,N_3722);
xnor U4077 (N_4077,N_3929,N_3866);
nand U4078 (N_4078,N_3786,N_3524);
and U4079 (N_4079,N_3897,N_3759);
xnor U4080 (N_4080,N_3650,N_3896);
nand U4081 (N_4081,N_3543,N_3574);
and U4082 (N_4082,N_3928,N_3653);
nor U4083 (N_4083,N_3582,N_3839);
nor U4084 (N_4084,N_3906,N_3973);
xnor U4085 (N_4085,N_3646,N_3891);
xor U4086 (N_4086,N_3701,N_3666);
xnor U4087 (N_4087,N_3686,N_3796);
nor U4088 (N_4088,N_3610,N_3719);
or U4089 (N_4089,N_3976,N_3752);
and U4090 (N_4090,N_3763,N_3528);
nor U4091 (N_4091,N_3717,N_3547);
nor U4092 (N_4092,N_3954,N_3939);
or U4093 (N_4093,N_3862,N_3781);
nand U4094 (N_4094,N_3859,N_3678);
nand U4095 (N_4095,N_3659,N_3643);
nor U4096 (N_4096,N_3773,N_3598);
xnor U4097 (N_4097,N_3927,N_3860);
xnor U4098 (N_4098,N_3718,N_3875);
nor U4099 (N_4099,N_3749,N_3848);
xor U4100 (N_4100,N_3572,N_3785);
or U4101 (N_4101,N_3609,N_3811);
xnor U4102 (N_4102,N_3756,N_3871);
or U4103 (N_4103,N_3593,N_3567);
or U4104 (N_4104,N_3579,N_3780);
nor U4105 (N_4105,N_3733,N_3599);
xnor U4106 (N_4106,N_3842,N_3670);
or U4107 (N_4107,N_3673,N_3552);
or U4108 (N_4108,N_3913,N_3854);
xor U4109 (N_4109,N_3622,N_3948);
nand U4110 (N_4110,N_3560,N_3975);
or U4111 (N_4111,N_3849,N_3985);
nand U4112 (N_4112,N_3965,N_3504);
nor U4113 (N_4113,N_3964,N_3949);
xor U4114 (N_4114,N_3640,N_3545);
xnor U4115 (N_4115,N_3641,N_3783);
nand U4116 (N_4116,N_3603,N_3731);
or U4117 (N_4117,N_3632,N_3508);
nor U4118 (N_4118,N_3909,N_3825);
nand U4119 (N_4119,N_3867,N_3951);
nand U4120 (N_4120,N_3595,N_3629);
nand U4121 (N_4121,N_3675,N_3930);
or U4122 (N_4122,N_3726,N_3648);
nand U4123 (N_4123,N_3514,N_3691);
or U4124 (N_4124,N_3532,N_3974);
nor U4125 (N_4125,N_3647,N_3633);
xnor U4126 (N_4126,N_3924,N_3645);
and U4127 (N_4127,N_3688,N_3999);
and U4128 (N_4128,N_3987,N_3669);
or U4129 (N_4129,N_3794,N_3902);
or U4130 (N_4130,N_3998,N_3596);
nand U4131 (N_4131,N_3627,N_3992);
nor U4132 (N_4132,N_3615,N_3803);
nand U4133 (N_4133,N_3857,N_3505);
nor U4134 (N_4134,N_3748,N_3584);
nor U4135 (N_4135,N_3549,N_3919);
xor U4136 (N_4136,N_3820,N_3557);
or U4137 (N_4137,N_3630,N_3868);
or U4138 (N_4138,N_3958,N_3668);
xor U4139 (N_4139,N_3566,N_3683);
or U4140 (N_4140,N_3728,N_3575);
nor U4141 (N_4141,N_3916,N_3922);
or U4142 (N_4142,N_3624,N_3704);
nand U4143 (N_4143,N_3846,N_3905);
and U4144 (N_4144,N_3551,N_3872);
nor U4145 (N_4145,N_3940,N_3920);
or U4146 (N_4146,N_3758,N_3716);
and U4147 (N_4147,N_3835,N_3507);
and U4148 (N_4148,N_3815,N_3779);
xor U4149 (N_4149,N_3816,N_3606);
nand U4150 (N_4150,N_3530,N_3720);
nor U4151 (N_4151,N_3943,N_3952);
nor U4152 (N_4152,N_3626,N_3953);
nand U4153 (N_4153,N_3990,N_3880);
nand U4154 (N_4154,N_3834,N_3959);
and U4155 (N_4155,N_3822,N_3826);
nand U4156 (N_4156,N_3873,N_3725);
or U4157 (N_4157,N_3510,N_3978);
and U4158 (N_4158,N_3617,N_3925);
or U4159 (N_4159,N_3995,N_3870);
nor U4160 (N_4160,N_3819,N_3611);
or U4161 (N_4161,N_3537,N_3804);
and U4162 (N_4162,N_3904,N_3502);
nor U4163 (N_4163,N_3702,N_3676);
nor U4164 (N_4164,N_3960,N_3618);
and U4165 (N_4165,N_3587,N_3898);
nor U4166 (N_4166,N_3856,N_3519);
or U4167 (N_4167,N_3674,N_3569);
and U4168 (N_4168,N_3501,N_3544);
and U4169 (N_4169,N_3932,N_3564);
nand U4170 (N_4170,N_3585,N_3963);
nor U4171 (N_4171,N_3838,N_3917);
and U4172 (N_4172,N_3573,N_3961);
xor U4173 (N_4173,N_3775,N_3699);
and U4174 (N_4174,N_3654,N_3613);
and U4175 (N_4175,N_3895,N_3527);
and U4176 (N_4176,N_3738,N_3586);
or U4177 (N_4177,N_3807,N_3962);
xor U4178 (N_4178,N_3511,N_3946);
nand U4179 (N_4179,N_3536,N_3982);
or U4180 (N_4180,N_3636,N_3734);
xnor U4181 (N_4181,N_3746,N_3840);
or U4182 (N_4182,N_3980,N_3837);
nor U4183 (N_4183,N_3529,N_3655);
xnor U4184 (N_4184,N_3667,N_3715);
xor U4185 (N_4185,N_3855,N_3677);
nand U4186 (N_4186,N_3874,N_3885);
or U4187 (N_4187,N_3823,N_3672);
or U4188 (N_4188,N_3828,N_3531);
nor U4189 (N_4189,N_3684,N_3515);
nor U4190 (N_4190,N_3908,N_3933);
and U4191 (N_4191,N_3812,N_3810);
or U4192 (N_4192,N_3914,N_3649);
xor U4193 (N_4193,N_3590,N_3568);
and U4194 (N_4194,N_3894,N_3800);
and U4195 (N_4195,N_3520,N_3861);
nor U4196 (N_4196,N_3921,N_3631);
nor U4197 (N_4197,N_3638,N_3694);
nand U4198 (N_4198,N_3788,N_3805);
or U4199 (N_4199,N_3836,N_3589);
xor U4200 (N_4200,N_3817,N_3681);
or U4201 (N_4201,N_3696,N_3931);
and U4202 (N_4202,N_3879,N_3806);
nor U4203 (N_4203,N_3588,N_3869);
nand U4204 (N_4204,N_3592,N_3741);
or U4205 (N_4205,N_3889,N_3808);
and U4206 (N_4206,N_3882,N_3821);
xnor U4207 (N_4207,N_3912,N_3656);
xnor U4208 (N_4208,N_3623,N_3706);
xnor U4209 (N_4209,N_3977,N_3742);
nand U4210 (N_4210,N_3657,N_3755);
or U4211 (N_4211,N_3818,N_3739);
and U4212 (N_4212,N_3594,N_3901);
nand U4213 (N_4213,N_3988,N_3851);
nand U4214 (N_4214,N_3535,N_3576);
and U4215 (N_4215,N_3743,N_3829);
xor U4216 (N_4216,N_3832,N_3685);
or U4217 (N_4217,N_3767,N_3642);
and U4218 (N_4218,N_3700,N_3941);
xor U4219 (N_4219,N_3997,N_3792);
nor U4220 (N_4220,N_3753,N_3971);
or U4221 (N_4221,N_3600,N_3737);
nand U4222 (N_4222,N_3695,N_3523);
or U4223 (N_4223,N_3947,N_3934);
and U4224 (N_4224,N_3662,N_3723);
or U4225 (N_4225,N_3559,N_3697);
or U4226 (N_4226,N_3563,N_3689);
or U4227 (N_4227,N_3799,N_3571);
and U4228 (N_4228,N_3762,N_3768);
and U4229 (N_4229,N_3538,N_3500);
or U4230 (N_4230,N_3863,N_3827);
nand U4231 (N_4231,N_3732,N_3972);
xor U4232 (N_4232,N_3597,N_3710);
xor U4233 (N_4233,N_3581,N_3604);
and U4234 (N_4234,N_3886,N_3833);
xor U4235 (N_4235,N_3687,N_3776);
xnor U4236 (N_4236,N_3522,N_3602);
xor U4237 (N_4237,N_3703,N_3766);
nand U4238 (N_4238,N_3680,N_3983);
nor U4239 (N_4239,N_3570,N_3955);
or U4240 (N_4240,N_3793,N_3989);
nand U4241 (N_4241,N_3892,N_3809);
and U4242 (N_4242,N_3658,N_3876);
or U4243 (N_4243,N_3608,N_3750);
nand U4244 (N_4244,N_3789,N_3690);
or U4245 (N_4245,N_3938,N_3561);
nor U4246 (N_4246,N_3663,N_3565);
nor U4247 (N_4247,N_3937,N_3903);
nand U4248 (N_4248,N_3801,N_3526);
nor U4249 (N_4249,N_3926,N_3936);
nor U4250 (N_4250,N_3775,N_3908);
and U4251 (N_4251,N_3571,N_3827);
nand U4252 (N_4252,N_3946,N_3880);
nor U4253 (N_4253,N_3845,N_3933);
nor U4254 (N_4254,N_3600,N_3538);
and U4255 (N_4255,N_3535,N_3598);
nor U4256 (N_4256,N_3911,N_3874);
and U4257 (N_4257,N_3545,N_3960);
and U4258 (N_4258,N_3776,N_3823);
nand U4259 (N_4259,N_3700,N_3972);
or U4260 (N_4260,N_3720,N_3999);
nand U4261 (N_4261,N_3624,N_3785);
nand U4262 (N_4262,N_3605,N_3786);
or U4263 (N_4263,N_3860,N_3843);
xor U4264 (N_4264,N_3892,N_3580);
nand U4265 (N_4265,N_3989,N_3867);
nand U4266 (N_4266,N_3935,N_3933);
nor U4267 (N_4267,N_3684,N_3930);
and U4268 (N_4268,N_3884,N_3748);
nor U4269 (N_4269,N_3509,N_3712);
and U4270 (N_4270,N_3515,N_3911);
or U4271 (N_4271,N_3548,N_3609);
and U4272 (N_4272,N_3754,N_3690);
nor U4273 (N_4273,N_3779,N_3884);
nand U4274 (N_4274,N_3620,N_3529);
and U4275 (N_4275,N_3900,N_3656);
xor U4276 (N_4276,N_3765,N_3800);
and U4277 (N_4277,N_3979,N_3962);
nand U4278 (N_4278,N_3761,N_3784);
or U4279 (N_4279,N_3739,N_3873);
and U4280 (N_4280,N_3914,N_3770);
and U4281 (N_4281,N_3741,N_3964);
and U4282 (N_4282,N_3838,N_3958);
nor U4283 (N_4283,N_3691,N_3894);
nor U4284 (N_4284,N_3561,N_3681);
nand U4285 (N_4285,N_3607,N_3674);
nand U4286 (N_4286,N_3578,N_3986);
nor U4287 (N_4287,N_3508,N_3929);
and U4288 (N_4288,N_3644,N_3624);
or U4289 (N_4289,N_3870,N_3801);
nor U4290 (N_4290,N_3551,N_3661);
and U4291 (N_4291,N_3917,N_3550);
nand U4292 (N_4292,N_3521,N_3620);
or U4293 (N_4293,N_3946,N_3594);
or U4294 (N_4294,N_3974,N_3840);
nand U4295 (N_4295,N_3505,N_3519);
and U4296 (N_4296,N_3785,N_3936);
nor U4297 (N_4297,N_3694,N_3788);
nand U4298 (N_4298,N_3778,N_3962);
and U4299 (N_4299,N_3503,N_3608);
xnor U4300 (N_4300,N_3526,N_3983);
and U4301 (N_4301,N_3709,N_3968);
xnor U4302 (N_4302,N_3737,N_3552);
xnor U4303 (N_4303,N_3722,N_3654);
nor U4304 (N_4304,N_3696,N_3778);
xor U4305 (N_4305,N_3850,N_3729);
nor U4306 (N_4306,N_3670,N_3644);
xor U4307 (N_4307,N_3856,N_3654);
or U4308 (N_4308,N_3645,N_3880);
nor U4309 (N_4309,N_3717,N_3647);
nor U4310 (N_4310,N_3532,N_3733);
xor U4311 (N_4311,N_3573,N_3921);
or U4312 (N_4312,N_3803,N_3863);
xor U4313 (N_4313,N_3560,N_3874);
and U4314 (N_4314,N_3705,N_3518);
or U4315 (N_4315,N_3871,N_3697);
and U4316 (N_4316,N_3995,N_3883);
xnor U4317 (N_4317,N_3974,N_3748);
and U4318 (N_4318,N_3591,N_3873);
or U4319 (N_4319,N_3799,N_3995);
nor U4320 (N_4320,N_3729,N_3631);
nand U4321 (N_4321,N_3785,N_3858);
or U4322 (N_4322,N_3938,N_3632);
and U4323 (N_4323,N_3791,N_3893);
nor U4324 (N_4324,N_3542,N_3886);
and U4325 (N_4325,N_3565,N_3609);
and U4326 (N_4326,N_3749,N_3824);
or U4327 (N_4327,N_3843,N_3751);
or U4328 (N_4328,N_3546,N_3586);
nor U4329 (N_4329,N_3756,N_3787);
xor U4330 (N_4330,N_3654,N_3828);
and U4331 (N_4331,N_3806,N_3777);
or U4332 (N_4332,N_3918,N_3684);
xnor U4333 (N_4333,N_3998,N_3768);
xor U4334 (N_4334,N_3528,N_3564);
xor U4335 (N_4335,N_3568,N_3617);
and U4336 (N_4336,N_3599,N_3875);
or U4337 (N_4337,N_3569,N_3648);
xnor U4338 (N_4338,N_3933,N_3872);
or U4339 (N_4339,N_3952,N_3923);
nand U4340 (N_4340,N_3647,N_3547);
or U4341 (N_4341,N_3964,N_3553);
nor U4342 (N_4342,N_3861,N_3828);
nand U4343 (N_4343,N_3872,N_3944);
nor U4344 (N_4344,N_3855,N_3956);
and U4345 (N_4345,N_3679,N_3693);
xnor U4346 (N_4346,N_3679,N_3636);
nand U4347 (N_4347,N_3951,N_3553);
xnor U4348 (N_4348,N_3804,N_3846);
or U4349 (N_4349,N_3549,N_3757);
nor U4350 (N_4350,N_3747,N_3568);
nand U4351 (N_4351,N_3740,N_3647);
nor U4352 (N_4352,N_3757,N_3659);
nor U4353 (N_4353,N_3816,N_3522);
and U4354 (N_4354,N_3551,N_3910);
or U4355 (N_4355,N_3831,N_3926);
xnor U4356 (N_4356,N_3960,N_3752);
nand U4357 (N_4357,N_3507,N_3786);
nor U4358 (N_4358,N_3861,N_3913);
and U4359 (N_4359,N_3832,N_3817);
xor U4360 (N_4360,N_3546,N_3593);
or U4361 (N_4361,N_3836,N_3967);
and U4362 (N_4362,N_3593,N_3667);
and U4363 (N_4363,N_3902,N_3885);
and U4364 (N_4364,N_3770,N_3708);
nand U4365 (N_4365,N_3888,N_3841);
or U4366 (N_4366,N_3683,N_3632);
nand U4367 (N_4367,N_3857,N_3980);
nor U4368 (N_4368,N_3652,N_3860);
nand U4369 (N_4369,N_3986,N_3744);
nand U4370 (N_4370,N_3652,N_3782);
xor U4371 (N_4371,N_3997,N_3844);
nand U4372 (N_4372,N_3909,N_3578);
nor U4373 (N_4373,N_3648,N_3822);
nor U4374 (N_4374,N_3662,N_3978);
nand U4375 (N_4375,N_3719,N_3893);
or U4376 (N_4376,N_3767,N_3922);
nor U4377 (N_4377,N_3791,N_3535);
nand U4378 (N_4378,N_3575,N_3857);
nor U4379 (N_4379,N_3567,N_3653);
or U4380 (N_4380,N_3960,N_3903);
or U4381 (N_4381,N_3708,N_3543);
nand U4382 (N_4382,N_3949,N_3563);
or U4383 (N_4383,N_3675,N_3927);
xor U4384 (N_4384,N_3697,N_3577);
nand U4385 (N_4385,N_3564,N_3560);
nor U4386 (N_4386,N_3789,N_3860);
nand U4387 (N_4387,N_3709,N_3563);
nand U4388 (N_4388,N_3884,N_3592);
or U4389 (N_4389,N_3823,N_3554);
or U4390 (N_4390,N_3627,N_3868);
nand U4391 (N_4391,N_3710,N_3887);
or U4392 (N_4392,N_3977,N_3953);
nor U4393 (N_4393,N_3629,N_3879);
xnor U4394 (N_4394,N_3971,N_3900);
nand U4395 (N_4395,N_3680,N_3622);
nand U4396 (N_4396,N_3866,N_3959);
xnor U4397 (N_4397,N_3539,N_3920);
nand U4398 (N_4398,N_3838,N_3711);
nor U4399 (N_4399,N_3815,N_3836);
xnor U4400 (N_4400,N_3766,N_3568);
xnor U4401 (N_4401,N_3562,N_3972);
xnor U4402 (N_4402,N_3554,N_3691);
nand U4403 (N_4403,N_3622,N_3725);
xor U4404 (N_4404,N_3768,N_3836);
xor U4405 (N_4405,N_3680,N_3929);
and U4406 (N_4406,N_3989,N_3838);
or U4407 (N_4407,N_3645,N_3543);
nor U4408 (N_4408,N_3571,N_3672);
xnor U4409 (N_4409,N_3529,N_3959);
nor U4410 (N_4410,N_3537,N_3615);
nor U4411 (N_4411,N_3709,N_3768);
nor U4412 (N_4412,N_3993,N_3719);
nand U4413 (N_4413,N_3734,N_3514);
or U4414 (N_4414,N_3678,N_3881);
xnor U4415 (N_4415,N_3576,N_3682);
nor U4416 (N_4416,N_3748,N_3674);
nor U4417 (N_4417,N_3716,N_3753);
nand U4418 (N_4418,N_3842,N_3935);
or U4419 (N_4419,N_3987,N_3597);
and U4420 (N_4420,N_3624,N_3734);
or U4421 (N_4421,N_3629,N_3769);
nand U4422 (N_4422,N_3624,N_3899);
nor U4423 (N_4423,N_3932,N_3820);
xnor U4424 (N_4424,N_3760,N_3851);
xnor U4425 (N_4425,N_3877,N_3613);
xnor U4426 (N_4426,N_3546,N_3515);
or U4427 (N_4427,N_3562,N_3591);
nand U4428 (N_4428,N_3722,N_3560);
xor U4429 (N_4429,N_3756,N_3966);
and U4430 (N_4430,N_3607,N_3783);
or U4431 (N_4431,N_3644,N_3727);
and U4432 (N_4432,N_3877,N_3878);
nor U4433 (N_4433,N_3870,N_3662);
nand U4434 (N_4434,N_3965,N_3627);
nor U4435 (N_4435,N_3887,N_3992);
and U4436 (N_4436,N_3959,N_3760);
nand U4437 (N_4437,N_3849,N_3896);
and U4438 (N_4438,N_3960,N_3731);
and U4439 (N_4439,N_3504,N_3717);
nor U4440 (N_4440,N_3706,N_3990);
and U4441 (N_4441,N_3952,N_3893);
or U4442 (N_4442,N_3950,N_3925);
nand U4443 (N_4443,N_3877,N_3717);
xnor U4444 (N_4444,N_3805,N_3791);
nand U4445 (N_4445,N_3501,N_3537);
nand U4446 (N_4446,N_3895,N_3640);
or U4447 (N_4447,N_3643,N_3962);
xnor U4448 (N_4448,N_3532,N_3527);
xor U4449 (N_4449,N_3856,N_3768);
nand U4450 (N_4450,N_3897,N_3560);
nor U4451 (N_4451,N_3905,N_3765);
nand U4452 (N_4452,N_3696,N_3651);
xnor U4453 (N_4453,N_3628,N_3658);
or U4454 (N_4454,N_3937,N_3560);
nand U4455 (N_4455,N_3864,N_3685);
nand U4456 (N_4456,N_3770,N_3832);
nor U4457 (N_4457,N_3647,N_3905);
and U4458 (N_4458,N_3630,N_3607);
nor U4459 (N_4459,N_3958,N_3600);
or U4460 (N_4460,N_3577,N_3715);
nor U4461 (N_4461,N_3602,N_3540);
nand U4462 (N_4462,N_3999,N_3749);
nor U4463 (N_4463,N_3939,N_3642);
nor U4464 (N_4464,N_3787,N_3912);
and U4465 (N_4465,N_3552,N_3622);
nand U4466 (N_4466,N_3699,N_3872);
xor U4467 (N_4467,N_3619,N_3796);
nand U4468 (N_4468,N_3971,N_3623);
or U4469 (N_4469,N_3877,N_3501);
xnor U4470 (N_4470,N_3988,N_3938);
or U4471 (N_4471,N_3721,N_3678);
xnor U4472 (N_4472,N_3580,N_3916);
and U4473 (N_4473,N_3642,N_3870);
and U4474 (N_4474,N_3501,N_3801);
xor U4475 (N_4475,N_3815,N_3564);
nand U4476 (N_4476,N_3838,N_3667);
nor U4477 (N_4477,N_3710,N_3671);
xor U4478 (N_4478,N_3829,N_3802);
xnor U4479 (N_4479,N_3776,N_3789);
and U4480 (N_4480,N_3587,N_3669);
xnor U4481 (N_4481,N_3654,N_3927);
nand U4482 (N_4482,N_3990,N_3978);
xnor U4483 (N_4483,N_3672,N_3643);
xor U4484 (N_4484,N_3698,N_3536);
nand U4485 (N_4485,N_3966,N_3619);
nor U4486 (N_4486,N_3668,N_3622);
or U4487 (N_4487,N_3649,N_3913);
xor U4488 (N_4488,N_3971,N_3844);
or U4489 (N_4489,N_3631,N_3693);
nor U4490 (N_4490,N_3927,N_3717);
nor U4491 (N_4491,N_3580,N_3610);
xnor U4492 (N_4492,N_3546,N_3780);
nand U4493 (N_4493,N_3913,N_3552);
or U4494 (N_4494,N_3742,N_3913);
xnor U4495 (N_4495,N_3700,N_3887);
nand U4496 (N_4496,N_3653,N_3977);
or U4497 (N_4497,N_3734,N_3515);
xor U4498 (N_4498,N_3933,N_3733);
and U4499 (N_4499,N_3845,N_3749);
nand U4500 (N_4500,N_4055,N_4275);
or U4501 (N_4501,N_4145,N_4278);
xnor U4502 (N_4502,N_4262,N_4343);
nor U4503 (N_4503,N_4070,N_4164);
and U4504 (N_4504,N_4191,N_4288);
nor U4505 (N_4505,N_4381,N_4113);
or U4506 (N_4506,N_4233,N_4356);
or U4507 (N_4507,N_4468,N_4122);
xor U4508 (N_4508,N_4427,N_4230);
and U4509 (N_4509,N_4342,N_4413);
xor U4510 (N_4510,N_4081,N_4102);
and U4511 (N_4511,N_4240,N_4041);
xor U4512 (N_4512,N_4495,N_4267);
and U4513 (N_4513,N_4117,N_4260);
nand U4514 (N_4514,N_4083,N_4310);
nand U4515 (N_4515,N_4486,N_4076);
nand U4516 (N_4516,N_4211,N_4048);
nand U4517 (N_4517,N_4300,N_4163);
nand U4518 (N_4518,N_4058,N_4247);
or U4519 (N_4519,N_4183,N_4021);
nor U4520 (N_4520,N_4092,N_4454);
and U4521 (N_4521,N_4185,N_4440);
nand U4522 (N_4522,N_4303,N_4474);
xor U4523 (N_4523,N_4393,N_4143);
nand U4524 (N_4524,N_4098,N_4000);
or U4525 (N_4525,N_4232,N_4036);
nor U4526 (N_4526,N_4341,N_4057);
and U4527 (N_4527,N_4366,N_4004);
or U4528 (N_4528,N_4124,N_4373);
nor U4529 (N_4529,N_4101,N_4200);
nor U4530 (N_4530,N_4475,N_4008);
or U4531 (N_4531,N_4479,N_4452);
nor U4532 (N_4532,N_4089,N_4001);
nor U4533 (N_4533,N_4248,N_4223);
and U4534 (N_4534,N_4269,N_4388);
nor U4535 (N_4535,N_4321,N_4244);
nand U4536 (N_4536,N_4157,N_4481);
nor U4537 (N_4537,N_4390,N_4289);
xnor U4538 (N_4538,N_4075,N_4238);
nor U4539 (N_4539,N_4405,N_4144);
nand U4540 (N_4540,N_4359,N_4497);
nand U4541 (N_4541,N_4068,N_4125);
or U4542 (N_4542,N_4088,N_4190);
or U4543 (N_4543,N_4199,N_4298);
and U4544 (N_4544,N_4167,N_4226);
or U4545 (N_4545,N_4436,N_4069);
nand U4546 (N_4546,N_4496,N_4177);
xor U4547 (N_4547,N_4470,N_4014);
or U4548 (N_4548,N_4133,N_4423);
and U4549 (N_4549,N_4108,N_4439);
xor U4550 (N_4550,N_4027,N_4264);
nand U4551 (N_4551,N_4192,N_4123);
nor U4552 (N_4552,N_4339,N_4246);
or U4553 (N_4553,N_4332,N_4302);
and U4554 (N_4554,N_4139,N_4499);
or U4555 (N_4555,N_4309,N_4446);
xnor U4556 (N_4556,N_4445,N_4361);
or U4557 (N_4557,N_4112,N_4448);
xnor U4558 (N_4558,N_4324,N_4184);
nand U4559 (N_4559,N_4030,N_4311);
xor U4560 (N_4560,N_4338,N_4253);
xor U4561 (N_4561,N_4484,N_4241);
xnor U4562 (N_4562,N_4046,N_4400);
and U4563 (N_4563,N_4319,N_4451);
and U4564 (N_4564,N_4255,N_4480);
xor U4565 (N_4565,N_4268,N_4315);
or U4566 (N_4566,N_4426,N_4419);
nor U4567 (N_4567,N_4009,N_4152);
nand U4568 (N_4568,N_4354,N_4358);
or U4569 (N_4569,N_4418,N_4159);
or U4570 (N_4570,N_4179,N_4257);
nor U4571 (N_4571,N_4172,N_4218);
nor U4572 (N_4572,N_4103,N_4034);
or U4573 (N_4573,N_4097,N_4111);
and U4574 (N_4574,N_4044,N_4146);
and U4575 (N_4575,N_4442,N_4029);
nor U4576 (N_4576,N_4379,N_4051);
or U4577 (N_4577,N_4265,N_4417);
nand U4578 (N_4578,N_4369,N_4209);
nand U4579 (N_4579,N_4433,N_4035);
nand U4580 (N_4580,N_4437,N_4326);
nand U4581 (N_4581,N_4422,N_4162);
xor U4582 (N_4582,N_4498,N_4357);
and U4583 (N_4583,N_4472,N_4126);
and U4584 (N_4584,N_4449,N_4372);
xnor U4585 (N_4585,N_4205,N_4220);
nand U4586 (N_4586,N_4488,N_4476);
nor U4587 (N_4587,N_4313,N_4494);
or U4588 (N_4588,N_4424,N_4182);
xor U4589 (N_4589,N_4091,N_4224);
and U4590 (N_4590,N_4028,N_4147);
xor U4591 (N_4591,N_4401,N_4158);
nand U4592 (N_4592,N_4397,N_4296);
nand U4593 (N_4593,N_4493,N_4186);
and U4594 (N_4594,N_4064,N_4148);
nor U4595 (N_4595,N_4382,N_4049);
nand U4596 (N_4596,N_4120,N_4322);
nor U4597 (N_4597,N_4037,N_4385);
xor U4598 (N_4598,N_4271,N_4453);
or U4599 (N_4599,N_4237,N_4295);
xor U4600 (N_4600,N_4461,N_4290);
nor U4601 (N_4601,N_4215,N_4208);
xor U4602 (N_4602,N_4250,N_4165);
nand U4603 (N_4603,N_4325,N_4022);
nand U4604 (N_4604,N_4273,N_4207);
nand U4605 (N_4605,N_4198,N_4348);
nand U4606 (N_4606,N_4406,N_4175);
nand U4607 (N_4607,N_4317,N_4377);
xor U4608 (N_4608,N_4414,N_4378);
nand U4609 (N_4609,N_4438,N_4093);
nand U4610 (N_4610,N_4299,N_4084);
nand U4611 (N_4611,N_4181,N_4193);
nand U4612 (N_4612,N_4380,N_4040);
and U4613 (N_4613,N_4056,N_4428);
nand U4614 (N_4614,N_4478,N_4180);
or U4615 (N_4615,N_4333,N_4196);
and U4616 (N_4616,N_4314,N_4032);
nand U4617 (N_4617,N_4285,N_4217);
or U4618 (N_4618,N_4294,N_4121);
nor U4619 (N_4619,N_4258,N_4487);
nor U4620 (N_4620,N_4119,N_4411);
xnor U4621 (N_4621,N_4304,N_4047);
nor U4622 (N_4622,N_4160,N_4327);
nand U4623 (N_4623,N_4187,N_4371);
and U4624 (N_4624,N_4308,N_4429);
or U4625 (N_4625,N_4151,N_4012);
or U4626 (N_4626,N_4225,N_4463);
xor U4627 (N_4627,N_4039,N_4394);
and U4628 (N_4628,N_4020,N_4024);
xor U4629 (N_4629,N_4079,N_4231);
or U4630 (N_4630,N_4128,N_4249);
or U4631 (N_4631,N_4455,N_4099);
nand U4632 (N_4632,N_4153,N_4087);
nor U4633 (N_4633,N_4259,N_4293);
or U4634 (N_4634,N_4245,N_4490);
nor U4635 (N_4635,N_4432,N_4360);
xnor U4636 (N_4636,N_4067,N_4396);
or U4637 (N_4637,N_4280,N_4168);
and U4638 (N_4638,N_4483,N_4082);
xnor U4639 (N_4639,N_4078,N_4077);
nand U4640 (N_4640,N_4235,N_4210);
and U4641 (N_4641,N_4323,N_4297);
or U4642 (N_4642,N_4467,N_4094);
and U4643 (N_4643,N_4431,N_4462);
xor U4644 (N_4644,N_4015,N_4085);
or U4645 (N_4645,N_4005,N_4450);
xor U4646 (N_4646,N_4243,N_4189);
and U4647 (N_4647,N_4178,N_4473);
or U4648 (N_4648,N_4066,N_4307);
nand U4649 (N_4649,N_4105,N_4228);
nand U4650 (N_4650,N_4138,N_4367);
or U4651 (N_4651,N_4482,N_4239);
nor U4652 (N_4652,N_4090,N_4254);
nor U4653 (N_4653,N_4033,N_4252);
and U4654 (N_4654,N_4376,N_4061);
nor U4655 (N_4655,N_4227,N_4206);
xnor U4656 (N_4656,N_4194,N_4489);
xor U4657 (N_4657,N_4292,N_4142);
and U4658 (N_4658,N_4389,N_4010);
nand U4659 (N_4659,N_4318,N_4170);
or U4660 (N_4660,N_4404,N_4465);
and U4661 (N_4661,N_4256,N_4072);
or U4662 (N_4662,N_4363,N_4301);
xnor U4663 (N_4663,N_4312,N_4026);
and U4664 (N_4664,N_4197,N_4306);
xnor U4665 (N_4665,N_4320,N_4464);
nor U4666 (N_4666,N_4261,N_4364);
or U4667 (N_4667,N_4266,N_4287);
and U4668 (N_4668,N_4229,N_4176);
or U4669 (N_4669,N_4331,N_4161);
or U4670 (N_4670,N_4457,N_4050);
nor U4671 (N_4671,N_4130,N_4408);
xor U4672 (N_4672,N_4351,N_4201);
nand U4673 (N_4673,N_4169,N_4018);
nor U4674 (N_4674,N_4149,N_4007);
xor U4675 (N_4675,N_4127,N_4042);
nor U4676 (N_4676,N_4038,N_4236);
or U4677 (N_4677,N_4140,N_4469);
and U4678 (N_4678,N_4116,N_4110);
xor U4679 (N_4679,N_4071,N_4277);
or U4680 (N_4680,N_4387,N_4115);
nand U4681 (N_4681,N_4011,N_4063);
nor U4682 (N_4682,N_4174,N_4173);
and U4683 (N_4683,N_4222,N_4291);
xor U4684 (N_4684,N_4368,N_4013);
or U4685 (N_4685,N_4402,N_4374);
xor U4686 (N_4686,N_4392,N_4335);
and U4687 (N_4687,N_4219,N_4403);
nand U4688 (N_4688,N_4109,N_4272);
or U4689 (N_4689,N_4276,N_4386);
nor U4690 (N_4690,N_4107,N_4492);
nand U4691 (N_4691,N_4347,N_4234);
or U4692 (N_4692,N_4305,N_4100);
and U4693 (N_4693,N_4477,N_4086);
and U4694 (N_4694,N_4471,N_4213);
nor U4695 (N_4695,N_4444,N_4132);
xnor U4696 (N_4696,N_4095,N_4150);
nand U4697 (N_4697,N_4270,N_4137);
nor U4698 (N_4698,N_4131,N_4362);
nand U4699 (N_4699,N_4370,N_4420);
nor U4700 (N_4700,N_4156,N_4284);
or U4701 (N_4701,N_4052,N_4204);
nor U4702 (N_4702,N_4221,N_4134);
nor U4703 (N_4703,N_4349,N_4214);
nor U4704 (N_4704,N_4062,N_4006);
xnor U4705 (N_4705,N_4410,N_4283);
nand U4706 (N_4706,N_4135,N_4251);
nor U4707 (N_4707,N_4434,N_4340);
nand U4708 (N_4708,N_4060,N_4330);
xnor U4709 (N_4709,N_4263,N_4415);
nand U4710 (N_4710,N_4466,N_4074);
nand U4711 (N_4711,N_4242,N_4337);
or U4712 (N_4712,N_4346,N_4441);
and U4713 (N_4713,N_4136,N_4031);
nand U4714 (N_4714,N_4118,N_4421);
or U4715 (N_4715,N_4002,N_4054);
nor U4716 (N_4716,N_4447,N_4334);
nor U4717 (N_4717,N_4316,N_4416);
or U4718 (N_4718,N_4019,N_4096);
nor U4719 (N_4719,N_4023,N_4395);
nand U4720 (N_4720,N_4365,N_4459);
and U4721 (N_4721,N_4336,N_4274);
nand U4722 (N_4722,N_4491,N_4155);
xor U4723 (N_4723,N_4443,N_4286);
xor U4724 (N_4724,N_4391,N_4053);
and U4725 (N_4725,N_4329,N_4129);
nand U4726 (N_4726,N_4080,N_4045);
or U4727 (N_4727,N_4166,N_4017);
nor U4728 (N_4728,N_4458,N_4203);
and U4729 (N_4729,N_4188,N_4456);
nor U4730 (N_4730,N_4171,N_4202);
and U4731 (N_4731,N_4353,N_4384);
and U4732 (N_4732,N_4430,N_4141);
and U4733 (N_4733,N_4383,N_4328);
xnor U4734 (N_4734,N_4350,N_4435);
nand U4735 (N_4735,N_4352,N_4425);
nand U4736 (N_4736,N_4344,N_4106);
nand U4737 (N_4737,N_4216,N_4460);
nor U4738 (N_4738,N_4065,N_4104);
and U4739 (N_4739,N_4003,N_4154);
or U4740 (N_4740,N_4212,N_4398);
xnor U4741 (N_4741,N_4016,N_4412);
nor U4742 (N_4742,N_4345,N_4355);
nor U4743 (N_4743,N_4375,N_4279);
and U4744 (N_4744,N_4059,N_4043);
xnor U4745 (N_4745,N_4409,N_4399);
or U4746 (N_4746,N_4282,N_4073);
or U4747 (N_4747,N_4114,N_4025);
nand U4748 (N_4748,N_4195,N_4407);
xnor U4749 (N_4749,N_4485,N_4281);
or U4750 (N_4750,N_4216,N_4406);
xnor U4751 (N_4751,N_4278,N_4400);
nand U4752 (N_4752,N_4347,N_4192);
or U4753 (N_4753,N_4021,N_4162);
and U4754 (N_4754,N_4213,N_4142);
and U4755 (N_4755,N_4442,N_4110);
xnor U4756 (N_4756,N_4055,N_4203);
and U4757 (N_4757,N_4412,N_4457);
nor U4758 (N_4758,N_4417,N_4119);
nor U4759 (N_4759,N_4303,N_4129);
nand U4760 (N_4760,N_4016,N_4366);
nand U4761 (N_4761,N_4317,N_4257);
nor U4762 (N_4762,N_4138,N_4004);
nand U4763 (N_4763,N_4259,N_4002);
nand U4764 (N_4764,N_4030,N_4022);
nor U4765 (N_4765,N_4068,N_4189);
nor U4766 (N_4766,N_4274,N_4364);
and U4767 (N_4767,N_4165,N_4101);
nand U4768 (N_4768,N_4091,N_4174);
nand U4769 (N_4769,N_4364,N_4406);
nor U4770 (N_4770,N_4361,N_4102);
nand U4771 (N_4771,N_4298,N_4409);
nand U4772 (N_4772,N_4129,N_4433);
or U4773 (N_4773,N_4298,N_4465);
nor U4774 (N_4774,N_4094,N_4489);
nand U4775 (N_4775,N_4034,N_4312);
and U4776 (N_4776,N_4035,N_4493);
nor U4777 (N_4777,N_4263,N_4362);
nor U4778 (N_4778,N_4006,N_4431);
and U4779 (N_4779,N_4006,N_4196);
and U4780 (N_4780,N_4334,N_4044);
nand U4781 (N_4781,N_4119,N_4314);
nor U4782 (N_4782,N_4440,N_4482);
nor U4783 (N_4783,N_4422,N_4364);
nor U4784 (N_4784,N_4327,N_4178);
or U4785 (N_4785,N_4058,N_4370);
xnor U4786 (N_4786,N_4253,N_4220);
or U4787 (N_4787,N_4266,N_4020);
and U4788 (N_4788,N_4112,N_4318);
nand U4789 (N_4789,N_4263,N_4150);
xnor U4790 (N_4790,N_4355,N_4343);
nor U4791 (N_4791,N_4369,N_4439);
xor U4792 (N_4792,N_4230,N_4049);
or U4793 (N_4793,N_4318,N_4033);
or U4794 (N_4794,N_4035,N_4226);
nor U4795 (N_4795,N_4209,N_4034);
and U4796 (N_4796,N_4312,N_4422);
and U4797 (N_4797,N_4125,N_4170);
nand U4798 (N_4798,N_4400,N_4496);
nand U4799 (N_4799,N_4327,N_4130);
xnor U4800 (N_4800,N_4261,N_4295);
nor U4801 (N_4801,N_4322,N_4156);
or U4802 (N_4802,N_4205,N_4242);
nor U4803 (N_4803,N_4156,N_4184);
nor U4804 (N_4804,N_4078,N_4401);
and U4805 (N_4805,N_4424,N_4372);
nor U4806 (N_4806,N_4294,N_4278);
nor U4807 (N_4807,N_4107,N_4236);
xor U4808 (N_4808,N_4111,N_4285);
nand U4809 (N_4809,N_4001,N_4244);
nor U4810 (N_4810,N_4430,N_4202);
and U4811 (N_4811,N_4285,N_4126);
nand U4812 (N_4812,N_4330,N_4204);
or U4813 (N_4813,N_4210,N_4003);
and U4814 (N_4814,N_4134,N_4431);
or U4815 (N_4815,N_4137,N_4213);
nand U4816 (N_4816,N_4148,N_4332);
nand U4817 (N_4817,N_4272,N_4458);
nand U4818 (N_4818,N_4468,N_4034);
xnor U4819 (N_4819,N_4434,N_4143);
nand U4820 (N_4820,N_4100,N_4427);
nor U4821 (N_4821,N_4280,N_4037);
nor U4822 (N_4822,N_4341,N_4066);
nor U4823 (N_4823,N_4232,N_4074);
or U4824 (N_4824,N_4057,N_4337);
and U4825 (N_4825,N_4140,N_4461);
xor U4826 (N_4826,N_4169,N_4014);
or U4827 (N_4827,N_4442,N_4014);
xor U4828 (N_4828,N_4088,N_4129);
xnor U4829 (N_4829,N_4325,N_4130);
nor U4830 (N_4830,N_4105,N_4023);
nor U4831 (N_4831,N_4192,N_4111);
and U4832 (N_4832,N_4353,N_4401);
nand U4833 (N_4833,N_4423,N_4244);
xor U4834 (N_4834,N_4086,N_4368);
and U4835 (N_4835,N_4229,N_4401);
nor U4836 (N_4836,N_4237,N_4243);
or U4837 (N_4837,N_4267,N_4438);
and U4838 (N_4838,N_4162,N_4477);
and U4839 (N_4839,N_4047,N_4315);
nand U4840 (N_4840,N_4312,N_4146);
or U4841 (N_4841,N_4336,N_4279);
xnor U4842 (N_4842,N_4297,N_4183);
nor U4843 (N_4843,N_4223,N_4345);
nor U4844 (N_4844,N_4257,N_4288);
and U4845 (N_4845,N_4337,N_4439);
and U4846 (N_4846,N_4139,N_4128);
nor U4847 (N_4847,N_4233,N_4175);
nand U4848 (N_4848,N_4093,N_4016);
xnor U4849 (N_4849,N_4243,N_4035);
nor U4850 (N_4850,N_4404,N_4331);
and U4851 (N_4851,N_4055,N_4221);
xor U4852 (N_4852,N_4428,N_4236);
or U4853 (N_4853,N_4157,N_4002);
xor U4854 (N_4854,N_4221,N_4116);
or U4855 (N_4855,N_4364,N_4471);
and U4856 (N_4856,N_4375,N_4458);
nor U4857 (N_4857,N_4354,N_4405);
nand U4858 (N_4858,N_4401,N_4304);
or U4859 (N_4859,N_4233,N_4006);
or U4860 (N_4860,N_4131,N_4023);
nor U4861 (N_4861,N_4083,N_4076);
or U4862 (N_4862,N_4346,N_4141);
nand U4863 (N_4863,N_4001,N_4452);
or U4864 (N_4864,N_4413,N_4362);
xnor U4865 (N_4865,N_4499,N_4207);
nand U4866 (N_4866,N_4121,N_4138);
or U4867 (N_4867,N_4416,N_4080);
and U4868 (N_4868,N_4489,N_4430);
nor U4869 (N_4869,N_4127,N_4411);
nor U4870 (N_4870,N_4326,N_4274);
nand U4871 (N_4871,N_4047,N_4140);
xor U4872 (N_4872,N_4199,N_4363);
or U4873 (N_4873,N_4287,N_4392);
and U4874 (N_4874,N_4316,N_4020);
nand U4875 (N_4875,N_4376,N_4401);
xnor U4876 (N_4876,N_4021,N_4480);
nor U4877 (N_4877,N_4079,N_4378);
or U4878 (N_4878,N_4457,N_4027);
nor U4879 (N_4879,N_4141,N_4198);
or U4880 (N_4880,N_4431,N_4173);
or U4881 (N_4881,N_4481,N_4067);
and U4882 (N_4882,N_4026,N_4240);
nand U4883 (N_4883,N_4441,N_4436);
nor U4884 (N_4884,N_4036,N_4452);
and U4885 (N_4885,N_4395,N_4054);
xor U4886 (N_4886,N_4136,N_4408);
xor U4887 (N_4887,N_4374,N_4176);
or U4888 (N_4888,N_4177,N_4396);
nand U4889 (N_4889,N_4175,N_4256);
nand U4890 (N_4890,N_4435,N_4001);
nand U4891 (N_4891,N_4289,N_4199);
and U4892 (N_4892,N_4296,N_4111);
nor U4893 (N_4893,N_4325,N_4198);
xor U4894 (N_4894,N_4108,N_4321);
xor U4895 (N_4895,N_4015,N_4190);
nand U4896 (N_4896,N_4391,N_4190);
and U4897 (N_4897,N_4374,N_4062);
and U4898 (N_4898,N_4426,N_4281);
and U4899 (N_4899,N_4086,N_4177);
nor U4900 (N_4900,N_4104,N_4188);
and U4901 (N_4901,N_4087,N_4258);
and U4902 (N_4902,N_4386,N_4145);
or U4903 (N_4903,N_4143,N_4432);
or U4904 (N_4904,N_4278,N_4259);
nor U4905 (N_4905,N_4016,N_4183);
xor U4906 (N_4906,N_4239,N_4281);
xnor U4907 (N_4907,N_4356,N_4114);
or U4908 (N_4908,N_4314,N_4414);
or U4909 (N_4909,N_4144,N_4071);
or U4910 (N_4910,N_4334,N_4114);
xnor U4911 (N_4911,N_4219,N_4281);
nand U4912 (N_4912,N_4134,N_4187);
and U4913 (N_4913,N_4370,N_4294);
and U4914 (N_4914,N_4333,N_4151);
nor U4915 (N_4915,N_4481,N_4369);
xor U4916 (N_4916,N_4385,N_4085);
and U4917 (N_4917,N_4277,N_4480);
nor U4918 (N_4918,N_4252,N_4379);
nand U4919 (N_4919,N_4065,N_4323);
and U4920 (N_4920,N_4313,N_4076);
nor U4921 (N_4921,N_4303,N_4254);
nor U4922 (N_4922,N_4144,N_4339);
or U4923 (N_4923,N_4147,N_4412);
or U4924 (N_4924,N_4247,N_4182);
nor U4925 (N_4925,N_4319,N_4347);
nor U4926 (N_4926,N_4176,N_4020);
xnor U4927 (N_4927,N_4197,N_4405);
nor U4928 (N_4928,N_4485,N_4335);
nor U4929 (N_4929,N_4106,N_4108);
xor U4930 (N_4930,N_4434,N_4080);
nor U4931 (N_4931,N_4257,N_4440);
nand U4932 (N_4932,N_4466,N_4374);
nor U4933 (N_4933,N_4434,N_4317);
xnor U4934 (N_4934,N_4203,N_4341);
nor U4935 (N_4935,N_4265,N_4312);
and U4936 (N_4936,N_4201,N_4137);
nor U4937 (N_4937,N_4436,N_4119);
nor U4938 (N_4938,N_4374,N_4226);
or U4939 (N_4939,N_4312,N_4332);
xnor U4940 (N_4940,N_4070,N_4246);
or U4941 (N_4941,N_4242,N_4150);
or U4942 (N_4942,N_4019,N_4432);
and U4943 (N_4943,N_4041,N_4471);
xor U4944 (N_4944,N_4004,N_4298);
xnor U4945 (N_4945,N_4309,N_4480);
and U4946 (N_4946,N_4111,N_4392);
xor U4947 (N_4947,N_4070,N_4105);
nand U4948 (N_4948,N_4420,N_4127);
xnor U4949 (N_4949,N_4063,N_4496);
and U4950 (N_4950,N_4095,N_4231);
xnor U4951 (N_4951,N_4106,N_4211);
or U4952 (N_4952,N_4150,N_4048);
nor U4953 (N_4953,N_4169,N_4062);
xnor U4954 (N_4954,N_4407,N_4057);
and U4955 (N_4955,N_4143,N_4164);
xor U4956 (N_4956,N_4169,N_4008);
nand U4957 (N_4957,N_4210,N_4363);
nand U4958 (N_4958,N_4392,N_4360);
nor U4959 (N_4959,N_4277,N_4221);
xor U4960 (N_4960,N_4313,N_4184);
nor U4961 (N_4961,N_4284,N_4075);
nor U4962 (N_4962,N_4056,N_4088);
nor U4963 (N_4963,N_4088,N_4266);
and U4964 (N_4964,N_4434,N_4063);
xnor U4965 (N_4965,N_4228,N_4101);
and U4966 (N_4966,N_4438,N_4120);
nand U4967 (N_4967,N_4288,N_4428);
nand U4968 (N_4968,N_4397,N_4362);
nand U4969 (N_4969,N_4414,N_4222);
or U4970 (N_4970,N_4325,N_4340);
nand U4971 (N_4971,N_4425,N_4041);
or U4972 (N_4972,N_4463,N_4292);
or U4973 (N_4973,N_4050,N_4266);
and U4974 (N_4974,N_4465,N_4474);
and U4975 (N_4975,N_4033,N_4250);
or U4976 (N_4976,N_4499,N_4472);
nor U4977 (N_4977,N_4185,N_4114);
or U4978 (N_4978,N_4417,N_4376);
and U4979 (N_4979,N_4111,N_4356);
nand U4980 (N_4980,N_4367,N_4167);
and U4981 (N_4981,N_4336,N_4192);
and U4982 (N_4982,N_4459,N_4308);
xor U4983 (N_4983,N_4274,N_4311);
or U4984 (N_4984,N_4471,N_4329);
xnor U4985 (N_4985,N_4344,N_4064);
or U4986 (N_4986,N_4196,N_4332);
xnor U4987 (N_4987,N_4184,N_4315);
xnor U4988 (N_4988,N_4016,N_4083);
nand U4989 (N_4989,N_4138,N_4422);
or U4990 (N_4990,N_4217,N_4028);
and U4991 (N_4991,N_4456,N_4292);
nor U4992 (N_4992,N_4293,N_4170);
nand U4993 (N_4993,N_4229,N_4266);
or U4994 (N_4994,N_4055,N_4463);
or U4995 (N_4995,N_4189,N_4490);
and U4996 (N_4996,N_4425,N_4183);
nand U4997 (N_4997,N_4097,N_4060);
nand U4998 (N_4998,N_4270,N_4289);
nor U4999 (N_4999,N_4014,N_4381);
or U5000 (N_5000,N_4618,N_4711);
nand U5001 (N_5001,N_4690,N_4718);
or U5002 (N_5002,N_4517,N_4689);
nand U5003 (N_5003,N_4667,N_4547);
xor U5004 (N_5004,N_4930,N_4842);
or U5005 (N_5005,N_4642,N_4692);
nand U5006 (N_5006,N_4544,N_4817);
nand U5007 (N_5007,N_4830,N_4658);
nor U5008 (N_5008,N_4999,N_4661);
nand U5009 (N_5009,N_4870,N_4738);
nand U5010 (N_5010,N_4515,N_4601);
nor U5011 (N_5011,N_4778,N_4583);
and U5012 (N_5012,N_4635,N_4825);
nor U5013 (N_5013,N_4901,N_4972);
or U5014 (N_5014,N_4745,N_4827);
nor U5015 (N_5015,N_4864,N_4907);
and U5016 (N_5016,N_4501,N_4510);
or U5017 (N_5017,N_4984,N_4931);
or U5018 (N_5018,N_4740,N_4823);
nor U5019 (N_5019,N_4557,N_4571);
xnor U5020 (N_5020,N_4888,N_4813);
or U5021 (N_5021,N_4576,N_4669);
and U5022 (N_5022,N_4623,N_4525);
nor U5023 (N_5023,N_4921,N_4586);
or U5024 (N_5024,N_4857,N_4719);
nor U5025 (N_5025,N_4770,N_4596);
nor U5026 (N_5026,N_4620,N_4737);
and U5027 (N_5027,N_4906,N_4704);
xnor U5028 (N_5028,N_4874,N_4734);
nand U5029 (N_5029,N_4611,N_4569);
nand U5030 (N_5030,N_4573,N_4800);
xnor U5031 (N_5031,N_4795,N_4528);
nand U5032 (N_5032,N_4927,N_4687);
xor U5033 (N_5033,N_4575,N_4915);
or U5034 (N_5034,N_4565,N_4736);
or U5035 (N_5035,N_4772,N_4807);
nand U5036 (N_5036,N_4735,N_4881);
xnor U5037 (N_5037,N_4723,N_4810);
xnor U5038 (N_5038,N_4920,N_4793);
nand U5039 (N_5039,N_4574,N_4905);
or U5040 (N_5040,N_4929,N_4783);
or U5041 (N_5041,N_4732,N_4892);
nor U5042 (N_5042,N_4521,N_4945);
and U5043 (N_5043,N_4987,N_4861);
nand U5044 (N_5044,N_4524,N_4750);
xor U5045 (N_5045,N_4978,N_4943);
and U5046 (N_5046,N_4814,N_4647);
and U5047 (N_5047,N_4947,N_4784);
xnor U5048 (N_5048,N_4540,N_4578);
or U5049 (N_5049,N_4961,N_4638);
and U5050 (N_5050,N_4804,N_4725);
xor U5051 (N_5051,N_4808,N_4624);
nand U5052 (N_5052,N_4934,N_4616);
or U5053 (N_5053,N_4787,N_4971);
and U5054 (N_5054,N_4603,N_4568);
nor U5055 (N_5055,N_4964,N_4581);
nor U5056 (N_5056,N_4869,N_4598);
nor U5057 (N_5057,N_4832,N_4660);
nor U5058 (N_5058,N_4767,N_4913);
and U5059 (N_5059,N_4679,N_4634);
xnor U5060 (N_5060,N_4829,N_4791);
nand U5061 (N_5061,N_4577,N_4656);
xnor U5062 (N_5062,N_4854,N_4815);
nor U5063 (N_5063,N_4703,N_4998);
xor U5064 (N_5064,N_4739,N_4867);
and U5065 (N_5065,N_4756,N_4629);
nand U5066 (N_5066,N_4883,N_4952);
and U5067 (N_5067,N_4786,N_4776);
and U5068 (N_5068,N_4805,N_4744);
or U5069 (N_5069,N_4836,N_4760);
or U5070 (N_5070,N_4664,N_4500);
nor U5071 (N_5071,N_4503,N_4533);
or U5072 (N_5072,N_4965,N_4560);
or U5073 (N_5073,N_4944,N_4975);
nand U5074 (N_5074,N_4518,N_4922);
xor U5075 (N_5075,N_4946,N_4876);
and U5076 (N_5076,N_4564,N_4530);
nand U5077 (N_5077,N_4802,N_4588);
nand U5078 (N_5078,N_4685,N_4562);
nor U5079 (N_5079,N_4715,N_4539);
and U5080 (N_5080,N_4879,N_4712);
and U5081 (N_5081,N_4937,N_4672);
and U5082 (N_5082,N_4966,N_4741);
or U5083 (N_5083,N_4619,N_4923);
xnor U5084 (N_5084,N_4798,N_4654);
nor U5085 (N_5085,N_4849,N_4893);
or U5086 (N_5086,N_4622,N_4792);
xnor U5087 (N_5087,N_4597,N_4797);
xor U5088 (N_5088,N_4592,N_4537);
nand U5089 (N_5089,N_4866,N_4919);
xnor U5090 (N_5090,N_4651,N_4646);
and U5091 (N_5091,N_4731,N_4853);
nand U5092 (N_5092,N_4653,N_4749);
and U5093 (N_5093,N_4962,N_4582);
or U5094 (N_5094,N_4834,N_4591);
and U5095 (N_5095,N_4520,N_4790);
or U5096 (N_5096,N_4705,N_4785);
and U5097 (N_5097,N_4926,N_4639);
nand U5098 (N_5098,N_4506,N_4645);
nor U5099 (N_5099,N_4709,N_4650);
nor U5100 (N_5100,N_4774,N_4779);
nor U5101 (N_5101,N_4902,N_4567);
xnor U5102 (N_5102,N_4835,N_4608);
nand U5103 (N_5103,N_4755,N_4811);
nand U5104 (N_5104,N_4941,N_4753);
nand U5105 (N_5105,N_4796,N_4928);
nor U5106 (N_5106,N_4561,N_4722);
xor U5107 (N_5107,N_4585,N_4904);
xnor U5108 (N_5108,N_4911,N_4968);
nor U5109 (N_5109,N_4652,N_4511);
and U5110 (N_5110,N_4949,N_4694);
or U5111 (N_5111,N_4769,N_4681);
or U5112 (N_5112,N_4532,N_4789);
nor U5113 (N_5113,N_4974,N_4936);
nor U5114 (N_5114,N_4884,N_4855);
xnor U5115 (N_5115,N_4875,N_4512);
or U5116 (N_5116,N_4534,N_4665);
nand U5117 (N_5117,N_4543,N_4717);
xor U5118 (N_5118,N_4950,N_4863);
nand U5119 (N_5119,N_4566,N_4840);
nor U5120 (N_5120,N_4643,N_4914);
nand U5121 (N_5121,N_4579,N_4831);
or U5122 (N_5122,N_4555,N_4548);
and U5123 (N_5123,N_4746,N_4541);
nand U5124 (N_5124,N_4648,N_4673);
nor U5125 (N_5125,N_4886,N_4513);
or U5126 (N_5126,N_4880,N_4948);
nor U5127 (N_5127,N_4505,N_4916);
nand U5128 (N_5128,N_4986,N_4625);
nor U5129 (N_5129,N_4801,N_4860);
nand U5130 (N_5130,N_4841,N_4594);
xor U5131 (N_5131,N_4821,N_4878);
nand U5132 (N_5132,N_4605,N_4988);
or U5133 (N_5133,N_4730,N_4644);
nand U5134 (N_5134,N_4726,N_4678);
and U5135 (N_5135,N_4826,N_4542);
or U5136 (N_5136,N_4933,N_4885);
or U5137 (N_5137,N_4570,N_4742);
and U5138 (N_5138,N_4816,N_4994);
nand U5139 (N_5139,N_4762,N_4612);
and U5140 (N_5140,N_4871,N_4688);
or U5141 (N_5141,N_4535,N_4680);
nand U5142 (N_5142,N_4641,N_4761);
xor U5143 (N_5143,N_4889,N_4777);
and U5144 (N_5144,N_4806,N_4953);
nor U5145 (N_5145,N_4981,N_4636);
or U5146 (N_5146,N_4851,N_4630);
or U5147 (N_5147,N_4587,N_4768);
nor U5148 (N_5148,N_4925,N_4788);
nor U5149 (N_5149,N_4780,N_4676);
and U5150 (N_5150,N_4508,N_4955);
and U5151 (N_5151,N_4584,N_4982);
nand U5152 (N_5152,N_4663,N_4529);
nor U5153 (N_5153,N_4877,N_4626);
or U5154 (N_5154,N_4504,N_4852);
and U5155 (N_5155,N_4657,N_4764);
nor U5156 (N_5156,N_4729,N_4812);
xor U5157 (N_5157,N_4822,N_4590);
nor U5158 (N_5158,N_4935,N_4846);
nor U5159 (N_5159,N_4958,N_4765);
xnor U5160 (N_5160,N_4979,N_4918);
or U5161 (N_5161,N_4649,N_4683);
nand U5162 (N_5162,N_4527,N_4782);
and U5163 (N_5163,N_4803,N_4701);
and U5164 (N_5164,N_4833,N_4748);
or U5165 (N_5165,N_4819,N_4940);
and U5166 (N_5166,N_4628,N_4702);
nor U5167 (N_5167,N_4640,N_4552);
xnor U5168 (N_5168,N_4794,N_4706);
nor U5169 (N_5169,N_4708,N_4522);
nor U5170 (N_5170,N_4684,N_4662);
xnor U5171 (N_5171,N_4589,N_4848);
nand U5172 (N_5172,N_4607,N_4960);
nand U5173 (N_5173,N_4536,N_4695);
nor U5174 (N_5174,N_4896,N_4580);
and U5175 (N_5175,N_4824,N_4617);
nor U5176 (N_5176,N_4939,N_4997);
or U5177 (N_5177,N_4507,N_4752);
xnor U5178 (N_5178,N_4995,N_4593);
nor U5179 (N_5179,N_4951,N_4843);
or U5180 (N_5180,N_4682,N_4894);
xor U5181 (N_5181,N_4686,N_4938);
and U5182 (N_5182,N_4724,N_4655);
and U5183 (N_5183,N_4519,N_4710);
nand U5184 (N_5184,N_4599,N_4954);
xor U5185 (N_5185,N_4743,N_4775);
nor U5186 (N_5186,N_4991,N_4900);
xnor U5187 (N_5187,N_4728,N_4516);
nor U5188 (N_5188,N_4809,N_4912);
nor U5189 (N_5189,N_4526,N_4713);
or U5190 (N_5190,N_4858,N_4957);
nor U5191 (N_5191,N_4727,N_4675);
and U5192 (N_5192,N_4632,N_4609);
xnor U5193 (N_5193,N_4666,N_4983);
nor U5194 (N_5194,N_4845,N_4977);
nand U5195 (N_5195,N_4700,N_4872);
nand U5196 (N_5196,N_4970,N_4898);
or U5197 (N_5197,N_4847,N_4859);
and U5198 (N_5198,N_4766,N_4973);
nor U5199 (N_5199,N_4771,N_4670);
xor U5200 (N_5200,N_4844,N_4615);
nor U5201 (N_5201,N_4799,N_4759);
or U5202 (N_5202,N_4671,N_4606);
or U5203 (N_5203,N_4721,N_4637);
xnor U5204 (N_5204,N_4613,N_4838);
and U5205 (N_5205,N_4985,N_4621);
and U5206 (N_5206,N_4865,N_4716);
or U5207 (N_5207,N_4909,N_4903);
and U5208 (N_5208,N_4917,N_4509);
nand U5209 (N_5209,N_4747,N_4895);
nor U5210 (N_5210,N_4602,N_4758);
nand U5211 (N_5211,N_4932,N_4963);
or U5212 (N_5212,N_4549,N_4523);
nor U5213 (N_5213,N_4545,N_4856);
nand U5214 (N_5214,N_4828,N_4899);
and U5215 (N_5215,N_4754,N_4956);
or U5216 (N_5216,N_4707,N_4820);
or U5217 (N_5217,N_4757,N_4610);
nand U5218 (N_5218,N_4631,N_4980);
xor U5219 (N_5219,N_4763,N_4559);
nand U5220 (N_5220,N_4674,N_4996);
and U5221 (N_5221,N_4992,N_4633);
and U5222 (N_5222,N_4969,N_4538);
and U5223 (N_5223,N_4862,N_4699);
and U5224 (N_5224,N_4751,N_4693);
and U5225 (N_5225,N_4733,N_4553);
nor U5226 (N_5226,N_4668,N_4868);
or U5227 (N_5227,N_4890,N_4891);
and U5228 (N_5228,N_4554,N_4691);
or U5229 (N_5229,N_4908,N_4959);
nand U5230 (N_5230,N_4910,N_4595);
or U5231 (N_5231,N_4850,N_4546);
and U5232 (N_5232,N_4514,N_4714);
and U5233 (N_5233,N_4627,N_4698);
nor U5234 (N_5234,N_4556,N_4989);
nand U5235 (N_5235,N_4781,N_4697);
nand U5236 (N_5236,N_4604,N_4600);
nand U5237 (N_5237,N_4563,N_4897);
nand U5238 (N_5238,N_4531,N_4773);
xor U5239 (N_5239,N_4720,N_4942);
xnor U5240 (N_5240,N_4502,N_4887);
and U5241 (N_5241,N_4976,N_4818);
xnor U5242 (N_5242,N_4572,N_4696);
and U5243 (N_5243,N_4614,N_4990);
and U5244 (N_5244,N_4967,N_4873);
or U5245 (N_5245,N_4558,N_4924);
nor U5246 (N_5246,N_4839,N_4837);
or U5247 (N_5247,N_4677,N_4993);
or U5248 (N_5248,N_4882,N_4551);
or U5249 (N_5249,N_4659,N_4550);
or U5250 (N_5250,N_4802,N_4827);
or U5251 (N_5251,N_4623,N_4553);
nor U5252 (N_5252,N_4974,N_4575);
nor U5253 (N_5253,N_4759,N_4528);
and U5254 (N_5254,N_4826,N_4822);
or U5255 (N_5255,N_4779,N_4501);
and U5256 (N_5256,N_4803,N_4793);
xnor U5257 (N_5257,N_4935,N_4654);
nor U5258 (N_5258,N_4568,N_4614);
nand U5259 (N_5259,N_4786,N_4556);
nand U5260 (N_5260,N_4954,N_4918);
nor U5261 (N_5261,N_4769,N_4867);
or U5262 (N_5262,N_4774,N_4689);
nor U5263 (N_5263,N_4619,N_4975);
nor U5264 (N_5264,N_4714,N_4608);
nand U5265 (N_5265,N_4531,N_4939);
nor U5266 (N_5266,N_4530,N_4656);
nor U5267 (N_5267,N_4574,N_4520);
or U5268 (N_5268,N_4670,N_4883);
nand U5269 (N_5269,N_4730,N_4875);
or U5270 (N_5270,N_4868,N_4946);
or U5271 (N_5271,N_4703,N_4934);
nand U5272 (N_5272,N_4904,N_4859);
nand U5273 (N_5273,N_4923,N_4562);
or U5274 (N_5274,N_4754,N_4652);
and U5275 (N_5275,N_4654,N_4993);
and U5276 (N_5276,N_4619,N_4776);
nor U5277 (N_5277,N_4889,N_4848);
xor U5278 (N_5278,N_4920,N_4699);
nor U5279 (N_5279,N_4791,N_4645);
xnor U5280 (N_5280,N_4668,N_4683);
or U5281 (N_5281,N_4505,N_4711);
nand U5282 (N_5282,N_4574,N_4799);
and U5283 (N_5283,N_4970,N_4617);
nand U5284 (N_5284,N_4914,N_4679);
or U5285 (N_5285,N_4600,N_4605);
nor U5286 (N_5286,N_4951,N_4519);
and U5287 (N_5287,N_4783,N_4830);
or U5288 (N_5288,N_4560,N_4530);
nand U5289 (N_5289,N_4827,N_4790);
nor U5290 (N_5290,N_4997,N_4888);
and U5291 (N_5291,N_4987,N_4918);
xor U5292 (N_5292,N_4726,N_4906);
nand U5293 (N_5293,N_4827,N_4850);
xnor U5294 (N_5294,N_4611,N_4912);
or U5295 (N_5295,N_4772,N_4801);
or U5296 (N_5296,N_4814,N_4717);
nand U5297 (N_5297,N_4762,N_4614);
nor U5298 (N_5298,N_4994,N_4626);
nor U5299 (N_5299,N_4687,N_4549);
or U5300 (N_5300,N_4524,N_4650);
xnor U5301 (N_5301,N_4906,N_4873);
or U5302 (N_5302,N_4946,N_4900);
or U5303 (N_5303,N_4701,N_4683);
nor U5304 (N_5304,N_4621,N_4801);
xnor U5305 (N_5305,N_4656,N_4957);
nand U5306 (N_5306,N_4860,N_4579);
nand U5307 (N_5307,N_4996,N_4872);
xor U5308 (N_5308,N_4989,N_4673);
and U5309 (N_5309,N_4895,N_4631);
xnor U5310 (N_5310,N_4933,N_4818);
or U5311 (N_5311,N_4858,N_4854);
or U5312 (N_5312,N_4549,N_4824);
xor U5313 (N_5313,N_4865,N_4613);
and U5314 (N_5314,N_4660,N_4715);
nor U5315 (N_5315,N_4991,N_4872);
xor U5316 (N_5316,N_4768,N_4629);
nor U5317 (N_5317,N_4579,N_4910);
nor U5318 (N_5318,N_4563,N_4524);
or U5319 (N_5319,N_4682,N_4584);
xor U5320 (N_5320,N_4547,N_4848);
xnor U5321 (N_5321,N_4528,N_4806);
or U5322 (N_5322,N_4689,N_4946);
nand U5323 (N_5323,N_4596,N_4606);
xnor U5324 (N_5324,N_4631,N_4744);
and U5325 (N_5325,N_4618,N_4590);
and U5326 (N_5326,N_4654,N_4779);
xnor U5327 (N_5327,N_4986,N_4787);
xor U5328 (N_5328,N_4861,N_4531);
nor U5329 (N_5329,N_4760,N_4547);
nor U5330 (N_5330,N_4760,N_4761);
and U5331 (N_5331,N_4595,N_4630);
and U5332 (N_5332,N_4931,N_4769);
nand U5333 (N_5333,N_4745,N_4818);
and U5334 (N_5334,N_4831,N_4649);
nor U5335 (N_5335,N_4564,N_4718);
or U5336 (N_5336,N_4905,N_4730);
or U5337 (N_5337,N_4544,N_4871);
and U5338 (N_5338,N_4950,N_4762);
or U5339 (N_5339,N_4971,N_4930);
and U5340 (N_5340,N_4681,N_4933);
and U5341 (N_5341,N_4629,N_4717);
or U5342 (N_5342,N_4772,N_4768);
and U5343 (N_5343,N_4976,N_4727);
nor U5344 (N_5344,N_4684,N_4870);
nor U5345 (N_5345,N_4798,N_4874);
and U5346 (N_5346,N_4523,N_4796);
and U5347 (N_5347,N_4939,N_4751);
or U5348 (N_5348,N_4693,N_4569);
nor U5349 (N_5349,N_4798,N_4591);
xnor U5350 (N_5350,N_4629,N_4884);
and U5351 (N_5351,N_4839,N_4835);
nor U5352 (N_5352,N_4930,N_4580);
and U5353 (N_5353,N_4547,N_4588);
and U5354 (N_5354,N_4539,N_4940);
nand U5355 (N_5355,N_4623,N_4668);
and U5356 (N_5356,N_4845,N_4649);
nor U5357 (N_5357,N_4673,N_4637);
or U5358 (N_5358,N_4767,N_4664);
or U5359 (N_5359,N_4989,N_4802);
xnor U5360 (N_5360,N_4538,N_4658);
xor U5361 (N_5361,N_4575,N_4694);
nand U5362 (N_5362,N_4512,N_4931);
or U5363 (N_5363,N_4540,N_4642);
or U5364 (N_5364,N_4651,N_4715);
xnor U5365 (N_5365,N_4580,N_4538);
and U5366 (N_5366,N_4754,N_4551);
and U5367 (N_5367,N_4530,N_4979);
or U5368 (N_5368,N_4619,N_4799);
xnor U5369 (N_5369,N_4915,N_4824);
nor U5370 (N_5370,N_4511,N_4820);
or U5371 (N_5371,N_4815,N_4523);
or U5372 (N_5372,N_4902,N_4705);
or U5373 (N_5373,N_4767,N_4525);
nor U5374 (N_5374,N_4935,N_4881);
xor U5375 (N_5375,N_4593,N_4747);
nand U5376 (N_5376,N_4595,N_4820);
nor U5377 (N_5377,N_4851,N_4861);
nand U5378 (N_5378,N_4629,N_4671);
nor U5379 (N_5379,N_4872,N_4568);
or U5380 (N_5380,N_4564,N_4886);
xnor U5381 (N_5381,N_4881,N_4966);
and U5382 (N_5382,N_4947,N_4686);
xor U5383 (N_5383,N_4567,N_4883);
nand U5384 (N_5384,N_4787,N_4727);
and U5385 (N_5385,N_4792,N_4508);
nand U5386 (N_5386,N_4669,N_4845);
nor U5387 (N_5387,N_4908,N_4637);
nor U5388 (N_5388,N_4509,N_4786);
xnor U5389 (N_5389,N_4737,N_4711);
xnor U5390 (N_5390,N_4916,N_4817);
or U5391 (N_5391,N_4748,N_4776);
and U5392 (N_5392,N_4736,N_4572);
and U5393 (N_5393,N_4583,N_4801);
and U5394 (N_5394,N_4619,N_4660);
or U5395 (N_5395,N_4824,N_4822);
nand U5396 (N_5396,N_4651,N_4963);
xnor U5397 (N_5397,N_4938,N_4500);
nand U5398 (N_5398,N_4865,N_4906);
or U5399 (N_5399,N_4741,N_4599);
xnor U5400 (N_5400,N_4554,N_4926);
nor U5401 (N_5401,N_4750,N_4609);
or U5402 (N_5402,N_4852,N_4572);
nand U5403 (N_5403,N_4922,N_4930);
or U5404 (N_5404,N_4646,N_4978);
or U5405 (N_5405,N_4884,N_4989);
nand U5406 (N_5406,N_4846,N_4523);
or U5407 (N_5407,N_4948,N_4815);
nor U5408 (N_5408,N_4798,N_4954);
xnor U5409 (N_5409,N_4565,N_4748);
or U5410 (N_5410,N_4715,N_4557);
nand U5411 (N_5411,N_4794,N_4945);
nor U5412 (N_5412,N_4775,N_4930);
xnor U5413 (N_5413,N_4645,N_4671);
xor U5414 (N_5414,N_4755,N_4814);
nor U5415 (N_5415,N_4995,N_4819);
or U5416 (N_5416,N_4808,N_4781);
xnor U5417 (N_5417,N_4912,N_4994);
nor U5418 (N_5418,N_4796,N_4870);
and U5419 (N_5419,N_4556,N_4878);
nand U5420 (N_5420,N_4883,N_4797);
or U5421 (N_5421,N_4519,N_4588);
nand U5422 (N_5422,N_4571,N_4542);
nand U5423 (N_5423,N_4686,N_4892);
nor U5424 (N_5424,N_4966,N_4800);
and U5425 (N_5425,N_4891,N_4967);
xnor U5426 (N_5426,N_4888,N_4875);
nand U5427 (N_5427,N_4875,N_4765);
nor U5428 (N_5428,N_4885,N_4571);
xnor U5429 (N_5429,N_4741,N_4903);
nand U5430 (N_5430,N_4790,N_4502);
xor U5431 (N_5431,N_4849,N_4786);
nand U5432 (N_5432,N_4909,N_4640);
and U5433 (N_5433,N_4842,N_4831);
nand U5434 (N_5434,N_4685,N_4605);
nand U5435 (N_5435,N_4678,N_4728);
or U5436 (N_5436,N_4907,N_4826);
or U5437 (N_5437,N_4758,N_4858);
nor U5438 (N_5438,N_4653,N_4696);
or U5439 (N_5439,N_4666,N_4710);
xor U5440 (N_5440,N_4611,N_4958);
and U5441 (N_5441,N_4670,N_4635);
or U5442 (N_5442,N_4748,N_4892);
xor U5443 (N_5443,N_4660,N_4605);
nand U5444 (N_5444,N_4718,N_4840);
or U5445 (N_5445,N_4985,N_4524);
or U5446 (N_5446,N_4552,N_4668);
nor U5447 (N_5447,N_4715,N_4667);
nand U5448 (N_5448,N_4859,N_4649);
and U5449 (N_5449,N_4584,N_4810);
nand U5450 (N_5450,N_4833,N_4684);
and U5451 (N_5451,N_4822,N_4813);
and U5452 (N_5452,N_4521,N_4953);
xnor U5453 (N_5453,N_4798,N_4506);
xnor U5454 (N_5454,N_4788,N_4822);
and U5455 (N_5455,N_4958,N_4966);
and U5456 (N_5456,N_4785,N_4930);
nor U5457 (N_5457,N_4892,N_4715);
xor U5458 (N_5458,N_4587,N_4882);
or U5459 (N_5459,N_4985,N_4977);
or U5460 (N_5460,N_4719,N_4982);
xor U5461 (N_5461,N_4603,N_4541);
or U5462 (N_5462,N_4585,N_4598);
xnor U5463 (N_5463,N_4696,N_4753);
or U5464 (N_5464,N_4875,N_4555);
or U5465 (N_5465,N_4544,N_4597);
nand U5466 (N_5466,N_4633,N_4831);
and U5467 (N_5467,N_4915,N_4981);
and U5468 (N_5468,N_4951,N_4766);
or U5469 (N_5469,N_4796,N_4861);
xnor U5470 (N_5470,N_4797,N_4813);
and U5471 (N_5471,N_4972,N_4811);
nand U5472 (N_5472,N_4796,N_4708);
and U5473 (N_5473,N_4662,N_4541);
nor U5474 (N_5474,N_4974,N_4604);
and U5475 (N_5475,N_4741,N_4563);
nand U5476 (N_5476,N_4559,N_4926);
xor U5477 (N_5477,N_4924,N_4902);
nor U5478 (N_5478,N_4707,N_4501);
or U5479 (N_5479,N_4705,N_4572);
nand U5480 (N_5480,N_4782,N_4731);
or U5481 (N_5481,N_4847,N_4836);
and U5482 (N_5482,N_4832,N_4848);
or U5483 (N_5483,N_4589,N_4971);
or U5484 (N_5484,N_4792,N_4949);
nand U5485 (N_5485,N_4921,N_4889);
nand U5486 (N_5486,N_4670,N_4719);
xor U5487 (N_5487,N_4977,N_4561);
and U5488 (N_5488,N_4600,N_4566);
and U5489 (N_5489,N_4870,N_4662);
or U5490 (N_5490,N_4608,N_4552);
and U5491 (N_5491,N_4630,N_4614);
and U5492 (N_5492,N_4503,N_4557);
or U5493 (N_5493,N_4629,N_4861);
nor U5494 (N_5494,N_4669,N_4946);
nor U5495 (N_5495,N_4887,N_4874);
or U5496 (N_5496,N_4930,N_4946);
and U5497 (N_5497,N_4763,N_4760);
or U5498 (N_5498,N_4813,N_4757);
xor U5499 (N_5499,N_4999,N_4890);
nor U5500 (N_5500,N_5074,N_5177);
nor U5501 (N_5501,N_5473,N_5362);
or U5502 (N_5502,N_5301,N_5185);
or U5503 (N_5503,N_5332,N_5309);
xor U5504 (N_5504,N_5068,N_5495);
nand U5505 (N_5505,N_5337,N_5042);
nor U5506 (N_5506,N_5345,N_5475);
nor U5507 (N_5507,N_5207,N_5160);
and U5508 (N_5508,N_5147,N_5210);
xnor U5509 (N_5509,N_5357,N_5298);
xor U5510 (N_5510,N_5025,N_5150);
nand U5511 (N_5511,N_5391,N_5233);
nor U5512 (N_5512,N_5130,N_5053);
xnor U5513 (N_5513,N_5248,N_5272);
nor U5514 (N_5514,N_5215,N_5313);
nor U5515 (N_5515,N_5259,N_5013);
xor U5516 (N_5516,N_5398,N_5026);
xnor U5517 (N_5517,N_5111,N_5359);
or U5518 (N_5518,N_5224,N_5247);
or U5519 (N_5519,N_5153,N_5446);
nor U5520 (N_5520,N_5031,N_5269);
nand U5521 (N_5521,N_5331,N_5354);
and U5522 (N_5522,N_5209,N_5494);
nand U5523 (N_5523,N_5389,N_5034);
xor U5524 (N_5524,N_5285,N_5282);
or U5525 (N_5525,N_5452,N_5418);
and U5526 (N_5526,N_5484,N_5387);
nor U5527 (N_5527,N_5135,N_5087);
and U5528 (N_5528,N_5325,N_5465);
or U5529 (N_5529,N_5107,N_5024);
xnor U5530 (N_5530,N_5226,N_5208);
nor U5531 (N_5531,N_5214,N_5098);
or U5532 (N_5532,N_5374,N_5052);
nand U5533 (N_5533,N_5295,N_5411);
or U5534 (N_5534,N_5291,N_5463);
or U5535 (N_5535,N_5032,N_5275);
nor U5536 (N_5536,N_5134,N_5441);
and U5537 (N_5537,N_5403,N_5381);
xnor U5538 (N_5538,N_5496,N_5137);
or U5539 (N_5539,N_5008,N_5288);
nand U5540 (N_5540,N_5405,N_5334);
or U5541 (N_5541,N_5469,N_5430);
and U5542 (N_5542,N_5290,N_5459);
nor U5543 (N_5543,N_5448,N_5447);
and U5544 (N_5544,N_5300,N_5478);
or U5545 (N_5545,N_5343,N_5439);
or U5546 (N_5546,N_5193,N_5167);
xor U5547 (N_5547,N_5165,N_5280);
and U5548 (N_5548,N_5170,N_5457);
and U5549 (N_5549,N_5372,N_5219);
and U5550 (N_5550,N_5241,N_5262);
nand U5551 (N_5551,N_5318,N_5489);
and U5552 (N_5552,N_5302,N_5242);
and U5553 (N_5553,N_5162,N_5213);
or U5554 (N_5554,N_5133,N_5472);
or U5555 (N_5555,N_5234,N_5428);
nor U5556 (N_5556,N_5455,N_5218);
xor U5557 (N_5557,N_5483,N_5037);
nand U5558 (N_5558,N_5294,N_5283);
and U5559 (N_5559,N_5067,N_5148);
xor U5560 (N_5560,N_5270,N_5046);
xor U5561 (N_5561,N_5047,N_5183);
or U5562 (N_5562,N_5073,N_5278);
nand U5563 (N_5563,N_5279,N_5268);
nor U5564 (N_5564,N_5438,N_5474);
or U5565 (N_5565,N_5012,N_5471);
nand U5566 (N_5566,N_5349,N_5249);
nand U5567 (N_5567,N_5161,N_5485);
xnor U5568 (N_5568,N_5124,N_5456);
nand U5569 (N_5569,N_5079,N_5009);
or U5570 (N_5570,N_5492,N_5103);
or U5571 (N_5571,N_5036,N_5138);
nand U5572 (N_5572,N_5392,N_5344);
xor U5573 (N_5573,N_5450,N_5369);
or U5574 (N_5574,N_5432,N_5289);
and U5575 (N_5575,N_5159,N_5466);
and U5576 (N_5576,N_5144,N_5017);
xor U5577 (N_5577,N_5035,N_5368);
nor U5578 (N_5578,N_5329,N_5001);
xnor U5579 (N_5579,N_5149,N_5250);
or U5580 (N_5580,N_5297,N_5397);
nor U5581 (N_5581,N_5422,N_5314);
or U5582 (N_5582,N_5077,N_5018);
or U5583 (N_5583,N_5386,N_5184);
xnor U5584 (N_5584,N_5075,N_5099);
nand U5585 (N_5585,N_5253,N_5066);
nand U5586 (N_5586,N_5311,N_5276);
xnor U5587 (N_5587,N_5409,N_5376);
nor U5588 (N_5588,N_5102,N_5493);
nand U5589 (N_5589,N_5072,N_5257);
nand U5590 (N_5590,N_5022,N_5251);
nor U5591 (N_5591,N_5261,N_5190);
and U5592 (N_5592,N_5330,N_5277);
and U5593 (N_5593,N_5360,N_5015);
or U5594 (N_5594,N_5464,N_5058);
xnor U5595 (N_5595,N_5267,N_5142);
nand U5596 (N_5596,N_5129,N_5141);
or U5597 (N_5597,N_5188,N_5217);
nor U5598 (N_5598,N_5014,N_5027);
nand U5599 (N_5599,N_5019,N_5479);
or U5600 (N_5600,N_5481,N_5000);
nor U5601 (N_5601,N_5310,N_5429);
nand U5602 (N_5602,N_5399,N_5467);
or U5603 (N_5603,N_5400,N_5445);
xnor U5604 (N_5604,N_5069,N_5348);
xnor U5605 (N_5605,N_5361,N_5131);
or U5606 (N_5606,N_5462,N_5336);
and U5607 (N_5607,N_5238,N_5100);
xor U5608 (N_5608,N_5119,N_5341);
xnor U5609 (N_5609,N_5440,N_5086);
or U5610 (N_5610,N_5023,N_5151);
xnor U5611 (N_5611,N_5319,N_5179);
nor U5612 (N_5612,N_5090,N_5375);
and U5613 (N_5613,N_5181,N_5454);
nor U5614 (N_5614,N_5449,N_5394);
nand U5615 (N_5615,N_5002,N_5385);
and U5616 (N_5616,N_5342,N_5164);
or U5617 (N_5617,N_5211,N_5174);
xnor U5618 (N_5618,N_5007,N_5266);
xnor U5619 (N_5619,N_5114,N_5414);
nand U5620 (N_5620,N_5488,N_5155);
nand U5621 (N_5621,N_5132,N_5196);
nor U5622 (N_5622,N_5158,N_5194);
or U5623 (N_5623,N_5109,N_5338);
nand U5624 (N_5624,N_5021,N_5085);
nand U5625 (N_5625,N_5482,N_5029);
nand U5626 (N_5626,N_5306,N_5367);
nor U5627 (N_5627,N_5435,N_5444);
nand U5628 (N_5628,N_5486,N_5157);
nor U5629 (N_5629,N_5355,N_5237);
nor U5630 (N_5630,N_5358,N_5413);
nand U5631 (N_5631,N_5143,N_5117);
nor U5632 (N_5632,N_5062,N_5421);
and U5633 (N_5633,N_5323,N_5402);
nor U5634 (N_5634,N_5458,N_5433);
and U5635 (N_5635,N_5044,N_5078);
and U5636 (N_5636,N_5426,N_5083);
and U5637 (N_5637,N_5178,N_5121);
nand U5638 (N_5638,N_5120,N_5057);
or U5639 (N_5639,N_5470,N_5437);
xnor U5640 (N_5640,N_5168,N_5038);
and U5641 (N_5641,N_5407,N_5351);
nor U5642 (N_5642,N_5112,N_5113);
or U5643 (N_5643,N_5200,N_5171);
and U5644 (N_5644,N_5420,N_5145);
and U5645 (N_5645,N_5404,N_5419);
nor U5646 (N_5646,N_5118,N_5427);
xor U5647 (N_5647,N_5051,N_5384);
and U5648 (N_5648,N_5232,N_5461);
and U5649 (N_5649,N_5274,N_5222);
or U5650 (N_5650,N_5371,N_5223);
and U5651 (N_5651,N_5497,N_5287);
nor U5652 (N_5652,N_5380,N_5182);
xnor U5653 (N_5653,N_5216,N_5322);
nand U5654 (N_5654,N_5230,N_5070);
or U5655 (N_5655,N_5154,N_5401);
xnor U5656 (N_5656,N_5366,N_5108);
nor U5657 (N_5657,N_5095,N_5317);
and U5658 (N_5658,N_5240,N_5383);
or U5659 (N_5659,N_5056,N_5370);
or U5660 (N_5660,N_5030,N_5417);
or U5661 (N_5661,N_5408,N_5172);
xnor U5662 (N_5662,N_5228,N_5498);
xnor U5663 (N_5663,N_5415,N_5064);
and U5664 (N_5664,N_5186,N_5254);
and U5665 (N_5665,N_5442,N_5166);
nand U5666 (N_5666,N_5049,N_5097);
nor U5667 (N_5667,N_5229,N_5451);
or U5668 (N_5668,N_5378,N_5203);
xnor U5669 (N_5669,N_5156,N_5106);
nand U5670 (N_5670,N_5255,N_5239);
or U5671 (N_5671,N_5431,N_5252);
xnor U5672 (N_5672,N_5406,N_5333);
nand U5673 (N_5673,N_5221,N_5076);
and U5674 (N_5674,N_5122,N_5003);
xor U5675 (N_5675,N_5412,N_5101);
xnor U5676 (N_5676,N_5390,N_5220);
xor U5677 (N_5677,N_5041,N_5180);
xor U5678 (N_5678,N_5443,N_5416);
or U5679 (N_5679,N_5352,N_5199);
nor U5680 (N_5680,N_5006,N_5340);
nor U5681 (N_5681,N_5312,N_5246);
nand U5682 (N_5682,N_5243,N_5175);
or U5683 (N_5683,N_5296,N_5189);
nand U5684 (N_5684,N_5128,N_5080);
nand U5685 (N_5685,N_5096,N_5460);
nand U5686 (N_5686,N_5324,N_5225);
and U5687 (N_5687,N_5396,N_5191);
nand U5688 (N_5688,N_5263,N_5105);
nor U5689 (N_5689,N_5089,N_5010);
xor U5690 (N_5690,N_5045,N_5258);
and U5691 (N_5691,N_5163,N_5260);
and U5692 (N_5692,N_5011,N_5491);
nor U5693 (N_5693,N_5304,N_5476);
nor U5694 (N_5694,N_5126,N_5016);
and U5695 (N_5695,N_5264,N_5192);
nor U5696 (N_5696,N_5071,N_5088);
or U5697 (N_5697,N_5028,N_5212);
nor U5698 (N_5698,N_5245,N_5499);
and U5699 (N_5699,N_5227,N_5256);
nor U5700 (N_5700,N_5379,N_5365);
nand U5701 (N_5701,N_5307,N_5235);
nand U5702 (N_5702,N_5202,N_5423);
nor U5703 (N_5703,N_5265,N_5061);
or U5704 (N_5704,N_5326,N_5104);
nand U5705 (N_5705,N_5043,N_5315);
xnor U5706 (N_5706,N_5048,N_5286);
nor U5707 (N_5707,N_5020,N_5198);
nand U5708 (N_5708,N_5284,N_5335);
or U5709 (N_5709,N_5373,N_5356);
nor U5710 (N_5710,N_5139,N_5092);
and U5711 (N_5711,N_5115,N_5195);
or U5712 (N_5712,N_5173,N_5350);
and U5713 (N_5713,N_5271,N_5059);
or U5714 (N_5714,N_5039,N_5136);
nor U5715 (N_5715,N_5410,N_5346);
nand U5716 (N_5716,N_5093,N_5127);
or U5717 (N_5717,N_5377,N_5424);
xor U5718 (N_5718,N_5197,N_5110);
nor U5719 (N_5719,N_5084,N_5303);
nand U5720 (N_5720,N_5004,N_5205);
or U5721 (N_5721,N_5339,N_5204);
nor U5722 (N_5722,N_5065,N_5187);
nor U5723 (N_5723,N_5347,N_5328);
or U5724 (N_5724,N_5054,N_5395);
or U5725 (N_5725,N_5176,N_5244);
nand U5726 (N_5726,N_5055,N_5094);
and U5727 (N_5727,N_5382,N_5081);
and U5728 (N_5728,N_5363,N_5123);
nor U5729 (N_5729,N_5140,N_5434);
nor U5730 (N_5730,N_5453,N_5480);
and U5731 (N_5731,N_5468,N_5146);
or U5732 (N_5732,N_5425,N_5033);
xnor U5733 (N_5733,N_5321,N_5231);
xor U5734 (N_5734,N_5169,N_5236);
nor U5735 (N_5735,N_5281,N_5299);
nand U5736 (N_5736,N_5327,N_5353);
nand U5737 (N_5737,N_5125,N_5364);
xnor U5738 (N_5738,N_5091,N_5477);
and U5739 (N_5739,N_5082,N_5201);
or U5740 (N_5740,N_5436,N_5305);
or U5741 (N_5741,N_5206,N_5293);
nand U5742 (N_5742,N_5273,N_5320);
and U5743 (N_5743,N_5393,N_5152);
nor U5744 (N_5744,N_5292,N_5040);
and U5745 (N_5745,N_5116,N_5316);
and U5746 (N_5746,N_5005,N_5060);
xnor U5747 (N_5747,N_5388,N_5050);
and U5748 (N_5748,N_5063,N_5490);
or U5749 (N_5749,N_5487,N_5308);
nor U5750 (N_5750,N_5379,N_5262);
xor U5751 (N_5751,N_5342,N_5336);
or U5752 (N_5752,N_5090,N_5278);
nand U5753 (N_5753,N_5005,N_5462);
and U5754 (N_5754,N_5440,N_5057);
and U5755 (N_5755,N_5056,N_5472);
nand U5756 (N_5756,N_5358,N_5337);
nor U5757 (N_5757,N_5491,N_5216);
or U5758 (N_5758,N_5326,N_5144);
xnor U5759 (N_5759,N_5087,N_5219);
nand U5760 (N_5760,N_5141,N_5046);
and U5761 (N_5761,N_5123,N_5138);
nor U5762 (N_5762,N_5378,N_5466);
nor U5763 (N_5763,N_5313,N_5059);
or U5764 (N_5764,N_5241,N_5080);
xnor U5765 (N_5765,N_5360,N_5158);
or U5766 (N_5766,N_5026,N_5050);
nand U5767 (N_5767,N_5345,N_5494);
and U5768 (N_5768,N_5235,N_5423);
and U5769 (N_5769,N_5493,N_5458);
nor U5770 (N_5770,N_5333,N_5342);
and U5771 (N_5771,N_5183,N_5303);
nor U5772 (N_5772,N_5041,N_5108);
nor U5773 (N_5773,N_5004,N_5363);
nand U5774 (N_5774,N_5299,N_5056);
and U5775 (N_5775,N_5166,N_5279);
nor U5776 (N_5776,N_5014,N_5419);
or U5777 (N_5777,N_5153,N_5110);
and U5778 (N_5778,N_5225,N_5081);
and U5779 (N_5779,N_5317,N_5396);
xnor U5780 (N_5780,N_5398,N_5473);
xor U5781 (N_5781,N_5260,N_5065);
and U5782 (N_5782,N_5462,N_5205);
xnor U5783 (N_5783,N_5203,N_5093);
or U5784 (N_5784,N_5143,N_5355);
nand U5785 (N_5785,N_5100,N_5157);
or U5786 (N_5786,N_5273,N_5032);
and U5787 (N_5787,N_5268,N_5092);
nand U5788 (N_5788,N_5398,N_5063);
or U5789 (N_5789,N_5352,N_5407);
or U5790 (N_5790,N_5305,N_5116);
or U5791 (N_5791,N_5154,N_5261);
xnor U5792 (N_5792,N_5216,N_5129);
nor U5793 (N_5793,N_5165,N_5279);
or U5794 (N_5794,N_5398,N_5165);
nand U5795 (N_5795,N_5217,N_5011);
or U5796 (N_5796,N_5157,N_5150);
xor U5797 (N_5797,N_5153,N_5282);
or U5798 (N_5798,N_5037,N_5081);
nand U5799 (N_5799,N_5064,N_5418);
and U5800 (N_5800,N_5223,N_5249);
and U5801 (N_5801,N_5434,N_5300);
xor U5802 (N_5802,N_5081,N_5077);
or U5803 (N_5803,N_5025,N_5107);
xor U5804 (N_5804,N_5185,N_5429);
nand U5805 (N_5805,N_5294,N_5160);
nand U5806 (N_5806,N_5412,N_5348);
and U5807 (N_5807,N_5414,N_5037);
nor U5808 (N_5808,N_5365,N_5206);
or U5809 (N_5809,N_5405,N_5414);
nand U5810 (N_5810,N_5191,N_5375);
xnor U5811 (N_5811,N_5418,N_5073);
and U5812 (N_5812,N_5098,N_5494);
nand U5813 (N_5813,N_5416,N_5468);
nor U5814 (N_5814,N_5336,N_5124);
nand U5815 (N_5815,N_5258,N_5123);
nand U5816 (N_5816,N_5468,N_5108);
nand U5817 (N_5817,N_5011,N_5115);
xnor U5818 (N_5818,N_5300,N_5051);
and U5819 (N_5819,N_5384,N_5105);
and U5820 (N_5820,N_5387,N_5226);
nor U5821 (N_5821,N_5254,N_5304);
and U5822 (N_5822,N_5387,N_5194);
nand U5823 (N_5823,N_5486,N_5450);
nand U5824 (N_5824,N_5363,N_5239);
xor U5825 (N_5825,N_5160,N_5300);
or U5826 (N_5826,N_5163,N_5289);
nor U5827 (N_5827,N_5465,N_5378);
or U5828 (N_5828,N_5249,N_5014);
nand U5829 (N_5829,N_5059,N_5223);
or U5830 (N_5830,N_5245,N_5343);
xnor U5831 (N_5831,N_5331,N_5018);
nor U5832 (N_5832,N_5115,N_5448);
nor U5833 (N_5833,N_5299,N_5249);
xor U5834 (N_5834,N_5272,N_5402);
xor U5835 (N_5835,N_5100,N_5312);
nand U5836 (N_5836,N_5254,N_5311);
nand U5837 (N_5837,N_5284,N_5087);
or U5838 (N_5838,N_5465,N_5171);
xnor U5839 (N_5839,N_5440,N_5138);
xnor U5840 (N_5840,N_5376,N_5059);
nand U5841 (N_5841,N_5486,N_5329);
or U5842 (N_5842,N_5410,N_5162);
nor U5843 (N_5843,N_5044,N_5376);
xor U5844 (N_5844,N_5195,N_5104);
or U5845 (N_5845,N_5158,N_5196);
nand U5846 (N_5846,N_5454,N_5424);
xor U5847 (N_5847,N_5284,N_5494);
xor U5848 (N_5848,N_5309,N_5259);
xnor U5849 (N_5849,N_5379,N_5490);
nand U5850 (N_5850,N_5004,N_5031);
or U5851 (N_5851,N_5094,N_5481);
xor U5852 (N_5852,N_5444,N_5261);
and U5853 (N_5853,N_5136,N_5210);
and U5854 (N_5854,N_5377,N_5490);
or U5855 (N_5855,N_5417,N_5261);
nor U5856 (N_5856,N_5334,N_5286);
and U5857 (N_5857,N_5208,N_5214);
xnor U5858 (N_5858,N_5048,N_5182);
nor U5859 (N_5859,N_5177,N_5135);
nor U5860 (N_5860,N_5181,N_5227);
and U5861 (N_5861,N_5071,N_5365);
nor U5862 (N_5862,N_5406,N_5328);
nand U5863 (N_5863,N_5401,N_5159);
and U5864 (N_5864,N_5441,N_5060);
nand U5865 (N_5865,N_5302,N_5095);
and U5866 (N_5866,N_5069,N_5427);
nand U5867 (N_5867,N_5144,N_5204);
nand U5868 (N_5868,N_5174,N_5106);
or U5869 (N_5869,N_5009,N_5250);
xnor U5870 (N_5870,N_5365,N_5450);
or U5871 (N_5871,N_5377,N_5114);
or U5872 (N_5872,N_5129,N_5361);
nor U5873 (N_5873,N_5029,N_5256);
nand U5874 (N_5874,N_5003,N_5373);
nand U5875 (N_5875,N_5046,N_5452);
xor U5876 (N_5876,N_5088,N_5132);
nand U5877 (N_5877,N_5354,N_5272);
xor U5878 (N_5878,N_5003,N_5210);
nor U5879 (N_5879,N_5167,N_5434);
xor U5880 (N_5880,N_5442,N_5458);
and U5881 (N_5881,N_5322,N_5430);
xor U5882 (N_5882,N_5020,N_5291);
nor U5883 (N_5883,N_5407,N_5243);
xor U5884 (N_5884,N_5093,N_5083);
or U5885 (N_5885,N_5424,N_5194);
or U5886 (N_5886,N_5089,N_5020);
nand U5887 (N_5887,N_5021,N_5254);
or U5888 (N_5888,N_5209,N_5166);
nand U5889 (N_5889,N_5084,N_5328);
and U5890 (N_5890,N_5027,N_5491);
or U5891 (N_5891,N_5336,N_5067);
nor U5892 (N_5892,N_5191,N_5478);
nor U5893 (N_5893,N_5074,N_5001);
or U5894 (N_5894,N_5006,N_5014);
nor U5895 (N_5895,N_5345,N_5399);
xor U5896 (N_5896,N_5072,N_5108);
or U5897 (N_5897,N_5275,N_5139);
and U5898 (N_5898,N_5235,N_5358);
and U5899 (N_5899,N_5434,N_5050);
or U5900 (N_5900,N_5188,N_5229);
xnor U5901 (N_5901,N_5366,N_5493);
or U5902 (N_5902,N_5210,N_5046);
and U5903 (N_5903,N_5476,N_5391);
nand U5904 (N_5904,N_5434,N_5384);
nand U5905 (N_5905,N_5003,N_5206);
and U5906 (N_5906,N_5010,N_5212);
or U5907 (N_5907,N_5451,N_5361);
nor U5908 (N_5908,N_5183,N_5102);
nand U5909 (N_5909,N_5225,N_5420);
and U5910 (N_5910,N_5403,N_5407);
xnor U5911 (N_5911,N_5376,N_5372);
and U5912 (N_5912,N_5429,N_5450);
and U5913 (N_5913,N_5073,N_5072);
nor U5914 (N_5914,N_5013,N_5485);
nor U5915 (N_5915,N_5218,N_5056);
and U5916 (N_5916,N_5464,N_5133);
nand U5917 (N_5917,N_5301,N_5203);
and U5918 (N_5918,N_5243,N_5397);
or U5919 (N_5919,N_5422,N_5378);
nor U5920 (N_5920,N_5065,N_5327);
nand U5921 (N_5921,N_5483,N_5439);
or U5922 (N_5922,N_5014,N_5216);
or U5923 (N_5923,N_5256,N_5238);
nor U5924 (N_5924,N_5492,N_5479);
and U5925 (N_5925,N_5299,N_5278);
or U5926 (N_5926,N_5366,N_5135);
xor U5927 (N_5927,N_5232,N_5340);
nor U5928 (N_5928,N_5214,N_5106);
or U5929 (N_5929,N_5412,N_5330);
xor U5930 (N_5930,N_5272,N_5400);
nor U5931 (N_5931,N_5072,N_5097);
nor U5932 (N_5932,N_5393,N_5415);
or U5933 (N_5933,N_5357,N_5274);
xnor U5934 (N_5934,N_5279,N_5041);
and U5935 (N_5935,N_5104,N_5181);
nor U5936 (N_5936,N_5019,N_5062);
and U5937 (N_5937,N_5238,N_5411);
and U5938 (N_5938,N_5130,N_5332);
nor U5939 (N_5939,N_5458,N_5393);
xnor U5940 (N_5940,N_5265,N_5444);
nor U5941 (N_5941,N_5273,N_5248);
and U5942 (N_5942,N_5051,N_5261);
nor U5943 (N_5943,N_5492,N_5163);
and U5944 (N_5944,N_5238,N_5015);
nand U5945 (N_5945,N_5130,N_5423);
xnor U5946 (N_5946,N_5365,N_5349);
and U5947 (N_5947,N_5175,N_5487);
xor U5948 (N_5948,N_5023,N_5346);
xnor U5949 (N_5949,N_5239,N_5289);
xnor U5950 (N_5950,N_5187,N_5034);
xor U5951 (N_5951,N_5305,N_5106);
nor U5952 (N_5952,N_5477,N_5249);
nand U5953 (N_5953,N_5319,N_5239);
and U5954 (N_5954,N_5030,N_5170);
or U5955 (N_5955,N_5221,N_5228);
nor U5956 (N_5956,N_5463,N_5402);
nand U5957 (N_5957,N_5461,N_5158);
nand U5958 (N_5958,N_5202,N_5103);
xor U5959 (N_5959,N_5449,N_5483);
xnor U5960 (N_5960,N_5210,N_5275);
xnor U5961 (N_5961,N_5158,N_5179);
nand U5962 (N_5962,N_5187,N_5161);
nor U5963 (N_5963,N_5110,N_5240);
and U5964 (N_5964,N_5285,N_5003);
or U5965 (N_5965,N_5144,N_5309);
or U5966 (N_5966,N_5297,N_5017);
nand U5967 (N_5967,N_5107,N_5160);
nand U5968 (N_5968,N_5494,N_5479);
nand U5969 (N_5969,N_5210,N_5378);
nand U5970 (N_5970,N_5229,N_5107);
xor U5971 (N_5971,N_5195,N_5444);
xor U5972 (N_5972,N_5278,N_5114);
or U5973 (N_5973,N_5471,N_5445);
xor U5974 (N_5974,N_5269,N_5009);
or U5975 (N_5975,N_5060,N_5306);
xor U5976 (N_5976,N_5307,N_5398);
or U5977 (N_5977,N_5174,N_5130);
xor U5978 (N_5978,N_5337,N_5021);
nor U5979 (N_5979,N_5416,N_5007);
or U5980 (N_5980,N_5025,N_5363);
nand U5981 (N_5981,N_5267,N_5242);
xor U5982 (N_5982,N_5342,N_5039);
or U5983 (N_5983,N_5056,N_5102);
nand U5984 (N_5984,N_5255,N_5065);
xnor U5985 (N_5985,N_5150,N_5151);
or U5986 (N_5986,N_5359,N_5227);
nand U5987 (N_5987,N_5052,N_5107);
nand U5988 (N_5988,N_5321,N_5039);
and U5989 (N_5989,N_5466,N_5176);
nand U5990 (N_5990,N_5213,N_5011);
xnor U5991 (N_5991,N_5303,N_5160);
xnor U5992 (N_5992,N_5189,N_5019);
xor U5993 (N_5993,N_5107,N_5406);
and U5994 (N_5994,N_5345,N_5105);
or U5995 (N_5995,N_5198,N_5035);
nor U5996 (N_5996,N_5421,N_5462);
or U5997 (N_5997,N_5208,N_5410);
nand U5998 (N_5998,N_5444,N_5250);
xnor U5999 (N_5999,N_5209,N_5219);
nand U6000 (N_6000,N_5610,N_5981);
and U6001 (N_6001,N_5502,N_5760);
nor U6002 (N_6002,N_5511,N_5904);
or U6003 (N_6003,N_5975,N_5902);
nor U6004 (N_6004,N_5849,N_5688);
nand U6005 (N_6005,N_5879,N_5890);
and U6006 (N_6006,N_5757,N_5747);
nor U6007 (N_6007,N_5834,N_5977);
xor U6008 (N_6008,N_5785,N_5826);
or U6009 (N_6009,N_5664,N_5632);
or U6010 (N_6010,N_5952,N_5573);
nand U6011 (N_6011,N_5930,N_5889);
xor U6012 (N_6012,N_5940,N_5579);
or U6013 (N_6013,N_5651,N_5780);
nor U6014 (N_6014,N_5836,N_5711);
xor U6015 (N_6015,N_5583,N_5729);
nor U6016 (N_6016,N_5841,N_5983);
nand U6017 (N_6017,N_5698,N_5553);
nand U6018 (N_6018,N_5700,N_5779);
nand U6019 (N_6019,N_5876,N_5936);
and U6020 (N_6020,N_5860,N_5787);
and U6021 (N_6021,N_5717,N_5942);
nor U6022 (N_6022,N_5689,N_5964);
and U6023 (N_6023,N_5781,N_5675);
or U6024 (N_6024,N_5840,N_5907);
nor U6025 (N_6025,N_5997,N_5674);
nand U6026 (N_6026,N_5850,N_5925);
nor U6027 (N_6027,N_5799,N_5802);
nand U6028 (N_6028,N_5636,N_5772);
nor U6029 (N_6029,N_5784,N_5692);
nor U6030 (N_6030,N_5814,N_5533);
and U6031 (N_6031,N_5595,N_5775);
nor U6032 (N_6032,N_5974,N_5594);
nor U6033 (N_6033,N_5920,N_5527);
or U6034 (N_6034,N_5627,N_5833);
and U6035 (N_6035,N_5823,N_5629);
and U6036 (N_6036,N_5791,N_5869);
nand U6037 (N_6037,N_5807,N_5572);
and U6038 (N_6038,N_5909,N_5864);
nand U6039 (N_6039,N_5770,N_5678);
xnor U6040 (N_6040,N_5885,N_5846);
or U6041 (N_6041,N_5642,N_5880);
xor U6042 (N_6042,N_5819,N_5894);
nand U6043 (N_6043,N_5985,N_5600);
and U6044 (N_6044,N_5928,N_5835);
and U6045 (N_6045,N_5701,N_5788);
nand U6046 (N_6046,N_5559,N_5858);
xnor U6047 (N_6047,N_5822,N_5503);
and U6048 (N_6048,N_5910,N_5883);
xor U6049 (N_6049,N_5721,N_5662);
nor U6050 (N_6050,N_5980,N_5839);
and U6051 (N_6051,N_5914,N_5805);
and U6052 (N_6052,N_5815,N_5963);
xnor U6053 (N_6053,N_5665,N_5808);
or U6054 (N_6054,N_5545,N_5803);
nor U6055 (N_6055,N_5725,N_5953);
or U6056 (N_6056,N_5608,N_5580);
or U6057 (N_6057,N_5856,N_5599);
and U6058 (N_6058,N_5901,N_5626);
or U6059 (N_6059,N_5562,N_5602);
or U6060 (N_6060,N_5965,N_5640);
and U6061 (N_6061,N_5549,N_5882);
xor U6062 (N_6062,N_5565,N_5761);
xor U6063 (N_6063,N_5581,N_5796);
or U6064 (N_6064,N_5520,N_5794);
or U6065 (N_6065,N_5989,N_5857);
nor U6066 (N_6066,N_5946,N_5624);
and U6067 (N_6067,N_5704,N_5886);
and U6068 (N_6068,N_5500,N_5530);
and U6069 (N_6069,N_5638,N_5673);
and U6070 (N_6070,N_5749,N_5646);
and U6071 (N_6071,N_5881,N_5709);
or U6072 (N_6072,N_5793,N_5978);
xor U6073 (N_6073,N_5712,N_5877);
xnor U6074 (N_6074,N_5604,N_5871);
nand U6075 (N_6075,N_5995,N_5728);
nand U6076 (N_6076,N_5681,N_5738);
xor U6077 (N_6077,N_5617,N_5816);
xnor U6078 (N_6078,N_5903,N_5691);
and U6079 (N_6079,N_5552,N_5654);
nand U6080 (N_6080,N_5526,N_5777);
xor U6081 (N_6081,N_5515,N_5518);
nand U6082 (N_6082,N_5628,N_5534);
nand U6083 (N_6083,N_5702,N_5919);
and U6084 (N_6084,N_5843,N_5618);
nor U6085 (N_6085,N_5611,N_5911);
nand U6086 (N_6086,N_5862,N_5873);
nand U6087 (N_6087,N_5731,N_5897);
xnor U6088 (N_6088,N_5748,N_5750);
nand U6089 (N_6089,N_5842,N_5999);
and U6090 (N_6090,N_5888,N_5720);
nor U6091 (N_6091,N_5623,N_5756);
nand U6092 (N_6092,N_5751,N_5543);
nor U6093 (N_6093,N_5979,N_5744);
or U6094 (N_6094,N_5697,N_5943);
xor U6095 (N_6095,N_5926,N_5722);
nand U6096 (N_6096,N_5923,N_5743);
nand U6097 (N_6097,N_5507,N_5512);
and U6098 (N_6098,N_5955,N_5510);
nor U6099 (N_6099,N_5786,N_5609);
nand U6100 (N_6100,N_5848,N_5912);
nor U6101 (N_6101,N_5687,N_5811);
and U6102 (N_6102,N_5535,N_5648);
nor U6103 (N_6103,N_5951,N_5656);
nand U6104 (N_6104,N_5619,N_5812);
or U6105 (N_6105,N_5949,N_5598);
or U6106 (N_6106,N_5521,N_5564);
nand U6107 (N_6107,N_5504,N_5956);
xor U6108 (N_6108,N_5714,N_5766);
xor U6109 (N_6109,N_5874,N_5892);
nand U6110 (N_6110,N_5653,N_5906);
nand U6111 (N_6111,N_5536,N_5569);
xor U6112 (N_6112,N_5937,N_5658);
and U6113 (N_6113,N_5957,N_5893);
nand U6114 (N_6114,N_5996,N_5655);
or U6115 (N_6115,N_5539,N_5855);
nor U6116 (N_6116,N_5705,N_5991);
nand U6117 (N_6117,N_5551,N_5758);
and U6118 (N_6118,N_5915,N_5804);
nor U6119 (N_6119,N_5867,N_5896);
nor U6120 (N_6120,N_5968,N_5973);
xor U6121 (N_6121,N_5690,N_5567);
or U6122 (N_6122,N_5922,N_5560);
or U6123 (N_6123,N_5829,N_5950);
or U6124 (N_6124,N_5635,N_5630);
or U6125 (N_6125,N_5724,N_5554);
or U6126 (N_6126,N_5558,N_5767);
nor U6127 (N_6127,N_5538,N_5607);
nand U6128 (N_6128,N_5644,N_5878);
and U6129 (N_6129,N_5838,N_5908);
or U6130 (N_6130,N_5870,N_5612);
nand U6131 (N_6131,N_5671,N_5982);
xor U6132 (N_6132,N_5847,N_5972);
or U6133 (N_6133,N_5597,N_5501);
or U6134 (N_6134,N_5820,N_5967);
and U6135 (N_6135,N_5517,N_5593);
nor U6136 (N_6136,N_5601,N_5782);
nor U6137 (N_6137,N_5669,N_5916);
nor U6138 (N_6138,N_5754,N_5707);
and U6139 (N_6139,N_5557,N_5613);
nor U6140 (N_6140,N_5875,N_5596);
nor U6141 (N_6141,N_5944,N_5990);
or U6142 (N_6142,N_5800,N_5986);
and U6143 (N_6143,N_5514,N_5672);
or U6144 (N_6144,N_5830,N_5993);
nand U6145 (N_6145,N_5506,N_5776);
and U6146 (N_6146,N_5945,N_5868);
or U6147 (N_6147,N_5994,N_5859);
nand U6148 (N_6148,N_5586,N_5755);
nor U6149 (N_6149,N_5745,N_5742);
nand U6150 (N_6150,N_5686,N_5939);
xor U6151 (N_6151,N_5809,N_5854);
nor U6152 (N_6152,N_5789,N_5641);
nand U6153 (N_6153,N_5866,N_5710);
xor U6154 (N_6154,N_5577,N_5778);
and U6155 (N_6155,N_5828,N_5519);
and U6156 (N_6156,N_5865,N_5941);
nor U6157 (N_6157,N_5516,N_5933);
xnor U6158 (N_6158,N_5790,N_5578);
nand U6159 (N_6159,N_5966,N_5582);
nand U6160 (N_6160,N_5555,N_5683);
and U6161 (N_6161,N_5541,N_5934);
nand U6162 (N_6162,N_5620,N_5935);
or U6163 (N_6163,N_5898,N_5827);
nor U6164 (N_6164,N_5529,N_5762);
nor U6165 (N_6165,N_5676,N_5546);
and U6166 (N_6166,N_5715,N_5962);
or U6167 (N_6167,N_5798,N_5625);
xnor U6168 (N_6168,N_5542,N_5525);
nor U6169 (N_6169,N_5605,N_5584);
and U6170 (N_6170,N_5606,N_5548);
and U6171 (N_6171,N_5547,N_5753);
or U6172 (N_6172,N_5763,N_5540);
and U6173 (N_6173,N_5719,N_5726);
nor U6174 (N_6174,N_5650,N_5663);
xor U6175 (N_6175,N_5921,N_5984);
or U6176 (N_6176,N_5741,N_5694);
and U6177 (N_6177,N_5752,N_5544);
and U6178 (N_6178,N_5872,N_5639);
nand U6179 (N_6179,N_5592,N_5723);
and U6180 (N_6180,N_5773,N_5832);
nor U6181 (N_6181,N_5988,N_5677);
xor U6182 (N_6182,N_5769,N_5783);
nand U6183 (N_6183,N_5792,N_5764);
and U6184 (N_6184,N_5509,N_5587);
and U6185 (N_6185,N_5716,N_5958);
nor U6186 (N_6186,N_5708,N_5649);
nor U6187 (N_6187,N_5703,N_5969);
nand U6188 (N_6188,N_5603,N_5695);
nor U6189 (N_6189,N_5528,N_5806);
or U6190 (N_6190,N_5621,N_5861);
xor U6191 (N_6191,N_5817,N_5631);
nand U6192 (N_6192,N_5588,N_5696);
xnor U6193 (N_6193,N_5706,N_5661);
or U6194 (N_6194,N_5531,N_5905);
or U6195 (N_6195,N_5853,N_5590);
nand U6196 (N_6196,N_5585,N_5818);
xnor U6197 (N_6197,N_5666,N_5774);
or U6198 (N_6198,N_5522,N_5887);
nand U6199 (N_6199,N_5680,N_5576);
or U6200 (N_6200,N_5765,N_5615);
nand U6201 (N_6201,N_5929,N_5917);
xor U6202 (N_6202,N_5532,N_5699);
and U6203 (N_6203,N_5947,N_5837);
and U6204 (N_6204,N_5693,N_5685);
or U6205 (N_6205,N_5513,N_5821);
nor U6206 (N_6206,N_5660,N_5736);
xnor U6207 (N_6207,N_5948,N_5924);
nor U6208 (N_6208,N_5574,N_5730);
xor U6209 (N_6209,N_5961,N_5647);
xnor U6210 (N_6210,N_5824,N_5801);
nor U6211 (N_6211,N_5735,N_5759);
and U6212 (N_6212,N_5563,N_5550);
and U6213 (N_6213,N_5900,N_5575);
or U6214 (N_6214,N_5684,N_5960);
xnor U6215 (N_6215,N_5813,N_5954);
nor U6216 (N_6216,N_5505,N_5927);
nand U6217 (N_6217,N_5932,N_5571);
xor U6218 (N_6218,N_5637,N_5718);
nor U6219 (N_6219,N_5771,N_5884);
nand U6220 (N_6220,N_5616,N_5670);
nand U6221 (N_6221,N_5537,N_5732);
nor U6222 (N_6222,N_5831,N_5652);
nor U6223 (N_6223,N_5797,N_5899);
xor U6224 (N_6224,N_5657,N_5795);
nor U6225 (N_6225,N_5931,N_5987);
nor U6226 (N_6226,N_5727,N_5643);
or U6227 (N_6227,N_5614,N_5976);
and U6228 (N_6228,N_5768,N_5633);
nor U6229 (N_6229,N_5913,N_5998);
and U6230 (N_6230,N_5970,N_5895);
xor U6231 (N_6231,N_5556,N_5739);
xnor U6232 (N_6232,N_5570,N_5659);
xor U6233 (N_6233,N_5645,N_5508);
xor U6234 (N_6234,N_5845,N_5844);
nor U6235 (N_6235,N_5682,N_5568);
nor U6236 (N_6236,N_5971,N_5622);
nor U6237 (N_6237,N_5561,N_5713);
xor U6238 (N_6238,N_5566,N_5825);
nor U6239 (N_6239,N_5524,N_5938);
nand U6240 (N_6240,N_5746,N_5737);
nor U6241 (N_6241,N_5852,N_5810);
nor U6242 (N_6242,N_5589,N_5523);
or U6243 (N_6243,N_5667,N_5959);
nor U6244 (N_6244,N_5733,N_5863);
nor U6245 (N_6245,N_5734,N_5634);
nor U6246 (N_6246,N_5918,N_5891);
or U6247 (N_6247,N_5851,N_5740);
and U6248 (N_6248,N_5591,N_5992);
xnor U6249 (N_6249,N_5679,N_5668);
nand U6250 (N_6250,N_5750,N_5628);
nand U6251 (N_6251,N_5863,N_5903);
or U6252 (N_6252,N_5918,N_5869);
xnor U6253 (N_6253,N_5751,N_5570);
nand U6254 (N_6254,N_5620,N_5833);
and U6255 (N_6255,N_5763,N_5621);
or U6256 (N_6256,N_5790,N_5584);
xor U6257 (N_6257,N_5682,N_5720);
and U6258 (N_6258,N_5665,N_5645);
xor U6259 (N_6259,N_5662,N_5759);
or U6260 (N_6260,N_5989,N_5567);
xnor U6261 (N_6261,N_5979,N_5631);
xor U6262 (N_6262,N_5829,N_5874);
xnor U6263 (N_6263,N_5833,N_5999);
or U6264 (N_6264,N_5769,N_5744);
and U6265 (N_6265,N_5960,N_5543);
or U6266 (N_6266,N_5538,N_5823);
and U6267 (N_6267,N_5743,N_5901);
nor U6268 (N_6268,N_5773,N_5533);
nand U6269 (N_6269,N_5654,N_5811);
nand U6270 (N_6270,N_5950,N_5803);
nand U6271 (N_6271,N_5564,N_5640);
nor U6272 (N_6272,N_5736,N_5631);
or U6273 (N_6273,N_5931,N_5519);
nand U6274 (N_6274,N_5662,N_5973);
or U6275 (N_6275,N_5833,N_5832);
or U6276 (N_6276,N_5579,N_5653);
nor U6277 (N_6277,N_5742,N_5920);
and U6278 (N_6278,N_5636,N_5823);
nor U6279 (N_6279,N_5574,N_5644);
and U6280 (N_6280,N_5799,N_5926);
xnor U6281 (N_6281,N_5943,N_5894);
and U6282 (N_6282,N_5802,N_5506);
nor U6283 (N_6283,N_5714,N_5515);
nor U6284 (N_6284,N_5929,N_5620);
and U6285 (N_6285,N_5723,N_5985);
or U6286 (N_6286,N_5512,N_5776);
nand U6287 (N_6287,N_5706,N_5861);
nor U6288 (N_6288,N_5643,N_5607);
xor U6289 (N_6289,N_5569,N_5578);
and U6290 (N_6290,N_5927,N_5715);
nor U6291 (N_6291,N_5744,N_5703);
xnor U6292 (N_6292,N_5709,N_5980);
nand U6293 (N_6293,N_5604,N_5600);
xor U6294 (N_6294,N_5856,N_5949);
nor U6295 (N_6295,N_5992,N_5687);
xor U6296 (N_6296,N_5541,N_5574);
nor U6297 (N_6297,N_5751,N_5866);
nor U6298 (N_6298,N_5551,N_5824);
xor U6299 (N_6299,N_5581,N_5767);
or U6300 (N_6300,N_5822,N_5851);
nor U6301 (N_6301,N_5565,N_5559);
nand U6302 (N_6302,N_5698,N_5935);
nand U6303 (N_6303,N_5949,N_5813);
nand U6304 (N_6304,N_5969,N_5934);
and U6305 (N_6305,N_5770,N_5671);
nand U6306 (N_6306,N_5974,N_5827);
or U6307 (N_6307,N_5627,N_5800);
nor U6308 (N_6308,N_5657,N_5978);
and U6309 (N_6309,N_5802,N_5838);
nor U6310 (N_6310,N_5992,N_5786);
and U6311 (N_6311,N_5650,N_5932);
or U6312 (N_6312,N_5736,N_5873);
nand U6313 (N_6313,N_5672,N_5638);
xnor U6314 (N_6314,N_5697,N_5609);
nor U6315 (N_6315,N_5806,N_5804);
xor U6316 (N_6316,N_5687,N_5530);
nand U6317 (N_6317,N_5542,N_5806);
and U6318 (N_6318,N_5602,N_5979);
nor U6319 (N_6319,N_5739,N_5746);
and U6320 (N_6320,N_5836,N_5548);
and U6321 (N_6321,N_5531,N_5770);
xor U6322 (N_6322,N_5521,N_5813);
nand U6323 (N_6323,N_5608,N_5914);
nand U6324 (N_6324,N_5883,N_5828);
nand U6325 (N_6325,N_5664,N_5521);
nand U6326 (N_6326,N_5756,N_5649);
or U6327 (N_6327,N_5856,N_5888);
nor U6328 (N_6328,N_5846,N_5849);
and U6329 (N_6329,N_5784,N_5785);
nor U6330 (N_6330,N_5933,N_5595);
nand U6331 (N_6331,N_5644,N_5758);
nor U6332 (N_6332,N_5973,N_5946);
and U6333 (N_6333,N_5954,N_5549);
xnor U6334 (N_6334,N_5581,N_5720);
xnor U6335 (N_6335,N_5506,N_5644);
and U6336 (N_6336,N_5947,N_5765);
nor U6337 (N_6337,N_5911,N_5906);
nand U6338 (N_6338,N_5519,N_5663);
xor U6339 (N_6339,N_5843,N_5517);
nand U6340 (N_6340,N_5906,N_5835);
xnor U6341 (N_6341,N_5869,N_5524);
nor U6342 (N_6342,N_5930,N_5604);
nand U6343 (N_6343,N_5916,N_5527);
or U6344 (N_6344,N_5764,N_5896);
or U6345 (N_6345,N_5702,N_5995);
nand U6346 (N_6346,N_5987,N_5594);
xor U6347 (N_6347,N_5901,N_5871);
or U6348 (N_6348,N_5597,N_5969);
nand U6349 (N_6349,N_5619,N_5976);
or U6350 (N_6350,N_5972,N_5805);
xnor U6351 (N_6351,N_5858,N_5735);
nor U6352 (N_6352,N_5603,N_5514);
xor U6353 (N_6353,N_5592,N_5707);
or U6354 (N_6354,N_5918,N_5705);
nor U6355 (N_6355,N_5800,N_5994);
nand U6356 (N_6356,N_5955,N_5520);
nor U6357 (N_6357,N_5715,N_5567);
nor U6358 (N_6358,N_5990,N_5680);
nand U6359 (N_6359,N_5954,N_5823);
nand U6360 (N_6360,N_5765,N_5549);
and U6361 (N_6361,N_5553,N_5544);
xnor U6362 (N_6362,N_5805,N_5727);
and U6363 (N_6363,N_5978,N_5999);
or U6364 (N_6364,N_5889,N_5931);
nand U6365 (N_6365,N_5535,N_5599);
nand U6366 (N_6366,N_5945,N_5646);
xor U6367 (N_6367,N_5876,N_5757);
nor U6368 (N_6368,N_5569,N_5942);
xor U6369 (N_6369,N_5831,N_5524);
or U6370 (N_6370,N_5679,N_5828);
nand U6371 (N_6371,N_5658,N_5727);
xnor U6372 (N_6372,N_5805,N_5807);
xnor U6373 (N_6373,N_5814,N_5829);
nor U6374 (N_6374,N_5613,N_5998);
or U6375 (N_6375,N_5633,N_5884);
nor U6376 (N_6376,N_5718,N_5589);
xor U6377 (N_6377,N_5943,N_5547);
xnor U6378 (N_6378,N_5784,N_5865);
or U6379 (N_6379,N_5500,N_5880);
nor U6380 (N_6380,N_5796,N_5841);
nor U6381 (N_6381,N_5833,N_5877);
nand U6382 (N_6382,N_5880,N_5796);
and U6383 (N_6383,N_5896,N_5682);
nor U6384 (N_6384,N_5629,N_5964);
xnor U6385 (N_6385,N_5520,N_5855);
nor U6386 (N_6386,N_5684,N_5845);
and U6387 (N_6387,N_5906,N_5713);
and U6388 (N_6388,N_5597,N_5792);
or U6389 (N_6389,N_5525,N_5776);
and U6390 (N_6390,N_5514,N_5870);
nand U6391 (N_6391,N_5510,N_5834);
xnor U6392 (N_6392,N_5955,N_5954);
nor U6393 (N_6393,N_5660,N_5972);
or U6394 (N_6394,N_5703,N_5913);
and U6395 (N_6395,N_5828,N_5649);
nor U6396 (N_6396,N_5939,N_5617);
nand U6397 (N_6397,N_5735,N_5664);
nand U6398 (N_6398,N_5957,N_5647);
nand U6399 (N_6399,N_5559,N_5940);
nor U6400 (N_6400,N_5720,N_5570);
or U6401 (N_6401,N_5631,N_5625);
and U6402 (N_6402,N_5809,N_5871);
or U6403 (N_6403,N_5687,N_5780);
xnor U6404 (N_6404,N_5500,N_5698);
xor U6405 (N_6405,N_5824,N_5960);
and U6406 (N_6406,N_5686,N_5609);
nand U6407 (N_6407,N_5820,N_5543);
xor U6408 (N_6408,N_5983,N_5635);
nor U6409 (N_6409,N_5771,N_5500);
nand U6410 (N_6410,N_5644,N_5705);
or U6411 (N_6411,N_5950,N_5750);
xor U6412 (N_6412,N_5518,N_5915);
nor U6413 (N_6413,N_5730,N_5868);
nor U6414 (N_6414,N_5589,N_5532);
nor U6415 (N_6415,N_5831,N_5856);
nand U6416 (N_6416,N_5686,N_5738);
or U6417 (N_6417,N_5561,N_5615);
or U6418 (N_6418,N_5836,N_5713);
or U6419 (N_6419,N_5843,N_5722);
xor U6420 (N_6420,N_5842,N_5508);
and U6421 (N_6421,N_5550,N_5541);
and U6422 (N_6422,N_5976,N_5853);
xor U6423 (N_6423,N_5547,N_5565);
xnor U6424 (N_6424,N_5884,N_5915);
and U6425 (N_6425,N_5712,N_5693);
or U6426 (N_6426,N_5501,N_5552);
and U6427 (N_6427,N_5613,N_5869);
or U6428 (N_6428,N_5967,N_5762);
and U6429 (N_6429,N_5558,N_5863);
nor U6430 (N_6430,N_5530,N_5893);
or U6431 (N_6431,N_5632,N_5709);
xor U6432 (N_6432,N_5597,N_5562);
nor U6433 (N_6433,N_5691,N_5612);
nor U6434 (N_6434,N_5883,N_5776);
and U6435 (N_6435,N_5553,N_5745);
nand U6436 (N_6436,N_5993,N_5729);
and U6437 (N_6437,N_5603,N_5912);
or U6438 (N_6438,N_5639,N_5549);
or U6439 (N_6439,N_5740,N_5633);
nand U6440 (N_6440,N_5798,N_5908);
nand U6441 (N_6441,N_5991,N_5633);
or U6442 (N_6442,N_5830,N_5617);
or U6443 (N_6443,N_5610,N_5913);
or U6444 (N_6444,N_5809,N_5811);
and U6445 (N_6445,N_5914,N_5662);
or U6446 (N_6446,N_5871,N_5701);
nor U6447 (N_6447,N_5934,N_5739);
or U6448 (N_6448,N_5666,N_5828);
xor U6449 (N_6449,N_5773,N_5821);
nand U6450 (N_6450,N_5694,N_5969);
xor U6451 (N_6451,N_5619,N_5943);
nand U6452 (N_6452,N_5950,N_5500);
and U6453 (N_6453,N_5644,N_5680);
xor U6454 (N_6454,N_5642,N_5989);
nor U6455 (N_6455,N_5699,N_5531);
or U6456 (N_6456,N_5660,N_5982);
nand U6457 (N_6457,N_5646,N_5754);
nand U6458 (N_6458,N_5962,N_5794);
and U6459 (N_6459,N_5826,N_5804);
nor U6460 (N_6460,N_5897,N_5608);
nor U6461 (N_6461,N_5793,N_5515);
xnor U6462 (N_6462,N_5729,N_5977);
nand U6463 (N_6463,N_5951,N_5658);
and U6464 (N_6464,N_5956,N_5678);
xnor U6465 (N_6465,N_5874,N_5628);
and U6466 (N_6466,N_5991,N_5935);
xor U6467 (N_6467,N_5976,N_5903);
xor U6468 (N_6468,N_5859,N_5951);
or U6469 (N_6469,N_5694,N_5717);
xor U6470 (N_6470,N_5518,N_5927);
or U6471 (N_6471,N_5666,N_5517);
nor U6472 (N_6472,N_5576,N_5552);
and U6473 (N_6473,N_5915,N_5972);
xnor U6474 (N_6474,N_5555,N_5547);
xnor U6475 (N_6475,N_5945,N_5501);
or U6476 (N_6476,N_5893,N_5622);
nor U6477 (N_6477,N_5878,N_5951);
or U6478 (N_6478,N_5998,N_5568);
nor U6479 (N_6479,N_5946,N_5563);
or U6480 (N_6480,N_5672,N_5743);
or U6481 (N_6481,N_5832,N_5980);
and U6482 (N_6482,N_5917,N_5502);
xor U6483 (N_6483,N_5539,N_5881);
nor U6484 (N_6484,N_5786,N_5854);
xnor U6485 (N_6485,N_5522,N_5686);
nor U6486 (N_6486,N_5668,N_5757);
xor U6487 (N_6487,N_5641,N_5661);
nand U6488 (N_6488,N_5797,N_5694);
xor U6489 (N_6489,N_5882,N_5849);
nor U6490 (N_6490,N_5751,N_5554);
xnor U6491 (N_6491,N_5815,N_5718);
nor U6492 (N_6492,N_5585,N_5761);
nor U6493 (N_6493,N_5815,N_5530);
and U6494 (N_6494,N_5956,N_5805);
or U6495 (N_6495,N_5823,N_5510);
xnor U6496 (N_6496,N_5691,N_5710);
or U6497 (N_6497,N_5665,N_5512);
xnor U6498 (N_6498,N_5969,N_5508);
and U6499 (N_6499,N_5634,N_5867);
nor U6500 (N_6500,N_6216,N_6453);
nor U6501 (N_6501,N_6377,N_6008);
or U6502 (N_6502,N_6183,N_6392);
nor U6503 (N_6503,N_6026,N_6155);
nor U6504 (N_6504,N_6204,N_6047);
nor U6505 (N_6505,N_6298,N_6258);
nand U6506 (N_6506,N_6198,N_6031);
or U6507 (N_6507,N_6361,N_6219);
xor U6508 (N_6508,N_6161,N_6498);
nand U6509 (N_6509,N_6094,N_6412);
xnor U6510 (N_6510,N_6193,N_6404);
or U6511 (N_6511,N_6433,N_6281);
nor U6512 (N_6512,N_6253,N_6358);
xnor U6513 (N_6513,N_6291,N_6028);
or U6514 (N_6514,N_6066,N_6046);
xor U6515 (N_6515,N_6274,N_6076);
xnor U6516 (N_6516,N_6445,N_6259);
xor U6517 (N_6517,N_6370,N_6299);
or U6518 (N_6518,N_6472,N_6150);
or U6519 (N_6519,N_6061,N_6084);
and U6520 (N_6520,N_6049,N_6043);
xor U6521 (N_6521,N_6068,N_6019);
or U6522 (N_6522,N_6473,N_6201);
nand U6523 (N_6523,N_6380,N_6101);
xnor U6524 (N_6524,N_6439,N_6456);
and U6525 (N_6525,N_6207,N_6120);
and U6526 (N_6526,N_6181,N_6236);
nand U6527 (N_6527,N_6329,N_6295);
and U6528 (N_6528,N_6128,N_6231);
or U6529 (N_6529,N_6360,N_6293);
xnor U6530 (N_6530,N_6347,N_6420);
nand U6531 (N_6531,N_6427,N_6438);
and U6532 (N_6532,N_6162,N_6121);
nand U6533 (N_6533,N_6434,N_6264);
xor U6534 (N_6534,N_6273,N_6232);
or U6535 (N_6535,N_6288,N_6414);
nand U6536 (N_6536,N_6167,N_6174);
nor U6537 (N_6537,N_6312,N_6118);
or U6538 (N_6538,N_6202,N_6369);
or U6539 (N_6539,N_6304,N_6218);
nand U6540 (N_6540,N_6185,N_6323);
nand U6541 (N_6541,N_6071,N_6085);
nor U6542 (N_6542,N_6494,N_6217);
nand U6543 (N_6543,N_6206,N_6317);
nand U6544 (N_6544,N_6469,N_6172);
nor U6545 (N_6545,N_6177,N_6459);
xnor U6546 (N_6546,N_6126,N_6109);
nor U6547 (N_6547,N_6470,N_6330);
nor U6548 (N_6548,N_6062,N_6239);
and U6549 (N_6549,N_6243,N_6034);
nor U6550 (N_6550,N_6014,N_6444);
or U6551 (N_6551,N_6276,N_6322);
nand U6552 (N_6552,N_6309,N_6376);
xnor U6553 (N_6553,N_6333,N_6362);
xnor U6554 (N_6554,N_6192,N_6441);
xor U6555 (N_6555,N_6462,N_6223);
nand U6556 (N_6556,N_6214,N_6331);
xor U6557 (N_6557,N_6210,N_6484);
nor U6558 (N_6558,N_6039,N_6159);
nor U6559 (N_6559,N_6311,N_6203);
and U6560 (N_6560,N_6345,N_6373);
nor U6561 (N_6561,N_6107,N_6448);
nand U6562 (N_6562,N_6129,N_6242);
nand U6563 (N_6563,N_6344,N_6176);
nand U6564 (N_6564,N_6215,N_6411);
and U6565 (N_6565,N_6478,N_6179);
nor U6566 (N_6566,N_6266,N_6467);
nor U6567 (N_6567,N_6270,N_6247);
or U6568 (N_6568,N_6496,N_6033);
and U6569 (N_6569,N_6263,N_6447);
xnor U6570 (N_6570,N_6166,N_6222);
xnor U6571 (N_6571,N_6148,N_6386);
xnor U6572 (N_6572,N_6132,N_6211);
nand U6573 (N_6573,N_6135,N_6170);
and U6574 (N_6574,N_6136,N_6142);
nand U6575 (N_6575,N_6108,N_6488);
and U6576 (N_6576,N_6029,N_6446);
and U6577 (N_6577,N_6290,N_6237);
xnor U6578 (N_6578,N_6173,N_6391);
or U6579 (N_6579,N_6381,N_6067);
nor U6580 (N_6580,N_6036,N_6228);
nand U6581 (N_6581,N_6030,N_6226);
xnor U6582 (N_6582,N_6460,N_6105);
nand U6583 (N_6583,N_6093,N_6353);
xor U6584 (N_6584,N_6012,N_6015);
and U6585 (N_6585,N_6285,N_6475);
or U6586 (N_6586,N_6042,N_6278);
xor U6587 (N_6587,N_6005,N_6275);
nand U6588 (N_6588,N_6490,N_6079);
nand U6589 (N_6589,N_6319,N_6156);
or U6590 (N_6590,N_6497,N_6397);
xor U6591 (N_6591,N_6096,N_6091);
nand U6592 (N_6592,N_6104,N_6078);
nor U6593 (N_6593,N_6131,N_6262);
xor U6594 (N_6594,N_6356,N_6251);
nand U6595 (N_6595,N_6082,N_6349);
and U6596 (N_6596,N_6286,N_6165);
or U6597 (N_6597,N_6209,N_6001);
nor U6598 (N_6598,N_6018,N_6440);
or U6599 (N_6599,N_6431,N_6424);
and U6600 (N_6600,N_6272,N_6044);
and U6601 (N_6601,N_6495,N_6442);
or U6602 (N_6602,N_6374,N_6325);
xor U6603 (N_6603,N_6038,N_6340);
or U6604 (N_6604,N_6149,N_6250);
or U6605 (N_6605,N_6419,N_6194);
xnor U6606 (N_6606,N_6205,N_6220);
and U6607 (N_6607,N_6188,N_6389);
and U6608 (N_6608,N_6316,N_6306);
nand U6609 (N_6609,N_6402,N_6393);
and U6610 (N_6610,N_6308,N_6310);
nor U6611 (N_6611,N_6010,N_6056);
nor U6612 (N_6612,N_6388,N_6385);
xor U6613 (N_6613,N_6463,N_6020);
and U6614 (N_6614,N_6267,N_6009);
and U6615 (N_6615,N_6007,N_6055);
and U6616 (N_6616,N_6423,N_6081);
or U6617 (N_6617,N_6413,N_6489);
xor U6618 (N_6618,N_6022,N_6338);
and U6619 (N_6619,N_6134,N_6261);
nand U6620 (N_6620,N_6169,N_6013);
and U6621 (N_6621,N_6147,N_6021);
and U6622 (N_6622,N_6408,N_6224);
xor U6623 (N_6623,N_6437,N_6059);
nand U6624 (N_6624,N_6378,N_6313);
nor U6625 (N_6625,N_6212,N_6152);
nand U6626 (N_6626,N_6100,N_6390);
nand U6627 (N_6627,N_6363,N_6271);
xor U6628 (N_6628,N_6297,N_6401);
nand U6629 (N_6629,N_6037,N_6372);
or U6630 (N_6630,N_6359,N_6301);
nand U6631 (N_6631,N_6127,N_6364);
and U6632 (N_6632,N_6016,N_6436);
nor U6633 (N_6633,N_6384,N_6058);
xor U6634 (N_6634,N_6171,N_6403);
nand U6635 (N_6635,N_6337,N_6450);
or U6636 (N_6636,N_6332,N_6075);
nand U6637 (N_6637,N_6035,N_6163);
or U6638 (N_6638,N_6083,N_6065);
xor U6639 (N_6639,N_6006,N_6480);
xnor U6640 (N_6640,N_6289,N_6334);
xor U6641 (N_6641,N_6328,N_6409);
nand U6642 (N_6642,N_6112,N_6294);
nand U6643 (N_6643,N_6417,N_6416);
nand U6644 (N_6644,N_6151,N_6095);
nor U6645 (N_6645,N_6199,N_6140);
nand U6646 (N_6646,N_6421,N_6057);
nor U6647 (N_6647,N_6023,N_6144);
nand U6648 (N_6648,N_6032,N_6352);
or U6649 (N_6649,N_6160,N_6196);
or U6650 (N_6650,N_6394,N_6367);
nor U6651 (N_6651,N_6341,N_6111);
and U6652 (N_6652,N_6244,N_6249);
nor U6653 (N_6653,N_6117,N_6195);
and U6654 (N_6654,N_6158,N_6164);
nor U6655 (N_6655,N_6189,N_6123);
nand U6656 (N_6656,N_6277,N_6230);
nand U6657 (N_6657,N_6466,N_6197);
and U6658 (N_6658,N_6415,N_6398);
or U6659 (N_6659,N_6077,N_6099);
and U6660 (N_6660,N_6284,N_6483);
xnor U6661 (N_6661,N_6110,N_6041);
or U6662 (N_6662,N_6305,N_6454);
and U6663 (N_6663,N_6400,N_6063);
nor U6664 (N_6664,N_6143,N_6474);
nor U6665 (N_6665,N_6300,N_6452);
nor U6666 (N_6666,N_6137,N_6269);
xnor U6667 (N_6667,N_6184,N_6418);
nor U6668 (N_6668,N_6233,N_6190);
nor U6669 (N_6669,N_6410,N_6115);
xnor U6670 (N_6670,N_6139,N_6200);
nor U6671 (N_6671,N_6339,N_6303);
xor U6672 (N_6672,N_6479,N_6060);
and U6673 (N_6673,N_6324,N_6141);
or U6674 (N_6674,N_6106,N_6265);
and U6675 (N_6675,N_6113,N_6375);
nor U6676 (N_6676,N_6070,N_6307);
and U6677 (N_6677,N_6255,N_6365);
or U6678 (N_6678,N_6103,N_6428);
nand U6679 (N_6679,N_6153,N_6241);
nor U6680 (N_6680,N_6130,N_6292);
nor U6681 (N_6681,N_6318,N_6133);
or U6682 (N_6682,N_6432,N_6011);
nand U6683 (N_6683,N_6114,N_6355);
or U6684 (N_6684,N_6074,N_6154);
and U6685 (N_6685,N_6025,N_6254);
or U6686 (N_6686,N_6396,N_6122);
nand U6687 (N_6687,N_6186,N_6168);
xor U6688 (N_6688,N_6451,N_6429);
and U6689 (N_6689,N_6296,N_6368);
and U6690 (N_6690,N_6465,N_6335);
and U6691 (N_6691,N_6138,N_6221);
nand U6692 (N_6692,N_6208,N_6157);
xor U6693 (N_6693,N_6405,N_6321);
nand U6694 (N_6694,N_6268,N_6482);
and U6695 (N_6695,N_6407,N_6464);
nor U6696 (N_6696,N_6248,N_6072);
xor U6697 (N_6697,N_6491,N_6125);
or U6698 (N_6698,N_6383,N_6346);
or U6699 (N_6699,N_6320,N_6234);
nand U6700 (N_6700,N_6098,N_6054);
and U6701 (N_6701,N_6090,N_6257);
nor U6702 (N_6702,N_6040,N_6000);
and U6703 (N_6703,N_6229,N_6245);
and U6704 (N_6704,N_6048,N_6282);
or U6705 (N_6705,N_6252,N_6145);
xor U6706 (N_6706,N_6348,N_6422);
nor U6707 (N_6707,N_6314,N_6182);
nor U6708 (N_6708,N_6260,N_6086);
nor U6709 (N_6709,N_6382,N_6050);
xnor U6710 (N_6710,N_6302,N_6351);
nand U6711 (N_6711,N_6477,N_6343);
nor U6712 (N_6712,N_6366,N_6283);
nand U6713 (N_6713,N_6092,N_6024);
nand U6714 (N_6714,N_6327,N_6175);
xor U6715 (N_6715,N_6004,N_6235);
or U6716 (N_6716,N_6492,N_6461);
nand U6717 (N_6717,N_6088,N_6213);
and U6718 (N_6718,N_6455,N_6045);
xnor U6719 (N_6719,N_6449,N_6256);
nor U6720 (N_6720,N_6187,N_6425);
nand U6721 (N_6721,N_6426,N_6087);
xnor U6722 (N_6722,N_6357,N_6240);
xnor U6723 (N_6723,N_6493,N_6180);
nor U6724 (N_6724,N_6485,N_6146);
xor U6725 (N_6725,N_6315,N_6051);
xnor U6726 (N_6726,N_6430,N_6102);
nor U6727 (N_6727,N_6080,N_6487);
xnor U6728 (N_6728,N_6471,N_6342);
and U6729 (N_6729,N_6435,N_6279);
nand U6730 (N_6730,N_6124,N_6178);
nor U6731 (N_6731,N_6069,N_6371);
and U6732 (N_6732,N_6073,N_6468);
or U6733 (N_6733,N_6395,N_6287);
or U6734 (N_6734,N_6191,N_6053);
xnor U6735 (N_6735,N_6486,N_6457);
nor U6736 (N_6736,N_6336,N_6027);
nor U6737 (N_6737,N_6064,N_6017);
xor U6738 (N_6738,N_6379,N_6116);
or U6739 (N_6739,N_6119,N_6354);
or U6740 (N_6740,N_6458,N_6225);
nor U6741 (N_6741,N_6326,N_6499);
nand U6742 (N_6742,N_6399,N_6097);
nand U6743 (N_6743,N_6003,N_6052);
or U6744 (N_6744,N_6089,N_6246);
and U6745 (N_6745,N_6406,N_6280);
xor U6746 (N_6746,N_6481,N_6387);
nand U6747 (N_6747,N_6238,N_6476);
nor U6748 (N_6748,N_6227,N_6443);
nor U6749 (N_6749,N_6002,N_6350);
and U6750 (N_6750,N_6208,N_6266);
or U6751 (N_6751,N_6413,N_6456);
nand U6752 (N_6752,N_6333,N_6317);
nor U6753 (N_6753,N_6074,N_6150);
xnor U6754 (N_6754,N_6251,N_6037);
nand U6755 (N_6755,N_6032,N_6280);
xnor U6756 (N_6756,N_6015,N_6082);
or U6757 (N_6757,N_6449,N_6104);
and U6758 (N_6758,N_6124,N_6371);
xnor U6759 (N_6759,N_6223,N_6225);
xor U6760 (N_6760,N_6186,N_6444);
xnor U6761 (N_6761,N_6363,N_6139);
and U6762 (N_6762,N_6477,N_6132);
nand U6763 (N_6763,N_6448,N_6456);
nand U6764 (N_6764,N_6422,N_6016);
nand U6765 (N_6765,N_6429,N_6124);
or U6766 (N_6766,N_6439,N_6269);
nor U6767 (N_6767,N_6226,N_6422);
nor U6768 (N_6768,N_6402,N_6083);
and U6769 (N_6769,N_6216,N_6008);
or U6770 (N_6770,N_6352,N_6266);
nor U6771 (N_6771,N_6494,N_6157);
xnor U6772 (N_6772,N_6028,N_6484);
nand U6773 (N_6773,N_6044,N_6054);
nor U6774 (N_6774,N_6139,N_6441);
and U6775 (N_6775,N_6454,N_6066);
xnor U6776 (N_6776,N_6462,N_6371);
and U6777 (N_6777,N_6214,N_6281);
and U6778 (N_6778,N_6339,N_6106);
or U6779 (N_6779,N_6281,N_6089);
nor U6780 (N_6780,N_6050,N_6087);
or U6781 (N_6781,N_6496,N_6161);
nor U6782 (N_6782,N_6391,N_6013);
nor U6783 (N_6783,N_6005,N_6470);
and U6784 (N_6784,N_6177,N_6015);
and U6785 (N_6785,N_6151,N_6029);
or U6786 (N_6786,N_6398,N_6237);
or U6787 (N_6787,N_6100,N_6312);
and U6788 (N_6788,N_6324,N_6077);
or U6789 (N_6789,N_6311,N_6288);
xor U6790 (N_6790,N_6055,N_6307);
and U6791 (N_6791,N_6283,N_6046);
nor U6792 (N_6792,N_6145,N_6007);
xor U6793 (N_6793,N_6399,N_6396);
xnor U6794 (N_6794,N_6473,N_6127);
and U6795 (N_6795,N_6172,N_6299);
nor U6796 (N_6796,N_6494,N_6386);
nand U6797 (N_6797,N_6435,N_6040);
nor U6798 (N_6798,N_6119,N_6281);
xnor U6799 (N_6799,N_6456,N_6202);
xor U6800 (N_6800,N_6483,N_6268);
and U6801 (N_6801,N_6258,N_6062);
and U6802 (N_6802,N_6468,N_6081);
nand U6803 (N_6803,N_6354,N_6275);
nand U6804 (N_6804,N_6257,N_6188);
nor U6805 (N_6805,N_6118,N_6493);
nand U6806 (N_6806,N_6114,N_6307);
nand U6807 (N_6807,N_6027,N_6364);
and U6808 (N_6808,N_6451,N_6480);
nor U6809 (N_6809,N_6273,N_6055);
nand U6810 (N_6810,N_6009,N_6334);
nor U6811 (N_6811,N_6172,N_6079);
and U6812 (N_6812,N_6037,N_6114);
or U6813 (N_6813,N_6192,N_6183);
and U6814 (N_6814,N_6210,N_6426);
nand U6815 (N_6815,N_6344,N_6387);
or U6816 (N_6816,N_6136,N_6018);
or U6817 (N_6817,N_6064,N_6259);
nor U6818 (N_6818,N_6312,N_6411);
and U6819 (N_6819,N_6260,N_6223);
or U6820 (N_6820,N_6224,N_6006);
nand U6821 (N_6821,N_6421,N_6114);
nand U6822 (N_6822,N_6200,N_6061);
or U6823 (N_6823,N_6316,N_6491);
nor U6824 (N_6824,N_6292,N_6187);
xnor U6825 (N_6825,N_6388,N_6178);
and U6826 (N_6826,N_6209,N_6401);
and U6827 (N_6827,N_6152,N_6407);
xnor U6828 (N_6828,N_6227,N_6358);
and U6829 (N_6829,N_6085,N_6134);
nor U6830 (N_6830,N_6317,N_6340);
and U6831 (N_6831,N_6214,N_6420);
or U6832 (N_6832,N_6362,N_6170);
or U6833 (N_6833,N_6244,N_6132);
nand U6834 (N_6834,N_6466,N_6408);
nor U6835 (N_6835,N_6063,N_6226);
and U6836 (N_6836,N_6033,N_6088);
and U6837 (N_6837,N_6000,N_6055);
or U6838 (N_6838,N_6161,N_6332);
nor U6839 (N_6839,N_6029,N_6326);
nor U6840 (N_6840,N_6457,N_6083);
xor U6841 (N_6841,N_6182,N_6441);
or U6842 (N_6842,N_6190,N_6386);
or U6843 (N_6843,N_6327,N_6401);
nor U6844 (N_6844,N_6149,N_6067);
nor U6845 (N_6845,N_6405,N_6318);
and U6846 (N_6846,N_6009,N_6410);
and U6847 (N_6847,N_6426,N_6370);
nand U6848 (N_6848,N_6252,N_6163);
and U6849 (N_6849,N_6040,N_6476);
nand U6850 (N_6850,N_6238,N_6433);
nand U6851 (N_6851,N_6401,N_6155);
and U6852 (N_6852,N_6185,N_6437);
nor U6853 (N_6853,N_6272,N_6131);
nand U6854 (N_6854,N_6445,N_6144);
and U6855 (N_6855,N_6025,N_6153);
and U6856 (N_6856,N_6214,N_6126);
xnor U6857 (N_6857,N_6189,N_6384);
nor U6858 (N_6858,N_6331,N_6173);
nand U6859 (N_6859,N_6323,N_6094);
and U6860 (N_6860,N_6479,N_6193);
xnor U6861 (N_6861,N_6025,N_6028);
xor U6862 (N_6862,N_6223,N_6421);
or U6863 (N_6863,N_6161,N_6018);
or U6864 (N_6864,N_6335,N_6054);
nand U6865 (N_6865,N_6291,N_6132);
and U6866 (N_6866,N_6424,N_6328);
and U6867 (N_6867,N_6410,N_6313);
xnor U6868 (N_6868,N_6314,N_6206);
nand U6869 (N_6869,N_6042,N_6239);
nand U6870 (N_6870,N_6374,N_6485);
nand U6871 (N_6871,N_6132,N_6130);
xnor U6872 (N_6872,N_6089,N_6393);
and U6873 (N_6873,N_6488,N_6037);
or U6874 (N_6874,N_6224,N_6360);
or U6875 (N_6875,N_6354,N_6059);
or U6876 (N_6876,N_6015,N_6377);
xnor U6877 (N_6877,N_6380,N_6361);
and U6878 (N_6878,N_6270,N_6491);
nand U6879 (N_6879,N_6279,N_6069);
or U6880 (N_6880,N_6356,N_6346);
nand U6881 (N_6881,N_6038,N_6384);
xnor U6882 (N_6882,N_6027,N_6277);
or U6883 (N_6883,N_6495,N_6323);
nor U6884 (N_6884,N_6028,N_6237);
and U6885 (N_6885,N_6113,N_6023);
or U6886 (N_6886,N_6411,N_6428);
nand U6887 (N_6887,N_6453,N_6458);
or U6888 (N_6888,N_6137,N_6151);
and U6889 (N_6889,N_6399,N_6045);
and U6890 (N_6890,N_6380,N_6366);
and U6891 (N_6891,N_6263,N_6343);
nand U6892 (N_6892,N_6492,N_6468);
nand U6893 (N_6893,N_6290,N_6078);
nor U6894 (N_6894,N_6221,N_6098);
or U6895 (N_6895,N_6113,N_6318);
xor U6896 (N_6896,N_6496,N_6173);
or U6897 (N_6897,N_6224,N_6387);
nand U6898 (N_6898,N_6245,N_6026);
and U6899 (N_6899,N_6477,N_6168);
nand U6900 (N_6900,N_6250,N_6494);
or U6901 (N_6901,N_6062,N_6484);
nor U6902 (N_6902,N_6127,N_6376);
nand U6903 (N_6903,N_6332,N_6008);
nand U6904 (N_6904,N_6077,N_6275);
nand U6905 (N_6905,N_6054,N_6316);
and U6906 (N_6906,N_6077,N_6098);
or U6907 (N_6907,N_6310,N_6259);
and U6908 (N_6908,N_6466,N_6249);
and U6909 (N_6909,N_6250,N_6202);
or U6910 (N_6910,N_6369,N_6487);
xor U6911 (N_6911,N_6025,N_6172);
xnor U6912 (N_6912,N_6193,N_6044);
nor U6913 (N_6913,N_6206,N_6427);
and U6914 (N_6914,N_6197,N_6165);
xor U6915 (N_6915,N_6453,N_6320);
nand U6916 (N_6916,N_6300,N_6216);
nand U6917 (N_6917,N_6316,N_6194);
xor U6918 (N_6918,N_6197,N_6044);
nor U6919 (N_6919,N_6181,N_6229);
or U6920 (N_6920,N_6205,N_6182);
or U6921 (N_6921,N_6297,N_6088);
nand U6922 (N_6922,N_6442,N_6436);
nor U6923 (N_6923,N_6076,N_6167);
or U6924 (N_6924,N_6302,N_6258);
xor U6925 (N_6925,N_6192,N_6233);
xor U6926 (N_6926,N_6333,N_6337);
nor U6927 (N_6927,N_6120,N_6036);
xnor U6928 (N_6928,N_6131,N_6399);
nand U6929 (N_6929,N_6454,N_6005);
or U6930 (N_6930,N_6245,N_6406);
xnor U6931 (N_6931,N_6488,N_6340);
or U6932 (N_6932,N_6016,N_6348);
and U6933 (N_6933,N_6182,N_6019);
nor U6934 (N_6934,N_6400,N_6279);
nor U6935 (N_6935,N_6491,N_6131);
nor U6936 (N_6936,N_6093,N_6120);
or U6937 (N_6937,N_6137,N_6478);
xnor U6938 (N_6938,N_6491,N_6363);
nor U6939 (N_6939,N_6242,N_6444);
nand U6940 (N_6940,N_6348,N_6299);
xor U6941 (N_6941,N_6123,N_6425);
or U6942 (N_6942,N_6054,N_6124);
and U6943 (N_6943,N_6118,N_6464);
xnor U6944 (N_6944,N_6045,N_6164);
or U6945 (N_6945,N_6034,N_6310);
nand U6946 (N_6946,N_6341,N_6473);
nand U6947 (N_6947,N_6476,N_6042);
nand U6948 (N_6948,N_6408,N_6445);
and U6949 (N_6949,N_6181,N_6027);
xnor U6950 (N_6950,N_6436,N_6136);
xor U6951 (N_6951,N_6342,N_6419);
nor U6952 (N_6952,N_6032,N_6015);
and U6953 (N_6953,N_6361,N_6451);
or U6954 (N_6954,N_6204,N_6055);
or U6955 (N_6955,N_6371,N_6083);
nor U6956 (N_6956,N_6184,N_6252);
and U6957 (N_6957,N_6499,N_6392);
nand U6958 (N_6958,N_6026,N_6423);
or U6959 (N_6959,N_6071,N_6475);
or U6960 (N_6960,N_6437,N_6431);
nor U6961 (N_6961,N_6390,N_6470);
nand U6962 (N_6962,N_6287,N_6314);
nand U6963 (N_6963,N_6046,N_6040);
nor U6964 (N_6964,N_6156,N_6467);
nand U6965 (N_6965,N_6095,N_6158);
nand U6966 (N_6966,N_6383,N_6126);
or U6967 (N_6967,N_6295,N_6040);
xor U6968 (N_6968,N_6181,N_6133);
nor U6969 (N_6969,N_6019,N_6288);
nor U6970 (N_6970,N_6016,N_6216);
nor U6971 (N_6971,N_6066,N_6292);
xor U6972 (N_6972,N_6389,N_6281);
nor U6973 (N_6973,N_6308,N_6039);
xnor U6974 (N_6974,N_6432,N_6186);
xor U6975 (N_6975,N_6175,N_6142);
nor U6976 (N_6976,N_6469,N_6470);
or U6977 (N_6977,N_6429,N_6231);
or U6978 (N_6978,N_6254,N_6278);
nand U6979 (N_6979,N_6314,N_6283);
nand U6980 (N_6980,N_6218,N_6319);
or U6981 (N_6981,N_6481,N_6139);
xor U6982 (N_6982,N_6306,N_6145);
nand U6983 (N_6983,N_6384,N_6304);
nor U6984 (N_6984,N_6471,N_6362);
and U6985 (N_6985,N_6144,N_6393);
or U6986 (N_6986,N_6318,N_6326);
and U6987 (N_6987,N_6290,N_6368);
and U6988 (N_6988,N_6119,N_6258);
and U6989 (N_6989,N_6383,N_6400);
or U6990 (N_6990,N_6228,N_6473);
nor U6991 (N_6991,N_6459,N_6369);
and U6992 (N_6992,N_6415,N_6078);
or U6993 (N_6993,N_6258,N_6057);
xnor U6994 (N_6994,N_6058,N_6324);
and U6995 (N_6995,N_6423,N_6133);
and U6996 (N_6996,N_6211,N_6479);
nor U6997 (N_6997,N_6383,N_6245);
nand U6998 (N_6998,N_6341,N_6258);
xnor U6999 (N_6999,N_6378,N_6122);
or U7000 (N_7000,N_6776,N_6881);
and U7001 (N_7001,N_6779,N_6733);
or U7002 (N_7002,N_6859,N_6511);
and U7003 (N_7003,N_6633,N_6685);
xnor U7004 (N_7004,N_6599,N_6508);
xnor U7005 (N_7005,N_6564,N_6600);
and U7006 (N_7006,N_6557,N_6801);
and U7007 (N_7007,N_6762,N_6648);
and U7008 (N_7008,N_6874,N_6954);
and U7009 (N_7009,N_6837,N_6532);
xor U7010 (N_7010,N_6937,N_6763);
and U7011 (N_7011,N_6899,N_6939);
and U7012 (N_7012,N_6690,N_6624);
and U7013 (N_7013,N_6549,N_6840);
or U7014 (N_7014,N_6616,N_6635);
or U7015 (N_7015,N_6523,N_6867);
or U7016 (N_7016,N_6876,N_6702);
xor U7017 (N_7017,N_6868,N_6521);
nand U7018 (N_7018,N_6670,N_6646);
nor U7019 (N_7019,N_6584,N_6816);
or U7020 (N_7020,N_6975,N_6655);
nor U7021 (N_7021,N_6796,N_6767);
and U7022 (N_7022,N_6673,N_6585);
nor U7023 (N_7023,N_6577,N_6922);
nand U7024 (N_7024,N_6708,N_6669);
nand U7025 (N_7025,N_6955,N_6548);
and U7026 (N_7026,N_6788,N_6632);
and U7027 (N_7027,N_6649,N_6977);
and U7028 (N_7028,N_6713,N_6596);
or U7029 (N_7029,N_6674,N_6927);
nor U7030 (N_7030,N_6808,N_6663);
and U7031 (N_7031,N_6567,N_6880);
nor U7032 (N_7032,N_6964,N_6550);
nand U7033 (N_7033,N_6643,N_6565);
nor U7034 (N_7034,N_6513,N_6810);
nor U7035 (N_7035,N_6902,N_6667);
nor U7036 (N_7036,N_6765,N_6684);
nand U7037 (N_7037,N_6652,N_6895);
xnor U7038 (N_7038,N_6898,N_6593);
or U7039 (N_7039,N_6682,N_6651);
and U7040 (N_7040,N_6869,N_6798);
or U7041 (N_7041,N_6724,N_6891);
nand U7042 (N_7042,N_6501,N_6835);
nor U7043 (N_7043,N_6625,N_6510);
xor U7044 (N_7044,N_6985,N_6570);
or U7045 (N_7045,N_6631,N_6996);
or U7046 (N_7046,N_6642,N_6709);
or U7047 (N_7047,N_6863,N_6664);
and U7048 (N_7048,N_6871,N_6644);
nand U7049 (N_7049,N_6589,N_6901);
or U7050 (N_7050,N_6700,N_6780);
and U7051 (N_7051,N_6703,N_6858);
and U7052 (N_7052,N_6615,N_6877);
xor U7053 (N_7053,N_6785,N_6935);
nand U7054 (N_7054,N_6768,N_6744);
or U7055 (N_7055,N_6998,N_6572);
xor U7056 (N_7056,N_6919,N_6515);
nor U7057 (N_7057,N_6750,N_6614);
nor U7058 (N_7058,N_6875,N_6806);
nor U7059 (N_7059,N_6719,N_6936);
nand U7060 (N_7060,N_6647,N_6541);
and U7061 (N_7061,N_6830,N_6607);
nor U7062 (N_7062,N_6571,N_6578);
and U7063 (N_7063,N_6842,N_6759);
or U7064 (N_7064,N_6710,N_6587);
xnor U7065 (N_7065,N_6883,N_6712);
nand U7066 (N_7066,N_6591,N_6626);
and U7067 (N_7067,N_6974,N_6641);
nor U7068 (N_7068,N_6793,N_6752);
nor U7069 (N_7069,N_6561,N_6732);
nor U7070 (N_7070,N_6925,N_6637);
nand U7071 (N_7071,N_6993,N_6848);
nand U7072 (N_7072,N_6535,N_6604);
and U7073 (N_7073,N_6613,N_6654);
nor U7074 (N_7074,N_6911,N_6660);
and U7075 (N_7075,N_6952,N_6560);
nor U7076 (N_7076,N_6723,N_6745);
and U7077 (N_7077,N_6849,N_6617);
and U7078 (N_7078,N_6672,N_6562);
nor U7079 (N_7079,N_6915,N_6524);
xnor U7080 (N_7080,N_6980,N_6692);
nand U7081 (N_7081,N_6804,N_6928);
or U7082 (N_7082,N_6802,N_6807);
nand U7083 (N_7083,N_6695,N_6716);
and U7084 (N_7084,N_6857,N_6675);
or U7085 (N_7085,N_6971,N_6558);
or U7086 (N_7086,N_6543,N_6687);
or U7087 (N_7087,N_6630,N_6887);
nor U7088 (N_7088,N_6627,N_6742);
nand U7089 (N_7089,N_6892,N_6997);
nand U7090 (N_7090,N_6951,N_6963);
and U7091 (N_7091,N_6882,N_6686);
nor U7092 (N_7092,N_6976,N_6729);
nor U7093 (N_7093,N_6934,N_6610);
xor U7094 (N_7094,N_6579,N_6966);
and U7095 (N_7095,N_6984,N_6846);
xnor U7096 (N_7096,N_6705,N_6715);
or U7097 (N_7097,N_6525,N_6845);
nand U7098 (N_7098,N_6896,N_6870);
nand U7099 (N_7099,N_6539,N_6989);
and U7100 (N_7100,N_6872,N_6605);
nor U7101 (N_7101,N_6847,N_6906);
or U7102 (N_7102,N_6711,N_6706);
or U7103 (N_7103,N_6965,N_6961);
nand U7104 (N_7104,N_6754,N_6988);
or U7105 (N_7105,N_6897,N_6661);
xnor U7106 (N_7106,N_6833,N_6940);
or U7107 (N_7107,N_6799,N_6540);
or U7108 (N_7108,N_6755,N_6926);
xor U7109 (N_7109,N_6512,N_6739);
nand U7110 (N_7110,N_6638,N_6582);
or U7111 (N_7111,N_6812,N_6611);
or U7112 (N_7112,N_6517,N_6653);
or U7113 (N_7113,N_6753,N_6597);
and U7114 (N_7114,N_6693,N_6516);
and U7115 (N_7115,N_6628,N_6932);
and U7116 (N_7116,N_6553,N_6916);
or U7117 (N_7117,N_6666,N_6778);
and U7118 (N_7118,N_6677,N_6990);
nand U7119 (N_7119,N_6618,N_6884);
or U7120 (N_7120,N_6865,N_6789);
or U7121 (N_7121,N_6691,N_6978);
nor U7122 (N_7122,N_6608,N_6878);
or U7123 (N_7123,N_6639,N_6592);
xnor U7124 (N_7124,N_6844,N_6995);
or U7125 (N_7125,N_6931,N_6533);
nor U7126 (N_7126,N_6791,N_6542);
nor U7127 (N_7127,N_6757,N_6609);
nor U7128 (N_7128,N_6656,N_6679);
nor U7129 (N_7129,N_6736,N_6590);
xnor U7130 (N_7130,N_6683,N_6576);
and U7131 (N_7131,N_6718,N_6790);
xor U7132 (N_7132,N_6629,N_6770);
nand U7133 (N_7133,N_6960,N_6853);
nor U7134 (N_7134,N_6894,N_6914);
nor U7135 (N_7135,N_6900,N_6601);
nor U7136 (N_7136,N_6697,N_6879);
and U7137 (N_7137,N_6938,N_6634);
nand U7138 (N_7138,N_6738,N_6886);
nor U7139 (N_7139,N_6657,N_6817);
nor U7140 (N_7140,N_6529,N_6509);
or U7141 (N_7141,N_6764,N_6851);
nor U7142 (N_7142,N_6982,N_6544);
xnor U7143 (N_7143,N_6704,N_6586);
or U7144 (N_7144,N_6740,N_6559);
or U7145 (N_7145,N_6820,N_6773);
nor U7146 (N_7146,N_6502,N_6803);
nor U7147 (N_7147,N_6813,N_6930);
nand U7148 (N_7148,N_6566,N_6825);
nand U7149 (N_7149,N_6786,N_6968);
and U7150 (N_7150,N_6536,N_6749);
nand U7151 (N_7151,N_6782,N_6504);
nand U7152 (N_7152,N_6531,N_6546);
or U7153 (N_7153,N_6743,N_6956);
nand U7154 (N_7154,N_6580,N_6507);
xor U7155 (N_7155,N_6819,N_6575);
nor U7156 (N_7156,N_6747,N_6866);
xor U7157 (N_7157,N_6962,N_6522);
xor U7158 (N_7158,N_6621,N_6904);
nor U7159 (N_7159,N_6979,N_6707);
xor U7160 (N_7160,N_6717,N_6855);
or U7161 (N_7161,N_6574,N_6918);
nand U7162 (N_7162,N_6603,N_6760);
or U7163 (N_7163,N_6885,N_6689);
and U7164 (N_7164,N_6699,N_6841);
xnor U7165 (N_7165,N_6727,N_6766);
nand U7166 (N_7166,N_6843,N_6698);
xnor U7167 (N_7167,N_6714,N_6973);
or U7168 (N_7168,N_6528,N_6772);
nand U7169 (N_7169,N_6581,N_6944);
or U7170 (N_7170,N_6573,N_6720);
nor U7171 (N_7171,N_6838,N_6983);
and U7172 (N_7172,N_6913,N_6889);
or U7173 (N_7173,N_6924,N_6726);
and U7174 (N_7174,N_6505,N_6828);
or U7175 (N_7175,N_6545,N_6781);
and U7176 (N_7176,N_6805,N_6769);
or U7177 (N_7177,N_6551,N_6506);
or U7178 (N_7178,N_6758,N_6751);
nand U7179 (N_7179,N_6795,N_6933);
or U7180 (N_7180,N_6731,N_6537);
or U7181 (N_7181,N_6734,N_6834);
xnor U7182 (N_7182,N_6905,N_6862);
nand U7183 (N_7183,N_6598,N_6994);
or U7184 (N_7184,N_6595,N_6777);
or U7185 (N_7185,N_6696,N_6622);
xor U7186 (N_7186,N_6526,N_6948);
nand U7187 (N_7187,N_6722,N_6908);
and U7188 (N_7188,N_6568,N_6873);
xnor U7189 (N_7189,N_6999,N_6518);
xor U7190 (N_7190,N_6829,N_6917);
nand U7191 (N_7191,N_6730,N_6864);
nand U7192 (N_7192,N_6890,N_6893);
and U7193 (N_7193,N_6678,N_6823);
xnor U7194 (N_7194,N_6556,N_6921);
or U7195 (N_7195,N_6746,N_6991);
xor U7196 (N_7196,N_6583,N_6694);
or U7197 (N_7197,N_6784,N_6552);
nor U7198 (N_7198,N_6671,N_6688);
nand U7199 (N_7199,N_6721,N_6821);
or U7200 (N_7200,N_6903,N_6809);
or U7201 (N_7201,N_6554,N_6792);
nor U7202 (N_7202,N_6555,N_6662);
nand U7203 (N_7203,N_6594,N_6665);
or U7204 (N_7204,N_6668,N_6981);
or U7205 (N_7205,N_6748,N_6958);
xnor U7206 (N_7206,N_6826,N_6815);
nand U7207 (N_7207,N_6923,N_6602);
nand U7208 (N_7208,N_6907,N_6645);
xor U7209 (N_7209,N_6850,N_6527);
nor U7210 (N_7210,N_6854,N_6910);
or U7211 (N_7211,N_6623,N_6852);
nor U7212 (N_7212,N_6827,N_6658);
nand U7213 (N_7213,N_6619,N_6503);
and U7214 (N_7214,N_6839,N_6860);
or U7215 (N_7215,N_6500,N_6728);
nor U7216 (N_7216,N_6945,N_6969);
nor U7217 (N_7217,N_6588,N_6681);
nor U7218 (N_7218,N_6797,N_6929);
or U7219 (N_7219,N_6676,N_6972);
or U7220 (N_7220,N_6831,N_6970);
nor U7221 (N_7221,N_6774,N_6912);
or U7222 (N_7222,N_6650,N_6836);
xnor U7223 (N_7223,N_6538,N_6761);
nand U7224 (N_7224,N_6606,N_6959);
xor U7225 (N_7225,N_6992,N_6741);
and U7226 (N_7226,N_6950,N_6701);
or U7227 (N_7227,N_6640,N_6547);
and U7228 (N_7228,N_6680,N_6856);
xnor U7229 (N_7229,N_6953,N_6800);
nand U7230 (N_7230,N_6947,N_6957);
or U7231 (N_7231,N_6775,N_6659);
or U7232 (N_7232,N_6949,N_6756);
nand U7233 (N_7233,N_6987,N_6818);
or U7234 (N_7234,N_6920,N_6519);
and U7235 (N_7235,N_6620,N_6530);
nor U7236 (N_7236,N_6824,N_6771);
or U7237 (N_7237,N_6946,N_6737);
or U7238 (N_7238,N_6725,N_6811);
xor U7239 (N_7239,N_6612,N_6942);
and U7240 (N_7240,N_6814,N_6735);
xnor U7241 (N_7241,N_6822,N_6888);
nand U7242 (N_7242,N_6909,N_6794);
or U7243 (N_7243,N_6520,N_6943);
xnor U7244 (N_7244,N_6986,N_6787);
xnor U7245 (N_7245,N_6783,N_6636);
nor U7246 (N_7246,N_6967,N_6534);
xor U7247 (N_7247,N_6832,N_6514);
nor U7248 (N_7248,N_6941,N_6563);
and U7249 (N_7249,N_6861,N_6569);
and U7250 (N_7250,N_6968,N_6719);
nor U7251 (N_7251,N_6664,N_6875);
and U7252 (N_7252,N_6840,N_6508);
and U7253 (N_7253,N_6647,N_6813);
and U7254 (N_7254,N_6616,N_6516);
nor U7255 (N_7255,N_6984,N_6729);
nor U7256 (N_7256,N_6516,N_6939);
nor U7257 (N_7257,N_6872,N_6526);
nand U7258 (N_7258,N_6803,N_6967);
and U7259 (N_7259,N_6995,N_6736);
xor U7260 (N_7260,N_6850,N_6914);
or U7261 (N_7261,N_6507,N_6626);
or U7262 (N_7262,N_6870,N_6731);
xnor U7263 (N_7263,N_6722,N_6522);
nand U7264 (N_7264,N_6672,N_6797);
nand U7265 (N_7265,N_6625,N_6931);
xor U7266 (N_7266,N_6982,N_6832);
and U7267 (N_7267,N_6948,N_6987);
xor U7268 (N_7268,N_6511,N_6587);
nand U7269 (N_7269,N_6639,N_6748);
and U7270 (N_7270,N_6510,N_6671);
and U7271 (N_7271,N_6527,N_6650);
xor U7272 (N_7272,N_6983,N_6775);
nand U7273 (N_7273,N_6901,N_6687);
nand U7274 (N_7274,N_6861,N_6896);
xnor U7275 (N_7275,N_6635,N_6883);
nor U7276 (N_7276,N_6535,N_6813);
nand U7277 (N_7277,N_6697,N_6680);
nor U7278 (N_7278,N_6906,N_6793);
nor U7279 (N_7279,N_6916,N_6687);
nand U7280 (N_7280,N_6666,N_6625);
xor U7281 (N_7281,N_6926,N_6943);
xnor U7282 (N_7282,N_6601,N_6668);
xnor U7283 (N_7283,N_6650,N_6861);
or U7284 (N_7284,N_6719,N_6515);
and U7285 (N_7285,N_6679,N_6739);
or U7286 (N_7286,N_6628,N_6533);
or U7287 (N_7287,N_6911,N_6800);
or U7288 (N_7288,N_6615,N_6571);
xor U7289 (N_7289,N_6630,N_6515);
or U7290 (N_7290,N_6824,N_6525);
xor U7291 (N_7291,N_6515,N_6903);
or U7292 (N_7292,N_6623,N_6835);
or U7293 (N_7293,N_6833,N_6784);
nor U7294 (N_7294,N_6959,N_6662);
and U7295 (N_7295,N_6521,N_6690);
nor U7296 (N_7296,N_6605,N_6791);
and U7297 (N_7297,N_6855,N_6711);
xor U7298 (N_7298,N_6522,N_6866);
or U7299 (N_7299,N_6693,N_6843);
or U7300 (N_7300,N_6703,N_6822);
and U7301 (N_7301,N_6959,N_6625);
nor U7302 (N_7302,N_6955,N_6780);
nor U7303 (N_7303,N_6527,N_6859);
xnor U7304 (N_7304,N_6544,N_6697);
xor U7305 (N_7305,N_6901,N_6831);
or U7306 (N_7306,N_6582,N_6526);
or U7307 (N_7307,N_6629,N_6724);
and U7308 (N_7308,N_6564,N_6511);
nand U7309 (N_7309,N_6734,N_6896);
or U7310 (N_7310,N_6900,N_6851);
nor U7311 (N_7311,N_6763,N_6902);
nor U7312 (N_7312,N_6710,N_6980);
and U7313 (N_7313,N_6645,N_6935);
nand U7314 (N_7314,N_6823,N_6580);
nand U7315 (N_7315,N_6624,N_6563);
nand U7316 (N_7316,N_6531,N_6610);
xor U7317 (N_7317,N_6656,N_6994);
nor U7318 (N_7318,N_6639,N_6665);
xnor U7319 (N_7319,N_6836,N_6626);
xor U7320 (N_7320,N_6728,N_6874);
nand U7321 (N_7321,N_6579,N_6891);
nor U7322 (N_7322,N_6887,N_6712);
and U7323 (N_7323,N_6900,N_6724);
xor U7324 (N_7324,N_6649,N_6934);
nand U7325 (N_7325,N_6556,N_6886);
or U7326 (N_7326,N_6630,N_6682);
nor U7327 (N_7327,N_6590,N_6729);
nor U7328 (N_7328,N_6931,N_6666);
nand U7329 (N_7329,N_6954,N_6790);
or U7330 (N_7330,N_6747,N_6814);
and U7331 (N_7331,N_6828,N_6678);
nand U7332 (N_7332,N_6869,N_6857);
and U7333 (N_7333,N_6728,N_6557);
xor U7334 (N_7334,N_6589,N_6619);
or U7335 (N_7335,N_6588,N_6601);
and U7336 (N_7336,N_6711,N_6761);
xor U7337 (N_7337,N_6547,N_6854);
nor U7338 (N_7338,N_6796,N_6603);
nand U7339 (N_7339,N_6559,N_6510);
and U7340 (N_7340,N_6714,N_6512);
xor U7341 (N_7341,N_6510,N_6868);
nand U7342 (N_7342,N_6638,N_6846);
or U7343 (N_7343,N_6615,N_6631);
xor U7344 (N_7344,N_6527,N_6836);
nand U7345 (N_7345,N_6537,N_6861);
nand U7346 (N_7346,N_6943,N_6677);
nand U7347 (N_7347,N_6650,N_6749);
and U7348 (N_7348,N_6649,N_6764);
and U7349 (N_7349,N_6890,N_6620);
and U7350 (N_7350,N_6697,N_6918);
xnor U7351 (N_7351,N_6902,N_6976);
nor U7352 (N_7352,N_6682,N_6718);
xor U7353 (N_7353,N_6628,N_6794);
nor U7354 (N_7354,N_6517,N_6659);
or U7355 (N_7355,N_6681,N_6855);
and U7356 (N_7356,N_6921,N_6842);
or U7357 (N_7357,N_6965,N_6523);
or U7358 (N_7358,N_6621,N_6934);
nor U7359 (N_7359,N_6611,N_6596);
nand U7360 (N_7360,N_6774,N_6656);
xor U7361 (N_7361,N_6565,N_6764);
and U7362 (N_7362,N_6820,N_6774);
and U7363 (N_7363,N_6655,N_6956);
xnor U7364 (N_7364,N_6861,N_6967);
or U7365 (N_7365,N_6644,N_6638);
or U7366 (N_7366,N_6731,N_6728);
or U7367 (N_7367,N_6812,N_6981);
nor U7368 (N_7368,N_6543,N_6851);
nor U7369 (N_7369,N_6555,N_6966);
nor U7370 (N_7370,N_6735,N_6726);
and U7371 (N_7371,N_6752,N_6667);
or U7372 (N_7372,N_6540,N_6776);
or U7373 (N_7373,N_6778,N_6524);
nor U7374 (N_7374,N_6764,N_6807);
nand U7375 (N_7375,N_6590,N_6997);
xor U7376 (N_7376,N_6701,N_6926);
xor U7377 (N_7377,N_6621,N_6850);
nor U7378 (N_7378,N_6688,N_6928);
nor U7379 (N_7379,N_6720,N_6835);
and U7380 (N_7380,N_6685,N_6907);
and U7381 (N_7381,N_6551,N_6784);
nand U7382 (N_7382,N_6849,N_6952);
xor U7383 (N_7383,N_6981,N_6990);
nor U7384 (N_7384,N_6691,N_6717);
nor U7385 (N_7385,N_6548,N_6779);
nand U7386 (N_7386,N_6572,N_6700);
nor U7387 (N_7387,N_6980,N_6850);
and U7388 (N_7388,N_6941,N_6910);
nand U7389 (N_7389,N_6779,N_6571);
or U7390 (N_7390,N_6519,N_6924);
nor U7391 (N_7391,N_6867,N_6578);
xnor U7392 (N_7392,N_6735,N_6783);
or U7393 (N_7393,N_6741,N_6578);
nor U7394 (N_7394,N_6888,N_6993);
nand U7395 (N_7395,N_6564,N_6594);
nand U7396 (N_7396,N_6726,N_6712);
nand U7397 (N_7397,N_6703,N_6984);
nand U7398 (N_7398,N_6790,N_6871);
nand U7399 (N_7399,N_6827,N_6638);
xor U7400 (N_7400,N_6871,N_6830);
and U7401 (N_7401,N_6662,N_6778);
nand U7402 (N_7402,N_6955,N_6528);
and U7403 (N_7403,N_6676,N_6819);
or U7404 (N_7404,N_6980,N_6724);
xor U7405 (N_7405,N_6556,N_6566);
nand U7406 (N_7406,N_6757,N_6812);
nand U7407 (N_7407,N_6628,N_6661);
nor U7408 (N_7408,N_6632,N_6865);
xnor U7409 (N_7409,N_6892,N_6840);
or U7410 (N_7410,N_6751,N_6520);
and U7411 (N_7411,N_6553,N_6938);
nor U7412 (N_7412,N_6532,N_6975);
nand U7413 (N_7413,N_6678,N_6925);
nor U7414 (N_7414,N_6772,N_6815);
nor U7415 (N_7415,N_6667,N_6595);
or U7416 (N_7416,N_6965,N_6702);
nand U7417 (N_7417,N_6640,N_6552);
and U7418 (N_7418,N_6578,N_6616);
nand U7419 (N_7419,N_6645,N_6975);
nor U7420 (N_7420,N_6874,N_6584);
and U7421 (N_7421,N_6994,N_6995);
nor U7422 (N_7422,N_6900,N_6529);
nor U7423 (N_7423,N_6642,N_6688);
and U7424 (N_7424,N_6698,N_6830);
nand U7425 (N_7425,N_6624,N_6813);
xnor U7426 (N_7426,N_6907,N_6737);
nor U7427 (N_7427,N_6923,N_6670);
or U7428 (N_7428,N_6852,N_6797);
and U7429 (N_7429,N_6613,N_6735);
nand U7430 (N_7430,N_6671,N_6664);
nor U7431 (N_7431,N_6648,N_6747);
and U7432 (N_7432,N_6793,N_6820);
xor U7433 (N_7433,N_6787,N_6703);
nand U7434 (N_7434,N_6952,N_6847);
xnor U7435 (N_7435,N_6785,N_6831);
and U7436 (N_7436,N_6970,N_6529);
and U7437 (N_7437,N_6887,N_6813);
nand U7438 (N_7438,N_6871,N_6502);
xnor U7439 (N_7439,N_6962,N_6882);
nor U7440 (N_7440,N_6550,N_6982);
nand U7441 (N_7441,N_6991,N_6642);
xor U7442 (N_7442,N_6514,N_6549);
nand U7443 (N_7443,N_6567,N_6873);
xnor U7444 (N_7444,N_6572,N_6766);
and U7445 (N_7445,N_6861,N_6689);
and U7446 (N_7446,N_6879,N_6944);
and U7447 (N_7447,N_6732,N_6558);
nand U7448 (N_7448,N_6851,N_6517);
nand U7449 (N_7449,N_6878,N_6789);
nor U7450 (N_7450,N_6760,N_6860);
nand U7451 (N_7451,N_6592,N_6912);
nor U7452 (N_7452,N_6887,N_6732);
or U7453 (N_7453,N_6816,N_6990);
xor U7454 (N_7454,N_6950,N_6699);
nand U7455 (N_7455,N_6606,N_6561);
and U7456 (N_7456,N_6857,N_6688);
or U7457 (N_7457,N_6625,N_6925);
xnor U7458 (N_7458,N_6971,N_6515);
or U7459 (N_7459,N_6781,N_6842);
and U7460 (N_7460,N_6991,N_6617);
and U7461 (N_7461,N_6791,N_6975);
nand U7462 (N_7462,N_6661,N_6691);
nor U7463 (N_7463,N_6634,N_6501);
nor U7464 (N_7464,N_6520,N_6876);
xor U7465 (N_7465,N_6695,N_6737);
nor U7466 (N_7466,N_6531,N_6938);
xnor U7467 (N_7467,N_6786,N_6855);
and U7468 (N_7468,N_6828,N_6778);
nand U7469 (N_7469,N_6828,N_6999);
and U7470 (N_7470,N_6647,N_6629);
nand U7471 (N_7471,N_6550,N_6838);
and U7472 (N_7472,N_6526,N_6687);
and U7473 (N_7473,N_6537,N_6551);
nor U7474 (N_7474,N_6612,N_6751);
or U7475 (N_7475,N_6980,N_6502);
or U7476 (N_7476,N_6547,N_6985);
and U7477 (N_7477,N_6592,N_6616);
nand U7478 (N_7478,N_6596,N_6598);
nand U7479 (N_7479,N_6957,N_6861);
and U7480 (N_7480,N_6657,N_6562);
xor U7481 (N_7481,N_6811,N_6852);
or U7482 (N_7482,N_6746,N_6878);
and U7483 (N_7483,N_6513,N_6818);
xnor U7484 (N_7484,N_6820,N_6545);
and U7485 (N_7485,N_6562,N_6917);
or U7486 (N_7486,N_6740,N_6802);
and U7487 (N_7487,N_6678,N_6887);
and U7488 (N_7488,N_6693,N_6895);
xnor U7489 (N_7489,N_6588,N_6555);
nor U7490 (N_7490,N_6831,N_6838);
nor U7491 (N_7491,N_6982,N_6873);
nor U7492 (N_7492,N_6835,N_6761);
xor U7493 (N_7493,N_6629,N_6707);
nor U7494 (N_7494,N_6887,N_6940);
nor U7495 (N_7495,N_6686,N_6518);
nor U7496 (N_7496,N_6676,N_6750);
xnor U7497 (N_7497,N_6707,N_6777);
and U7498 (N_7498,N_6707,N_6502);
and U7499 (N_7499,N_6778,N_6510);
nor U7500 (N_7500,N_7336,N_7494);
nor U7501 (N_7501,N_7146,N_7477);
nand U7502 (N_7502,N_7415,N_7362);
xnor U7503 (N_7503,N_7103,N_7000);
nor U7504 (N_7504,N_7124,N_7021);
nor U7505 (N_7505,N_7212,N_7402);
nand U7506 (N_7506,N_7358,N_7045);
or U7507 (N_7507,N_7126,N_7025);
nor U7508 (N_7508,N_7440,N_7384);
xnor U7509 (N_7509,N_7241,N_7291);
and U7510 (N_7510,N_7267,N_7339);
nor U7511 (N_7511,N_7098,N_7423);
and U7512 (N_7512,N_7024,N_7275);
nand U7513 (N_7513,N_7343,N_7314);
nand U7514 (N_7514,N_7227,N_7006);
nor U7515 (N_7515,N_7054,N_7132);
or U7516 (N_7516,N_7180,N_7020);
nand U7517 (N_7517,N_7127,N_7359);
nor U7518 (N_7518,N_7004,N_7217);
xor U7519 (N_7519,N_7398,N_7156);
and U7520 (N_7520,N_7473,N_7374);
and U7521 (N_7521,N_7026,N_7283);
nand U7522 (N_7522,N_7478,N_7068);
nor U7523 (N_7523,N_7176,N_7226);
and U7524 (N_7524,N_7209,N_7207);
nor U7525 (N_7525,N_7194,N_7095);
nand U7526 (N_7526,N_7173,N_7138);
nor U7527 (N_7527,N_7058,N_7495);
nand U7528 (N_7528,N_7121,N_7438);
xnor U7529 (N_7529,N_7118,N_7360);
nand U7530 (N_7530,N_7282,N_7247);
xor U7531 (N_7531,N_7222,N_7076);
and U7532 (N_7532,N_7040,N_7347);
nand U7533 (N_7533,N_7178,N_7493);
and U7534 (N_7534,N_7220,N_7181);
nand U7535 (N_7535,N_7168,N_7465);
nor U7536 (N_7536,N_7102,N_7299);
nor U7537 (N_7537,N_7412,N_7294);
nor U7538 (N_7538,N_7163,N_7329);
nand U7539 (N_7539,N_7381,N_7462);
or U7540 (N_7540,N_7424,N_7310);
and U7541 (N_7541,N_7376,N_7235);
or U7542 (N_7542,N_7039,N_7104);
or U7543 (N_7543,N_7380,N_7052);
nor U7544 (N_7544,N_7334,N_7474);
nor U7545 (N_7545,N_7453,N_7206);
or U7546 (N_7546,N_7112,N_7169);
and U7547 (N_7547,N_7386,N_7388);
or U7548 (N_7548,N_7298,N_7221);
xnor U7549 (N_7549,N_7147,N_7140);
or U7550 (N_7550,N_7285,N_7117);
or U7551 (N_7551,N_7201,N_7182);
or U7552 (N_7552,N_7466,N_7364);
xnor U7553 (N_7553,N_7165,N_7391);
nor U7554 (N_7554,N_7369,N_7028);
nand U7555 (N_7555,N_7033,N_7136);
nand U7556 (N_7556,N_7489,N_7428);
and U7557 (N_7557,N_7367,N_7481);
nand U7558 (N_7558,N_7332,N_7361);
and U7559 (N_7559,N_7061,N_7430);
and U7560 (N_7560,N_7413,N_7320);
nand U7561 (N_7561,N_7306,N_7442);
nor U7562 (N_7562,N_7010,N_7394);
nand U7563 (N_7563,N_7346,N_7253);
or U7564 (N_7564,N_7326,N_7274);
and U7565 (N_7565,N_7188,N_7036);
or U7566 (N_7566,N_7083,N_7213);
nand U7567 (N_7567,N_7099,N_7301);
nor U7568 (N_7568,N_7436,N_7093);
nor U7569 (N_7569,N_7145,N_7151);
and U7570 (N_7570,N_7480,N_7096);
or U7571 (N_7571,N_7107,N_7086);
nor U7572 (N_7572,N_7189,N_7309);
nor U7573 (N_7573,N_7308,N_7321);
xnor U7574 (N_7574,N_7234,N_7419);
or U7575 (N_7575,N_7268,N_7370);
and U7576 (N_7576,N_7001,N_7342);
and U7577 (N_7577,N_7447,N_7337);
xnor U7578 (N_7578,N_7353,N_7433);
or U7579 (N_7579,N_7479,N_7260);
nor U7580 (N_7580,N_7385,N_7105);
xnor U7581 (N_7581,N_7008,N_7407);
xor U7582 (N_7582,N_7085,N_7292);
nor U7583 (N_7583,N_7141,N_7354);
and U7584 (N_7584,N_7075,N_7435);
or U7585 (N_7585,N_7317,N_7219);
or U7586 (N_7586,N_7200,N_7081);
xnor U7587 (N_7587,N_7451,N_7248);
nand U7588 (N_7588,N_7273,N_7059);
nor U7589 (N_7589,N_7225,N_7312);
nor U7590 (N_7590,N_7431,N_7044);
or U7591 (N_7591,N_7101,N_7390);
nor U7592 (N_7592,N_7202,N_7256);
xor U7593 (N_7593,N_7373,N_7160);
nor U7594 (N_7594,N_7483,N_7457);
nand U7595 (N_7595,N_7452,N_7199);
nand U7596 (N_7596,N_7186,N_7114);
xor U7597 (N_7597,N_7411,N_7356);
and U7598 (N_7598,N_7377,N_7315);
or U7599 (N_7599,N_7257,N_7281);
xor U7600 (N_7600,N_7115,N_7072);
nand U7601 (N_7601,N_7074,N_7456);
nand U7602 (N_7602,N_7497,N_7486);
nand U7603 (N_7603,N_7417,N_7092);
or U7604 (N_7604,N_7392,N_7137);
and U7605 (N_7605,N_7254,N_7322);
and U7606 (N_7606,N_7422,N_7414);
nand U7607 (N_7607,N_7345,N_7454);
or U7608 (N_7608,N_7240,N_7047);
xnor U7609 (N_7609,N_7230,N_7444);
and U7610 (N_7610,N_7149,N_7154);
or U7611 (N_7611,N_7300,N_7064);
and U7612 (N_7612,N_7463,N_7236);
and U7613 (N_7613,N_7327,N_7475);
nor U7614 (N_7614,N_7170,N_7158);
nor U7615 (N_7615,N_7284,N_7249);
xor U7616 (N_7616,N_7122,N_7302);
nor U7617 (N_7617,N_7097,N_7043);
and U7618 (N_7618,N_7079,N_7009);
nor U7619 (N_7619,N_7263,N_7041);
nand U7620 (N_7620,N_7191,N_7077);
and U7621 (N_7621,N_7175,N_7197);
nor U7622 (N_7622,N_7205,N_7153);
and U7623 (N_7623,N_7445,N_7368);
xor U7624 (N_7624,N_7066,N_7437);
and U7625 (N_7625,N_7499,N_7065);
nor U7626 (N_7626,N_7034,N_7090);
or U7627 (N_7627,N_7016,N_7190);
and U7628 (N_7628,N_7379,N_7128);
or U7629 (N_7629,N_7297,N_7461);
nand U7630 (N_7630,N_7100,N_7152);
xnor U7631 (N_7631,N_7211,N_7289);
nand U7632 (N_7632,N_7296,N_7459);
or U7633 (N_7633,N_7303,N_7464);
and U7634 (N_7634,N_7293,N_7214);
xor U7635 (N_7635,N_7401,N_7017);
nand U7636 (N_7636,N_7476,N_7023);
and U7637 (N_7637,N_7488,N_7406);
xor U7638 (N_7638,N_7397,N_7243);
xnor U7639 (N_7639,N_7073,N_7338);
or U7640 (N_7640,N_7487,N_7223);
and U7641 (N_7641,N_7005,N_7266);
or U7642 (N_7642,N_7179,N_7070);
or U7643 (N_7643,N_7088,N_7242);
nand U7644 (N_7644,N_7421,N_7019);
nor U7645 (N_7645,N_7305,N_7426);
xnor U7646 (N_7646,N_7148,N_7166);
and U7647 (N_7647,N_7174,N_7408);
nand U7648 (N_7648,N_7276,N_7049);
xor U7649 (N_7649,N_7255,N_7251);
or U7650 (N_7650,N_7133,N_7144);
nand U7651 (N_7651,N_7395,N_7239);
nand U7652 (N_7652,N_7348,N_7279);
or U7653 (N_7653,N_7113,N_7304);
or U7654 (N_7654,N_7427,N_7371);
and U7655 (N_7655,N_7157,N_7071);
and U7656 (N_7656,N_7446,N_7003);
nand U7657 (N_7657,N_7491,N_7449);
nor U7658 (N_7658,N_7231,N_7011);
nand U7659 (N_7659,N_7027,N_7094);
nand U7660 (N_7660,N_7229,N_7192);
and U7661 (N_7661,N_7051,N_7443);
nor U7662 (N_7662,N_7035,N_7187);
nand U7663 (N_7663,N_7286,N_7029);
and U7664 (N_7664,N_7265,N_7404);
xnor U7665 (N_7665,N_7498,N_7139);
xnor U7666 (N_7666,N_7131,N_7069);
nand U7667 (N_7667,N_7238,N_7307);
nor U7668 (N_7668,N_7484,N_7492);
nor U7669 (N_7669,N_7224,N_7335);
nor U7670 (N_7670,N_7400,N_7375);
xnor U7671 (N_7671,N_7389,N_7357);
nor U7672 (N_7672,N_7272,N_7318);
or U7673 (N_7673,N_7448,N_7067);
xnor U7674 (N_7674,N_7037,N_7172);
nand U7675 (N_7675,N_7429,N_7396);
nor U7676 (N_7676,N_7496,N_7108);
and U7677 (N_7677,N_7387,N_7116);
and U7678 (N_7678,N_7420,N_7363);
xnor U7679 (N_7679,N_7142,N_7366);
or U7680 (N_7680,N_7472,N_7123);
or U7681 (N_7681,N_7167,N_7203);
xor U7682 (N_7682,N_7215,N_7460);
nand U7683 (N_7683,N_7135,N_7485);
xor U7684 (N_7684,N_7164,N_7013);
nand U7685 (N_7685,N_7405,N_7259);
xnor U7686 (N_7686,N_7110,N_7434);
and U7687 (N_7687,N_7355,N_7130);
nand U7688 (N_7688,N_7277,N_7340);
and U7689 (N_7689,N_7288,N_7311);
nor U7690 (N_7690,N_7063,N_7490);
and U7691 (N_7691,N_7204,N_7271);
nand U7692 (N_7692,N_7233,N_7319);
or U7693 (N_7693,N_7055,N_7134);
or U7694 (N_7694,N_7458,N_7007);
xnor U7695 (N_7695,N_7002,N_7014);
xnor U7696 (N_7696,N_7091,N_7393);
nand U7697 (N_7697,N_7352,N_7080);
or U7698 (N_7698,N_7365,N_7150);
nor U7699 (N_7699,N_7171,N_7482);
nand U7700 (N_7700,N_7250,N_7125);
xnor U7701 (N_7701,N_7232,N_7060);
xnor U7702 (N_7702,N_7261,N_7316);
nor U7703 (N_7703,N_7280,N_7210);
or U7704 (N_7704,N_7228,N_7062);
nor U7705 (N_7705,N_7089,N_7295);
and U7706 (N_7706,N_7258,N_7399);
nor U7707 (N_7707,N_7432,N_7469);
nor U7708 (N_7708,N_7198,N_7410);
nand U7709 (N_7709,N_7084,N_7450);
nand U7710 (N_7710,N_7409,N_7031);
nand U7711 (N_7711,N_7159,N_7022);
xor U7712 (N_7712,N_7468,N_7264);
nor U7713 (N_7713,N_7439,N_7120);
or U7714 (N_7714,N_7184,N_7078);
or U7715 (N_7715,N_7046,N_7416);
or U7716 (N_7716,N_7328,N_7030);
nor U7717 (N_7717,N_7341,N_7333);
xnor U7718 (N_7718,N_7467,N_7143);
nand U7719 (N_7719,N_7218,N_7470);
nor U7720 (N_7720,N_7244,N_7050);
nand U7721 (N_7721,N_7042,N_7325);
xnor U7722 (N_7722,N_7425,N_7262);
and U7723 (N_7723,N_7270,N_7441);
or U7724 (N_7724,N_7161,N_7378);
nor U7725 (N_7725,N_7269,N_7109);
xor U7726 (N_7726,N_7313,N_7183);
or U7727 (N_7727,N_7246,N_7290);
nor U7728 (N_7728,N_7349,N_7208);
nor U7729 (N_7729,N_7111,N_7382);
nand U7730 (N_7730,N_7106,N_7119);
or U7731 (N_7731,N_7129,N_7418);
or U7732 (N_7732,N_7252,N_7455);
or U7733 (N_7733,N_7177,N_7018);
nor U7734 (N_7734,N_7185,N_7350);
nand U7735 (N_7735,N_7344,N_7032);
xor U7736 (N_7736,N_7057,N_7155);
or U7737 (N_7737,N_7471,N_7012);
or U7738 (N_7738,N_7351,N_7216);
nand U7739 (N_7739,N_7330,N_7162);
and U7740 (N_7740,N_7323,N_7403);
nand U7741 (N_7741,N_7056,N_7048);
xnor U7742 (N_7742,N_7287,N_7372);
xor U7743 (N_7743,N_7015,N_7324);
nor U7744 (N_7744,N_7237,N_7053);
xor U7745 (N_7745,N_7195,N_7082);
nor U7746 (N_7746,N_7196,N_7087);
and U7747 (N_7747,N_7193,N_7038);
and U7748 (N_7748,N_7245,N_7278);
nor U7749 (N_7749,N_7383,N_7331);
and U7750 (N_7750,N_7173,N_7465);
or U7751 (N_7751,N_7110,N_7048);
xnor U7752 (N_7752,N_7469,N_7070);
nor U7753 (N_7753,N_7320,N_7372);
and U7754 (N_7754,N_7255,N_7379);
nand U7755 (N_7755,N_7433,N_7464);
nand U7756 (N_7756,N_7072,N_7176);
nand U7757 (N_7757,N_7204,N_7477);
nor U7758 (N_7758,N_7017,N_7477);
nand U7759 (N_7759,N_7199,N_7063);
nand U7760 (N_7760,N_7295,N_7152);
nand U7761 (N_7761,N_7217,N_7058);
and U7762 (N_7762,N_7225,N_7425);
or U7763 (N_7763,N_7190,N_7306);
xor U7764 (N_7764,N_7157,N_7451);
nor U7765 (N_7765,N_7154,N_7084);
nand U7766 (N_7766,N_7300,N_7124);
and U7767 (N_7767,N_7166,N_7201);
nand U7768 (N_7768,N_7060,N_7256);
nor U7769 (N_7769,N_7359,N_7399);
nand U7770 (N_7770,N_7494,N_7124);
and U7771 (N_7771,N_7158,N_7047);
or U7772 (N_7772,N_7117,N_7299);
or U7773 (N_7773,N_7185,N_7120);
nor U7774 (N_7774,N_7284,N_7040);
or U7775 (N_7775,N_7040,N_7319);
xnor U7776 (N_7776,N_7495,N_7230);
nor U7777 (N_7777,N_7014,N_7062);
and U7778 (N_7778,N_7134,N_7473);
and U7779 (N_7779,N_7305,N_7422);
and U7780 (N_7780,N_7313,N_7432);
or U7781 (N_7781,N_7232,N_7114);
nand U7782 (N_7782,N_7457,N_7365);
and U7783 (N_7783,N_7394,N_7192);
nand U7784 (N_7784,N_7483,N_7151);
nand U7785 (N_7785,N_7352,N_7163);
xnor U7786 (N_7786,N_7241,N_7298);
nor U7787 (N_7787,N_7096,N_7398);
nand U7788 (N_7788,N_7459,N_7156);
nand U7789 (N_7789,N_7343,N_7089);
xor U7790 (N_7790,N_7201,N_7399);
nand U7791 (N_7791,N_7035,N_7012);
nand U7792 (N_7792,N_7163,N_7083);
and U7793 (N_7793,N_7086,N_7333);
and U7794 (N_7794,N_7002,N_7064);
nand U7795 (N_7795,N_7050,N_7430);
or U7796 (N_7796,N_7227,N_7013);
or U7797 (N_7797,N_7253,N_7379);
and U7798 (N_7798,N_7227,N_7051);
nor U7799 (N_7799,N_7314,N_7232);
or U7800 (N_7800,N_7093,N_7433);
xor U7801 (N_7801,N_7017,N_7375);
and U7802 (N_7802,N_7026,N_7239);
or U7803 (N_7803,N_7108,N_7081);
nand U7804 (N_7804,N_7399,N_7388);
xor U7805 (N_7805,N_7470,N_7314);
or U7806 (N_7806,N_7327,N_7153);
nand U7807 (N_7807,N_7076,N_7179);
nor U7808 (N_7808,N_7022,N_7418);
and U7809 (N_7809,N_7118,N_7346);
nor U7810 (N_7810,N_7214,N_7077);
and U7811 (N_7811,N_7222,N_7201);
nor U7812 (N_7812,N_7221,N_7013);
and U7813 (N_7813,N_7223,N_7434);
or U7814 (N_7814,N_7461,N_7261);
nor U7815 (N_7815,N_7074,N_7335);
nor U7816 (N_7816,N_7387,N_7371);
xnor U7817 (N_7817,N_7287,N_7282);
xor U7818 (N_7818,N_7190,N_7388);
nand U7819 (N_7819,N_7461,N_7223);
or U7820 (N_7820,N_7140,N_7113);
nand U7821 (N_7821,N_7350,N_7016);
xnor U7822 (N_7822,N_7002,N_7327);
nor U7823 (N_7823,N_7358,N_7071);
or U7824 (N_7824,N_7259,N_7420);
nand U7825 (N_7825,N_7296,N_7149);
or U7826 (N_7826,N_7339,N_7095);
and U7827 (N_7827,N_7482,N_7491);
or U7828 (N_7828,N_7289,N_7364);
nand U7829 (N_7829,N_7449,N_7128);
and U7830 (N_7830,N_7039,N_7190);
nor U7831 (N_7831,N_7112,N_7197);
nand U7832 (N_7832,N_7133,N_7052);
or U7833 (N_7833,N_7127,N_7154);
xnor U7834 (N_7834,N_7339,N_7491);
or U7835 (N_7835,N_7250,N_7431);
nor U7836 (N_7836,N_7393,N_7369);
nor U7837 (N_7837,N_7146,N_7387);
or U7838 (N_7838,N_7462,N_7128);
nor U7839 (N_7839,N_7316,N_7305);
nand U7840 (N_7840,N_7235,N_7424);
xor U7841 (N_7841,N_7223,N_7033);
and U7842 (N_7842,N_7040,N_7245);
nor U7843 (N_7843,N_7100,N_7345);
or U7844 (N_7844,N_7246,N_7024);
xor U7845 (N_7845,N_7491,N_7370);
and U7846 (N_7846,N_7212,N_7140);
xor U7847 (N_7847,N_7355,N_7097);
xnor U7848 (N_7848,N_7197,N_7018);
nor U7849 (N_7849,N_7142,N_7145);
or U7850 (N_7850,N_7107,N_7265);
xor U7851 (N_7851,N_7217,N_7266);
or U7852 (N_7852,N_7241,N_7494);
xnor U7853 (N_7853,N_7296,N_7003);
nand U7854 (N_7854,N_7163,N_7172);
nor U7855 (N_7855,N_7126,N_7472);
and U7856 (N_7856,N_7008,N_7257);
nor U7857 (N_7857,N_7370,N_7299);
or U7858 (N_7858,N_7022,N_7464);
or U7859 (N_7859,N_7233,N_7075);
nor U7860 (N_7860,N_7395,N_7343);
nor U7861 (N_7861,N_7067,N_7431);
and U7862 (N_7862,N_7337,N_7355);
or U7863 (N_7863,N_7223,N_7147);
xnor U7864 (N_7864,N_7229,N_7204);
nor U7865 (N_7865,N_7360,N_7057);
xnor U7866 (N_7866,N_7274,N_7028);
or U7867 (N_7867,N_7109,N_7328);
or U7868 (N_7868,N_7121,N_7426);
xnor U7869 (N_7869,N_7114,N_7319);
or U7870 (N_7870,N_7011,N_7158);
or U7871 (N_7871,N_7095,N_7408);
and U7872 (N_7872,N_7414,N_7382);
nand U7873 (N_7873,N_7146,N_7024);
or U7874 (N_7874,N_7138,N_7279);
xnor U7875 (N_7875,N_7297,N_7122);
xnor U7876 (N_7876,N_7420,N_7450);
and U7877 (N_7877,N_7069,N_7032);
nand U7878 (N_7878,N_7328,N_7180);
xor U7879 (N_7879,N_7308,N_7391);
or U7880 (N_7880,N_7205,N_7041);
and U7881 (N_7881,N_7400,N_7069);
nand U7882 (N_7882,N_7258,N_7214);
nor U7883 (N_7883,N_7386,N_7262);
or U7884 (N_7884,N_7328,N_7396);
nand U7885 (N_7885,N_7142,N_7361);
nor U7886 (N_7886,N_7142,N_7255);
nand U7887 (N_7887,N_7217,N_7056);
and U7888 (N_7888,N_7093,N_7349);
nor U7889 (N_7889,N_7349,N_7047);
nand U7890 (N_7890,N_7119,N_7398);
and U7891 (N_7891,N_7090,N_7252);
nor U7892 (N_7892,N_7209,N_7237);
nor U7893 (N_7893,N_7114,N_7202);
nand U7894 (N_7894,N_7286,N_7300);
or U7895 (N_7895,N_7195,N_7070);
nand U7896 (N_7896,N_7048,N_7422);
nor U7897 (N_7897,N_7424,N_7451);
nand U7898 (N_7898,N_7493,N_7266);
or U7899 (N_7899,N_7077,N_7493);
or U7900 (N_7900,N_7106,N_7130);
xnor U7901 (N_7901,N_7004,N_7027);
nor U7902 (N_7902,N_7222,N_7467);
or U7903 (N_7903,N_7013,N_7476);
xnor U7904 (N_7904,N_7024,N_7222);
nand U7905 (N_7905,N_7184,N_7129);
or U7906 (N_7906,N_7036,N_7392);
nor U7907 (N_7907,N_7438,N_7269);
xor U7908 (N_7908,N_7350,N_7402);
xnor U7909 (N_7909,N_7463,N_7402);
nand U7910 (N_7910,N_7035,N_7120);
nand U7911 (N_7911,N_7219,N_7265);
nor U7912 (N_7912,N_7376,N_7099);
and U7913 (N_7913,N_7049,N_7057);
and U7914 (N_7914,N_7428,N_7258);
xor U7915 (N_7915,N_7036,N_7289);
nand U7916 (N_7916,N_7217,N_7462);
or U7917 (N_7917,N_7390,N_7070);
or U7918 (N_7918,N_7064,N_7473);
or U7919 (N_7919,N_7401,N_7121);
xnor U7920 (N_7920,N_7376,N_7170);
and U7921 (N_7921,N_7261,N_7335);
or U7922 (N_7922,N_7478,N_7279);
nand U7923 (N_7923,N_7031,N_7341);
xor U7924 (N_7924,N_7024,N_7153);
and U7925 (N_7925,N_7487,N_7038);
xor U7926 (N_7926,N_7100,N_7029);
or U7927 (N_7927,N_7297,N_7487);
xnor U7928 (N_7928,N_7083,N_7275);
nor U7929 (N_7929,N_7181,N_7167);
nor U7930 (N_7930,N_7095,N_7151);
or U7931 (N_7931,N_7218,N_7247);
or U7932 (N_7932,N_7298,N_7480);
nor U7933 (N_7933,N_7292,N_7007);
xnor U7934 (N_7934,N_7463,N_7406);
nor U7935 (N_7935,N_7079,N_7224);
or U7936 (N_7936,N_7190,N_7348);
nor U7937 (N_7937,N_7060,N_7106);
nor U7938 (N_7938,N_7203,N_7213);
or U7939 (N_7939,N_7129,N_7462);
nor U7940 (N_7940,N_7159,N_7180);
xnor U7941 (N_7941,N_7272,N_7229);
nor U7942 (N_7942,N_7078,N_7352);
xor U7943 (N_7943,N_7422,N_7140);
and U7944 (N_7944,N_7270,N_7242);
or U7945 (N_7945,N_7447,N_7245);
nor U7946 (N_7946,N_7352,N_7246);
nor U7947 (N_7947,N_7027,N_7409);
nor U7948 (N_7948,N_7356,N_7085);
and U7949 (N_7949,N_7381,N_7063);
nand U7950 (N_7950,N_7023,N_7115);
and U7951 (N_7951,N_7284,N_7245);
nor U7952 (N_7952,N_7207,N_7023);
and U7953 (N_7953,N_7163,N_7440);
nor U7954 (N_7954,N_7362,N_7452);
xor U7955 (N_7955,N_7073,N_7317);
xnor U7956 (N_7956,N_7073,N_7242);
nor U7957 (N_7957,N_7430,N_7415);
nor U7958 (N_7958,N_7146,N_7119);
or U7959 (N_7959,N_7159,N_7395);
and U7960 (N_7960,N_7439,N_7483);
xor U7961 (N_7961,N_7121,N_7428);
nand U7962 (N_7962,N_7391,N_7118);
or U7963 (N_7963,N_7370,N_7344);
xor U7964 (N_7964,N_7139,N_7162);
xnor U7965 (N_7965,N_7215,N_7277);
and U7966 (N_7966,N_7136,N_7184);
nor U7967 (N_7967,N_7242,N_7026);
xnor U7968 (N_7968,N_7102,N_7127);
xor U7969 (N_7969,N_7093,N_7319);
or U7970 (N_7970,N_7064,N_7365);
nor U7971 (N_7971,N_7469,N_7338);
or U7972 (N_7972,N_7484,N_7361);
or U7973 (N_7973,N_7167,N_7294);
nand U7974 (N_7974,N_7216,N_7362);
nand U7975 (N_7975,N_7037,N_7131);
and U7976 (N_7976,N_7498,N_7300);
and U7977 (N_7977,N_7270,N_7303);
nand U7978 (N_7978,N_7266,N_7252);
or U7979 (N_7979,N_7467,N_7402);
xor U7980 (N_7980,N_7488,N_7189);
xnor U7981 (N_7981,N_7093,N_7053);
and U7982 (N_7982,N_7258,N_7224);
xor U7983 (N_7983,N_7115,N_7038);
nand U7984 (N_7984,N_7319,N_7293);
and U7985 (N_7985,N_7422,N_7366);
and U7986 (N_7986,N_7144,N_7141);
nand U7987 (N_7987,N_7099,N_7233);
or U7988 (N_7988,N_7079,N_7393);
or U7989 (N_7989,N_7364,N_7134);
xnor U7990 (N_7990,N_7216,N_7241);
nor U7991 (N_7991,N_7015,N_7494);
xor U7992 (N_7992,N_7282,N_7241);
nor U7993 (N_7993,N_7277,N_7363);
nor U7994 (N_7994,N_7178,N_7293);
or U7995 (N_7995,N_7487,N_7457);
nand U7996 (N_7996,N_7446,N_7451);
and U7997 (N_7997,N_7075,N_7492);
nand U7998 (N_7998,N_7437,N_7159);
or U7999 (N_7999,N_7223,N_7385);
or U8000 (N_8000,N_7843,N_7970);
and U8001 (N_8001,N_7599,N_7602);
and U8002 (N_8002,N_7889,N_7900);
or U8003 (N_8003,N_7824,N_7858);
and U8004 (N_8004,N_7543,N_7532);
nor U8005 (N_8005,N_7790,N_7693);
or U8006 (N_8006,N_7964,N_7617);
nand U8007 (N_8007,N_7878,N_7513);
and U8008 (N_8008,N_7819,N_7573);
and U8009 (N_8009,N_7991,N_7833);
or U8010 (N_8010,N_7933,N_7547);
and U8011 (N_8011,N_7590,N_7890);
or U8012 (N_8012,N_7612,N_7868);
xor U8013 (N_8013,N_7982,N_7909);
or U8014 (N_8014,N_7713,N_7511);
or U8015 (N_8015,N_7886,N_7697);
nor U8016 (N_8016,N_7848,N_7540);
and U8017 (N_8017,N_7704,N_7812);
and U8018 (N_8018,N_7947,N_7972);
nand U8019 (N_8019,N_7550,N_7853);
or U8020 (N_8020,N_7649,N_7606);
or U8021 (N_8021,N_7510,N_7971);
and U8022 (N_8022,N_7977,N_7897);
nor U8023 (N_8023,N_7902,N_7891);
nand U8024 (N_8024,N_7930,N_7773);
nand U8025 (N_8025,N_7892,N_7791);
and U8026 (N_8026,N_7944,N_7847);
xnor U8027 (N_8027,N_7870,N_7524);
and U8028 (N_8028,N_7595,N_7554);
nor U8029 (N_8029,N_7685,N_7657);
xor U8030 (N_8030,N_7643,N_7631);
and U8031 (N_8031,N_7894,N_7711);
xor U8032 (N_8032,N_7952,N_7718);
and U8033 (N_8033,N_7586,N_7701);
nand U8034 (N_8034,N_7954,N_7683);
nor U8035 (N_8035,N_7743,N_7899);
xor U8036 (N_8036,N_7572,N_7814);
and U8037 (N_8037,N_7607,N_7968);
nor U8038 (N_8038,N_7929,N_7839);
xor U8039 (N_8039,N_7611,N_7938);
or U8040 (N_8040,N_7915,N_7585);
and U8041 (N_8041,N_7624,N_7809);
or U8042 (N_8042,N_7912,N_7852);
nor U8043 (N_8043,N_7798,N_7598);
xnor U8044 (N_8044,N_7750,N_7605);
nor U8045 (N_8045,N_7733,N_7821);
and U8046 (N_8046,N_7854,N_7862);
nand U8047 (N_8047,N_7731,N_7916);
or U8048 (N_8048,N_7978,N_7951);
nor U8049 (N_8049,N_7741,N_7807);
or U8050 (N_8050,N_7642,N_7725);
or U8051 (N_8051,N_7559,N_7721);
nand U8052 (N_8052,N_7761,N_7734);
nor U8053 (N_8053,N_7776,N_7665);
nor U8054 (N_8054,N_7645,N_7989);
nor U8055 (N_8055,N_7981,N_7580);
and U8056 (N_8056,N_7619,N_7517);
xor U8057 (N_8057,N_7608,N_7804);
nand U8058 (N_8058,N_7980,N_7792);
xor U8059 (N_8059,N_7680,N_7961);
nand U8060 (N_8060,N_7594,N_7647);
or U8061 (N_8061,N_7560,N_7896);
xor U8062 (N_8062,N_7509,N_7566);
or U8063 (N_8063,N_7724,N_7910);
nand U8064 (N_8064,N_7735,N_7615);
or U8065 (N_8065,N_7682,N_7674);
nand U8066 (N_8066,N_7696,N_7652);
nor U8067 (N_8067,N_7635,N_7946);
nand U8068 (N_8068,N_7765,N_7562);
or U8069 (N_8069,N_7775,N_7996);
nor U8070 (N_8070,N_7931,N_7830);
nor U8071 (N_8071,N_7508,N_7687);
nand U8072 (N_8072,N_7739,N_7784);
or U8073 (N_8073,N_7544,N_7815);
or U8074 (N_8074,N_7908,N_7626);
xor U8075 (N_8075,N_7613,N_7770);
or U8076 (N_8076,N_7873,N_7553);
and U8077 (N_8077,N_7979,N_7568);
nor U8078 (N_8078,N_7832,N_7706);
and U8079 (N_8079,N_7575,N_7677);
nor U8080 (N_8080,N_7918,N_7698);
nand U8081 (N_8081,N_7542,N_7849);
xor U8082 (N_8082,N_7884,N_7620);
nand U8083 (N_8083,N_7986,N_7670);
or U8084 (N_8084,N_7905,N_7764);
and U8085 (N_8085,N_7633,N_7831);
nor U8086 (N_8086,N_7686,N_7623);
nand U8087 (N_8087,N_7935,N_7907);
xor U8088 (N_8088,N_7747,N_7926);
or U8089 (N_8089,N_7800,N_7576);
or U8090 (N_8090,N_7692,N_7730);
and U8091 (N_8091,N_7551,N_7880);
and U8092 (N_8092,N_7584,N_7666);
or U8093 (N_8093,N_7936,N_7604);
or U8094 (N_8094,N_7866,N_7529);
nand U8095 (N_8095,N_7879,N_7638);
or U8096 (N_8096,N_7719,N_7563);
xor U8097 (N_8097,N_7664,N_7667);
and U8098 (N_8098,N_7826,N_7537);
and U8099 (N_8099,N_7969,N_7808);
nor U8100 (N_8100,N_7828,N_7835);
nand U8101 (N_8101,N_7766,N_7548);
and U8102 (N_8102,N_7850,N_7787);
xnor U8103 (N_8103,N_7521,N_7903);
nand U8104 (N_8104,N_7588,N_7924);
and U8105 (N_8105,N_7885,N_7882);
nor U8106 (N_8106,N_7813,N_7751);
xor U8107 (N_8107,N_7875,N_7778);
xnor U8108 (N_8108,N_7914,N_7565);
nor U8109 (N_8109,N_7549,N_7834);
or U8110 (N_8110,N_7745,N_7836);
or U8111 (N_8111,N_7581,N_7661);
nand U8112 (N_8112,N_7782,N_7874);
xnor U8113 (N_8113,N_7714,N_7917);
and U8114 (N_8114,N_7934,N_7803);
nor U8115 (N_8115,N_7941,N_7793);
xnor U8116 (N_8116,N_7740,N_7712);
and U8117 (N_8117,N_7520,N_7690);
or U8118 (N_8118,N_7992,N_7865);
and U8119 (N_8119,N_7583,N_7998);
nand U8120 (N_8120,N_7911,N_7653);
nor U8121 (N_8121,N_7597,N_7771);
or U8122 (N_8122,N_7950,N_7997);
and U8123 (N_8123,N_7906,N_7641);
nand U8124 (N_8124,N_7748,N_7956);
nor U8125 (N_8125,N_7558,N_7514);
xnor U8126 (N_8126,N_7700,N_7709);
or U8127 (N_8127,N_7629,N_7546);
xor U8128 (N_8128,N_7987,N_7569);
nor U8129 (N_8129,N_7856,N_7519);
nand U8130 (N_8130,N_7522,N_7837);
xnor U8131 (N_8131,N_7694,N_7654);
and U8132 (N_8132,N_7736,N_7959);
xnor U8133 (N_8133,N_7863,N_7579);
nand U8134 (N_8134,N_7571,N_7867);
xnor U8135 (N_8135,N_7669,N_7846);
and U8136 (N_8136,N_7610,N_7990);
xor U8137 (N_8137,N_7525,N_7772);
nor U8138 (N_8138,N_7715,N_7592);
nor U8139 (N_8139,N_7726,N_7675);
xor U8140 (N_8140,N_7601,N_7634);
xnor U8141 (N_8141,N_7659,N_7855);
or U8142 (N_8142,N_7545,N_7500);
xor U8143 (N_8143,N_7920,N_7744);
xnor U8144 (N_8144,N_7962,N_7753);
xnor U8145 (N_8145,N_7928,N_7769);
nand U8146 (N_8146,N_7561,N_7552);
xor U8147 (N_8147,N_7533,N_7945);
xnor U8148 (N_8148,N_7805,N_7913);
and U8149 (N_8149,N_7636,N_7759);
nand U8150 (N_8150,N_7796,N_7923);
xnor U8151 (N_8151,N_7788,N_7589);
xnor U8152 (N_8152,N_7518,N_7842);
nor U8153 (N_8153,N_7786,N_7948);
nor U8154 (N_8154,N_7555,N_7672);
and U8155 (N_8155,N_7515,N_7976);
xnor U8156 (N_8156,N_7646,N_7795);
nor U8157 (N_8157,N_7707,N_7506);
nand U8158 (N_8158,N_7760,N_7838);
and U8159 (N_8159,N_7816,N_7919);
or U8160 (N_8160,N_7932,N_7628);
nor U8161 (N_8161,N_7527,N_7596);
or U8162 (N_8162,N_7502,N_7621);
xnor U8163 (N_8163,N_7955,N_7671);
and U8164 (N_8164,N_7723,N_7658);
nand U8165 (N_8165,N_7627,N_7785);
and U8166 (N_8166,N_7722,N_7940);
nand U8167 (N_8167,N_7995,N_7966);
nand U8168 (N_8168,N_7869,N_7904);
and U8169 (N_8169,N_7679,N_7802);
xnor U8170 (N_8170,N_7503,N_7799);
and U8171 (N_8171,N_7827,N_7591);
or U8172 (N_8172,N_7818,N_7738);
or U8173 (N_8173,N_7895,N_7825);
nand U8174 (N_8174,N_7953,N_7587);
nand U8175 (N_8175,N_7648,N_7844);
nor U8176 (N_8176,N_7582,N_7681);
nor U8177 (N_8177,N_7660,N_7789);
nor U8178 (N_8178,N_7810,N_7663);
nand U8179 (N_8179,N_7662,N_7777);
and U8180 (N_8180,N_7717,N_7530);
or U8181 (N_8181,N_7535,N_7516);
nor U8182 (N_8182,N_7655,N_7557);
nor U8183 (N_8183,N_7541,N_7603);
xor U8184 (N_8184,N_7767,N_7512);
and U8185 (N_8185,N_7716,N_7942);
nand U8186 (N_8186,N_7994,N_7609);
or U8187 (N_8187,N_7822,N_7965);
xnor U8188 (N_8188,N_7676,N_7746);
nand U8189 (N_8189,N_7806,N_7921);
nor U8190 (N_8190,N_7877,N_7691);
xor U8191 (N_8191,N_7708,N_7673);
nor U8192 (N_8192,N_7695,N_7507);
nor U8193 (N_8193,N_7534,N_7859);
nor U8194 (N_8194,N_7616,N_7531);
nor U8195 (N_8195,N_7757,N_7829);
nand U8196 (N_8196,N_7988,N_7949);
nand U8197 (N_8197,N_7538,N_7539);
nand U8198 (N_8198,N_7556,N_7960);
nor U8199 (N_8199,N_7574,N_7668);
xor U8200 (N_8200,N_7749,N_7630);
or U8201 (N_8201,N_7999,N_7811);
xor U8202 (N_8202,N_7644,N_7857);
and U8203 (N_8203,N_7614,N_7754);
nand U8204 (N_8204,N_7871,N_7689);
or U8205 (N_8205,N_7993,N_7864);
nor U8206 (N_8206,N_7984,N_7567);
nand U8207 (N_8207,N_7876,N_7600);
xor U8208 (N_8208,N_7983,N_7985);
and U8209 (N_8209,N_7505,N_7794);
xor U8210 (N_8210,N_7758,N_7729);
or U8211 (N_8211,N_7841,N_7650);
nand U8212 (N_8212,N_7774,N_7898);
nand U8213 (N_8213,N_7570,N_7887);
xor U8214 (N_8214,N_7779,N_7763);
and U8215 (N_8215,N_7893,N_7737);
or U8216 (N_8216,N_7640,N_7536);
nand U8217 (N_8217,N_7705,N_7922);
or U8218 (N_8218,N_7963,N_7943);
nor U8219 (N_8219,N_7564,N_7925);
nor U8220 (N_8220,N_7501,N_7637);
nand U8221 (N_8221,N_7958,N_7817);
nand U8222 (N_8222,N_7752,N_7861);
or U8223 (N_8223,N_7840,N_7781);
and U8224 (N_8224,N_7688,N_7937);
nand U8225 (N_8225,N_7528,N_7823);
nand U8226 (N_8226,N_7927,N_7768);
and U8227 (N_8227,N_7732,N_7888);
nor U8228 (N_8228,N_7577,N_7756);
nand U8229 (N_8229,N_7703,N_7957);
and U8230 (N_8230,N_7632,N_7578);
and U8231 (N_8231,N_7860,N_7820);
and U8232 (N_8232,N_7625,N_7526);
or U8233 (N_8233,N_7851,N_7523);
or U8234 (N_8234,N_7618,N_7678);
nor U8235 (N_8235,N_7742,N_7710);
nor U8236 (N_8236,N_7762,N_7797);
or U8237 (N_8237,N_7699,N_7720);
xnor U8238 (N_8238,N_7656,N_7639);
xnor U8239 (N_8239,N_7783,N_7684);
nand U8240 (N_8240,N_7755,N_7504);
or U8241 (N_8241,N_7974,N_7973);
and U8242 (N_8242,N_7881,N_7967);
and U8243 (N_8243,N_7872,N_7651);
xor U8244 (N_8244,N_7975,N_7727);
or U8245 (N_8245,N_7780,N_7801);
xnor U8246 (N_8246,N_7939,N_7728);
or U8247 (N_8247,N_7593,N_7622);
or U8248 (N_8248,N_7883,N_7901);
nor U8249 (N_8249,N_7845,N_7702);
and U8250 (N_8250,N_7906,N_7862);
xnor U8251 (N_8251,N_7714,N_7998);
xor U8252 (N_8252,N_7800,N_7586);
and U8253 (N_8253,N_7544,N_7899);
nor U8254 (N_8254,N_7511,N_7978);
xor U8255 (N_8255,N_7648,N_7959);
nand U8256 (N_8256,N_7672,N_7807);
nor U8257 (N_8257,N_7653,N_7773);
nor U8258 (N_8258,N_7614,N_7780);
and U8259 (N_8259,N_7544,N_7834);
or U8260 (N_8260,N_7538,N_7901);
nor U8261 (N_8261,N_7824,N_7685);
and U8262 (N_8262,N_7626,N_7682);
nand U8263 (N_8263,N_7850,N_7635);
or U8264 (N_8264,N_7620,N_7600);
xnor U8265 (N_8265,N_7976,N_7984);
or U8266 (N_8266,N_7950,N_7967);
nor U8267 (N_8267,N_7964,N_7644);
nor U8268 (N_8268,N_7984,N_7834);
and U8269 (N_8269,N_7566,N_7757);
nor U8270 (N_8270,N_7714,N_7609);
nor U8271 (N_8271,N_7947,N_7959);
nand U8272 (N_8272,N_7586,N_7872);
nand U8273 (N_8273,N_7718,N_7613);
and U8274 (N_8274,N_7791,N_7939);
and U8275 (N_8275,N_7583,N_7715);
xor U8276 (N_8276,N_7934,N_7861);
xnor U8277 (N_8277,N_7849,N_7754);
and U8278 (N_8278,N_7965,N_7836);
nor U8279 (N_8279,N_7517,N_7941);
xnor U8280 (N_8280,N_7598,N_7655);
xor U8281 (N_8281,N_7900,N_7678);
nand U8282 (N_8282,N_7543,N_7973);
or U8283 (N_8283,N_7959,N_7776);
xor U8284 (N_8284,N_7628,N_7843);
nand U8285 (N_8285,N_7757,N_7643);
and U8286 (N_8286,N_7611,N_7534);
and U8287 (N_8287,N_7864,N_7544);
xnor U8288 (N_8288,N_7838,N_7973);
nand U8289 (N_8289,N_7688,N_7781);
nand U8290 (N_8290,N_7983,N_7659);
nor U8291 (N_8291,N_7708,N_7769);
or U8292 (N_8292,N_7934,N_7896);
xor U8293 (N_8293,N_7912,N_7842);
nor U8294 (N_8294,N_7854,N_7859);
xnor U8295 (N_8295,N_7656,N_7957);
and U8296 (N_8296,N_7561,N_7575);
or U8297 (N_8297,N_7654,N_7849);
and U8298 (N_8298,N_7793,N_7907);
nand U8299 (N_8299,N_7861,N_7577);
and U8300 (N_8300,N_7507,N_7964);
and U8301 (N_8301,N_7893,N_7545);
and U8302 (N_8302,N_7808,N_7899);
nand U8303 (N_8303,N_7698,N_7652);
or U8304 (N_8304,N_7686,N_7566);
or U8305 (N_8305,N_7984,N_7694);
nand U8306 (N_8306,N_7617,N_7758);
and U8307 (N_8307,N_7579,N_7850);
and U8308 (N_8308,N_7560,N_7605);
xnor U8309 (N_8309,N_7769,N_7681);
and U8310 (N_8310,N_7815,N_7664);
and U8311 (N_8311,N_7515,N_7992);
nor U8312 (N_8312,N_7605,N_7969);
or U8313 (N_8313,N_7838,N_7952);
and U8314 (N_8314,N_7850,N_7512);
nor U8315 (N_8315,N_7541,N_7902);
xnor U8316 (N_8316,N_7626,N_7886);
or U8317 (N_8317,N_7998,N_7621);
xor U8318 (N_8318,N_7938,N_7654);
xnor U8319 (N_8319,N_7671,N_7726);
nand U8320 (N_8320,N_7891,N_7664);
xor U8321 (N_8321,N_7924,N_7993);
xnor U8322 (N_8322,N_7619,N_7504);
xor U8323 (N_8323,N_7874,N_7727);
xnor U8324 (N_8324,N_7889,N_7947);
or U8325 (N_8325,N_7788,N_7654);
nor U8326 (N_8326,N_7759,N_7850);
and U8327 (N_8327,N_7684,N_7903);
nor U8328 (N_8328,N_7976,N_7503);
xor U8329 (N_8329,N_7649,N_7705);
xor U8330 (N_8330,N_7757,N_7854);
nor U8331 (N_8331,N_7813,N_7855);
or U8332 (N_8332,N_7647,N_7986);
and U8333 (N_8333,N_7504,N_7875);
nor U8334 (N_8334,N_7605,N_7895);
or U8335 (N_8335,N_7556,N_7753);
and U8336 (N_8336,N_7647,N_7558);
xnor U8337 (N_8337,N_7796,N_7931);
or U8338 (N_8338,N_7998,N_7568);
nor U8339 (N_8339,N_7753,N_7637);
or U8340 (N_8340,N_7876,N_7525);
or U8341 (N_8341,N_7800,N_7605);
xnor U8342 (N_8342,N_7802,N_7962);
nand U8343 (N_8343,N_7572,N_7549);
and U8344 (N_8344,N_7710,N_7658);
nand U8345 (N_8345,N_7723,N_7696);
xnor U8346 (N_8346,N_7943,N_7683);
or U8347 (N_8347,N_7994,N_7693);
nor U8348 (N_8348,N_7876,N_7568);
and U8349 (N_8349,N_7736,N_7599);
or U8350 (N_8350,N_7843,N_7571);
nand U8351 (N_8351,N_7777,N_7864);
nand U8352 (N_8352,N_7765,N_7924);
and U8353 (N_8353,N_7827,N_7630);
and U8354 (N_8354,N_7733,N_7977);
xnor U8355 (N_8355,N_7944,N_7695);
and U8356 (N_8356,N_7721,N_7852);
nand U8357 (N_8357,N_7907,N_7640);
nor U8358 (N_8358,N_7996,N_7985);
nand U8359 (N_8359,N_7779,N_7982);
nand U8360 (N_8360,N_7980,N_7940);
and U8361 (N_8361,N_7642,N_7695);
or U8362 (N_8362,N_7984,N_7956);
nand U8363 (N_8363,N_7569,N_7681);
or U8364 (N_8364,N_7860,N_7868);
nand U8365 (N_8365,N_7982,N_7927);
or U8366 (N_8366,N_7759,N_7564);
and U8367 (N_8367,N_7572,N_7979);
nand U8368 (N_8368,N_7530,N_7741);
nand U8369 (N_8369,N_7698,N_7829);
or U8370 (N_8370,N_7842,N_7881);
xnor U8371 (N_8371,N_7611,N_7748);
nand U8372 (N_8372,N_7994,N_7533);
nand U8373 (N_8373,N_7970,N_7542);
nor U8374 (N_8374,N_7841,N_7726);
nand U8375 (N_8375,N_7994,N_7687);
xnor U8376 (N_8376,N_7626,N_7599);
nand U8377 (N_8377,N_7686,N_7621);
and U8378 (N_8378,N_7590,N_7865);
nor U8379 (N_8379,N_7702,N_7915);
nand U8380 (N_8380,N_7873,N_7538);
nor U8381 (N_8381,N_7696,N_7978);
nand U8382 (N_8382,N_7648,N_7785);
nor U8383 (N_8383,N_7568,N_7719);
xnor U8384 (N_8384,N_7848,N_7599);
nand U8385 (N_8385,N_7600,N_7763);
xor U8386 (N_8386,N_7811,N_7849);
nand U8387 (N_8387,N_7941,N_7557);
nor U8388 (N_8388,N_7982,N_7730);
or U8389 (N_8389,N_7566,N_7658);
and U8390 (N_8390,N_7974,N_7736);
or U8391 (N_8391,N_7729,N_7763);
or U8392 (N_8392,N_7858,N_7506);
xor U8393 (N_8393,N_7633,N_7788);
nor U8394 (N_8394,N_7875,N_7577);
nor U8395 (N_8395,N_7703,N_7915);
xor U8396 (N_8396,N_7766,N_7925);
or U8397 (N_8397,N_7887,N_7807);
xnor U8398 (N_8398,N_7707,N_7935);
and U8399 (N_8399,N_7632,N_7603);
xnor U8400 (N_8400,N_7886,N_7521);
xnor U8401 (N_8401,N_7946,N_7716);
and U8402 (N_8402,N_7948,N_7546);
and U8403 (N_8403,N_7812,N_7775);
and U8404 (N_8404,N_7518,N_7813);
xnor U8405 (N_8405,N_7522,N_7998);
or U8406 (N_8406,N_7722,N_7607);
or U8407 (N_8407,N_7663,N_7622);
or U8408 (N_8408,N_7605,N_7950);
or U8409 (N_8409,N_7909,N_7834);
and U8410 (N_8410,N_7902,N_7737);
xnor U8411 (N_8411,N_7830,N_7868);
nand U8412 (N_8412,N_7804,N_7705);
xor U8413 (N_8413,N_7564,N_7561);
nand U8414 (N_8414,N_7545,N_7943);
and U8415 (N_8415,N_7588,N_7914);
or U8416 (N_8416,N_7547,N_7789);
or U8417 (N_8417,N_7659,N_7973);
and U8418 (N_8418,N_7987,N_7833);
nand U8419 (N_8419,N_7615,N_7556);
nand U8420 (N_8420,N_7644,N_7565);
nand U8421 (N_8421,N_7991,N_7911);
nor U8422 (N_8422,N_7899,N_7654);
and U8423 (N_8423,N_7918,N_7847);
or U8424 (N_8424,N_7663,N_7528);
xnor U8425 (N_8425,N_7999,N_7730);
or U8426 (N_8426,N_7751,N_7650);
xor U8427 (N_8427,N_7521,N_7508);
and U8428 (N_8428,N_7545,N_7629);
nand U8429 (N_8429,N_7568,N_7926);
and U8430 (N_8430,N_7537,N_7643);
xor U8431 (N_8431,N_7580,N_7770);
and U8432 (N_8432,N_7932,N_7528);
xnor U8433 (N_8433,N_7604,N_7516);
nor U8434 (N_8434,N_7853,N_7811);
or U8435 (N_8435,N_7982,N_7585);
xnor U8436 (N_8436,N_7912,N_7977);
and U8437 (N_8437,N_7520,N_7858);
or U8438 (N_8438,N_7993,N_7698);
xnor U8439 (N_8439,N_7719,N_7726);
xor U8440 (N_8440,N_7850,N_7950);
and U8441 (N_8441,N_7867,N_7542);
nand U8442 (N_8442,N_7867,N_7773);
xnor U8443 (N_8443,N_7686,N_7536);
and U8444 (N_8444,N_7712,N_7892);
or U8445 (N_8445,N_7647,N_7552);
nor U8446 (N_8446,N_7883,N_7900);
nor U8447 (N_8447,N_7796,N_7932);
xor U8448 (N_8448,N_7742,N_7532);
xor U8449 (N_8449,N_7555,N_7841);
xnor U8450 (N_8450,N_7519,N_7954);
or U8451 (N_8451,N_7918,N_7549);
or U8452 (N_8452,N_7576,N_7693);
xor U8453 (N_8453,N_7520,N_7677);
nor U8454 (N_8454,N_7615,N_7899);
and U8455 (N_8455,N_7868,N_7942);
xor U8456 (N_8456,N_7516,N_7767);
nand U8457 (N_8457,N_7847,N_7856);
nor U8458 (N_8458,N_7632,N_7924);
and U8459 (N_8459,N_7532,N_7608);
nor U8460 (N_8460,N_7848,N_7845);
and U8461 (N_8461,N_7506,N_7975);
and U8462 (N_8462,N_7943,N_7840);
nand U8463 (N_8463,N_7660,N_7832);
or U8464 (N_8464,N_7532,N_7511);
nor U8465 (N_8465,N_7782,N_7911);
and U8466 (N_8466,N_7994,N_7769);
xor U8467 (N_8467,N_7617,N_7688);
nand U8468 (N_8468,N_7987,N_7508);
nand U8469 (N_8469,N_7931,N_7619);
nand U8470 (N_8470,N_7544,N_7988);
nand U8471 (N_8471,N_7524,N_7926);
or U8472 (N_8472,N_7830,N_7637);
and U8473 (N_8473,N_7637,N_7654);
and U8474 (N_8474,N_7641,N_7642);
and U8475 (N_8475,N_7533,N_7841);
and U8476 (N_8476,N_7673,N_7519);
nand U8477 (N_8477,N_7779,N_7759);
nor U8478 (N_8478,N_7881,N_7846);
or U8479 (N_8479,N_7727,N_7671);
or U8480 (N_8480,N_7930,N_7747);
and U8481 (N_8481,N_7965,N_7738);
nand U8482 (N_8482,N_7790,N_7789);
nand U8483 (N_8483,N_7856,N_7678);
or U8484 (N_8484,N_7654,N_7962);
or U8485 (N_8485,N_7665,N_7659);
nor U8486 (N_8486,N_7851,N_7612);
xnor U8487 (N_8487,N_7577,N_7592);
or U8488 (N_8488,N_7530,N_7938);
nor U8489 (N_8489,N_7591,N_7656);
nand U8490 (N_8490,N_7820,N_7843);
nor U8491 (N_8491,N_7691,N_7983);
nand U8492 (N_8492,N_7660,N_7643);
nand U8493 (N_8493,N_7950,N_7785);
xor U8494 (N_8494,N_7911,N_7724);
or U8495 (N_8495,N_7679,N_7685);
and U8496 (N_8496,N_7694,N_7768);
xor U8497 (N_8497,N_7533,N_7706);
nor U8498 (N_8498,N_7851,N_7927);
nor U8499 (N_8499,N_7905,N_7594);
xor U8500 (N_8500,N_8343,N_8428);
or U8501 (N_8501,N_8149,N_8277);
or U8502 (N_8502,N_8010,N_8132);
and U8503 (N_8503,N_8136,N_8247);
nor U8504 (N_8504,N_8098,N_8158);
xnor U8505 (N_8505,N_8028,N_8274);
or U8506 (N_8506,N_8232,N_8363);
nor U8507 (N_8507,N_8006,N_8401);
or U8508 (N_8508,N_8390,N_8154);
xnor U8509 (N_8509,N_8494,N_8474);
nor U8510 (N_8510,N_8359,N_8301);
nand U8511 (N_8511,N_8042,N_8325);
and U8512 (N_8512,N_8252,N_8241);
xnor U8513 (N_8513,N_8074,N_8330);
or U8514 (N_8514,N_8342,N_8203);
and U8515 (N_8515,N_8016,N_8129);
nand U8516 (N_8516,N_8271,N_8285);
nor U8517 (N_8517,N_8444,N_8372);
and U8518 (N_8518,N_8204,N_8397);
nor U8519 (N_8519,N_8472,N_8282);
nor U8520 (N_8520,N_8346,N_8105);
xnor U8521 (N_8521,N_8115,N_8059);
nor U8522 (N_8522,N_8293,N_8226);
or U8523 (N_8523,N_8446,N_8067);
nand U8524 (N_8524,N_8045,N_8322);
nand U8525 (N_8525,N_8462,N_8395);
and U8526 (N_8526,N_8255,N_8114);
nor U8527 (N_8527,N_8174,N_8200);
nand U8528 (N_8528,N_8066,N_8336);
nor U8529 (N_8529,N_8235,N_8469);
nand U8530 (N_8530,N_8213,N_8464);
xor U8531 (N_8531,N_8141,N_8003);
or U8532 (N_8532,N_8254,N_8097);
nand U8533 (N_8533,N_8032,N_8036);
or U8534 (N_8534,N_8058,N_8447);
or U8535 (N_8535,N_8170,N_8125);
nand U8536 (N_8536,N_8075,N_8092);
or U8537 (N_8537,N_8086,N_8374);
nand U8538 (N_8538,N_8048,N_8224);
nand U8539 (N_8539,N_8157,N_8454);
xor U8540 (N_8540,N_8068,N_8439);
xor U8541 (N_8541,N_8261,N_8292);
nor U8542 (N_8542,N_8205,N_8162);
nand U8543 (N_8543,N_8055,N_8117);
or U8544 (N_8544,N_8485,N_8169);
nor U8545 (N_8545,N_8243,N_8187);
nand U8546 (N_8546,N_8240,N_8137);
or U8547 (N_8547,N_8034,N_8366);
nand U8548 (N_8548,N_8418,N_8423);
nand U8549 (N_8549,N_8442,N_8465);
nand U8550 (N_8550,N_8451,N_8477);
and U8551 (N_8551,N_8297,N_8202);
and U8552 (N_8552,N_8100,N_8299);
and U8553 (N_8553,N_8345,N_8371);
nand U8554 (N_8554,N_8014,N_8287);
and U8555 (N_8555,N_8049,N_8410);
nor U8556 (N_8556,N_8278,N_8393);
or U8557 (N_8557,N_8121,N_8361);
nand U8558 (N_8558,N_8031,N_8217);
xnor U8559 (N_8559,N_8171,N_8238);
xnor U8560 (N_8560,N_8239,N_8193);
nor U8561 (N_8561,N_8425,N_8348);
or U8562 (N_8562,N_8470,N_8272);
xor U8563 (N_8563,N_8267,N_8269);
and U8564 (N_8564,N_8402,N_8142);
and U8565 (N_8565,N_8176,N_8384);
or U8566 (N_8566,N_8147,N_8107);
nor U8567 (N_8567,N_8391,N_8248);
or U8568 (N_8568,N_8093,N_8113);
nand U8569 (N_8569,N_8222,N_8072);
nor U8570 (N_8570,N_8354,N_8103);
xnor U8571 (N_8571,N_8030,N_8087);
or U8572 (N_8572,N_8094,N_8168);
or U8573 (N_8573,N_8318,N_8284);
nor U8574 (N_8574,N_8473,N_8122);
nand U8575 (N_8575,N_8190,N_8064);
nor U8576 (N_8576,N_8436,N_8090);
nand U8577 (N_8577,N_8275,N_8338);
xnor U8578 (N_8578,N_8327,N_8483);
or U8579 (N_8579,N_8134,N_8478);
or U8580 (N_8580,N_8312,N_8151);
or U8581 (N_8581,N_8073,N_8091);
nand U8582 (N_8582,N_8022,N_8166);
and U8583 (N_8583,N_8258,N_8381);
or U8584 (N_8584,N_8047,N_8373);
or U8585 (N_8585,N_8298,N_8025);
xnor U8586 (N_8586,N_8419,N_8110);
nand U8587 (N_8587,N_8427,N_8043);
and U8588 (N_8588,N_8340,N_8289);
and U8589 (N_8589,N_8279,N_8368);
and U8590 (N_8590,N_8400,N_8405);
or U8591 (N_8591,N_8482,N_8357);
nand U8592 (N_8592,N_8146,N_8159);
nor U8593 (N_8593,N_8233,N_8367);
nand U8594 (N_8594,N_8455,N_8286);
and U8595 (N_8595,N_8399,N_8040);
or U8596 (N_8596,N_8290,N_8440);
xor U8597 (N_8597,N_8228,N_8013);
and U8598 (N_8598,N_8294,N_8063);
nand U8599 (N_8599,N_8457,N_8347);
or U8600 (N_8600,N_8076,N_8081);
nand U8601 (N_8601,N_8452,N_8080);
and U8602 (N_8602,N_8408,N_8054);
xnor U8603 (N_8603,N_8186,N_8430);
and U8604 (N_8604,N_8128,N_8253);
nor U8605 (N_8605,N_8172,N_8488);
or U8606 (N_8606,N_8281,N_8356);
xor U8607 (N_8607,N_8331,N_8265);
nor U8608 (N_8608,N_8362,N_8260);
nor U8609 (N_8609,N_8018,N_8460);
nor U8610 (N_8610,N_8225,N_8029);
nand U8611 (N_8611,N_8424,N_8388);
and U8612 (N_8612,N_8387,N_8386);
nand U8613 (N_8613,N_8484,N_8314);
and U8614 (N_8614,N_8406,N_8050);
nand U8615 (N_8615,N_8037,N_8421);
or U8616 (N_8616,N_8223,N_8270);
xor U8617 (N_8617,N_8459,N_8324);
nand U8618 (N_8618,N_8052,N_8433);
and U8619 (N_8619,N_8351,N_8078);
or U8620 (N_8620,N_8138,N_8127);
or U8621 (N_8621,N_8104,N_8133);
or U8622 (N_8622,N_8001,N_8412);
xor U8623 (N_8623,N_8320,N_8209);
xnor U8624 (N_8624,N_8481,N_8116);
nor U8625 (N_8625,N_8178,N_8046);
and U8626 (N_8626,N_8341,N_8216);
or U8627 (N_8627,N_8196,N_8065);
nor U8628 (N_8628,N_8414,N_8246);
nor U8629 (N_8629,N_8041,N_8008);
and U8630 (N_8630,N_8135,N_8335);
nand U8631 (N_8631,N_8389,N_8139);
nor U8632 (N_8632,N_8156,N_8329);
nor U8633 (N_8633,N_8112,N_8438);
and U8634 (N_8634,N_8012,N_8199);
xor U8635 (N_8635,N_8244,N_8208);
or U8636 (N_8636,N_8140,N_8323);
nand U8637 (N_8637,N_8120,N_8291);
or U8638 (N_8638,N_8130,N_8349);
and U8639 (N_8639,N_8417,N_8035);
nor U8640 (N_8640,N_8307,N_8015);
xor U8641 (N_8641,N_8475,N_8449);
or U8642 (N_8642,N_8355,N_8360);
or U8643 (N_8643,N_8060,N_8306);
nand U8644 (N_8644,N_8334,N_8227);
or U8645 (N_8645,N_8313,N_8242);
and U8646 (N_8646,N_8358,N_8184);
and U8647 (N_8647,N_8163,N_8005);
or U8648 (N_8648,N_8420,N_8353);
nand U8649 (N_8649,N_8300,N_8394);
xor U8650 (N_8650,N_8328,N_8434);
nand U8651 (N_8651,N_8332,N_8195);
nor U8652 (N_8652,N_8053,N_8165);
xnor U8653 (N_8653,N_8296,N_8411);
nor U8654 (N_8654,N_8375,N_8221);
or U8655 (N_8655,N_8020,N_8364);
nor U8656 (N_8656,N_8079,N_8422);
or U8657 (N_8657,N_8497,N_8144);
and U8658 (N_8658,N_8085,N_8118);
and U8659 (N_8659,N_8183,N_8276);
nor U8660 (N_8660,N_8370,N_8480);
nand U8661 (N_8661,N_8326,N_8038);
nor U8662 (N_8662,N_8153,N_8378);
nand U8663 (N_8663,N_8316,N_8295);
and U8664 (N_8664,N_8007,N_8061);
xnor U8665 (N_8665,N_8099,N_8197);
xnor U8666 (N_8666,N_8167,N_8229);
nand U8667 (N_8667,N_8317,N_8493);
nand U8668 (N_8668,N_8207,N_8131);
and U8669 (N_8669,N_8148,N_8056);
nand U8670 (N_8670,N_8160,N_8017);
nor U8671 (N_8671,N_8413,N_8185);
xor U8672 (N_8672,N_8376,N_8264);
xor U8673 (N_8673,N_8311,N_8304);
nor U8674 (N_8674,N_8212,N_8182);
xnor U8675 (N_8675,N_8069,N_8237);
nor U8676 (N_8676,N_8453,N_8051);
and U8677 (N_8677,N_8380,N_8004);
or U8678 (N_8678,N_8206,N_8344);
and U8679 (N_8679,N_8429,N_8407);
xnor U8680 (N_8680,N_8310,N_8441);
nand U8681 (N_8681,N_8431,N_8234);
or U8682 (N_8682,N_8396,N_8236);
nand U8683 (N_8683,N_8435,N_8152);
xor U8684 (N_8684,N_8445,N_8188);
or U8685 (N_8685,N_8309,N_8218);
nand U8686 (N_8686,N_8467,N_8259);
or U8687 (N_8687,N_8403,N_8077);
and U8688 (N_8688,N_8230,N_8256);
and U8689 (N_8689,N_8011,N_8164);
and U8690 (N_8690,N_8303,N_8145);
xor U8691 (N_8691,N_8492,N_8491);
and U8692 (N_8692,N_8095,N_8432);
nor U8693 (N_8693,N_8249,N_8487);
xnor U8694 (N_8694,N_8339,N_8161);
or U8695 (N_8695,N_8398,N_8215);
xnor U8696 (N_8696,N_8479,N_8201);
nand U8697 (N_8697,N_8211,N_8471);
xor U8698 (N_8698,N_8179,N_8251);
nor U8699 (N_8699,N_8083,N_8124);
or U8700 (N_8700,N_8392,N_8245);
or U8701 (N_8701,N_8415,N_8119);
and U8702 (N_8702,N_8071,N_8111);
xnor U8703 (N_8703,N_8257,N_8385);
nand U8704 (N_8704,N_8173,N_8021);
nor U8705 (N_8705,N_8437,N_8382);
or U8706 (N_8706,N_8194,N_8023);
nand U8707 (N_8707,N_8365,N_8499);
or U8708 (N_8708,N_8192,N_8191);
and U8709 (N_8709,N_8369,N_8250);
or U8710 (N_8710,N_8321,N_8495);
and U8711 (N_8711,N_8490,N_8333);
nand U8712 (N_8712,N_8024,N_8057);
or U8713 (N_8713,N_8143,N_8352);
and U8714 (N_8714,N_8379,N_8096);
nor U8715 (N_8715,N_8283,N_8476);
and U8716 (N_8716,N_8000,N_8033);
and U8717 (N_8717,N_8102,N_8126);
xor U8718 (N_8718,N_8443,N_8315);
xnor U8719 (N_8719,N_8288,N_8039);
nand U8720 (N_8720,N_8019,N_8109);
or U8721 (N_8721,N_8280,N_8404);
xor U8722 (N_8722,N_8155,N_8266);
nor U8723 (N_8723,N_8496,N_8489);
xor U8724 (N_8724,N_8319,N_8498);
or U8725 (N_8725,N_8044,N_8108);
or U8726 (N_8726,N_8210,N_8377);
and U8727 (N_8727,N_8273,N_8177);
and U8728 (N_8728,N_8305,N_8101);
nor U8729 (N_8729,N_8070,N_8219);
nand U8730 (N_8730,N_8231,N_8062);
or U8731 (N_8731,N_8383,N_8486);
and U8732 (N_8732,N_8089,N_8106);
and U8733 (N_8733,N_8268,N_8263);
nor U8734 (N_8734,N_8198,N_8468);
nor U8735 (N_8735,N_8082,N_8466);
and U8736 (N_8736,N_8409,N_8175);
nand U8737 (N_8737,N_8002,N_8262);
xor U8738 (N_8738,N_8084,N_8426);
nand U8739 (N_8739,N_8026,N_8337);
and U8740 (N_8740,N_8180,N_8150);
nor U8741 (N_8741,N_8302,N_8456);
nand U8742 (N_8742,N_8027,N_8448);
xnor U8743 (N_8743,N_8458,N_8416);
nor U8744 (N_8744,N_8214,N_8308);
nand U8745 (N_8745,N_8463,N_8450);
nand U8746 (N_8746,N_8461,N_8181);
xnor U8747 (N_8747,N_8189,N_8220);
xnor U8748 (N_8748,N_8350,N_8123);
nand U8749 (N_8749,N_8088,N_8009);
nand U8750 (N_8750,N_8490,N_8160);
nand U8751 (N_8751,N_8284,N_8184);
nor U8752 (N_8752,N_8181,N_8409);
or U8753 (N_8753,N_8106,N_8379);
nor U8754 (N_8754,N_8426,N_8281);
and U8755 (N_8755,N_8014,N_8383);
nand U8756 (N_8756,N_8012,N_8096);
and U8757 (N_8757,N_8271,N_8092);
or U8758 (N_8758,N_8478,N_8179);
nor U8759 (N_8759,N_8372,N_8352);
and U8760 (N_8760,N_8081,N_8010);
nor U8761 (N_8761,N_8153,N_8054);
and U8762 (N_8762,N_8186,N_8479);
xnor U8763 (N_8763,N_8316,N_8081);
or U8764 (N_8764,N_8061,N_8090);
nor U8765 (N_8765,N_8287,N_8025);
and U8766 (N_8766,N_8313,N_8081);
and U8767 (N_8767,N_8016,N_8195);
or U8768 (N_8768,N_8127,N_8293);
xor U8769 (N_8769,N_8487,N_8453);
nor U8770 (N_8770,N_8367,N_8035);
or U8771 (N_8771,N_8009,N_8309);
or U8772 (N_8772,N_8139,N_8094);
and U8773 (N_8773,N_8415,N_8407);
xor U8774 (N_8774,N_8012,N_8008);
nor U8775 (N_8775,N_8100,N_8233);
or U8776 (N_8776,N_8248,N_8179);
nor U8777 (N_8777,N_8396,N_8382);
nor U8778 (N_8778,N_8406,N_8156);
or U8779 (N_8779,N_8097,N_8141);
xor U8780 (N_8780,N_8461,N_8078);
or U8781 (N_8781,N_8398,N_8063);
or U8782 (N_8782,N_8073,N_8064);
and U8783 (N_8783,N_8400,N_8382);
nor U8784 (N_8784,N_8050,N_8201);
and U8785 (N_8785,N_8489,N_8110);
xor U8786 (N_8786,N_8005,N_8057);
xor U8787 (N_8787,N_8427,N_8316);
and U8788 (N_8788,N_8022,N_8478);
nor U8789 (N_8789,N_8192,N_8099);
xor U8790 (N_8790,N_8468,N_8462);
xor U8791 (N_8791,N_8165,N_8458);
and U8792 (N_8792,N_8475,N_8313);
nor U8793 (N_8793,N_8026,N_8192);
xor U8794 (N_8794,N_8376,N_8155);
and U8795 (N_8795,N_8019,N_8394);
or U8796 (N_8796,N_8139,N_8317);
nand U8797 (N_8797,N_8205,N_8426);
nand U8798 (N_8798,N_8111,N_8322);
nor U8799 (N_8799,N_8195,N_8234);
nor U8800 (N_8800,N_8495,N_8397);
and U8801 (N_8801,N_8152,N_8021);
xor U8802 (N_8802,N_8182,N_8368);
and U8803 (N_8803,N_8029,N_8396);
and U8804 (N_8804,N_8364,N_8203);
xor U8805 (N_8805,N_8408,N_8412);
and U8806 (N_8806,N_8059,N_8076);
nand U8807 (N_8807,N_8394,N_8059);
or U8808 (N_8808,N_8105,N_8430);
or U8809 (N_8809,N_8463,N_8384);
nand U8810 (N_8810,N_8294,N_8021);
and U8811 (N_8811,N_8415,N_8173);
and U8812 (N_8812,N_8368,N_8180);
and U8813 (N_8813,N_8280,N_8065);
and U8814 (N_8814,N_8369,N_8168);
nand U8815 (N_8815,N_8215,N_8011);
nor U8816 (N_8816,N_8068,N_8038);
nor U8817 (N_8817,N_8251,N_8002);
or U8818 (N_8818,N_8351,N_8365);
or U8819 (N_8819,N_8332,N_8216);
nor U8820 (N_8820,N_8126,N_8281);
nor U8821 (N_8821,N_8154,N_8385);
and U8822 (N_8822,N_8313,N_8169);
nor U8823 (N_8823,N_8133,N_8008);
xor U8824 (N_8824,N_8065,N_8146);
nor U8825 (N_8825,N_8262,N_8125);
and U8826 (N_8826,N_8409,N_8111);
nand U8827 (N_8827,N_8469,N_8203);
or U8828 (N_8828,N_8035,N_8349);
nand U8829 (N_8829,N_8298,N_8390);
nor U8830 (N_8830,N_8274,N_8259);
nand U8831 (N_8831,N_8251,N_8278);
nand U8832 (N_8832,N_8131,N_8459);
nand U8833 (N_8833,N_8213,N_8408);
nor U8834 (N_8834,N_8142,N_8087);
and U8835 (N_8835,N_8237,N_8103);
and U8836 (N_8836,N_8378,N_8425);
and U8837 (N_8837,N_8435,N_8388);
nor U8838 (N_8838,N_8416,N_8283);
nor U8839 (N_8839,N_8304,N_8366);
xnor U8840 (N_8840,N_8463,N_8169);
and U8841 (N_8841,N_8172,N_8355);
or U8842 (N_8842,N_8325,N_8287);
xor U8843 (N_8843,N_8189,N_8437);
nand U8844 (N_8844,N_8331,N_8197);
xor U8845 (N_8845,N_8133,N_8129);
nand U8846 (N_8846,N_8360,N_8151);
nand U8847 (N_8847,N_8406,N_8329);
xor U8848 (N_8848,N_8471,N_8420);
nor U8849 (N_8849,N_8466,N_8288);
nor U8850 (N_8850,N_8013,N_8059);
nor U8851 (N_8851,N_8041,N_8113);
or U8852 (N_8852,N_8083,N_8397);
nor U8853 (N_8853,N_8111,N_8335);
nand U8854 (N_8854,N_8012,N_8250);
and U8855 (N_8855,N_8327,N_8152);
xnor U8856 (N_8856,N_8282,N_8367);
xnor U8857 (N_8857,N_8313,N_8080);
and U8858 (N_8858,N_8351,N_8172);
or U8859 (N_8859,N_8362,N_8047);
nand U8860 (N_8860,N_8111,N_8374);
nand U8861 (N_8861,N_8034,N_8398);
or U8862 (N_8862,N_8229,N_8063);
and U8863 (N_8863,N_8406,N_8319);
nand U8864 (N_8864,N_8264,N_8092);
and U8865 (N_8865,N_8275,N_8317);
nand U8866 (N_8866,N_8214,N_8309);
nand U8867 (N_8867,N_8357,N_8164);
or U8868 (N_8868,N_8054,N_8078);
nand U8869 (N_8869,N_8187,N_8396);
and U8870 (N_8870,N_8109,N_8489);
nand U8871 (N_8871,N_8114,N_8116);
and U8872 (N_8872,N_8163,N_8058);
and U8873 (N_8873,N_8490,N_8195);
nor U8874 (N_8874,N_8168,N_8054);
and U8875 (N_8875,N_8471,N_8007);
nand U8876 (N_8876,N_8032,N_8267);
and U8877 (N_8877,N_8440,N_8102);
xor U8878 (N_8878,N_8435,N_8493);
nand U8879 (N_8879,N_8189,N_8112);
nand U8880 (N_8880,N_8407,N_8089);
or U8881 (N_8881,N_8116,N_8227);
nor U8882 (N_8882,N_8249,N_8406);
xor U8883 (N_8883,N_8346,N_8198);
nand U8884 (N_8884,N_8324,N_8478);
nand U8885 (N_8885,N_8415,N_8141);
nand U8886 (N_8886,N_8303,N_8267);
nand U8887 (N_8887,N_8341,N_8104);
or U8888 (N_8888,N_8492,N_8054);
nand U8889 (N_8889,N_8042,N_8262);
nor U8890 (N_8890,N_8482,N_8465);
and U8891 (N_8891,N_8253,N_8308);
nand U8892 (N_8892,N_8374,N_8345);
or U8893 (N_8893,N_8450,N_8268);
nand U8894 (N_8894,N_8098,N_8345);
nand U8895 (N_8895,N_8066,N_8047);
or U8896 (N_8896,N_8377,N_8493);
and U8897 (N_8897,N_8082,N_8275);
or U8898 (N_8898,N_8024,N_8039);
and U8899 (N_8899,N_8353,N_8342);
xnor U8900 (N_8900,N_8207,N_8115);
nor U8901 (N_8901,N_8328,N_8197);
nand U8902 (N_8902,N_8026,N_8395);
and U8903 (N_8903,N_8129,N_8479);
or U8904 (N_8904,N_8431,N_8185);
nand U8905 (N_8905,N_8127,N_8371);
or U8906 (N_8906,N_8436,N_8346);
xnor U8907 (N_8907,N_8181,N_8447);
xor U8908 (N_8908,N_8428,N_8275);
nor U8909 (N_8909,N_8403,N_8456);
nor U8910 (N_8910,N_8444,N_8024);
nor U8911 (N_8911,N_8460,N_8228);
nor U8912 (N_8912,N_8226,N_8062);
or U8913 (N_8913,N_8359,N_8383);
or U8914 (N_8914,N_8168,N_8073);
xnor U8915 (N_8915,N_8254,N_8430);
xnor U8916 (N_8916,N_8381,N_8499);
nand U8917 (N_8917,N_8169,N_8228);
or U8918 (N_8918,N_8018,N_8480);
or U8919 (N_8919,N_8378,N_8260);
nand U8920 (N_8920,N_8188,N_8069);
nand U8921 (N_8921,N_8369,N_8458);
nand U8922 (N_8922,N_8092,N_8246);
xnor U8923 (N_8923,N_8062,N_8366);
or U8924 (N_8924,N_8092,N_8398);
xnor U8925 (N_8925,N_8072,N_8357);
or U8926 (N_8926,N_8383,N_8470);
and U8927 (N_8927,N_8143,N_8378);
nand U8928 (N_8928,N_8379,N_8196);
nand U8929 (N_8929,N_8433,N_8419);
nor U8930 (N_8930,N_8141,N_8204);
and U8931 (N_8931,N_8211,N_8107);
nor U8932 (N_8932,N_8034,N_8428);
nor U8933 (N_8933,N_8268,N_8322);
xor U8934 (N_8934,N_8003,N_8317);
nor U8935 (N_8935,N_8268,N_8038);
and U8936 (N_8936,N_8067,N_8097);
nor U8937 (N_8937,N_8148,N_8223);
nor U8938 (N_8938,N_8087,N_8192);
and U8939 (N_8939,N_8064,N_8273);
or U8940 (N_8940,N_8479,N_8224);
xnor U8941 (N_8941,N_8409,N_8164);
nor U8942 (N_8942,N_8456,N_8078);
nand U8943 (N_8943,N_8050,N_8132);
and U8944 (N_8944,N_8114,N_8320);
and U8945 (N_8945,N_8357,N_8494);
or U8946 (N_8946,N_8323,N_8366);
and U8947 (N_8947,N_8205,N_8436);
nand U8948 (N_8948,N_8217,N_8409);
or U8949 (N_8949,N_8004,N_8414);
xor U8950 (N_8950,N_8030,N_8343);
nor U8951 (N_8951,N_8127,N_8288);
or U8952 (N_8952,N_8085,N_8365);
or U8953 (N_8953,N_8133,N_8335);
xnor U8954 (N_8954,N_8160,N_8031);
and U8955 (N_8955,N_8187,N_8130);
xor U8956 (N_8956,N_8090,N_8104);
xor U8957 (N_8957,N_8350,N_8140);
or U8958 (N_8958,N_8334,N_8068);
nor U8959 (N_8959,N_8336,N_8235);
nand U8960 (N_8960,N_8287,N_8257);
and U8961 (N_8961,N_8142,N_8483);
xor U8962 (N_8962,N_8360,N_8378);
nor U8963 (N_8963,N_8314,N_8434);
or U8964 (N_8964,N_8453,N_8305);
nand U8965 (N_8965,N_8047,N_8065);
nand U8966 (N_8966,N_8374,N_8003);
nor U8967 (N_8967,N_8144,N_8270);
nor U8968 (N_8968,N_8107,N_8094);
xor U8969 (N_8969,N_8254,N_8135);
nand U8970 (N_8970,N_8220,N_8239);
nand U8971 (N_8971,N_8339,N_8336);
or U8972 (N_8972,N_8411,N_8145);
nor U8973 (N_8973,N_8347,N_8352);
xor U8974 (N_8974,N_8214,N_8136);
and U8975 (N_8975,N_8421,N_8316);
nand U8976 (N_8976,N_8466,N_8033);
nand U8977 (N_8977,N_8087,N_8146);
or U8978 (N_8978,N_8265,N_8231);
and U8979 (N_8979,N_8352,N_8049);
nor U8980 (N_8980,N_8276,N_8337);
and U8981 (N_8981,N_8335,N_8417);
nand U8982 (N_8982,N_8492,N_8136);
nand U8983 (N_8983,N_8441,N_8425);
xnor U8984 (N_8984,N_8303,N_8120);
xnor U8985 (N_8985,N_8085,N_8075);
and U8986 (N_8986,N_8182,N_8363);
xnor U8987 (N_8987,N_8259,N_8472);
nand U8988 (N_8988,N_8308,N_8008);
or U8989 (N_8989,N_8384,N_8421);
nor U8990 (N_8990,N_8057,N_8099);
nand U8991 (N_8991,N_8262,N_8336);
and U8992 (N_8992,N_8082,N_8459);
or U8993 (N_8993,N_8430,N_8013);
nand U8994 (N_8994,N_8319,N_8435);
nand U8995 (N_8995,N_8201,N_8376);
nand U8996 (N_8996,N_8254,N_8074);
xnor U8997 (N_8997,N_8036,N_8026);
xnor U8998 (N_8998,N_8409,N_8339);
xor U8999 (N_8999,N_8164,N_8479);
xor U9000 (N_9000,N_8658,N_8963);
nand U9001 (N_9001,N_8836,N_8773);
or U9002 (N_9002,N_8670,N_8810);
nand U9003 (N_9003,N_8664,N_8881);
and U9004 (N_9004,N_8536,N_8555);
xor U9005 (N_9005,N_8705,N_8924);
and U9006 (N_9006,N_8977,N_8807);
nor U9007 (N_9007,N_8790,N_8759);
nor U9008 (N_9008,N_8743,N_8798);
xor U9009 (N_9009,N_8824,N_8776);
nor U9010 (N_9010,N_8579,N_8838);
nand U9011 (N_9011,N_8597,N_8765);
and U9012 (N_9012,N_8632,N_8696);
nor U9013 (N_9013,N_8827,N_8591);
or U9014 (N_9014,N_8746,N_8806);
or U9015 (N_9015,N_8638,N_8882);
xor U9016 (N_9016,N_8805,N_8930);
xor U9017 (N_9017,N_8546,N_8851);
nand U9018 (N_9018,N_8572,N_8926);
and U9019 (N_9019,N_8995,N_8512);
or U9020 (N_9020,N_8648,N_8586);
or U9021 (N_9021,N_8662,N_8989);
or U9022 (N_9022,N_8764,N_8966);
and U9023 (N_9023,N_8745,N_8573);
or U9024 (N_9024,N_8630,N_8869);
nand U9025 (N_9025,N_8792,N_8825);
nand U9026 (N_9026,N_8797,N_8699);
nand U9027 (N_9027,N_8593,N_8858);
and U9028 (N_9028,N_8950,N_8800);
or U9029 (N_9029,N_8668,N_8719);
nand U9030 (N_9030,N_8642,N_8808);
xor U9031 (N_9031,N_8721,N_8679);
xor U9032 (N_9032,N_8657,N_8799);
nand U9033 (N_9033,N_8590,N_8880);
and U9034 (N_9034,N_8636,N_8713);
xnor U9035 (N_9035,N_8617,N_8994);
and U9036 (N_9036,N_8667,N_8785);
or U9037 (N_9037,N_8928,N_8606);
nand U9038 (N_9038,N_8929,N_8643);
nor U9039 (N_9039,N_8535,N_8828);
nand U9040 (N_9040,N_8949,N_8955);
and U9041 (N_9041,N_8871,N_8844);
nand U9042 (N_9042,N_8973,N_8980);
or U9043 (N_9043,N_8526,N_8751);
nor U9044 (N_9044,N_8707,N_8985);
and U9045 (N_9045,N_8716,N_8940);
nand U9046 (N_9046,N_8849,N_8976);
or U9047 (N_9047,N_8616,N_8513);
xnor U9048 (N_9048,N_8506,N_8770);
xnor U9049 (N_9049,N_8523,N_8508);
nand U9050 (N_9050,N_8684,N_8917);
xnor U9051 (N_9051,N_8725,N_8850);
or U9052 (N_9052,N_8631,N_8706);
nor U9053 (N_9053,N_8961,N_8848);
xor U9054 (N_9054,N_8500,N_8704);
and U9055 (N_9055,N_8520,N_8672);
nor U9056 (N_9056,N_8511,N_8974);
or U9057 (N_9057,N_8819,N_8548);
nor U9058 (N_9058,N_8766,N_8567);
nor U9059 (N_9059,N_8558,N_8916);
nor U9060 (N_9060,N_8783,N_8730);
nand U9061 (N_9061,N_8556,N_8525);
nand U9062 (N_9062,N_8644,N_8560);
nor U9063 (N_9063,N_8821,N_8757);
nand U9064 (N_9064,N_8677,N_8912);
xor U9065 (N_9065,N_8964,N_8674);
nand U9066 (N_9066,N_8864,N_8729);
nor U9067 (N_9067,N_8709,N_8522);
nand U9068 (N_9068,N_8996,N_8875);
xor U9069 (N_9069,N_8703,N_8519);
xor U9070 (N_9070,N_8564,N_8602);
nand U9071 (N_9071,N_8660,N_8780);
nor U9072 (N_9072,N_8649,N_8866);
or U9073 (N_9073,N_8641,N_8655);
and U9074 (N_9074,N_8620,N_8507);
xnor U9075 (N_9075,N_8576,N_8829);
nor U9076 (N_9076,N_8942,N_8634);
xor U9077 (N_9077,N_8998,N_8698);
nor U9078 (N_9078,N_8551,N_8767);
and U9079 (N_9079,N_8561,N_8999);
or U9080 (N_9080,N_8943,N_8600);
nand U9081 (N_9081,N_8544,N_8585);
or U9082 (N_9082,N_8900,N_8768);
xnor U9083 (N_9083,N_8531,N_8760);
xor U9084 (N_9084,N_8727,N_8692);
and U9085 (N_9085,N_8865,N_8575);
nand U9086 (N_9086,N_8599,N_8794);
or U9087 (N_9087,N_8610,N_8744);
xnor U9088 (N_9088,N_8505,N_8758);
nor U9089 (N_9089,N_8907,N_8921);
nor U9090 (N_9090,N_8681,N_8565);
nor U9091 (N_9091,N_8893,N_8515);
nor U9092 (N_9092,N_8609,N_8854);
nand U9093 (N_9093,N_8971,N_8659);
xor U9094 (N_9094,N_8663,N_8877);
nand U9095 (N_9095,N_8583,N_8899);
and U9096 (N_9096,N_8802,N_8510);
xor U9097 (N_9097,N_8835,N_8883);
nand U9098 (N_9098,N_8876,N_8504);
nor U9099 (N_9099,N_8922,N_8603);
nand U9100 (N_9100,N_8627,N_8615);
xor U9101 (N_9101,N_8813,N_8733);
nor U9102 (N_9102,N_8629,N_8761);
and U9103 (N_9103,N_8981,N_8958);
and U9104 (N_9104,N_8736,N_8762);
nand U9105 (N_9105,N_8686,N_8997);
and U9106 (N_9106,N_8934,N_8968);
and U9107 (N_9107,N_8749,N_8863);
xor U9108 (N_9108,N_8710,N_8748);
xor U9109 (N_9109,N_8902,N_8771);
xor U9110 (N_9110,N_8534,N_8554);
nand U9111 (N_9111,N_8936,N_8784);
nor U9112 (N_9112,N_8509,N_8817);
nand U9113 (N_9113,N_8624,N_8502);
nor U9114 (N_9114,N_8932,N_8789);
nand U9115 (N_9115,N_8584,N_8847);
nor U9116 (N_9116,N_8781,N_8820);
and U9117 (N_9117,N_8688,N_8656);
nor U9118 (N_9118,N_8991,N_8925);
nand U9119 (N_9119,N_8892,N_8682);
nand U9120 (N_9120,N_8952,N_8803);
nor U9121 (N_9121,N_8661,N_8633);
or U9122 (N_9122,N_8840,N_8984);
or U9123 (N_9123,N_8666,N_8524);
or U9124 (N_9124,N_8589,N_8647);
nor U9125 (N_9125,N_8547,N_8690);
or U9126 (N_9126,N_8793,N_8683);
nand U9127 (N_9127,N_8946,N_8685);
and U9128 (N_9128,N_8975,N_8972);
xor U9129 (N_9129,N_8755,N_8872);
nand U9130 (N_9130,N_8947,N_8532);
nor U9131 (N_9131,N_8853,N_8712);
nor U9132 (N_9132,N_8516,N_8860);
nand U9133 (N_9133,N_8884,N_8954);
nor U9134 (N_9134,N_8697,N_8957);
nand U9135 (N_9135,N_8889,N_8652);
xor U9136 (N_9136,N_8960,N_8528);
or U9137 (N_9137,N_8935,N_8896);
and U9138 (N_9138,N_8846,N_8687);
or U9139 (N_9139,N_8752,N_8607);
or U9140 (N_9140,N_8675,N_8774);
and U9141 (N_9141,N_8628,N_8913);
nor U9142 (N_9142,N_8804,N_8578);
nand U9143 (N_9143,N_8618,N_8862);
nand U9144 (N_9144,N_8969,N_8941);
nor U9145 (N_9145,N_8693,N_8914);
and U9146 (N_9146,N_8557,N_8689);
xnor U9147 (N_9147,N_8538,N_8953);
and U9148 (N_9148,N_8605,N_8574);
xor U9149 (N_9149,N_8718,N_8738);
or U9150 (N_9150,N_8637,N_8592);
or U9151 (N_9151,N_8694,N_8959);
and U9152 (N_9152,N_8779,N_8569);
or U9153 (N_9153,N_8540,N_8521);
xor U9154 (N_9154,N_8986,N_8728);
nand U9155 (N_9155,N_8678,N_8903);
or U9156 (N_9156,N_8868,N_8948);
xor U9157 (N_9157,N_8908,N_8772);
and U9158 (N_9158,N_8734,N_8587);
nor U9159 (N_9159,N_8801,N_8811);
xor U9160 (N_9160,N_8938,N_8816);
nor U9161 (N_9161,N_8830,N_8787);
nor U9162 (N_9162,N_8639,N_8653);
xor U9163 (N_9163,N_8612,N_8834);
nor U9164 (N_9164,N_8867,N_8927);
and U9165 (N_9165,N_8814,N_8708);
nor U9166 (N_9166,N_8753,N_8987);
and U9167 (N_9167,N_8897,N_8650);
and U9168 (N_9168,N_8887,N_8553);
or U9169 (N_9169,N_8669,N_8852);
nor U9170 (N_9170,N_8901,N_8861);
or U9171 (N_9171,N_8856,N_8542);
and U9172 (N_9172,N_8640,N_8918);
nor U9173 (N_9173,N_8537,N_8777);
nor U9174 (N_9174,N_8665,N_8711);
and U9175 (N_9175,N_8782,N_8501);
nor U9176 (N_9176,N_8671,N_8933);
or U9177 (N_9177,N_8832,N_8823);
or U9178 (N_9178,N_8756,N_8735);
nand U9179 (N_9179,N_8724,N_8993);
nand U9180 (N_9180,N_8791,N_8855);
or U9181 (N_9181,N_8552,N_8812);
and U9182 (N_9182,N_8625,N_8621);
xnor U9183 (N_9183,N_8559,N_8894);
xnor U9184 (N_9184,N_8701,N_8895);
nand U9185 (N_9185,N_8530,N_8747);
nand U9186 (N_9186,N_8951,N_8904);
or U9187 (N_9187,N_8691,N_8737);
and U9188 (N_9188,N_8601,N_8598);
nand U9189 (N_9189,N_8945,N_8962);
nor U9190 (N_9190,N_8740,N_8931);
xor U9191 (N_9191,N_8731,N_8885);
or U9192 (N_9192,N_8978,N_8786);
nor U9193 (N_9193,N_8970,N_8539);
xor U9194 (N_9194,N_8619,N_8608);
xnor U9195 (N_9195,N_8550,N_8541);
and U9196 (N_9196,N_8841,N_8680);
or U9197 (N_9197,N_8614,N_8622);
xnor U9198 (N_9198,N_8910,N_8839);
xnor U9199 (N_9199,N_8965,N_8992);
nor U9200 (N_9200,N_8714,N_8596);
xnor U9201 (N_9201,N_8911,N_8988);
xnor U9202 (N_9202,N_8857,N_8909);
nand U9203 (N_9203,N_8545,N_8571);
or U9204 (N_9204,N_8645,N_8613);
and U9205 (N_9205,N_8580,N_8543);
xnor U9206 (N_9206,N_8886,N_8611);
nor U9207 (N_9207,N_8939,N_8732);
or U9208 (N_9208,N_8722,N_8635);
or U9209 (N_9209,N_8845,N_8873);
xor U9210 (N_9210,N_8588,N_8582);
or U9211 (N_9211,N_8604,N_8944);
or U9212 (N_9212,N_8676,N_8570);
nand U9213 (N_9213,N_8529,N_8919);
xnor U9214 (N_9214,N_8723,N_8818);
or U9215 (N_9215,N_8870,N_8967);
and U9216 (N_9216,N_8796,N_8750);
or U9217 (N_9217,N_8518,N_8837);
xnor U9218 (N_9218,N_8879,N_8715);
xnor U9219 (N_9219,N_8905,N_8874);
and U9220 (N_9220,N_8623,N_8654);
nand U9221 (N_9221,N_8568,N_8503);
or U9222 (N_9222,N_8920,N_8888);
nor U9223 (N_9223,N_8700,N_8741);
xnor U9224 (N_9224,N_8809,N_8906);
or U9225 (N_9225,N_8562,N_8826);
nand U9226 (N_9226,N_8527,N_8514);
xor U9227 (N_9227,N_8595,N_8726);
xor U9228 (N_9228,N_8651,N_8982);
nand U9229 (N_9229,N_8695,N_8915);
and U9230 (N_9230,N_8742,N_8673);
nand U9231 (N_9231,N_8775,N_8533);
or U9232 (N_9232,N_8843,N_8842);
or U9233 (N_9233,N_8763,N_8769);
xnor U9234 (N_9234,N_8890,N_8577);
and U9235 (N_9235,N_8646,N_8990);
nor U9236 (N_9236,N_8822,N_8795);
nand U9237 (N_9237,N_8566,N_8626);
nand U9238 (N_9238,N_8891,N_8898);
xor U9239 (N_9239,N_8702,N_8581);
nand U9240 (N_9240,N_8594,N_8859);
nor U9241 (N_9241,N_8878,N_8717);
or U9242 (N_9242,N_8831,N_8563);
and U9243 (N_9243,N_8923,N_8517);
nor U9244 (N_9244,N_8833,N_8754);
nand U9245 (N_9245,N_8778,N_8788);
nand U9246 (N_9246,N_8549,N_8739);
nand U9247 (N_9247,N_8979,N_8956);
nand U9248 (N_9248,N_8815,N_8937);
nor U9249 (N_9249,N_8983,N_8720);
and U9250 (N_9250,N_8974,N_8786);
xor U9251 (N_9251,N_8825,N_8635);
and U9252 (N_9252,N_8845,N_8711);
and U9253 (N_9253,N_8741,N_8501);
nand U9254 (N_9254,N_8909,N_8793);
xor U9255 (N_9255,N_8781,N_8993);
nor U9256 (N_9256,N_8510,N_8759);
nand U9257 (N_9257,N_8611,N_8679);
nor U9258 (N_9258,N_8739,N_8845);
and U9259 (N_9259,N_8823,N_8698);
nand U9260 (N_9260,N_8677,N_8631);
and U9261 (N_9261,N_8738,N_8503);
and U9262 (N_9262,N_8677,N_8916);
or U9263 (N_9263,N_8882,N_8654);
nand U9264 (N_9264,N_8641,N_8747);
xnor U9265 (N_9265,N_8752,N_8870);
and U9266 (N_9266,N_8755,N_8914);
xnor U9267 (N_9267,N_8707,N_8820);
xnor U9268 (N_9268,N_8863,N_8833);
and U9269 (N_9269,N_8903,N_8869);
nor U9270 (N_9270,N_8870,N_8529);
nand U9271 (N_9271,N_8731,N_8837);
and U9272 (N_9272,N_8836,N_8521);
and U9273 (N_9273,N_8980,N_8914);
or U9274 (N_9274,N_8884,N_8579);
xnor U9275 (N_9275,N_8578,N_8820);
or U9276 (N_9276,N_8554,N_8890);
xnor U9277 (N_9277,N_8781,N_8591);
nand U9278 (N_9278,N_8595,N_8950);
nand U9279 (N_9279,N_8574,N_8643);
and U9280 (N_9280,N_8897,N_8538);
nand U9281 (N_9281,N_8911,N_8970);
xor U9282 (N_9282,N_8590,N_8730);
nand U9283 (N_9283,N_8686,N_8897);
nor U9284 (N_9284,N_8941,N_8746);
and U9285 (N_9285,N_8516,N_8656);
xor U9286 (N_9286,N_8885,N_8974);
and U9287 (N_9287,N_8638,N_8762);
or U9288 (N_9288,N_8897,N_8760);
nor U9289 (N_9289,N_8912,N_8990);
xnor U9290 (N_9290,N_8935,N_8941);
xnor U9291 (N_9291,N_8751,N_8934);
nand U9292 (N_9292,N_8905,N_8695);
nand U9293 (N_9293,N_8919,N_8526);
xnor U9294 (N_9294,N_8706,N_8510);
nor U9295 (N_9295,N_8743,N_8823);
and U9296 (N_9296,N_8723,N_8578);
and U9297 (N_9297,N_8792,N_8906);
nand U9298 (N_9298,N_8593,N_8842);
xnor U9299 (N_9299,N_8864,N_8537);
and U9300 (N_9300,N_8593,N_8825);
and U9301 (N_9301,N_8688,N_8596);
nand U9302 (N_9302,N_8876,N_8799);
and U9303 (N_9303,N_8748,N_8869);
nand U9304 (N_9304,N_8610,N_8816);
nor U9305 (N_9305,N_8955,N_8926);
or U9306 (N_9306,N_8504,N_8531);
nand U9307 (N_9307,N_8805,N_8512);
and U9308 (N_9308,N_8510,N_8812);
nor U9309 (N_9309,N_8711,N_8923);
nor U9310 (N_9310,N_8673,N_8976);
nand U9311 (N_9311,N_8535,N_8545);
nor U9312 (N_9312,N_8984,N_8634);
xnor U9313 (N_9313,N_8730,N_8577);
or U9314 (N_9314,N_8966,N_8822);
or U9315 (N_9315,N_8838,N_8567);
nor U9316 (N_9316,N_8747,N_8719);
xor U9317 (N_9317,N_8819,N_8517);
or U9318 (N_9318,N_8947,N_8771);
nor U9319 (N_9319,N_8595,N_8763);
nand U9320 (N_9320,N_8885,N_8829);
and U9321 (N_9321,N_8743,N_8769);
or U9322 (N_9322,N_8630,N_8893);
nor U9323 (N_9323,N_8867,N_8593);
nor U9324 (N_9324,N_8591,N_8717);
or U9325 (N_9325,N_8728,N_8821);
and U9326 (N_9326,N_8784,N_8660);
xnor U9327 (N_9327,N_8611,N_8728);
nor U9328 (N_9328,N_8928,N_8834);
xnor U9329 (N_9329,N_8582,N_8540);
or U9330 (N_9330,N_8896,N_8987);
and U9331 (N_9331,N_8791,N_8869);
and U9332 (N_9332,N_8701,N_8532);
nand U9333 (N_9333,N_8507,N_8576);
or U9334 (N_9334,N_8944,N_8665);
xor U9335 (N_9335,N_8770,N_8987);
and U9336 (N_9336,N_8875,N_8964);
and U9337 (N_9337,N_8579,N_8933);
nand U9338 (N_9338,N_8834,N_8970);
or U9339 (N_9339,N_8996,N_8602);
xnor U9340 (N_9340,N_8536,N_8752);
xnor U9341 (N_9341,N_8528,N_8919);
or U9342 (N_9342,N_8533,N_8866);
and U9343 (N_9343,N_8645,N_8833);
xnor U9344 (N_9344,N_8671,N_8854);
and U9345 (N_9345,N_8859,N_8787);
nand U9346 (N_9346,N_8822,N_8730);
xor U9347 (N_9347,N_8617,N_8770);
nand U9348 (N_9348,N_8781,N_8567);
nand U9349 (N_9349,N_8987,N_8503);
and U9350 (N_9350,N_8710,N_8657);
or U9351 (N_9351,N_8899,N_8633);
and U9352 (N_9352,N_8707,N_8625);
nor U9353 (N_9353,N_8657,N_8895);
nand U9354 (N_9354,N_8770,N_8660);
nand U9355 (N_9355,N_8996,N_8679);
nand U9356 (N_9356,N_8972,N_8668);
or U9357 (N_9357,N_8814,N_8936);
nand U9358 (N_9358,N_8508,N_8832);
nand U9359 (N_9359,N_8776,N_8737);
nand U9360 (N_9360,N_8738,N_8722);
nand U9361 (N_9361,N_8691,N_8623);
xor U9362 (N_9362,N_8752,N_8692);
xor U9363 (N_9363,N_8935,N_8547);
and U9364 (N_9364,N_8939,N_8784);
or U9365 (N_9365,N_8755,N_8936);
nand U9366 (N_9366,N_8763,N_8984);
nand U9367 (N_9367,N_8859,N_8917);
nand U9368 (N_9368,N_8737,N_8550);
nand U9369 (N_9369,N_8549,N_8851);
and U9370 (N_9370,N_8984,N_8561);
and U9371 (N_9371,N_8652,N_8844);
nand U9372 (N_9372,N_8908,N_8792);
nand U9373 (N_9373,N_8710,N_8560);
nand U9374 (N_9374,N_8874,N_8963);
nor U9375 (N_9375,N_8925,N_8582);
xnor U9376 (N_9376,N_8963,N_8722);
xnor U9377 (N_9377,N_8536,N_8961);
and U9378 (N_9378,N_8880,N_8556);
and U9379 (N_9379,N_8902,N_8698);
nor U9380 (N_9380,N_8690,N_8688);
nand U9381 (N_9381,N_8577,N_8845);
nor U9382 (N_9382,N_8586,N_8679);
or U9383 (N_9383,N_8610,N_8758);
nand U9384 (N_9384,N_8686,N_8887);
or U9385 (N_9385,N_8835,N_8803);
and U9386 (N_9386,N_8927,N_8934);
and U9387 (N_9387,N_8752,N_8821);
nor U9388 (N_9388,N_8618,N_8870);
and U9389 (N_9389,N_8996,N_8740);
xor U9390 (N_9390,N_8500,N_8633);
xor U9391 (N_9391,N_8543,N_8789);
nor U9392 (N_9392,N_8620,N_8875);
nor U9393 (N_9393,N_8784,N_8860);
nor U9394 (N_9394,N_8839,N_8502);
or U9395 (N_9395,N_8737,N_8570);
and U9396 (N_9396,N_8753,N_8668);
xnor U9397 (N_9397,N_8680,N_8944);
or U9398 (N_9398,N_8683,N_8998);
nand U9399 (N_9399,N_8906,N_8942);
xnor U9400 (N_9400,N_8922,N_8633);
xor U9401 (N_9401,N_8737,N_8650);
and U9402 (N_9402,N_8580,N_8740);
nor U9403 (N_9403,N_8632,N_8872);
nor U9404 (N_9404,N_8902,N_8533);
xnor U9405 (N_9405,N_8859,N_8655);
xor U9406 (N_9406,N_8783,N_8507);
and U9407 (N_9407,N_8883,N_8656);
nand U9408 (N_9408,N_8691,N_8538);
nand U9409 (N_9409,N_8745,N_8506);
nand U9410 (N_9410,N_8543,N_8716);
nand U9411 (N_9411,N_8949,N_8638);
nor U9412 (N_9412,N_8987,N_8855);
nand U9413 (N_9413,N_8508,N_8985);
and U9414 (N_9414,N_8983,N_8793);
nand U9415 (N_9415,N_8707,N_8764);
and U9416 (N_9416,N_8777,N_8734);
or U9417 (N_9417,N_8914,N_8875);
or U9418 (N_9418,N_8829,N_8627);
and U9419 (N_9419,N_8883,N_8593);
nor U9420 (N_9420,N_8611,N_8536);
and U9421 (N_9421,N_8756,N_8873);
xnor U9422 (N_9422,N_8715,N_8770);
nand U9423 (N_9423,N_8503,N_8931);
and U9424 (N_9424,N_8530,N_8845);
and U9425 (N_9425,N_8517,N_8798);
xnor U9426 (N_9426,N_8537,N_8741);
nand U9427 (N_9427,N_8801,N_8874);
or U9428 (N_9428,N_8677,N_8925);
nor U9429 (N_9429,N_8681,N_8625);
or U9430 (N_9430,N_8926,N_8980);
nor U9431 (N_9431,N_8581,N_8567);
xnor U9432 (N_9432,N_8685,N_8627);
and U9433 (N_9433,N_8540,N_8996);
nand U9434 (N_9434,N_8546,N_8577);
xor U9435 (N_9435,N_8872,N_8986);
nor U9436 (N_9436,N_8543,N_8934);
nor U9437 (N_9437,N_8849,N_8877);
nand U9438 (N_9438,N_8758,N_8877);
nor U9439 (N_9439,N_8968,N_8801);
xnor U9440 (N_9440,N_8974,N_8743);
and U9441 (N_9441,N_8640,N_8697);
xnor U9442 (N_9442,N_8570,N_8960);
and U9443 (N_9443,N_8628,N_8776);
xnor U9444 (N_9444,N_8572,N_8728);
xor U9445 (N_9445,N_8880,N_8857);
xnor U9446 (N_9446,N_8641,N_8625);
or U9447 (N_9447,N_8642,N_8990);
or U9448 (N_9448,N_8723,N_8684);
nor U9449 (N_9449,N_8820,N_8751);
xor U9450 (N_9450,N_8797,N_8822);
nor U9451 (N_9451,N_8923,N_8770);
nand U9452 (N_9452,N_8859,N_8709);
or U9453 (N_9453,N_8834,N_8951);
nand U9454 (N_9454,N_8709,N_8523);
or U9455 (N_9455,N_8587,N_8855);
nor U9456 (N_9456,N_8903,N_8832);
nand U9457 (N_9457,N_8946,N_8901);
or U9458 (N_9458,N_8642,N_8823);
and U9459 (N_9459,N_8566,N_8622);
nor U9460 (N_9460,N_8633,N_8667);
xor U9461 (N_9461,N_8814,N_8971);
xnor U9462 (N_9462,N_8691,N_8863);
or U9463 (N_9463,N_8743,N_8678);
nor U9464 (N_9464,N_8832,N_8816);
nor U9465 (N_9465,N_8669,N_8800);
nor U9466 (N_9466,N_8642,N_8811);
or U9467 (N_9467,N_8730,N_8721);
nor U9468 (N_9468,N_8623,N_8937);
and U9469 (N_9469,N_8966,N_8802);
and U9470 (N_9470,N_8641,N_8782);
nor U9471 (N_9471,N_8765,N_8549);
nand U9472 (N_9472,N_8544,N_8538);
xor U9473 (N_9473,N_8742,N_8558);
nand U9474 (N_9474,N_8708,N_8804);
xor U9475 (N_9475,N_8892,N_8647);
and U9476 (N_9476,N_8709,N_8596);
nand U9477 (N_9477,N_8684,N_8639);
or U9478 (N_9478,N_8704,N_8587);
and U9479 (N_9479,N_8528,N_8856);
xnor U9480 (N_9480,N_8794,N_8508);
nand U9481 (N_9481,N_8506,N_8924);
xnor U9482 (N_9482,N_8912,N_8692);
or U9483 (N_9483,N_8799,N_8964);
xnor U9484 (N_9484,N_8506,N_8738);
and U9485 (N_9485,N_8622,N_8819);
xnor U9486 (N_9486,N_8818,N_8541);
nor U9487 (N_9487,N_8600,N_8625);
nand U9488 (N_9488,N_8948,N_8598);
nor U9489 (N_9489,N_8633,N_8727);
nor U9490 (N_9490,N_8659,N_8579);
xnor U9491 (N_9491,N_8837,N_8909);
and U9492 (N_9492,N_8682,N_8829);
and U9493 (N_9493,N_8953,N_8853);
or U9494 (N_9494,N_8793,N_8516);
xor U9495 (N_9495,N_8749,N_8750);
or U9496 (N_9496,N_8782,N_8874);
or U9497 (N_9497,N_8681,N_8813);
or U9498 (N_9498,N_8778,N_8909);
xor U9499 (N_9499,N_8654,N_8903);
xor U9500 (N_9500,N_9149,N_9125);
and U9501 (N_9501,N_9304,N_9392);
nor U9502 (N_9502,N_9394,N_9129);
xor U9503 (N_9503,N_9439,N_9245);
xor U9504 (N_9504,N_9353,N_9088);
or U9505 (N_9505,N_9223,N_9481);
or U9506 (N_9506,N_9424,N_9135);
and U9507 (N_9507,N_9253,N_9179);
xnor U9508 (N_9508,N_9431,N_9073);
and U9509 (N_9509,N_9087,N_9209);
nand U9510 (N_9510,N_9446,N_9458);
nor U9511 (N_9511,N_9013,N_9367);
nand U9512 (N_9512,N_9117,N_9146);
and U9513 (N_9513,N_9473,N_9200);
and U9514 (N_9514,N_9410,N_9077);
and U9515 (N_9515,N_9123,N_9252);
or U9516 (N_9516,N_9463,N_9427);
nand U9517 (N_9517,N_9346,N_9264);
nor U9518 (N_9518,N_9051,N_9413);
nor U9519 (N_9519,N_9398,N_9406);
or U9520 (N_9520,N_9169,N_9444);
nor U9521 (N_9521,N_9495,N_9277);
and U9522 (N_9522,N_9315,N_9079);
or U9523 (N_9523,N_9379,N_9488);
xor U9524 (N_9524,N_9216,N_9498);
nor U9525 (N_9525,N_9342,N_9303);
and U9526 (N_9526,N_9229,N_9474);
nor U9527 (N_9527,N_9081,N_9181);
nand U9528 (N_9528,N_9449,N_9005);
xor U9529 (N_9529,N_9151,N_9355);
nor U9530 (N_9530,N_9261,N_9199);
nor U9531 (N_9531,N_9015,N_9138);
nor U9532 (N_9532,N_9065,N_9409);
xor U9533 (N_9533,N_9365,N_9349);
nor U9534 (N_9534,N_9034,N_9066);
nor U9535 (N_9535,N_9140,N_9113);
and U9536 (N_9536,N_9395,N_9174);
nand U9537 (N_9537,N_9150,N_9399);
nor U9538 (N_9538,N_9064,N_9256);
xnor U9539 (N_9539,N_9244,N_9322);
or U9540 (N_9540,N_9120,N_9247);
nor U9541 (N_9541,N_9496,N_9468);
nand U9542 (N_9542,N_9197,N_9335);
and U9543 (N_9543,N_9075,N_9376);
nor U9544 (N_9544,N_9457,N_9320);
nand U9545 (N_9545,N_9327,N_9499);
nand U9546 (N_9546,N_9196,N_9471);
or U9547 (N_9547,N_9071,N_9221);
nand U9548 (N_9548,N_9311,N_9428);
or U9549 (N_9549,N_9106,N_9483);
or U9550 (N_9550,N_9144,N_9348);
nand U9551 (N_9551,N_9275,N_9130);
or U9552 (N_9552,N_9175,N_9121);
xor U9553 (N_9553,N_9103,N_9262);
or U9554 (N_9554,N_9132,N_9198);
nand U9555 (N_9555,N_9340,N_9260);
nor U9556 (N_9556,N_9308,N_9053);
or U9557 (N_9557,N_9152,N_9239);
or U9558 (N_9558,N_9302,N_9313);
xnor U9559 (N_9559,N_9194,N_9494);
nand U9560 (N_9560,N_9105,N_9435);
or U9561 (N_9561,N_9212,N_9257);
xnor U9562 (N_9562,N_9116,N_9419);
xnor U9563 (N_9563,N_9300,N_9434);
and U9564 (N_9564,N_9141,N_9270);
nor U9565 (N_9565,N_9094,N_9301);
xor U9566 (N_9566,N_9234,N_9345);
xnor U9567 (N_9567,N_9241,N_9272);
nor U9568 (N_9568,N_9085,N_9204);
nor U9569 (N_9569,N_9017,N_9233);
xor U9570 (N_9570,N_9203,N_9102);
or U9571 (N_9571,N_9442,N_9237);
or U9572 (N_9572,N_9432,N_9029);
xor U9573 (N_9573,N_9180,N_9248);
or U9574 (N_9574,N_9287,N_9238);
nor U9575 (N_9575,N_9067,N_9372);
and U9576 (N_9576,N_9030,N_9389);
xnor U9577 (N_9577,N_9014,N_9492);
nor U9578 (N_9578,N_9405,N_9470);
nor U9579 (N_9579,N_9267,N_9069);
nor U9580 (N_9580,N_9288,N_9265);
nor U9581 (N_9581,N_9326,N_9091);
nand U9582 (N_9582,N_9447,N_9222);
xor U9583 (N_9583,N_9385,N_9182);
xnor U9584 (N_9584,N_9210,N_9191);
and U9585 (N_9585,N_9154,N_9176);
and U9586 (N_9586,N_9039,N_9416);
and U9587 (N_9587,N_9321,N_9429);
and U9588 (N_9588,N_9329,N_9050);
or U9589 (N_9589,N_9018,N_9273);
and U9590 (N_9590,N_9477,N_9185);
nand U9591 (N_9591,N_9258,N_9104);
nor U9592 (N_9592,N_9041,N_9004);
nor U9593 (N_9593,N_9478,N_9192);
nor U9594 (N_9594,N_9453,N_9083);
or U9595 (N_9595,N_9299,N_9173);
xor U9596 (N_9596,N_9049,N_9207);
or U9597 (N_9597,N_9019,N_9323);
nand U9598 (N_9598,N_9430,N_9250);
nor U9599 (N_9599,N_9309,N_9297);
nand U9600 (N_9600,N_9225,N_9070);
or U9601 (N_9601,N_9023,N_9358);
xor U9602 (N_9602,N_9437,N_9168);
or U9603 (N_9603,N_9443,N_9084);
nand U9604 (N_9604,N_9040,N_9354);
xnor U9605 (N_9605,N_9324,N_9112);
nor U9606 (N_9606,N_9415,N_9111);
or U9607 (N_9607,N_9027,N_9373);
or U9608 (N_9608,N_9178,N_9008);
xnor U9609 (N_9609,N_9356,N_9080);
xor U9610 (N_9610,N_9156,N_9279);
nor U9611 (N_9611,N_9128,N_9240);
nand U9612 (N_9612,N_9361,N_9161);
and U9613 (N_9613,N_9386,N_9134);
xnor U9614 (N_9614,N_9285,N_9167);
or U9615 (N_9615,N_9206,N_9171);
or U9616 (N_9616,N_9391,N_9158);
or U9617 (N_9617,N_9318,N_9452);
and U9618 (N_9618,N_9246,N_9445);
xnor U9619 (N_9619,N_9086,N_9371);
or U9620 (N_9620,N_9193,N_9314);
or U9621 (N_9621,N_9296,N_9284);
or U9622 (N_9622,N_9290,N_9189);
or U9623 (N_9623,N_9145,N_9126);
and U9624 (N_9624,N_9336,N_9352);
xnor U9625 (N_9625,N_9251,N_9114);
xor U9626 (N_9626,N_9160,N_9078);
nand U9627 (N_9627,N_9139,N_9387);
nor U9628 (N_9628,N_9357,N_9142);
nor U9629 (N_9629,N_9215,N_9426);
nand U9630 (N_9630,N_9031,N_9487);
and U9631 (N_9631,N_9057,N_9440);
nand U9632 (N_9632,N_9407,N_9164);
xnor U9633 (N_9633,N_9059,N_9025);
or U9634 (N_9634,N_9054,N_9006);
nor U9635 (N_9635,N_9016,N_9119);
nor U9636 (N_9636,N_9307,N_9062);
or U9637 (N_9637,N_9289,N_9096);
nor U9638 (N_9638,N_9100,N_9107);
and U9639 (N_9639,N_9363,N_9208);
xnor U9640 (N_9640,N_9166,N_9411);
nor U9641 (N_9641,N_9249,N_9047);
or U9642 (N_9642,N_9131,N_9147);
nor U9643 (N_9643,N_9032,N_9186);
nand U9644 (N_9644,N_9493,N_9400);
nor U9645 (N_9645,N_9375,N_9101);
nor U9646 (N_9646,N_9421,N_9020);
nand U9647 (N_9647,N_9089,N_9092);
or U9648 (N_9648,N_9339,N_9118);
or U9649 (N_9649,N_9045,N_9479);
nor U9650 (N_9650,N_9157,N_9475);
or U9651 (N_9651,N_9343,N_9026);
and U9652 (N_9652,N_9305,N_9072);
nand U9653 (N_9653,N_9042,N_9286);
nor U9654 (N_9654,N_9384,N_9122);
nor U9655 (N_9655,N_9162,N_9009);
and U9656 (N_9656,N_9362,N_9044);
and U9657 (N_9657,N_9382,N_9063);
or U9658 (N_9658,N_9211,N_9124);
nor U9659 (N_9659,N_9055,N_9317);
or U9660 (N_9660,N_9095,N_9422);
nand U9661 (N_9661,N_9283,N_9414);
nor U9662 (N_9662,N_9451,N_9282);
nand U9663 (N_9663,N_9011,N_9060);
nand U9664 (N_9664,N_9331,N_9390);
or U9665 (N_9665,N_9058,N_9010);
nor U9666 (N_9666,N_9485,N_9404);
or U9667 (N_9667,N_9364,N_9456);
and U9668 (N_9668,N_9061,N_9330);
xnor U9669 (N_9669,N_9201,N_9316);
and U9670 (N_9670,N_9374,N_9450);
or U9671 (N_9671,N_9155,N_9377);
nand U9672 (N_9672,N_9338,N_9219);
or U9673 (N_9673,N_9441,N_9480);
and U9674 (N_9674,N_9347,N_9036);
xnor U9675 (N_9675,N_9417,N_9076);
nand U9676 (N_9676,N_9369,N_9337);
nor U9677 (N_9677,N_9035,N_9022);
nor U9678 (N_9678,N_9214,N_9436);
xor U9679 (N_9679,N_9403,N_9127);
nor U9680 (N_9680,N_9002,N_9412);
nor U9681 (N_9681,N_9325,N_9046);
or U9682 (N_9682,N_9438,N_9388);
and U9683 (N_9683,N_9205,N_9213);
nor U9684 (N_9684,N_9108,N_9467);
nand U9685 (N_9685,N_9228,N_9136);
xor U9686 (N_9686,N_9271,N_9217);
xnor U9687 (N_9687,N_9295,N_9202);
xor U9688 (N_9688,N_9266,N_9052);
nand U9689 (N_9689,N_9469,N_9466);
and U9690 (N_9690,N_9484,N_9235);
or U9691 (N_9691,N_9236,N_9056);
nor U9692 (N_9692,N_9226,N_9098);
nand U9693 (N_9693,N_9269,N_9489);
and U9694 (N_9694,N_9433,N_9291);
xor U9695 (N_9695,N_9243,N_9263);
and U9696 (N_9696,N_9274,N_9190);
and U9697 (N_9697,N_9038,N_9418);
nor U9698 (N_9698,N_9328,N_9153);
nand U9699 (N_9699,N_9276,N_9278);
nor U9700 (N_9700,N_9227,N_9230);
nor U9701 (N_9701,N_9048,N_9177);
xnor U9702 (N_9702,N_9007,N_9195);
nand U9703 (N_9703,N_9242,N_9082);
nand U9704 (N_9704,N_9133,N_9159);
or U9705 (N_9705,N_9280,N_9137);
nand U9706 (N_9706,N_9401,N_9043);
nand U9707 (N_9707,N_9491,N_9490);
xor U9708 (N_9708,N_9380,N_9464);
nand U9709 (N_9709,N_9000,N_9420);
nand U9710 (N_9710,N_9319,N_9455);
nor U9711 (N_9711,N_9184,N_9218);
nor U9712 (N_9712,N_9187,N_9381);
nor U9713 (N_9713,N_9143,N_9028);
or U9714 (N_9714,N_9482,N_9472);
xnor U9715 (N_9715,N_9097,N_9110);
nand U9716 (N_9716,N_9476,N_9099);
and U9717 (N_9717,N_9220,N_9462);
or U9718 (N_9718,N_9344,N_9170);
nand U9719 (N_9719,N_9460,N_9334);
and U9720 (N_9720,N_9090,N_9459);
and U9721 (N_9721,N_9093,N_9231);
xor U9722 (N_9722,N_9366,N_9312);
nand U9723 (N_9723,N_9281,N_9359);
nor U9724 (N_9724,N_9292,N_9293);
or U9725 (N_9725,N_9306,N_9074);
nand U9726 (N_9726,N_9341,N_9448);
and U9727 (N_9727,N_9012,N_9497);
nor U9728 (N_9728,N_9294,N_9454);
nand U9729 (N_9729,N_9232,N_9332);
and U9730 (N_9730,N_9024,N_9259);
or U9731 (N_9731,N_9172,N_9461);
nor U9732 (N_9732,N_9383,N_9350);
nand U9733 (N_9733,N_9370,N_9360);
nand U9734 (N_9734,N_9115,N_9310);
and U9735 (N_9735,N_9423,N_9001);
nand U9736 (N_9736,N_9425,N_9068);
and U9737 (N_9737,N_9254,N_9465);
or U9738 (N_9738,N_9165,N_9396);
nand U9739 (N_9739,N_9333,N_9298);
and U9740 (N_9740,N_9268,N_9037);
nand U9741 (N_9741,N_9183,N_9163);
or U9742 (N_9742,N_9148,N_9021);
or U9743 (N_9743,N_9255,N_9378);
and U9744 (N_9744,N_9368,N_9402);
nor U9745 (N_9745,N_9393,N_9486);
and U9746 (N_9746,N_9109,N_9224);
or U9747 (N_9747,N_9188,N_9351);
and U9748 (N_9748,N_9408,N_9003);
or U9749 (N_9749,N_9397,N_9033);
nand U9750 (N_9750,N_9044,N_9312);
xnor U9751 (N_9751,N_9486,N_9451);
xnor U9752 (N_9752,N_9018,N_9132);
and U9753 (N_9753,N_9337,N_9018);
nor U9754 (N_9754,N_9054,N_9287);
and U9755 (N_9755,N_9196,N_9053);
nand U9756 (N_9756,N_9277,N_9171);
and U9757 (N_9757,N_9023,N_9364);
nor U9758 (N_9758,N_9173,N_9233);
nand U9759 (N_9759,N_9348,N_9000);
nand U9760 (N_9760,N_9113,N_9310);
nor U9761 (N_9761,N_9006,N_9246);
xor U9762 (N_9762,N_9325,N_9428);
or U9763 (N_9763,N_9043,N_9310);
or U9764 (N_9764,N_9290,N_9035);
xnor U9765 (N_9765,N_9002,N_9493);
xor U9766 (N_9766,N_9412,N_9052);
xnor U9767 (N_9767,N_9169,N_9335);
xor U9768 (N_9768,N_9337,N_9131);
or U9769 (N_9769,N_9386,N_9079);
and U9770 (N_9770,N_9218,N_9302);
and U9771 (N_9771,N_9367,N_9391);
nor U9772 (N_9772,N_9118,N_9319);
or U9773 (N_9773,N_9105,N_9027);
nor U9774 (N_9774,N_9266,N_9064);
or U9775 (N_9775,N_9474,N_9359);
xor U9776 (N_9776,N_9008,N_9398);
or U9777 (N_9777,N_9457,N_9243);
or U9778 (N_9778,N_9100,N_9430);
and U9779 (N_9779,N_9002,N_9009);
nand U9780 (N_9780,N_9173,N_9161);
nand U9781 (N_9781,N_9194,N_9466);
and U9782 (N_9782,N_9360,N_9308);
xnor U9783 (N_9783,N_9184,N_9286);
xnor U9784 (N_9784,N_9434,N_9212);
nor U9785 (N_9785,N_9426,N_9126);
and U9786 (N_9786,N_9184,N_9401);
nor U9787 (N_9787,N_9018,N_9455);
nand U9788 (N_9788,N_9025,N_9085);
or U9789 (N_9789,N_9294,N_9360);
nor U9790 (N_9790,N_9351,N_9286);
nor U9791 (N_9791,N_9486,N_9392);
and U9792 (N_9792,N_9155,N_9070);
nor U9793 (N_9793,N_9398,N_9052);
or U9794 (N_9794,N_9320,N_9343);
nand U9795 (N_9795,N_9225,N_9456);
nand U9796 (N_9796,N_9137,N_9191);
and U9797 (N_9797,N_9069,N_9321);
nand U9798 (N_9798,N_9197,N_9309);
xnor U9799 (N_9799,N_9474,N_9083);
nor U9800 (N_9800,N_9155,N_9450);
nor U9801 (N_9801,N_9304,N_9434);
nor U9802 (N_9802,N_9047,N_9165);
nor U9803 (N_9803,N_9240,N_9134);
xor U9804 (N_9804,N_9491,N_9141);
nand U9805 (N_9805,N_9352,N_9293);
nand U9806 (N_9806,N_9165,N_9067);
nor U9807 (N_9807,N_9140,N_9479);
nor U9808 (N_9808,N_9350,N_9495);
nand U9809 (N_9809,N_9482,N_9208);
xor U9810 (N_9810,N_9104,N_9425);
nor U9811 (N_9811,N_9002,N_9437);
or U9812 (N_9812,N_9120,N_9353);
nor U9813 (N_9813,N_9273,N_9483);
xor U9814 (N_9814,N_9065,N_9353);
xnor U9815 (N_9815,N_9146,N_9220);
or U9816 (N_9816,N_9473,N_9407);
nand U9817 (N_9817,N_9378,N_9463);
xor U9818 (N_9818,N_9282,N_9159);
or U9819 (N_9819,N_9003,N_9351);
xor U9820 (N_9820,N_9012,N_9438);
and U9821 (N_9821,N_9390,N_9399);
xor U9822 (N_9822,N_9016,N_9286);
or U9823 (N_9823,N_9256,N_9030);
or U9824 (N_9824,N_9442,N_9142);
and U9825 (N_9825,N_9201,N_9044);
or U9826 (N_9826,N_9277,N_9084);
nor U9827 (N_9827,N_9385,N_9097);
xor U9828 (N_9828,N_9283,N_9351);
nor U9829 (N_9829,N_9146,N_9369);
nand U9830 (N_9830,N_9178,N_9168);
nand U9831 (N_9831,N_9105,N_9080);
nand U9832 (N_9832,N_9218,N_9162);
nor U9833 (N_9833,N_9102,N_9425);
xnor U9834 (N_9834,N_9202,N_9482);
nor U9835 (N_9835,N_9436,N_9276);
or U9836 (N_9836,N_9323,N_9105);
nor U9837 (N_9837,N_9306,N_9399);
nand U9838 (N_9838,N_9080,N_9082);
xnor U9839 (N_9839,N_9003,N_9360);
nand U9840 (N_9840,N_9194,N_9081);
nand U9841 (N_9841,N_9208,N_9146);
and U9842 (N_9842,N_9010,N_9336);
nand U9843 (N_9843,N_9464,N_9141);
nand U9844 (N_9844,N_9282,N_9280);
nand U9845 (N_9845,N_9230,N_9129);
and U9846 (N_9846,N_9378,N_9381);
and U9847 (N_9847,N_9160,N_9342);
nor U9848 (N_9848,N_9176,N_9288);
and U9849 (N_9849,N_9076,N_9159);
and U9850 (N_9850,N_9257,N_9027);
and U9851 (N_9851,N_9357,N_9475);
nor U9852 (N_9852,N_9252,N_9186);
xnor U9853 (N_9853,N_9177,N_9374);
nor U9854 (N_9854,N_9176,N_9128);
or U9855 (N_9855,N_9044,N_9222);
and U9856 (N_9856,N_9324,N_9448);
nand U9857 (N_9857,N_9479,N_9474);
nand U9858 (N_9858,N_9312,N_9036);
and U9859 (N_9859,N_9149,N_9497);
and U9860 (N_9860,N_9394,N_9272);
and U9861 (N_9861,N_9105,N_9385);
xor U9862 (N_9862,N_9485,N_9123);
and U9863 (N_9863,N_9378,N_9406);
nand U9864 (N_9864,N_9071,N_9199);
and U9865 (N_9865,N_9273,N_9121);
and U9866 (N_9866,N_9242,N_9431);
or U9867 (N_9867,N_9466,N_9359);
xor U9868 (N_9868,N_9065,N_9018);
or U9869 (N_9869,N_9200,N_9282);
nand U9870 (N_9870,N_9118,N_9140);
xor U9871 (N_9871,N_9416,N_9180);
nand U9872 (N_9872,N_9009,N_9008);
xor U9873 (N_9873,N_9230,N_9008);
xnor U9874 (N_9874,N_9482,N_9111);
nand U9875 (N_9875,N_9282,N_9477);
or U9876 (N_9876,N_9120,N_9266);
and U9877 (N_9877,N_9069,N_9141);
xnor U9878 (N_9878,N_9073,N_9165);
xor U9879 (N_9879,N_9066,N_9107);
nand U9880 (N_9880,N_9058,N_9130);
or U9881 (N_9881,N_9499,N_9498);
nand U9882 (N_9882,N_9368,N_9182);
or U9883 (N_9883,N_9324,N_9040);
nand U9884 (N_9884,N_9009,N_9098);
nor U9885 (N_9885,N_9436,N_9273);
xor U9886 (N_9886,N_9206,N_9316);
xnor U9887 (N_9887,N_9285,N_9359);
or U9888 (N_9888,N_9196,N_9215);
nand U9889 (N_9889,N_9002,N_9286);
xor U9890 (N_9890,N_9326,N_9391);
nand U9891 (N_9891,N_9257,N_9390);
and U9892 (N_9892,N_9223,N_9186);
nor U9893 (N_9893,N_9316,N_9349);
and U9894 (N_9894,N_9350,N_9160);
nor U9895 (N_9895,N_9147,N_9375);
and U9896 (N_9896,N_9449,N_9023);
nor U9897 (N_9897,N_9391,N_9215);
or U9898 (N_9898,N_9081,N_9058);
or U9899 (N_9899,N_9382,N_9051);
and U9900 (N_9900,N_9223,N_9122);
xnor U9901 (N_9901,N_9030,N_9272);
nor U9902 (N_9902,N_9205,N_9098);
nor U9903 (N_9903,N_9121,N_9478);
xnor U9904 (N_9904,N_9148,N_9446);
or U9905 (N_9905,N_9299,N_9418);
xor U9906 (N_9906,N_9043,N_9426);
or U9907 (N_9907,N_9294,N_9422);
xor U9908 (N_9908,N_9257,N_9351);
nor U9909 (N_9909,N_9324,N_9483);
and U9910 (N_9910,N_9498,N_9436);
or U9911 (N_9911,N_9242,N_9208);
nor U9912 (N_9912,N_9304,N_9474);
xnor U9913 (N_9913,N_9389,N_9253);
and U9914 (N_9914,N_9473,N_9437);
nand U9915 (N_9915,N_9280,N_9377);
nor U9916 (N_9916,N_9275,N_9083);
xnor U9917 (N_9917,N_9006,N_9339);
nand U9918 (N_9918,N_9093,N_9205);
and U9919 (N_9919,N_9135,N_9448);
nand U9920 (N_9920,N_9385,N_9107);
nand U9921 (N_9921,N_9140,N_9016);
xnor U9922 (N_9922,N_9420,N_9271);
nor U9923 (N_9923,N_9016,N_9481);
xnor U9924 (N_9924,N_9470,N_9352);
or U9925 (N_9925,N_9156,N_9384);
and U9926 (N_9926,N_9077,N_9130);
xor U9927 (N_9927,N_9377,N_9175);
nor U9928 (N_9928,N_9008,N_9060);
and U9929 (N_9929,N_9180,N_9262);
nor U9930 (N_9930,N_9214,N_9155);
xor U9931 (N_9931,N_9205,N_9032);
xor U9932 (N_9932,N_9422,N_9191);
xnor U9933 (N_9933,N_9464,N_9060);
or U9934 (N_9934,N_9364,N_9353);
nand U9935 (N_9935,N_9204,N_9493);
and U9936 (N_9936,N_9437,N_9170);
and U9937 (N_9937,N_9181,N_9050);
xnor U9938 (N_9938,N_9062,N_9084);
nand U9939 (N_9939,N_9304,N_9329);
nor U9940 (N_9940,N_9097,N_9310);
and U9941 (N_9941,N_9251,N_9259);
xnor U9942 (N_9942,N_9359,N_9320);
or U9943 (N_9943,N_9170,N_9076);
nor U9944 (N_9944,N_9219,N_9007);
or U9945 (N_9945,N_9246,N_9332);
and U9946 (N_9946,N_9259,N_9371);
nor U9947 (N_9947,N_9049,N_9234);
and U9948 (N_9948,N_9281,N_9439);
nor U9949 (N_9949,N_9248,N_9076);
nand U9950 (N_9950,N_9498,N_9470);
nand U9951 (N_9951,N_9279,N_9385);
and U9952 (N_9952,N_9383,N_9289);
xor U9953 (N_9953,N_9487,N_9243);
nor U9954 (N_9954,N_9257,N_9399);
or U9955 (N_9955,N_9490,N_9254);
nor U9956 (N_9956,N_9073,N_9096);
and U9957 (N_9957,N_9299,N_9479);
or U9958 (N_9958,N_9494,N_9149);
nand U9959 (N_9959,N_9266,N_9380);
or U9960 (N_9960,N_9468,N_9416);
and U9961 (N_9961,N_9494,N_9420);
nor U9962 (N_9962,N_9282,N_9350);
nand U9963 (N_9963,N_9011,N_9268);
and U9964 (N_9964,N_9340,N_9013);
nand U9965 (N_9965,N_9272,N_9346);
nand U9966 (N_9966,N_9465,N_9268);
nor U9967 (N_9967,N_9474,N_9084);
xnor U9968 (N_9968,N_9322,N_9330);
and U9969 (N_9969,N_9426,N_9493);
or U9970 (N_9970,N_9466,N_9316);
nand U9971 (N_9971,N_9375,N_9287);
or U9972 (N_9972,N_9218,N_9074);
nand U9973 (N_9973,N_9357,N_9416);
nand U9974 (N_9974,N_9262,N_9351);
xnor U9975 (N_9975,N_9089,N_9180);
or U9976 (N_9976,N_9059,N_9037);
nor U9977 (N_9977,N_9070,N_9433);
and U9978 (N_9978,N_9315,N_9365);
or U9979 (N_9979,N_9438,N_9409);
and U9980 (N_9980,N_9391,N_9132);
and U9981 (N_9981,N_9465,N_9058);
xnor U9982 (N_9982,N_9257,N_9085);
nor U9983 (N_9983,N_9355,N_9050);
nor U9984 (N_9984,N_9041,N_9495);
nand U9985 (N_9985,N_9305,N_9462);
xor U9986 (N_9986,N_9213,N_9080);
and U9987 (N_9987,N_9355,N_9264);
and U9988 (N_9988,N_9494,N_9118);
xnor U9989 (N_9989,N_9205,N_9498);
xor U9990 (N_9990,N_9294,N_9139);
nor U9991 (N_9991,N_9146,N_9079);
and U9992 (N_9992,N_9443,N_9105);
and U9993 (N_9993,N_9290,N_9463);
nand U9994 (N_9994,N_9073,N_9409);
nand U9995 (N_9995,N_9338,N_9422);
or U9996 (N_9996,N_9325,N_9068);
and U9997 (N_9997,N_9234,N_9078);
xnor U9998 (N_9998,N_9076,N_9324);
xnor U9999 (N_9999,N_9046,N_9181);
nand U10000 (N_10000,N_9740,N_9979);
nor U10001 (N_10001,N_9853,N_9588);
xnor U10002 (N_10002,N_9548,N_9777);
nor U10003 (N_10003,N_9678,N_9667);
xnor U10004 (N_10004,N_9507,N_9929);
nand U10005 (N_10005,N_9623,N_9876);
nor U10006 (N_10006,N_9883,N_9844);
nand U10007 (N_10007,N_9640,N_9556);
and U10008 (N_10008,N_9659,N_9601);
nor U10009 (N_10009,N_9970,N_9945);
nand U10010 (N_10010,N_9734,N_9753);
nor U10011 (N_10011,N_9502,N_9782);
or U10012 (N_10012,N_9531,N_9975);
nand U10013 (N_10013,N_9882,N_9660);
nand U10014 (N_10014,N_9878,N_9893);
nor U10015 (N_10015,N_9772,N_9969);
nor U10016 (N_10016,N_9616,N_9928);
and U10017 (N_10017,N_9527,N_9717);
and U10018 (N_10018,N_9907,N_9776);
xnor U10019 (N_10019,N_9506,N_9936);
or U10020 (N_10020,N_9808,N_9511);
or U10021 (N_10021,N_9791,N_9804);
or U10022 (N_10022,N_9626,N_9741);
nand U10023 (N_10023,N_9879,N_9838);
or U10024 (N_10024,N_9875,N_9578);
nand U10025 (N_10025,N_9648,N_9504);
or U10026 (N_10026,N_9957,N_9728);
nand U10027 (N_10027,N_9747,N_9976);
nand U10028 (N_10028,N_9811,N_9520);
and U10029 (N_10029,N_9888,N_9915);
and U10030 (N_10030,N_9580,N_9974);
or U10031 (N_10031,N_9637,N_9523);
nand U10032 (N_10032,N_9553,N_9916);
nor U10033 (N_10033,N_9906,N_9670);
or U10034 (N_10034,N_9505,N_9650);
or U10035 (N_10035,N_9864,N_9737);
xor U10036 (N_10036,N_9651,N_9971);
nand U10037 (N_10037,N_9887,N_9769);
xor U10038 (N_10038,N_9614,N_9518);
or U10039 (N_10039,N_9503,N_9603);
nor U10040 (N_10040,N_9763,N_9767);
and U10041 (N_10041,N_9951,N_9886);
nand U10042 (N_10042,N_9542,N_9559);
nor U10043 (N_10043,N_9770,N_9942);
and U10044 (N_10044,N_9687,N_9571);
and U10045 (N_10045,N_9829,N_9788);
and U10046 (N_10046,N_9952,N_9819);
and U10047 (N_10047,N_9833,N_9681);
and U10048 (N_10048,N_9733,N_9856);
nand U10049 (N_10049,N_9989,N_9694);
and U10050 (N_10050,N_9963,N_9690);
nor U10051 (N_10051,N_9848,N_9863);
or U10052 (N_10052,N_9644,N_9710);
and U10053 (N_10053,N_9561,N_9684);
and U10054 (N_10054,N_9744,N_9709);
xor U10055 (N_10055,N_9718,N_9865);
xnor U10056 (N_10056,N_9547,N_9755);
xor U10057 (N_10057,N_9999,N_9619);
nand U10058 (N_10058,N_9993,N_9810);
or U10059 (N_10059,N_9815,N_9943);
nand U10060 (N_10060,N_9743,N_9519);
xor U10061 (N_10061,N_9778,N_9742);
nor U10062 (N_10062,N_9587,N_9572);
nand U10063 (N_10063,N_9837,N_9536);
nand U10064 (N_10064,N_9760,N_9600);
or U10065 (N_10065,N_9884,N_9630);
xnor U10066 (N_10066,N_9977,N_9628);
or U10067 (N_10067,N_9522,N_9797);
nand U10068 (N_10068,N_9890,N_9568);
and U10069 (N_10069,N_9754,N_9719);
nand U10070 (N_10070,N_9939,N_9799);
nor U10071 (N_10071,N_9720,N_9521);
and U10072 (N_10072,N_9579,N_9596);
and U10073 (N_10073,N_9908,N_9947);
nor U10074 (N_10074,N_9953,N_9714);
or U10075 (N_10075,N_9570,N_9765);
and U10076 (N_10076,N_9867,N_9533);
and U10077 (N_10077,N_9639,N_9510);
nand U10078 (N_10078,N_9968,N_9849);
nor U10079 (N_10079,N_9857,N_9850);
xnor U10080 (N_10080,N_9780,N_9941);
xnor U10081 (N_10081,N_9679,N_9558);
or U10082 (N_10082,N_9735,N_9983);
or U10083 (N_10083,N_9918,N_9618);
or U10084 (N_10084,N_9610,N_9583);
nor U10085 (N_10085,N_9826,N_9708);
nor U10086 (N_10086,N_9545,N_9560);
xnor U10087 (N_10087,N_9723,N_9529);
nand U10088 (N_10088,N_9792,N_9688);
xor U10089 (N_10089,N_9862,N_9896);
and U10090 (N_10090,N_9698,N_9880);
nand U10091 (N_10091,N_9924,N_9569);
xnor U10092 (N_10092,N_9909,N_9794);
nand U10093 (N_10093,N_9940,N_9736);
nor U10094 (N_10094,N_9784,N_9746);
or U10095 (N_10095,N_9910,N_9814);
and U10096 (N_10096,N_9738,N_9912);
and U10097 (N_10097,N_9582,N_9987);
nor U10098 (N_10098,N_9834,N_9995);
nor U10099 (N_10099,N_9551,N_9972);
and U10100 (N_10100,N_9930,N_9901);
nand U10101 (N_10101,N_9573,N_9696);
xnor U10102 (N_10102,N_9686,N_9635);
or U10103 (N_10103,N_9593,N_9641);
xor U10104 (N_10104,N_9775,N_9988);
xor U10105 (N_10105,N_9855,N_9552);
xnor U10106 (N_10106,N_9994,N_9615);
or U10107 (N_10107,N_9996,N_9665);
and U10108 (N_10108,N_9576,N_9567);
nand U10109 (N_10109,N_9591,N_9549);
or U10110 (N_10110,N_9661,N_9956);
xor U10111 (N_10111,N_9955,N_9801);
nor U10112 (N_10112,N_9731,N_9828);
or U10113 (N_10113,N_9873,N_9611);
nor U10114 (N_10114,N_9962,N_9795);
nand U10115 (N_10115,N_9807,N_9858);
nor U10116 (N_10116,N_9509,N_9786);
or U10117 (N_10117,N_9535,N_9689);
nor U10118 (N_10118,N_9745,N_9960);
nand U10119 (N_10119,N_9816,N_9701);
nor U10120 (N_10120,N_9897,N_9827);
nand U10121 (N_10121,N_9885,N_9851);
nor U10122 (N_10122,N_9861,N_9805);
or U10123 (N_10123,N_9779,N_9725);
nand U10124 (N_10124,N_9564,N_9721);
nand U10125 (N_10125,N_9562,N_9716);
nor U10126 (N_10126,N_9715,N_9904);
xor U10127 (N_10127,N_9866,N_9557);
or U10128 (N_10128,N_9500,N_9980);
xnor U10129 (N_10129,N_9676,N_9802);
or U10130 (N_10130,N_9697,N_9913);
xor U10131 (N_10131,N_9664,N_9544);
xnor U10132 (N_10132,N_9868,N_9830);
or U10133 (N_10133,N_9599,N_9624);
nand U10134 (N_10134,N_9981,N_9605);
or U10135 (N_10135,N_9647,N_9806);
nor U10136 (N_10136,N_9724,N_9563);
nor U10137 (N_10137,N_9666,N_9675);
and U10138 (N_10138,N_9654,N_9704);
nor U10139 (N_10139,N_9900,N_9575);
nand U10140 (N_10140,N_9729,N_9606);
nand U10141 (N_10141,N_9847,N_9602);
xnor U10142 (N_10142,N_9852,N_9817);
xor U10143 (N_10143,N_9656,N_9998);
or U10144 (N_10144,N_9954,N_9949);
nand U10145 (N_10145,N_9860,N_9541);
nand U10146 (N_10146,N_9931,N_9756);
nor U10147 (N_10147,N_9622,N_9543);
xnor U10148 (N_10148,N_9809,N_9514);
xor U10149 (N_10149,N_9700,N_9663);
nand U10150 (N_10150,N_9768,N_9649);
and U10151 (N_10151,N_9613,N_9984);
or U10152 (N_10152,N_9584,N_9793);
nor U10153 (N_10153,N_9835,N_9566);
or U10154 (N_10154,N_9712,N_9764);
nor U10155 (N_10155,N_9693,N_9517);
and U10156 (N_10156,N_9516,N_9699);
or U10157 (N_10157,N_9683,N_9978);
or U10158 (N_10158,N_9668,N_9964);
and U10159 (N_10159,N_9530,N_9662);
and U10160 (N_10160,N_9933,N_9726);
xor U10161 (N_10161,N_9796,N_9997);
nand U10162 (N_10162,N_9774,N_9766);
nor U10163 (N_10163,N_9672,N_9625);
xor U10164 (N_10164,N_9761,N_9967);
and U10165 (N_10165,N_9652,N_9629);
nor U10166 (N_10166,N_9937,N_9903);
nor U10167 (N_10167,N_9895,N_9825);
and U10168 (N_10168,N_9524,N_9617);
or U10169 (N_10169,N_9959,N_9739);
or U10170 (N_10170,N_9598,N_9950);
nand U10171 (N_10171,N_9537,N_9594);
xnor U10172 (N_10172,N_9870,N_9713);
nand U10173 (N_10173,N_9550,N_9508);
nor U10174 (N_10174,N_9525,N_9771);
or U10175 (N_10175,N_9845,N_9555);
nand U10176 (N_10176,N_9682,N_9934);
or U10177 (N_10177,N_9691,N_9633);
nand U10178 (N_10178,N_9966,N_9758);
nand U10179 (N_10179,N_9586,N_9642);
nor U10180 (N_10180,N_9927,N_9991);
xor U10181 (N_10181,N_9905,N_9585);
and U10182 (N_10182,N_9922,N_9680);
nor U10183 (N_10183,N_9592,N_9702);
and U10184 (N_10184,N_9839,N_9528);
nor U10185 (N_10185,N_9706,N_9653);
nand U10186 (N_10186,N_9932,N_9917);
nand U10187 (N_10187,N_9899,N_9711);
nand U10188 (N_10188,N_9926,N_9982);
nor U10189 (N_10189,N_9581,N_9973);
nor U10190 (N_10190,N_9781,N_9539);
or U10191 (N_10191,N_9773,N_9958);
xnor U10192 (N_10192,N_9919,N_9526);
and U10193 (N_10193,N_9824,N_9512);
nor U10194 (N_10194,N_9920,N_9751);
and U10195 (N_10195,N_9923,N_9846);
xor U10196 (N_10196,N_9859,N_9609);
nor U10197 (N_10197,N_9874,N_9894);
nor U10198 (N_10198,N_9759,N_9532);
nor U10199 (N_10199,N_9538,N_9871);
and U10200 (N_10200,N_9589,N_9612);
or U10201 (N_10201,N_9677,N_9822);
or U10202 (N_10202,N_9707,N_9800);
and U10203 (N_10203,N_9832,N_9818);
and U10204 (N_10204,N_9748,N_9554);
and U10205 (N_10205,N_9546,N_9534);
xnor U10206 (N_10206,N_9877,N_9787);
nor U10207 (N_10207,N_9597,N_9803);
xor U10208 (N_10208,N_9540,N_9590);
xnor U10209 (N_10209,N_9634,N_9925);
or U10210 (N_10210,N_9935,N_9620);
and U10211 (N_10211,N_9902,N_9658);
or U10212 (N_10212,N_9632,N_9911);
or U10213 (N_10213,N_9938,N_9841);
xor U10214 (N_10214,N_9722,N_9608);
and U10215 (N_10215,N_9785,N_9948);
or U10216 (N_10216,N_9577,N_9757);
and U10217 (N_10217,N_9515,N_9921);
nor U10218 (N_10218,N_9840,N_9705);
xor U10219 (N_10219,N_9985,N_9965);
and U10220 (N_10220,N_9783,N_9671);
and U10221 (N_10221,N_9685,N_9836);
nor U10222 (N_10222,N_9732,N_9892);
nand U10223 (N_10223,N_9674,N_9636);
nand U10224 (N_10224,N_9645,N_9604);
nand U10225 (N_10225,N_9730,N_9513);
xor U10226 (N_10226,N_9762,N_9813);
or U10227 (N_10227,N_9631,N_9842);
and U10228 (N_10228,N_9790,N_9752);
xor U10229 (N_10229,N_9946,N_9673);
nand U10230 (N_10230,N_9501,N_9750);
and U10231 (N_10231,N_9657,N_9821);
or U10232 (N_10232,N_9992,N_9627);
nor U10233 (N_10233,N_9831,N_9854);
or U10234 (N_10234,N_9891,N_9869);
or U10235 (N_10235,N_9812,N_9703);
or U10236 (N_10236,N_9574,N_9944);
or U10237 (N_10237,N_9961,N_9889);
xnor U10238 (N_10238,N_9695,N_9990);
and U10239 (N_10239,N_9565,N_9872);
nand U10240 (N_10240,N_9655,N_9646);
nor U10241 (N_10241,N_9820,N_9881);
or U10242 (N_10242,N_9727,N_9607);
nand U10243 (N_10243,N_9823,N_9986);
xor U10244 (N_10244,N_9914,N_9621);
xor U10245 (N_10245,N_9595,N_9843);
nor U10246 (N_10246,N_9638,N_9789);
nor U10247 (N_10247,N_9898,N_9749);
nand U10248 (N_10248,N_9692,N_9669);
xnor U10249 (N_10249,N_9643,N_9798);
nor U10250 (N_10250,N_9682,N_9995);
or U10251 (N_10251,N_9738,N_9669);
nor U10252 (N_10252,N_9844,N_9796);
nor U10253 (N_10253,N_9506,N_9666);
nand U10254 (N_10254,N_9529,N_9660);
nand U10255 (N_10255,N_9846,N_9876);
and U10256 (N_10256,N_9826,N_9834);
and U10257 (N_10257,N_9576,N_9960);
nor U10258 (N_10258,N_9510,N_9749);
or U10259 (N_10259,N_9830,N_9889);
and U10260 (N_10260,N_9809,N_9530);
nand U10261 (N_10261,N_9746,N_9611);
nand U10262 (N_10262,N_9973,N_9517);
and U10263 (N_10263,N_9775,N_9771);
nor U10264 (N_10264,N_9774,N_9592);
or U10265 (N_10265,N_9792,N_9823);
xnor U10266 (N_10266,N_9617,N_9826);
nor U10267 (N_10267,N_9677,N_9862);
nor U10268 (N_10268,N_9588,N_9691);
and U10269 (N_10269,N_9943,N_9861);
nand U10270 (N_10270,N_9765,N_9825);
nor U10271 (N_10271,N_9557,N_9891);
or U10272 (N_10272,N_9690,N_9929);
nor U10273 (N_10273,N_9788,N_9849);
or U10274 (N_10274,N_9863,N_9904);
or U10275 (N_10275,N_9657,N_9575);
nand U10276 (N_10276,N_9621,N_9808);
or U10277 (N_10277,N_9929,N_9662);
nand U10278 (N_10278,N_9572,N_9815);
nand U10279 (N_10279,N_9675,N_9787);
nand U10280 (N_10280,N_9602,N_9766);
nand U10281 (N_10281,N_9936,N_9504);
or U10282 (N_10282,N_9610,N_9710);
and U10283 (N_10283,N_9938,N_9720);
nor U10284 (N_10284,N_9822,N_9989);
and U10285 (N_10285,N_9902,N_9952);
xor U10286 (N_10286,N_9732,N_9675);
or U10287 (N_10287,N_9601,N_9945);
nor U10288 (N_10288,N_9707,N_9883);
nand U10289 (N_10289,N_9580,N_9796);
or U10290 (N_10290,N_9509,N_9952);
or U10291 (N_10291,N_9765,N_9658);
or U10292 (N_10292,N_9637,N_9738);
nor U10293 (N_10293,N_9627,N_9575);
nor U10294 (N_10294,N_9506,N_9706);
nor U10295 (N_10295,N_9935,N_9963);
and U10296 (N_10296,N_9609,N_9914);
xor U10297 (N_10297,N_9838,N_9806);
xor U10298 (N_10298,N_9798,N_9951);
nand U10299 (N_10299,N_9670,N_9975);
and U10300 (N_10300,N_9587,N_9679);
or U10301 (N_10301,N_9870,N_9578);
xnor U10302 (N_10302,N_9970,N_9822);
nor U10303 (N_10303,N_9874,N_9831);
and U10304 (N_10304,N_9513,N_9789);
nor U10305 (N_10305,N_9813,N_9684);
nor U10306 (N_10306,N_9770,N_9790);
or U10307 (N_10307,N_9629,N_9831);
or U10308 (N_10308,N_9901,N_9610);
nand U10309 (N_10309,N_9677,N_9642);
xnor U10310 (N_10310,N_9647,N_9653);
and U10311 (N_10311,N_9660,N_9597);
xnor U10312 (N_10312,N_9958,N_9942);
or U10313 (N_10313,N_9576,N_9770);
and U10314 (N_10314,N_9629,N_9867);
or U10315 (N_10315,N_9681,N_9958);
and U10316 (N_10316,N_9697,N_9577);
nand U10317 (N_10317,N_9768,N_9512);
and U10318 (N_10318,N_9972,N_9923);
xnor U10319 (N_10319,N_9685,N_9595);
or U10320 (N_10320,N_9693,N_9861);
xnor U10321 (N_10321,N_9581,N_9958);
and U10322 (N_10322,N_9992,N_9739);
and U10323 (N_10323,N_9722,N_9786);
nor U10324 (N_10324,N_9594,N_9786);
xnor U10325 (N_10325,N_9909,N_9620);
nor U10326 (N_10326,N_9591,N_9511);
nor U10327 (N_10327,N_9743,N_9608);
nand U10328 (N_10328,N_9855,N_9536);
and U10329 (N_10329,N_9549,N_9811);
xor U10330 (N_10330,N_9783,N_9977);
nor U10331 (N_10331,N_9763,N_9545);
or U10332 (N_10332,N_9619,N_9639);
nor U10333 (N_10333,N_9541,N_9708);
nand U10334 (N_10334,N_9982,N_9753);
nand U10335 (N_10335,N_9700,N_9968);
xnor U10336 (N_10336,N_9570,N_9749);
nor U10337 (N_10337,N_9697,N_9687);
and U10338 (N_10338,N_9910,N_9915);
and U10339 (N_10339,N_9864,N_9619);
xnor U10340 (N_10340,N_9758,N_9719);
nand U10341 (N_10341,N_9634,N_9708);
xnor U10342 (N_10342,N_9562,N_9711);
or U10343 (N_10343,N_9844,N_9773);
nand U10344 (N_10344,N_9715,N_9774);
nand U10345 (N_10345,N_9918,N_9922);
xor U10346 (N_10346,N_9555,N_9608);
xnor U10347 (N_10347,N_9799,N_9539);
and U10348 (N_10348,N_9949,N_9765);
nor U10349 (N_10349,N_9557,N_9783);
xnor U10350 (N_10350,N_9976,N_9988);
or U10351 (N_10351,N_9755,N_9563);
and U10352 (N_10352,N_9505,N_9657);
xor U10353 (N_10353,N_9630,N_9518);
xnor U10354 (N_10354,N_9649,N_9773);
xnor U10355 (N_10355,N_9934,N_9583);
or U10356 (N_10356,N_9559,N_9730);
xor U10357 (N_10357,N_9719,N_9789);
or U10358 (N_10358,N_9604,N_9783);
or U10359 (N_10359,N_9654,N_9582);
or U10360 (N_10360,N_9919,N_9857);
or U10361 (N_10361,N_9662,N_9665);
nand U10362 (N_10362,N_9869,N_9707);
or U10363 (N_10363,N_9539,N_9996);
xnor U10364 (N_10364,N_9978,N_9571);
nand U10365 (N_10365,N_9715,N_9868);
or U10366 (N_10366,N_9808,N_9708);
nand U10367 (N_10367,N_9969,N_9592);
nand U10368 (N_10368,N_9926,N_9906);
xnor U10369 (N_10369,N_9828,N_9747);
nand U10370 (N_10370,N_9918,N_9711);
or U10371 (N_10371,N_9963,N_9654);
or U10372 (N_10372,N_9982,N_9835);
nor U10373 (N_10373,N_9856,N_9835);
nor U10374 (N_10374,N_9983,N_9713);
nand U10375 (N_10375,N_9965,N_9756);
and U10376 (N_10376,N_9581,N_9967);
nor U10377 (N_10377,N_9728,N_9761);
or U10378 (N_10378,N_9968,N_9621);
xor U10379 (N_10379,N_9692,N_9840);
or U10380 (N_10380,N_9711,N_9732);
and U10381 (N_10381,N_9725,N_9892);
nand U10382 (N_10382,N_9939,N_9586);
or U10383 (N_10383,N_9976,N_9635);
nor U10384 (N_10384,N_9638,N_9718);
and U10385 (N_10385,N_9838,N_9723);
nand U10386 (N_10386,N_9691,N_9551);
and U10387 (N_10387,N_9962,N_9908);
and U10388 (N_10388,N_9698,N_9789);
nor U10389 (N_10389,N_9926,N_9538);
or U10390 (N_10390,N_9718,N_9576);
nand U10391 (N_10391,N_9562,N_9896);
or U10392 (N_10392,N_9904,N_9745);
xor U10393 (N_10393,N_9798,N_9732);
nand U10394 (N_10394,N_9596,N_9520);
xor U10395 (N_10395,N_9623,N_9516);
nand U10396 (N_10396,N_9836,N_9650);
nor U10397 (N_10397,N_9826,N_9662);
xnor U10398 (N_10398,N_9844,N_9761);
xnor U10399 (N_10399,N_9811,N_9658);
nand U10400 (N_10400,N_9883,N_9957);
nand U10401 (N_10401,N_9728,N_9827);
xnor U10402 (N_10402,N_9873,N_9588);
or U10403 (N_10403,N_9784,N_9596);
xor U10404 (N_10404,N_9908,N_9677);
nand U10405 (N_10405,N_9635,N_9871);
nor U10406 (N_10406,N_9917,N_9793);
nand U10407 (N_10407,N_9787,N_9799);
and U10408 (N_10408,N_9763,N_9853);
nand U10409 (N_10409,N_9745,N_9701);
nand U10410 (N_10410,N_9622,N_9915);
nor U10411 (N_10411,N_9641,N_9642);
nand U10412 (N_10412,N_9903,N_9705);
and U10413 (N_10413,N_9724,N_9752);
and U10414 (N_10414,N_9528,N_9841);
xor U10415 (N_10415,N_9990,N_9831);
xnor U10416 (N_10416,N_9532,N_9731);
nor U10417 (N_10417,N_9651,N_9933);
nor U10418 (N_10418,N_9714,N_9875);
or U10419 (N_10419,N_9960,N_9660);
nand U10420 (N_10420,N_9954,N_9697);
nor U10421 (N_10421,N_9857,N_9830);
or U10422 (N_10422,N_9533,N_9742);
or U10423 (N_10423,N_9843,N_9929);
and U10424 (N_10424,N_9892,N_9864);
xnor U10425 (N_10425,N_9657,N_9814);
nand U10426 (N_10426,N_9573,N_9548);
xor U10427 (N_10427,N_9873,N_9737);
nand U10428 (N_10428,N_9599,N_9502);
nand U10429 (N_10429,N_9507,N_9745);
nand U10430 (N_10430,N_9819,N_9955);
xor U10431 (N_10431,N_9702,N_9546);
nand U10432 (N_10432,N_9663,N_9812);
and U10433 (N_10433,N_9674,N_9817);
nor U10434 (N_10434,N_9795,N_9553);
and U10435 (N_10435,N_9854,N_9675);
xor U10436 (N_10436,N_9860,N_9605);
nor U10437 (N_10437,N_9825,N_9500);
or U10438 (N_10438,N_9889,N_9954);
or U10439 (N_10439,N_9912,N_9737);
or U10440 (N_10440,N_9720,N_9894);
or U10441 (N_10441,N_9692,N_9661);
xor U10442 (N_10442,N_9910,N_9877);
nor U10443 (N_10443,N_9553,N_9587);
nand U10444 (N_10444,N_9847,N_9689);
nor U10445 (N_10445,N_9547,N_9834);
nand U10446 (N_10446,N_9970,N_9844);
nor U10447 (N_10447,N_9981,N_9787);
and U10448 (N_10448,N_9865,N_9688);
and U10449 (N_10449,N_9789,N_9940);
nand U10450 (N_10450,N_9692,N_9601);
nand U10451 (N_10451,N_9818,N_9558);
xor U10452 (N_10452,N_9954,N_9797);
and U10453 (N_10453,N_9699,N_9832);
or U10454 (N_10454,N_9587,N_9501);
or U10455 (N_10455,N_9678,N_9805);
xor U10456 (N_10456,N_9733,N_9590);
or U10457 (N_10457,N_9850,N_9564);
nor U10458 (N_10458,N_9733,N_9984);
or U10459 (N_10459,N_9895,N_9539);
nor U10460 (N_10460,N_9701,N_9658);
or U10461 (N_10461,N_9829,N_9862);
nor U10462 (N_10462,N_9916,N_9851);
and U10463 (N_10463,N_9967,N_9660);
nand U10464 (N_10464,N_9934,N_9630);
or U10465 (N_10465,N_9642,N_9634);
xnor U10466 (N_10466,N_9854,N_9747);
nand U10467 (N_10467,N_9955,N_9621);
nor U10468 (N_10468,N_9563,N_9639);
nor U10469 (N_10469,N_9936,N_9502);
nor U10470 (N_10470,N_9598,N_9685);
nor U10471 (N_10471,N_9582,N_9780);
nor U10472 (N_10472,N_9828,N_9917);
nor U10473 (N_10473,N_9623,N_9843);
nor U10474 (N_10474,N_9600,N_9867);
nor U10475 (N_10475,N_9766,N_9594);
xor U10476 (N_10476,N_9564,N_9804);
nor U10477 (N_10477,N_9688,N_9916);
nor U10478 (N_10478,N_9685,N_9716);
xnor U10479 (N_10479,N_9908,N_9749);
and U10480 (N_10480,N_9939,N_9661);
xor U10481 (N_10481,N_9686,N_9894);
xor U10482 (N_10482,N_9815,N_9511);
nand U10483 (N_10483,N_9633,N_9875);
and U10484 (N_10484,N_9947,N_9955);
and U10485 (N_10485,N_9814,N_9988);
or U10486 (N_10486,N_9805,N_9849);
nor U10487 (N_10487,N_9540,N_9934);
nand U10488 (N_10488,N_9764,N_9755);
and U10489 (N_10489,N_9564,N_9927);
xor U10490 (N_10490,N_9941,N_9938);
or U10491 (N_10491,N_9674,N_9977);
nor U10492 (N_10492,N_9879,N_9502);
nand U10493 (N_10493,N_9763,N_9671);
nand U10494 (N_10494,N_9920,N_9510);
nor U10495 (N_10495,N_9638,N_9589);
nand U10496 (N_10496,N_9804,N_9677);
nand U10497 (N_10497,N_9603,N_9715);
or U10498 (N_10498,N_9696,N_9980);
and U10499 (N_10499,N_9818,N_9794);
nand U10500 (N_10500,N_10081,N_10355);
nor U10501 (N_10501,N_10255,N_10436);
xnor U10502 (N_10502,N_10137,N_10219);
nor U10503 (N_10503,N_10031,N_10442);
xor U10504 (N_10504,N_10102,N_10015);
xnor U10505 (N_10505,N_10211,N_10498);
nand U10506 (N_10506,N_10133,N_10095);
nand U10507 (N_10507,N_10462,N_10154);
nand U10508 (N_10508,N_10431,N_10492);
nand U10509 (N_10509,N_10477,N_10068);
nor U10510 (N_10510,N_10340,N_10106);
or U10511 (N_10511,N_10076,N_10495);
or U10512 (N_10512,N_10252,N_10455);
or U10513 (N_10513,N_10062,N_10132);
or U10514 (N_10514,N_10315,N_10411);
nand U10515 (N_10515,N_10329,N_10259);
nand U10516 (N_10516,N_10171,N_10108);
and U10517 (N_10517,N_10275,N_10346);
or U10518 (N_10518,N_10096,N_10342);
xor U10519 (N_10519,N_10307,N_10478);
and U10520 (N_10520,N_10144,N_10395);
nand U10521 (N_10521,N_10080,N_10451);
and U10522 (N_10522,N_10045,N_10088);
nand U10523 (N_10523,N_10217,N_10286);
or U10524 (N_10524,N_10333,N_10011);
nor U10525 (N_10525,N_10248,N_10371);
nand U10526 (N_10526,N_10290,N_10380);
xnor U10527 (N_10527,N_10309,N_10463);
xnor U10528 (N_10528,N_10469,N_10225);
nor U10529 (N_10529,N_10051,N_10231);
or U10530 (N_10530,N_10405,N_10204);
nor U10531 (N_10531,N_10203,N_10196);
xor U10532 (N_10532,N_10141,N_10020);
nand U10533 (N_10533,N_10099,N_10400);
and U10534 (N_10534,N_10409,N_10152);
xnor U10535 (N_10535,N_10341,N_10375);
nand U10536 (N_10536,N_10325,N_10326);
nand U10537 (N_10537,N_10302,N_10454);
nand U10538 (N_10538,N_10033,N_10130);
nor U10539 (N_10539,N_10291,N_10056);
or U10540 (N_10540,N_10456,N_10120);
nor U10541 (N_10541,N_10337,N_10317);
xor U10542 (N_10542,N_10446,N_10321);
nand U10543 (N_10543,N_10364,N_10304);
or U10544 (N_10544,N_10330,N_10287);
nand U10545 (N_10545,N_10403,N_10335);
nor U10546 (N_10546,N_10267,N_10491);
xor U10547 (N_10547,N_10114,N_10336);
or U10548 (N_10548,N_10457,N_10294);
nor U10549 (N_10549,N_10202,N_10303);
or U10550 (N_10550,N_10282,N_10098);
xor U10551 (N_10551,N_10271,N_10301);
or U10552 (N_10552,N_10421,N_10432);
and U10553 (N_10553,N_10151,N_10205);
or U10554 (N_10554,N_10245,N_10097);
nor U10555 (N_10555,N_10209,N_10028);
xor U10556 (N_10556,N_10288,N_10453);
nand U10557 (N_10557,N_10087,N_10420);
nand U10558 (N_10558,N_10393,N_10058);
and U10559 (N_10559,N_10003,N_10496);
xnor U10560 (N_10560,N_10072,N_10254);
nand U10561 (N_10561,N_10361,N_10418);
nor U10562 (N_10562,N_10273,N_10150);
nand U10563 (N_10563,N_10348,N_10377);
xor U10564 (N_10564,N_10048,N_10055);
nand U10565 (N_10565,N_10353,N_10128);
nand U10566 (N_10566,N_10206,N_10401);
and U10567 (N_10567,N_10433,N_10136);
and U10568 (N_10568,N_10366,N_10192);
nor U10569 (N_10569,N_10310,N_10308);
or U10570 (N_10570,N_10201,N_10178);
nor U10571 (N_10571,N_10124,N_10042);
nor U10572 (N_10572,N_10390,N_10032);
and U10573 (N_10573,N_10264,N_10189);
xnor U10574 (N_10574,N_10373,N_10066);
nor U10575 (N_10575,N_10413,N_10283);
xor U10576 (N_10576,N_10212,N_10482);
or U10577 (N_10577,N_10473,N_10163);
nor U10578 (N_10578,N_10193,N_10358);
xor U10579 (N_10579,N_10197,N_10232);
nand U10580 (N_10580,N_10417,N_10018);
and U10581 (N_10581,N_10109,N_10181);
and U10582 (N_10582,N_10448,N_10314);
nand U10583 (N_10583,N_10372,N_10430);
nor U10584 (N_10584,N_10292,N_10170);
xnor U10585 (N_10585,N_10334,N_10316);
nand U10586 (N_10586,N_10265,N_10021);
and U10587 (N_10587,N_10157,N_10155);
or U10588 (N_10588,N_10458,N_10117);
or U10589 (N_10589,N_10253,N_10161);
nor U10590 (N_10590,N_10470,N_10240);
nor U10591 (N_10591,N_10429,N_10338);
and U10592 (N_10592,N_10001,N_10391);
and U10593 (N_10593,N_10422,N_10261);
or U10594 (N_10594,N_10350,N_10063);
nor U10595 (N_10595,N_10268,N_10044);
nor U10596 (N_10596,N_10298,N_10179);
nor U10597 (N_10597,N_10386,N_10075);
nor U10598 (N_10598,N_10370,N_10440);
nand U10599 (N_10599,N_10323,N_10296);
and U10600 (N_10600,N_10138,N_10388);
nor U10601 (N_10601,N_10183,N_10119);
xor U10602 (N_10602,N_10121,N_10069);
xnor U10603 (N_10603,N_10200,N_10419);
or U10604 (N_10604,N_10262,N_10194);
nor U10605 (N_10605,N_10452,N_10030);
nor U10606 (N_10606,N_10297,N_10399);
or U10607 (N_10607,N_10057,N_10199);
or U10608 (N_10608,N_10289,N_10177);
and U10609 (N_10609,N_10332,N_10378);
or U10610 (N_10610,N_10357,N_10047);
or U10611 (N_10611,N_10131,N_10093);
and U10612 (N_10612,N_10035,N_10083);
xnor U10613 (N_10613,N_10276,N_10019);
nor U10614 (N_10614,N_10347,N_10184);
nand U10615 (N_10615,N_10443,N_10174);
and U10616 (N_10616,N_10312,N_10230);
and U10617 (N_10617,N_10190,N_10459);
xor U10618 (N_10618,N_10414,N_10236);
nand U10619 (N_10619,N_10143,N_10071);
nand U10620 (N_10620,N_10423,N_10159);
nor U10621 (N_10621,N_10256,N_10165);
xor U10622 (N_10622,N_10300,N_10319);
nor U10623 (N_10623,N_10382,N_10438);
xnor U10624 (N_10624,N_10016,N_10490);
nand U10625 (N_10625,N_10284,N_10173);
and U10626 (N_10626,N_10249,N_10160);
xor U10627 (N_10627,N_10392,N_10424);
and U10628 (N_10628,N_10369,N_10367);
and U10629 (N_10629,N_10147,N_10295);
and U10630 (N_10630,N_10127,N_10241);
nand U10631 (N_10631,N_10322,N_10339);
nand U10632 (N_10632,N_10101,N_10243);
xor U10633 (N_10633,N_10140,N_10135);
nand U10634 (N_10634,N_10260,N_10054);
or U10635 (N_10635,N_10280,N_10100);
nor U10636 (N_10636,N_10084,N_10029);
or U10637 (N_10637,N_10486,N_10356);
or U10638 (N_10638,N_10331,N_10113);
nor U10639 (N_10639,N_10238,N_10277);
nand U10640 (N_10640,N_10354,N_10207);
nand U10641 (N_10641,N_10049,N_10387);
nor U10642 (N_10642,N_10471,N_10352);
xnor U10643 (N_10643,N_10077,N_10213);
nor U10644 (N_10644,N_10434,N_10406);
xor U10645 (N_10645,N_10461,N_10060);
nand U10646 (N_10646,N_10416,N_10168);
and U10647 (N_10647,N_10092,N_10006);
nand U10648 (N_10648,N_10224,N_10475);
nor U10649 (N_10649,N_10318,N_10182);
and U10650 (N_10650,N_10198,N_10176);
or U10651 (N_10651,N_10125,N_10464);
nand U10652 (N_10652,N_10126,N_10123);
nand U10653 (N_10653,N_10220,N_10191);
xor U10654 (N_10654,N_10383,N_10266);
and U10655 (N_10655,N_10129,N_10234);
or U10656 (N_10656,N_10112,N_10064);
or U10657 (N_10657,N_10269,N_10024);
or U10658 (N_10658,N_10164,N_10142);
nor U10659 (N_10659,N_10368,N_10246);
nor U10660 (N_10660,N_10017,N_10476);
nor U10661 (N_10661,N_10270,N_10105);
nand U10662 (N_10662,N_10065,N_10285);
xor U10663 (N_10663,N_10214,N_10376);
nand U10664 (N_10664,N_10404,N_10484);
and U10665 (N_10665,N_10328,N_10474);
xnor U10666 (N_10666,N_10235,N_10293);
nand U10667 (N_10667,N_10480,N_10445);
nor U10668 (N_10668,N_10094,N_10145);
xnor U10669 (N_10669,N_10002,N_10188);
nor U10670 (N_10670,N_10233,N_10449);
or U10671 (N_10671,N_10494,N_10435);
nand U10672 (N_10672,N_10208,N_10359);
or U10673 (N_10673,N_10483,N_10043);
and U10674 (N_10674,N_10122,N_10110);
or U10675 (N_10675,N_10465,N_10036);
nand U10676 (N_10676,N_10493,N_10311);
and U10677 (N_10677,N_10082,N_10360);
xnor U10678 (N_10678,N_10008,N_10180);
xor U10679 (N_10679,N_10229,N_10365);
and U10680 (N_10680,N_10023,N_10085);
nor U10681 (N_10681,N_10223,N_10488);
nand U10682 (N_10682,N_10439,N_10195);
or U10683 (N_10683,N_10251,N_10441);
and U10684 (N_10684,N_10007,N_10038);
xnor U10685 (N_10685,N_10408,N_10379);
nand U10686 (N_10686,N_10070,N_10107);
and U10687 (N_10687,N_10139,N_10073);
nand U10688 (N_10688,N_10226,N_10381);
nor U10689 (N_10689,N_10103,N_10467);
and U10690 (N_10690,N_10010,N_10116);
or U10691 (N_10691,N_10022,N_10450);
or U10692 (N_10692,N_10175,N_10444);
or U10693 (N_10693,N_10079,N_10374);
or U10694 (N_10694,N_10447,N_10000);
xor U10695 (N_10695,N_10258,N_10215);
and U10696 (N_10696,N_10086,N_10059);
or U10697 (N_10697,N_10025,N_10146);
nand U10698 (N_10698,N_10153,N_10428);
xnor U10699 (N_10699,N_10009,N_10239);
nand U10700 (N_10700,N_10362,N_10250);
nand U10701 (N_10701,N_10320,N_10013);
nand U10702 (N_10702,N_10345,N_10472);
or U10703 (N_10703,N_10158,N_10394);
nand U10704 (N_10704,N_10426,N_10104);
or U10705 (N_10705,N_10040,N_10274);
nand U10706 (N_10706,N_10039,N_10427);
xor U10707 (N_10707,N_10499,N_10156);
and U10708 (N_10708,N_10415,N_10487);
or U10709 (N_10709,N_10410,N_10050);
or U10710 (N_10710,N_10384,N_10244);
nor U10711 (N_10711,N_10037,N_10041);
nand U10712 (N_10712,N_10412,N_10272);
or U10713 (N_10713,N_10166,N_10460);
and U10714 (N_10714,N_10227,N_10489);
nor U10715 (N_10715,N_10004,N_10061);
and U10716 (N_10716,N_10149,N_10026);
or U10717 (N_10717,N_10027,N_10034);
nor U10718 (N_10718,N_10118,N_10324);
or U10719 (N_10719,N_10185,N_10407);
nor U10720 (N_10720,N_10005,N_10306);
nand U10721 (N_10721,N_10257,N_10111);
xnor U10722 (N_10722,N_10278,N_10221);
nor U10723 (N_10723,N_10237,N_10468);
and U10724 (N_10724,N_10305,N_10090);
xor U10725 (N_10725,N_10279,N_10115);
and U10726 (N_10726,N_10344,N_10351);
xnor U10727 (N_10727,N_10052,N_10397);
and U10728 (N_10728,N_10363,N_10385);
and U10729 (N_10729,N_10014,N_10481);
xor U10730 (N_10730,N_10343,N_10053);
nor U10731 (N_10731,N_10299,N_10263);
nand U10732 (N_10732,N_10186,N_10216);
and U10733 (N_10733,N_10497,N_10479);
or U10734 (N_10734,N_10425,N_10228);
nand U10735 (N_10735,N_10172,N_10327);
nor U10736 (N_10736,N_10046,N_10167);
nand U10737 (N_10737,N_10169,N_10218);
and U10738 (N_10738,N_10281,N_10466);
nor U10739 (N_10739,N_10210,N_10134);
and U10740 (N_10740,N_10091,N_10012);
nand U10741 (N_10741,N_10078,N_10437);
and U10742 (N_10742,N_10148,N_10242);
nand U10743 (N_10743,N_10222,N_10402);
xor U10744 (N_10744,N_10389,N_10074);
nand U10745 (N_10745,N_10398,N_10349);
xnor U10746 (N_10746,N_10247,N_10187);
nor U10747 (N_10747,N_10396,N_10067);
xnor U10748 (N_10748,N_10162,N_10089);
or U10749 (N_10749,N_10313,N_10485);
nand U10750 (N_10750,N_10101,N_10231);
and U10751 (N_10751,N_10160,N_10345);
xor U10752 (N_10752,N_10186,N_10083);
xnor U10753 (N_10753,N_10317,N_10175);
or U10754 (N_10754,N_10008,N_10056);
or U10755 (N_10755,N_10044,N_10199);
or U10756 (N_10756,N_10299,N_10470);
nor U10757 (N_10757,N_10191,N_10146);
or U10758 (N_10758,N_10492,N_10129);
and U10759 (N_10759,N_10417,N_10180);
or U10760 (N_10760,N_10074,N_10098);
xor U10761 (N_10761,N_10432,N_10245);
nor U10762 (N_10762,N_10249,N_10278);
or U10763 (N_10763,N_10269,N_10013);
xor U10764 (N_10764,N_10406,N_10413);
or U10765 (N_10765,N_10101,N_10429);
nor U10766 (N_10766,N_10341,N_10113);
xnor U10767 (N_10767,N_10121,N_10453);
and U10768 (N_10768,N_10303,N_10044);
and U10769 (N_10769,N_10388,N_10080);
and U10770 (N_10770,N_10363,N_10447);
nand U10771 (N_10771,N_10446,N_10126);
xnor U10772 (N_10772,N_10456,N_10436);
nor U10773 (N_10773,N_10354,N_10438);
and U10774 (N_10774,N_10333,N_10444);
nor U10775 (N_10775,N_10452,N_10261);
nor U10776 (N_10776,N_10090,N_10146);
xnor U10777 (N_10777,N_10374,N_10446);
or U10778 (N_10778,N_10214,N_10079);
and U10779 (N_10779,N_10047,N_10314);
xor U10780 (N_10780,N_10133,N_10250);
xnor U10781 (N_10781,N_10314,N_10449);
and U10782 (N_10782,N_10422,N_10200);
nand U10783 (N_10783,N_10379,N_10483);
xnor U10784 (N_10784,N_10219,N_10281);
nor U10785 (N_10785,N_10333,N_10215);
nand U10786 (N_10786,N_10145,N_10446);
xnor U10787 (N_10787,N_10271,N_10210);
and U10788 (N_10788,N_10266,N_10057);
or U10789 (N_10789,N_10460,N_10023);
and U10790 (N_10790,N_10134,N_10075);
xnor U10791 (N_10791,N_10014,N_10085);
or U10792 (N_10792,N_10063,N_10107);
nor U10793 (N_10793,N_10039,N_10475);
xor U10794 (N_10794,N_10264,N_10498);
xor U10795 (N_10795,N_10274,N_10392);
and U10796 (N_10796,N_10368,N_10343);
xnor U10797 (N_10797,N_10471,N_10485);
xnor U10798 (N_10798,N_10248,N_10337);
nor U10799 (N_10799,N_10104,N_10427);
nand U10800 (N_10800,N_10323,N_10128);
xnor U10801 (N_10801,N_10336,N_10235);
nand U10802 (N_10802,N_10485,N_10393);
nor U10803 (N_10803,N_10003,N_10108);
nand U10804 (N_10804,N_10475,N_10385);
xor U10805 (N_10805,N_10468,N_10273);
nor U10806 (N_10806,N_10203,N_10492);
xor U10807 (N_10807,N_10475,N_10130);
nand U10808 (N_10808,N_10097,N_10053);
nand U10809 (N_10809,N_10252,N_10099);
nand U10810 (N_10810,N_10432,N_10053);
nand U10811 (N_10811,N_10243,N_10392);
nand U10812 (N_10812,N_10107,N_10412);
nand U10813 (N_10813,N_10488,N_10390);
xor U10814 (N_10814,N_10463,N_10483);
or U10815 (N_10815,N_10485,N_10397);
or U10816 (N_10816,N_10282,N_10210);
xor U10817 (N_10817,N_10495,N_10144);
or U10818 (N_10818,N_10347,N_10386);
or U10819 (N_10819,N_10410,N_10163);
or U10820 (N_10820,N_10177,N_10365);
xor U10821 (N_10821,N_10466,N_10268);
xor U10822 (N_10822,N_10324,N_10271);
xnor U10823 (N_10823,N_10422,N_10476);
and U10824 (N_10824,N_10432,N_10024);
nor U10825 (N_10825,N_10126,N_10191);
and U10826 (N_10826,N_10174,N_10324);
nor U10827 (N_10827,N_10375,N_10207);
nor U10828 (N_10828,N_10475,N_10078);
nand U10829 (N_10829,N_10318,N_10034);
nand U10830 (N_10830,N_10353,N_10222);
or U10831 (N_10831,N_10412,N_10330);
xor U10832 (N_10832,N_10241,N_10279);
nand U10833 (N_10833,N_10157,N_10078);
and U10834 (N_10834,N_10296,N_10420);
nand U10835 (N_10835,N_10235,N_10205);
nor U10836 (N_10836,N_10077,N_10033);
or U10837 (N_10837,N_10470,N_10347);
or U10838 (N_10838,N_10051,N_10353);
and U10839 (N_10839,N_10103,N_10358);
nand U10840 (N_10840,N_10082,N_10445);
nor U10841 (N_10841,N_10339,N_10384);
xnor U10842 (N_10842,N_10283,N_10222);
nand U10843 (N_10843,N_10176,N_10277);
xnor U10844 (N_10844,N_10124,N_10099);
or U10845 (N_10845,N_10241,N_10036);
xnor U10846 (N_10846,N_10486,N_10362);
nor U10847 (N_10847,N_10068,N_10232);
nor U10848 (N_10848,N_10356,N_10321);
and U10849 (N_10849,N_10279,N_10495);
nand U10850 (N_10850,N_10073,N_10318);
xor U10851 (N_10851,N_10466,N_10115);
and U10852 (N_10852,N_10019,N_10420);
or U10853 (N_10853,N_10398,N_10317);
nor U10854 (N_10854,N_10314,N_10261);
or U10855 (N_10855,N_10025,N_10095);
xnor U10856 (N_10856,N_10498,N_10047);
and U10857 (N_10857,N_10235,N_10247);
or U10858 (N_10858,N_10334,N_10206);
nor U10859 (N_10859,N_10024,N_10071);
nand U10860 (N_10860,N_10462,N_10351);
nor U10861 (N_10861,N_10154,N_10157);
or U10862 (N_10862,N_10169,N_10484);
and U10863 (N_10863,N_10224,N_10370);
and U10864 (N_10864,N_10157,N_10165);
nor U10865 (N_10865,N_10336,N_10152);
nand U10866 (N_10866,N_10063,N_10292);
nand U10867 (N_10867,N_10081,N_10173);
xor U10868 (N_10868,N_10433,N_10112);
or U10869 (N_10869,N_10078,N_10252);
xor U10870 (N_10870,N_10252,N_10427);
or U10871 (N_10871,N_10365,N_10426);
nand U10872 (N_10872,N_10374,N_10134);
nand U10873 (N_10873,N_10126,N_10205);
nor U10874 (N_10874,N_10039,N_10403);
and U10875 (N_10875,N_10171,N_10014);
or U10876 (N_10876,N_10499,N_10466);
and U10877 (N_10877,N_10463,N_10315);
nor U10878 (N_10878,N_10401,N_10204);
nor U10879 (N_10879,N_10413,N_10268);
and U10880 (N_10880,N_10317,N_10147);
xnor U10881 (N_10881,N_10188,N_10121);
nand U10882 (N_10882,N_10117,N_10254);
nor U10883 (N_10883,N_10314,N_10100);
or U10884 (N_10884,N_10074,N_10426);
nand U10885 (N_10885,N_10076,N_10009);
nor U10886 (N_10886,N_10083,N_10256);
or U10887 (N_10887,N_10479,N_10225);
and U10888 (N_10888,N_10066,N_10423);
or U10889 (N_10889,N_10241,N_10299);
and U10890 (N_10890,N_10416,N_10273);
nor U10891 (N_10891,N_10398,N_10358);
xnor U10892 (N_10892,N_10148,N_10000);
nor U10893 (N_10893,N_10043,N_10006);
xnor U10894 (N_10894,N_10076,N_10144);
or U10895 (N_10895,N_10304,N_10329);
and U10896 (N_10896,N_10345,N_10077);
nand U10897 (N_10897,N_10254,N_10220);
nor U10898 (N_10898,N_10048,N_10249);
and U10899 (N_10899,N_10291,N_10157);
and U10900 (N_10900,N_10188,N_10283);
and U10901 (N_10901,N_10011,N_10026);
xor U10902 (N_10902,N_10251,N_10296);
nor U10903 (N_10903,N_10092,N_10425);
xnor U10904 (N_10904,N_10288,N_10258);
nor U10905 (N_10905,N_10267,N_10424);
nor U10906 (N_10906,N_10469,N_10193);
nand U10907 (N_10907,N_10187,N_10217);
and U10908 (N_10908,N_10392,N_10327);
or U10909 (N_10909,N_10103,N_10252);
nor U10910 (N_10910,N_10052,N_10086);
nand U10911 (N_10911,N_10453,N_10367);
nand U10912 (N_10912,N_10163,N_10037);
nor U10913 (N_10913,N_10266,N_10019);
or U10914 (N_10914,N_10120,N_10399);
or U10915 (N_10915,N_10479,N_10297);
xor U10916 (N_10916,N_10078,N_10381);
or U10917 (N_10917,N_10469,N_10472);
nand U10918 (N_10918,N_10289,N_10208);
nand U10919 (N_10919,N_10335,N_10364);
xor U10920 (N_10920,N_10184,N_10434);
xor U10921 (N_10921,N_10055,N_10128);
nor U10922 (N_10922,N_10278,N_10065);
xor U10923 (N_10923,N_10049,N_10291);
nand U10924 (N_10924,N_10488,N_10371);
nor U10925 (N_10925,N_10203,N_10123);
nand U10926 (N_10926,N_10014,N_10178);
nor U10927 (N_10927,N_10114,N_10463);
or U10928 (N_10928,N_10149,N_10090);
nand U10929 (N_10929,N_10166,N_10478);
xor U10930 (N_10930,N_10242,N_10036);
nor U10931 (N_10931,N_10008,N_10192);
or U10932 (N_10932,N_10222,N_10173);
xnor U10933 (N_10933,N_10176,N_10064);
and U10934 (N_10934,N_10125,N_10036);
xor U10935 (N_10935,N_10044,N_10058);
or U10936 (N_10936,N_10120,N_10380);
xnor U10937 (N_10937,N_10107,N_10443);
nor U10938 (N_10938,N_10345,N_10377);
and U10939 (N_10939,N_10329,N_10244);
and U10940 (N_10940,N_10380,N_10092);
and U10941 (N_10941,N_10301,N_10361);
nor U10942 (N_10942,N_10289,N_10479);
and U10943 (N_10943,N_10451,N_10182);
and U10944 (N_10944,N_10172,N_10268);
nand U10945 (N_10945,N_10236,N_10295);
nand U10946 (N_10946,N_10376,N_10052);
xor U10947 (N_10947,N_10275,N_10270);
and U10948 (N_10948,N_10439,N_10438);
or U10949 (N_10949,N_10055,N_10346);
nor U10950 (N_10950,N_10065,N_10410);
nand U10951 (N_10951,N_10497,N_10395);
nand U10952 (N_10952,N_10339,N_10414);
nand U10953 (N_10953,N_10114,N_10457);
or U10954 (N_10954,N_10490,N_10160);
or U10955 (N_10955,N_10006,N_10197);
nor U10956 (N_10956,N_10073,N_10163);
xnor U10957 (N_10957,N_10299,N_10104);
and U10958 (N_10958,N_10096,N_10213);
or U10959 (N_10959,N_10362,N_10471);
or U10960 (N_10960,N_10048,N_10262);
nor U10961 (N_10961,N_10413,N_10272);
xor U10962 (N_10962,N_10023,N_10372);
or U10963 (N_10963,N_10177,N_10362);
nand U10964 (N_10964,N_10126,N_10113);
and U10965 (N_10965,N_10487,N_10176);
and U10966 (N_10966,N_10319,N_10028);
nor U10967 (N_10967,N_10064,N_10146);
and U10968 (N_10968,N_10036,N_10244);
nor U10969 (N_10969,N_10411,N_10043);
xnor U10970 (N_10970,N_10155,N_10020);
or U10971 (N_10971,N_10372,N_10031);
nand U10972 (N_10972,N_10070,N_10144);
nand U10973 (N_10973,N_10302,N_10220);
and U10974 (N_10974,N_10380,N_10071);
nor U10975 (N_10975,N_10429,N_10131);
and U10976 (N_10976,N_10274,N_10128);
nor U10977 (N_10977,N_10059,N_10375);
and U10978 (N_10978,N_10111,N_10062);
nand U10979 (N_10979,N_10104,N_10402);
and U10980 (N_10980,N_10466,N_10493);
nand U10981 (N_10981,N_10014,N_10400);
or U10982 (N_10982,N_10460,N_10102);
and U10983 (N_10983,N_10023,N_10333);
xnor U10984 (N_10984,N_10096,N_10132);
xnor U10985 (N_10985,N_10495,N_10080);
nand U10986 (N_10986,N_10059,N_10069);
xor U10987 (N_10987,N_10005,N_10437);
and U10988 (N_10988,N_10079,N_10399);
nor U10989 (N_10989,N_10322,N_10094);
and U10990 (N_10990,N_10184,N_10269);
xor U10991 (N_10991,N_10491,N_10061);
nand U10992 (N_10992,N_10038,N_10355);
and U10993 (N_10993,N_10264,N_10107);
nor U10994 (N_10994,N_10281,N_10098);
nand U10995 (N_10995,N_10374,N_10332);
nor U10996 (N_10996,N_10096,N_10236);
xnor U10997 (N_10997,N_10028,N_10383);
nand U10998 (N_10998,N_10277,N_10099);
xor U10999 (N_10999,N_10046,N_10187);
or U11000 (N_11000,N_10663,N_10604);
and U11001 (N_11001,N_10632,N_10820);
xor U11002 (N_11002,N_10550,N_10584);
nand U11003 (N_11003,N_10645,N_10573);
xor U11004 (N_11004,N_10644,N_10588);
nand U11005 (N_11005,N_10967,N_10574);
xor U11006 (N_11006,N_10891,N_10672);
xor U11007 (N_11007,N_10850,N_10762);
xor U11008 (N_11008,N_10991,N_10928);
or U11009 (N_11009,N_10887,N_10923);
nand U11010 (N_11010,N_10936,N_10767);
nand U11011 (N_11011,N_10543,N_10565);
or U11012 (N_11012,N_10782,N_10873);
xor U11013 (N_11013,N_10610,N_10987);
and U11014 (N_11014,N_10770,N_10680);
nor U11015 (N_11015,N_10559,N_10970);
nand U11016 (N_11016,N_10557,N_10599);
or U11017 (N_11017,N_10611,N_10654);
or U11018 (N_11018,N_10979,N_10552);
and U11019 (N_11019,N_10913,N_10576);
or U11020 (N_11020,N_10867,N_10640);
nand U11021 (N_11021,N_10638,N_10854);
xor U11022 (N_11022,N_10798,N_10882);
nor U11023 (N_11023,N_10839,N_10947);
nand U11024 (N_11024,N_10833,N_10639);
nand U11025 (N_11025,N_10617,N_10514);
nand U11026 (N_11026,N_10577,N_10907);
nand U11027 (N_11027,N_10908,N_10501);
xor U11028 (N_11028,N_10622,N_10626);
and U11029 (N_11029,N_10972,N_10558);
nor U11030 (N_11030,N_10684,N_10919);
and U11031 (N_11031,N_10927,N_10821);
or U11032 (N_11032,N_10720,N_10951);
nand U11033 (N_11033,N_10546,N_10834);
xor U11034 (N_11034,N_10661,N_10615);
nor U11035 (N_11035,N_10875,N_10747);
or U11036 (N_11036,N_10563,N_10773);
xnor U11037 (N_11037,N_10502,N_10929);
and U11038 (N_11038,N_10825,N_10667);
nor U11039 (N_11039,N_10731,N_10556);
nor U11040 (N_11040,N_10709,N_10505);
nor U11041 (N_11041,N_10549,N_10669);
xnor U11042 (N_11042,N_10816,N_10539);
nor U11043 (N_11043,N_10740,N_10902);
or U11044 (N_11044,N_10636,N_10569);
xor U11045 (N_11045,N_10959,N_10695);
xnor U11046 (N_11046,N_10790,N_10560);
or U11047 (N_11047,N_10724,N_10796);
nor U11048 (N_11048,N_10692,N_10792);
xor U11049 (N_11049,N_10789,N_10500);
xor U11050 (N_11050,N_10884,N_10838);
nor U11051 (N_11051,N_10630,N_10534);
xor U11052 (N_11052,N_10718,N_10736);
or U11053 (N_11053,N_10733,N_10517);
or U11054 (N_11054,N_10957,N_10542);
xnor U11055 (N_11055,N_10705,N_10993);
and U11056 (N_11056,N_10671,N_10749);
xnor U11057 (N_11057,N_10859,N_10656);
nand U11058 (N_11058,N_10879,N_10723);
and U11059 (N_11059,N_10739,N_10688);
nor U11060 (N_11060,N_10968,N_10949);
and U11061 (N_11061,N_10944,N_10570);
or U11062 (N_11062,N_10912,N_10594);
nand U11063 (N_11063,N_10541,N_10600);
or U11064 (N_11064,N_10781,N_10930);
nand U11065 (N_11065,N_10682,N_10730);
nand U11066 (N_11066,N_10532,N_10948);
nor U11067 (N_11067,N_10862,N_10870);
nor U11068 (N_11068,N_10886,N_10710);
nand U11069 (N_11069,N_10809,N_10974);
and U11070 (N_11070,N_10978,N_10677);
and U11071 (N_11071,N_10648,N_10634);
and U11072 (N_11072,N_10612,N_10871);
nand U11073 (N_11073,N_10826,N_10900);
and U11074 (N_11074,N_10575,N_10535);
or U11075 (N_11075,N_10659,N_10727);
xor U11076 (N_11076,N_10614,N_10771);
nand U11077 (N_11077,N_10605,N_10571);
xnor U11078 (N_11078,N_10503,N_10732);
nand U11079 (N_11079,N_10608,N_10803);
or U11080 (N_11080,N_10738,N_10868);
nor U11081 (N_11081,N_10544,N_10775);
nand U11082 (N_11082,N_10765,N_10579);
nor U11083 (N_11083,N_10980,N_10960);
nand U11084 (N_11084,N_10704,N_10872);
nor U11085 (N_11085,N_10819,N_10774);
and U11086 (N_11086,N_10830,N_10531);
and U11087 (N_11087,N_10931,N_10547);
nand U11088 (N_11088,N_10601,N_10642);
or U11089 (N_11089,N_10933,N_10598);
xor U11090 (N_11090,N_10937,N_10863);
and U11091 (N_11091,N_10609,N_10787);
and U11092 (N_11092,N_10603,N_10679);
xnor U11093 (N_11093,N_10842,N_10580);
nand U11094 (N_11094,N_10624,N_10811);
nand U11095 (N_11095,N_10898,N_10866);
nand U11096 (N_11096,N_10805,N_10742);
or U11097 (N_11097,N_10697,N_10986);
nand U11098 (N_11098,N_10904,N_10845);
nand U11099 (N_11099,N_10650,N_10917);
nand U11100 (N_11100,N_10646,N_10916);
nand U11101 (N_11101,N_10751,N_10647);
xnor U11102 (N_11102,N_10795,N_10651);
xor U11103 (N_11103,N_10837,N_10613);
or U11104 (N_11104,N_10529,N_10606);
nor U11105 (N_11105,N_10776,N_10969);
xnor U11106 (N_11106,N_10797,N_10523);
and U11107 (N_11107,N_10851,N_10956);
or U11108 (N_11108,N_10880,N_10513);
and U11109 (N_11109,N_10566,N_10548);
or U11110 (N_11110,N_10800,N_10701);
nor U11111 (N_11111,N_10623,N_10681);
and U11112 (N_11112,N_10678,N_10920);
or U11113 (N_11113,N_10629,N_10725);
and U11114 (N_11114,N_10888,N_10625);
or U11115 (N_11115,N_10585,N_10766);
nand U11116 (N_11116,N_10719,N_10707);
nor U11117 (N_11117,N_10621,N_10988);
xor U11118 (N_11118,N_10832,N_10618);
and U11119 (N_11119,N_10779,N_10761);
nand U11120 (N_11120,N_10652,N_10509);
or U11121 (N_11121,N_10637,N_10561);
nand U11122 (N_11122,N_10855,N_10756);
nand U11123 (N_11123,N_10712,N_10746);
nand U11124 (N_11124,N_10966,N_10828);
xor U11125 (N_11125,N_10990,N_10734);
or U11126 (N_11126,N_10844,N_10856);
nor U11127 (N_11127,N_10586,N_10932);
or U11128 (N_11128,N_10938,N_10939);
nor U11129 (N_11129,N_10780,N_10649);
or U11130 (N_11130,N_10943,N_10665);
and U11131 (N_11131,N_10578,N_10537);
and U11132 (N_11132,N_10946,N_10883);
nor U11133 (N_11133,N_10591,N_10530);
nand U11134 (N_11134,N_10914,N_10668);
nand U11135 (N_11135,N_10675,N_10769);
and U11136 (N_11136,N_10953,N_10962);
nand U11137 (N_11137,N_10894,N_10568);
nor U11138 (N_11138,N_10587,N_10999);
nand U11139 (N_11139,N_10683,N_10996);
xor U11140 (N_11140,N_10596,N_10759);
xnor U11141 (N_11141,N_10722,N_10744);
nand U11142 (N_11142,N_10903,N_10975);
and U11143 (N_11143,N_10983,N_10597);
xor U11144 (N_11144,N_10674,N_10890);
nand U11145 (N_11145,N_10522,N_10687);
nor U11146 (N_11146,N_10905,N_10940);
or U11147 (N_11147,N_10686,N_10799);
and U11148 (N_11148,N_10673,N_10961);
and U11149 (N_11149,N_10909,N_10950);
nand U11150 (N_11150,N_10997,N_10892);
nand U11151 (N_11151,N_10555,N_10864);
xnor U11152 (N_11152,N_10858,N_10926);
nand U11153 (N_11153,N_10620,N_10602);
xnor U11154 (N_11154,N_10525,N_10516);
or U11155 (N_11155,N_10985,N_10728);
or U11156 (N_11156,N_10847,N_10589);
nor U11157 (N_11157,N_10976,N_10527);
nor U11158 (N_11158,N_10818,N_10593);
nand U11159 (N_11159,N_10802,N_10924);
or U11160 (N_11160,N_10595,N_10757);
xnor U11161 (N_11161,N_10786,N_10753);
and U11162 (N_11162,N_10590,N_10785);
and U11163 (N_11163,N_10876,N_10752);
xor U11164 (N_11164,N_10982,N_10981);
and U11165 (N_11165,N_10817,N_10504);
and U11166 (N_11166,N_10965,N_10696);
or U11167 (N_11167,N_10693,N_10760);
nor U11168 (N_11168,N_10843,N_10783);
nor U11169 (N_11169,N_10526,N_10750);
xnor U11170 (N_11170,N_10690,N_10653);
nand U11171 (N_11171,N_10564,N_10804);
xnor U11172 (N_11172,N_10524,N_10538);
nor U11173 (N_11173,N_10881,N_10852);
xnor U11174 (N_11174,N_10942,N_10758);
nor U11175 (N_11175,N_10554,N_10694);
and U11176 (N_11176,N_10754,N_10941);
or U11177 (N_11177,N_10829,N_10910);
nand U11178 (N_11178,N_10860,N_10801);
and U11179 (N_11179,N_10810,N_10553);
and U11180 (N_11180,N_10921,N_10995);
and U11181 (N_11181,N_10893,N_10567);
and U11182 (N_11182,N_10840,N_10657);
nand U11183 (N_11183,N_10635,N_10735);
and U11184 (N_11184,N_10813,N_10631);
xnor U11185 (N_11185,N_10633,N_10715);
and U11186 (N_11186,N_10964,N_10521);
nor U11187 (N_11187,N_10741,N_10592);
nor U11188 (N_11188,N_10791,N_10743);
or U11189 (N_11189,N_10877,N_10583);
and U11190 (N_11190,N_10662,N_10835);
xnor U11191 (N_11191,N_10551,N_10520);
nand U11192 (N_11192,N_10691,N_10831);
nand U11193 (N_11193,N_10515,N_10655);
nor U11194 (N_11194,N_10510,N_10628);
or U11195 (N_11195,N_10992,N_10998);
or U11196 (N_11196,N_10807,N_10528);
xor U11197 (N_11197,N_10643,N_10853);
xor U11198 (N_11198,N_10676,N_10827);
nand U11199 (N_11199,N_10699,N_10562);
nor U11200 (N_11200,N_10607,N_10519);
or U11201 (N_11201,N_10954,N_10660);
xnor U11202 (N_11202,N_10973,N_10512);
nor U11203 (N_11203,N_10989,N_10714);
and U11204 (N_11204,N_10945,N_10878);
nor U11205 (N_11205,N_10717,N_10806);
nand U11206 (N_11206,N_10689,N_10616);
nor U11207 (N_11207,N_10778,N_10963);
or U11208 (N_11208,N_10822,N_10984);
nand U11209 (N_11209,N_10511,N_10971);
nor U11210 (N_11210,N_10506,N_10823);
or U11211 (N_11211,N_10934,N_10627);
or U11212 (N_11212,N_10777,N_10658);
or U11213 (N_11213,N_10619,N_10918);
nand U11214 (N_11214,N_10582,N_10906);
or U11215 (N_11215,N_10540,N_10729);
or U11216 (N_11216,N_10533,N_10935);
or U11217 (N_11217,N_10706,N_10536);
xnor U11218 (N_11218,N_10713,N_10849);
nor U11219 (N_11219,N_10925,N_10885);
xor U11220 (N_11220,N_10793,N_10812);
nand U11221 (N_11221,N_10664,N_10572);
or U11222 (N_11222,N_10716,N_10922);
and U11223 (N_11223,N_10952,N_10841);
and U11224 (N_11224,N_10915,N_10698);
xor U11225 (N_11225,N_10895,N_10702);
and U11226 (N_11226,N_10755,N_10768);
and U11227 (N_11227,N_10846,N_10824);
xor U11228 (N_11228,N_10721,N_10977);
and U11229 (N_11229,N_10518,N_10703);
and U11230 (N_11230,N_10911,N_10737);
nand U11231 (N_11231,N_10857,N_10865);
nor U11232 (N_11232,N_10581,N_10794);
xnor U11233 (N_11233,N_10848,N_10763);
and U11234 (N_11234,N_10958,N_10700);
and U11235 (N_11235,N_10508,N_10666);
and U11236 (N_11236,N_10748,N_10889);
nand U11237 (N_11237,N_10897,N_10711);
nand U11238 (N_11238,N_10899,N_10955);
xnor U11239 (N_11239,N_10896,N_10545);
and U11240 (N_11240,N_10874,N_10670);
nor U11241 (N_11241,N_10901,N_10814);
xor U11242 (N_11242,N_10685,N_10861);
xnor U11243 (N_11243,N_10772,N_10507);
or U11244 (N_11244,N_10815,N_10708);
nand U11245 (N_11245,N_10784,N_10808);
nand U11246 (N_11246,N_10745,N_10994);
and U11247 (N_11247,N_10764,N_10869);
and U11248 (N_11248,N_10726,N_10641);
or U11249 (N_11249,N_10788,N_10836);
and U11250 (N_11250,N_10956,N_10758);
nand U11251 (N_11251,N_10968,N_10784);
and U11252 (N_11252,N_10898,N_10616);
nand U11253 (N_11253,N_10895,N_10649);
nor U11254 (N_11254,N_10877,N_10770);
or U11255 (N_11255,N_10653,N_10638);
or U11256 (N_11256,N_10760,N_10964);
or U11257 (N_11257,N_10536,N_10850);
and U11258 (N_11258,N_10841,N_10700);
nor U11259 (N_11259,N_10503,N_10926);
or U11260 (N_11260,N_10625,N_10908);
nand U11261 (N_11261,N_10691,N_10606);
nand U11262 (N_11262,N_10773,N_10874);
nand U11263 (N_11263,N_10963,N_10782);
nand U11264 (N_11264,N_10944,N_10997);
nor U11265 (N_11265,N_10606,N_10936);
nand U11266 (N_11266,N_10945,N_10851);
xnor U11267 (N_11267,N_10915,N_10916);
nand U11268 (N_11268,N_10599,N_10870);
nand U11269 (N_11269,N_10972,N_10574);
or U11270 (N_11270,N_10909,N_10585);
nor U11271 (N_11271,N_10534,N_10515);
nor U11272 (N_11272,N_10838,N_10918);
and U11273 (N_11273,N_10998,N_10752);
nand U11274 (N_11274,N_10919,N_10670);
or U11275 (N_11275,N_10675,N_10964);
nor U11276 (N_11276,N_10607,N_10763);
nor U11277 (N_11277,N_10889,N_10724);
nor U11278 (N_11278,N_10709,N_10543);
or U11279 (N_11279,N_10818,N_10934);
or U11280 (N_11280,N_10853,N_10691);
or U11281 (N_11281,N_10906,N_10721);
or U11282 (N_11282,N_10702,N_10526);
nand U11283 (N_11283,N_10766,N_10790);
or U11284 (N_11284,N_10838,N_10801);
xor U11285 (N_11285,N_10921,N_10693);
nor U11286 (N_11286,N_10824,N_10982);
xnor U11287 (N_11287,N_10662,N_10533);
or U11288 (N_11288,N_10886,N_10860);
or U11289 (N_11289,N_10744,N_10784);
and U11290 (N_11290,N_10793,N_10591);
and U11291 (N_11291,N_10732,N_10859);
and U11292 (N_11292,N_10964,N_10954);
nor U11293 (N_11293,N_10645,N_10897);
or U11294 (N_11294,N_10561,N_10816);
nor U11295 (N_11295,N_10627,N_10972);
nor U11296 (N_11296,N_10696,N_10976);
nand U11297 (N_11297,N_10873,N_10916);
xnor U11298 (N_11298,N_10902,N_10593);
nor U11299 (N_11299,N_10539,N_10594);
or U11300 (N_11300,N_10648,N_10516);
nand U11301 (N_11301,N_10974,N_10783);
nor U11302 (N_11302,N_10735,N_10785);
xnor U11303 (N_11303,N_10567,N_10823);
xor U11304 (N_11304,N_10714,N_10581);
or U11305 (N_11305,N_10800,N_10506);
xor U11306 (N_11306,N_10774,N_10644);
or U11307 (N_11307,N_10802,N_10754);
nand U11308 (N_11308,N_10837,N_10685);
and U11309 (N_11309,N_10601,N_10906);
nand U11310 (N_11310,N_10862,N_10851);
and U11311 (N_11311,N_10716,N_10640);
nor U11312 (N_11312,N_10504,N_10503);
nor U11313 (N_11313,N_10734,N_10704);
xor U11314 (N_11314,N_10869,N_10967);
nand U11315 (N_11315,N_10599,N_10635);
xor U11316 (N_11316,N_10999,N_10566);
or U11317 (N_11317,N_10718,N_10822);
or U11318 (N_11318,N_10918,N_10900);
and U11319 (N_11319,N_10983,N_10869);
and U11320 (N_11320,N_10804,N_10707);
or U11321 (N_11321,N_10780,N_10635);
or U11322 (N_11322,N_10600,N_10865);
nand U11323 (N_11323,N_10874,N_10727);
xor U11324 (N_11324,N_10999,N_10585);
and U11325 (N_11325,N_10712,N_10536);
nand U11326 (N_11326,N_10629,N_10908);
or U11327 (N_11327,N_10793,N_10849);
and U11328 (N_11328,N_10852,N_10544);
and U11329 (N_11329,N_10737,N_10981);
xor U11330 (N_11330,N_10544,N_10755);
nand U11331 (N_11331,N_10688,N_10936);
xnor U11332 (N_11332,N_10605,N_10948);
or U11333 (N_11333,N_10651,N_10586);
or U11334 (N_11334,N_10811,N_10525);
xor U11335 (N_11335,N_10667,N_10928);
xnor U11336 (N_11336,N_10555,N_10988);
and U11337 (N_11337,N_10506,N_10905);
nand U11338 (N_11338,N_10546,N_10630);
xnor U11339 (N_11339,N_10718,N_10920);
xor U11340 (N_11340,N_10777,N_10893);
xnor U11341 (N_11341,N_10796,N_10659);
and U11342 (N_11342,N_10541,N_10565);
nand U11343 (N_11343,N_10923,N_10760);
or U11344 (N_11344,N_10533,N_10778);
and U11345 (N_11345,N_10850,N_10751);
or U11346 (N_11346,N_10868,N_10683);
xor U11347 (N_11347,N_10561,N_10792);
nand U11348 (N_11348,N_10844,N_10987);
or U11349 (N_11349,N_10500,N_10836);
and U11350 (N_11350,N_10661,N_10795);
nand U11351 (N_11351,N_10697,N_10716);
and U11352 (N_11352,N_10927,N_10619);
or U11353 (N_11353,N_10719,N_10887);
and U11354 (N_11354,N_10764,N_10987);
and U11355 (N_11355,N_10638,N_10924);
nand U11356 (N_11356,N_10757,N_10741);
or U11357 (N_11357,N_10911,N_10556);
nor U11358 (N_11358,N_10518,N_10663);
xor U11359 (N_11359,N_10798,N_10739);
nand U11360 (N_11360,N_10841,N_10965);
or U11361 (N_11361,N_10955,N_10581);
nor U11362 (N_11362,N_10882,N_10531);
nor U11363 (N_11363,N_10846,N_10997);
xnor U11364 (N_11364,N_10560,N_10929);
and U11365 (N_11365,N_10915,N_10510);
nor U11366 (N_11366,N_10808,N_10526);
and U11367 (N_11367,N_10879,N_10680);
nand U11368 (N_11368,N_10845,N_10841);
nor U11369 (N_11369,N_10822,N_10580);
nand U11370 (N_11370,N_10599,N_10540);
nor U11371 (N_11371,N_10626,N_10979);
or U11372 (N_11372,N_10811,N_10519);
nand U11373 (N_11373,N_10614,N_10666);
xnor U11374 (N_11374,N_10937,N_10508);
or U11375 (N_11375,N_10868,N_10511);
or U11376 (N_11376,N_10916,N_10697);
nand U11377 (N_11377,N_10839,N_10569);
nand U11378 (N_11378,N_10799,N_10622);
nand U11379 (N_11379,N_10932,N_10644);
nor U11380 (N_11380,N_10517,N_10641);
or U11381 (N_11381,N_10517,N_10528);
and U11382 (N_11382,N_10967,N_10722);
nor U11383 (N_11383,N_10667,N_10784);
and U11384 (N_11384,N_10892,N_10942);
xnor U11385 (N_11385,N_10823,N_10817);
nand U11386 (N_11386,N_10734,N_10702);
nand U11387 (N_11387,N_10896,N_10656);
xnor U11388 (N_11388,N_10611,N_10612);
and U11389 (N_11389,N_10663,N_10653);
or U11390 (N_11390,N_10990,N_10899);
xnor U11391 (N_11391,N_10710,N_10764);
and U11392 (N_11392,N_10571,N_10807);
nand U11393 (N_11393,N_10961,N_10878);
or U11394 (N_11394,N_10737,N_10618);
nand U11395 (N_11395,N_10505,N_10737);
or U11396 (N_11396,N_10989,N_10863);
nand U11397 (N_11397,N_10977,N_10533);
and U11398 (N_11398,N_10572,N_10899);
xor U11399 (N_11399,N_10534,N_10850);
xnor U11400 (N_11400,N_10857,N_10875);
xnor U11401 (N_11401,N_10858,N_10807);
and U11402 (N_11402,N_10937,N_10933);
xnor U11403 (N_11403,N_10569,N_10977);
xnor U11404 (N_11404,N_10768,N_10614);
nor U11405 (N_11405,N_10623,N_10711);
nor U11406 (N_11406,N_10984,N_10946);
xnor U11407 (N_11407,N_10539,N_10984);
and U11408 (N_11408,N_10703,N_10904);
xnor U11409 (N_11409,N_10529,N_10789);
and U11410 (N_11410,N_10959,N_10912);
and U11411 (N_11411,N_10703,N_10934);
or U11412 (N_11412,N_10607,N_10936);
xnor U11413 (N_11413,N_10706,N_10654);
or U11414 (N_11414,N_10969,N_10959);
and U11415 (N_11415,N_10683,N_10858);
xnor U11416 (N_11416,N_10788,N_10799);
or U11417 (N_11417,N_10854,N_10673);
or U11418 (N_11418,N_10708,N_10791);
xor U11419 (N_11419,N_10737,N_10597);
and U11420 (N_11420,N_10742,N_10856);
nor U11421 (N_11421,N_10818,N_10594);
nor U11422 (N_11422,N_10633,N_10814);
nor U11423 (N_11423,N_10986,N_10928);
xor U11424 (N_11424,N_10756,N_10810);
nor U11425 (N_11425,N_10662,N_10650);
nand U11426 (N_11426,N_10924,N_10857);
or U11427 (N_11427,N_10910,N_10840);
xnor U11428 (N_11428,N_10869,N_10683);
nand U11429 (N_11429,N_10726,N_10649);
or U11430 (N_11430,N_10884,N_10898);
xor U11431 (N_11431,N_10871,N_10827);
nor U11432 (N_11432,N_10943,N_10721);
nand U11433 (N_11433,N_10986,N_10932);
nand U11434 (N_11434,N_10979,N_10757);
nand U11435 (N_11435,N_10967,N_10979);
xnor U11436 (N_11436,N_10554,N_10815);
xnor U11437 (N_11437,N_10931,N_10511);
xnor U11438 (N_11438,N_10831,N_10714);
and U11439 (N_11439,N_10618,N_10710);
nor U11440 (N_11440,N_10754,N_10957);
nand U11441 (N_11441,N_10901,N_10529);
and U11442 (N_11442,N_10770,N_10605);
or U11443 (N_11443,N_10737,N_10701);
xnor U11444 (N_11444,N_10646,N_10955);
nand U11445 (N_11445,N_10609,N_10928);
nor U11446 (N_11446,N_10558,N_10730);
and U11447 (N_11447,N_10830,N_10915);
xor U11448 (N_11448,N_10923,N_10604);
xnor U11449 (N_11449,N_10648,N_10782);
nand U11450 (N_11450,N_10777,N_10588);
nand U11451 (N_11451,N_10751,N_10797);
or U11452 (N_11452,N_10598,N_10597);
or U11453 (N_11453,N_10679,N_10670);
xnor U11454 (N_11454,N_10663,N_10906);
nor U11455 (N_11455,N_10592,N_10666);
nor U11456 (N_11456,N_10525,N_10913);
xor U11457 (N_11457,N_10662,N_10661);
xor U11458 (N_11458,N_10639,N_10819);
nor U11459 (N_11459,N_10561,N_10744);
or U11460 (N_11460,N_10553,N_10600);
nor U11461 (N_11461,N_10989,N_10591);
nand U11462 (N_11462,N_10914,N_10732);
nor U11463 (N_11463,N_10869,N_10560);
nor U11464 (N_11464,N_10705,N_10661);
or U11465 (N_11465,N_10583,N_10555);
and U11466 (N_11466,N_10819,N_10781);
nor U11467 (N_11467,N_10996,N_10928);
or U11468 (N_11468,N_10889,N_10910);
xnor U11469 (N_11469,N_10912,N_10524);
and U11470 (N_11470,N_10751,N_10800);
and U11471 (N_11471,N_10929,N_10703);
xor U11472 (N_11472,N_10506,N_10995);
nor U11473 (N_11473,N_10619,N_10593);
or U11474 (N_11474,N_10539,N_10886);
xnor U11475 (N_11475,N_10569,N_10778);
and U11476 (N_11476,N_10701,N_10576);
and U11477 (N_11477,N_10822,N_10823);
nand U11478 (N_11478,N_10547,N_10846);
nor U11479 (N_11479,N_10944,N_10903);
nor U11480 (N_11480,N_10684,N_10773);
and U11481 (N_11481,N_10807,N_10640);
nor U11482 (N_11482,N_10768,N_10564);
xnor U11483 (N_11483,N_10668,N_10929);
or U11484 (N_11484,N_10689,N_10945);
or U11485 (N_11485,N_10596,N_10780);
or U11486 (N_11486,N_10556,N_10851);
or U11487 (N_11487,N_10727,N_10732);
nand U11488 (N_11488,N_10523,N_10724);
nand U11489 (N_11489,N_10588,N_10942);
nor U11490 (N_11490,N_10570,N_10990);
nor U11491 (N_11491,N_10781,N_10870);
nand U11492 (N_11492,N_10999,N_10920);
and U11493 (N_11493,N_10997,N_10914);
xor U11494 (N_11494,N_10986,N_10813);
xor U11495 (N_11495,N_10812,N_10867);
xnor U11496 (N_11496,N_10810,N_10559);
and U11497 (N_11497,N_10966,N_10993);
nand U11498 (N_11498,N_10631,N_10720);
xnor U11499 (N_11499,N_10934,N_10784);
nor U11500 (N_11500,N_11317,N_11487);
nor U11501 (N_11501,N_11026,N_11373);
nand U11502 (N_11502,N_11061,N_11389);
nand U11503 (N_11503,N_11367,N_11442);
nand U11504 (N_11504,N_11104,N_11233);
nand U11505 (N_11505,N_11129,N_11368);
nand U11506 (N_11506,N_11440,N_11215);
nor U11507 (N_11507,N_11036,N_11451);
nor U11508 (N_11508,N_11286,N_11460);
xor U11509 (N_11509,N_11006,N_11485);
xnor U11510 (N_11510,N_11292,N_11459);
nand U11511 (N_11511,N_11092,N_11477);
nor U11512 (N_11512,N_11366,N_11113);
or U11513 (N_11513,N_11302,N_11280);
or U11514 (N_11514,N_11322,N_11353);
nor U11515 (N_11515,N_11467,N_11076);
nor U11516 (N_11516,N_11393,N_11143);
nor U11517 (N_11517,N_11196,N_11169);
nand U11518 (N_11518,N_11141,N_11381);
nor U11519 (N_11519,N_11334,N_11193);
nor U11520 (N_11520,N_11152,N_11380);
nor U11521 (N_11521,N_11136,N_11240);
and U11522 (N_11522,N_11374,N_11333);
xor U11523 (N_11523,N_11320,N_11438);
or U11524 (N_11524,N_11218,N_11157);
xnor U11525 (N_11525,N_11032,N_11007);
nor U11526 (N_11526,N_11035,N_11391);
nand U11527 (N_11527,N_11078,N_11452);
nand U11528 (N_11528,N_11100,N_11384);
nand U11529 (N_11529,N_11254,N_11172);
xnor U11530 (N_11530,N_11179,N_11156);
xor U11531 (N_11531,N_11465,N_11262);
xnor U11532 (N_11532,N_11133,N_11432);
nor U11533 (N_11533,N_11038,N_11103);
and U11534 (N_11534,N_11147,N_11028);
or U11535 (N_11535,N_11120,N_11344);
nor U11536 (N_11536,N_11230,N_11247);
nor U11537 (N_11537,N_11361,N_11093);
xnor U11538 (N_11538,N_11029,N_11017);
xnor U11539 (N_11539,N_11064,N_11225);
or U11540 (N_11540,N_11050,N_11114);
xnor U11541 (N_11541,N_11189,N_11355);
or U11542 (N_11542,N_11276,N_11447);
nand U11543 (N_11543,N_11101,N_11070);
nand U11544 (N_11544,N_11345,N_11063);
or U11545 (N_11545,N_11168,N_11425);
nor U11546 (N_11546,N_11370,N_11107);
or U11547 (N_11547,N_11111,N_11060);
and U11548 (N_11548,N_11144,N_11273);
and U11549 (N_11549,N_11171,N_11117);
nor U11550 (N_11550,N_11229,N_11135);
or U11551 (N_11551,N_11080,N_11476);
xnor U11552 (N_11552,N_11263,N_11140);
or U11553 (N_11553,N_11019,N_11269);
nor U11554 (N_11554,N_11191,N_11095);
or U11555 (N_11555,N_11245,N_11318);
or U11556 (N_11556,N_11200,N_11174);
or U11557 (N_11557,N_11204,N_11031);
nor U11558 (N_11558,N_11148,N_11348);
and U11559 (N_11559,N_11255,N_11416);
and U11560 (N_11560,N_11206,N_11347);
nor U11561 (N_11561,N_11058,N_11216);
or U11562 (N_11562,N_11219,N_11307);
or U11563 (N_11563,N_11358,N_11072);
and U11564 (N_11564,N_11237,N_11242);
nor U11565 (N_11565,N_11332,N_11201);
nor U11566 (N_11566,N_11155,N_11371);
xor U11567 (N_11567,N_11372,N_11112);
nand U11568 (N_11568,N_11359,N_11375);
and U11569 (N_11569,N_11162,N_11088);
or U11570 (N_11570,N_11034,N_11354);
xnor U11571 (N_11571,N_11000,N_11085);
nor U11572 (N_11572,N_11160,N_11102);
nor U11573 (N_11573,N_11024,N_11183);
and U11574 (N_11574,N_11453,N_11119);
nand U11575 (N_11575,N_11441,N_11411);
and U11576 (N_11576,N_11491,N_11398);
and U11577 (N_11577,N_11079,N_11470);
and U11578 (N_11578,N_11426,N_11249);
and U11579 (N_11579,N_11409,N_11258);
or U11580 (N_11580,N_11335,N_11291);
xnor U11581 (N_11581,N_11468,N_11296);
nand U11582 (N_11582,N_11131,N_11122);
or U11583 (N_11583,N_11264,N_11443);
or U11584 (N_11584,N_11082,N_11110);
xnor U11585 (N_11585,N_11421,N_11455);
or U11586 (N_11586,N_11331,N_11486);
nand U11587 (N_11587,N_11068,N_11257);
and U11588 (N_11588,N_11436,N_11349);
and U11589 (N_11589,N_11473,N_11134);
nand U11590 (N_11590,N_11021,N_11271);
xnor U11591 (N_11591,N_11256,N_11422);
nor U11592 (N_11592,N_11239,N_11163);
and U11593 (N_11593,N_11170,N_11313);
or U11594 (N_11594,N_11378,N_11016);
or U11595 (N_11595,N_11327,N_11096);
nor U11596 (N_11596,N_11410,N_11434);
nand U11597 (N_11597,N_11338,N_11464);
or U11598 (N_11598,N_11165,N_11294);
and U11599 (N_11599,N_11175,N_11265);
xnor U11600 (N_11600,N_11091,N_11118);
xnor U11601 (N_11601,N_11176,N_11243);
nand U11602 (N_11602,N_11192,N_11362);
or U11603 (N_11603,N_11472,N_11494);
nor U11604 (N_11604,N_11462,N_11329);
nand U11605 (N_11605,N_11083,N_11306);
or U11606 (N_11606,N_11207,N_11126);
nand U11607 (N_11607,N_11044,N_11252);
and U11608 (N_11608,N_11417,N_11402);
nand U11609 (N_11609,N_11444,N_11020);
xor U11610 (N_11610,N_11047,N_11385);
nand U11611 (N_11611,N_11221,N_11304);
xor U11612 (N_11612,N_11356,N_11309);
and U11613 (N_11613,N_11084,N_11180);
nand U11614 (N_11614,N_11167,N_11469);
nand U11615 (N_11615,N_11316,N_11337);
nor U11616 (N_11616,N_11159,N_11446);
or U11617 (N_11617,N_11458,N_11151);
nor U11618 (N_11618,N_11153,N_11051);
nor U11619 (N_11619,N_11301,N_11098);
xnor U11620 (N_11620,N_11281,N_11161);
nor U11621 (N_11621,N_11379,N_11405);
and U11622 (N_11622,N_11399,N_11097);
xnor U11623 (N_11623,N_11445,N_11369);
or U11624 (N_11624,N_11099,N_11094);
nor U11625 (N_11625,N_11392,N_11423);
or U11626 (N_11626,N_11115,N_11275);
nand U11627 (N_11627,N_11124,N_11489);
and U11628 (N_11628,N_11213,N_11203);
and U11629 (N_11629,N_11430,N_11323);
and U11630 (N_11630,N_11346,N_11224);
and U11631 (N_11631,N_11270,N_11057);
and U11632 (N_11632,N_11339,N_11238);
nor U11633 (N_11633,N_11289,N_11182);
nor U11634 (N_11634,N_11043,N_11395);
or U11635 (N_11635,N_11074,N_11138);
and U11636 (N_11636,N_11069,N_11435);
and U11637 (N_11637,N_11001,N_11360);
xor U11638 (N_11638,N_11056,N_11315);
or U11639 (N_11639,N_11277,N_11437);
and U11640 (N_11640,N_11431,N_11283);
and U11641 (N_11641,N_11266,N_11282);
nor U11642 (N_11642,N_11042,N_11420);
and U11643 (N_11643,N_11414,N_11041);
nor U11644 (N_11644,N_11033,N_11412);
nand U11645 (N_11645,N_11212,N_11382);
xor U11646 (N_11646,N_11186,N_11456);
or U11647 (N_11647,N_11295,N_11298);
nand U11648 (N_11648,N_11478,N_11363);
xor U11649 (N_11649,N_11012,N_11383);
xnor U11650 (N_11650,N_11128,N_11211);
and U11651 (N_11651,N_11177,N_11222);
xnor U11652 (N_11652,N_11474,N_11045);
xor U11653 (N_11653,N_11299,N_11279);
and U11654 (N_11654,N_11433,N_11198);
or U11655 (N_11655,N_11387,N_11077);
nor U11656 (N_11656,N_11241,N_11178);
nor U11657 (N_11657,N_11228,N_11261);
nand U11658 (N_11658,N_11108,N_11413);
or U11659 (N_11659,N_11287,N_11268);
xor U11660 (N_11660,N_11272,N_11429);
xnor U11661 (N_11661,N_11246,N_11397);
nand U11662 (N_11662,N_11483,N_11448);
xnor U11663 (N_11663,N_11227,N_11428);
nand U11664 (N_11664,N_11482,N_11340);
nor U11665 (N_11665,N_11008,N_11154);
and U11666 (N_11666,N_11314,N_11439);
nand U11667 (N_11667,N_11054,N_11208);
and U11668 (N_11668,N_11052,N_11259);
xnor U11669 (N_11669,N_11014,N_11025);
and U11670 (N_11670,N_11146,N_11199);
xor U11671 (N_11671,N_11415,N_11197);
nor U11672 (N_11672,N_11493,N_11010);
or U11673 (N_11673,N_11449,N_11496);
or U11674 (N_11674,N_11018,N_11173);
or U11675 (N_11675,N_11300,N_11454);
nor U11676 (N_11676,N_11002,N_11343);
nand U11677 (N_11677,N_11022,N_11365);
and U11678 (N_11678,N_11009,N_11116);
nand U11679 (N_11679,N_11461,N_11466);
xnor U11680 (N_11680,N_11231,N_11303);
xor U11681 (N_11681,N_11086,N_11293);
and U11682 (N_11682,N_11181,N_11226);
nand U11683 (N_11683,N_11424,N_11125);
and U11684 (N_11684,N_11040,N_11284);
and U11685 (N_11685,N_11336,N_11325);
nand U11686 (N_11686,N_11142,N_11404);
and U11687 (N_11687,N_11342,N_11364);
nand U11688 (N_11688,N_11067,N_11390);
nand U11689 (N_11689,N_11351,N_11046);
or U11690 (N_11690,N_11190,N_11495);
xor U11691 (N_11691,N_11039,N_11013);
nor U11692 (N_11692,N_11075,N_11223);
or U11693 (N_11693,N_11400,N_11150);
or U11694 (N_11694,N_11475,N_11187);
nand U11695 (N_11695,N_11248,N_11406);
xnor U11696 (N_11696,N_11130,N_11324);
xnor U11697 (N_11697,N_11048,N_11403);
xnor U11698 (N_11698,N_11419,N_11066);
xor U11699 (N_11699,N_11023,N_11109);
xnor U11700 (N_11700,N_11184,N_11499);
or U11701 (N_11701,N_11260,N_11278);
and U11702 (N_11702,N_11087,N_11401);
xor U11703 (N_11703,N_11326,N_11005);
or U11704 (N_11704,N_11071,N_11090);
nand U11705 (N_11705,N_11049,N_11484);
nor U11706 (N_11706,N_11105,N_11127);
xnor U11707 (N_11707,N_11352,N_11463);
and U11708 (N_11708,N_11202,N_11376);
xnor U11709 (N_11709,N_11328,N_11418);
or U11710 (N_11710,N_11386,N_11194);
xor U11711 (N_11711,N_11062,N_11205);
and U11712 (N_11712,N_11235,N_11220);
or U11713 (N_11713,N_11471,N_11004);
and U11714 (N_11714,N_11188,N_11003);
and U11715 (N_11715,N_11288,N_11274);
xnor U11716 (N_11716,N_11308,N_11166);
nor U11717 (N_11717,N_11479,N_11350);
and U11718 (N_11718,N_11065,N_11195);
and U11719 (N_11719,N_11234,N_11037);
or U11720 (N_11720,N_11121,N_11015);
and U11721 (N_11721,N_11158,N_11055);
or U11722 (N_11722,N_11053,N_11232);
nor U11723 (N_11723,N_11388,N_11145);
and U11724 (N_11724,N_11209,N_11490);
or U11725 (N_11725,N_11137,N_11377);
and U11726 (N_11726,N_11267,N_11396);
nor U11727 (N_11727,N_11149,N_11321);
xor U11728 (N_11728,N_11311,N_11488);
or U11729 (N_11729,N_11059,N_11210);
or U11730 (N_11730,N_11185,N_11250);
and U11731 (N_11731,N_11139,N_11244);
nand U11732 (N_11732,N_11312,N_11285);
xor U11733 (N_11733,N_11305,N_11027);
or U11734 (N_11734,N_11253,N_11427);
and U11735 (N_11735,N_11217,N_11123);
nor U11736 (N_11736,N_11073,N_11106);
and U11737 (N_11737,N_11290,N_11492);
nor U11738 (N_11738,N_11357,N_11251);
nand U11739 (N_11739,N_11497,N_11341);
nand U11740 (N_11740,N_11089,N_11214);
nor U11741 (N_11741,N_11394,N_11310);
nand U11742 (N_11742,N_11319,N_11498);
nor U11743 (N_11743,N_11450,N_11480);
or U11744 (N_11744,N_11164,N_11481);
nand U11745 (N_11745,N_11457,N_11297);
nand U11746 (N_11746,N_11081,N_11407);
nand U11747 (N_11747,N_11132,N_11030);
or U11748 (N_11748,N_11236,N_11330);
nand U11749 (N_11749,N_11011,N_11408);
nand U11750 (N_11750,N_11007,N_11075);
nand U11751 (N_11751,N_11303,N_11240);
nor U11752 (N_11752,N_11397,N_11451);
nor U11753 (N_11753,N_11212,N_11120);
nor U11754 (N_11754,N_11152,N_11206);
xnor U11755 (N_11755,N_11416,N_11294);
nand U11756 (N_11756,N_11432,N_11100);
xnor U11757 (N_11757,N_11120,N_11291);
nand U11758 (N_11758,N_11008,N_11371);
nor U11759 (N_11759,N_11048,N_11479);
xnor U11760 (N_11760,N_11055,N_11067);
xnor U11761 (N_11761,N_11477,N_11466);
nor U11762 (N_11762,N_11157,N_11305);
and U11763 (N_11763,N_11288,N_11011);
nor U11764 (N_11764,N_11428,N_11221);
or U11765 (N_11765,N_11179,N_11192);
and U11766 (N_11766,N_11368,N_11080);
xnor U11767 (N_11767,N_11217,N_11486);
xor U11768 (N_11768,N_11404,N_11382);
nand U11769 (N_11769,N_11353,N_11260);
and U11770 (N_11770,N_11494,N_11421);
nand U11771 (N_11771,N_11299,N_11239);
or U11772 (N_11772,N_11248,N_11417);
xnor U11773 (N_11773,N_11317,N_11281);
xnor U11774 (N_11774,N_11122,N_11473);
xor U11775 (N_11775,N_11087,N_11408);
nand U11776 (N_11776,N_11221,N_11043);
or U11777 (N_11777,N_11388,N_11009);
xor U11778 (N_11778,N_11191,N_11348);
nor U11779 (N_11779,N_11360,N_11013);
nand U11780 (N_11780,N_11000,N_11240);
nand U11781 (N_11781,N_11117,N_11266);
and U11782 (N_11782,N_11186,N_11311);
xnor U11783 (N_11783,N_11420,N_11214);
xor U11784 (N_11784,N_11394,N_11081);
or U11785 (N_11785,N_11468,N_11279);
xor U11786 (N_11786,N_11404,N_11310);
or U11787 (N_11787,N_11036,N_11377);
xor U11788 (N_11788,N_11000,N_11374);
or U11789 (N_11789,N_11392,N_11311);
nor U11790 (N_11790,N_11491,N_11248);
and U11791 (N_11791,N_11197,N_11055);
or U11792 (N_11792,N_11387,N_11091);
nand U11793 (N_11793,N_11027,N_11124);
nand U11794 (N_11794,N_11491,N_11143);
and U11795 (N_11795,N_11142,N_11266);
xnor U11796 (N_11796,N_11235,N_11270);
nor U11797 (N_11797,N_11121,N_11198);
xnor U11798 (N_11798,N_11152,N_11365);
or U11799 (N_11799,N_11077,N_11403);
or U11800 (N_11800,N_11397,N_11308);
or U11801 (N_11801,N_11260,N_11183);
or U11802 (N_11802,N_11359,N_11332);
nand U11803 (N_11803,N_11093,N_11314);
nand U11804 (N_11804,N_11410,N_11183);
or U11805 (N_11805,N_11141,N_11430);
nor U11806 (N_11806,N_11391,N_11102);
nand U11807 (N_11807,N_11009,N_11485);
or U11808 (N_11808,N_11084,N_11178);
nand U11809 (N_11809,N_11317,N_11097);
nand U11810 (N_11810,N_11054,N_11400);
xor U11811 (N_11811,N_11461,N_11152);
nand U11812 (N_11812,N_11466,N_11036);
and U11813 (N_11813,N_11093,N_11373);
xor U11814 (N_11814,N_11479,N_11195);
nor U11815 (N_11815,N_11124,N_11011);
nand U11816 (N_11816,N_11131,N_11329);
and U11817 (N_11817,N_11159,N_11332);
or U11818 (N_11818,N_11300,N_11460);
xor U11819 (N_11819,N_11491,N_11150);
nand U11820 (N_11820,N_11301,N_11220);
xnor U11821 (N_11821,N_11044,N_11397);
nand U11822 (N_11822,N_11493,N_11337);
nand U11823 (N_11823,N_11320,N_11220);
xnor U11824 (N_11824,N_11471,N_11289);
or U11825 (N_11825,N_11066,N_11091);
nor U11826 (N_11826,N_11400,N_11314);
and U11827 (N_11827,N_11029,N_11412);
nor U11828 (N_11828,N_11148,N_11175);
and U11829 (N_11829,N_11170,N_11015);
xnor U11830 (N_11830,N_11495,N_11464);
nand U11831 (N_11831,N_11139,N_11229);
nor U11832 (N_11832,N_11016,N_11358);
nand U11833 (N_11833,N_11297,N_11473);
nand U11834 (N_11834,N_11132,N_11305);
xor U11835 (N_11835,N_11354,N_11183);
and U11836 (N_11836,N_11194,N_11261);
nand U11837 (N_11837,N_11147,N_11063);
nand U11838 (N_11838,N_11246,N_11006);
xor U11839 (N_11839,N_11200,N_11196);
or U11840 (N_11840,N_11437,N_11077);
xnor U11841 (N_11841,N_11065,N_11414);
nand U11842 (N_11842,N_11336,N_11461);
nand U11843 (N_11843,N_11115,N_11064);
or U11844 (N_11844,N_11099,N_11163);
or U11845 (N_11845,N_11011,N_11317);
nor U11846 (N_11846,N_11412,N_11351);
nand U11847 (N_11847,N_11261,N_11112);
nor U11848 (N_11848,N_11286,N_11454);
and U11849 (N_11849,N_11239,N_11465);
and U11850 (N_11850,N_11072,N_11287);
nand U11851 (N_11851,N_11218,N_11476);
nor U11852 (N_11852,N_11142,N_11466);
xor U11853 (N_11853,N_11418,N_11392);
or U11854 (N_11854,N_11312,N_11353);
or U11855 (N_11855,N_11319,N_11035);
nor U11856 (N_11856,N_11169,N_11162);
nand U11857 (N_11857,N_11054,N_11489);
nor U11858 (N_11858,N_11205,N_11220);
nand U11859 (N_11859,N_11369,N_11089);
xor U11860 (N_11860,N_11150,N_11232);
nor U11861 (N_11861,N_11030,N_11091);
or U11862 (N_11862,N_11156,N_11313);
nand U11863 (N_11863,N_11095,N_11099);
or U11864 (N_11864,N_11257,N_11247);
and U11865 (N_11865,N_11353,N_11066);
xnor U11866 (N_11866,N_11080,N_11389);
nand U11867 (N_11867,N_11011,N_11256);
and U11868 (N_11868,N_11263,N_11335);
nand U11869 (N_11869,N_11077,N_11384);
nor U11870 (N_11870,N_11497,N_11176);
nor U11871 (N_11871,N_11385,N_11202);
nand U11872 (N_11872,N_11418,N_11431);
xor U11873 (N_11873,N_11078,N_11339);
or U11874 (N_11874,N_11187,N_11140);
nor U11875 (N_11875,N_11180,N_11284);
or U11876 (N_11876,N_11336,N_11048);
nor U11877 (N_11877,N_11170,N_11065);
nand U11878 (N_11878,N_11345,N_11350);
or U11879 (N_11879,N_11176,N_11238);
nand U11880 (N_11880,N_11022,N_11107);
or U11881 (N_11881,N_11470,N_11221);
nor U11882 (N_11882,N_11395,N_11072);
nor U11883 (N_11883,N_11395,N_11402);
nand U11884 (N_11884,N_11452,N_11451);
nor U11885 (N_11885,N_11436,N_11196);
or U11886 (N_11886,N_11064,N_11162);
nor U11887 (N_11887,N_11161,N_11492);
and U11888 (N_11888,N_11294,N_11305);
nor U11889 (N_11889,N_11050,N_11275);
or U11890 (N_11890,N_11147,N_11318);
nor U11891 (N_11891,N_11437,N_11220);
xnor U11892 (N_11892,N_11160,N_11022);
nor U11893 (N_11893,N_11414,N_11112);
or U11894 (N_11894,N_11460,N_11384);
and U11895 (N_11895,N_11480,N_11240);
and U11896 (N_11896,N_11284,N_11292);
and U11897 (N_11897,N_11325,N_11312);
nand U11898 (N_11898,N_11214,N_11052);
xor U11899 (N_11899,N_11448,N_11062);
xor U11900 (N_11900,N_11032,N_11150);
or U11901 (N_11901,N_11093,N_11370);
xnor U11902 (N_11902,N_11360,N_11416);
nand U11903 (N_11903,N_11004,N_11038);
nand U11904 (N_11904,N_11399,N_11157);
xor U11905 (N_11905,N_11455,N_11498);
and U11906 (N_11906,N_11216,N_11245);
nor U11907 (N_11907,N_11366,N_11401);
or U11908 (N_11908,N_11139,N_11472);
nand U11909 (N_11909,N_11098,N_11457);
and U11910 (N_11910,N_11376,N_11287);
nand U11911 (N_11911,N_11467,N_11342);
or U11912 (N_11912,N_11023,N_11359);
and U11913 (N_11913,N_11003,N_11042);
nor U11914 (N_11914,N_11232,N_11070);
xor U11915 (N_11915,N_11091,N_11291);
and U11916 (N_11916,N_11018,N_11116);
nor U11917 (N_11917,N_11215,N_11293);
and U11918 (N_11918,N_11344,N_11225);
or U11919 (N_11919,N_11022,N_11487);
nand U11920 (N_11920,N_11255,N_11309);
nand U11921 (N_11921,N_11442,N_11113);
xor U11922 (N_11922,N_11186,N_11257);
and U11923 (N_11923,N_11387,N_11090);
and U11924 (N_11924,N_11400,N_11397);
or U11925 (N_11925,N_11166,N_11246);
xnor U11926 (N_11926,N_11179,N_11100);
nor U11927 (N_11927,N_11261,N_11428);
nand U11928 (N_11928,N_11276,N_11209);
and U11929 (N_11929,N_11399,N_11232);
or U11930 (N_11930,N_11098,N_11219);
xnor U11931 (N_11931,N_11037,N_11001);
nor U11932 (N_11932,N_11227,N_11194);
or U11933 (N_11933,N_11038,N_11068);
xnor U11934 (N_11934,N_11237,N_11452);
xor U11935 (N_11935,N_11047,N_11418);
nand U11936 (N_11936,N_11101,N_11309);
xor U11937 (N_11937,N_11359,N_11256);
nor U11938 (N_11938,N_11227,N_11186);
xnor U11939 (N_11939,N_11226,N_11051);
and U11940 (N_11940,N_11100,N_11178);
or U11941 (N_11941,N_11260,N_11085);
nand U11942 (N_11942,N_11496,N_11150);
nand U11943 (N_11943,N_11390,N_11296);
nor U11944 (N_11944,N_11120,N_11206);
or U11945 (N_11945,N_11444,N_11052);
or U11946 (N_11946,N_11359,N_11051);
xor U11947 (N_11947,N_11137,N_11246);
nor U11948 (N_11948,N_11393,N_11075);
nand U11949 (N_11949,N_11447,N_11110);
and U11950 (N_11950,N_11474,N_11108);
or U11951 (N_11951,N_11136,N_11426);
or U11952 (N_11952,N_11177,N_11329);
and U11953 (N_11953,N_11036,N_11457);
xnor U11954 (N_11954,N_11037,N_11317);
and U11955 (N_11955,N_11311,N_11023);
nor U11956 (N_11956,N_11458,N_11463);
and U11957 (N_11957,N_11378,N_11407);
and U11958 (N_11958,N_11057,N_11200);
or U11959 (N_11959,N_11456,N_11276);
or U11960 (N_11960,N_11366,N_11375);
nand U11961 (N_11961,N_11005,N_11453);
nand U11962 (N_11962,N_11444,N_11352);
nor U11963 (N_11963,N_11384,N_11450);
nor U11964 (N_11964,N_11087,N_11441);
xnor U11965 (N_11965,N_11156,N_11285);
and U11966 (N_11966,N_11328,N_11033);
nor U11967 (N_11967,N_11108,N_11318);
and U11968 (N_11968,N_11119,N_11444);
nand U11969 (N_11969,N_11348,N_11462);
or U11970 (N_11970,N_11178,N_11302);
nor U11971 (N_11971,N_11120,N_11319);
and U11972 (N_11972,N_11136,N_11253);
nor U11973 (N_11973,N_11448,N_11343);
nand U11974 (N_11974,N_11245,N_11008);
xnor U11975 (N_11975,N_11265,N_11290);
and U11976 (N_11976,N_11349,N_11407);
or U11977 (N_11977,N_11251,N_11267);
xnor U11978 (N_11978,N_11282,N_11360);
nor U11979 (N_11979,N_11132,N_11057);
or U11980 (N_11980,N_11314,N_11021);
nand U11981 (N_11981,N_11444,N_11181);
xnor U11982 (N_11982,N_11311,N_11250);
or U11983 (N_11983,N_11399,N_11142);
and U11984 (N_11984,N_11282,N_11263);
xnor U11985 (N_11985,N_11497,N_11410);
or U11986 (N_11986,N_11421,N_11309);
or U11987 (N_11987,N_11435,N_11380);
nor U11988 (N_11988,N_11073,N_11403);
nor U11989 (N_11989,N_11465,N_11331);
nand U11990 (N_11990,N_11305,N_11064);
nor U11991 (N_11991,N_11380,N_11306);
nor U11992 (N_11992,N_11001,N_11096);
and U11993 (N_11993,N_11450,N_11148);
nor U11994 (N_11994,N_11319,N_11436);
and U11995 (N_11995,N_11280,N_11155);
xor U11996 (N_11996,N_11269,N_11053);
or U11997 (N_11997,N_11342,N_11354);
xor U11998 (N_11998,N_11062,N_11262);
nand U11999 (N_11999,N_11219,N_11226);
nor U12000 (N_12000,N_11839,N_11986);
nand U12001 (N_12001,N_11500,N_11727);
or U12002 (N_12002,N_11878,N_11693);
nor U12003 (N_12003,N_11554,N_11646);
xnor U12004 (N_12004,N_11725,N_11502);
xnor U12005 (N_12005,N_11989,N_11962);
and U12006 (N_12006,N_11755,N_11843);
and U12007 (N_12007,N_11606,N_11864);
nand U12008 (N_12008,N_11783,N_11598);
and U12009 (N_12009,N_11972,N_11967);
nor U12010 (N_12010,N_11726,N_11649);
xor U12011 (N_12011,N_11935,N_11737);
nand U12012 (N_12012,N_11776,N_11604);
or U12013 (N_12013,N_11719,N_11671);
or U12014 (N_12014,N_11885,N_11564);
nor U12015 (N_12015,N_11634,N_11603);
nor U12016 (N_12016,N_11516,N_11684);
nand U12017 (N_12017,N_11888,N_11668);
or U12018 (N_12018,N_11542,N_11552);
or U12019 (N_12019,N_11589,N_11653);
nor U12020 (N_12020,N_11907,N_11617);
xor U12021 (N_12021,N_11581,N_11541);
nand U12022 (N_12022,N_11505,N_11764);
nor U12023 (N_12023,N_11922,N_11501);
and U12024 (N_12024,N_11995,N_11645);
or U12025 (N_12025,N_11512,N_11510);
and U12026 (N_12026,N_11580,N_11774);
xnor U12027 (N_12027,N_11520,N_11840);
nor U12028 (N_12028,N_11681,N_11909);
and U12029 (N_12029,N_11584,N_11752);
nor U12030 (N_12030,N_11627,N_11696);
nand U12031 (N_12031,N_11615,N_11712);
xnor U12032 (N_12032,N_11970,N_11673);
nand U12033 (N_12033,N_11539,N_11526);
or U12034 (N_12034,N_11728,N_11994);
and U12035 (N_12035,N_11924,N_11999);
nor U12036 (N_12036,N_11622,N_11988);
and U12037 (N_12037,N_11705,N_11574);
nand U12038 (N_12038,N_11829,N_11561);
xor U12039 (N_12039,N_11810,N_11555);
xnor U12040 (N_12040,N_11895,N_11915);
and U12041 (N_12041,N_11631,N_11619);
and U12042 (N_12042,N_11704,N_11889);
and U12043 (N_12043,N_11716,N_11641);
or U12044 (N_12044,N_11896,N_11954);
xnor U12045 (N_12045,N_11969,N_11964);
or U12046 (N_12046,N_11533,N_11934);
nand U12047 (N_12047,N_11770,N_11666);
xnor U12048 (N_12048,N_11971,N_11593);
and U12049 (N_12049,N_11744,N_11953);
nor U12050 (N_12050,N_11578,N_11754);
nand U12051 (N_12051,N_11957,N_11587);
nor U12052 (N_12052,N_11858,N_11626);
or U12053 (N_12053,N_11700,N_11694);
nor U12054 (N_12054,N_11799,N_11675);
nand U12055 (N_12055,N_11659,N_11921);
and U12056 (N_12056,N_11750,N_11530);
and U12057 (N_12057,N_11515,N_11819);
nand U12058 (N_12058,N_11960,N_11644);
or U12059 (N_12059,N_11871,N_11767);
nand U12060 (N_12060,N_11674,N_11656);
nand U12061 (N_12061,N_11630,N_11911);
xnor U12062 (N_12062,N_11718,N_11600);
xnor U12063 (N_12063,N_11883,N_11944);
and U12064 (N_12064,N_11943,N_11794);
and U12065 (N_12065,N_11607,N_11929);
nor U12066 (N_12066,N_11820,N_11812);
nand U12067 (N_12067,N_11525,N_11789);
nor U12068 (N_12068,N_11602,N_11551);
and U12069 (N_12069,N_11667,N_11601);
nor U12070 (N_12070,N_11879,N_11761);
xor U12071 (N_12071,N_11594,N_11628);
nor U12072 (N_12072,N_11798,N_11872);
xor U12073 (N_12073,N_11762,N_11570);
and U12074 (N_12074,N_11816,N_11865);
and U12075 (N_12075,N_11629,N_11746);
and U12076 (N_12076,N_11660,N_11753);
and U12077 (N_12077,N_11766,N_11874);
nor U12078 (N_12078,N_11528,N_11648);
nand U12079 (N_12079,N_11850,N_11679);
nand U12080 (N_12080,N_11984,N_11847);
or U12081 (N_12081,N_11625,N_11811);
nand U12082 (N_12082,N_11723,N_11866);
nand U12083 (N_12083,N_11663,N_11832);
nor U12084 (N_12084,N_11939,N_11608);
or U12085 (N_12085,N_11688,N_11747);
and U12086 (N_12086,N_11886,N_11519);
and U12087 (N_12087,N_11857,N_11848);
nor U12088 (N_12088,N_11524,N_11790);
nand U12089 (N_12089,N_11758,N_11612);
or U12090 (N_12090,N_11855,N_11639);
xor U12091 (N_12091,N_11796,N_11546);
or U12092 (N_12092,N_11662,N_11956);
or U12093 (N_12093,N_11821,N_11860);
or U12094 (N_12094,N_11773,N_11958);
or U12095 (N_12095,N_11562,N_11738);
nor U12096 (N_12096,N_11894,N_11749);
nand U12097 (N_12097,N_11527,N_11565);
and U12098 (N_12098,N_11740,N_11950);
nor U12099 (N_12099,N_11784,N_11788);
xnor U12100 (N_12100,N_11987,N_11532);
or U12101 (N_12101,N_11813,N_11881);
nand U12102 (N_12102,N_11509,N_11707);
nand U12103 (N_12103,N_11805,N_11624);
xor U12104 (N_12104,N_11852,N_11635);
and U12105 (N_12105,N_11677,N_11765);
or U12106 (N_12106,N_11717,N_11916);
and U12107 (N_12107,N_11926,N_11948);
nor U12108 (N_12108,N_11529,N_11701);
nand U12109 (N_12109,N_11946,N_11592);
or U12110 (N_12110,N_11913,N_11538);
nor U12111 (N_12111,N_11993,N_11504);
and U12112 (N_12112,N_11898,N_11891);
nor U12113 (N_12113,N_11535,N_11835);
or U12114 (N_12114,N_11616,N_11801);
nand U12115 (N_12115,N_11951,N_11664);
or U12116 (N_12116,N_11997,N_11611);
or U12117 (N_12117,N_11743,N_11920);
or U12118 (N_12118,N_11632,N_11869);
and U12119 (N_12119,N_11787,N_11678);
and U12120 (N_12120,N_11672,N_11748);
and U12121 (N_12121,N_11806,N_11521);
or U12122 (N_12122,N_11928,N_11556);
nand U12123 (N_12123,N_11685,N_11730);
or U12124 (N_12124,N_11825,N_11779);
nor U12125 (N_12125,N_11724,N_11807);
or U12126 (N_12126,N_11808,N_11523);
xnor U12127 (N_12127,N_11853,N_11563);
xnor U12128 (N_12128,N_11975,N_11669);
nor U12129 (N_12129,N_11837,N_11949);
or U12130 (N_12130,N_11751,N_11623);
nand U12131 (N_12131,N_11834,N_11591);
or U12132 (N_12132,N_11938,N_11817);
or U12133 (N_12133,N_11933,N_11560);
xnor U12134 (N_12134,N_11899,N_11518);
and U12135 (N_12135,N_11536,N_11595);
and U12136 (N_12136,N_11809,N_11877);
and U12137 (N_12137,N_11609,N_11867);
xnor U12138 (N_12138,N_11937,N_11577);
nor U12139 (N_12139,N_11550,N_11522);
or U12140 (N_12140,N_11711,N_11952);
or U12141 (N_12141,N_11976,N_11981);
or U12142 (N_12142,N_11793,N_11769);
or U12143 (N_12143,N_11978,N_11729);
and U12144 (N_12144,N_11849,N_11508);
nor U12145 (N_12145,N_11912,N_11880);
nand U12146 (N_12146,N_11768,N_11559);
nor U12147 (N_12147,N_11540,N_11985);
nor U12148 (N_12148,N_11698,N_11780);
xor U12149 (N_12149,N_11804,N_11585);
nor U12150 (N_12150,N_11586,N_11873);
nand U12151 (N_12151,N_11941,N_11683);
nand U12152 (N_12152,N_11710,N_11859);
nor U12153 (N_12153,N_11545,N_11823);
nor U12154 (N_12154,N_11513,N_11637);
xnor U12155 (N_12155,N_11618,N_11945);
nor U12156 (N_12156,N_11680,N_11590);
nand U12157 (N_12157,N_11745,N_11936);
and U12158 (N_12158,N_11573,N_11983);
and U12159 (N_12159,N_11961,N_11661);
and U12160 (N_12160,N_11919,N_11982);
or U12161 (N_12161,N_11695,N_11980);
xnor U12162 (N_12162,N_11868,N_11965);
or U12163 (N_12163,N_11721,N_11687);
xor U12164 (N_12164,N_11854,N_11905);
or U12165 (N_12165,N_11955,N_11763);
or U12166 (N_12166,N_11741,N_11582);
and U12167 (N_12167,N_11733,N_11537);
and U12168 (N_12168,N_11826,N_11633);
xnor U12169 (N_12169,N_11651,N_11781);
xnor U12170 (N_12170,N_11549,N_11566);
and U12171 (N_12171,N_11670,N_11697);
nand U12172 (N_12172,N_11599,N_11771);
nor U12173 (N_12173,N_11507,N_11918);
or U12174 (N_12174,N_11947,N_11786);
or U12175 (N_12175,N_11568,N_11818);
xor U12176 (N_12176,N_11640,N_11890);
nor U12177 (N_12177,N_11692,N_11931);
and U12178 (N_12178,N_11824,N_11792);
xnor U12179 (N_12179,N_11803,N_11914);
nor U12180 (N_12180,N_11828,N_11567);
nand U12181 (N_12181,N_11511,N_11990);
nand U12182 (N_12182,N_11517,N_11547);
and U12183 (N_12183,N_11605,N_11917);
and U12184 (N_12184,N_11991,N_11543);
or U12185 (N_12185,N_11650,N_11802);
xnor U12186 (N_12186,N_11652,N_11887);
and U12187 (N_12187,N_11884,N_11772);
or U12188 (N_12188,N_11657,N_11734);
nor U12189 (N_12189,N_11557,N_11709);
and U12190 (N_12190,N_11963,N_11940);
or U12191 (N_12191,N_11875,N_11572);
nand U12192 (N_12192,N_11930,N_11966);
nor U12193 (N_12193,N_11757,N_11882);
nand U12194 (N_12194,N_11910,N_11756);
xor U12195 (N_12195,N_11610,N_11862);
or U12196 (N_12196,N_11815,N_11553);
nor U12197 (N_12197,N_11760,N_11703);
nor U12198 (N_12198,N_11548,N_11979);
and U12199 (N_12199,N_11569,N_11827);
or U12200 (N_12200,N_11699,N_11676);
nor U12201 (N_12201,N_11842,N_11583);
or U12202 (N_12202,N_11742,N_11851);
xor U12203 (N_12203,N_11841,N_11782);
and U12204 (N_12204,N_11702,N_11778);
and U12205 (N_12205,N_11706,N_11814);
and U12206 (N_12206,N_11658,N_11998);
nor U12207 (N_12207,N_11731,N_11797);
nand U12208 (N_12208,N_11932,N_11613);
nand U12209 (N_12209,N_11836,N_11708);
or U12210 (N_12210,N_11791,N_11900);
nand U12211 (N_12211,N_11654,N_11643);
xnor U12212 (N_12212,N_11691,N_11777);
nor U12213 (N_12213,N_11892,N_11588);
and U12214 (N_12214,N_11996,N_11714);
or U12215 (N_12215,N_11534,N_11925);
nand U12216 (N_12216,N_11621,N_11785);
nand U12217 (N_12217,N_11893,N_11636);
xor U12218 (N_12218,N_11973,N_11992);
xnor U12219 (N_12219,N_11795,N_11923);
nor U12220 (N_12220,N_11904,N_11838);
or U12221 (N_12221,N_11642,N_11576);
nand U12222 (N_12222,N_11739,N_11735);
nand U12223 (N_12223,N_11503,N_11908);
nand U12224 (N_12224,N_11647,N_11596);
nor U12225 (N_12225,N_11686,N_11514);
nor U12226 (N_12226,N_11856,N_11977);
or U12227 (N_12227,N_11597,N_11531);
and U12228 (N_12228,N_11863,N_11876);
or U12229 (N_12229,N_11846,N_11775);
nand U12230 (N_12230,N_11800,N_11614);
nand U12231 (N_12231,N_11831,N_11506);
nand U12232 (N_12232,N_11620,N_11690);
and U12233 (N_12233,N_11732,N_11720);
xor U12234 (N_12234,N_11897,N_11736);
or U12235 (N_12235,N_11558,N_11655);
and U12236 (N_12236,N_11822,N_11722);
nor U12237 (N_12237,N_11575,N_11902);
or U12238 (N_12238,N_11544,N_11713);
nor U12239 (N_12239,N_11579,N_11833);
or U12240 (N_12240,N_11906,N_11844);
nand U12241 (N_12241,N_11974,N_11689);
and U12242 (N_12242,N_11845,N_11959);
nand U12243 (N_12243,N_11638,N_11665);
nor U12244 (N_12244,N_11861,N_11901);
nand U12245 (N_12245,N_11870,N_11715);
xor U12246 (N_12246,N_11759,N_11682);
nand U12247 (N_12247,N_11968,N_11942);
and U12248 (N_12248,N_11903,N_11571);
nor U12249 (N_12249,N_11927,N_11830);
nor U12250 (N_12250,N_11545,N_11728);
nor U12251 (N_12251,N_11633,N_11901);
or U12252 (N_12252,N_11832,N_11771);
and U12253 (N_12253,N_11898,N_11820);
and U12254 (N_12254,N_11774,N_11871);
xnor U12255 (N_12255,N_11533,N_11684);
xor U12256 (N_12256,N_11768,N_11868);
or U12257 (N_12257,N_11774,N_11504);
and U12258 (N_12258,N_11695,N_11681);
nand U12259 (N_12259,N_11907,N_11625);
nand U12260 (N_12260,N_11639,N_11567);
or U12261 (N_12261,N_11794,N_11903);
nand U12262 (N_12262,N_11798,N_11568);
xor U12263 (N_12263,N_11607,N_11755);
xnor U12264 (N_12264,N_11541,N_11844);
or U12265 (N_12265,N_11609,N_11537);
or U12266 (N_12266,N_11588,N_11733);
nor U12267 (N_12267,N_11604,N_11944);
nand U12268 (N_12268,N_11689,N_11538);
xnor U12269 (N_12269,N_11584,N_11969);
xnor U12270 (N_12270,N_11683,N_11541);
and U12271 (N_12271,N_11936,N_11541);
nor U12272 (N_12272,N_11675,N_11680);
and U12273 (N_12273,N_11691,N_11594);
or U12274 (N_12274,N_11620,N_11873);
or U12275 (N_12275,N_11844,N_11890);
nand U12276 (N_12276,N_11571,N_11559);
nor U12277 (N_12277,N_11831,N_11948);
or U12278 (N_12278,N_11835,N_11589);
xor U12279 (N_12279,N_11528,N_11891);
nand U12280 (N_12280,N_11856,N_11971);
xor U12281 (N_12281,N_11728,N_11707);
xnor U12282 (N_12282,N_11538,N_11632);
or U12283 (N_12283,N_11540,N_11718);
and U12284 (N_12284,N_11780,N_11631);
and U12285 (N_12285,N_11637,N_11717);
nor U12286 (N_12286,N_11836,N_11777);
or U12287 (N_12287,N_11965,N_11643);
nor U12288 (N_12288,N_11507,N_11803);
or U12289 (N_12289,N_11636,N_11688);
xnor U12290 (N_12290,N_11932,N_11591);
nor U12291 (N_12291,N_11950,N_11835);
and U12292 (N_12292,N_11672,N_11837);
nor U12293 (N_12293,N_11609,N_11758);
or U12294 (N_12294,N_11911,N_11592);
nand U12295 (N_12295,N_11998,N_11987);
nor U12296 (N_12296,N_11857,N_11513);
nand U12297 (N_12297,N_11917,N_11564);
nor U12298 (N_12298,N_11717,N_11705);
xnor U12299 (N_12299,N_11759,N_11544);
and U12300 (N_12300,N_11722,N_11823);
or U12301 (N_12301,N_11721,N_11949);
and U12302 (N_12302,N_11999,N_11518);
and U12303 (N_12303,N_11895,N_11604);
and U12304 (N_12304,N_11802,N_11720);
or U12305 (N_12305,N_11798,N_11815);
and U12306 (N_12306,N_11681,N_11626);
and U12307 (N_12307,N_11509,N_11540);
nor U12308 (N_12308,N_11704,N_11720);
xnor U12309 (N_12309,N_11804,N_11504);
and U12310 (N_12310,N_11921,N_11700);
and U12311 (N_12311,N_11754,N_11700);
and U12312 (N_12312,N_11515,N_11814);
nand U12313 (N_12313,N_11611,N_11674);
and U12314 (N_12314,N_11661,N_11869);
or U12315 (N_12315,N_11601,N_11640);
and U12316 (N_12316,N_11577,N_11617);
and U12317 (N_12317,N_11529,N_11737);
nor U12318 (N_12318,N_11948,N_11525);
or U12319 (N_12319,N_11500,N_11502);
or U12320 (N_12320,N_11839,N_11955);
nand U12321 (N_12321,N_11936,N_11509);
nand U12322 (N_12322,N_11638,N_11535);
xnor U12323 (N_12323,N_11545,N_11974);
xnor U12324 (N_12324,N_11526,N_11735);
or U12325 (N_12325,N_11762,N_11590);
nand U12326 (N_12326,N_11541,N_11860);
nor U12327 (N_12327,N_11716,N_11661);
or U12328 (N_12328,N_11606,N_11710);
nand U12329 (N_12329,N_11827,N_11772);
nand U12330 (N_12330,N_11847,N_11991);
nand U12331 (N_12331,N_11998,N_11677);
or U12332 (N_12332,N_11961,N_11632);
and U12333 (N_12333,N_11823,N_11776);
xor U12334 (N_12334,N_11548,N_11625);
xor U12335 (N_12335,N_11983,N_11609);
nor U12336 (N_12336,N_11591,N_11581);
and U12337 (N_12337,N_11902,N_11514);
and U12338 (N_12338,N_11579,N_11519);
and U12339 (N_12339,N_11810,N_11636);
nor U12340 (N_12340,N_11771,N_11554);
xor U12341 (N_12341,N_11840,N_11543);
nand U12342 (N_12342,N_11794,N_11739);
nor U12343 (N_12343,N_11821,N_11559);
and U12344 (N_12344,N_11748,N_11562);
xor U12345 (N_12345,N_11779,N_11727);
xor U12346 (N_12346,N_11709,N_11803);
or U12347 (N_12347,N_11672,N_11997);
or U12348 (N_12348,N_11611,N_11841);
nand U12349 (N_12349,N_11512,N_11975);
nor U12350 (N_12350,N_11509,N_11923);
nand U12351 (N_12351,N_11880,N_11801);
xnor U12352 (N_12352,N_11857,N_11771);
xnor U12353 (N_12353,N_11955,N_11767);
nand U12354 (N_12354,N_11846,N_11854);
nand U12355 (N_12355,N_11662,N_11731);
nand U12356 (N_12356,N_11750,N_11653);
nor U12357 (N_12357,N_11878,N_11871);
nor U12358 (N_12358,N_11788,N_11830);
and U12359 (N_12359,N_11831,N_11676);
nor U12360 (N_12360,N_11529,N_11519);
xnor U12361 (N_12361,N_11527,N_11728);
or U12362 (N_12362,N_11909,N_11670);
and U12363 (N_12363,N_11817,N_11996);
and U12364 (N_12364,N_11569,N_11677);
nor U12365 (N_12365,N_11897,N_11978);
nand U12366 (N_12366,N_11863,N_11626);
nand U12367 (N_12367,N_11654,N_11750);
xnor U12368 (N_12368,N_11896,N_11776);
xnor U12369 (N_12369,N_11749,N_11571);
xor U12370 (N_12370,N_11720,N_11795);
xnor U12371 (N_12371,N_11506,N_11512);
nor U12372 (N_12372,N_11727,N_11781);
nand U12373 (N_12373,N_11759,N_11785);
and U12374 (N_12374,N_11518,N_11907);
and U12375 (N_12375,N_11673,N_11909);
xor U12376 (N_12376,N_11765,N_11921);
nand U12377 (N_12377,N_11904,N_11749);
xnor U12378 (N_12378,N_11812,N_11810);
and U12379 (N_12379,N_11791,N_11623);
or U12380 (N_12380,N_11722,N_11584);
or U12381 (N_12381,N_11558,N_11716);
nor U12382 (N_12382,N_11669,N_11824);
or U12383 (N_12383,N_11598,N_11642);
and U12384 (N_12384,N_11874,N_11691);
nand U12385 (N_12385,N_11699,N_11605);
or U12386 (N_12386,N_11500,N_11880);
nand U12387 (N_12387,N_11964,N_11837);
or U12388 (N_12388,N_11767,N_11775);
nor U12389 (N_12389,N_11849,N_11949);
xor U12390 (N_12390,N_11527,N_11913);
nand U12391 (N_12391,N_11818,N_11978);
and U12392 (N_12392,N_11983,N_11927);
nor U12393 (N_12393,N_11675,N_11644);
or U12394 (N_12394,N_11901,N_11731);
and U12395 (N_12395,N_11806,N_11640);
or U12396 (N_12396,N_11957,N_11863);
nor U12397 (N_12397,N_11620,N_11676);
or U12398 (N_12398,N_11572,N_11508);
and U12399 (N_12399,N_11801,N_11521);
xnor U12400 (N_12400,N_11926,N_11722);
xor U12401 (N_12401,N_11948,N_11805);
and U12402 (N_12402,N_11640,N_11924);
xnor U12403 (N_12403,N_11546,N_11640);
and U12404 (N_12404,N_11802,N_11976);
xor U12405 (N_12405,N_11544,N_11911);
or U12406 (N_12406,N_11900,N_11699);
or U12407 (N_12407,N_11742,N_11952);
nor U12408 (N_12408,N_11671,N_11551);
or U12409 (N_12409,N_11516,N_11872);
xor U12410 (N_12410,N_11793,N_11690);
and U12411 (N_12411,N_11516,N_11703);
or U12412 (N_12412,N_11915,N_11673);
nor U12413 (N_12413,N_11893,N_11700);
and U12414 (N_12414,N_11592,N_11618);
xor U12415 (N_12415,N_11895,N_11570);
or U12416 (N_12416,N_11575,N_11939);
nand U12417 (N_12417,N_11585,N_11876);
nor U12418 (N_12418,N_11880,N_11709);
nand U12419 (N_12419,N_11950,N_11876);
or U12420 (N_12420,N_11547,N_11696);
and U12421 (N_12421,N_11525,N_11973);
nor U12422 (N_12422,N_11570,N_11733);
nor U12423 (N_12423,N_11780,N_11520);
nor U12424 (N_12424,N_11684,N_11826);
and U12425 (N_12425,N_11585,N_11862);
nand U12426 (N_12426,N_11955,N_11642);
xor U12427 (N_12427,N_11927,N_11794);
nor U12428 (N_12428,N_11873,N_11697);
nand U12429 (N_12429,N_11693,N_11659);
nor U12430 (N_12430,N_11501,N_11573);
and U12431 (N_12431,N_11617,N_11641);
and U12432 (N_12432,N_11702,N_11619);
xnor U12433 (N_12433,N_11557,N_11589);
nand U12434 (N_12434,N_11537,N_11695);
nor U12435 (N_12435,N_11701,N_11861);
nand U12436 (N_12436,N_11854,N_11900);
nor U12437 (N_12437,N_11949,N_11553);
nor U12438 (N_12438,N_11831,N_11638);
and U12439 (N_12439,N_11758,N_11680);
xor U12440 (N_12440,N_11960,N_11904);
xnor U12441 (N_12441,N_11746,N_11891);
or U12442 (N_12442,N_11658,N_11814);
or U12443 (N_12443,N_11528,N_11828);
nand U12444 (N_12444,N_11742,N_11553);
and U12445 (N_12445,N_11749,N_11645);
or U12446 (N_12446,N_11925,N_11911);
or U12447 (N_12447,N_11635,N_11931);
or U12448 (N_12448,N_11779,N_11929);
nand U12449 (N_12449,N_11913,N_11845);
nand U12450 (N_12450,N_11821,N_11989);
and U12451 (N_12451,N_11598,N_11691);
or U12452 (N_12452,N_11914,N_11558);
nor U12453 (N_12453,N_11720,N_11678);
or U12454 (N_12454,N_11646,N_11538);
nand U12455 (N_12455,N_11884,N_11530);
and U12456 (N_12456,N_11746,N_11887);
and U12457 (N_12457,N_11629,N_11879);
or U12458 (N_12458,N_11551,N_11651);
xnor U12459 (N_12459,N_11968,N_11548);
and U12460 (N_12460,N_11814,N_11783);
xor U12461 (N_12461,N_11875,N_11672);
xnor U12462 (N_12462,N_11577,N_11621);
and U12463 (N_12463,N_11854,N_11890);
nand U12464 (N_12464,N_11778,N_11908);
xor U12465 (N_12465,N_11696,N_11729);
nor U12466 (N_12466,N_11966,N_11958);
nand U12467 (N_12467,N_11513,N_11842);
xor U12468 (N_12468,N_11974,N_11927);
or U12469 (N_12469,N_11993,N_11647);
nor U12470 (N_12470,N_11613,N_11700);
nor U12471 (N_12471,N_11897,N_11513);
nand U12472 (N_12472,N_11969,N_11785);
xor U12473 (N_12473,N_11857,N_11706);
or U12474 (N_12474,N_11524,N_11952);
or U12475 (N_12475,N_11501,N_11602);
nor U12476 (N_12476,N_11720,N_11823);
nor U12477 (N_12477,N_11787,N_11725);
xnor U12478 (N_12478,N_11778,N_11790);
xnor U12479 (N_12479,N_11511,N_11854);
or U12480 (N_12480,N_11743,N_11681);
nor U12481 (N_12481,N_11981,N_11931);
xnor U12482 (N_12482,N_11753,N_11918);
or U12483 (N_12483,N_11735,N_11642);
or U12484 (N_12484,N_11629,N_11786);
nand U12485 (N_12485,N_11553,N_11814);
or U12486 (N_12486,N_11665,N_11568);
nor U12487 (N_12487,N_11877,N_11951);
nor U12488 (N_12488,N_11981,N_11882);
or U12489 (N_12489,N_11774,N_11776);
nor U12490 (N_12490,N_11750,N_11540);
nor U12491 (N_12491,N_11892,N_11780);
xor U12492 (N_12492,N_11798,N_11551);
xnor U12493 (N_12493,N_11965,N_11675);
or U12494 (N_12494,N_11607,N_11940);
xor U12495 (N_12495,N_11720,N_11898);
nor U12496 (N_12496,N_11917,N_11612);
or U12497 (N_12497,N_11928,N_11720);
nor U12498 (N_12498,N_11760,N_11660);
and U12499 (N_12499,N_11546,N_11725);
xnor U12500 (N_12500,N_12122,N_12276);
and U12501 (N_12501,N_12283,N_12065);
xnor U12502 (N_12502,N_12129,N_12491);
or U12503 (N_12503,N_12192,N_12001);
nand U12504 (N_12504,N_12102,N_12105);
or U12505 (N_12505,N_12115,N_12238);
nand U12506 (N_12506,N_12255,N_12052);
nand U12507 (N_12507,N_12304,N_12332);
nor U12508 (N_12508,N_12143,N_12068);
nand U12509 (N_12509,N_12013,N_12070);
xor U12510 (N_12510,N_12084,N_12054);
or U12511 (N_12511,N_12447,N_12412);
xor U12512 (N_12512,N_12214,N_12027);
or U12513 (N_12513,N_12226,N_12346);
and U12514 (N_12514,N_12212,N_12152);
xnor U12515 (N_12515,N_12133,N_12179);
and U12516 (N_12516,N_12303,N_12337);
nor U12517 (N_12517,N_12082,N_12480);
xor U12518 (N_12518,N_12302,N_12374);
xnor U12519 (N_12519,N_12221,N_12058);
or U12520 (N_12520,N_12063,N_12009);
nand U12521 (N_12521,N_12430,N_12003);
xor U12522 (N_12522,N_12112,N_12395);
and U12523 (N_12523,N_12316,N_12484);
and U12524 (N_12524,N_12467,N_12217);
or U12525 (N_12525,N_12089,N_12064);
xor U12526 (N_12526,N_12388,N_12023);
xor U12527 (N_12527,N_12146,N_12470);
and U12528 (N_12528,N_12477,N_12130);
and U12529 (N_12529,N_12178,N_12140);
nand U12530 (N_12530,N_12116,N_12088);
nand U12531 (N_12531,N_12478,N_12229);
nand U12532 (N_12532,N_12244,N_12322);
and U12533 (N_12533,N_12021,N_12028);
and U12534 (N_12534,N_12160,N_12444);
xor U12535 (N_12535,N_12440,N_12072);
xor U12536 (N_12536,N_12326,N_12461);
nand U12537 (N_12537,N_12149,N_12465);
or U12538 (N_12538,N_12053,N_12452);
nor U12539 (N_12539,N_12279,N_12370);
or U12540 (N_12540,N_12498,N_12085);
xnor U12541 (N_12541,N_12010,N_12131);
xor U12542 (N_12542,N_12142,N_12284);
xor U12543 (N_12543,N_12016,N_12004);
nor U12544 (N_12544,N_12067,N_12442);
nor U12545 (N_12545,N_12181,N_12017);
nor U12546 (N_12546,N_12485,N_12047);
nor U12547 (N_12547,N_12489,N_12005);
nor U12548 (N_12548,N_12087,N_12367);
and U12549 (N_12549,N_12301,N_12051);
xor U12550 (N_12550,N_12231,N_12358);
and U12551 (N_12551,N_12331,N_12459);
and U12552 (N_12552,N_12202,N_12096);
or U12553 (N_12553,N_12435,N_12425);
nor U12554 (N_12554,N_12039,N_12032);
nor U12555 (N_12555,N_12166,N_12030);
nor U12556 (N_12556,N_12278,N_12482);
and U12557 (N_12557,N_12111,N_12277);
or U12558 (N_12558,N_12090,N_12256);
or U12559 (N_12559,N_12134,N_12205);
nand U12560 (N_12560,N_12315,N_12294);
or U12561 (N_12561,N_12191,N_12135);
and U12562 (N_12562,N_12250,N_12300);
nor U12563 (N_12563,N_12055,N_12247);
or U12564 (N_12564,N_12488,N_12138);
nor U12565 (N_12565,N_12376,N_12394);
nand U12566 (N_12566,N_12443,N_12445);
xor U12567 (N_12567,N_12069,N_12264);
xnor U12568 (N_12568,N_12479,N_12185);
or U12569 (N_12569,N_12455,N_12237);
nand U12570 (N_12570,N_12210,N_12310);
and U12571 (N_12571,N_12392,N_12495);
nor U12572 (N_12572,N_12168,N_12363);
xor U12573 (N_12573,N_12271,N_12057);
or U12574 (N_12574,N_12422,N_12014);
or U12575 (N_12575,N_12432,N_12319);
nand U12576 (N_12576,N_12081,N_12383);
nor U12577 (N_12577,N_12073,N_12273);
or U12578 (N_12578,N_12213,N_12171);
xnor U12579 (N_12579,N_12106,N_12145);
nor U12580 (N_12580,N_12311,N_12243);
and U12581 (N_12581,N_12078,N_12126);
and U12582 (N_12582,N_12233,N_12163);
nand U12583 (N_12583,N_12196,N_12483);
or U12584 (N_12584,N_12409,N_12263);
or U12585 (N_12585,N_12037,N_12492);
or U12586 (N_12586,N_12416,N_12093);
xor U12587 (N_12587,N_12353,N_12026);
nor U12588 (N_12588,N_12306,N_12359);
or U12589 (N_12589,N_12463,N_12282);
or U12590 (N_12590,N_12270,N_12469);
and U12591 (N_12591,N_12289,N_12448);
or U12592 (N_12592,N_12399,N_12352);
nor U12593 (N_12593,N_12297,N_12329);
or U12594 (N_12594,N_12471,N_12476);
or U12595 (N_12595,N_12313,N_12012);
nor U12596 (N_12596,N_12060,N_12103);
nor U12597 (N_12597,N_12187,N_12481);
or U12598 (N_12598,N_12104,N_12338);
and U12599 (N_12599,N_12259,N_12373);
xnor U12600 (N_12600,N_12219,N_12147);
nand U12601 (N_12601,N_12274,N_12265);
xor U12602 (N_12602,N_12426,N_12074);
and U12603 (N_12603,N_12195,N_12366);
or U12604 (N_12604,N_12019,N_12101);
xor U12605 (N_12605,N_12439,N_12071);
xnor U12606 (N_12606,N_12132,N_12401);
and U12607 (N_12607,N_12288,N_12473);
or U12608 (N_12608,N_12197,N_12257);
nor U12609 (N_12609,N_12371,N_12127);
nor U12610 (N_12610,N_12049,N_12204);
and U12611 (N_12611,N_12113,N_12266);
nand U12612 (N_12612,N_12232,N_12268);
or U12613 (N_12613,N_12299,N_12043);
and U12614 (N_12614,N_12296,N_12086);
xor U12615 (N_12615,N_12364,N_12227);
nor U12616 (N_12616,N_12177,N_12453);
xor U12617 (N_12617,N_12059,N_12208);
xnor U12618 (N_12618,N_12354,N_12050);
xor U12619 (N_12619,N_12080,N_12083);
nand U12620 (N_12620,N_12228,N_12345);
or U12621 (N_12621,N_12397,N_12293);
xor U12622 (N_12622,N_12100,N_12262);
nand U12623 (N_12623,N_12493,N_12114);
and U12624 (N_12624,N_12333,N_12025);
nor U12625 (N_12625,N_12184,N_12155);
xnor U12626 (N_12626,N_12437,N_12117);
and U12627 (N_12627,N_12123,N_12144);
nor U12628 (N_12628,N_12159,N_12029);
nor U12629 (N_12629,N_12077,N_12380);
nand U12630 (N_12630,N_12061,N_12251);
or U12631 (N_12631,N_12218,N_12006);
xor U12632 (N_12632,N_12234,N_12391);
xnor U12633 (N_12633,N_12245,N_12389);
nor U12634 (N_12634,N_12407,N_12167);
xnor U12635 (N_12635,N_12375,N_12235);
or U12636 (N_12636,N_12421,N_12169);
nor U12637 (N_12637,N_12230,N_12285);
and U12638 (N_12638,N_12406,N_12324);
nand U12639 (N_12639,N_12434,N_12468);
nor U12640 (N_12640,N_12487,N_12361);
xor U12641 (N_12641,N_12258,N_12109);
nand U12642 (N_12642,N_12041,N_12206);
or U12643 (N_12643,N_12048,N_12327);
nand U12644 (N_12644,N_12239,N_12120);
or U12645 (N_12645,N_12330,N_12248);
or U12646 (N_12646,N_12249,N_12173);
or U12647 (N_12647,N_12280,N_12454);
nand U12648 (N_12648,N_12308,N_12497);
nand U12649 (N_12649,N_12355,N_12305);
nor U12650 (N_12650,N_12220,N_12141);
nor U12651 (N_12651,N_12099,N_12404);
or U12652 (N_12652,N_12449,N_12224);
and U12653 (N_12653,N_12044,N_12349);
nand U12654 (N_12654,N_12351,N_12098);
and U12655 (N_12655,N_12314,N_12151);
nand U12656 (N_12656,N_12034,N_12203);
and U12657 (N_12657,N_12446,N_12387);
or U12658 (N_12658,N_12298,N_12036);
xor U12659 (N_12659,N_12292,N_12198);
nand U12660 (N_12660,N_12170,N_12040);
and U12661 (N_12661,N_12225,N_12024);
xnor U12662 (N_12662,N_12420,N_12403);
xnor U12663 (N_12663,N_12460,N_12415);
nor U12664 (N_12664,N_12408,N_12119);
nor U12665 (N_12665,N_12200,N_12417);
nand U12666 (N_12666,N_12433,N_12287);
nand U12667 (N_12667,N_12382,N_12148);
nand U12668 (N_12668,N_12431,N_12405);
or U12669 (N_12669,N_12475,N_12121);
or U12670 (N_12670,N_12398,N_12325);
nor U12671 (N_12671,N_12118,N_12318);
nor U12672 (N_12672,N_12261,N_12400);
or U12673 (N_12673,N_12496,N_12348);
nor U12674 (N_12674,N_12384,N_12267);
xnor U12675 (N_12675,N_12194,N_12396);
and U12676 (N_12676,N_12031,N_12153);
xor U12677 (N_12677,N_12079,N_12334);
or U12678 (N_12678,N_12182,N_12342);
xor U12679 (N_12679,N_12457,N_12386);
nand U12680 (N_12680,N_12428,N_12362);
xor U12681 (N_12681,N_12490,N_12253);
and U12682 (N_12682,N_12360,N_12207);
or U12683 (N_12683,N_12175,N_12161);
xor U12684 (N_12684,N_12494,N_12464);
and U12685 (N_12685,N_12260,N_12472);
or U12686 (N_12686,N_12336,N_12307);
nand U12687 (N_12687,N_12008,N_12357);
and U12688 (N_12688,N_12164,N_12002);
or U12689 (N_12689,N_12450,N_12107);
or U12690 (N_12690,N_12372,N_12419);
or U12691 (N_12691,N_12018,N_12042);
xnor U12692 (N_12692,N_12189,N_12393);
nand U12693 (N_12693,N_12411,N_12413);
nand U12694 (N_12694,N_12223,N_12022);
or U12695 (N_12695,N_12451,N_12124);
and U12696 (N_12696,N_12154,N_12436);
or U12697 (N_12697,N_12272,N_12075);
xor U12698 (N_12698,N_12246,N_12240);
nand U12699 (N_12699,N_12209,N_12377);
and U12700 (N_12700,N_12418,N_12254);
nor U12701 (N_12701,N_12091,N_12344);
xnor U12702 (N_12702,N_12328,N_12176);
or U12703 (N_12703,N_12410,N_12312);
xnor U12704 (N_12704,N_12158,N_12424);
xnor U12705 (N_12705,N_12020,N_12015);
nor U12706 (N_12706,N_12381,N_12056);
xnor U12707 (N_12707,N_12365,N_12295);
nor U12708 (N_12708,N_12341,N_12222);
or U12709 (N_12709,N_12462,N_12286);
nor U12710 (N_12710,N_12199,N_12190);
xnor U12711 (N_12711,N_12320,N_12188);
and U12712 (N_12712,N_12139,N_12499);
nand U12713 (N_12713,N_12035,N_12242);
and U12714 (N_12714,N_12137,N_12339);
nor U12715 (N_12715,N_12157,N_12066);
nand U12716 (N_12716,N_12429,N_12108);
xnor U12717 (N_12717,N_12046,N_12456);
nor U12718 (N_12718,N_12290,N_12281);
and U12719 (N_12719,N_12165,N_12172);
or U12720 (N_12720,N_12347,N_12156);
xnor U12721 (N_12721,N_12215,N_12458);
nor U12722 (N_12722,N_12216,N_12174);
xnor U12723 (N_12723,N_12241,N_12486);
xnor U12724 (N_12724,N_12275,N_12125);
nor U12725 (N_12725,N_12466,N_12201);
nand U12726 (N_12726,N_12097,N_12356);
nand U12727 (N_12727,N_12180,N_12000);
and U12728 (N_12728,N_12309,N_12186);
nand U12729 (N_12729,N_12438,N_12269);
nand U12730 (N_12730,N_12402,N_12369);
nor U12731 (N_12731,N_12076,N_12414);
and U12732 (N_12732,N_12162,N_12423);
xor U12733 (N_12733,N_12011,N_12390);
nand U12734 (N_12734,N_12323,N_12378);
and U12735 (N_12735,N_12062,N_12033);
xor U12736 (N_12736,N_12045,N_12427);
nand U12737 (N_12737,N_12474,N_12321);
or U12738 (N_12738,N_12092,N_12441);
and U12739 (N_12739,N_12094,N_12150);
or U12740 (N_12740,N_12379,N_12007);
nand U12741 (N_12741,N_12128,N_12350);
and U12742 (N_12742,N_12183,N_12335);
and U12743 (N_12743,N_12317,N_12236);
nor U12744 (N_12744,N_12038,N_12136);
and U12745 (N_12745,N_12252,N_12291);
and U12746 (N_12746,N_12343,N_12340);
nor U12747 (N_12747,N_12211,N_12368);
nor U12748 (N_12748,N_12110,N_12095);
or U12749 (N_12749,N_12193,N_12385);
xor U12750 (N_12750,N_12057,N_12495);
and U12751 (N_12751,N_12215,N_12315);
xor U12752 (N_12752,N_12317,N_12084);
and U12753 (N_12753,N_12080,N_12204);
xnor U12754 (N_12754,N_12411,N_12002);
xnor U12755 (N_12755,N_12230,N_12493);
or U12756 (N_12756,N_12403,N_12395);
or U12757 (N_12757,N_12186,N_12459);
and U12758 (N_12758,N_12085,N_12173);
or U12759 (N_12759,N_12076,N_12352);
xnor U12760 (N_12760,N_12201,N_12196);
or U12761 (N_12761,N_12423,N_12138);
and U12762 (N_12762,N_12016,N_12206);
and U12763 (N_12763,N_12043,N_12045);
nand U12764 (N_12764,N_12176,N_12157);
or U12765 (N_12765,N_12220,N_12181);
nor U12766 (N_12766,N_12359,N_12264);
nand U12767 (N_12767,N_12466,N_12193);
or U12768 (N_12768,N_12171,N_12097);
and U12769 (N_12769,N_12301,N_12247);
or U12770 (N_12770,N_12175,N_12471);
nor U12771 (N_12771,N_12486,N_12283);
and U12772 (N_12772,N_12061,N_12262);
nor U12773 (N_12773,N_12136,N_12009);
nand U12774 (N_12774,N_12002,N_12236);
or U12775 (N_12775,N_12285,N_12265);
nor U12776 (N_12776,N_12331,N_12247);
xnor U12777 (N_12777,N_12276,N_12135);
nor U12778 (N_12778,N_12129,N_12394);
nand U12779 (N_12779,N_12341,N_12169);
nand U12780 (N_12780,N_12378,N_12085);
nand U12781 (N_12781,N_12420,N_12349);
xnor U12782 (N_12782,N_12040,N_12387);
or U12783 (N_12783,N_12268,N_12027);
nor U12784 (N_12784,N_12446,N_12482);
or U12785 (N_12785,N_12256,N_12037);
or U12786 (N_12786,N_12375,N_12367);
nand U12787 (N_12787,N_12398,N_12218);
nand U12788 (N_12788,N_12033,N_12147);
nor U12789 (N_12789,N_12265,N_12485);
nor U12790 (N_12790,N_12347,N_12001);
nor U12791 (N_12791,N_12374,N_12207);
nor U12792 (N_12792,N_12369,N_12268);
or U12793 (N_12793,N_12212,N_12089);
and U12794 (N_12794,N_12465,N_12492);
xor U12795 (N_12795,N_12188,N_12401);
xor U12796 (N_12796,N_12018,N_12193);
nand U12797 (N_12797,N_12317,N_12108);
xnor U12798 (N_12798,N_12058,N_12114);
and U12799 (N_12799,N_12291,N_12470);
and U12800 (N_12800,N_12371,N_12345);
or U12801 (N_12801,N_12256,N_12491);
nor U12802 (N_12802,N_12386,N_12265);
and U12803 (N_12803,N_12269,N_12156);
xor U12804 (N_12804,N_12475,N_12031);
xor U12805 (N_12805,N_12440,N_12426);
or U12806 (N_12806,N_12024,N_12236);
nor U12807 (N_12807,N_12397,N_12059);
nor U12808 (N_12808,N_12401,N_12219);
and U12809 (N_12809,N_12143,N_12044);
nand U12810 (N_12810,N_12307,N_12449);
nand U12811 (N_12811,N_12287,N_12104);
or U12812 (N_12812,N_12194,N_12452);
xnor U12813 (N_12813,N_12053,N_12189);
nand U12814 (N_12814,N_12201,N_12465);
and U12815 (N_12815,N_12491,N_12150);
xor U12816 (N_12816,N_12162,N_12260);
or U12817 (N_12817,N_12177,N_12371);
nand U12818 (N_12818,N_12173,N_12020);
xnor U12819 (N_12819,N_12460,N_12096);
or U12820 (N_12820,N_12000,N_12260);
nand U12821 (N_12821,N_12249,N_12135);
xor U12822 (N_12822,N_12165,N_12470);
nor U12823 (N_12823,N_12080,N_12019);
xor U12824 (N_12824,N_12379,N_12243);
nor U12825 (N_12825,N_12083,N_12419);
xor U12826 (N_12826,N_12210,N_12163);
and U12827 (N_12827,N_12065,N_12027);
nand U12828 (N_12828,N_12155,N_12194);
or U12829 (N_12829,N_12101,N_12116);
xnor U12830 (N_12830,N_12164,N_12165);
xnor U12831 (N_12831,N_12065,N_12287);
and U12832 (N_12832,N_12019,N_12414);
nor U12833 (N_12833,N_12081,N_12322);
and U12834 (N_12834,N_12359,N_12476);
and U12835 (N_12835,N_12440,N_12336);
or U12836 (N_12836,N_12356,N_12295);
and U12837 (N_12837,N_12143,N_12260);
and U12838 (N_12838,N_12082,N_12153);
or U12839 (N_12839,N_12446,N_12124);
xor U12840 (N_12840,N_12338,N_12406);
or U12841 (N_12841,N_12147,N_12074);
nand U12842 (N_12842,N_12028,N_12132);
nor U12843 (N_12843,N_12467,N_12398);
xor U12844 (N_12844,N_12384,N_12319);
and U12845 (N_12845,N_12361,N_12272);
and U12846 (N_12846,N_12020,N_12483);
xnor U12847 (N_12847,N_12003,N_12425);
or U12848 (N_12848,N_12354,N_12218);
xor U12849 (N_12849,N_12301,N_12356);
or U12850 (N_12850,N_12068,N_12315);
or U12851 (N_12851,N_12268,N_12013);
nor U12852 (N_12852,N_12012,N_12417);
xor U12853 (N_12853,N_12498,N_12342);
and U12854 (N_12854,N_12187,N_12282);
or U12855 (N_12855,N_12362,N_12443);
and U12856 (N_12856,N_12126,N_12248);
xor U12857 (N_12857,N_12257,N_12015);
nand U12858 (N_12858,N_12343,N_12264);
nor U12859 (N_12859,N_12328,N_12324);
and U12860 (N_12860,N_12443,N_12185);
and U12861 (N_12861,N_12427,N_12193);
nor U12862 (N_12862,N_12165,N_12494);
xnor U12863 (N_12863,N_12453,N_12261);
xnor U12864 (N_12864,N_12369,N_12032);
nand U12865 (N_12865,N_12010,N_12181);
nor U12866 (N_12866,N_12005,N_12181);
nor U12867 (N_12867,N_12015,N_12238);
nor U12868 (N_12868,N_12492,N_12191);
and U12869 (N_12869,N_12482,N_12000);
and U12870 (N_12870,N_12455,N_12408);
and U12871 (N_12871,N_12449,N_12370);
nand U12872 (N_12872,N_12062,N_12402);
nor U12873 (N_12873,N_12366,N_12030);
and U12874 (N_12874,N_12489,N_12145);
and U12875 (N_12875,N_12214,N_12290);
and U12876 (N_12876,N_12055,N_12465);
xnor U12877 (N_12877,N_12259,N_12276);
nor U12878 (N_12878,N_12141,N_12170);
nor U12879 (N_12879,N_12315,N_12409);
nand U12880 (N_12880,N_12393,N_12402);
or U12881 (N_12881,N_12314,N_12358);
xor U12882 (N_12882,N_12331,N_12321);
nand U12883 (N_12883,N_12325,N_12223);
nor U12884 (N_12884,N_12269,N_12352);
or U12885 (N_12885,N_12311,N_12005);
xor U12886 (N_12886,N_12352,N_12307);
xnor U12887 (N_12887,N_12442,N_12383);
xor U12888 (N_12888,N_12164,N_12296);
xor U12889 (N_12889,N_12270,N_12194);
nor U12890 (N_12890,N_12177,N_12276);
nand U12891 (N_12891,N_12042,N_12493);
nand U12892 (N_12892,N_12435,N_12332);
and U12893 (N_12893,N_12123,N_12105);
and U12894 (N_12894,N_12206,N_12495);
xnor U12895 (N_12895,N_12375,N_12061);
xor U12896 (N_12896,N_12379,N_12392);
and U12897 (N_12897,N_12310,N_12412);
and U12898 (N_12898,N_12468,N_12120);
xnor U12899 (N_12899,N_12428,N_12161);
nor U12900 (N_12900,N_12063,N_12072);
or U12901 (N_12901,N_12437,N_12041);
nor U12902 (N_12902,N_12045,N_12196);
nand U12903 (N_12903,N_12155,N_12423);
nand U12904 (N_12904,N_12040,N_12116);
xnor U12905 (N_12905,N_12385,N_12331);
and U12906 (N_12906,N_12151,N_12085);
xnor U12907 (N_12907,N_12205,N_12378);
or U12908 (N_12908,N_12475,N_12484);
and U12909 (N_12909,N_12425,N_12235);
and U12910 (N_12910,N_12325,N_12495);
or U12911 (N_12911,N_12213,N_12223);
xor U12912 (N_12912,N_12311,N_12414);
or U12913 (N_12913,N_12044,N_12090);
and U12914 (N_12914,N_12016,N_12349);
nand U12915 (N_12915,N_12441,N_12079);
and U12916 (N_12916,N_12146,N_12208);
nand U12917 (N_12917,N_12071,N_12045);
or U12918 (N_12918,N_12485,N_12434);
xor U12919 (N_12919,N_12062,N_12377);
and U12920 (N_12920,N_12156,N_12246);
xnor U12921 (N_12921,N_12441,N_12078);
or U12922 (N_12922,N_12025,N_12390);
or U12923 (N_12923,N_12103,N_12005);
and U12924 (N_12924,N_12029,N_12489);
and U12925 (N_12925,N_12194,N_12148);
and U12926 (N_12926,N_12019,N_12283);
or U12927 (N_12927,N_12096,N_12446);
and U12928 (N_12928,N_12029,N_12037);
and U12929 (N_12929,N_12101,N_12211);
nand U12930 (N_12930,N_12109,N_12218);
xnor U12931 (N_12931,N_12337,N_12080);
and U12932 (N_12932,N_12042,N_12456);
xor U12933 (N_12933,N_12187,N_12145);
xnor U12934 (N_12934,N_12435,N_12478);
nor U12935 (N_12935,N_12286,N_12235);
xnor U12936 (N_12936,N_12449,N_12004);
nor U12937 (N_12937,N_12306,N_12446);
and U12938 (N_12938,N_12306,N_12158);
nand U12939 (N_12939,N_12220,N_12353);
or U12940 (N_12940,N_12495,N_12052);
nor U12941 (N_12941,N_12046,N_12335);
xnor U12942 (N_12942,N_12456,N_12459);
and U12943 (N_12943,N_12472,N_12232);
nand U12944 (N_12944,N_12413,N_12225);
and U12945 (N_12945,N_12364,N_12171);
xnor U12946 (N_12946,N_12302,N_12322);
nor U12947 (N_12947,N_12431,N_12400);
xor U12948 (N_12948,N_12101,N_12030);
xnor U12949 (N_12949,N_12308,N_12400);
nor U12950 (N_12950,N_12266,N_12359);
and U12951 (N_12951,N_12143,N_12365);
or U12952 (N_12952,N_12053,N_12047);
and U12953 (N_12953,N_12210,N_12355);
and U12954 (N_12954,N_12024,N_12287);
and U12955 (N_12955,N_12274,N_12183);
xnor U12956 (N_12956,N_12196,N_12271);
xnor U12957 (N_12957,N_12078,N_12437);
xnor U12958 (N_12958,N_12244,N_12151);
and U12959 (N_12959,N_12343,N_12303);
or U12960 (N_12960,N_12205,N_12013);
xor U12961 (N_12961,N_12017,N_12438);
xor U12962 (N_12962,N_12286,N_12000);
nand U12963 (N_12963,N_12133,N_12161);
or U12964 (N_12964,N_12273,N_12154);
or U12965 (N_12965,N_12023,N_12055);
or U12966 (N_12966,N_12420,N_12452);
or U12967 (N_12967,N_12415,N_12395);
xnor U12968 (N_12968,N_12432,N_12416);
nand U12969 (N_12969,N_12390,N_12388);
xor U12970 (N_12970,N_12453,N_12222);
nand U12971 (N_12971,N_12205,N_12119);
or U12972 (N_12972,N_12416,N_12000);
and U12973 (N_12973,N_12017,N_12436);
or U12974 (N_12974,N_12118,N_12329);
or U12975 (N_12975,N_12211,N_12168);
nor U12976 (N_12976,N_12297,N_12075);
and U12977 (N_12977,N_12063,N_12187);
or U12978 (N_12978,N_12343,N_12373);
nor U12979 (N_12979,N_12096,N_12235);
nor U12980 (N_12980,N_12291,N_12398);
nor U12981 (N_12981,N_12358,N_12494);
and U12982 (N_12982,N_12217,N_12341);
xnor U12983 (N_12983,N_12391,N_12136);
or U12984 (N_12984,N_12280,N_12165);
nand U12985 (N_12985,N_12245,N_12391);
or U12986 (N_12986,N_12055,N_12030);
nand U12987 (N_12987,N_12400,N_12045);
nor U12988 (N_12988,N_12199,N_12329);
xor U12989 (N_12989,N_12484,N_12169);
nor U12990 (N_12990,N_12453,N_12205);
and U12991 (N_12991,N_12255,N_12400);
and U12992 (N_12992,N_12176,N_12100);
and U12993 (N_12993,N_12173,N_12172);
and U12994 (N_12994,N_12048,N_12441);
xor U12995 (N_12995,N_12009,N_12092);
nor U12996 (N_12996,N_12388,N_12146);
xor U12997 (N_12997,N_12444,N_12477);
xnor U12998 (N_12998,N_12129,N_12352);
nor U12999 (N_12999,N_12249,N_12200);
nand U13000 (N_13000,N_12658,N_12589);
xnor U13001 (N_13001,N_12749,N_12574);
xor U13002 (N_13002,N_12513,N_12529);
xor U13003 (N_13003,N_12588,N_12794);
nor U13004 (N_13004,N_12910,N_12888);
nor U13005 (N_13005,N_12925,N_12986);
nor U13006 (N_13006,N_12772,N_12659);
nor U13007 (N_13007,N_12531,N_12859);
or U13008 (N_13008,N_12965,N_12846);
or U13009 (N_13009,N_12867,N_12510);
xnor U13010 (N_13010,N_12985,N_12792);
nand U13011 (N_13011,N_12676,N_12604);
nor U13012 (N_13012,N_12524,N_12569);
xnor U13013 (N_13013,N_12753,N_12603);
or U13014 (N_13014,N_12537,N_12801);
or U13015 (N_13015,N_12804,N_12864);
xnor U13016 (N_13016,N_12826,N_12972);
and U13017 (N_13017,N_12698,N_12626);
nor U13018 (N_13018,N_12543,N_12776);
or U13019 (N_13019,N_12692,N_12743);
and U13020 (N_13020,N_12863,N_12705);
nor U13021 (N_13021,N_12545,N_12530);
xor U13022 (N_13022,N_12670,N_12728);
nor U13023 (N_13023,N_12739,N_12982);
nor U13024 (N_13024,N_12605,N_12642);
or U13025 (N_13025,N_12517,N_12722);
and U13026 (N_13026,N_12766,N_12778);
xor U13027 (N_13027,N_12761,N_12756);
or U13028 (N_13028,N_12861,N_12704);
or U13029 (N_13029,N_12602,N_12909);
nand U13030 (N_13030,N_12702,N_12695);
xor U13031 (N_13031,N_12538,N_12686);
nor U13032 (N_13032,N_12587,N_12713);
nor U13033 (N_13033,N_12850,N_12539);
nand U13034 (N_13034,N_12503,N_12819);
xnor U13035 (N_13035,N_12979,N_12549);
nor U13036 (N_13036,N_12854,N_12601);
nor U13037 (N_13037,N_12842,N_12940);
xor U13038 (N_13038,N_12976,N_12565);
xor U13039 (N_13039,N_12662,N_12639);
nand U13040 (N_13040,N_12652,N_12783);
xor U13041 (N_13041,N_12696,N_12798);
nand U13042 (N_13042,N_12673,N_12532);
and U13043 (N_13043,N_12782,N_12526);
or U13044 (N_13044,N_12620,N_12777);
or U13045 (N_13045,N_12632,N_12664);
nor U13046 (N_13046,N_12520,N_12619);
or U13047 (N_13047,N_12715,N_12701);
xnor U13048 (N_13048,N_12806,N_12636);
and U13049 (N_13049,N_12727,N_12667);
and U13050 (N_13050,N_12820,N_12677);
and U13051 (N_13051,N_12546,N_12745);
and U13052 (N_13052,N_12596,N_12998);
or U13053 (N_13053,N_12915,N_12708);
nand U13054 (N_13054,N_12735,N_12822);
nand U13055 (N_13055,N_12580,N_12841);
nand U13056 (N_13056,N_12941,N_12577);
or U13057 (N_13057,N_12651,N_12871);
xnor U13058 (N_13058,N_12638,N_12895);
xor U13059 (N_13059,N_12991,N_12990);
or U13060 (N_13060,N_12599,N_12897);
or U13061 (N_13061,N_12898,N_12844);
xor U13062 (N_13062,N_12678,N_12614);
nor U13063 (N_13063,N_12679,N_12901);
nand U13064 (N_13064,N_12672,N_12875);
nand U13065 (N_13065,N_12827,N_12711);
xor U13066 (N_13066,N_12629,N_12784);
and U13067 (N_13067,N_12561,N_12916);
and U13068 (N_13068,N_12558,N_12879);
or U13069 (N_13069,N_12902,N_12641);
and U13070 (N_13070,N_12880,N_12855);
nand U13071 (N_13071,N_12942,N_12535);
nand U13072 (N_13072,N_12865,N_12911);
nand U13073 (N_13073,N_12928,N_12560);
nand U13074 (N_13074,N_12969,N_12576);
nor U13075 (N_13075,N_12866,N_12912);
and U13076 (N_13076,N_12694,N_12858);
nand U13077 (N_13077,N_12765,N_12683);
nor U13078 (N_13078,N_12750,N_12556);
and U13079 (N_13079,N_12689,N_12885);
xnor U13080 (N_13080,N_12829,N_12555);
nand U13081 (N_13081,N_12729,N_12790);
and U13082 (N_13082,N_12693,N_12697);
nand U13083 (N_13083,N_12807,N_12786);
or U13084 (N_13084,N_12548,N_12958);
and U13085 (N_13085,N_12547,N_12994);
xnor U13086 (N_13086,N_12892,N_12920);
and U13087 (N_13087,N_12917,N_12968);
nand U13088 (N_13088,N_12762,N_12824);
or U13089 (N_13089,N_12763,N_12980);
nor U13090 (N_13090,N_12734,N_12809);
and U13091 (N_13091,N_12950,N_12847);
xor U13092 (N_13092,N_12738,N_12868);
and U13093 (N_13093,N_12607,N_12703);
nand U13094 (N_13094,N_12506,N_12723);
or U13095 (N_13095,N_12802,N_12997);
nor U13096 (N_13096,N_12877,N_12624);
xor U13097 (N_13097,N_12685,N_12815);
nor U13098 (N_13098,N_12514,N_12852);
xnor U13099 (N_13099,N_12700,N_12592);
and U13100 (N_13100,N_12906,N_12907);
and U13101 (N_13101,N_12984,N_12881);
and U13102 (N_13102,N_12839,N_12785);
or U13103 (N_13103,N_12680,N_12769);
or U13104 (N_13104,N_12954,N_12821);
and U13105 (N_13105,N_12712,N_12564);
xor U13106 (N_13106,N_12813,N_12963);
nand U13107 (N_13107,N_12598,N_12780);
xnor U13108 (N_13108,N_12961,N_12648);
or U13109 (N_13109,N_12665,N_12876);
xor U13110 (N_13110,N_12828,N_12578);
nand U13111 (N_13111,N_12710,N_12742);
nand U13112 (N_13112,N_12903,N_12869);
and U13113 (N_13113,N_12618,N_12554);
nor U13114 (N_13114,N_12657,N_12699);
xnor U13115 (N_13115,N_12525,N_12924);
or U13116 (N_13116,N_12611,N_12643);
nor U13117 (N_13117,N_12656,N_12609);
nand U13118 (N_13118,N_12817,N_12860);
nor U13119 (N_13119,N_12688,N_12812);
xnor U13120 (N_13120,N_12760,N_12585);
and U13121 (N_13121,N_12527,N_12567);
and U13122 (N_13122,N_12518,N_12936);
nor U13123 (N_13123,N_12774,N_12967);
xor U13124 (N_13124,N_12719,N_12878);
nand U13125 (N_13125,N_12966,N_12996);
or U13126 (N_13126,N_12977,N_12833);
xor U13127 (N_13127,N_12631,N_12949);
or U13128 (N_13128,N_12899,N_12721);
nor U13129 (N_13129,N_12691,N_12737);
nand U13130 (N_13130,N_12690,N_12758);
xnor U13131 (N_13131,N_12811,N_12586);
nand U13132 (N_13132,N_12927,N_12674);
xnor U13133 (N_13133,N_12889,N_12504);
xnor U13134 (N_13134,N_12521,N_12610);
nand U13135 (N_13135,N_12922,N_12736);
xnor U13136 (N_13136,N_12709,N_12835);
or U13137 (N_13137,N_12717,N_12793);
nand U13138 (N_13138,N_12971,N_12523);
nor U13139 (N_13139,N_12573,N_12542);
and U13140 (N_13140,N_12779,N_12791);
or U13141 (N_13141,N_12836,N_12956);
and U13142 (N_13142,N_12988,N_12788);
and U13143 (N_13143,N_12856,N_12845);
or U13144 (N_13144,N_12945,N_12796);
nor U13145 (N_13145,N_12724,N_12725);
xnor U13146 (N_13146,N_12947,N_12617);
nor U13147 (N_13147,N_12787,N_12654);
and U13148 (N_13148,N_12551,N_12934);
and U13149 (N_13149,N_12550,N_12516);
and U13150 (N_13150,N_12533,N_12730);
nor U13151 (N_13151,N_12507,N_12647);
nor U13152 (N_13152,N_12849,N_12952);
or U13153 (N_13153,N_12764,N_12832);
nor U13154 (N_13154,N_12568,N_12810);
nor U13155 (N_13155,N_12595,N_12502);
and U13156 (N_13156,N_12744,N_12933);
and U13157 (N_13157,N_12570,N_12628);
nand U13158 (N_13158,N_12834,N_12935);
and U13159 (N_13159,N_12884,N_12773);
and U13160 (N_13160,N_12640,N_12944);
and U13161 (N_13161,N_12853,N_12757);
nand U13162 (N_13162,N_12660,N_12706);
nor U13163 (N_13163,N_12661,N_12501);
or U13164 (N_13164,N_12748,N_12775);
or U13165 (N_13165,N_12714,N_12978);
or U13166 (N_13166,N_12843,N_12590);
nand U13167 (N_13167,N_12768,N_12883);
nand U13168 (N_13168,N_12575,N_12767);
nor U13169 (N_13169,N_12515,N_12974);
and U13170 (N_13170,N_12816,N_12939);
nor U13171 (N_13171,N_12579,N_12621);
nor U13172 (N_13172,N_12716,N_12999);
and U13173 (N_13173,N_12509,N_12755);
or U13174 (N_13174,N_12951,N_12752);
nand U13175 (N_13175,N_12593,N_12771);
nand U13176 (N_13176,N_12908,N_12600);
nor U13177 (N_13177,N_12633,N_12781);
nand U13178 (N_13178,N_12930,N_12894);
and U13179 (N_13179,N_12655,N_12622);
nand U13180 (N_13180,N_12644,N_12919);
or U13181 (N_13181,N_12534,N_12630);
nand U13182 (N_13182,N_12663,N_12615);
or U13183 (N_13183,N_12953,N_12606);
nand U13184 (N_13184,N_12886,N_12571);
or U13185 (N_13185,N_12987,N_12741);
xnor U13186 (N_13186,N_12726,N_12754);
and U13187 (N_13187,N_12946,N_12682);
nand U13188 (N_13188,N_12720,N_12582);
and U13189 (N_13189,N_12918,N_12552);
xor U13190 (N_13190,N_12962,N_12937);
and U13191 (N_13191,N_12932,N_12973);
xnor U13192 (N_13192,N_12795,N_12668);
xnor U13193 (N_13193,N_12584,N_12914);
and U13194 (N_13194,N_12684,N_12650);
xnor U13195 (N_13195,N_12536,N_12970);
and U13196 (N_13196,N_12522,N_12838);
or U13197 (N_13197,N_12649,N_12808);
or U13198 (N_13198,N_12666,N_12964);
xnor U13199 (N_13199,N_12675,N_12563);
xor U13200 (N_13200,N_12823,N_12789);
nor U13201 (N_13201,N_12740,N_12904);
xnor U13202 (N_13202,N_12989,N_12825);
nor U13203 (N_13203,N_12653,N_12751);
or U13204 (N_13204,N_12805,N_12562);
nand U13205 (N_13205,N_12637,N_12519);
nand U13206 (N_13206,N_12896,N_12623);
xor U13207 (N_13207,N_12800,N_12851);
or U13208 (N_13208,N_12893,N_12926);
nor U13209 (N_13209,N_12613,N_12541);
nand U13210 (N_13210,N_12572,N_12957);
xnor U13211 (N_13211,N_12625,N_12687);
xnor U13212 (N_13212,N_12874,N_12959);
xnor U13213 (N_13213,N_12731,N_12747);
or U13214 (N_13214,N_12929,N_12818);
nand U13215 (N_13215,N_12505,N_12797);
nand U13216 (N_13216,N_12882,N_12671);
and U13217 (N_13217,N_12923,N_12646);
xor U13218 (N_13218,N_12645,N_12581);
nand U13219 (N_13219,N_12913,N_12993);
xnor U13220 (N_13220,N_12983,N_12732);
nand U13221 (N_13221,N_12943,N_12837);
and U13222 (N_13222,N_12981,N_12921);
and U13223 (N_13223,N_12992,N_12553);
xor U13224 (N_13224,N_12870,N_12594);
xor U13225 (N_13225,N_12559,N_12830);
nand U13226 (N_13226,N_12890,N_12759);
and U13227 (N_13227,N_12528,N_12511);
nor U13228 (N_13228,N_12591,N_12681);
nor U13229 (N_13229,N_12905,N_12831);
or U13230 (N_13230,N_12635,N_12848);
nor U13231 (N_13231,N_12840,N_12612);
xnor U13232 (N_13232,N_12746,N_12803);
nand U13233 (N_13233,N_12770,N_12857);
or U13234 (N_13234,N_12887,N_12960);
or U13235 (N_13235,N_12508,N_12669);
nor U13236 (N_13236,N_12608,N_12995);
or U13237 (N_13237,N_12975,N_12512);
and U13238 (N_13238,N_12872,N_12862);
nand U13239 (N_13239,N_12707,N_12955);
xnor U13240 (N_13240,N_12873,N_12814);
and U13241 (N_13241,N_12718,N_12627);
and U13242 (N_13242,N_12948,N_12544);
xor U13243 (N_13243,N_12891,N_12583);
or U13244 (N_13244,N_12634,N_12557);
xor U13245 (N_13245,N_12733,N_12931);
nor U13246 (N_13246,N_12799,N_12900);
xnor U13247 (N_13247,N_12616,N_12540);
xnor U13248 (N_13248,N_12500,N_12938);
nand U13249 (N_13249,N_12566,N_12597);
and U13250 (N_13250,N_12580,N_12523);
nand U13251 (N_13251,N_12975,N_12945);
or U13252 (N_13252,N_12880,N_12862);
and U13253 (N_13253,N_12895,N_12734);
nor U13254 (N_13254,N_12731,N_12702);
or U13255 (N_13255,N_12979,N_12998);
or U13256 (N_13256,N_12578,N_12972);
and U13257 (N_13257,N_12559,N_12827);
nand U13258 (N_13258,N_12763,N_12670);
or U13259 (N_13259,N_12776,N_12645);
and U13260 (N_13260,N_12519,N_12761);
nand U13261 (N_13261,N_12734,N_12785);
and U13262 (N_13262,N_12568,N_12750);
nor U13263 (N_13263,N_12654,N_12613);
or U13264 (N_13264,N_12665,N_12659);
or U13265 (N_13265,N_12999,N_12802);
xnor U13266 (N_13266,N_12637,N_12529);
or U13267 (N_13267,N_12504,N_12510);
or U13268 (N_13268,N_12508,N_12739);
nand U13269 (N_13269,N_12948,N_12850);
or U13270 (N_13270,N_12515,N_12897);
xor U13271 (N_13271,N_12742,N_12637);
nand U13272 (N_13272,N_12864,N_12872);
or U13273 (N_13273,N_12707,N_12728);
nand U13274 (N_13274,N_12587,N_12894);
or U13275 (N_13275,N_12940,N_12532);
xnor U13276 (N_13276,N_12645,N_12659);
xor U13277 (N_13277,N_12826,N_12764);
nor U13278 (N_13278,N_12769,N_12971);
or U13279 (N_13279,N_12699,N_12763);
nor U13280 (N_13280,N_12981,N_12555);
nor U13281 (N_13281,N_12848,N_12512);
nand U13282 (N_13282,N_12967,N_12521);
xor U13283 (N_13283,N_12831,N_12751);
xnor U13284 (N_13284,N_12973,N_12944);
or U13285 (N_13285,N_12665,N_12897);
nor U13286 (N_13286,N_12723,N_12537);
xor U13287 (N_13287,N_12861,N_12936);
nand U13288 (N_13288,N_12689,N_12846);
nor U13289 (N_13289,N_12917,N_12609);
and U13290 (N_13290,N_12759,N_12962);
nor U13291 (N_13291,N_12938,N_12809);
and U13292 (N_13292,N_12980,N_12894);
or U13293 (N_13293,N_12987,N_12753);
xor U13294 (N_13294,N_12684,N_12654);
or U13295 (N_13295,N_12990,N_12721);
nor U13296 (N_13296,N_12563,N_12755);
or U13297 (N_13297,N_12621,N_12975);
xor U13298 (N_13298,N_12690,N_12863);
xnor U13299 (N_13299,N_12683,N_12754);
and U13300 (N_13300,N_12599,N_12951);
nand U13301 (N_13301,N_12747,N_12901);
xor U13302 (N_13302,N_12719,N_12888);
and U13303 (N_13303,N_12847,N_12940);
nand U13304 (N_13304,N_12703,N_12930);
nand U13305 (N_13305,N_12519,N_12638);
nand U13306 (N_13306,N_12645,N_12601);
nor U13307 (N_13307,N_12684,N_12930);
xnor U13308 (N_13308,N_12704,N_12808);
and U13309 (N_13309,N_12521,N_12724);
and U13310 (N_13310,N_12696,N_12743);
and U13311 (N_13311,N_12934,N_12917);
xnor U13312 (N_13312,N_12796,N_12604);
nor U13313 (N_13313,N_12616,N_12740);
and U13314 (N_13314,N_12819,N_12769);
or U13315 (N_13315,N_12843,N_12762);
nor U13316 (N_13316,N_12527,N_12781);
xnor U13317 (N_13317,N_12613,N_12888);
nand U13318 (N_13318,N_12626,N_12668);
nor U13319 (N_13319,N_12730,N_12616);
or U13320 (N_13320,N_12719,N_12749);
and U13321 (N_13321,N_12924,N_12845);
nor U13322 (N_13322,N_12576,N_12536);
nand U13323 (N_13323,N_12887,N_12746);
and U13324 (N_13324,N_12961,N_12528);
nand U13325 (N_13325,N_12520,N_12849);
xor U13326 (N_13326,N_12517,N_12636);
xnor U13327 (N_13327,N_12632,N_12612);
or U13328 (N_13328,N_12871,N_12885);
nand U13329 (N_13329,N_12813,N_12920);
or U13330 (N_13330,N_12608,N_12635);
nand U13331 (N_13331,N_12519,N_12801);
xor U13332 (N_13332,N_12826,N_12732);
nor U13333 (N_13333,N_12851,N_12569);
nor U13334 (N_13334,N_12732,N_12579);
or U13335 (N_13335,N_12932,N_12592);
nor U13336 (N_13336,N_12502,N_12820);
or U13337 (N_13337,N_12879,N_12730);
and U13338 (N_13338,N_12838,N_12599);
and U13339 (N_13339,N_12787,N_12572);
or U13340 (N_13340,N_12820,N_12883);
nand U13341 (N_13341,N_12925,N_12508);
nor U13342 (N_13342,N_12667,N_12608);
nand U13343 (N_13343,N_12866,N_12631);
and U13344 (N_13344,N_12702,N_12540);
nor U13345 (N_13345,N_12540,N_12614);
or U13346 (N_13346,N_12961,N_12589);
and U13347 (N_13347,N_12876,N_12529);
or U13348 (N_13348,N_12871,N_12962);
xor U13349 (N_13349,N_12716,N_12809);
nand U13350 (N_13350,N_12677,N_12737);
and U13351 (N_13351,N_12546,N_12761);
or U13352 (N_13352,N_12650,N_12940);
xnor U13353 (N_13353,N_12695,N_12518);
xor U13354 (N_13354,N_12910,N_12859);
or U13355 (N_13355,N_12879,N_12684);
or U13356 (N_13356,N_12597,N_12786);
nand U13357 (N_13357,N_12500,N_12944);
xor U13358 (N_13358,N_12883,N_12802);
and U13359 (N_13359,N_12853,N_12723);
xnor U13360 (N_13360,N_12700,N_12518);
nand U13361 (N_13361,N_12741,N_12722);
nor U13362 (N_13362,N_12550,N_12695);
xnor U13363 (N_13363,N_12697,N_12837);
nor U13364 (N_13364,N_12537,N_12747);
or U13365 (N_13365,N_12602,N_12949);
nor U13366 (N_13366,N_12920,N_12607);
and U13367 (N_13367,N_12586,N_12964);
xor U13368 (N_13368,N_12821,N_12969);
or U13369 (N_13369,N_12532,N_12856);
nand U13370 (N_13370,N_12572,N_12703);
nor U13371 (N_13371,N_12998,N_12657);
nor U13372 (N_13372,N_12658,N_12713);
xor U13373 (N_13373,N_12994,N_12619);
nand U13374 (N_13374,N_12960,N_12951);
and U13375 (N_13375,N_12732,N_12896);
or U13376 (N_13376,N_12925,N_12517);
nor U13377 (N_13377,N_12675,N_12811);
xor U13378 (N_13378,N_12783,N_12755);
or U13379 (N_13379,N_12941,N_12615);
nor U13380 (N_13380,N_12905,N_12666);
nand U13381 (N_13381,N_12986,N_12634);
nand U13382 (N_13382,N_12707,N_12576);
nor U13383 (N_13383,N_12768,N_12727);
and U13384 (N_13384,N_12813,N_12562);
nand U13385 (N_13385,N_12526,N_12705);
and U13386 (N_13386,N_12795,N_12535);
and U13387 (N_13387,N_12835,N_12639);
nand U13388 (N_13388,N_12911,N_12754);
nand U13389 (N_13389,N_12965,N_12948);
nand U13390 (N_13390,N_12877,N_12737);
xnor U13391 (N_13391,N_12508,N_12778);
nor U13392 (N_13392,N_12801,N_12919);
nand U13393 (N_13393,N_12990,N_12803);
nor U13394 (N_13394,N_12811,N_12773);
and U13395 (N_13395,N_12993,N_12581);
or U13396 (N_13396,N_12654,N_12539);
xor U13397 (N_13397,N_12979,N_12746);
or U13398 (N_13398,N_12648,N_12914);
xor U13399 (N_13399,N_12891,N_12879);
nand U13400 (N_13400,N_12708,N_12629);
or U13401 (N_13401,N_12962,N_12672);
nand U13402 (N_13402,N_12685,N_12825);
and U13403 (N_13403,N_12740,N_12982);
and U13404 (N_13404,N_12960,N_12617);
xnor U13405 (N_13405,N_12861,N_12582);
or U13406 (N_13406,N_12828,N_12800);
nor U13407 (N_13407,N_12937,N_12849);
xnor U13408 (N_13408,N_12597,N_12757);
nand U13409 (N_13409,N_12731,N_12941);
nand U13410 (N_13410,N_12665,N_12627);
nor U13411 (N_13411,N_12941,N_12781);
xnor U13412 (N_13412,N_12986,N_12922);
and U13413 (N_13413,N_12934,N_12762);
nor U13414 (N_13414,N_12710,N_12640);
xor U13415 (N_13415,N_12797,N_12724);
and U13416 (N_13416,N_12836,N_12829);
nand U13417 (N_13417,N_12899,N_12733);
xnor U13418 (N_13418,N_12616,N_12824);
or U13419 (N_13419,N_12812,N_12795);
xor U13420 (N_13420,N_12519,N_12508);
and U13421 (N_13421,N_12608,N_12682);
and U13422 (N_13422,N_12730,N_12963);
or U13423 (N_13423,N_12702,N_12854);
nand U13424 (N_13424,N_12569,N_12560);
or U13425 (N_13425,N_12526,N_12893);
xor U13426 (N_13426,N_12822,N_12639);
or U13427 (N_13427,N_12717,N_12700);
or U13428 (N_13428,N_12500,N_12939);
or U13429 (N_13429,N_12515,N_12721);
and U13430 (N_13430,N_12876,N_12664);
and U13431 (N_13431,N_12662,N_12744);
nand U13432 (N_13432,N_12702,N_12572);
and U13433 (N_13433,N_12813,N_12958);
and U13434 (N_13434,N_12619,N_12502);
or U13435 (N_13435,N_12657,N_12975);
nor U13436 (N_13436,N_12785,N_12841);
nand U13437 (N_13437,N_12629,N_12886);
or U13438 (N_13438,N_12599,N_12513);
and U13439 (N_13439,N_12523,N_12500);
nand U13440 (N_13440,N_12917,N_12671);
nand U13441 (N_13441,N_12832,N_12803);
and U13442 (N_13442,N_12771,N_12944);
nor U13443 (N_13443,N_12925,N_12759);
xor U13444 (N_13444,N_12676,N_12947);
nand U13445 (N_13445,N_12960,N_12690);
xnor U13446 (N_13446,N_12671,N_12717);
and U13447 (N_13447,N_12643,N_12645);
xor U13448 (N_13448,N_12644,N_12973);
and U13449 (N_13449,N_12525,N_12588);
xor U13450 (N_13450,N_12517,N_12936);
and U13451 (N_13451,N_12916,N_12969);
xor U13452 (N_13452,N_12848,N_12665);
nor U13453 (N_13453,N_12771,N_12617);
xor U13454 (N_13454,N_12771,N_12551);
or U13455 (N_13455,N_12702,N_12942);
or U13456 (N_13456,N_12553,N_12780);
xnor U13457 (N_13457,N_12857,N_12586);
or U13458 (N_13458,N_12906,N_12555);
nor U13459 (N_13459,N_12639,N_12604);
and U13460 (N_13460,N_12555,N_12741);
xnor U13461 (N_13461,N_12955,N_12692);
nor U13462 (N_13462,N_12617,N_12660);
or U13463 (N_13463,N_12598,N_12600);
xnor U13464 (N_13464,N_12873,N_12971);
nand U13465 (N_13465,N_12563,N_12676);
xnor U13466 (N_13466,N_12693,N_12640);
xnor U13467 (N_13467,N_12541,N_12788);
nor U13468 (N_13468,N_12543,N_12819);
xnor U13469 (N_13469,N_12990,N_12877);
and U13470 (N_13470,N_12595,N_12602);
xor U13471 (N_13471,N_12575,N_12758);
nor U13472 (N_13472,N_12592,N_12666);
nand U13473 (N_13473,N_12896,N_12739);
and U13474 (N_13474,N_12841,N_12584);
nor U13475 (N_13475,N_12911,N_12730);
and U13476 (N_13476,N_12839,N_12813);
or U13477 (N_13477,N_12830,N_12936);
nor U13478 (N_13478,N_12914,N_12735);
xnor U13479 (N_13479,N_12563,N_12969);
or U13480 (N_13480,N_12718,N_12898);
or U13481 (N_13481,N_12519,N_12997);
and U13482 (N_13482,N_12897,N_12743);
or U13483 (N_13483,N_12751,N_12877);
and U13484 (N_13484,N_12853,N_12948);
xnor U13485 (N_13485,N_12855,N_12541);
nand U13486 (N_13486,N_12941,N_12646);
nand U13487 (N_13487,N_12600,N_12617);
and U13488 (N_13488,N_12674,N_12997);
xor U13489 (N_13489,N_12809,N_12551);
or U13490 (N_13490,N_12719,N_12532);
nand U13491 (N_13491,N_12502,N_12693);
and U13492 (N_13492,N_12543,N_12968);
or U13493 (N_13493,N_12548,N_12654);
nand U13494 (N_13494,N_12962,N_12752);
xnor U13495 (N_13495,N_12987,N_12701);
nor U13496 (N_13496,N_12806,N_12914);
or U13497 (N_13497,N_12727,N_12813);
or U13498 (N_13498,N_12769,N_12948);
xnor U13499 (N_13499,N_12810,N_12734);
nand U13500 (N_13500,N_13202,N_13480);
or U13501 (N_13501,N_13274,N_13302);
or U13502 (N_13502,N_13270,N_13330);
and U13503 (N_13503,N_13460,N_13285);
or U13504 (N_13504,N_13450,N_13421);
xnor U13505 (N_13505,N_13346,N_13391);
nor U13506 (N_13506,N_13322,N_13030);
xor U13507 (N_13507,N_13019,N_13101);
xor U13508 (N_13508,N_13200,N_13357);
and U13509 (N_13509,N_13241,N_13212);
xnor U13510 (N_13510,N_13208,N_13482);
nand U13511 (N_13511,N_13224,N_13052);
xnor U13512 (N_13512,N_13328,N_13429);
and U13513 (N_13513,N_13141,N_13121);
or U13514 (N_13514,N_13010,N_13182);
nor U13515 (N_13515,N_13418,N_13281);
xnor U13516 (N_13516,N_13031,N_13159);
nand U13517 (N_13517,N_13237,N_13265);
nor U13518 (N_13518,N_13117,N_13493);
nor U13519 (N_13519,N_13289,N_13446);
or U13520 (N_13520,N_13057,N_13492);
nor U13521 (N_13521,N_13283,N_13111);
nand U13522 (N_13522,N_13044,N_13228);
xnor U13523 (N_13523,N_13275,N_13110);
or U13524 (N_13524,N_13015,N_13012);
xnor U13525 (N_13525,N_13254,N_13222);
nor U13526 (N_13526,N_13350,N_13298);
nand U13527 (N_13527,N_13297,N_13428);
nor U13528 (N_13528,N_13478,N_13286);
and U13529 (N_13529,N_13223,N_13412);
xnor U13530 (N_13530,N_13175,N_13171);
and U13531 (N_13531,N_13261,N_13252);
nor U13532 (N_13532,N_13308,N_13307);
nand U13533 (N_13533,N_13143,N_13005);
and U13534 (N_13534,N_13156,N_13234);
nand U13535 (N_13535,N_13310,N_13292);
nand U13536 (N_13536,N_13444,N_13454);
nor U13537 (N_13537,N_13321,N_13045);
nand U13538 (N_13538,N_13487,N_13282);
xnor U13539 (N_13539,N_13469,N_13253);
or U13540 (N_13540,N_13128,N_13449);
nor U13541 (N_13541,N_13299,N_13495);
or U13542 (N_13542,N_13001,N_13414);
and U13543 (N_13543,N_13100,N_13189);
or U13544 (N_13544,N_13293,N_13024);
and U13545 (N_13545,N_13116,N_13055);
nand U13546 (N_13546,N_13186,N_13040);
or U13547 (N_13547,N_13406,N_13173);
xnor U13548 (N_13548,N_13023,N_13259);
nor U13549 (N_13549,N_13161,N_13301);
nand U13550 (N_13550,N_13191,N_13435);
nand U13551 (N_13551,N_13433,N_13476);
or U13552 (N_13552,N_13471,N_13071);
and U13553 (N_13553,N_13074,N_13432);
or U13554 (N_13554,N_13351,N_13017);
xor U13555 (N_13555,N_13213,N_13407);
xor U13556 (N_13556,N_13066,N_13436);
and U13557 (N_13557,N_13356,N_13473);
or U13558 (N_13558,N_13472,N_13287);
or U13559 (N_13559,N_13250,N_13375);
or U13560 (N_13560,N_13483,N_13073);
nor U13561 (N_13561,N_13392,N_13020);
nand U13562 (N_13562,N_13344,N_13205);
or U13563 (N_13563,N_13185,N_13154);
nand U13564 (N_13564,N_13046,N_13388);
xnor U13565 (N_13565,N_13104,N_13405);
xor U13566 (N_13566,N_13148,N_13437);
nor U13567 (N_13567,N_13164,N_13147);
xnor U13568 (N_13568,N_13341,N_13304);
xnor U13569 (N_13569,N_13135,N_13439);
or U13570 (N_13570,N_13124,N_13149);
and U13571 (N_13571,N_13174,N_13086);
or U13572 (N_13572,N_13268,N_13196);
and U13573 (N_13573,N_13059,N_13342);
xor U13574 (N_13574,N_13235,N_13009);
or U13575 (N_13575,N_13422,N_13312);
and U13576 (N_13576,N_13144,N_13003);
nand U13577 (N_13577,N_13221,N_13177);
and U13578 (N_13578,N_13078,N_13459);
xor U13579 (N_13579,N_13353,N_13236);
or U13580 (N_13580,N_13489,N_13188);
xnor U13581 (N_13581,N_13393,N_13376);
nor U13582 (N_13582,N_13199,N_13361);
and U13583 (N_13583,N_13324,N_13158);
nor U13584 (N_13584,N_13319,N_13070);
and U13585 (N_13585,N_13063,N_13399);
nor U13586 (N_13586,N_13430,N_13163);
nand U13587 (N_13587,N_13207,N_13458);
nor U13588 (N_13588,N_13413,N_13440);
and U13589 (N_13589,N_13220,N_13337);
xnor U13590 (N_13590,N_13457,N_13036);
and U13591 (N_13591,N_13008,N_13263);
or U13592 (N_13592,N_13484,N_13314);
or U13593 (N_13593,N_13166,N_13134);
or U13594 (N_13594,N_13033,N_13379);
or U13595 (N_13595,N_13425,N_13417);
or U13596 (N_13596,N_13214,N_13358);
nor U13597 (N_13597,N_13317,N_13119);
or U13598 (N_13598,N_13474,N_13363);
nor U13599 (N_13599,N_13348,N_13233);
nand U13600 (N_13600,N_13455,N_13318);
or U13601 (N_13601,N_13230,N_13088);
nor U13602 (N_13602,N_13076,N_13096);
nor U13603 (N_13603,N_13021,N_13043);
nand U13604 (N_13604,N_13258,N_13231);
nand U13605 (N_13605,N_13056,N_13061);
nand U13606 (N_13606,N_13386,N_13087);
xor U13607 (N_13607,N_13332,N_13131);
or U13608 (N_13608,N_13466,N_13416);
nor U13609 (N_13609,N_13278,N_13146);
nand U13610 (N_13610,N_13349,N_13380);
xor U13611 (N_13611,N_13452,N_13080);
xnor U13612 (N_13612,N_13145,N_13176);
nand U13613 (N_13613,N_13039,N_13113);
nor U13614 (N_13614,N_13465,N_13069);
nor U13615 (N_13615,N_13400,N_13083);
or U13616 (N_13616,N_13338,N_13058);
xor U13617 (N_13617,N_13419,N_13256);
or U13618 (N_13618,N_13443,N_13095);
or U13619 (N_13619,N_13127,N_13215);
or U13620 (N_13620,N_13226,N_13178);
and U13621 (N_13621,N_13306,N_13227);
nor U13622 (N_13622,N_13402,N_13309);
nor U13623 (N_13623,N_13099,N_13403);
xnor U13624 (N_13624,N_13384,N_13120);
and U13625 (N_13625,N_13211,N_13294);
nor U13626 (N_13626,N_13150,N_13497);
xnor U13627 (N_13627,N_13260,N_13387);
and U13628 (N_13628,N_13132,N_13242);
nand U13629 (N_13629,N_13053,N_13467);
xnor U13630 (N_13630,N_13248,N_13273);
nor U13631 (N_13631,N_13303,N_13198);
or U13632 (N_13632,N_13288,N_13415);
nand U13633 (N_13633,N_13206,N_13075);
xor U13634 (N_13634,N_13032,N_13142);
xnor U13635 (N_13635,N_13102,N_13038);
nor U13636 (N_13636,N_13169,N_13257);
and U13637 (N_13637,N_13369,N_13092);
and U13638 (N_13638,N_13225,N_13354);
and U13639 (N_13639,N_13067,N_13165);
xnor U13640 (N_13640,N_13204,N_13000);
or U13641 (N_13641,N_13448,N_13034);
and U13642 (N_13642,N_13323,N_13442);
nand U13643 (N_13643,N_13445,N_13180);
or U13644 (N_13644,N_13491,N_13456);
and U13645 (N_13645,N_13168,N_13496);
or U13646 (N_13646,N_13300,N_13488);
xnor U13647 (N_13647,N_13336,N_13105);
and U13648 (N_13648,N_13468,N_13389);
nand U13649 (N_13649,N_13160,N_13382);
xor U13650 (N_13650,N_13271,N_13002);
and U13651 (N_13651,N_13049,N_13272);
and U13652 (N_13652,N_13232,N_13155);
and U13653 (N_13653,N_13395,N_13434);
or U13654 (N_13654,N_13249,N_13329);
nand U13655 (N_13655,N_13431,N_13245);
xnor U13656 (N_13656,N_13172,N_13264);
xor U13657 (N_13657,N_13079,N_13360);
xor U13658 (N_13658,N_13453,N_13193);
and U13659 (N_13659,N_13410,N_13084);
xnor U13660 (N_13660,N_13219,N_13153);
nand U13661 (N_13661,N_13423,N_13451);
nand U13662 (N_13662,N_13006,N_13093);
and U13663 (N_13663,N_13162,N_13126);
and U13664 (N_13664,N_13401,N_13028);
or U13665 (N_13665,N_13404,N_13331);
and U13666 (N_13666,N_13463,N_13374);
or U13667 (N_13667,N_13359,N_13130);
and U13668 (N_13668,N_13136,N_13368);
nor U13669 (N_13669,N_13409,N_13209);
nor U13670 (N_13670,N_13438,N_13464);
and U13671 (N_13671,N_13364,N_13118);
xnor U13672 (N_13672,N_13262,N_13094);
or U13673 (N_13673,N_13152,N_13295);
nand U13674 (N_13674,N_13390,N_13305);
or U13675 (N_13675,N_13441,N_13279);
and U13676 (N_13676,N_13197,N_13378);
xor U13677 (N_13677,N_13026,N_13477);
and U13678 (N_13678,N_13335,N_13247);
or U13679 (N_13679,N_13426,N_13398);
xor U13680 (N_13680,N_13201,N_13485);
nor U13681 (N_13681,N_13139,N_13112);
nand U13682 (N_13682,N_13097,N_13427);
and U13683 (N_13683,N_13103,N_13107);
nand U13684 (N_13684,N_13123,N_13068);
or U13685 (N_13685,N_13133,N_13313);
xor U13686 (N_13686,N_13267,N_13396);
xor U13687 (N_13687,N_13089,N_13424);
and U13688 (N_13688,N_13187,N_13372);
or U13689 (N_13689,N_13284,N_13470);
nor U13690 (N_13690,N_13397,N_13371);
nand U13691 (N_13691,N_13064,N_13420);
nor U13692 (N_13692,N_13042,N_13311);
nand U13693 (N_13693,N_13138,N_13183);
nand U13694 (N_13694,N_13229,N_13109);
xor U13695 (N_13695,N_13238,N_13461);
xnor U13696 (N_13696,N_13246,N_13355);
and U13697 (N_13697,N_13479,N_13352);
xnor U13698 (N_13698,N_13106,N_13315);
nand U13699 (N_13699,N_13266,N_13326);
nor U13700 (N_13700,N_13025,N_13085);
and U13701 (N_13701,N_13081,N_13373);
and U13702 (N_13702,N_13016,N_13037);
and U13703 (N_13703,N_13217,N_13362);
nor U13704 (N_13704,N_13098,N_13377);
and U13705 (N_13705,N_13327,N_13255);
xor U13706 (N_13706,N_13027,N_13157);
nor U13707 (N_13707,N_13210,N_13269);
nor U13708 (N_13708,N_13022,N_13345);
xor U13709 (N_13709,N_13462,N_13447);
xor U13710 (N_13710,N_13486,N_13190);
xnor U13711 (N_13711,N_13218,N_13394);
and U13712 (N_13712,N_13498,N_13243);
xnor U13713 (N_13713,N_13475,N_13276);
or U13714 (N_13714,N_13339,N_13029);
xnor U13715 (N_13715,N_13333,N_13240);
nand U13716 (N_13716,N_13151,N_13125);
xor U13717 (N_13717,N_13320,N_13408);
nor U13718 (N_13718,N_13347,N_13291);
xor U13719 (N_13719,N_13490,N_13054);
nor U13720 (N_13720,N_13050,N_13411);
and U13721 (N_13721,N_13239,N_13343);
or U13722 (N_13722,N_13060,N_13122);
and U13723 (N_13723,N_13090,N_13137);
nor U13724 (N_13724,N_13325,N_13035);
nor U13725 (N_13725,N_13316,N_13129);
and U13726 (N_13726,N_13203,N_13011);
and U13727 (N_13727,N_13048,N_13366);
nand U13728 (N_13728,N_13072,N_13014);
nand U13729 (N_13729,N_13370,N_13184);
and U13730 (N_13730,N_13381,N_13082);
and U13731 (N_13731,N_13065,N_13091);
nand U13732 (N_13732,N_13077,N_13244);
nand U13733 (N_13733,N_13004,N_13340);
xor U13734 (N_13734,N_13296,N_13179);
nand U13735 (N_13735,N_13051,N_13167);
and U13736 (N_13736,N_13277,N_13385);
nand U13737 (N_13737,N_13194,N_13062);
or U13738 (N_13738,N_13290,N_13018);
nand U13739 (N_13739,N_13280,N_13181);
nor U13740 (N_13740,N_13365,N_13251);
or U13741 (N_13741,N_13013,N_13007);
nor U13742 (N_13742,N_13041,N_13383);
nand U13743 (N_13743,N_13140,N_13115);
nor U13744 (N_13744,N_13192,N_13114);
nor U13745 (N_13745,N_13499,N_13481);
or U13746 (N_13746,N_13216,N_13047);
or U13747 (N_13747,N_13334,N_13108);
xor U13748 (N_13748,N_13170,N_13195);
and U13749 (N_13749,N_13494,N_13367);
nand U13750 (N_13750,N_13067,N_13198);
or U13751 (N_13751,N_13265,N_13383);
nand U13752 (N_13752,N_13203,N_13451);
xor U13753 (N_13753,N_13138,N_13470);
or U13754 (N_13754,N_13398,N_13295);
and U13755 (N_13755,N_13007,N_13225);
and U13756 (N_13756,N_13024,N_13282);
nor U13757 (N_13757,N_13161,N_13230);
nand U13758 (N_13758,N_13243,N_13342);
and U13759 (N_13759,N_13307,N_13365);
xor U13760 (N_13760,N_13052,N_13264);
nand U13761 (N_13761,N_13035,N_13491);
nor U13762 (N_13762,N_13129,N_13445);
xor U13763 (N_13763,N_13312,N_13166);
or U13764 (N_13764,N_13404,N_13140);
nand U13765 (N_13765,N_13054,N_13415);
nand U13766 (N_13766,N_13249,N_13288);
xor U13767 (N_13767,N_13096,N_13142);
nor U13768 (N_13768,N_13146,N_13270);
nor U13769 (N_13769,N_13093,N_13425);
xor U13770 (N_13770,N_13193,N_13277);
or U13771 (N_13771,N_13130,N_13312);
nand U13772 (N_13772,N_13085,N_13070);
or U13773 (N_13773,N_13484,N_13225);
and U13774 (N_13774,N_13302,N_13429);
xor U13775 (N_13775,N_13163,N_13484);
nand U13776 (N_13776,N_13371,N_13437);
or U13777 (N_13777,N_13243,N_13235);
xor U13778 (N_13778,N_13287,N_13257);
and U13779 (N_13779,N_13378,N_13236);
or U13780 (N_13780,N_13033,N_13353);
and U13781 (N_13781,N_13397,N_13292);
nor U13782 (N_13782,N_13127,N_13294);
and U13783 (N_13783,N_13457,N_13264);
nand U13784 (N_13784,N_13167,N_13470);
and U13785 (N_13785,N_13205,N_13068);
or U13786 (N_13786,N_13419,N_13326);
nand U13787 (N_13787,N_13394,N_13109);
or U13788 (N_13788,N_13075,N_13040);
or U13789 (N_13789,N_13204,N_13492);
or U13790 (N_13790,N_13330,N_13114);
xor U13791 (N_13791,N_13342,N_13179);
xnor U13792 (N_13792,N_13468,N_13079);
xor U13793 (N_13793,N_13429,N_13215);
or U13794 (N_13794,N_13226,N_13310);
and U13795 (N_13795,N_13268,N_13004);
nand U13796 (N_13796,N_13340,N_13245);
nor U13797 (N_13797,N_13481,N_13204);
and U13798 (N_13798,N_13366,N_13078);
nand U13799 (N_13799,N_13488,N_13229);
xnor U13800 (N_13800,N_13435,N_13365);
nand U13801 (N_13801,N_13128,N_13231);
nor U13802 (N_13802,N_13237,N_13080);
or U13803 (N_13803,N_13053,N_13446);
nand U13804 (N_13804,N_13389,N_13460);
and U13805 (N_13805,N_13154,N_13474);
nor U13806 (N_13806,N_13340,N_13218);
nand U13807 (N_13807,N_13290,N_13091);
nand U13808 (N_13808,N_13418,N_13023);
xnor U13809 (N_13809,N_13458,N_13389);
nor U13810 (N_13810,N_13311,N_13028);
nand U13811 (N_13811,N_13036,N_13054);
nand U13812 (N_13812,N_13357,N_13277);
and U13813 (N_13813,N_13247,N_13256);
or U13814 (N_13814,N_13494,N_13272);
nor U13815 (N_13815,N_13466,N_13348);
xor U13816 (N_13816,N_13234,N_13274);
or U13817 (N_13817,N_13216,N_13114);
or U13818 (N_13818,N_13189,N_13245);
nand U13819 (N_13819,N_13331,N_13364);
and U13820 (N_13820,N_13008,N_13404);
xnor U13821 (N_13821,N_13183,N_13295);
and U13822 (N_13822,N_13086,N_13444);
nand U13823 (N_13823,N_13184,N_13054);
nand U13824 (N_13824,N_13384,N_13018);
xor U13825 (N_13825,N_13056,N_13306);
nand U13826 (N_13826,N_13496,N_13341);
or U13827 (N_13827,N_13432,N_13282);
and U13828 (N_13828,N_13439,N_13282);
nand U13829 (N_13829,N_13089,N_13397);
nand U13830 (N_13830,N_13214,N_13242);
nand U13831 (N_13831,N_13361,N_13367);
and U13832 (N_13832,N_13407,N_13372);
xnor U13833 (N_13833,N_13308,N_13345);
nor U13834 (N_13834,N_13483,N_13299);
nand U13835 (N_13835,N_13209,N_13289);
or U13836 (N_13836,N_13114,N_13259);
nor U13837 (N_13837,N_13087,N_13399);
nand U13838 (N_13838,N_13416,N_13057);
nor U13839 (N_13839,N_13149,N_13390);
nor U13840 (N_13840,N_13172,N_13110);
nand U13841 (N_13841,N_13164,N_13467);
xor U13842 (N_13842,N_13285,N_13198);
xor U13843 (N_13843,N_13328,N_13207);
nor U13844 (N_13844,N_13367,N_13458);
nand U13845 (N_13845,N_13100,N_13049);
and U13846 (N_13846,N_13082,N_13211);
or U13847 (N_13847,N_13114,N_13292);
and U13848 (N_13848,N_13043,N_13165);
xor U13849 (N_13849,N_13071,N_13051);
and U13850 (N_13850,N_13185,N_13193);
and U13851 (N_13851,N_13203,N_13119);
xor U13852 (N_13852,N_13458,N_13285);
xnor U13853 (N_13853,N_13197,N_13231);
or U13854 (N_13854,N_13050,N_13140);
xnor U13855 (N_13855,N_13405,N_13079);
or U13856 (N_13856,N_13416,N_13282);
xnor U13857 (N_13857,N_13282,N_13392);
nand U13858 (N_13858,N_13338,N_13427);
or U13859 (N_13859,N_13063,N_13044);
nor U13860 (N_13860,N_13220,N_13474);
xor U13861 (N_13861,N_13361,N_13157);
nor U13862 (N_13862,N_13125,N_13011);
xor U13863 (N_13863,N_13065,N_13082);
xnor U13864 (N_13864,N_13100,N_13337);
and U13865 (N_13865,N_13245,N_13133);
and U13866 (N_13866,N_13270,N_13095);
and U13867 (N_13867,N_13402,N_13366);
and U13868 (N_13868,N_13168,N_13136);
and U13869 (N_13869,N_13392,N_13117);
nand U13870 (N_13870,N_13408,N_13413);
and U13871 (N_13871,N_13219,N_13204);
nand U13872 (N_13872,N_13127,N_13457);
nand U13873 (N_13873,N_13344,N_13182);
xnor U13874 (N_13874,N_13198,N_13075);
and U13875 (N_13875,N_13451,N_13239);
or U13876 (N_13876,N_13190,N_13116);
nor U13877 (N_13877,N_13017,N_13428);
xnor U13878 (N_13878,N_13472,N_13177);
or U13879 (N_13879,N_13044,N_13079);
xnor U13880 (N_13880,N_13445,N_13393);
xor U13881 (N_13881,N_13050,N_13348);
xnor U13882 (N_13882,N_13202,N_13101);
or U13883 (N_13883,N_13412,N_13007);
or U13884 (N_13884,N_13116,N_13196);
nor U13885 (N_13885,N_13117,N_13001);
xnor U13886 (N_13886,N_13231,N_13461);
xnor U13887 (N_13887,N_13207,N_13481);
xor U13888 (N_13888,N_13311,N_13344);
or U13889 (N_13889,N_13081,N_13340);
or U13890 (N_13890,N_13197,N_13465);
and U13891 (N_13891,N_13345,N_13178);
and U13892 (N_13892,N_13228,N_13000);
nand U13893 (N_13893,N_13344,N_13498);
nor U13894 (N_13894,N_13164,N_13136);
and U13895 (N_13895,N_13120,N_13351);
xor U13896 (N_13896,N_13281,N_13159);
or U13897 (N_13897,N_13035,N_13308);
xor U13898 (N_13898,N_13404,N_13004);
nor U13899 (N_13899,N_13047,N_13023);
and U13900 (N_13900,N_13013,N_13076);
or U13901 (N_13901,N_13045,N_13008);
nor U13902 (N_13902,N_13399,N_13202);
nand U13903 (N_13903,N_13102,N_13371);
nor U13904 (N_13904,N_13323,N_13435);
or U13905 (N_13905,N_13051,N_13016);
or U13906 (N_13906,N_13308,N_13335);
nand U13907 (N_13907,N_13198,N_13099);
and U13908 (N_13908,N_13280,N_13249);
xor U13909 (N_13909,N_13042,N_13025);
nand U13910 (N_13910,N_13173,N_13295);
xnor U13911 (N_13911,N_13167,N_13248);
xor U13912 (N_13912,N_13138,N_13323);
and U13913 (N_13913,N_13447,N_13016);
nand U13914 (N_13914,N_13341,N_13445);
nor U13915 (N_13915,N_13494,N_13434);
or U13916 (N_13916,N_13461,N_13170);
nor U13917 (N_13917,N_13096,N_13344);
nand U13918 (N_13918,N_13411,N_13065);
or U13919 (N_13919,N_13135,N_13145);
and U13920 (N_13920,N_13495,N_13157);
and U13921 (N_13921,N_13474,N_13303);
and U13922 (N_13922,N_13168,N_13137);
nand U13923 (N_13923,N_13286,N_13088);
and U13924 (N_13924,N_13236,N_13046);
or U13925 (N_13925,N_13357,N_13084);
nor U13926 (N_13926,N_13343,N_13366);
or U13927 (N_13927,N_13360,N_13298);
nand U13928 (N_13928,N_13482,N_13130);
nand U13929 (N_13929,N_13034,N_13287);
xor U13930 (N_13930,N_13446,N_13213);
nand U13931 (N_13931,N_13276,N_13158);
xnor U13932 (N_13932,N_13379,N_13293);
or U13933 (N_13933,N_13022,N_13264);
nor U13934 (N_13934,N_13498,N_13475);
nor U13935 (N_13935,N_13253,N_13318);
or U13936 (N_13936,N_13141,N_13115);
and U13937 (N_13937,N_13474,N_13494);
and U13938 (N_13938,N_13449,N_13016);
nor U13939 (N_13939,N_13180,N_13030);
xnor U13940 (N_13940,N_13260,N_13454);
nor U13941 (N_13941,N_13102,N_13246);
and U13942 (N_13942,N_13192,N_13023);
or U13943 (N_13943,N_13035,N_13009);
nor U13944 (N_13944,N_13214,N_13444);
xnor U13945 (N_13945,N_13402,N_13434);
xor U13946 (N_13946,N_13274,N_13460);
and U13947 (N_13947,N_13422,N_13100);
nor U13948 (N_13948,N_13366,N_13471);
nand U13949 (N_13949,N_13298,N_13081);
xor U13950 (N_13950,N_13237,N_13267);
xor U13951 (N_13951,N_13295,N_13279);
xor U13952 (N_13952,N_13209,N_13200);
nor U13953 (N_13953,N_13341,N_13024);
or U13954 (N_13954,N_13030,N_13224);
nor U13955 (N_13955,N_13022,N_13089);
xnor U13956 (N_13956,N_13394,N_13308);
nor U13957 (N_13957,N_13426,N_13153);
nor U13958 (N_13958,N_13187,N_13171);
or U13959 (N_13959,N_13028,N_13272);
nand U13960 (N_13960,N_13268,N_13236);
nor U13961 (N_13961,N_13028,N_13161);
or U13962 (N_13962,N_13056,N_13117);
nor U13963 (N_13963,N_13377,N_13178);
xor U13964 (N_13964,N_13275,N_13071);
xnor U13965 (N_13965,N_13174,N_13006);
or U13966 (N_13966,N_13071,N_13078);
or U13967 (N_13967,N_13048,N_13317);
xor U13968 (N_13968,N_13295,N_13145);
or U13969 (N_13969,N_13331,N_13197);
nor U13970 (N_13970,N_13496,N_13177);
or U13971 (N_13971,N_13210,N_13053);
and U13972 (N_13972,N_13479,N_13474);
nand U13973 (N_13973,N_13167,N_13185);
nand U13974 (N_13974,N_13481,N_13167);
and U13975 (N_13975,N_13199,N_13012);
and U13976 (N_13976,N_13476,N_13424);
xnor U13977 (N_13977,N_13010,N_13233);
nand U13978 (N_13978,N_13008,N_13362);
xnor U13979 (N_13979,N_13499,N_13148);
nor U13980 (N_13980,N_13127,N_13011);
nand U13981 (N_13981,N_13136,N_13120);
and U13982 (N_13982,N_13383,N_13423);
nand U13983 (N_13983,N_13052,N_13019);
and U13984 (N_13984,N_13380,N_13437);
or U13985 (N_13985,N_13189,N_13337);
nand U13986 (N_13986,N_13191,N_13453);
or U13987 (N_13987,N_13323,N_13167);
xnor U13988 (N_13988,N_13289,N_13410);
nor U13989 (N_13989,N_13168,N_13185);
xor U13990 (N_13990,N_13077,N_13296);
nor U13991 (N_13991,N_13497,N_13222);
nand U13992 (N_13992,N_13410,N_13340);
nand U13993 (N_13993,N_13368,N_13325);
and U13994 (N_13994,N_13426,N_13017);
nand U13995 (N_13995,N_13346,N_13381);
or U13996 (N_13996,N_13278,N_13263);
xnor U13997 (N_13997,N_13370,N_13122);
nor U13998 (N_13998,N_13157,N_13193);
xor U13999 (N_13999,N_13100,N_13349);
or U14000 (N_14000,N_13763,N_13884);
and U14001 (N_14001,N_13759,N_13794);
nand U14002 (N_14002,N_13738,N_13924);
nor U14003 (N_14003,N_13556,N_13880);
or U14004 (N_14004,N_13604,N_13964);
xnor U14005 (N_14005,N_13595,N_13955);
xor U14006 (N_14006,N_13576,N_13740);
and U14007 (N_14007,N_13878,N_13693);
xnor U14008 (N_14008,N_13666,N_13834);
or U14009 (N_14009,N_13939,N_13607);
nor U14010 (N_14010,N_13558,N_13781);
xor U14011 (N_14011,N_13718,N_13697);
and U14012 (N_14012,N_13546,N_13761);
nor U14013 (N_14013,N_13755,N_13678);
and U14014 (N_14014,N_13743,N_13862);
xor U14015 (N_14015,N_13831,N_13599);
or U14016 (N_14016,N_13935,N_13977);
xor U14017 (N_14017,N_13629,N_13904);
nor U14018 (N_14018,N_13901,N_13704);
nor U14019 (N_14019,N_13968,N_13571);
nand U14020 (N_14020,N_13797,N_13573);
nand U14021 (N_14021,N_13848,N_13766);
and U14022 (N_14022,N_13916,N_13757);
or U14023 (N_14023,N_13729,N_13575);
and U14024 (N_14024,N_13852,N_13992);
nand U14025 (N_14025,N_13510,N_13900);
nand U14026 (N_14026,N_13804,N_13512);
nand U14027 (N_14027,N_13849,N_13934);
nand U14028 (N_14028,N_13696,N_13787);
nor U14029 (N_14029,N_13502,N_13543);
and U14030 (N_14030,N_13758,N_13663);
nor U14031 (N_14031,N_13875,N_13997);
or U14032 (N_14032,N_13597,N_13555);
nand U14033 (N_14033,N_13756,N_13768);
and U14034 (N_14034,N_13530,N_13744);
nand U14035 (N_14035,N_13658,N_13933);
nand U14036 (N_14036,N_13717,N_13819);
or U14037 (N_14037,N_13507,N_13898);
nand U14038 (N_14038,N_13847,N_13855);
nor U14039 (N_14039,N_13568,N_13715);
nand U14040 (N_14040,N_13918,N_13810);
nor U14041 (N_14041,N_13679,N_13646);
and U14042 (N_14042,N_13559,N_13990);
nor U14043 (N_14043,N_13917,N_13726);
nor U14044 (N_14044,N_13713,N_13586);
xor U14045 (N_14045,N_13942,N_13619);
or U14046 (N_14046,N_13722,N_13865);
xor U14047 (N_14047,N_13680,N_13820);
nor U14048 (N_14048,N_13951,N_13504);
or U14049 (N_14049,N_13605,N_13813);
xor U14050 (N_14050,N_13998,N_13868);
nand U14051 (N_14051,N_13866,N_13554);
xnor U14052 (N_14052,N_13922,N_13822);
and U14053 (N_14053,N_13879,N_13683);
nor U14054 (N_14054,N_13513,N_13850);
nand U14055 (N_14055,N_13577,N_13579);
and U14056 (N_14056,N_13505,N_13843);
nor U14057 (N_14057,N_13653,N_13927);
and U14058 (N_14058,N_13881,N_13585);
nand U14059 (N_14059,N_13945,N_13527);
nand U14060 (N_14060,N_13692,N_13953);
nor U14061 (N_14061,N_13592,N_13617);
or U14062 (N_14062,N_13739,N_13937);
nor U14063 (N_14063,N_13814,N_13538);
or U14064 (N_14064,N_13603,N_13669);
nand U14065 (N_14065,N_13824,N_13973);
and U14066 (N_14066,N_13903,N_13811);
and U14067 (N_14067,N_13832,N_13562);
or U14068 (N_14068,N_13520,N_13701);
nor U14069 (N_14069,N_13869,N_13882);
nor U14070 (N_14070,N_13565,N_13549);
nor U14071 (N_14071,N_13695,N_13836);
nor U14072 (N_14072,N_13963,N_13703);
xor U14073 (N_14073,N_13642,N_13611);
xor U14074 (N_14074,N_13888,N_13932);
nand U14075 (N_14075,N_13788,N_13533);
xnor U14076 (N_14076,N_13796,N_13681);
nand U14077 (N_14077,N_13754,N_13566);
nor U14078 (N_14078,N_13838,N_13976);
and U14079 (N_14079,N_13574,N_13989);
xor U14080 (N_14080,N_13514,N_13615);
and U14081 (N_14081,N_13638,N_13550);
nor U14082 (N_14082,N_13521,N_13508);
nor U14083 (N_14083,N_13765,N_13730);
and U14084 (N_14084,N_13863,N_13890);
nand U14085 (N_14085,N_13802,N_13632);
or U14086 (N_14086,N_13539,N_13913);
or U14087 (N_14087,N_13800,N_13630);
nand U14088 (N_14088,N_13641,N_13639);
and U14089 (N_14089,N_13652,N_13987);
or U14090 (N_14090,N_13694,N_13517);
nand U14091 (N_14091,N_13594,N_13971);
and U14092 (N_14092,N_13570,N_13612);
nor U14093 (N_14093,N_13957,N_13979);
or U14094 (N_14094,N_13747,N_13691);
xor U14095 (N_14095,N_13816,N_13775);
nand U14096 (N_14096,N_13689,N_13910);
or U14097 (N_14097,N_13833,N_13857);
nand U14098 (N_14098,N_13503,N_13938);
xnor U14099 (N_14099,N_13867,N_13628);
or U14100 (N_14100,N_13567,N_13661);
or U14101 (N_14101,N_13561,N_13534);
nor U14102 (N_14102,N_13501,N_13516);
xnor U14103 (N_14103,N_13870,N_13515);
nand U14104 (N_14104,N_13557,N_13777);
xor U14105 (N_14105,N_13776,N_13805);
and U14106 (N_14106,N_13902,N_13706);
or U14107 (N_14107,N_13786,N_13807);
nor U14108 (N_14108,N_13943,N_13801);
nand U14109 (N_14109,N_13829,N_13986);
nor U14110 (N_14110,N_13705,N_13753);
nand U14111 (N_14111,N_13782,N_13853);
nand U14112 (N_14112,N_13798,N_13966);
or U14113 (N_14113,N_13529,N_13974);
and U14114 (N_14114,N_13608,N_13885);
xor U14115 (N_14115,N_13792,N_13899);
or U14116 (N_14116,N_13908,N_13789);
xnor U14117 (N_14117,N_13541,N_13780);
xnor U14118 (N_14118,N_13828,N_13660);
xor U14119 (N_14119,N_13746,N_13644);
xor U14120 (N_14120,N_13839,N_13941);
xor U14121 (N_14121,N_13818,N_13896);
or U14122 (N_14122,N_13877,N_13894);
xnor U14123 (N_14123,N_13978,N_13626);
nand U14124 (N_14124,N_13914,N_13544);
or U14125 (N_14125,N_13731,N_13621);
or U14126 (N_14126,N_13821,N_13817);
xor U14127 (N_14127,N_13873,N_13690);
or U14128 (N_14128,N_13688,N_13654);
and U14129 (N_14129,N_13581,N_13664);
nand U14130 (N_14130,N_13672,N_13522);
nand U14131 (N_14131,N_13795,N_13837);
xor U14132 (N_14132,N_13736,N_13871);
and U14133 (N_14133,N_13700,N_13634);
or U14134 (N_14134,N_13686,N_13657);
nand U14135 (N_14135,N_13648,N_13827);
nand U14136 (N_14136,N_13921,N_13600);
and U14137 (N_14137,N_13676,N_13809);
or U14138 (N_14138,N_13785,N_13699);
nand U14139 (N_14139,N_13685,N_13985);
xor U14140 (N_14140,N_13928,N_13716);
nand U14141 (N_14141,N_13708,N_13511);
xor U14142 (N_14142,N_13840,N_13564);
nand U14143 (N_14143,N_13636,N_13742);
nand U14144 (N_14144,N_13961,N_13655);
and U14145 (N_14145,N_13844,N_13674);
and U14146 (N_14146,N_13825,N_13732);
nor U14147 (N_14147,N_13545,N_13772);
nand U14148 (N_14148,N_13889,N_13734);
or U14149 (N_14149,N_13925,N_13682);
nand U14150 (N_14150,N_13996,N_13640);
nor U14151 (N_14151,N_13712,N_13948);
nor U14152 (N_14152,N_13624,N_13733);
xor U14153 (N_14153,N_13969,N_13861);
nand U14154 (N_14154,N_13946,N_13506);
xor U14155 (N_14155,N_13856,N_13725);
or U14156 (N_14156,N_13650,N_13892);
nand U14157 (N_14157,N_13752,N_13967);
and U14158 (N_14158,N_13525,N_13665);
nor U14159 (N_14159,N_13911,N_13893);
and U14160 (N_14160,N_13687,N_13891);
and U14161 (N_14161,N_13931,N_13774);
nand U14162 (N_14162,N_13618,N_13883);
xor U14163 (N_14163,N_13906,N_13930);
nor U14164 (N_14164,N_13872,N_13773);
and U14165 (N_14165,N_13659,N_13727);
nand U14166 (N_14166,N_13609,N_13764);
and U14167 (N_14167,N_13553,N_13656);
and U14168 (N_14168,N_13588,N_13684);
xnor U14169 (N_14169,N_13846,N_13926);
xnor U14170 (N_14170,N_13960,N_13649);
nor U14171 (N_14171,N_13728,N_13723);
nand U14172 (N_14172,N_13509,N_13735);
nand U14173 (N_14173,N_13601,N_13815);
nand U14174 (N_14174,N_13923,N_13623);
or U14175 (N_14175,N_13671,N_13959);
xnor U14176 (N_14176,N_13531,N_13950);
or U14177 (N_14177,N_13698,N_13859);
xnor U14178 (N_14178,N_13719,N_13526);
nor U14179 (N_14179,N_13988,N_13587);
nor U14180 (N_14180,N_13711,N_13769);
or U14181 (N_14181,N_13952,N_13637);
and U14182 (N_14182,N_13548,N_13647);
nand U14183 (N_14183,N_13572,N_13675);
and U14184 (N_14184,N_13949,N_13835);
nand U14185 (N_14185,N_13591,N_13826);
and U14186 (N_14186,N_13984,N_13536);
nor U14187 (N_14187,N_13860,N_13995);
or U14188 (N_14188,N_13830,N_13803);
nand U14189 (N_14189,N_13806,N_13677);
and U14190 (N_14190,N_13524,N_13583);
or U14191 (N_14191,N_13993,N_13741);
nand U14192 (N_14192,N_13750,N_13793);
nand U14193 (N_14193,N_13940,N_13907);
nand U14194 (N_14194,N_13542,N_13560);
and U14195 (N_14195,N_13702,N_13970);
xnor U14196 (N_14196,N_13622,N_13631);
nor U14197 (N_14197,N_13547,N_13905);
and U14198 (N_14198,N_13707,N_13762);
and U14199 (N_14199,N_13912,N_13842);
or U14200 (N_14200,N_13745,N_13994);
and U14201 (N_14201,N_13709,N_13929);
or U14202 (N_14202,N_13962,N_13598);
nor U14203 (N_14203,N_13633,N_13651);
or U14204 (N_14204,N_13851,N_13858);
and U14205 (N_14205,N_13721,N_13919);
and U14206 (N_14206,N_13783,N_13551);
nand U14207 (N_14207,N_13981,N_13580);
and U14208 (N_14208,N_13799,N_13737);
and U14209 (N_14209,N_13770,N_13610);
and U14210 (N_14210,N_13920,N_13552);
nand U14211 (N_14211,N_13645,N_13540);
nand U14212 (N_14212,N_13535,N_13519);
nor U14213 (N_14213,N_13895,N_13983);
and U14214 (N_14214,N_13841,N_13500);
nand U14215 (N_14215,N_13532,N_13613);
nand U14216 (N_14216,N_13668,N_13779);
and U14217 (N_14217,N_13748,N_13602);
nor U14218 (N_14218,N_13808,N_13673);
nand U14219 (N_14219,N_13710,N_13874);
nand U14220 (N_14220,N_13965,N_13537);
and U14221 (N_14221,N_13714,N_13643);
nor U14222 (N_14222,N_13915,N_13584);
and U14223 (N_14223,N_13760,N_13578);
nand U14224 (N_14224,N_13590,N_13947);
xor U14225 (N_14225,N_13845,N_13569);
or U14226 (N_14226,N_13956,N_13999);
and U14227 (N_14227,N_13635,N_13982);
nand U14228 (N_14228,N_13667,N_13662);
nor U14229 (N_14229,N_13593,N_13954);
nor U14230 (N_14230,N_13589,N_13864);
xor U14231 (N_14231,N_13991,N_13823);
nor U14232 (N_14232,N_13975,N_13909);
xor U14233 (N_14233,N_13791,N_13749);
nand U14234 (N_14234,N_13751,N_13876);
nor U14235 (N_14235,N_13784,N_13958);
and U14236 (N_14236,N_13980,N_13627);
or U14237 (N_14237,N_13670,N_13886);
or U14238 (N_14238,N_13582,N_13936);
nor U14239 (N_14239,N_13778,N_13563);
xnor U14240 (N_14240,N_13620,N_13812);
nor U14241 (N_14241,N_13518,N_13523);
nor U14242 (N_14242,N_13972,N_13854);
nor U14243 (N_14243,N_13625,N_13720);
nand U14244 (N_14244,N_13606,N_13944);
nor U14245 (N_14245,N_13724,N_13790);
nand U14246 (N_14246,N_13771,N_13616);
and U14247 (N_14247,N_13887,N_13528);
and U14248 (N_14248,N_13596,N_13767);
xnor U14249 (N_14249,N_13614,N_13897);
or U14250 (N_14250,N_13990,N_13868);
and U14251 (N_14251,N_13710,N_13609);
xor U14252 (N_14252,N_13694,N_13865);
and U14253 (N_14253,N_13785,N_13940);
and U14254 (N_14254,N_13505,N_13610);
xnor U14255 (N_14255,N_13635,N_13643);
nand U14256 (N_14256,N_13965,N_13840);
xnor U14257 (N_14257,N_13678,N_13567);
nor U14258 (N_14258,N_13666,N_13979);
xor U14259 (N_14259,N_13611,N_13571);
nand U14260 (N_14260,N_13741,N_13526);
nor U14261 (N_14261,N_13873,N_13895);
or U14262 (N_14262,N_13742,N_13897);
nand U14263 (N_14263,N_13920,N_13629);
nor U14264 (N_14264,N_13827,N_13739);
nor U14265 (N_14265,N_13866,N_13583);
nand U14266 (N_14266,N_13506,N_13736);
nand U14267 (N_14267,N_13566,N_13573);
xnor U14268 (N_14268,N_13994,N_13747);
nand U14269 (N_14269,N_13698,N_13597);
and U14270 (N_14270,N_13597,N_13718);
xnor U14271 (N_14271,N_13708,N_13564);
or U14272 (N_14272,N_13666,N_13827);
nor U14273 (N_14273,N_13547,N_13887);
xor U14274 (N_14274,N_13990,N_13717);
or U14275 (N_14275,N_13680,N_13920);
or U14276 (N_14276,N_13656,N_13510);
nor U14277 (N_14277,N_13684,N_13736);
nor U14278 (N_14278,N_13676,N_13930);
nor U14279 (N_14279,N_13502,N_13888);
nand U14280 (N_14280,N_13857,N_13691);
or U14281 (N_14281,N_13839,N_13784);
or U14282 (N_14282,N_13973,N_13710);
or U14283 (N_14283,N_13516,N_13719);
nand U14284 (N_14284,N_13595,N_13722);
xnor U14285 (N_14285,N_13781,N_13938);
nor U14286 (N_14286,N_13736,N_13781);
or U14287 (N_14287,N_13556,N_13976);
and U14288 (N_14288,N_13553,N_13978);
and U14289 (N_14289,N_13564,N_13504);
and U14290 (N_14290,N_13637,N_13533);
xor U14291 (N_14291,N_13885,N_13548);
or U14292 (N_14292,N_13980,N_13594);
and U14293 (N_14293,N_13838,N_13844);
nor U14294 (N_14294,N_13959,N_13749);
or U14295 (N_14295,N_13503,N_13645);
xor U14296 (N_14296,N_13957,N_13720);
and U14297 (N_14297,N_13547,N_13839);
nand U14298 (N_14298,N_13605,N_13517);
nand U14299 (N_14299,N_13998,N_13681);
nor U14300 (N_14300,N_13987,N_13953);
or U14301 (N_14301,N_13789,N_13666);
and U14302 (N_14302,N_13750,N_13922);
nor U14303 (N_14303,N_13602,N_13940);
nand U14304 (N_14304,N_13915,N_13967);
and U14305 (N_14305,N_13858,N_13643);
nor U14306 (N_14306,N_13951,N_13999);
or U14307 (N_14307,N_13711,N_13934);
nor U14308 (N_14308,N_13558,N_13958);
nor U14309 (N_14309,N_13523,N_13985);
nor U14310 (N_14310,N_13625,N_13782);
or U14311 (N_14311,N_13983,N_13909);
nand U14312 (N_14312,N_13761,N_13784);
nor U14313 (N_14313,N_13920,N_13937);
xor U14314 (N_14314,N_13725,N_13890);
nor U14315 (N_14315,N_13597,N_13508);
or U14316 (N_14316,N_13525,N_13858);
xor U14317 (N_14317,N_13914,N_13850);
nand U14318 (N_14318,N_13699,N_13914);
xor U14319 (N_14319,N_13982,N_13954);
or U14320 (N_14320,N_13509,N_13518);
xor U14321 (N_14321,N_13664,N_13642);
nand U14322 (N_14322,N_13889,N_13801);
nor U14323 (N_14323,N_13713,N_13964);
nor U14324 (N_14324,N_13690,N_13758);
and U14325 (N_14325,N_13807,N_13880);
nor U14326 (N_14326,N_13652,N_13785);
nand U14327 (N_14327,N_13655,N_13797);
or U14328 (N_14328,N_13831,N_13533);
or U14329 (N_14329,N_13619,N_13512);
xor U14330 (N_14330,N_13683,N_13924);
nand U14331 (N_14331,N_13641,N_13922);
and U14332 (N_14332,N_13645,N_13774);
nand U14333 (N_14333,N_13963,N_13990);
xor U14334 (N_14334,N_13855,N_13976);
nand U14335 (N_14335,N_13676,N_13907);
and U14336 (N_14336,N_13852,N_13646);
nand U14337 (N_14337,N_13545,N_13649);
xnor U14338 (N_14338,N_13873,N_13663);
and U14339 (N_14339,N_13927,N_13917);
or U14340 (N_14340,N_13859,N_13922);
xor U14341 (N_14341,N_13608,N_13612);
nand U14342 (N_14342,N_13656,N_13557);
nand U14343 (N_14343,N_13807,N_13924);
and U14344 (N_14344,N_13561,N_13888);
nor U14345 (N_14345,N_13823,N_13955);
or U14346 (N_14346,N_13984,N_13665);
or U14347 (N_14347,N_13795,N_13619);
and U14348 (N_14348,N_13500,N_13939);
or U14349 (N_14349,N_13588,N_13610);
xor U14350 (N_14350,N_13736,N_13747);
nand U14351 (N_14351,N_13763,N_13705);
and U14352 (N_14352,N_13957,N_13824);
or U14353 (N_14353,N_13822,N_13860);
and U14354 (N_14354,N_13530,N_13845);
nor U14355 (N_14355,N_13832,N_13790);
or U14356 (N_14356,N_13790,N_13915);
nand U14357 (N_14357,N_13940,N_13680);
nor U14358 (N_14358,N_13552,N_13910);
nand U14359 (N_14359,N_13742,N_13996);
nor U14360 (N_14360,N_13738,N_13833);
or U14361 (N_14361,N_13663,N_13555);
nand U14362 (N_14362,N_13886,N_13643);
or U14363 (N_14363,N_13745,N_13837);
nand U14364 (N_14364,N_13520,N_13542);
nand U14365 (N_14365,N_13639,N_13900);
nor U14366 (N_14366,N_13733,N_13773);
nor U14367 (N_14367,N_13504,N_13521);
xnor U14368 (N_14368,N_13609,N_13645);
nor U14369 (N_14369,N_13912,N_13629);
nor U14370 (N_14370,N_13736,N_13776);
nand U14371 (N_14371,N_13681,N_13857);
nor U14372 (N_14372,N_13685,N_13825);
xor U14373 (N_14373,N_13968,N_13771);
and U14374 (N_14374,N_13998,N_13743);
or U14375 (N_14375,N_13687,N_13801);
or U14376 (N_14376,N_13546,N_13717);
nand U14377 (N_14377,N_13907,N_13629);
or U14378 (N_14378,N_13946,N_13887);
nand U14379 (N_14379,N_13706,N_13675);
nand U14380 (N_14380,N_13782,N_13674);
nand U14381 (N_14381,N_13583,N_13994);
nor U14382 (N_14382,N_13663,N_13802);
xnor U14383 (N_14383,N_13855,N_13997);
nor U14384 (N_14384,N_13922,N_13996);
or U14385 (N_14385,N_13905,N_13595);
xnor U14386 (N_14386,N_13856,N_13716);
and U14387 (N_14387,N_13942,N_13559);
xnor U14388 (N_14388,N_13826,N_13945);
xnor U14389 (N_14389,N_13784,N_13729);
or U14390 (N_14390,N_13877,N_13971);
or U14391 (N_14391,N_13865,N_13977);
or U14392 (N_14392,N_13717,N_13621);
nor U14393 (N_14393,N_13635,N_13971);
and U14394 (N_14394,N_13979,N_13708);
nor U14395 (N_14395,N_13505,N_13501);
and U14396 (N_14396,N_13880,N_13668);
and U14397 (N_14397,N_13687,N_13802);
nor U14398 (N_14398,N_13812,N_13528);
or U14399 (N_14399,N_13562,N_13926);
nand U14400 (N_14400,N_13916,N_13576);
and U14401 (N_14401,N_13963,N_13663);
xor U14402 (N_14402,N_13910,N_13578);
xor U14403 (N_14403,N_13769,N_13872);
nor U14404 (N_14404,N_13679,N_13852);
and U14405 (N_14405,N_13677,N_13665);
and U14406 (N_14406,N_13785,N_13864);
or U14407 (N_14407,N_13781,N_13954);
nand U14408 (N_14408,N_13650,N_13973);
nor U14409 (N_14409,N_13724,N_13822);
nor U14410 (N_14410,N_13649,N_13987);
and U14411 (N_14411,N_13562,N_13979);
nand U14412 (N_14412,N_13683,N_13668);
xor U14413 (N_14413,N_13743,N_13529);
and U14414 (N_14414,N_13569,N_13626);
and U14415 (N_14415,N_13981,N_13675);
xnor U14416 (N_14416,N_13874,N_13696);
and U14417 (N_14417,N_13655,N_13865);
xor U14418 (N_14418,N_13762,N_13741);
or U14419 (N_14419,N_13641,N_13773);
or U14420 (N_14420,N_13838,N_13754);
and U14421 (N_14421,N_13761,N_13637);
and U14422 (N_14422,N_13604,N_13656);
nand U14423 (N_14423,N_13683,N_13985);
or U14424 (N_14424,N_13512,N_13625);
xnor U14425 (N_14425,N_13547,N_13514);
or U14426 (N_14426,N_13647,N_13588);
nor U14427 (N_14427,N_13725,N_13702);
xnor U14428 (N_14428,N_13826,N_13777);
nor U14429 (N_14429,N_13786,N_13803);
nor U14430 (N_14430,N_13522,N_13932);
and U14431 (N_14431,N_13905,N_13774);
nand U14432 (N_14432,N_13728,N_13627);
nor U14433 (N_14433,N_13649,N_13901);
nor U14434 (N_14434,N_13691,N_13670);
nand U14435 (N_14435,N_13661,N_13700);
or U14436 (N_14436,N_13849,N_13891);
xor U14437 (N_14437,N_13944,N_13774);
or U14438 (N_14438,N_13765,N_13582);
or U14439 (N_14439,N_13790,N_13919);
and U14440 (N_14440,N_13673,N_13878);
nor U14441 (N_14441,N_13923,N_13983);
nor U14442 (N_14442,N_13907,N_13543);
nand U14443 (N_14443,N_13698,N_13638);
xnor U14444 (N_14444,N_13681,N_13886);
xor U14445 (N_14445,N_13884,N_13518);
xnor U14446 (N_14446,N_13684,N_13623);
xnor U14447 (N_14447,N_13802,N_13537);
and U14448 (N_14448,N_13947,N_13791);
nor U14449 (N_14449,N_13961,N_13918);
xnor U14450 (N_14450,N_13722,N_13676);
or U14451 (N_14451,N_13682,N_13516);
nand U14452 (N_14452,N_13733,N_13576);
or U14453 (N_14453,N_13860,N_13890);
or U14454 (N_14454,N_13877,N_13525);
nand U14455 (N_14455,N_13536,N_13992);
or U14456 (N_14456,N_13718,N_13794);
or U14457 (N_14457,N_13878,N_13766);
and U14458 (N_14458,N_13709,N_13746);
and U14459 (N_14459,N_13510,N_13663);
or U14460 (N_14460,N_13815,N_13620);
xnor U14461 (N_14461,N_13597,N_13994);
or U14462 (N_14462,N_13688,N_13987);
and U14463 (N_14463,N_13726,N_13977);
nor U14464 (N_14464,N_13623,N_13711);
nand U14465 (N_14465,N_13826,N_13771);
nand U14466 (N_14466,N_13516,N_13693);
or U14467 (N_14467,N_13673,N_13908);
nor U14468 (N_14468,N_13545,N_13500);
xnor U14469 (N_14469,N_13676,N_13708);
nor U14470 (N_14470,N_13976,N_13503);
nand U14471 (N_14471,N_13669,N_13548);
nand U14472 (N_14472,N_13694,N_13657);
xnor U14473 (N_14473,N_13532,N_13991);
and U14474 (N_14474,N_13569,N_13791);
and U14475 (N_14475,N_13641,N_13505);
nor U14476 (N_14476,N_13673,N_13906);
nand U14477 (N_14477,N_13965,N_13766);
and U14478 (N_14478,N_13948,N_13526);
nor U14479 (N_14479,N_13700,N_13605);
nand U14480 (N_14480,N_13740,N_13725);
nand U14481 (N_14481,N_13928,N_13505);
nor U14482 (N_14482,N_13841,N_13956);
or U14483 (N_14483,N_13547,N_13549);
nor U14484 (N_14484,N_13608,N_13973);
or U14485 (N_14485,N_13588,N_13698);
and U14486 (N_14486,N_13859,N_13681);
nand U14487 (N_14487,N_13716,N_13746);
or U14488 (N_14488,N_13628,N_13956);
or U14489 (N_14489,N_13548,N_13625);
nor U14490 (N_14490,N_13676,N_13807);
nor U14491 (N_14491,N_13536,N_13600);
nor U14492 (N_14492,N_13611,N_13600);
xnor U14493 (N_14493,N_13650,N_13867);
nand U14494 (N_14494,N_13849,N_13834);
xor U14495 (N_14495,N_13658,N_13749);
and U14496 (N_14496,N_13819,N_13634);
nor U14497 (N_14497,N_13554,N_13651);
xor U14498 (N_14498,N_13535,N_13717);
nand U14499 (N_14499,N_13824,N_13975);
or U14500 (N_14500,N_14049,N_14431);
or U14501 (N_14501,N_14210,N_14305);
xor U14502 (N_14502,N_14393,N_14332);
and U14503 (N_14503,N_14430,N_14159);
or U14504 (N_14504,N_14373,N_14415);
and U14505 (N_14505,N_14356,N_14196);
or U14506 (N_14506,N_14339,N_14232);
nor U14507 (N_14507,N_14152,N_14486);
xnor U14508 (N_14508,N_14138,N_14452);
or U14509 (N_14509,N_14336,N_14046);
xnor U14510 (N_14510,N_14398,N_14437);
and U14511 (N_14511,N_14429,N_14456);
or U14512 (N_14512,N_14064,N_14307);
or U14513 (N_14513,N_14278,N_14166);
or U14514 (N_14514,N_14280,N_14033);
nand U14515 (N_14515,N_14099,N_14117);
or U14516 (N_14516,N_14198,N_14403);
nor U14517 (N_14517,N_14247,N_14438);
xor U14518 (N_14518,N_14017,N_14227);
or U14519 (N_14519,N_14281,N_14193);
and U14520 (N_14520,N_14459,N_14112);
and U14521 (N_14521,N_14069,N_14228);
nor U14522 (N_14522,N_14241,N_14182);
nand U14523 (N_14523,N_14239,N_14480);
or U14524 (N_14524,N_14086,N_14105);
nand U14525 (N_14525,N_14122,N_14255);
nand U14526 (N_14526,N_14291,N_14355);
and U14527 (N_14527,N_14286,N_14318);
xnor U14528 (N_14528,N_14412,N_14026);
nand U14529 (N_14529,N_14482,N_14229);
and U14530 (N_14530,N_14365,N_14254);
or U14531 (N_14531,N_14016,N_14218);
nor U14532 (N_14532,N_14208,N_14400);
nand U14533 (N_14533,N_14436,N_14110);
or U14534 (N_14534,N_14370,N_14235);
nor U14535 (N_14535,N_14475,N_14071);
xor U14536 (N_14536,N_14157,N_14382);
or U14537 (N_14537,N_14334,N_14207);
nor U14538 (N_14538,N_14472,N_14055);
nand U14539 (N_14539,N_14192,N_14076);
nor U14540 (N_14540,N_14427,N_14406);
and U14541 (N_14541,N_14184,N_14283);
or U14542 (N_14542,N_14432,N_14168);
xor U14543 (N_14543,N_14333,N_14005);
xor U14544 (N_14544,N_14113,N_14097);
or U14545 (N_14545,N_14092,N_14484);
xnor U14546 (N_14546,N_14290,N_14455);
xor U14547 (N_14547,N_14317,N_14156);
nor U14548 (N_14548,N_14111,N_14006);
nor U14549 (N_14549,N_14267,N_14119);
xnor U14550 (N_14550,N_14380,N_14357);
and U14551 (N_14551,N_14024,N_14129);
xnor U14552 (N_14552,N_14203,N_14428);
xor U14553 (N_14553,N_14478,N_14185);
nand U14554 (N_14554,N_14367,N_14223);
xnor U14555 (N_14555,N_14359,N_14375);
or U14556 (N_14556,N_14053,N_14433);
xnor U14557 (N_14557,N_14108,N_14195);
and U14558 (N_14558,N_14376,N_14288);
nand U14559 (N_14559,N_14411,N_14036);
nand U14560 (N_14560,N_14217,N_14287);
nand U14561 (N_14561,N_14153,N_14421);
xnor U14562 (N_14562,N_14042,N_14128);
or U14563 (N_14563,N_14021,N_14065);
and U14564 (N_14564,N_14491,N_14029);
xnor U14565 (N_14565,N_14466,N_14186);
and U14566 (N_14566,N_14141,N_14023);
xnor U14567 (N_14567,N_14404,N_14424);
nor U14568 (N_14568,N_14230,N_14088);
xor U14569 (N_14569,N_14018,N_14199);
and U14570 (N_14570,N_14409,N_14037);
nand U14571 (N_14571,N_14212,N_14276);
or U14572 (N_14572,N_14084,N_14324);
and U14573 (N_14573,N_14214,N_14014);
or U14574 (N_14574,N_14030,N_14008);
nor U14575 (N_14575,N_14385,N_14078);
or U14576 (N_14576,N_14183,N_14109);
xor U14577 (N_14577,N_14360,N_14272);
or U14578 (N_14578,N_14449,N_14352);
or U14579 (N_14579,N_14137,N_14450);
xnor U14580 (N_14580,N_14273,N_14487);
xor U14581 (N_14581,N_14350,N_14143);
nor U14582 (N_14582,N_14261,N_14224);
nor U14583 (N_14583,N_14003,N_14170);
nor U14584 (N_14584,N_14298,N_14209);
nor U14585 (N_14585,N_14384,N_14263);
and U14586 (N_14586,N_14440,N_14469);
nand U14587 (N_14587,N_14392,N_14050);
and U14588 (N_14588,N_14419,N_14041);
and U14589 (N_14589,N_14454,N_14399);
nor U14590 (N_14590,N_14066,N_14204);
and U14591 (N_14591,N_14171,N_14163);
nor U14592 (N_14592,N_14426,N_14351);
or U14593 (N_14593,N_14463,N_14158);
nor U14594 (N_14594,N_14022,N_14057);
or U14595 (N_14595,N_14091,N_14100);
nand U14596 (N_14596,N_14221,N_14354);
nand U14597 (N_14597,N_14031,N_14443);
xor U14598 (N_14598,N_14107,N_14330);
or U14599 (N_14599,N_14397,N_14251);
or U14600 (N_14600,N_14101,N_14079);
nor U14601 (N_14601,N_14222,N_14175);
nor U14602 (N_14602,N_14087,N_14338);
nand U14603 (N_14603,N_14059,N_14446);
nand U14604 (N_14604,N_14151,N_14048);
and U14605 (N_14605,N_14481,N_14114);
or U14606 (N_14606,N_14106,N_14477);
nand U14607 (N_14607,N_14180,N_14306);
xnor U14608 (N_14608,N_14345,N_14483);
and U14609 (N_14609,N_14173,N_14445);
or U14610 (N_14610,N_14314,N_14083);
or U14611 (N_14611,N_14162,N_14028);
nor U14612 (N_14612,N_14134,N_14001);
or U14613 (N_14613,N_14147,N_14448);
xnor U14614 (N_14614,N_14249,N_14269);
xnor U14615 (N_14615,N_14342,N_14172);
and U14616 (N_14616,N_14169,N_14407);
and U14617 (N_14617,N_14377,N_14139);
nor U14618 (N_14618,N_14231,N_14270);
or U14619 (N_14619,N_14019,N_14479);
xnor U14620 (N_14620,N_14335,N_14374);
or U14621 (N_14621,N_14002,N_14225);
nand U14622 (N_14622,N_14346,N_14371);
nor U14623 (N_14623,N_14341,N_14009);
and U14624 (N_14624,N_14067,N_14040);
and U14625 (N_14625,N_14045,N_14118);
or U14626 (N_14626,N_14361,N_14080);
or U14627 (N_14627,N_14468,N_14379);
and U14628 (N_14628,N_14020,N_14073);
nand U14629 (N_14629,N_14155,N_14289);
xor U14630 (N_14630,N_14090,N_14476);
nand U14631 (N_14631,N_14387,N_14242);
xor U14632 (N_14632,N_14148,N_14420);
and U14633 (N_14633,N_14369,N_14416);
or U14634 (N_14634,N_14275,N_14328);
nand U14635 (N_14635,N_14326,N_14439);
nor U14636 (N_14636,N_14451,N_14081);
or U14637 (N_14637,N_14343,N_14226);
or U14638 (N_14638,N_14102,N_14259);
and U14639 (N_14639,N_14015,N_14285);
nand U14640 (N_14640,N_14442,N_14142);
and U14641 (N_14641,N_14165,N_14130);
nand U14642 (N_14642,N_14401,N_14258);
nor U14643 (N_14643,N_14039,N_14423);
and U14644 (N_14644,N_14124,N_14197);
or U14645 (N_14645,N_14274,N_14123);
xnor U14646 (N_14646,N_14062,N_14095);
and U14647 (N_14647,N_14394,N_14304);
xor U14648 (N_14648,N_14444,N_14136);
or U14649 (N_14649,N_14312,N_14489);
and U14650 (N_14650,N_14160,N_14434);
and U14651 (N_14651,N_14191,N_14211);
nand U14652 (N_14652,N_14457,N_14070);
and U14653 (N_14653,N_14331,N_14068);
and U14654 (N_14654,N_14093,N_14043);
xor U14655 (N_14655,N_14051,N_14120);
or U14656 (N_14656,N_14297,N_14414);
nand U14657 (N_14657,N_14292,N_14441);
nor U14658 (N_14658,N_14311,N_14140);
or U14659 (N_14659,N_14310,N_14188);
or U14660 (N_14660,N_14320,N_14150);
or U14661 (N_14661,N_14115,N_14381);
nor U14662 (N_14662,N_14245,N_14422);
xor U14663 (N_14663,N_14104,N_14490);
xor U14664 (N_14664,N_14389,N_14103);
nor U14665 (N_14665,N_14219,N_14471);
xnor U14666 (N_14666,N_14497,N_14368);
or U14667 (N_14667,N_14220,N_14194);
and U14668 (N_14668,N_14052,N_14492);
or U14669 (N_14669,N_14319,N_14453);
xor U14670 (N_14670,N_14047,N_14265);
xnor U14671 (N_14671,N_14072,N_14190);
nand U14672 (N_14672,N_14300,N_14202);
or U14673 (N_14673,N_14327,N_14145);
nand U14674 (N_14674,N_14200,N_14116);
xnor U14675 (N_14675,N_14418,N_14322);
nand U14676 (N_14676,N_14205,N_14098);
and U14677 (N_14677,N_14233,N_14144);
or U14678 (N_14678,N_14362,N_14027);
and U14679 (N_14679,N_14238,N_14154);
nor U14680 (N_14680,N_14234,N_14296);
nand U14681 (N_14681,N_14262,N_14464);
and U14682 (N_14682,N_14253,N_14284);
nor U14683 (N_14683,N_14013,N_14282);
or U14684 (N_14684,N_14473,N_14408);
and U14685 (N_14685,N_14316,N_14063);
or U14686 (N_14686,N_14164,N_14126);
xor U14687 (N_14687,N_14495,N_14363);
nand U14688 (N_14688,N_14294,N_14237);
or U14689 (N_14689,N_14149,N_14060);
xor U14690 (N_14690,N_14058,N_14044);
or U14691 (N_14691,N_14461,N_14189);
nor U14692 (N_14692,N_14256,N_14075);
nor U14693 (N_14693,N_14321,N_14250);
nand U14694 (N_14694,N_14178,N_14038);
and U14695 (N_14695,N_14447,N_14271);
xnor U14696 (N_14696,N_14131,N_14146);
xnor U14697 (N_14697,N_14074,N_14012);
nand U14698 (N_14698,N_14243,N_14395);
nor U14699 (N_14699,N_14007,N_14094);
and U14700 (N_14700,N_14056,N_14435);
and U14701 (N_14701,N_14465,N_14488);
xor U14702 (N_14702,N_14413,N_14187);
and U14703 (N_14703,N_14011,N_14206);
nor U14704 (N_14704,N_14244,N_14176);
and U14705 (N_14705,N_14494,N_14348);
xor U14706 (N_14706,N_14004,N_14010);
or U14707 (N_14707,N_14496,N_14299);
nor U14708 (N_14708,N_14295,N_14460);
or U14709 (N_14709,N_14127,N_14293);
and U14710 (N_14710,N_14061,N_14493);
nand U14711 (N_14711,N_14467,N_14347);
nor U14712 (N_14712,N_14215,N_14279);
nand U14713 (N_14713,N_14301,N_14266);
nor U14714 (N_14714,N_14313,N_14396);
xor U14715 (N_14715,N_14386,N_14366);
xnor U14716 (N_14716,N_14213,N_14133);
nand U14717 (N_14717,N_14405,N_14388);
and U14718 (N_14718,N_14498,N_14372);
xor U14719 (N_14719,N_14390,N_14035);
nand U14720 (N_14720,N_14121,N_14358);
nor U14721 (N_14721,N_14309,N_14308);
or U14722 (N_14722,N_14054,N_14485);
nor U14723 (N_14723,N_14000,N_14303);
or U14724 (N_14724,N_14462,N_14364);
or U14725 (N_14725,N_14034,N_14277);
or U14726 (N_14726,N_14268,N_14179);
xnor U14727 (N_14727,N_14174,N_14135);
nand U14728 (N_14728,N_14085,N_14167);
and U14729 (N_14729,N_14329,N_14032);
xnor U14730 (N_14730,N_14201,N_14216);
xnor U14731 (N_14731,N_14383,N_14246);
or U14732 (N_14732,N_14264,N_14458);
or U14733 (N_14733,N_14077,N_14323);
nand U14734 (N_14734,N_14132,N_14499);
or U14735 (N_14735,N_14470,N_14391);
nor U14736 (N_14736,N_14248,N_14402);
nor U14737 (N_14737,N_14161,N_14315);
nand U14738 (N_14738,N_14236,N_14177);
and U14739 (N_14739,N_14089,N_14096);
nor U14740 (N_14740,N_14410,N_14082);
and U14741 (N_14741,N_14337,N_14340);
nor U14742 (N_14742,N_14125,N_14302);
and U14743 (N_14743,N_14025,N_14425);
or U14744 (N_14744,N_14378,N_14474);
nor U14745 (N_14745,N_14240,N_14325);
or U14746 (N_14746,N_14344,N_14252);
or U14747 (N_14747,N_14257,N_14181);
nand U14748 (N_14748,N_14349,N_14417);
and U14749 (N_14749,N_14260,N_14353);
nor U14750 (N_14750,N_14454,N_14451);
nor U14751 (N_14751,N_14415,N_14142);
nor U14752 (N_14752,N_14113,N_14029);
or U14753 (N_14753,N_14453,N_14493);
or U14754 (N_14754,N_14316,N_14134);
xor U14755 (N_14755,N_14048,N_14383);
nor U14756 (N_14756,N_14382,N_14411);
nor U14757 (N_14757,N_14438,N_14375);
xnor U14758 (N_14758,N_14128,N_14299);
or U14759 (N_14759,N_14281,N_14117);
xnor U14760 (N_14760,N_14278,N_14405);
nand U14761 (N_14761,N_14249,N_14125);
or U14762 (N_14762,N_14434,N_14037);
xnor U14763 (N_14763,N_14365,N_14106);
and U14764 (N_14764,N_14082,N_14141);
or U14765 (N_14765,N_14083,N_14210);
nand U14766 (N_14766,N_14189,N_14111);
and U14767 (N_14767,N_14378,N_14064);
xor U14768 (N_14768,N_14225,N_14140);
xnor U14769 (N_14769,N_14416,N_14317);
nor U14770 (N_14770,N_14337,N_14008);
xnor U14771 (N_14771,N_14142,N_14013);
nor U14772 (N_14772,N_14288,N_14254);
or U14773 (N_14773,N_14396,N_14399);
or U14774 (N_14774,N_14327,N_14236);
xnor U14775 (N_14775,N_14316,N_14179);
xor U14776 (N_14776,N_14393,N_14371);
xnor U14777 (N_14777,N_14435,N_14162);
xor U14778 (N_14778,N_14151,N_14060);
xor U14779 (N_14779,N_14211,N_14318);
and U14780 (N_14780,N_14353,N_14251);
and U14781 (N_14781,N_14116,N_14315);
nand U14782 (N_14782,N_14416,N_14021);
and U14783 (N_14783,N_14361,N_14038);
nand U14784 (N_14784,N_14164,N_14177);
xnor U14785 (N_14785,N_14166,N_14080);
or U14786 (N_14786,N_14113,N_14198);
xor U14787 (N_14787,N_14338,N_14133);
or U14788 (N_14788,N_14093,N_14224);
and U14789 (N_14789,N_14041,N_14430);
nand U14790 (N_14790,N_14171,N_14144);
and U14791 (N_14791,N_14223,N_14327);
nor U14792 (N_14792,N_14412,N_14183);
or U14793 (N_14793,N_14167,N_14457);
and U14794 (N_14794,N_14184,N_14403);
and U14795 (N_14795,N_14021,N_14342);
xor U14796 (N_14796,N_14299,N_14350);
and U14797 (N_14797,N_14482,N_14270);
nor U14798 (N_14798,N_14312,N_14076);
xnor U14799 (N_14799,N_14254,N_14209);
or U14800 (N_14800,N_14428,N_14204);
nor U14801 (N_14801,N_14331,N_14114);
and U14802 (N_14802,N_14179,N_14497);
or U14803 (N_14803,N_14064,N_14036);
and U14804 (N_14804,N_14105,N_14114);
or U14805 (N_14805,N_14460,N_14225);
xnor U14806 (N_14806,N_14414,N_14365);
nand U14807 (N_14807,N_14203,N_14212);
and U14808 (N_14808,N_14083,N_14076);
nor U14809 (N_14809,N_14472,N_14177);
nor U14810 (N_14810,N_14311,N_14352);
nand U14811 (N_14811,N_14076,N_14067);
and U14812 (N_14812,N_14462,N_14341);
nor U14813 (N_14813,N_14371,N_14223);
or U14814 (N_14814,N_14198,N_14300);
nand U14815 (N_14815,N_14295,N_14031);
and U14816 (N_14816,N_14262,N_14294);
or U14817 (N_14817,N_14099,N_14209);
or U14818 (N_14818,N_14224,N_14185);
nor U14819 (N_14819,N_14378,N_14241);
or U14820 (N_14820,N_14143,N_14038);
or U14821 (N_14821,N_14278,N_14491);
xor U14822 (N_14822,N_14309,N_14407);
nand U14823 (N_14823,N_14010,N_14050);
or U14824 (N_14824,N_14415,N_14086);
or U14825 (N_14825,N_14280,N_14368);
and U14826 (N_14826,N_14398,N_14394);
and U14827 (N_14827,N_14080,N_14028);
xnor U14828 (N_14828,N_14002,N_14413);
or U14829 (N_14829,N_14116,N_14155);
xnor U14830 (N_14830,N_14150,N_14109);
and U14831 (N_14831,N_14365,N_14218);
nor U14832 (N_14832,N_14378,N_14374);
nand U14833 (N_14833,N_14229,N_14224);
xor U14834 (N_14834,N_14463,N_14369);
xnor U14835 (N_14835,N_14429,N_14279);
or U14836 (N_14836,N_14051,N_14391);
nor U14837 (N_14837,N_14097,N_14202);
nor U14838 (N_14838,N_14272,N_14129);
and U14839 (N_14839,N_14468,N_14235);
or U14840 (N_14840,N_14350,N_14409);
nor U14841 (N_14841,N_14101,N_14421);
nand U14842 (N_14842,N_14219,N_14250);
xor U14843 (N_14843,N_14410,N_14246);
and U14844 (N_14844,N_14321,N_14393);
or U14845 (N_14845,N_14105,N_14207);
or U14846 (N_14846,N_14395,N_14269);
xnor U14847 (N_14847,N_14080,N_14211);
or U14848 (N_14848,N_14139,N_14432);
and U14849 (N_14849,N_14322,N_14318);
nor U14850 (N_14850,N_14367,N_14311);
and U14851 (N_14851,N_14318,N_14136);
xnor U14852 (N_14852,N_14048,N_14420);
and U14853 (N_14853,N_14329,N_14205);
or U14854 (N_14854,N_14246,N_14249);
or U14855 (N_14855,N_14310,N_14117);
xor U14856 (N_14856,N_14071,N_14492);
nor U14857 (N_14857,N_14288,N_14088);
and U14858 (N_14858,N_14124,N_14217);
or U14859 (N_14859,N_14410,N_14400);
xor U14860 (N_14860,N_14203,N_14141);
or U14861 (N_14861,N_14114,N_14076);
nor U14862 (N_14862,N_14422,N_14018);
xor U14863 (N_14863,N_14005,N_14184);
xor U14864 (N_14864,N_14050,N_14167);
nand U14865 (N_14865,N_14243,N_14161);
nand U14866 (N_14866,N_14214,N_14396);
nor U14867 (N_14867,N_14423,N_14158);
xor U14868 (N_14868,N_14416,N_14253);
nor U14869 (N_14869,N_14367,N_14271);
or U14870 (N_14870,N_14397,N_14432);
or U14871 (N_14871,N_14198,N_14032);
or U14872 (N_14872,N_14051,N_14008);
and U14873 (N_14873,N_14233,N_14412);
or U14874 (N_14874,N_14447,N_14360);
nor U14875 (N_14875,N_14495,N_14073);
nor U14876 (N_14876,N_14360,N_14394);
xor U14877 (N_14877,N_14240,N_14170);
nand U14878 (N_14878,N_14196,N_14071);
nor U14879 (N_14879,N_14232,N_14388);
or U14880 (N_14880,N_14304,N_14119);
or U14881 (N_14881,N_14492,N_14158);
and U14882 (N_14882,N_14358,N_14261);
and U14883 (N_14883,N_14112,N_14061);
or U14884 (N_14884,N_14424,N_14050);
nand U14885 (N_14885,N_14098,N_14151);
nand U14886 (N_14886,N_14354,N_14383);
nand U14887 (N_14887,N_14197,N_14439);
nand U14888 (N_14888,N_14060,N_14412);
and U14889 (N_14889,N_14356,N_14185);
xor U14890 (N_14890,N_14224,N_14048);
xnor U14891 (N_14891,N_14334,N_14199);
nand U14892 (N_14892,N_14148,N_14223);
and U14893 (N_14893,N_14239,N_14301);
xor U14894 (N_14894,N_14254,N_14107);
nor U14895 (N_14895,N_14115,N_14081);
nand U14896 (N_14896,N_14350,N_14265);
nor U14897 (N_14897,N_14318,N_14012);
nor U14898 (N_14898,N_14225,N_14404);
xor U14899 (N_14899,N_14286,N_14051);
and U14900 (N_14900,N_14391,N_14499);
or U14901 (N_14901,N_14446,N_14063);
nand U14902 (N_14902,N_14022,N_14191);
xnor U14903 (N_14903,N_14005,N_14292);
xor U14904 (N_14904,N_14014,N_14127);
xor U14905 (N_14905,N_14079,N_14284);
nand U14906 (N_14906,N_14413,N_14105);
nor U14907 (N_14907,N_14440,N_14116);
nor U14908 (N_14908,N_14087,N_14368);
xnor U14909 (N_14909,N_14220,N_14179);
xnor U14910 (N_14910,N_14136,N_14311);
or U14911 (N_14911,N_14166,N_14358);
nand U14912 (N_14912,N_14153,N_14266);
and U14913 (N_14913,N_14183,N_14268);
and U14914 (N_14914,N_14362,N_14225);
xor U14915 (N_14915,N_14368,N_14269);
and U14916 (N_14916,N_14128,N_14421);
and U14917 (N_14917,N_14203,N_14430);
nand U14918 (N_14918,N_14320,N_14462);
or U14919 (N_14919,N_14419,N_14174);
nand U14920 (N_14920,N_14471,N_14069);
or U14921 (N_14921,N_14272,N_14421);
or U14922 (N_14922,N_14438,N_14086);
nor U14923 (N_14923,N_14111,N_14399);
or U14924 (N_14924,N_14098,N_14107);
nand U14925 (N_14925,N_14486,N_14253);
nand U14926 (N_14926,N_14153,N_14440);
and U14927 (N_14927,N_14062,N_14251);
xnor U14928 (N_14928,N_14092,N_14306);
and U14929 (N_14929,N_14080,N_14240);
nor U14930 (N_14930,N_14183,N_14013);
nand U14931 (N_14931,N_14149,N_14215);
nand U14932 (N_14932,N_14435,N_14335);
and U14933 (N_14933,N_14226,N_14458);
and U14934 (N_14934,N_14283,N_14273);
nor U14935 (N_14935,N_14490,N_14135);
nand U14936 (N_14936,N_14439,N_14026);
nand U14937 (N_14937,N_14369,N_14432);
nand U14938 (N_14938,N_14297,N_14185);
and U14939 (N_14939,N_14128,N_14492);
xor U14940 (N_14940,N_14446,N_14280);
and U14941 (N_14941,N_14365,N_14451);
and U14942 (N_14942,N_14440,N_14338);
and U14943 (N_14943,N_14300,N_14135);
xor U14944 (N_14944,N_14275,N_14011);
and U14945 (N_14945,N_14329,N_14491);
and U14946 (N_14946,N_14221,N_14377);
or U14947 (N_14947,N_14121,N_14125);
xnor U14948 (N_14948,N_14011,N_14182);
and U14949 (N_14949,N_14297,N_14256);
xor U14950 (N_14950,N_14467,N_14335);
nand U14951 (N_14951,N_14085,N_14155);
and U14952 (N_14952,N_14096,N_14139);
and U14953 (N_14953,N_14180,N_14246);
nand U14954 (N_14954,N_14048,N_14203);
and U14955 (N_14955,N_14086,N_14338);
nor U14956 (N_14956,N_14097,N_14127);
nor U14957 (N_14957,N_14074,N_14318);
nand U14958 (N_14958,N_14317,N_14000);
xor U14959 (N_14959,N_14429,N_14241);
or U14960 (N_14960,N_14103,N_14114);
xnor U14961 (N_14961,N_14051,N_14477);
or U14962 (N_14962,N_14214,N_14009);
xnor U14963 (N_14963,N_14345,N_14030);
xor U14964 (N_14964,N_14132,N_14308);
nand U14965 (N_14965,N_14118,N_14405);
nand U14966 (N_14966,N_14018,N_14483);
and U14967 (N_14967,N_14453,N_14412);
and U14968 (N_14968,N_14346,N_14122);
nand U14969 (N_14969,N_14341,N_14221);
nand U14970 (N_14970,N_14442,N_14233);
or U14971 (N_14971,N_14176,N_14441);
or U14972 (N_14972,N_14443,N_14135);
or U14973 (N_14973,N_14309,N_14366);
nand U14974 (N_14974,N_14094,N_14299);
xnor U14975 (N_14975,N_14228,N_14278);
xor U14976 (N_14976,N_14496,N_14465);
and U14977 (N_14977,N_14492,N_14497);
nor U14978 (N_14978,N_14385,N_14424);
nor U14979 (N_14979,N_14247,N_14342);
nand U14980 (N_14980,N_14396,N_14477);
or U14981 (N_14981,N_14150,N_14378);
nand U14982 (N_14982,N_14061,N_14003);
nand U14983 (N_14983,N_14200,N_14093);
or U14984 (N_14984,N_14463,N_14303);
nand U14985 (N_14985,N_14250,N_14116);
nor U14986 (N_14986,N_14278,N_14355);
nand U14987 (N_14987,N_14083,N_14169);
xor U14988 (N_14988,N_14316,N_14303);
nand U14989 (N_14989,N_14309,N_14222);
xor U14990 (N_14990,N_14252,N_14064);
nand U14991 (N_14991,N_14075,N_14311);
and U14992 (N_14992,N_14025,N_14105);
xor U14993 (N_14993,N_14496,N_14270);
nor U14994 (N_14994,N_14444,N_14206);
or U14995 (N_14995,N_14143,N_14455);
and U14996 (N_14996,N_14328,N_14456);
xor U14997 (N_14997,N_14117,N_14297);
and U14998 (N_14998,N_14206,N_14270);
nand U14999 (N_14999,N_14176,N_14315);
or UO_0 (O_0,N_14970,N_14687);
xnor UO_1 (O_1,N_14545,N_14636);
nand UO_2 (O_2,N_14582,N_14624);
xor UO_3 (O_3,N_14853,N_14862);
xor UO_4 (O_4,N_14888,N_14891);
and UO_5 (O_5,N_14851,N_14659);
nor UO_6 (O_6,N_14897,N_14592);
nor UO_7 (O_7,N_14773,N_14701);
and UO_8 (O_8,N_14657,N_14625);
xnor UO_9 (O_9,N_14716,N_14777);
nor UO_10 (O_10,N_14560,N_14571);
xnor UO_11 (O_11,N_14858,N_14892);
xnor UO_12 (O_12,N_14904,N_14641);
and UO_13 (O_13,N_14983,N_14867);
xnor UO_14 (O_14,N_14623,N_14693);
nor UO_15 (O_15,N_14935,N_14981);
nor UO_16 (O_16,N_14845,N_14815);
or UO_17 (O_17,N_14588,N_14916);
nand UO_18 (O_18,N_14943,N_14570);
xnor UO_19 (O_19,N_14748,N_14667);
nand UO_20 (O_20,N_14802,N_14534);
nor UO_21 (O_21,N_14756,N_14686);
xor UO_22 (O_22,N_14562,N_14599);
nand UO_23 (O_23,N_14835,N_14601);
xor UO_24 (O_24,N_14979,N_14895);
nor UO_25 (O_25,N_14648,N_14722);
nand UO_26 (O_26,N_14512,N_14913);
or UO_27 (O_27,N_14663,N_14603);
xnor UO_28 (O_28,N_14880,N_14600);
xnor UO_29 (O_29,N_14967,N_14776);
xor UO_30 (O_30,N_14695,N_14549);
or UO_31 (O_31,N_14676,N_14989);
nor UO_32 (O_32,N_14741,N_14666);
nor UO_33 (O_33,N_14922,N_14712);
xor UO_34 (O_34,N_14850,N_14863);
xor UO_35 (O_35,N_14902,N_14555);
and UO_36 (O_36,N_14665,N_14679);
nor UO_37 (O_37,N_14515,N_14804);
or UO_38 (O_38,N_14841,N_14668);
nor UO_39 (O_39,N_14957,N_14501);
nand UO_40 (O_40,N_14511,N_14627);
xor UO_41 (O_41,N_14865,N_14807);
xor UO_42 (O_42,N_14813,N_14567);
or UO_43 (O_43,N_14610,N_14972);
xor UO_44 (O_44,N_14608,N_14889);
and UO_45 (O_45,N_14751,N_14682);
or UO_46 (O_46,N_14994,N_14612);
xnor UO_47 (O_47,N_14921,N_14569);
nor UO_48 (O_48,N_14514,N_14925);
or UO_49 (O_49,N_14951,N_14558);
xnor UO_50 (O_50,N_14525,N_14688);
nor UO_51 (O_51,N_14597,N_14763);
xor UO_52 (O_52,N_14803,N_14689);
nor UO_53 (O_53,N_14816,N_14842);
and UO_54 (O_54,N_14932,N_14953);
xor UO_55 (O_55,N_14596,N_14540);
and UO_56 (O_56,N_14868,N_14557);
or UO_57 (O_57,N_14505,N_14517);
and UO_58 (O_58,N_14664,N_14723);
and UO_59 (O_59,N_14531,N_14772);
xor UO_60 (O_60,N_14926,N_14528);
nand UO_61 (O_61,N_14946,N_14632);
or UO_62 (O_62,N_14546,N_14556);
or UO_63 (O_63,N_14566,N_14702);
nor UO_64 (O_64,N_14767,N_14878);
xor UO_65 (O_65,N_14640,N_14854);
or UO_66 (O_66,N_14784,N_14912);
or UO_67 (O_67,N_14616,N_14621);
nand UO_68 (O_68,N_14905,N_14948);
or UO_69 (O_69,N_14662,N_14919);
xor UO_70 (O_70,N_14982,N_14931);
nor UO_71 (O_71,N_14780,N_14585);
xor UO_72 (O_72,N_14530,N_14734);
nand UO_73 (O_73,N_14990,N_14604);
nand UO_74 (O_74,N_14898,N_14728);
nor UO_75 (O_75,N_14911,N_14626);
nand UO_76 (O_76,N_14848,N_14633);
xor UO_77 (O_77,N_14532,N_14575);
nor UO_78 (O_78,N_14876,N_14749);
xnor UO_79 (O_79,N_14602,N_14713);
nor UO_80 (O_80,N_14811,N_14826);
and UO_81 (O_81,N_14565,N_14580);
or UO_82 (O_82,N_14730,N_14928);
or UO_83 (O_83,N_14699,N_14870);
xor UO_84 (O_84,N_14832,N_14955);
nor UO_85 (O_85,N_14934,N_14759);
nand UO_86 (O_86,N_14704,N_14538);
nand UO_87 (O_87,N_14903,N_14731);
nand UO_88 (O_88,N_14881,N_14890);
xor UO_89 (O_89,N_14718,N_14579);
xor UO_90 (O_90,N_14521,N_14944);
and UO_91 (O_91,N_14942,N_14871);
nand UO_92 (O_92,N_14980,N_14812);
xnor UO_93 (O_93,N_14875,N_14615);
nand UO_94 (O_94,N_14987,N_14586);
nand UO_95 (O_95,N_14938,N_14568);
nor UO_96 (O_96,N_14508,N_14866);
xor UO_97 (O_97,N_14824,N_14522);
nand UO_98 (O_98,N_14527,N_14707);
nor UO_99 (O_99,N_14869,N_14945);
and UO_100 (O_100,N_14852,N_14859);
xor UO_101 (O_101,N_14809,N_14752);
nand UO_102 (O_102,N_14769,N_14790);
nand UO_103 (O_103,N_14651,N_14598);
xnor UO_104 (O_104,N_14743,N_14793);
or UO_105 (O_105,N_14761,N_14960);
and UO_106 (O_106,N_14893,N_14680);
or UO_107 (O_107,N_14638,N_14618);
and UO_108 (O_108,N_14894,N_14703);
or UO_109 (O_109,N_14744,N_14705);
nor UO_110 (O_110,N_14768,N_14634);
xnor UO_111 (O_111,N_14739,N_14721);
nor UO_112 (O_112,N_14978,N_14954);
nor UO_113 (O_113,N_14860,N_14553);
or UO_114 (O_114,N_14573,N_14649);
nand UO_115 (O_115,N_14940,N_14698);
nand UO_116 (O_116,N_14593,N_14786);
and UO_117 (O_117,N_14988,N_14520);
nand UO_118 (O_118,N_14840,N_14963);
nand UO_119 (O_119,N_14941,N_14821);
nand UO_120 (O_120,N_14918,N_14681);
nand UO_121 (O_121,N_14678,N_14537);
nand UO_122 (O_122,N_14690,N_14855);
or UO_123 (O_123,N_14754,N_14552);
nand UO_124 (O_124,N_14559,N_14643);
xor UO_125 (O_125,N_14827,N_14991);
xor UO_126 (O_126,N_14877,N_14986);
xor UO_127 (O_127,N_14736,N_14965);
and UO_128 (O_128,N_14781,N_14828);
or UO_129 (O_129,N_14823,N_14923);
nor UO_130 (O_130,N_14766,N_14746);
or UO_131 (O_131,N_14849,N_14509);
nand UO_132 (O_132,N_14639,N_14874);
nor UO_133 (O_133,N_14727,N_14765);
and UO_134 (O_134,N_14544,N_14714);
nand UO_135 (O_135,N_14645,N_14795);
and UO_136 (O_136,N_14720,N_14536);
or UO_137 (O_137,N_14920,N_14740);
and UO_138 (O_138,N_14952,N_14959);
and UO_139 (O_139,N_14782,N_14861);
nand UO_140 (O_140,N_14783,N_14770);
nor UO_141 (O_141,N_14884,N_14958);
nor UO_142 (O_142,N_14882,N_14885);
nor UO_143 (O_143,N_14587,N_14726);
nand UO_144 (O_144,N_14785,N_14864);
nor UO_145 (O_145,N_14900,N_14886);
xor UO_146 (O_146,N_14937,N_14629);
nor UO_147 (O_147,N_14654,N_14798);
and UO_148 (O_148,N_14755,N_14594);
nor UO_149 (O_149,N_14605,N_14924);
nand UO_150 (O_150,N_14735,N_14995);
nor UO_151 (O_151,N_14706,N_14561);
nor UO_152 (O_152,N_14578,N_14810);
or UO_153 (O_153,N_14622,N_14516);
and UO_154 (O_154,N_14791,N_14529);
nor UO_155 (O_155,N_14523,N_14883);
nor UO_156 (O_156,N_14822,N_14825);
xnor UO_157 (O_157,N_14694,N_14539);
nor UO_158 (O_158,N_14742,N_14507);
or UO_159 (O_159,N_14787,N_14669);
xor UO_160 (O_160,N_14611,N_14844);
nand UO_161 (O_161,N_14647,N_14677);
nand UO_162 (O_162,N_14652,N_14576);
and UO_163 (O_163,N_14554,N_14590);
or UO_164 (O_164,N_14907,N_14541);
nand UO_165 (O_165,N_14819,N_14563);
xor UO_166 (O_166,N_14917,N_14500);
nor UO_167 (O_167,N_14843,N_14502);
nand UO_168 (O_168,N_14646,N_14901);
nand UO_169 (O_169,N_14733,N_14595);
and UO_170 (O_170,N_14760,N_14831);
xor UO_171 (O_171,N_14543,N_14533);
nand UO_172 (O_172,N_14504,N_14614);
nand UO_173 (O_173,N_14909,N_14789);
xor UO_174 (O_174,N_14887,N_14985);
xnor UO_175 (O_175,N_14591,N_14830);
xor UO_176 (O_176,N_14933,N_14758);
nor UO_177 (O_177,N_14974,N_14656);
nor UO_178 (O_178,N_14839,N_14794);
and UO_179 (O_179,N_14535,N_14673);
nor UO_180 (O_180,N_14631,N_14856);
nor UO_181 (O_181,N_14674,N_14750);
nand UO_182 (O_182,N_14797,N_14799);
xor UO_183 (O_183,N_14910,N_14607);
xnor UO_184 (O_184,N_14998,N_14524);
and UO_185 (O_185,N_14915,N_14729);
and UO_186 (O_186,N_14962,N_14606);
xor UO_187 (O_187,N_14550,N_14619);
and UO_188 (O_188,N_14992,N_14817);
and UO_189 (O_189,N_14717,N_14655);
xor UO_190 (O_190,N_14719,N_14589);
nand UO_191 (O_191,N_14513,N_14642);
or UO_192 (O_192,N_14929,N_14745);
nand UO_193 (O_193,N_14617,N_14834);
nor UO_194 (O_194,N_14732,N_14930);
or UO_195 (O_195,N_14738,N_14757);
nor UO_196 (O_196,N_14950,N_14711);
nor UO_197 (O_197,N_14526,N_14684);
and UO_198 (O_198,N_14838,N_14996);
or UO_199 (O_199,N_14966,N_14753);
xor UO_200 (O_200,N_14683,N_14961);
or UO_201 (O_201,N_14939,N_14542);
or UO_202 (O_202,N_14806,N_14650);
xnor UO_203 (O_203,N_14872,N_14700);
and UO_204 (O_204,N_14778,N_14964);
nor UO_205 (O_205,N_14691,N_14837);
or UO_206 (O_206,N_14653,N_14792);
nor UO_207 (O_207,N_14914,N_14697);
xnor UO_208 (O_208,N_14947,N_14788);
and UO_209 (O_209,N_14801,N_14975);
xnor UO_210 (O_210,N_14997,N_14908);
xor UO_211 (O_211,N_14637,N_14808);
nand UO_212 (O_212,N_14628,N_14692);
nor UO_213 (O_213,N_14936,N_14969);
nor UO_214 (O_214,N_14779,N_14581);
nand UO_215 (O_215,N_14899,N_14661);
or UO_216 (O_216,N_14609,N_14747);
nor UO_217 (O_217,N_14548,N_14724);
nand UO_218 (O_218,N_14572,N_14685);
nor UO_219 (O_219,N_14503,N_14956);
nor UO_220 (O_220,N_14630,N_14708);
nor UO_221 (O_221,N_14993,N_14820);
nand UO_222 (O_222,N_14675,N_14949);
or UO_223 (O_223,N_14577,N_14574);
nor UO_224 (O_224,N_14518,N_14510);
xor UO_225 (O_225,N_14564,N_14818);
xor UO_226 (O_226,N_14971,N_14771);
or UO_227 (O_227,N_14999,N_14800);
nor UO_228 (O_228,N_14805,N_14984);
or UO_229 (O_229,N_14846,N_14879);
and UO_230 (O_230,N_14762,N_14774);
xor UO_231 (O_231,N_14670,N_14613);
nor UO_232 (O_232,N_14906,N_14709);
and UO_233 (O_233,N_14506,N_14658);
or UO_234 (O_234,N_14829,N_14519);
xor UO_235 (O_235,N_14671,N_14977);
nand UO_236 (O_236,N_14715,N_14644);
and UO_237 (O_237,N_14836,N_14547);
and UO_238 (O_238,N_14896,N_14660);
nor UO_239 (O_239,N_14976,N_14973);
or UO_240 (O_240,N_14847,N_14927);
xnor UO_241 (O_241,N_14725,N_14635);
and UO_242 (O_242,N_14857,N_14620);
and UO_243 (O_243,N_14873,N_14968);
xnor UO_244 (O_244,N_14583,N_14775);
nor UO_245 (O_245,N_14584,N_14814);
and UO_246 (O_246,N_14551,N_14710);
and UO_247 (O_247,N_14696,N_14737);
and UO_248 (O_248,N_14796,N_14672);
nand UO_249 (O_249,N_14764,N_14833);
xor UO_250 (O_250,N_14693,N_14710);
and UO_251 (O_251,N_14788,N_14769);
or UO_252 (O_252,N_14887,N_14722);
nor UO_253 (O_253,N_14625,N_14631);
and UO_254 (O_254,N_14758,N_14501);
nand UO_255 (O_255,N_14661,N_14681);
or UO_256 (O_256,N_14992,N_14872);
nor UO_257 (O_257,N_14726,N_14802);
or UO_258 (O_258,N_14979,N_14562);
or UO_259 (O_259,N_14829,N_14773);
nor UO_260 (O_260,N_14540,N_14717);
nor UO_261 (O_261,N_14860,N_14847);
and UO_262 (O_262,N_14853,N_14917);
xor UO_263 (O_263,N_14997,N_14628);
or UO_264 (O_264,N_14787,N_14796);
xnor UO_265 (O_265,N_14610,N_14524);
or UO_266 (O_266,N_14582,N_14993);
or UO_267 (O_267,N_14743,N_14738);
nand UO_268 (O_268,N_14824,N_14539);
nand UO_269 (O_269,N_14941,N_14935);
or UO_270 (O_270,N_14665,N_14732);
nor UO_271 (O_271,N_14806,N_14966);
and UO_272 (O_272,N_14702,N_14618);
nor UO_273 (O_273,N_14928,N_14752);
nand UO_274 (O_274,N_14844,N_14786);
nor UO_275 (O_275,N_14846,N_14896);
nor UO_276 (O_276,N_14641,N_14618);
and UO_277 (O_277,N_14866,N_14954);
nor UO_278 (O_278,N_14826,N_14521);
and UO_279 (O_279,N_14681,N_14546);
xnor UO_280 (O_280,N_14582,N_14859);
nor UO_281 (O_281,N_14720,N_14503);
and UO_282 (O_282,N_14977,N_14688);
and UO_283 (O_283,N_14663,N_14943);
xor UO_284 (O_284,N_14979,N_14576);
xor UO_285 (O_285,N_14960,N_14685);
and UO_286 (O_286,N_14860,N_14887);
nand UO_287 (O_287,N_14925,N_14795);
nor UO_288 (O_288,N_14943,N_14786);
and UO_289 (O_289,N_14741,N_14890);
xor UO_290 (O_290,N_14804,N_14817);
and UO_291 (O_291,N_14727,N_14916);
xor UO_292 (O_292,N_14557,N_14631);
and UO_293 (O_293,N_14731,N_14818);
xor UO_294 (O_294,N_14891,N_14772);
nor UO_295 (O_295,N_14505,N_14547);
xnor UO_296 (O_296,N_14731,N_14797);
nor UO_297 (O_297,N_14829,N_14767);
nor UO_298 (O_298,N_14542,N_14735);
or UO_299 (O_299,N_14787,N_14559);
nand UO_300 (O_300,N_14705,N_14599);
and UO_301 (O_301,N_14549,N_14511);
and UO_302 (O_302,N_14692,N_14912);
or UO_303 (O_303,N_14805,N_14843);
and UO_304 (O_304,N_14582,N_14724);
and UO_305 (O_305,N_14605,N_14773);
nand UO_306 (O_306,N_14873,N_14897);
xor UO_307 (O_307,N_14853,N_14825);
nor UO_308 (O_308,N_14719,N_14529);
xor UO_309 (O_309,N_14731,N_14926);
or UO_310 (O_310,N_14580,N_14540);
nor UO_311 (O_311,N_14566,N_14705);
or UO_312 (O_312,N_14651,N_14599);
xnor UO_313 (O_313,N_14714,N_14660);
nand UO_314 (O_314,N_14785,N_14882);
or UO_315 (O_315,N_14620,N_14934);
nor UO_316 (O_316,N_14629,N_14687);
nand UO_317 (O_317,N_14677,N_14798);
nor UO_318 (O_318,N_14854,N_14790);
and UO_319 (O_319,N_14770,N_14586);
nand UO_320 (O_320,N_14951,N_14535);
nor UO_321 (O_321,N_14749,N_14899);
and UO_322 (O_322,N_14881,N_14616);
or UO_323 (O_323,N_14750,N_14777);
or UO_324 (O_324,N_14853,N_14514);
and UO_325 (O_325,N_14823,N_14560);
and UO_326 (O_326,N_14706,N_14992);
nor UO_327 (O_327,N_14721,N_14753);
nor UO_328 (O_328,N_14776,N_14815);
xor UO_329 (O_329,N_14710,N_14608);
nand UO_330 (O_330,N_14926,N_14761);
nand UO_331 (O_331,N_14626,N_14693);
nor UO_332 (O_332,N_14983,N_14742);
nor UO_333 (O_333,N_14753,N_14904);
xnor UO_334 (O_334,N_14806,N_14701);
xor UO_335 (O_335,N_14625,N_14596);
and UO_336 (O_336,N_14610,N_14821);
or UO_337 (O_337,N_14815,N_14953);
nand UO_338 (O_338,N_14701,N_14532);
and UO_339 (O_339,N_14829,N_14718);
and UO_340 (O_340,N_14959,N_14895);
xnor UO_341 (O_341,N_14542,N_14723);
or UO_342 (O_342,N_14528,N_14802);
xor UO_343 (O_343,N_14636,N_14881);
or UO_344 (O_344,N_14918,N_14884);
nor UO_345 (O_345,N_14879,N_14940);
nor UO_346 (O_346,N_14513,N_14841);
or UO_347 (O_347,N_14826,N_14673);
or UO_348 (O_348,N_14998,N_14552);
nand UO_349 (O_349,N_14757,N_14943);
xor UO_350 (O_350,N_14542,N_14962);
or UO_351 (O_351,N_14957,N_14846);
and UO_352 (O_352,N_14624,N_14751);
nand UO_353 (O_353,N_14604,N_14502);
or UO_354 (O_354,N_14855,N_14718);
nor UO_355 (O_355,N_14958,N_14607);
or UO_356 (O_356,N_14633,N_14802);
nand UO_357 (O_357,N_14777,N_14744);
or UO_358 (O_358,N_14629,N_14993);
or UO_359 (O_359,N_14868,N_14861);
xnor UO_360 (O_360,N_14555,N_14795);
or UO_361 (O_361,N_14762,N_14647);
xor UO_362 (O_362,N_14994,N_14504);
or UO_363 (O_363,N_14572,N_14832);
nor UO_364 (O_364,N_14840,N_14519);
xnor UO_365 (O_365,N_14692,N_14774);
or UO_366 (O_366,N_14796,N_14722);
nor UO_367 (O_367,N_14737,N_14623);
nand UO_368 (O_368,N_14856,N_14698);
or UO_369 (O_369,N_14986,N_14893);
and UO_370 (O_370,N_14962,N_14620);
or UO_371 (O_371,N_14678,N_14524);
or UO_372 (O_372,N_14943,N_14751);
nand UO_373 (O_373,N_14516,N_14962);
nand UO_374 (O_374,N_14720,N_14829);
or UO_375 (O_375,N_14709,N_14502);
nor UO_376 (O_376,N_14829,N_14590);
xor UO_377 (O_377,N_14509,N_14784);
nor UO_378 (O_378,N_14648,N_14644);
nor UO_379 (O_379,N_14842,N_14995);
nand UO_380 (O_380,N_14795,N_14949);
or UO_381 (O_381,N_14952,N_14572);
xnor UO_382 (O_382,N_14661,N_14721);
nand UO_383 (O_383,N_14514,N_14545);
and UO_384 (O_384,N_14815,N_14996);
xnor UO_385 (O_385,N_14789,N_14663);
xnor UO_386 (O_386,N_14538,N_14549);
nor UO_387 (O_387,N_14884,N_14803);
xor UO_388 (O_388,N_14969,N_14527);
and UO_389 (O_389,N_14759,N_14711);
or UO_390 (O_390,N_14885,N_14946);
or UO_391 (O_391,N_14959,N_14793);
xor UO_392 (O_392,N_14696,N_14556);
xor UO_393 (O_393,N_14632,N_14699);
xnor UO_394 (O_394,N_14692,N_14694);
or UO_395 (O_395,N_14693,N_14845);
or UO_396 (O_396,N_14766,N_14542);
xor UO_397 (O_397,N_14598,N_14771);
nand UO_398 (O_398,N_14539,N_14609);
nand UO_399 (O_399,N_14583,N_14563);
nand UO_400 (O_400,N_14693,N_14514);
or UO_401 (O_401,N_14785,N_14892);
nor UO_402 (O_402,N_14988,N_14511);
and UO_403 (O_403,N_14587,N_14912);
nand UO_404 (O_404,N_14966,N_14730);
nor UO_405 (O_405,N_14844,N_14979);
xor UO_406 (O_406,N_14647,N_14778);
and UO_407 (O_407,N_14899,N_14573);
or UO_408 (O_408,N_14779,N_14523);
and UO_409 (O_409,N_14688,N_14627);
nand UO_410 (O_410,N_14582,N_14605);
or UO_411 (O_411,N_14500,N_14952);
xor UO_412 (O_412,N_14693,N_14848);
xor UO_413 (O_413,N_14577,N_14657);
nor UO_414 (O_414,N_14968,N_14527);
xnor UO_415 (O_415,N_14558,N_14750);
nand UO_416 (O_416,N_14727,N_14628);
xnor UO_417 (O_417,N_14869,N_14677);
or UO_418 (O_418,N_14823,N_14975);
nor UO_419 (O_419,N_14649,N_14608);
nor UO_420 (O_420,N_14837,N_14530);
xor UO_421 (O_421,N_14768,N_14824);
and UO_422 (O_422,N_14872,N_14675);
nand UO_423 (O_423,N_14764,N_14711);
or UO_424 (O_424,N_14507,N_14706);
and UO_425 (O_425,N_14794,N_14942);
xor UO_426 (O_426,N_14770,N_14551);
and UO_427 (O_427,N_14631,N_14530);
or UO_428 (O_428,N_14677,N_14930);
nor UO_429 (O_429,N_14854,N_14867);
nor UO_430 (O_430,N_14819,N_14891);
nor UO_431 (O_431,N_14597,N_14831);
xor UO_432 (O_432,N_14984,N_14897);
and UO_433 (O_433,N_14873,N_14685);
or UO_434 (O_434,N_14828,N_14608);
and UO_435 (O_435,N_14541,N_14900);
xnor UO_436 (O_436,N_14924,N_14576);
xnor UO_437 (O_437,N_14542,N_14546);
xnor UO_438 (O_438,N_14523,N_14893);
and UO_439 (O_439,N_14703,N_14504);
or UO_440 (O_440,N_14967,N_14959);
or UO_441 (O_441,N_14556,N_14875);
nand UO_442 (O_442,N_14993,N_14623);
and UO_443 (O_443,N_14805,N_14914);
and UO_444 (O_444,N_14942,N_14877);
or UO_445 (O_445,N_14931,N_14501);
nor UO_446 (O_446,N_14938,N_14998);
nor UO_447 (O_447,N_14530,N_14758);
nand UO_448 (O_448,N_14797,N_14958);
nor UO_449 (O_449,N_14677,N_14712);
nor UO_450 (O_450,N_14847,N_14656);
nor UO_451 (O_451,N_14855,N_14757);
nor UO_452 (O_452,N_14782,N_14731);
or UO_453 (O_453,N_14786,N_14516);
and UO_454 (O_454,N_14519,N_14999);
xor UO_455 (O_455,N_14717,N_14768);
and UO_456 (O_456,N_14648,N_14779);
nand UO_457 (O_457,N_14503,N_14698);
or UO_458 (O_458,N_14972,N_14548);
and UO_459 (O_459,N_14701,N_14996);
or UO_460 (O_460,N_14928,N_14664);
nor UO_461 (O_461,N_14732,N_14597);
xnor UO_462 (O_462,N_14977,N_14997);
or UO_463 (O_463,N_14708,N_14936);
nor UO_464 (O_464,N_14723,N_14817);
xnor UO_465 (O_465,N_14746,N_14691);
or UO_466 (O_466,N_14908,N_14521);
and UO_467 (O_467,N_14767,N_14904);
and UO_468 (O_468,N_14600,N_14759);
and UO_469 (O_469,N_14595,N_14511);
nor UO_470 (O_470,N_14713,N_14974);
nand UO_471 (O_471,N_14614,N_14846);
and UO_472 (O_472,N_14856,N_14566);
nand UO_473 (O_473,N_14935,N_14533);
nor UO_474 (O_474,N_14760,N_14776);
and UO_475 (O_475,N_14582,N_14840);
nand UO_476 (O_476,N_14794,N_14657);
nand UO_477 (O_477,N_14632,N_14828);
and UO_478 (O_478,N_14504,N_14624);
xor UO_479 (O_479,N_14508,N_14940);
or UO_480 (O_480,N_14742,N_14547);
nand UO_481 (O_481,N_14899,N_14897);
nor UO_482 (O_482,N_14535,N_14501);
nand UO_483 (O_483,N_14554,N_14549);
xnor UO_484 (O_484,N_14635,N_14952);
nor UO_485 (O_485,N_14706,N_14604);
xnor UO_486 (O_486,N_14909,N_14577);
nand UO_487 (O_487,N_14503,N_14746);
nand UO_488 (O_488,N_14639,N_14554);
and UO_489 (O_489,N_14884,N_14587);
or UO_490 (O_490,N_14514,N_14615);
nor UO_491 (O_491,N_14886,N_14717);
or UO_492 (O_492,N_14530,N_14520);
nand UO_493 (O_493,N_14914,N_14880);
nand UO_494 (O_494,N_14977,N_14996);
or UO_495 (O_495,N_14949,N_14621);
or UO_496 (O_496,N_14630,N_14559);
xnor UO_497 (O_497,N_14749,N_14954);
xnor UO_498 (O_498,N_14853,N_14506);
xnor UO_499 (O_499,N_14623,N_14974);
nor UO_500 (O_500,N_14602,N_14975);
xnor UO_501 (O_501,N_14924,N_14751);
and UO_502 (O_502,N_14528,N_14542);
nand UO_503 (O_503,N_14707,N_14882);
or UO_504 (O_504,N_14887,N_14645);
nand UO_505 (O_505,N_14861,N_14685);
nand UO_506 (O_506,N_14972,N_14853);
xor UO_507 (O_507,N_14865,N_14877);
nand UO_508 (O_508,N_14789,N_14884);
nand UO_509 (O_509,N_14809,N_14797);
and UO_510 (O_510,N_14653,N_14924);
xnor UO_511 (O_511,N_14526,N_14881);
and UO_512 (O_512,N_14755,N_14901);
or UO_513 (O_513,N_14830,N_14659);
nand UO_514 (O_514,N_14858,N_14793);
nor UO_515 (O_515,N_14894,N_14680);
nor UO_516 (O_516,N_14539,N_14560);
and UO_517 (O_517,N_14517,N_14891);
nand UO_518 (O_518,N_14647,N_14513);
nand UO_519 (O_519,N_14562,N_14870);
nand UO_520 (O_520,N_14500,N_14995);
nand UO_521 (O_521,N_14757,N_14947);
or UO_522 (O_522,N_14719,N_14967);
nand UO_523 (O_523,N_14938,N_14895);
or UO_524 (O_524,N_14950,N_14673);
or UO_525 (O_525,N_14680,N_14573);
and UO_526 (O_526,N_14970,N_14815);
nor UO_527 (O_527,N_14925,N_14876);
nand UO_528 (O_528,N_14662,N_14664);
or UO_529 (O_529,N_14570,N_14895);
xor UO_530 (O_530,N_14623,N_14733);
nor UO_531 (O_531,N_14782,N_14879);
nand UO_532 (O_532,N_14910,N_14682);
nand UO_533 (O_533,N_14605,N_14947);
and UO_534 (O_534,N_14981,N_14739);
nand UO_535 (O_535,N_14540,N_14586);
nand UO_536 (O_536,N_14760,N_14521);
nand UO_537 (O_537,N_14698,N_14574);
and UO_538 (O_538,N_14521,N_14935);
nor UO_539 (O_539,N_14796,N_14781);
nor UO_540 (O_540,N_14810,N_14666);
and UO_541 (O_541,N_14584,N_14743);
xnor UO_542 (O_542,N_14668,N_14942);
or UO_543 (O_543,N_14658,N_14623);
and UO_544 (O_544,N_14854,N_14831);
and UO_545 (O_545,N_14742,N_14872);
or UO_546 (O_546,N_14787,N_14694);
xor UO_547 (O_547,N_14873,N_14622);
and UO_548 (O_548,N_14601,N_14898);
nand UO_549 (O_549,N_14933,N_14562);
or UO_550 (O_550,N_14678,N_14520);
or UO_551 (O_551,N_14675,N_14640);
and UO_552 (O_552,N_14941,N_14962);
nor UO_553 (O_553,N_14662,N_14863);
xnor UO_554 (O_554,N_14554,N_14879);
or UO_555 (O_555,N_14751,N_14944);
and UO_556 (O_556,N_14712,N_14615);
nand UO_557 (O_557,N_14698,N_14713);
nand UO_558 (O_558,N_14522,N_14768);
and UO_559 (O_559,N_14693,N_14838);
nor UO_560 (O_560,N_14798,N_14507);
nor UO_561 (O_561,N_14917,N_14817);
or UO_562 (O_562,N_14773,N_14573);
or UO_563 (O_563,N_14865,N_14500);
or UO_564 (O_564,N_14705,N_14963);
xor UO_565 (O_565,N_14662,N_14766);
nor UO_566 (O_566,N_14590,N_14896);
and UO_567 (O_567,N_14784,N_14595);
and UO_568 (O_568,N_14757,N_14573);
nor UO_569 (O_569,N_14605,N_14624);
nand UO_570 (O_570,N_14774,N_14781);
nor UO_571 (O_571,N_14614,N_14722);
xnor UO_572 (O_572,N_14736,N_14523);
and UO_573 (O_573,N_14957,N_14795);
nand UO_574 (O_574,N_14601,N_14759);
nand UO_575 (O_575,N_14728,N_14558);
xor UO_576 (O_576,N_14987,N_14777);
nand UO_577 (O_577,N_14577,N_14781);
or UO_578 (O_578,N_14974,N_14680);
nor UO_579 (O_579,N_14667,N_14533);
nand UO_580 (O_580,N_14661,N_14915);
or UO_581 (O_581,N_14988,N_14711);
nor UO_582 (O_582,N_14583,N_14630);
nand UO_583 (O_583,N_14876,N_14603);
xor UO_584 (O_584,N_14985,N_14586);
or UO_585 (O_585,N_14743,N_14662);
nand UO_586 (O_586,N_14816,N_14864);
nor UO_587 (O_587,N_14898,N_14781);
nand UO_588 (O_588,N_14705,N_14993);
or UO_589 (O_589,N_14887,N_14688);
or UO_590 (O_590,N_14535,N_14626);
nor UO_591 (O_591,N_14704,N_14507);
and UO_592 (O_592,N_14539,N_14808);
or UO_593 (O_593,N_14825,N_14816);
xor UO_594 (O_594,N_14946,N_14534);
or UO_595 (O_595,N_14886,N_14799);
xnor UO_596 (O_596,N_14771,N_14841);
and UO_597 (O_597,N_14788,N_14648);
nor UO_598 (O_598,N_14666,N_14866);
xor UO_599 (O_599,N_14797,N_14847);
nor UO_600 (O_600,N_14589,N_14841);
or UO_601 (O_601,N_14523,N_14841);
nor UO_602 (O_602,N_14971,N_14554);
or UO_603 (O_603,N_14567,N_14696);
nor UO_604 (O_604,N_14697,N_14646);
xor UO_605 (O_605,N_14652,N_14601);
nand UO_606 (O_606,N_14684,N_14530);
or UO_607 (O_607,N_14958,N_14842);
or UO_608 (O_608,N_14944,N_14744);
nand UO_609 (O_609,N_14507,N_14913);
and UO_610 (O_610,N_14941,N_14517);
nand UO_611 (O_611,N_14560,N_14656);
or UO_612 (O_612,N_14768,N_14797);
nor UO_613 (O_613,N_14728,N_14926);
nand UO_614 (O_614,N_14894,N_14638);
and UO_615 (O_615,N_14925,N_14630);
nor UO_616 (O_616,N_14586,N_14973);
or UO_617 (O_617,N_14940,N_14694);
xor UO_618 (O_618,N_14775,N_14939);
nor UO_619 (O_619,N_14531,N_14998);
nand UO_620 (O_620,N_14871,N_14838);
and UO_621 (O_621,N_14989,N_14721);
or UO_622 (O_622,N_14563,N_14704);
and UO_623 (O_623,N_14508,N_14799);
and UO_624 (O_624,N_14565,N_14522);
xnor UO_625 (O_625,N_14594,N_14934);
or UO_626 (O_626,N_14723,N_14655);
nor UO_627 (O_627,N_14599,N_14510);
nand UO_628 (O_628,N_14644,N_14613);
or UO_629 (O_629,N_14911,N_14539);
or UO_630 (O_630,N_14629,N_14586);
nor UO_631 (O_631,N_14640,N_14637);
or UO_632 (O_632,N_14656,N_14703);
or UO_633 (O_633,N_14659,N_14609);
and UO_634 (O_634,N_14735,N_14724);
nor UO_635 (O_635,N_14918,N_14617);
and UO_636 (O_636,N_14572,N_14547);
xor UO_637 (O_637,N_14749,N_14865);
nor UO_638 (O_638,N_14850,N_14618);
and UO_639 (O_639,N_14705,N_14575);
nand UO_640 (O_640,N_14674,N_14807);
xnor UO_641 (O_641,N_14715,N_14588);
nor UO_642 (O_642,N_14748,N_14825);
nor UO_643 (O_643,N_14747,N_14611);
or UO_644 (O_644,N_14569,N_14597);
and UO_645 (O_645,N_14882,N_14905);
or UO_646 (O_646,N_14726,N_14825);
nor UO_647 (O_647,N_14542,N_14910);
or UO_648 (O_648,N_14809,N_14796);
and UO_649 (O_649,N_14825,N_14750);
nand UO_650 (O_650,N_14661,N_14548);
or UO_651 (O_651,N_14645,N_14665);
or UO_652 (O_652,N_14728,N_14678);
and UO_653 (O_653,N_14890,N_14601);
and UO_654 (O_654,N_14725,N_14882);
xnor UO_655 (O_655,N_14833,N_14572);
nand UO_656 (O_656,N_14642,N_14953);
nand UO_657 (O_657,N_14857,N_14519);
nand UO_658 (O_658,N_14722,N_14741);
nor UO_659 (O_659,N_14799,N_14997);
or UO_660 (O_660,N_14844,N_14567);
and UO_661 (O_661,N_14840,N_14654);
or UO_662 (O_662,N_14545,N_14942);
xor UO_663 (O_663,N_14613,N_14997);
or UO_664 (O_664,N_14560,N_14968);
nor UO_665 (O_665,N_14515,N_14831);
and UO_666 (O_666,N_14779,N_14687);
xnor UO_667 (O_667,N_14845,N_14939);
xnor UO_668 (O_668,N_14517,N_14843);
xor UO_669 (O_669,N_14635,N_14742);
or UO_670 (O_670,N_14687,N_14550);
and UO_671 (O_671,N_14893,N_14752);
and UO_672 (O_672,N_14614,N_14760);
nor UO_673 (O_673,N_14661,N_14651);
and UO_674 (O_674,N_14948,N_14818);
nand UO_675 (O_675,N_14696,N_14791);
xor UO_676 (O_676,N_14987,N_14789);
xnor UO_677 (O_677,N_14926,N_14756);
or UO_678 (O_678,N_14672,N_14899);
and UO_679 (O_679,N_14993,N_14650);
nand UO_680 (O_680,N_14979,N_14952);
nor UO_681 (O_681,N_14932,N_14550);
nor UO_682 (O_682,N_14591,N_14988);
and UO_683 (O_683,N_14644,N_14684);
and UO_684 (O_684,N_14850,N_14700);
nand UO_685 (O_685,N_14981,N_14755);
xnor UO_686 (O_686,N_14760,N_14531);
and UO_687 (O_687,N_14967,N_14615);
xor UO_688 (O_688,N_14510,N_14801);
and UO_689 (O_689,N_14619,N_14555);
nand UO_690 (O_690,N_14990,N_14632);
xnor UO_691 (O_691,N_14759,N_14938);
or UO_692 (O_692,N_14599,N_14746);
or UO_693 (O_693,N_14561,N_14564);
or UO_694 (O_694,N_14534,N_14824);
or UO_695 (O_695,N_14765,N_14595);
nor UO_696 (O_696,N_14876,N_14907);
nor UO_697 (O_697,N_14911,N_14541);
and UO_698 (O_698,N_14665,N_14675);
nor UO_699 (O_699,N_14770,N_14547);
nor UO_700 (O_700,N_14996,N_14511);
or UO_701 (O_701,N_14633,N_14824);
nand UO_702 (O_702,N_14747,N_14540);
and UO_703 (O_703,N_14685,N_14835);
xnor UO_704 (O_704,N_14560,N_14727);
nand UO_705 (O_705,N_14820,N_14943);
or UO_706 (O_706,N_14616,N_14826);
nand UO_707 (O_707,N_14812,N_14814);
nor UO_708 (O_708,N_14718,N_14719);
xor UO_709 (O_709,N_14693,N_14906);
and UO_710 (O_710,N_14573,N_14783);
nor UO_711 (O_711,N_14942,N_14644);
and UO_712 (O_712,N_14612,N_14529);
nor UO_713 (O_713,N_14592,N_14963);
or UO_714 (O_714,N_14715,N_14584);
nand UO_715 (O_715,N_14772,N_14996);
xnor UO_716 (O_716,N_14978,N_14693);
nor UO_717 (O_717,N_14900,N_14754);
or UO_718 (O_718,N_14976,N_14966);
or UO_719 (O_719,N_14661,N_14578);
nor UO_720 (O_720,N_14965,N_14514);
nor UO_721 (O_721,N_14943,N_14579);
and UO_722 (O_722,N_14695,N_14760);
nor UO_723 (O_723,N_14732,N_14531);
or UO_724 (O_724,N_14590,N_14650);
and UO_725 (O_725,N_14793,N_14649);
nand UO_726 (O_726,N_14797,N_14563);
and UO_727 (O_727,N_14688,N_14698);
or UO_728 (O_728,N_14948,N_14536);
and UO_729 (O_729,N_14970,N_14844);
xor UO_730 (O_730,N_14798,N_14751);
or UO_731 (O_731,N_14662,N_14939);
nor UO_732 (O_732,N_14810,N_14882);
nand UO_733 (O_733,N_14558,N_14876);
or UO_734 (O_734,N_14528,N_14918);
nand UO_735 (O_735,N_14993,N_14812);
and UO_736 (O_736,N_14504,N_14679);
nor UO_737 (O_737,N_14590,N_14632);
or UO_738 (O_738,N_14505,N_14838);
nor UO_739 (O_739,N_14659,N_14799);
nor UO_740 (O_740,N_14594,N_14764);
nand UO_741 (O_741,N_14543,N_14622);
or UO_742 (O_742,N_14604,N_14803);
xor UO_743 (O_743,N_14713,N_14592);
and UO_744 (O_744,N_14796,N_14891);
nand UO_745 (O_745,N_14545,N_14674);
or UO_746 (O_746,N_14603,N_14877);
or UO_747 (O_747,N_14740,N_14543);
xor UO_748 (O_748,N_14700,N_14680);
or UO_749 (O_749,N_14982,N_14589);
xnor UO_750 (O_750,N_14612,N_14561);
or UO_751 (O_751,N_14909,N_14813);
xor UO_752 (O_752,N_14648,N_14893);
nor UO_753 (O_753,N_14748,N_14874);
xnor UO_754 (O_754,N_14950,N_14764);
nand UO_755 (O_755,N_14739,N_14621);
xor UO_756 (O_756,N_14865,N_14979);
xnor UO_757 (O_757,N_14647,N_14810);
nand UO_758 (O_758,N_14885,N_14743);
and UO_759 (O_759,N_14755,N_14874);
nand UO_760 (O_760,N_14907,N_14971);
nand UO_761 (O_761,N_14830,N_14655);
xor UO_762 (O_762,N_14915,N_14816);
nand UO_763 (O_763,N_14792,N_14747);
and UO_764 (O_764,N_14545,N_14665);
nand UO_765 (O_765,N_14990,N_14795);
and UO_766 (O_766,N_14561,N_14835);
nor UO_767 (O_767,N_14549,N_14833);
or UO_768 (O_768,N_14829,N_14592);
nor UO_769 (O_769,N_14799,N_14752);
and UO_770 (O_770,N_14660,N_14940);
nand UO_771 (O_771,N_14677,N_14801);
xnor UO_772 (O_772,N_14583,N_14785);
nor UO_773 (O_773,N_14971,N_14535);
nor UO_774 (O_774,N_14991,N_14946);
or UO_775 (O_775,N_14645,N_14854);
or UO_776 (O_776,N_14599,N_14849);
nor UO_777 (O_777,N_14606,N_14707);
or UO_778 (O_778,N_14527,N_14699);
and UO_779 (O_779,N_14645,N_14538);
or UO_780 (O_780,N_14623,N_14543);
and UO_781 (O_781,N_14996,N_14741);
and UO_782 (O_782,N_14528,N_14601);
nor UO_783 (O_783,N_14909,N_14660);
or UO_784 (O_784,N_14747,N_14692);
xor UO_785 (O_785,N_14778,N_14563);
nor UO_786 (O_786,N_14764,N_14947);
nand UO_787 (O_787,N_14618,N_14788);
nor UO_788 (O_788,N_14942,N_14557);
or UO_789 (O_789,N_14578,N_14942);
and UO_790 (O_790,N_14818,N_14530);
nor UO_791 (O_791,N_14730,N_14919);
nor UO_792 (O_792,N_14750,N_14955);
nand UO_793 (O_793,N_14544,N_14768);
or UO_794 (O_794,N_14551,N_14744);
or UO_795 (O_795,N_14509,N_14840);
xnor UO_796 (O_796,N_14521,N_14548);
and UO_797 (O_797,N_14917,N_14524);
and UO_798 (O_798,N_14817,N_14639);
and UO_799 (O_799,N_14852,N_14690);
xnor UO_800 (O_800,N_14727,N_14718);
and UO_801 (O_801,N_14500,N_14573);
or UO_802 (O_802,N_14834,N_14601);
and UO_803 (O_803,N_14513,N_14990);
xnor UO_804 (O_804,N_14726,N_14554);
and UO_805 (O_805,N_14596,N_14650);
xor UO_806 (O_806,N_14830,N_14750);
xor UO_807 (O_807,N_14649,N_14774);
xnor UO_808 (O_808,N_14788,N_14720);
nor UO_809 (O_809,N_14734,N_14668);
nor UO_810 (O_810,N_14834,N_14790);
and UO_811 (O_811,N_14593,N_14877);
nor UO_812 (O_812,N_14660,N_14634);
nor UO_813 (O_813,N_14894,N_14877);
nand UO_814 (O_814,N_14538,N_14747);
and UO_815 (O_815,N_14553,N_14743);
nand UO_816 (O_816,N_14718,N_14922);
nor UO_817 (O_817,N_14579,N_14830);
nand UO_818 (O_818,N_14860,N_14944);
or UO_819 (O_819,N_14936,N_14718);
xnor UO_820 (O_820,N_14765,N_14674);
xnor UO_821 (O_821,N_14546,N_14651);
nand UO_822 (O_822,N_14608,N_14835);
nor UO_823 (O_823,N_14874,N_14593);
xor UO_824 (O_824,N_14616,N_14698);
and UO_825 (O_825,N_14689,N_14521);
or UO_826 (O_826,N_14583,N_14814);
nor UO_827 (O_827,N_14906,N_14732);
xnor UO_828 (O_828,N_14739,N_14707);
nand UO_829 (O_829,N_14628,N_14779);
nor UO_830 (O_830,N_14889,N_14887);
xor UO_831 (O_831,N_14627,N_14774);
nor UO_832 (O_832,N_14715,N_14723);
xor UO_833 (O_833,N_14828,N_14647);
or UO_834 (O_834,N_14798,N_14881);
nor UO_835 (O_835,N_14582,N_14782);
nor UO_836 (O_836,N_14858,N_14559);
or UO_837 (O_837,N_14569,N_14766);
or UO_838 (O_838,N_14906,N_14787);
nand UO_839 (O_839,N_14926,N_14720);
xor UO_840 (O_840,N_14756,N_14649);
or UO_841 (O_841,N_14751,N_14611);
xor UO_842 (O_842,N_14723,N_14919);
nor UO_843 (O_843,N_14815,N_14963);
nor UO_844 (O_844,N_14956,N_14600);
and UO_845 (O_845,N_14763,N_14632);
and UO_846 (O_846,N_14710,N_14961);
nor UO_847 (O_847,N_14826,N_14995);
or UO_848 (O_848,N_14654,N_14500);
or UO_849 (O_849,N_14627,N_14903);
nor UO_850 (O_850,N_14564,N_14757);
xor UO_851 (O_851,N_14648,N_14566);
nor UO_852 (O_852,N_14545,N_14549);
xnor UO_853 (O_853,N_14624,N_14518);
nor UO_854 (O_854,N_14926,N_14962);
or UO_855 (O_855,N_14664,N_14551);
and UO_856 (O_856,N_14923,N_14694);
nor UO_857 (O_857,N_14633,N_14876);
and UO_858 (O_858,N_14679,N_14759);
nand UO_859 (O_859,N_14574,N_14537);
or UO_860 (O_860,N_14663,N_14656);
or UO_861 (O_861,N_14828,N_14916);
nand UO_862 (O_862,N_14820,N_14911);
nand UO_863 (O_863,N_14963,N_14804);
and UO_864 (O_864,N_14718,N_14780);
and UO_865 (O_865,N_14859,N_14790);
xor UO_866 (O_866,N_14538,N_14719);
nand UO_867 (O_867,N_14781,N_14591);
and UO_868 (O_868,N_14636,N_14997);
or UO_869 (O_869,N_14982,N_14705);
or UO_870 (O_870,N_14996,N_14918);
nand UO_871 (O_871,N_14664,N_14754);
and UO_872 (O_872,N_14974,N_14756);
and UO_873 (O_873,N_14576,N_14977);
xor UO_874 (O_874,N_14803,N_14800);
xnor UO_875 (O_875,N_14959,N_14766);
or UO_876 (O_876,N_14720,N_14831);
xnor UO_877 (O_877,N_14855,N_14742);
nand UO_878 (O_878,N_14829,N_14609);
nor UO_879 (O_879,N_14718,N_14960);
nor UO_880 (O_880,N_14589,N_14542);
xor UO_881 (O_881,N_14956,N_14891);
xor UO_882 (O_882,N_14527,N_14952);
nor UO_883 (O_883,N_14519,N_14706);
and UO_884 (O_884,N_14775,N_14592);
nor UO_885 (O_885,N_14945,N_14753);
nor UO_886 (O_886,N_14979,N_14684);
nor UO_887 (O_887,N_14893,N_14867);
nand UO_888 (O_888,N_14691,N_14980);
and UO_889 (O_889,N_14702,N_14711);
nor UO_890 (O_890,N_14984,N_14954);
or UO_891 (O_891,N_14804,N_14826);
nand UO_892 (O_892,N_14536,N_14940);
and UO_893 (O_893,N_14909,N_14559);
nor UO_894 (O_894,N_14501,N_14909);
and UO_895 (O_895,N_14884,N_14935);
and UO_896 (O_896,N_14839,N_14565);
nor UO_897 (O_897,N_14586,N_14751);
nand UO_898 (O_898,N_14983,N_14763);
and UO_899 (O_899,N_14731,N_14927);
nand UO_900 (O_900,N_14713,N_14522);
and UO_901 (O_901,N_14859,N_14912);
nor UO_902 (O_902,N_14650,N_14992);
or UO_903 (O_903,N_14827,N_14529);
and UO_904 (O_904,N_14849,N_14566);
xor UO_905 (O_905,N_14610,N_14530);
and UO_906 (O_906,N_14982,N_14935);
or UO_907 (O_907,N_14692,N_14878);
nand UO_908 (O_908,N_14863,N_14868);
nor UO_909 (O_909,N_14961,N_14891);
nor UO_910 (O_910,N_14966,N_14919);
or UO_911 (O_911,N_14571,N_14806);
and UO_912 (O_912,N_14610,N_14934);
nor UO_913 (O_913,N_14758,N_14695);
xnor UO_914 (O_914,N_14859,N_14915);
nor UO_915 (O_915,N_14883,N_14504);
nor UO_916 (O_916,N_14810,N_14988);
xnor UO_917 (O_917,N_14861,N_14857);
and UO_918 (O_918,N_14883,N_14869);
and UO_919 (O_919,N_14537,N_14794);
nor UO_920 (O_920,N_14790,N_14890);
nand UO_921 (O_921,N_14784,N_14890);
and UO_922 (O_922,N_14653,N_14995);
nand UO_923 (O_923,N_14618,N_14507);
xor UO_924 (O_924,N_14868,N_14884);
nor UO_925 (O_925,N_14898,N_14566);
or UO_926 (O_926,N_14732,N_14625);
or UO_927 (O_927,N_14922,N_14931);
or UO_928 (O_928,N_14803,N_14658);
nor UO_929 (O_929,N_14514,N_14608);
and UO_930 (O_930,N_14837,N_14761);
or UO_931 (O_931,N_14976,N_14592);
xnor UO_932 (O_932,N_14751,N_14524);
or UO_933 (O_933,N_14971,N_14888);
or UO_934 (O_934,N_14763,N_14899);
xor UO_935 (O_935,N_14597,N_14646);
and UO_936 (O_936,N_14843,N_14686);
xnor UO_937 (O_937,N_14558,N_14752);
xor UO_938 (O_938,N_14763,N_14878);
or UO_939 (O_939,N_14563,N_14911);
xnor UO_940 (O_940,N_14739,N_14559);
nor UO_941 (O_941,N_14823,N_14895);
nand UO_942 (O_942,N_14727,N_14687);
or UO_943 (O_943,N_14617,N_14888);
or UO_944 (O_944,N_14544,N_14633);
or UO_945 (O_945,N_14728,N_14664);
nand UO_946 (O_946,N_14500,N_14868);
nand UO_947 (O_947,N_14707,N_14924);
or UO_948 (O_948,N_14968,N_14977);
and UO_949 (O_949,N_14908,N_14540);
or UO_950 (O_950,N_14514,N_14606);
nand UO_951 (O_951,N_14717,N_14622);
and UO_952 (O_952,N_14576,N_14849);
xor UO_953 (O_953,N_14742,N_14687);
nor UO_954 (O_954,N_14665,N_14673);
nor UO_955 (O_955,N_14770,N_14722);
nand UO_956 (O_956,N_14709,N_14698);
and UO_957 (O_957,N_14568,N_14514);
or UO_958 (O_958,N_14575,N_14552);
nand UO_959 (O_959,N_14679,N_14661);
or UO_960 (O_960,N_14796,N_14543);
xnor UO_961 (O_961,N_14855,N_14919);
or UO_962 (O_962,N_14567,N_14523);
nor UO_963 (O_963,N_14608,N_14893);
nor UO_964 (O_964,N_14960,N_14812);
and UO_965 (O_965,N_14598,N_14721);
nand UO_966 (O_966,N_14560,N_14515);
nand UO_967 (O_967,N_14798,N_14554);
and UO_968 (O_968,N_14948,N_14886);
nor UO_969 (O_969,N_14655,N_14508);
or UO_970 (O_970,N_14855,N_14587);
nor UO_971 (O_971,N_14533,N_14767);
or UO_972 (O_972,N_14733,N_14550);
xor UO_973 (O_973,N_14803,N_14869);
or UO_974 (O_974,N_14808,N_14666);
or UO_975 (O_975,N_14923,N_14680);
xor UO_976 (O_976,N_14807,N_14606);
xor UO_977 (O_977,N_14784,N_14571);
and UO_978 (O_978,N_14818,N_14955);
or UO_979 (O_979,N_14643,N_14965);
nand UO_980 (O_980,N_14624,N_14533);
and UO_981 (O_981,N_14661,N_14633);
nor UO_982 (O_982,N_14770,N_14805);
nand UO_983 (O_983,N_14861,N_14900);
or UO_984 (O_984,N_14718,N_14854);
and UO_985 (O_985,N_14556,N_14874);
nor UO_986 (O_986,N_14503,N_14739);
xnor UO_987 (O_987,N_14849,N_14649);
nand UO_988 (O_988,N_14941,N_14662);
xor UO_989 (O_989,N_14521,N_14569);
and UO_990 (O_990,N_14855,N_14668);
and UO_991 (O_991,N_14904,N_14513);
nor UO_992 (O_992,N_14724,N_14885);
or UO_993 (O_993,N_14643,N_14902);
nand UO_994 (O_994,N_14690,N_14877);
and UO_995 (O_995,N_14716,N_14683);
nor UO_996 (O_996,N_14851,N_14665);
and UO_997 (O_997,N_14835,N_14735);
nand UO_998 (O_998,N_14954,N_14751);
nor UO_999 (O_999,N_14704,N_14631);
nand UO_1000 (O_1000,N_14709,N_14809);
or UO_1001 (O_1001,N_14640,N_14824);
nor UO_1002 (O_1002,N_14512,N_14571);
nand UO_1003 (O_1003,N_14941,N_14719);
and UO_1004 (O_1004,N_14525,N_14882);
and UO_1005 (O_1005,N_14687,N_14603);
and UO_1006 (O_1006,N_14901,N_14953);
and UO_1007 (O_1007,N_14568,N_14675);
xnor UO_1008 (O_1008,N_14757,N_14515);
nor UO_1009 (O_1009,N_14590,N_14624);
nor UO_1010 (O_1010,N_14587,N_14937);
nor UO_1011 (O_1011,N_14948,N_14640);
or UO_1012 (O_1012,N_14901,N_14511);
or UO_1013 (O_1013,N_14767,N_14658);
and UO_1014 (O_1014,N_14691,N_14824);
xor UO_1015 (O_1015,N_14532,N_14850);
and UO_1016 (O_1016,N_14833,N_14560);
nor UO_1017 (O_1017,N_14654,N_14871);
nor UO_1018 (O_1018,N_14857,N_14568);
or UO_1019 (O_1019,N_14686,N_14873);
nor UO_1020 (O_1020,N_14924,N_14553);
and UO_1021 (O_1021,N_14868,N_14567);
nand UO_1022 (O_1022,N_14837,N_14993);
nand UO_1023 (O_1023,N_14612,N_14703);
and UO_1024 (O_1024,N_14570,N_14941);
or UO_1025 (O_1025,N_14552,N_14682);
xor UO_1026 (O_1026,N_14522,N_14873);
or UO_1027 (O_1027,N_14713,N_14865);
and UO_1028 (O_1028,N_14681,N_14500);
or UO_1029 (O_1029,N_14576,N_14737);
or UO_1030 (O_1030,N_14561,N_14801);
nand UO_1031 (O_1031,N_14927,N_14749);
nor UO_1032 (O_1032,N_14526,N_14634);
or UO_1033 (O_1033,N_14876,N_14905);
or UO_1034 (O_1034,N_14683,N_14809);
xor UO_1035 (O_1035,N_14839,N_14741);
nand UO_1036 (O_1036,N_14687,N_14685);
or UO_1037 (O_1037,N_14755,N_14985);
nor UO_1038 (O_1038,N_14767,N_14963);
nor UO_1039 (O_1039,N_14752,N_14845);
xor UO_1040 (O_1040,N_14715,N_14933);
or UO_1041 (O_1041,N_14698,N_14850);
xnor UO_1042 (O_1042,N_14852,N_14812);
nor UO_1043 (O_1043,N_14654,N_14999);
and UO_1044 (O_1044,N_14590,N_14766);
xor UO_1045 (O_1045,N_14736,N_14971);
and UO_1046 (O_1046,N_14529,N_14570);
nand UO_1047 (O_1047,N_14980,N_14714);
or UO_1048 (O_1048,N_14608,N_14775);
nand UO_1049 (O_1049,N_14779,N_14594);
and UO_1050 (O_1050,N_14652,N_14721);
and UO_1051 (O_1051,N_14598,N_14797);
and UO_1052 (O_1052,N_14902,N_14970);
xor UO_1053 (O_1053,N_14807,N_14501);
nor UO_1054 (O_1054,N_14502,N_14730);
or UO_1055 (O_1055,N_14963,N_14663);
nor UO_1056 (O_1056,N_14685,N_14553);
and UO_1057 (O_1057,N_14886,N_14665);
or UO_1058 (O_1058,N_14558,N_14802);
xor UO_1059 (O_1059,N_14519,N_14883);
nor UO_1060 (O_1060,N_14522,N_14849);
and UO_1061 (O_1061,N_14900,N_14937);
and UO_1062 (O_1062,N_14616,N_14638);
and UO_1063 (O_1063,N_14802,N_14705);
nand UO_1064 (O_1064,N_14638,N_14589);
xor UO_1065 (O_1065,N_14829,N_14651);
and UO_1066 (O_1066,N_14918,N_14815);
nand UO_1067 (O_1067,N_14807,N_14899);
nor UO_1068 (O_1068,N_14607,N_14759);
xnor UO_1069 (O_1069,N_14548,N_14882);
or UO_1070 (O_1070,N_14648,N_14543);
nand UO_1071 (O_1071,N_14769,N_14678);
or UO_1072 (O_1072,N_14642,N_14949);
or UO_1073 (O_1073,N_14615,N_14718);
nor UO_1074 (O_1074,N_14745,N_14561);
or UO_1075 (O_1075,N_14750,N_14935);
or UO_1076 (O_1076,N_14515,N_14702);
nand UO_1077 (O_1077,N_14672,N_14634);
nand UO_1078 (O_1078,N_14634,N_14806);
nand UO_1079 (O_1079,N_14987,N_14521);
nor UO_1080 (O_1080,N_14584,N_14915);
nand UO_1081 (O_1081,N_14874,N_14940);
and UO_1082 (O_1082,N_14819,N_14809);
xor UO_1083 (O_1083,N_14892,N_14839);
xor UO_1084 (O_1084,N_14756,N_14657);
or UO_1085 (O_1085,N_14677,N_14817);
and UO_1086 (O_1086,N_14522,N_14848);
nor UO_1087 (O_1087,N_14671,N_14521);
nand UO_1088 (O_1088,N_14865,N_14858);
xor UO_1089 (O_1089,N_14535,N_14603);
nand UO_1090 (O_1090,N_14787,N_14734);
and UO_1091 (O_1091,N_14773,N_14933);
xor UO_1092 (O_1092,N_14512,N_14726);
or UO_1093 (O_1093,N_14964,N_14935);
xor UO_1094 (O_1094,N_14932,N_14527);
nand UO_1095 (O_1095,N_14516,N_14592);
and UO_1096 (O_1096,N_14755,N_14561);
or UO_1097 (O_1097,N_14895,N_14896);
xor UO_1098 (O_1098,N_14738,N_14777);
or UO_1099 (O_1099,N_14668,N_14599);
nor UO_1100 (O_1100,N_14628,N_14742);
nor UO_1101 (O_1101,N_14503,N_14858);
xor UO_1102 (O_1102,N_14574,N_14823);
nand UO_1103 (O_1103,N_14658,N_14877);
nor UO_1104 (O_1104,N_14514,N_14689);
nand UO_1105 (O_1105,N_14575,N_14510);
xnor UO_1106 (O_1106,N_14539,N_14688);
nand UO_1107 (O_1107,N_14697,N_14990);
nor UO_1108 (O_1108,N_14991,N_14762);
nor UO_1109 (O_1109,N_14571,N_14692);
nand UO_1110 (O_1110,N_14905,N_14989);
nand UO_1111 (O_1111,N_14550,N_14965);
nor UO_1112 (O_1112,N_14911,N_14977);
and UO_1113 (O_1113,N_14509,N_14577);
nand UO_1114 (O_1114,N_14956,N_14663);
nor UO_1115 (O_1115,N_14927,N_14809);
nand UO_1116 (O_1116,N_14501,N_14517);
nand UO_1117 (O_1117,N_14775,N_14531);
and UO_1118 (O_1118,N_14829,N_14917);
and UO_1119 (O_1119,N_14739,N_14856);
xor UO_1120 (O_1120,N_14707,N_14826);
nor UO_1121 (O_1121,N_14841,N_14738);
nand UO_1122 (O_1122,N_14713,N_14869);
or UO_1123 (O_1123,N_14884,N_14942);
and UO_1124 (O_1124,N_14627,N_14652);
nor UO_1125 (O_1125,N_14877,N_14837);
xnor UO_1126 (O_1126,N_14548,N_14620);
nor UO_1127 (O_1127,N_14532,N_14915);
or UO_1128 (O_1128,N_14885,N_14572);
xor UO_1129 (O_1129,N_14883,N_14607);
xor UO_1130 (O_1130,N_14925,N_14649);
xnor UO_1131 (O_1131,N_14851,N_14552);
or UO_1132 (O_1132,N_14534,N_14697);
xnor UO_1133 (O_1133,N_14843,N_14510);
nand UO_1134 (O_1134,N_14680,N_14501);
nand UO_1135 (O_1135,N_14993,N_14697);
xnor UO_1136 (O_1136,N_14995,N_14947);
and UO_1137 (O_1137,N_14921,N_14946);
or UO_1138 (O_1138,N_14810,N_14640);
or UO_1139 (O_1139,N_14738,N_14690);
nand UO_1140 (O_1140,N_14946,N_14795);
or UO_1141 (O_1141,N_14791,N_14673);
or UO_1142 (O_1142,N_14973,N_14756);
nand UO_1143 (O_1143,N_14833,N_14678);
nand UO_1144 (O_1144,N_14768,N_14605);
or UO_1145 (O_1145,N_14527,N_14794);
nor UO_1146 (O_1146,N_14889,N_14823);
nand UO_1147 (O_1147,N_14674,N_14998);
or UO_1148 (O_1148,N_14652,N_14687);
nand UO_1149 (O_1149,N_14729,N_14575);
or UO_1150 (O_1150,N_14822,N_14808);
nand UO_1151 (O_1151,N_14780,N_14631);
nor UO_1152 (O_1152,N_14756,N_14776);
and UO_1153 (O_1153,N_14617,N_14743);
or UO_1154 (O_1154,N_14566,N_14807);
nor UO_1155 (O_1155,N_14691,N_14839);
and UO_1156 (O_1156,N_14873,N_14691);
nand UO_1157 (O_1157,N_14603,N_14802);
nor UO_1158 (O_1158,N_14559,N_14821);
nand UO_1159 (O_1159,N_14501,N_14657);
nand UO_1160 (O_1160,N_14713,N_14921);
nand UO_1161 (O_1161,N_14570,N_14544);
nor UO_1162 (O_1162,N_14954,N_14572);
and UO_1163 (O_1163,N_14648,N_14519);
xnor UO_1164 (O_1164,N_14541,N_14589);
nor UO_1165 (O_1165,N_14518,N_14921);
nor UO_1166 (O_1166,N_14626,N_14719);
nand UO_1167 (O_1167,N_14642,N_14664);
and UO_1168 (O_1168,N_14728,N_14634);
nand UO_1169 (O_1169,N_14927,N_14590);
xor UO_1170 (O_1170,N_14739,N_14909);
xnor UO_1171 (O_1171,N_14898,N_14754);
xor UO_1172 (O_1172,N_14805,N_14533);
and UO_1173 (O_1173,N_14925,N_14629);
and UO_1174 (O_1174,N_14534,N_14570);
nor UO_1175 (O_1175,N_14921,N_14532);
nor UO_1176 (O_1176,N_14699,N_14604);
nand UO_1177 (O_1177,N_14900,N_14926);
nor UO_1178 (O_1178,N_14801,N_14884);
or UO_1179 (O_1179,N_14819,N_14554);
or UO_1180 (O_1180,N_14708,N_14641);
and UO_1181 (O_1181,N_14894,N_14901);
xnor UO_1182 (O_1182,N_14835,N_14796);
and UO_1183 (O_1183,N_14667,N_14976);
and UO_1184 (O_1184,N_14961,N_14742);
nand UO_1185 (O_1185,N_14595,N_14589);
or UO_1186 (O_1186,N_14603,N_14544);
xor UO_1187 (O_1187,N_14745,N_14749);
and UO_1188 (O_1188,N_14591,N_14809);
nor UO_1189 (O_1189,N_14539,N_14633);
nor UO_1190 (O_1190,N_14955,N_14953);
xor UO_1191 (O_1191,N_14816,N_14698);
or UO_1192 (O_1192,N_14795,N_14892);
or UO_1193 (O_1193,N_14718,N_14503);
or UO_1194 (O_1194,N_14916,N_14742);
nor UO_1195 (O_1195,N_14936,N_14906);
xnor UO_1196 (O_1196,N_14799,N_14986);
and UO_1197 (O_1197,N_14990,N_14723);
or UO_1198 (O_1198,N_14997,N_14714);
and UO_1199 (O_1199,N_14915,N_14677);
nor UO_1200 (O_1200,N_14943,N_14890);
nor UO_1201 (O_1201,N_14874,N_14689);
and UO_1202 (O_1202,N_14760,N_14803);
nand UO_1203 (O_1203,N_14713,N_14646);
or UO_1204 (O_1204,N_14577,N_14870);
or UO_1205 (O_1205,N_14967,N_14520);
and UO_1206 (O_1206,N_14740,N_14575);
and UO_1207 (O_1207,N_14732,N_14931);
and UO_1208 (O_1208,N_14599,N_14819);
or UO_1209 (O_1209,N_14872,N_14686);
xor UO_1210 (O_1210,N_14505,N_14667);
nor UO_1211 (O_1211,N_14597,N_14823);
xnor UO_1212 (O_1212,N_14965,N_14767);
and UO_1213 (O_1213,N_14919,N_14780);
nand UO_1214 (O_1214,N_14597,N_14564);
xnor UO_1215 (O_1215,N_14953,N_14726);
and UO_1216 (O_1216,N_14878,N_14860);
or UO_1217 (O_1217,N_14703,N_14560);
nor UO_1218 (O_1218,N_14911,N_14710);
nor UO_1219 (O_1219,N_14662,N_14906);
xor UO_1220 (O_1220,N_14934,N_14507);
xnor UO_1221 (O_1221,N_14500,N_14589);
or UO_1222 (O_1222,N_14718,N_14812);
nand UO_1223 (O_1223,N_14786,N_14603);
nor UO_1224 (O_1224,N_14846,N_14606);
nor UO_1225 (O_1225,N_14930,N_14985);
nor UO_1226 (O_1226,N_14820,N_14805);
nand UO_1227 (O_1227,N_14965,N_14691);
xor UO_1228 (O_1228,N_14732,N_14621);
xnor UO_1229 (O_1229,N_14575,N_14975);
nand UO_1230 (O_1230,N_14715,N_14550);
and UO_1231 (O_1231,N_14840,N_14860);
xnor UO_1232 (O_1232,N_14837,N_14960);
or UO_1233 (O_1233,N_14886,N_14965);
nand UO_1234 (O_1234,N_14896,N_14720);
or UO_1235 (O_1235,N_14678,N_14595);
and UO_1236 (O_1236,N_14657,N_14800);
nand UO_1237 (O_1237,N_14596,N_14899);
nor UO_1238 (O_1238,N_14551,N_14916);
and UO_1239 (O_1239,N_14552,N_14871);
xor UO_1240 (O_1240,N_14860,N_14600);
or UO_1241 (O_1241,N_14745,N_14923);
nand UO_1242 (O_1242,N_14717,N_14955);
xor UO_1243 (O_1243,N_14651,N_14919);
and UO_1244 (O_1244,N_14731,N_14615);
nand UO_1245 (O_1245,N_14846,N_14868);
nor UO_1246 (O_1246,N_14867,N_14580);
and UO_1247 (O_1247,N_14840,N_14613);
xnor UO_1248 (O_1248,N_14901,N_14691);
nand UO_1249 (O_1249,N_14924,N_14764);
nor UO_1250 (O_1250,N_14972,N_14747);
or UO_1251 (O_1251,N_14986,N_14926);
or UO_1252 (O_1252,N_14555,N_14920);
nor UO_1253 (O_1253,N_14804,N_14923);
xor UO_1254 (O_1254,N_14894,N_14974);
or UO_1255 (O_1255,N_14830,N_14647);
nand UO_1256 (O_1256,N_14965,N_14524);
and UO_1257 (O_1257,N_14626,N_14596);
nand UO_1258 (O_1258,N_14881,N_14589);
or UO_1259 (O_1259,N_14810,N_14961);
nor UO_1260 (O_1260,N_14999,N_14545);
nor UO_1261 (O_1261,N_14843,N_14771);
or UO_1262 (O_1262,N_14823,N_14511);
or UO_1263 (O_1263,N_14688,N_14825);
xor UO_1264 (O_1264,N_14892,N_14631);
nor UO_1265 (O_1265,N_14704,N_14671);
nand UO_1266 (O_1266,N_14723,N_14696);
nand UO_1267 (O_1267,N_14948,N_14974);
nor UO_1268 (O_1268,N_14807,N_14805);
xor UO_1269 (O_1269,N_14811,N_14835);
or UO_1270 (O_1270,N_14748,N_14683);
nand UO_1271 (O_1271,N_14770,N_14675);
nand UO_1272 (O_1272,N_14596,N_14672);
or UO_1273 (O_1273,N_14975,N_14711);
xnor UO_1274 (O_1274,N_14749,N_14917);
xnor UO_1275 (O_1275,N_14914,N_14925);
and UO_1276 (O_1276,N_14945,N_14507);
xor UO_1277 (O_1277,N_14571,N_14738);
nand UO_1278 (O_1278,N_14759,N_14694);
nand UO_1279 (O_1279,N_14519,N_14656);
and UO_1280 (O_1280,N_14528,N_14566);
nor UO_1281 (O_1281,N_14793,N_14659);
or UO_1282 (O_1282,N_14656,N_14698);
and UO_1283 (O_1283,N_14777,N_14585);
and UO_1284 (O_1284,N_14981,N_14608);
xor UO_1285 (O_1285,N_14810,N_14864);
nand UO_1286 (O_1286,N_14829,N_14652);
xor UO_1287 (O_1287,N_14698,N_14718);
nor UO_1288 (O_1288,N_14841,N_14527);
or UO_1289 (O_1289,N_14962,N_14570);
nor UO_1290 (O_1290,N_14983,N_14594);
or UO_1291 (O_1291,N_14517,N_14898);
nand UO_1292 (O_1292,N_14963,N_14648);
xnor UO_1293 (O_1293,N_14779,N_14707);
and UO_1294 (O_1294,N_14874,N_14885);
and UO_1295 (O_1295,N_14959,N_14560);
and UO_1296 (O_1296,N_14607,N_14786);
nor UO_1297 (O_1297,N_14888,N_14923);
xor UO_1298 (O_1298,N_14993,N_14688);
xor UO_1299 (O_1299,N_14642,N_14994);
xnor UO_1300 (O_1300,N_14998,N_14680);
or UO_1301 (O_1301,N_14544,N_14729);
nor UO_1302 (O_1302,N_14697,N_14660);
xnor UO_1303 (O_1303,N_14900,N_14510);
nand UO_1304 (O_1304,N_14807,N_14909);
xnor UO_1305 (O_1305,N_14728,N_14836);
and UO_1306 (O_1306,N_14532,N_14750);
xnor UO_1307 (O_1307,N_14951,N_14755);
xor UO_1308 (O_1308,N_14795,N_14902);
and UO_1309 (O_1309,N_14592,N_14873);
nand UO_1310 (O_1310,N_14569,N_14613);
xor UO_1311 (O_1311,N_14512,N_14654);
and UO_1312 (O_1312,N_14675,N_14549);
and UO_1313 (O_1313,N_14681,N_14592);
xnor UO_1314 (O_1314,N_14972,N_14745);
xnor UO_1315 (O_1315,N_14682,N_14975);
nor UO_1316 (O_1316,N_14514,N_14776);
xor UO_1317 (O_1317,N_14782,N_14859);
or UO_1318 (O_1318,N_14995,N_14503);
xnor UO_1319 (O_1319,N_14532,N_14647);
and UO_1320 (O_1320,N_14591,N_14910);
and UO_1321 (O_1321,N_14838,N_14884);
nor UO_1322 (O_1322,N_14562,N_14813);
xnor UO_1323 (O_1323,N_14896,N_14938);
or UO_1324 (O_1324,N_14700,N_14815);
nor UO_1325 (O_1325,N_14648,N_14789);
nand UO_1326 (O_1326,N_14773,N_14580);
nand UO_1327 (O_1327,N_14687,N_14936);
nor UO_1328 (O_1328,N_14550,N_14621);
or UO_1329 (O_1329,N_14552,N_14737);
nor UO_1330 (O_1330,N_14715,N_14954);
and UO_1331 (O_1331,N_14987,N_14900);
nor UO_1332 (O_1332,N_14531,N_14574);
nor UO_1333 (O_1333,N_14967,N_14957);
nor UO_1334 (O_1334,N_14749,N_14911);
xor UO_1335 (O_1335,N_14772,N_14563);
nor UO_1336 (O_1336,N_14988,N_14502);
xnor UO_1337 (O_1337,N_14830,N_14670);
and UO_1338 (O_1338,N_14709,N_14886);
xnor UO_1339 (O_1339,N_14871,N_14826);
nand UO_1340 (O_1340,N_14574,N_14536);
nand UO_1341 (O_1341,N_14993,N_14721);
xor UO_1342 (O_1342,N_14616,N_14717);
nor UO_1343 (O_1343,N_14826,N_14900);
nor UO_1344 (O_1344,N_14577,N_14718);
or UO_1345 (O_1345,N_14661,N_14741);
and UO_1346 (O_1346,N_14643,N_14622);
nand UO_1347 (O_1347,N_14513,N_14999);
nand UO_1348 (O_1348,N_14982,N_14795);
and UO_1349 (O_1349,N_14973,N_14595);
and UO_1350 (O_1350,N_14966,N_14819);
nand UO_1351 (O_1351,N_14706,N_14739);
nor UO_1352 (O_1352,N_14539,N_14970);
xor UO_1353 (O_1353,N_14608,N_14506);
and UO_1354 (O_1354,N_14603,N_14533);
xnor UO_1355 (O_1355,N_14604,N_14849);
nor UO_1356 (O_1356,N_14500,N_14523);
or UO_1357 (O_1357,N_14892,N_14726);
xnor UO_1358 (O_1358,N_14602,N_14993);
nor UO_1359 (O_1359,N_14889,N_14661);
nand UO_1360 (O_1360,N_14525,N_14874);
nand UO_1361 (O_1361,N_14750,N_14578);
xnor UO_1362 (O_1362,N_14706,N_14713);
or UO_1363 (O_1363,N_14539,N_14516);
or UO_1364 (O_1364,N_14846,N_14540);
nor UO_1365 (O_1365,N_14662,N_14826);
or UO_1366 (O_1366,N_14903,N_14807);
or UO_1367 (O_1367,N_14540,N_14567);
nand UO_1368 (O_1368,N_14965,N_14566);
or UO_1369 (O_1369,N_14693,N_14999);
and UO_1370 (O_1370,N_14637,N_14626);
nor UO_1371 (O_1371,N_14726,N_14525);
xor UO_1372 (O_1372,N_14934,N_14587);
nor UO_1373 (O_1373,N_14595,N_14776);
or UO_1374 (O_1374,N_14971,N_14574);
xnor UO_1375 (O_1375,N_14999,N_14753);
nor UO_1376 (O_1376,N_14995,N_14836);
or UO_1377 (O_1377,N_14732,N_14859);
or UO_1378 (O_1378,N_14533,N_14942);
nor UO_1379 (O_1379,N_14774,N_14666);
nand UO_1380 (O_1380,N_14674,N_14888);
nand UO_1381 (O_1381,N_14815,N_14507);
xor UO_1382 (O_1382,N_14887,N_14626);
xor UO_1383 (O_1383,N_14558,N_14598);
and UO_1384 (O_1384,N_14739,N_14796);
nor UO_1385 (O_1385,N_14949,N_14898);
nor UO_1386 (O_1386,N_14640,N_14732);
nand UO_1387 (O_1387,N_14738,N_14619);
and UO_1388 (O_1388,N_14926,N_14620);
nor UO_1389 (O_1389,N_14716,N_14947);
xor UO_1390 (O_1390,N_14842,N_14768);
and UO_1391 (O_1391,N_14842,N_14513);
nand UO_1392 (O_1392,N_14767,N_14559);
nor UO_1393 (O_1393,N_14586,N_14922);
nor UO_1394 (O_1394,N_14943,N_14983);
xor UO_1395 (O_1395,N_14804,N_14904);
and UO_1396 (O_1396,N_14852,N_14965);
nand UO_1397 (O_1397,N_14532,N_14513);
nand UO_1398 (O_1398,N_14756,N_14654);
xor UO_1399 (O_1399,N_14878,N_14646);
or UO_1400 (O_1400,N_14554,N_14866);
nand UO_1401 (O_1401,N_14786,N_14504);
nand UO_1402 (O_1402,N_14567,N_14709);
xor UO_1403 (O_1403,N_14987,N_14507);
and UO_1404 (O_1404,N_14784,N_14504);
and UO_1405 (O_1405,N_14683,N_14677);
xor UO_1406 (O_1406,N_14937,N_14570);
nand UO_1407 (O_1407,N_14617,N_14748);
or UO_1408 (O_1408,N_14748,N_14769);
nand UO_1409 (O_1409,N_14979,N_14783);
nor UO_1410 (O_1410,N_14826,N_14581);
and UO_1411 (O_1411,N_14890,N_14932);
nor UO_1412 (O_1412,N_14997,N_14562);
or UO_1413 (O_1413,N_14812,N_14690);
xor UO_1414 (O_1414,N_14662,N_14757);
xor UO_1415 (O_1415,N_14520,N_14681);
nor UO_1416 (O_1416,N_14886,N_14651);
or UO_1417 (O_1417,N_14623,N_14875);
nor UO_1418 (O_1418,N_14935,N_14816);
nand UO_1419 (O_1419,N_14721,N_14557);
nand UO_1420 (O_1420,N_14532,N_14889);
or UO_1421 (O_1421,N_14931,N_14785);
or UO_1422 (O_1422,N_14742,N_14750);
nand UO_1423 (O_1423,N_14798,N_14775);
nand UO_1424 (O_1424,N_14796,N_14656);
nor UO_1425 (O_1425,N_14767,N_14691);
nor UO_1426 (O_1426,N_14687,N_14921);
nor UO_1427 (O_1427,N_14855,N_14735);
or UO_1428 (O_1428,N_14529,N_14517);
nand UO_1429 (O_1429,N_14610,N_14876);
nor UO_1430 (O_1430,N_14674,N_14580);
and UO_1431 (O_1431,N_14825,N_14833);
or UO_1432 (O_1432,N_14627,N_14806);
and UO_1433 (O_1433,N_14895,N_14891);
or UO_1434 (O_1434,N_14581,N_14875);
and UO_1435 (O_1435,N_14668,N_14700);
xor UO_1436 (O_1436,N_14694,N_14620);
and UO_1437 (O_1437,N_14930,N_14596);
nor UO_1438 (O_1438,N_14876,N_14555);
or UO_1439 (O_1439,N_14806,N_14958);
or UO_1440 (O_1440,N_14526,N_14941);
or UO_1441 (O_1441,N_14830,N_14836);
and UO_1442 (O_1442,N_14815,N_14669);
nor UO_1443 (O_1443,N_14537,N_14844);
nand UO_1444 (O_1444,N_14931,N_14677);
and UO_1445 (O_1445,N_14573,N_14508);
or UO_1446 (O_1446,N_14613,N_14803);
or UO_1447 (O_1447,N_14850,N_14891);
and UO_1448 (O_1448,N_14919,N_14903);
nand UO_1449 (O_1449,N_14654,N_14839);
and UO_1450 (O_1450,N_14763,N_14821);
nand UO_1451 (O_1451,N_14961,N_14640);
nand UO_1452 (O_1452,N_14924,N_14686);
or UO_1453 (O_1453,N_14773,N_14844);
nor UO_1454 (O_1454,N_14857,N_14745);
nand UO_1455 (O_1455,N_14559,N_14738);
or UO_1456 (O_1456,N_14718,N_14895);
nor UO_1457 (O_1457,N_14979,N_14611);
nor UO_1458 (O_1458,N_14541,N_14909);
and UO_1459 (O_1459,N_14630,N_14979);
nand UO_1460 (O_1460,N_14693,N_14921);
or UO_1461 (O_1461,N_14979,N_14730);
nand UO_1462 (O_1462,N_14542,N_14840);
xnor UO_1463 (O_1463,N_14920,N_14553);
nand UO_1464 (O_1464,N_14904,N_14562);
xor UO_1465 (O_1465,N_14738,N_14620);
nor UO_1466 (O_1466,N_14964,N_14776);
xnor UO_1467 (O_1467,N_14758,N_14690);
xor UO_1468 (O_1468,N_14971,N_14610);
and UO_1469 (O_1469,N_14928,N_14853);
nand UO_1470 (O_1470,N_14737,N_14515);
nor UO_1471 (O_1471,N_14805,N_14778);
nand UO_1472 (O_1472,N_14559,N_14656);
nor UO_1473 (O_1473,N_14535,N_14787);
nand UO_1474 (O_1474,N_14763,N_14759);
xor UO_1475 (O_1475,N_14809,N_14696);
nand UO_1476 (O_1476,N_14610,N_14704);
nand UO_1477 (O_1477,N_14836,N_14937);
nor UO_1478 (O_1478,N_14937,N_14723);
xnor UO_1479 (O_1479,N_14913,N_14800);
and UO_1480 (O_1480,N_14511,N_14534);
xor UO_1481 (O_1481,N_14789,N_14630);
and UO_1482 (O_1482,N_14557,N_14517);
nand UO_1483 (O_1483,N_14614,N_14900);
nor UO_1484 (O_1484,N_14501,N_14630);
nor UO_1485 (O_1485,N_14965,N_14712);
and UO_1486 (O_1486,N_14767,N_14625);
nor UO_1487 (O_1487,N_14937,N_14517);
and UO_1488 (O_1488,N_14944,N_14560);
or UO_1489 (O_1489,N_14631,N_14987);
xor UO_1490 (O_1490,N_14666,N_14566);
xnor UO_1491 (O_1491,N_14640,N_14666);
and UO_1492 (O_1492,N_14706,N_14937);
xor UO_1493 (O_1493,N_14600,N_14760);
and UO_1494 (O_1494,N_14563,N_14697);
and UO_1495 (O_1495,N_14899,N_14568);
xnor UO_1496 (O_1496,N_14878,N_14713);
and UO_1497 (O_1497,N_14960,N_14596);
nor UO_1498 (O_1498,N_14544,N_14510);
nand UO_1499 (O_1499,N_14991,N_14795);
xor UO_1500 (O_1500,N_14567,N_14570);
xor UO_1501 (O_1501,N_14522,N_14748);
or UO_1502 (O_1502,N_14562,N_14678);
and UO_1503 (O_1503,N_14566,N_14501);
and UO_1504 (O_1504,N_14727,N_14797);
nor UO_1505 (O_1505,N_14712,N_14519);
xor UO_1506 (O_1506,N_14552,N_14631);
nor UO_1507 (O_1507,N_14973,N_14831);
xor UO_1508 (O_1508,N_14700,N_14703);
nor UO_1509 (O_1509,N_14629,N_14571);
xor UO_1510 (O_1510,N_14576,N_14925);
or UO_1511 (O_1511,N_14823,N_14581);
xor UO_1512 (O_1512,N_14932,N_14584);
or UO_1513 (O_1513,N_14761,N_14856);
xor UO_1514 (O_1514,N_14694,N_14580);
nor UO_1515 (O_1515,N_14643,N_14797);
xnor UO_1516 (O_1516,N_14644,N_14752);
xor UO_1517 (O_1517,N_14811,N_14563);
xnor UO_1518 (O_1518,N_14758,N_14947);
or UO_1519 (O_1519,N_14963,N_14566);
xor UO_1520 (O_1520,N_14752,N_14926);
nand UO_1521 (O_1521,N_14626,N_14761);
and UO_1522 (O_1522,N_14766,N_14532);
and UO_1523 (O_1523,N_14692,N_14800);
xnor UO_1524 (O_1524,N_14798,N_14847);
and UO_1525 (O_1525,N_14835,N_14628);
or UO_1526 (O_1526,N_14796,N_14704);
nor UO_1527 (O_1527,N_14885,N_14790);
nand UO_1528 (O_1528,N_14729,N_14846);
nand UO_1529 (O_1529,N_14632,N_14676);
nor UO_1530 (O_1530,N_14852,N_14961);
and UO_1531 (O_1531,N_14947,N_14739);
nand UO_1532 (O_1532,N_14847,N_14520);
xor UO_1533 (O_1533,N_14758,N_14891);
or UO_1534 (O_1534,N_14709,N_14742);
or UO_1535 (O_1535,N_14936,N_14741);
or UO_1536 (O_1536,N_14670,N_14757);
or UO_1537 (O_1537,N_14815,N_14886);
xor UO_1538 (O_1538,N_14925,N_14915);
xnor UO_1539 (O_1539,N_14664,N_14894);
nor UO_1540 (O_1540,N_14603,N_14895);
nor UO_1541 (O_1541,N_14680,N_14512);
xnor UO_1542 (O_1542,N_14972,N_14650);
or UO_1543 (O_1543,N_14777,N_14876);
and UO_1544 (O_1544,N_14563,N_14572);
nor UO_1545 (O_1545,N_14897,N_14939);
or UO_1546 (O_1546,N_14837,N_14709);
nand UO_1547 (O_1547,N_14833,N_14651);
xor UO_1548 (O_1548,N_14777,N_14898);
xor UO_1549 (O_1549,N_14854,N_14758);
nor UO_1550 (O_1550,N_14911,N_14594);
nand UO_1551 (O_1551,N_14554,N_14614);
nand UO_1552 (O_1552,N_14682,N_14926);
nand UO_1553 (O_1553,N_14530,N_14751);
nand UO_1554 (O_1554,N_14724,N_14973);
nor UO_1555 (O_1555,N_14818,N_14609);
or UO_1556 (O_1556,N_14800,N_14617);
xor UO_1557 (O_1557,N_14769,N_14507);
or UO_1558 (O_1558,N_14525,N_14919);
or UO_1559 (O_1559,N_14789,N_14801);
or UO_1560 (O_1560,N_14704,N_14688);
nor UO_1561 (O_1561,N_14831,N_14658);
or UO_1562 (O_1562,N_14592,N_14813);
or UO_1563 (O_1563,N_14530,N_14528);
and UO_1564 (O_1564,N_14893,N_14800);
nor UO_1565 (O_1565,N_14895,N_14795);
nand UO_1566 (O_1566,N_14840,N_14867);
and UO_1567 (O_1567,N_14752,N_14899);
or UO_1568 (O_1568,N_14892,N_14963);
xnor UO_1569 (O_1569,N_14910,N_14665);
or UO_1570 (O_1570,N_14972,N_14897);
nor UO_1571 (O_1571,N_14962,N_14907);
or UO_1572 (O_1572,N_14977,N_14862);
nor UO_1573 (O_1573,N_14771,N_14629);
and UO_1574 (O_1574,N_14944,N_14707);
and UO_1575 (O_1575,N_14992,N_14654);
nor UO_1576 (O_1576,N_14931,N_14755);
or UO_1577 (O_1577,N_14687,N_14625);
xor UO_1578 (O_1578,N_14695,N_14991);
xnor UO_1579 (O_1579,N_14850,N_14834);
nand UO_1580 (O_1580,N_14769,N_14861);
or UO_1581 (O_1581,N_14694,N_14931);
xor UO_1582 (O_1582,N_14501,N_14833);
and UO_1583 (O_1583,N_14533,N_14768);
and UO_1584 (O_1584,N_14738,N_14721);
nand UO_1585 (O_1585,N_14547,N_14867);
nand UO_1586 (O_1586,N_14671,N_14530);
nand UO_1587 (O_1587,N_14600,N_14960);
or UO_1588 (O_1588,N_14663,N_14892);
or UO_1589 (O_1589,N_14965,N_14907);
or UO_1590 (O_1590,N_14945,N_14534);
nor UO_1591 (O_1591,N_14788,N_14608);
nor UO_1592 (O_1592,N_14969,N_14504);
nand UO_1593 (O_1593,N_14662,N_14783);
nor UO_1594 (O_1594,N_14763,N_14984);
or UO_1595 (O_1595,N_14562,N_14973);
nand UO_1596 (O_1596,N_14928,N_14622);
xor UO_1597 (O_1597,N_14551,N_14793);
or UO_1598 (O_1598,N_14745,N_14794);
or UO_1599 (O_1599,N_14963,N_14528);
and UO_1600 (O_1600,N_14936,N_14696);
or UO_1601 (O_1601,N_14686,N_14797);
xor UO_1602 (O_1602,N_14948,N_14771);
and UO_1603 (O_1603,N_14684,N_14960);
and UO_1604 (O_1604,N_14745,N_14613);
nand UO_1605 (O_1605,N_14545,N_14530);
nand UO_1606 (O_1606,N_14987,N_14793);
nor UO_1607 (O_1607,N_14942,N_14683);
nor UO_1608 (O_1608,N_14552,N_14931);
nor UO_1609 (O_1609,N_14864,N_14579);
nand UO_1610 (O_1610,N_14946,N_14657);
or UO_1611 (O_1611,N_14524,N_14833);
or UO_1612 (O_1612,N_14774,N_14973);
nor UO_1613 (O_1613,N_14593,N_14866);
nand UO_1614 (O_1614,N_14553,N_14981);
or UO_1615 (O_1615,N_14591,N_14578);
nor UO_1616 (O_1616,N_14850,N_14803);
or UO_1617 (O_1617,N_14802,N_14658);
and UO_1618 (O_1618,N_14708,N_14794);
xor UO_1619 (O_1619,N_14686,N_14755);
nand UO_1620 (O_1620,N_14906,N_14619);
or UO_1621 (O_1621,N_14507,N_14729);
nor UO_1622 (O_1622,N_14737,N_14845);
nor UO_1623 (O_1623,N_14996,N_14809);
nand UO_1624 (O_1624,N_14690,N_14527);
and UO_1625 (O_1625,N_14776,N_14972);
and UO_1626 (O_1626,N_14797,N_14614);
nor UO_1627 (O_1627,N_14930,N_14540);
xnor UO_1628 (O_1628,N_14732,N_14912);
or UO_1629 (O_1629,N_14862,N_14651);
xor UO_1630 (O_1630,N_14776,N_14686);
xor UO_1631 (O_1631,N_14544,N_14609);
and UO_1632 (O_1632,N_14727,N_14674);
or UO_1633 (O_1633,N_14946,N_14652);
nand UO_1634 (O_1634,N_14809,N_14901);
nand UO_1635 (O_1635,N_14588,N_14913);
nand UO_1636 (O_1636,N_14945,N_14751);
nand UO_1637 (O_1637,N_14985,N_14924);
nand UO_1638 (O_1638,N_14759,N_14686);
xnor UO_1639 (O_1639,N_14647,N_14728);
nor UO_1640 (O_1640,N_14941,N_14521);
or UO_1641 (O_1641,N_14588,N_14971);
nor UO_1642 (O_1642,N_14986,N_14673);
nor UO_1643 (O_1643,N_14963,N_14921);
nand UO_1644 (O_1644,N_14868,N_14759);
nor UO_1645 (O_1645,N_14724,N_14716);
xor UO_1646 (O_1646,N_14746,N_14892);
or UO_1647 (O_1647,N_14935,N_14798);
xnor UO_1648 (O_1648,N_14654,N_14676);
nor UO_1649 (O_1649,N_14676,N_14769);
nor UO_1650 (O_1650,N_14561,N_14863);
nand UO_1651 (O_1651,N_14954,N_14670);
nor UO_1652 (O_1652,N_14607,N_14908);
or UO_1653 (O_1653,N_14944,N_14552);
nand UO_1654 (O_1654,N_14667,N_14626);
nor UO_1655 (O_1655,N_14776,N_14558);
and UO_1656 (O_1656,N_14919,N_14834);
nor UO_1657 (O_1657,N_14926,N_14883);
or UO_1658 (O_1658,N_14704,N_14999);
nor UO_1659 (O_1659,N_14779,N_14998);
xnor UO_1660 (O_1660,N_14707,N_14555);
or UO_1661 (O_1661,N_14684,N_14926);
xnor UO_1662 (O_1662,N_14657,N_14719);
nor UO_1663 (O_1663,N_14796,N_14759);
or UO_1664 (O_1664,N_14742,N_14981);
nor UO_1665 (O_1665,N_14801,N_14869);
nor UO_1666 (O_1666,N_14865,N_14933);
nor UO_1667 (O_1667,N_14751,N_14574);
nand UO_1668 (O_1668,N_14607,N_14995);
and UO_1669 (O_1669,N_14502,N_14846);
nor UO_1670 (O_1670,N_14835,N_14651);
or UO_1671 (O_1671,N_14731,N_14812);
nand UO_1672 (O_1672,N_14936,N_14997);
nor UO_1673 (O_1673,N_14691,N_14649);
or UO_1674 (O_1674,N_14530,N_14845);
nand UO_1675 (O_1675,N_14786,N_14902);
xor UO_1676 (O_1676,N_14904,N_14868);
and UO_1677 (O_1677,N_14621,N_14910);
nor UO_1678 (O_1678,N_14751,N_14858);
and UO_1679 (O_1679,N_14594,N_14847);
nor UO_1680 (O_1680,N_14992,N_14613);
xnor UO_1681 (O_1681,N_14810,N_14601);
xor UO_1682 (O_1682,N_14860,N_14718);
or UO_1683 (O_1683,N_14645,N_14783);
and UO_1684 (O_1684,N_14917,N_14634);
and UO_1685 (O_1685,N_14555,N_14805);
nand UO_1686 (O_1686,N_14963,N_14622);
nand UO_1687 (O_1687,N_14929,N_14980);
and UO_1688 (O_1688,N_14853,N_14686);
nand UO_1689 (O_1689,N_14767,N_14609);
or UO_1690 (O_1690,N_14974,N_14985);
xor UO_1691 (O_1691,N_14792,N_14982);
or UO_1692 (O_1692,N_14729,N_14828);
and UO_1693 (O_1693,N_14953,N_14736);
nand UO_1694 (O_1694,N_14532,N_14974);
xor UO_1695 (O_1695,N_14898,N_14574);
or UO_1696 (O_1696,N_14541,N_14525);
nor UO_1697 (O_1697,N_14886,N_14688);
xor UO_1698 (O_1698,N_14855,N_14884);
xnor UO_1699 (O_1699,N_14587,N_14814);
or UO_1700 (O_1700,N_14737,N_14811);
and UO_1701 (O_1701,N_14730,N_14822);
xor UO_1702 (O_1702,N_14850,N_14781);
and UO_1703 (O_1703,N_14813,N_14820);
nor UO_1704 (O_1704,N_14937,N_14994);
xor UO_1705 (O_1705,N_14572,N_14679);
or UO_1706 (O_1706,N_14747,N_14877);
nor UO_1707 (O_1707,N_14586,N_14831);
nor UO_1708 (O_1708,N_14790,N_14883);
or UO_1709 (O_1709,N_14671,N_14864);
nor UO_1710 (O_1710,N_14636,N_14601);
nor UO_1711 (O_1711,N_14834,N_14511);
and UO_1712 (O_1712,N_14915,N_14905);
nand UO_1713 (O_1713,N_14989,N_14744);
nor UO_1714 (O_1714,N_14588,N_14953);
nor UO_1715 (O_1715,N_14672,N_14518);
and UO_1716 (O_1716,N_14844,N_14593);
nor UO_1717 (O_1717,N_14917,N_14664);
nor UO_1718 (O_1718,N_14706,N_14659);
nor UO_1719 (O_1719,N_14599,N_14825);
nor UO_1720 (O_1720,N_14701,N_14651);
or UO_1721 (O_1721,N_14933,N_14849);
nand UO_1722 (O_1722,N_14862,N_14896);
nand UO_1723 (O_1723,N_14553,N_14558);
or UO_1724 (O_1724,N_14546,N_14540);
nor UO_1725 (O_1725,N_14564,N_14974);
nor UO_1726 (O_1726,N_14984,N_14965);
nor UO_1727 (O_1727,N_14965,N_14664);
and UO_1728 (O_1728,N_14860,N_14966);
xnor UO_1729 (O_1729,N_14685,N_14520);
xnor UO_1730 (O_1730,N_14886,N_14767);
or UO_1731 (O_1731,N_14629,N_14721);
xnor UO_1732 (O_1732,N_14565,N_14950);
xor UO_1733 (O_1733,N_14579,N_14617);
and UO_1734 (O_1734,N_14556,N_14756);
nand UO_1735 (O_1735,N_14704,N_14733);
and UO_1736 (O_1736,N_14918,N_14831);
nand UO_1737 (O_1737,N_14969,N_14509);
nor UO_1738 (O_1738,N_14997,N_14843);
and UO_1739 (O_1739,N_14883,N_14867);
nor UO_1740 (O_1740,N_14544,N_14514);
or UO_1741 (O_1741,N_14716,N_14578);
nor UO_1742 (O_1742,N_14959,N_14701);
xor UO_1743 (O_1743,N_14999,N_14583);
nand UO_1744 (O_1744,N_14795,N_14704);
xor UO_1745 (O_1745,N_14639,N_14759);
nand UO_1746 (O_1746,N_14509,N_14592);
xor UO_1747 (O_1747,N_14553,N_14561);
nand UO_1748 (O_1748,N_14929,N_14693);
nand UO_1749 (O_1749,N_14946,N_14706);
and UO_1750 (O_1750,N_14864,N_14828);
nand UO_1751 (O_1751,N_14715,N_14904);
nand UO_1752 (O_1752,N_14993,N_14612);
nand UO_1753 (O_1753,N_14617,N_14854);
nor UO_1754 (O_1754,N_14810,N_14978);
nor UO_1755 (O_1755,N_14999,N_14720);
nor UO_1756 (O_1756,N_14876,N_14695);
and UO_1757 (O_1757,N_14863,N_14630);
xnor UO_1758 (O_1758,N_14651,N_14502);
and UO_1759 (O_1759,N_14834,N_14735);
xor UO_1760 (O_1760,N_14580,N_14820);
or UO_1761 (O_1761,N_14698,N_14764);
nor UO_1762 (O_1762,N_14810,N_14514);
nand UO_1763 (O_1763,N_14624,N_14853);
xnor UO_1764 (O_1764,N_14860,N_14786);
nor UO_1765 (O_1765,N_14571,N_14992);
or UO_1766 (O_1766,N_14780,N_14767);
xor UO_1767 (O_1767,N_14575,N_14825);
nor UO_1768 (O_1768,N_14864,N_14901);
xnor UO_1769 (O_1769,N_14925,N_14692);
nor UO_1770 (O_1770,N_14795,N_14662);
xor UO_1771 (O_1771,N_14852,N_14653);
xor UO_1772 (O_1772,N_14929,N_14799);
nor UO_1773 (O_1773,N_14934,N_14763);
nor UO_1774 (O_1774,N_14704,N_14692);
and UO_1775 (O_1775,N_14971,N_14757);
nand UO_1776 (O_1776,N_14935,N_14614);
and UO_1777 (O_1777,N_14942,N_14676);
xnor UO_1778 (O_1778,N_14950,N_14589);
or UO_1779 (O_1779,N_14618,N_14901);
or UO_1780 (O_1780,N_14697,N_14959);
and UO_1781 (O_1781,N_14720,N_14777);
xor UO_1782 (O_1782,N_14866,N_14937);
nand UO_1783 (O_1783,N_14885,N_14925);
xnor UO_1784 (O_1784,N_14591,N_14636);
nand UO_1785 (O_1785,N_14886,N_14797);
nor UO_1786 (O_1786,N_14750,N_14870);
nor UO_1787 (O_1787,N_14958,N_14957);
and UO_1788 (O_1788,N_14733,N_14971);
nor UO_1789 (O_1789,N_14634,N_14861);
nor UO_1790 (O_1790,N_14913,N_14783);
nor UO_1791 (O_1791,N_14593,N_14835);
nor UO_1792 (O_1792,N_14555,N_14647);
nor UO_1793 (O_1793,N_14543,N_14625);
and UO_1794 (O_1794,N_14540,N_14574);
and UO_1795 (O_1795,N_14813,N_14509);
nor UO_1796 (O_1796,N_14509,N_14943);
nand UO_1797 (O_1797,N_14865,N_14893);
nand UO_1798 (O_1798,N_14553,N_14605);
and UO_1799 (O_1799,N_14943,N_14774);
nor UO_1800 (O_1800,N_14857,N_14847);
xnor UO_1801 (O_1801,N_14672,N_14624);
nor UO_1802 (O_1802,N_14948,N_14556);
nor UO_1803 (O_1803,N_14846,N_14637);
or UO_1804 (O_1804,N_14825,N_14838);
nand UO_1805 (O_1805,N_14731,N_14935);
or UO_1806 (O_1806,N_14530,N_14889);
and UO_1807 (O_1807,N_14969,N_14679);
nor UO_1808 (O_1808,N_14503,N_14645);
or UO_1809 (O_1809,N_14928,N_14552);
or UO_1810 (O_1810,N_14620,N_14658);
nor UO_1811 (O_1811,N_14678,N_14502);
nor UO_1812 (O_1812,N_14602,N_14532);
nor UO_1813 (O_1813,N_14644,N_14791);
or UO_1814 (O_1814,N_14705,N_14550);
nor UO_1815 (O_1815,N_14985,N_14865);
xor UO_1816 (O_1816,N_14749,N_14877);
xor UO_1817 (O_1817,N_14636,N_14794);
nor UO_1818 (O_1818,N_14970,N_14858);
and UO_1819 (O_1819,N_14946,N_14741);
and UO_1820 (O_1820,N_14633,N_14668);
and UO_1821 (O_1821,N_14975,N_14505);
xor UO_1822 (O_1822,N_14845,N_14529);
xor UO_1823 (O_1823,N_14534,N_14734);
nand UO_1824 (O_1824,N_14891,N_14683);
and UO_1825 (O_1825,N_14622,N_14662);
nor UO_1826 (O_1826,N_14671,N_14578);
and UO_1827 (O_1827,N_14625,N_14511);
and UO_1828 (O_1828,N_14507,N_14814);
nand UO_1829 (O_1829,N_14594,N_14824);
nand UO_1830 (O_1830,N_14789,N_14924);
or UO_1831 (O_1831,N_14738,N_14661);
or UO_1832 (O_1832,N_14915,N_14991);
or UO_1833 (O_1833,N_14588,N_14851);
nand UO_1834 (O_1834,N_14935,N_14748);
nand UO_1835 (O_1835,N_14719,N_14883);
nor UO_1836 (O_1836,N_14829,N_14788);
xnor UO_1837 (O_1837,N_14769,N_14900);
nand UO_1838 (O_1838,N_14504,N_14678);
nand UO_1839 (O_1839,N_14865,N_14983);
nand UO_1840 (O_1840,N_14881,N_14907);
and UO_1841 (O_1841,N_14555,N_14913);
and UO_1842 (O_1842,N_14633,N_14627);
nand UO_1843 (O_1843,N_14831,N_14505);
and UO_1844 (O_1844,N_14699,N_14860);
nor UO_1845 (O_1845,N_14808,N_14558);
or UO_1846 (O_1846,N_14968,N_14674);
nor UO_1847 (O_1847,N_14771,N_14638);
nor UO_1848 (O_1848,N_14647,N_14716);
nand UO_1849 (O_1849,N_14797,N_14684);
xnor UO_1850 (O_1850,N_14926,N_14776);
or UO_1851 (O_1851,N_14515,N_14508);
nand UO_1852 (O_1852,N_14810,N_14692);
and UO_1853 (O_1853,N_14941,N_14678);
and UO_1854 (O_1854,N_14946,N_14839);
xor UO_1855 (O_1855,N_14538,N_14703);
or UO_1856 (O_1856,N_14712,N_14906);
nor UO_1857 (O_1857,N_14760,N_14522);
xor UO_1858 (O_1858,N_14723,N_14787);
nor UO_1859 (O_1859,N_14946,N_14717);
nand UO_1860 (O_1860,N_14736,N_14639);
xnor UO_1861 (O_1861,N_14595,N_14625);
nor UO_1862 (O_1862,N_14801,N_14850);
nand UO_1863 (O_1863,N_14524,N_14632);
nor UO_1864 (O_1864,N_14952,N_14965);
xor UO_1865 (O_1865,N_14587,N_14713);
or UO_1866 (O_1866,N_14784,N_14765);
xor UO_1867 (O_1867,N_14956,N_14939);
nor UO_1868 (O_1868,N_14882,N_14984);
nor UO_1869 (O_1869,N_14894,N_14852);
xor UO_1870 (O_1870,N_14710,N_14541);
and UO_1871 (O_1871,N_14888,N_14904);
nand UO_1872 (O_1872,N_14807,N_14720);
nor UO_1873 (O_1873,N_14814,N_14615);
nor UO_1874 (O_1874,N_14859,N_14976);
and UO_1875 (O_1875,N_14523,N_14898);
nand UO_1876 (O_1876,N_14944,N_14566);
xor UO_1877 (O_1877,N_14643,N_14748);
nand UO_1878 (O_1878,N_14848,N_14708);
xor UO_1879 (O_1879,N_14812,N_14593);
nor UO_1880 (O_1880,N_14795,N_14993);
nor UO_1881 (O_1881,N_14519,N_14828);
nand UO_1882 (O_1882,N_14522,N_14971);
nor UO_1883 (O_1883,N_14788,N_14843);
nor UO_1884 (O_1884,N_14884,N_14506);
and UO_1885 (O_1885,N_14557,N_14995);
nor UO_1886 (O_1886,N_14510,N_14640);
nand UO_1887 (O_1887,N_14676,N_14607);
and UO_1888 (O_1888,N_14838,N_14852);
or UO_1889 (O_1889,N_14860,N_14576);
nand UO_1890 (O_1890,N_14964,N_14532);
nand UO_1891 (O_1891,N_14609,N_14940);
or UO_1892 (O_1892,N_14798,N_14980);
nand UO_1893 (O_1893,N_14554,N_14706);
and UO_1894 (O_1894,N_14929,N_14835);
or UO_1895 (O_1895,N_14607,N_14673);
xnor UO_1896 (O_1896,N_14521,N_14752);
and UO_1897 (O_1897,N_14710,N_14728);
nand UO_1898 (O_1898,N_14992,N_14762);
nand UO_1899 (O_1899,N_14986,N_14771);
xor UO_1900 (O_1900,N_14783,N_14634);
nor UO_1901 (O_1901,N_14716,N_14885);
nor UO_1902 (O_1902,N_14595,N_14636);
nand UO_1903 (O_1903,N_14617,N_14742);
nand UO_1904 (O_1904,N_14551,N_14716);
and UO_1905 (O_1905,N_14670,N_14924);
or UO_1906 (O_1906,N_14753,N_14907);
nand UO_1907 (O_1907,N_14907,N_14872);
xnor UO_1908 (O_1908,N_14876,N_14680);
nand UO_1909 (O_1909,N_14728,N_14904);
xnor UO_1910 (O_1910,N_14644,N_14593);
or UO_1911 (O_1911,N_14704,N_14824);
or UO_1912 (O_1912,N_14667,N_14899);
and UO_1913 (O_1913,N_14662,N_14556);
nor UO_1914 (O_1914,N_14798,N_14559);
nor UO_1915 (O_1915,N_14818,N_14503);
nor UO_1916 (O_1916,N_14519,N_14692);
nor UO_1917 (O_1917,N_14644,N_14806);
and UO_1918 (O_1918,N_14752,N_14910);
and UO_1919 (O_1919,N_14703,N_14966);
nand UO_1920 (O_1920,N_14747,N_14853);
or UO_1921 (O_1921,N_14999,N_14812);
xnor UO_1922 (O_1922,N_14804,N_14566);
nand UO_1923 (O_1923,N_14609,N_14804);
nand UO_1924 (O_1924,N_14764,N_14797);
or UO_1925 (O_1925,N_14523,N_14847);
nor UO_1926 (O_1926,N_14984,N_14616);
xnor UO_1927 (O_1927,N_14983,N_14600);
or UO_1928 (O_1928,N_14587,N_14563);
xor UO_1929 (O_1929,N_14657,N_14565);
or UO_1930 (O_1930,N_14762,N_14823);
nor UO_1931 (O_1931,N_14702,N_14764);
xnor UO_1932 (O_1932,N_14592,N_14726);
or UO_1933 (O_1933,N_14553,N_14551);
xnor UO_1934 (O_1934,N_14714,N_14729);
or UO_1935 (O_1935,N_14775,N_14501);
nor UO_1936 (O_1936,N_14948,N_14567);
nor UO_1937 (O_1937,N_14955,N_14992);
or UO_1938 (O_1938,N_14962,N_14567);
nand UO_1939 (O_1939,N_14963,N_14839);
nor UO_1940 (O_1940,N_14849,N_14822);
nor UO_1941 (O_1941,N_14635,N_14562);
nor UO_1942 (O_1942,N_14941,N_14945);
nor UO_1943 (O_1943,N_14687,N_14942);
nor UO_1944 (O_1944,N_14639,N_14566);
nor UO_1945 (O_1945,N_14512,N_14614);
and UO_1946 (O_1946,N_14929,N_14811);
and UO_1947 (O_1947,N_14835,N_14904);
nor UO_1948 (O_1948,N_14823,N_14788);
and UO_1949 (O_1949,N_14947,N_14515);
xor UO_1950 (O_1950,N_14542,N_14605);
and UO_1951 (O_1951,N_14972,N_14959);
xor UO_1952 (O_1952,N_14722,N_14556);
nand UO_1953 (O_1953,N_14564,N_14764);
xor UO_1954 (O_1954,N_14716,N_14958);
and UO_1955 (O_1955,N_14748,N_14535);
or UO_1956 (O_1956,N_14587,N_14809);
and UO_1957 (O_1957,N_14719,N_14895);
xor UO_1958 (O_1958,N_14559,N_14683);
xor UO_1959 (O_1959,N_14657,N_14729);
nor UO_1960 (O_1960,N_14916,N_14651);
and UO_1961 (O_1961,N_14642,N_14839);
nand UO_1962 (O_1962,N_14718,N_14688);
xnor UO_1963 (O_1963,N_14763,N_14583);
xor UO_1964 (O_1964,N_14987,N_14625);
nand UO_1965 (O_1965,N_14707,N_14860);
xor UO_1966 (O_1966,N_14705,N_14708);
nor UO_1967 (O_1967,N_14802,N_14986);
nor UO_1968 (O_1968,N_14546,N_14953);
xor UO_1969 (O_1969,N_14897,N_14818);
nand UO_1970 (O_1970,N_14632,N_14618);
or UO_1971 (O_1971,N_14781,N_14807);
nand UO_1972 (O_1972,N_14854,N_14905);
or UO_1973 (O_1973,N_14984,N_14666);
nand UO_1974 (O_1974,N_14975,N_14872);
xor UO_1975 (O_1975,N_14890,N_14918);
and UO_1976 (O_1976,N_14632,N_14564);
nor UO_1977 (O_1977,N_14768,N_14560);
xnor UO_1978 (O_1978,N_14996,N_14819);
or UO_1979 (O_1979,N_14790,N_14686);
nor UO_1980 (O_1980,N_14746,N_14941);
or UO_1981 (O_1981,N_14852,N_14772);
nor UO_1982 (O_1982,N_14883,N_14529);
and UO_1983 (O_1983,N_14657,N_14798);
xor UO_1984 (O_1984,N_14894,N_14847);
or UO_1985 (O_1985,N_14540,N_14537);
nor UO_1986 (O_1986,N_14604,N_14858);
xor UO_1987 (O_1987,N_14635,N_14639);
xnor UO_1988 (O_1988,N_14767,N_14615);
nor UO_1989 (O_1989,N_14975,N_14628);
nand UO_1990 (O_1990,N_14821,N_14906);
and UO_1991 (O_1991,N_14947,N_14599);
xor UO_1992 (O_1992,N_14767,N_14553);
or UO_1993 (O_1993,N_14891,N_14617);
nand UO_1994 (O_1994,N_14991,N_14919);
or UO_1995 (O_1995,N_14825,N_14987);
nand UO_1996 (O_1996,N_14864,N_14988);
nor UO_1997 (O_1997,N_14505,N_14925);
nor UO_1998 (O_1998,N_14947,N_14679);
and UO_1999 (O_1999,N_14987,N_14795);
endmodule